PK
     mdZ �b=�' �'    cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0":["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_0","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_0","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_0"],"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1":["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_1","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_1","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_1"],"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2":["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"],"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3":["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_0":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_1":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_3":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_4":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_6":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_7":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_8":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_9":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_10":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_11":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_12":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_13":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_14":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_15":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_16":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_17":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_18":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_20":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_21":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_22":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_23":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_25":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28":["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_3"],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29":["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_3"],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_30":["pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_3"],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_31":["pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_2"],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32":["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_2","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_2"],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_33":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_34":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_35":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_36":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_37":[],"pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_0":[],"pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1":["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_6","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_6"],"pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2":["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3"],"pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_0":[],"pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1":["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_6","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_8"],"pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2":["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3"],"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0":["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"],"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1":["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"],"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0":["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0"],"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1":["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1"],"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2":["pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_4"],"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3":["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_5","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2"],"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0":["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0"],"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1":["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1"],"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2":["pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_5"],"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3":["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_5","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2"],"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_0":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"],"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_1":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"],"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_2":["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32"],"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_3":["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28"],"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4":["pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_9"],"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_5":["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3"],"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_6":["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1"],"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_0":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"],"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_1":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"],"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_2":["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32"],"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_3":["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29"],"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4":["pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_7"],"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_5":["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3"],"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_6":["pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1"],"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0":["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0"],"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1":["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1"],"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"],"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"],"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_0":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"],"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_1":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"],"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_2":["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_31"],"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_3":["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_30"],"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_4":["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2"],"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_5":["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2"],"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_6":["pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1"],"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_7":["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4"],"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_8":["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1"],"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_9":["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4"]},"pin_to_color":{"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0":"#005F39","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1":"#9E008E","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2":"#FF6E41","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3":"#00FFC6","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_0":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_1":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_3":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_4":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_6":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_7":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_8":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_9":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_10":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_11":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_12":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_13":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_14":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_15":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_16":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_17":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_18":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19":"#005F39","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_20":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_21":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_22":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_23":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24":"#9E008E","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_25":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28":"#001544","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29":"#91D0CB","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_30":"#FF029D","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_31":"#5FAD4E","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32":"#007DB5","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_33":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_34":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_35":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_36":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_37":"#000000","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_0":"#000000","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1":"#FFE502","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2":"#E85EBE","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_0":"#000000","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1":"#005F39","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2":"#010067","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0":"#0076FF","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1":"#85A900","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0":"#0076FF","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1":"#85A900","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2":"#683D3B","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3":"#E85EBE","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0":"#0076FF","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1":"#85A900","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2":"#98FF52","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3":"#010067","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_0":"#005F39","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_1":"#9E008E","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_2":"#007DB5","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_3":"#001544","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4":"#968AE8","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_5":"#010067","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_6":"#005F39","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_0":"#005F39","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_1":"#9E008E","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_2":"#007DB5","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_3":"#91D0CB","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4":"#FF74A3","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_5":"#E85EBE","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_6":"#FFE502","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0":"#0076FF","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1":"#85A900","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2":"#00FFC6","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3":"#FF6E41","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_0":"#005F39","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_1":"#9E008E","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_2":"#5FAD4E","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_3":"#FF029D","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_4":"#683D3B","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_5":"#98FF52","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_6":"#FFE502","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_7":"#FF74A3","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_8":"#005F39","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_9":"#968AE8"},"pin_to_state":{"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0":"neutral","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1":"neutral","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2":"neutral","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_0":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_1":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_3":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_4":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_6":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_7":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_8":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_9":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_10":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_11":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_12":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_13":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_14":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_15":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_16":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_17":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_18":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_20":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_21":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_22":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_23":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_25":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_30":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_31":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_33":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_34":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_35":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_36":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_37":"neutral","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_0":"neutral","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1":"neutral","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2":"neutral","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_0":"neutral","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1":"neutral","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2":"neutral","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0":"neutral","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1":"neutral","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0":"neutral","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1":"neutral","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2":"neutral","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3":"neutral","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0":"neutral","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1":"neutral","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2":"neutral","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3":"neutral","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_0":"neutral","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_1":"neutral","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_2":"neutral","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_3":"neutral","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4":"neutral","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_5":"neutral","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_6":"neutral","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_0":"neutral","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_1":"neutral","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_2":"neutral","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_3":"neutral","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4":"neutral","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_5":"neutral","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_6":"neutral","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0":"neutral","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1":"neutral","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2":"neutral","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3":"neutral","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_0":"neutral","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_1":"neutral","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_2":"neutral","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_3":"neutral","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_4":"neutral","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_5":"neutral","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_6":"neutral","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_7":"neutral","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_8":"neutral","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_9":"neutral"},"next_color_idx":20,"wires_placed_in_order":[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_29"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_28"],["pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_28","pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_1"],["pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_0","pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_15"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_29"],["pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_3"],["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_13"],["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_14"],["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_15"],["pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_36"],["pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5"],["pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_0"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_1"],["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_2","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_1"],["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_0","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_0"],["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_1","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_2"],["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_2","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_1"],["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_1","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_2"],["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_0","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_0"],["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_2","pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_1"],["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_1","pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_2"],["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_0","pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_0"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_4"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_4"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_4"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_5"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_5"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_5"],["pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_12"],["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_8"],["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_9"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_0"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_1"],["pin-type-component_a8221eb9-381c-43f6-a63c-1fa17c525231_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"],["pin-type-component_a8221eb9-381c-43f6-a63c-1fa17c525231_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"],["pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_23"],["pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_25"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_0"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_1"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_11"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_10"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_0"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_0"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_1"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_1"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1"],["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"],["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_0"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_3"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_3"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_0"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26"],["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_2"],["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27"],["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_1"],["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"],["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6"],["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_10","pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_0"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_9","pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_1"],["pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_0","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2"],["pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_1","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1"],["pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_0","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2"],["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"],["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"],["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"],["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2"],["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_0"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_1"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"],["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6"],["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4"],["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_5","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3"],["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_5"],["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4"],["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4"],["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2"],["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2"],["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_6","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1"],["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_6","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_7","pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_1"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_8","pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_0"],["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28"],["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29"],["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32"],["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_2"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_1"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_1"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_0"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_0"],["pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_0","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_5"],["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_7","pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_1"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_5","pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_0"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_7","pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_1"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"],["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"],["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"],["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"],["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"],["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"],["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"],["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"],["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_0"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_1"],["pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_31"],["pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_30"],["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_4"],["pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_6"],["pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_7","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4"],["pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_9","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4"],["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_5"],["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_8"]],"wires_removed_and_placed_in_order":[[[],[]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_29"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_28"]]],[[],[["pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_28","pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_1"]]],[[],[["pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_0","pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_15"]]],[[["pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_29","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_29"]]],[[],[]],[[["pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_15","pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_0"]],[]],[[["pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_28","pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_1"],["pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_28","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[["pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]]],[[["pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_29","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_3"]]],[[],[["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_13"]]],[[],[["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_14"]]],[[],[["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_15"]]],[[],[["pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_36"]]],[[],[["pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5"]]],[[],[["pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_0"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_1"]]],[[],[["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_2","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_1"]]],[[],[["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_0","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_0"]]],[[],[["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_1","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_2"]]],[[],[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_2","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_1"]]],[[],[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_1","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_2"]]],[[],[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_0","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_0"]]],[[],[["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_2","pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_1"]]],[[],[["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_1","pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_2"]]],[[],[["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_0","pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_0"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_4"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_4"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_4"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_5"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_5"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_5"]]],[[],[["pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_12"]]],[[],[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_8"]]],[[],[["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_9"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_0"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_1"]]],[[],[["pin-type-component_a8221eb9-381c-43f6-a63c-1fa17c525231_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]]],[[],[["pin-type-component_a8221eb9-381c-43f6-a63c-1fa17c525231_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]]],[[["pin-type-component_a8221eb9-381c-43f6-a63c-1fa17c525231_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]],[]],[[["pin-type-component_a8221eb9-381c-43f6-a63c-1fa17c525231_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]],[]],[[],[["pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_23"]]],[[],[["pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_25"]]],[[["pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_36"]],[]],[[["pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[["pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2"]],[]],[[["pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5"]],[]],[[["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_13"]],[]],[[["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_14"]],[]],[[["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_15"]],[]],[[["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_0","pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_0"]],[]],[[["pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_1","pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_2"]],[]],[[["pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_2","pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_1"]],[]],[[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_0","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_0"]],[]],[[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_2","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_1"]],[]],[[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_1","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_2"]],[]],[[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_8"]],[]],[[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_4","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_5","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_9"]],[]],[[["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_4","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_5","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_0","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_0"]],[]],[[["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_1","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_2"]],[]],[[["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_2","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_1"]],[]],[[["pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_12"]],[]],[[["pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_4","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[["pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_5","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[["pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_23"]],[]],[[["pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_25"]],[]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_0"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_1"]]],[[],[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_11"]]],[[],[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_10"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_0"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_0"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_1"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_1"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1"]]],[[],[["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]]],[[],[["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_0"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_3"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_3"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_0"]]],[[],[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26"]]],[[],[["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_2"]]],[[],[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27"]]],[[],[["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_1"]]],[[],[["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"]]],[[],[["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6"]]],[[],[["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"]]],[[],[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_10","pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_0"]]],[[],[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_9","pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_1"]]],[[],[["pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_0","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2"]]],[[],[["pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_1","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1"]]],[[],[["pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_0","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2"]]],[[["pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1","pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_1"]],[]],[[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1"]],[]],[[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6","pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0"],["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"],["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]],[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"],["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]]],[[["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"],["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]],[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]]],[[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_0"],["pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2","pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_0"]],[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2"]]],[[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_1"]],[]],[[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_0"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_0"]],[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0"]]],[[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_1"]],[]],[[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0"]],[]],[[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6"]],[]],[[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]],[]],[[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]],[]],[[],[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"]]],[[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"]],[]],[[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"]],[]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0"]]],[[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3"]],[]],[[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2"]],[]],[[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0"]],[]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_0"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_1"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"]]],[[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]],[]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"]]],[[],[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6"]]],[[],[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4"]]],[[],[["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_5","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3"]]],[[],[["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_5"]]],[[],[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4"]]],[[],[["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4"]]],[[],[["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2"]]],[[],[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2"]]],[[],[["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_6","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1"]]],[[],[["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_6","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1"]]],[[],[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_7","pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_1"]]],[[],[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_8","pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_0"]]],[[],[["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28"]]],[[],[["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29"]]],[[],[["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32"]]],[[],[["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_2"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_1"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_1"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_0"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_0"]]],[[],[["pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_0","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_5"]]],[[],[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_7","pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_1"]]],[[],[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_5","pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_0"]]],[[],[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_7","pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_1"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"]]],[[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_0","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"]],[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"]]],[[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_1","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"]],[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"]]],[[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]],[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"],["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]]],[[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]],[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"],["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]]],[[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]],[]],[[],[["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]]],[[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]],[]],[[],[["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]]],[[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"]],[]],[[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"]],[]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"]]],[[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27"]],[]],[[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26"]],[]],[[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"]],[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"]]],[[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_5","pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_0"]],[]],[[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"]],[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"]]],[[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_7","pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_1"]],[]],[[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27"]],[]],[[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26"]],[]],[[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"]],[]],[[["pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_0","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_5"]],[]],[[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"]],[]],[[["pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_1","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_7"]],[]],[[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_10"]],[]],[[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_11"]],[]],[[["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5"]],[]],[[["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6"]],[]],[[["pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_1","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_7"]],[]],[[["pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_0","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_8"]],[]],[[["pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_1","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_9"]],[]],[[["pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_0","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_10"]],[]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_0"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_1"]]],[[],[["pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_31"]]],[[],[["pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_30"]]],[[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4"]],[]],[[],[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_4"]]],[[],[["pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_6"]]],[[],[["pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_7","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4"]]],[[["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4"]],[]],[[],[["pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_9","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4"]]],[[],[["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_5"]]],[[],[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_8"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0":"0000000000000000","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1":"0000000000000001","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2":"0000000000000011","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3":"0000000000000010","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_0":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_1":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_3":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_4":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_6":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_7":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_8":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_9":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_10":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_11":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_12":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_13":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_14":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_15":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_16":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_17":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_18":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19":"0000000000000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_20":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_21":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_22":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_23":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24":"0000000000000001","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_25":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28":"0000000000000020","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29":"0000000000000021","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_30":"0000000000000003","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_31":"0000000000000002","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32":"0000000000000022","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_33":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_34":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_35":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_36":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_37":"_","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_0":"_","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1":"0000000000000016","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2":"0000000000000012","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_0":"_","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1":"0000000000000017","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2":"0000000000000013","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0":"0000000000000004","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1":"0000000000000005","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0":"0000000000000004","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1":"0000000000000005","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2":"0000000000000006","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3":"0000000000000012","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0":"0000000000000004","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1":"0000000000000005","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2":"0000000000000009","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3":"0000000000000013","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_0":"0000000000000000","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_1":"0000000000000001","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_2":"0000000000000022","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_3":"0000000000000020","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4":"0000000000000008","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_5":"0000000000000013","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_6":"0000000000000017","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_0":"0000000000000000","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_1":"0000000000000001","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_2":"0000000000000022","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_3":"0000000000000021","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4":"0000000000000007","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_5":"0000000000000012","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_6":"0000000000000016","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0":"0000000000000004","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1":"0000000000000005","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2":"0000000000000010","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3":"0000000000000011","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_0":"0000000000000000","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_1":"0000000000000001","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_2":"0000000000000002","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_3":"0000000000000003","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_4":"0000000000000006","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_5":"0000000000000009","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_6":"0000000000000016","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_7":"0000000000000007","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_8":"0000000000000017","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_9":"0000000000000008"},"component_id_to_pins":{"d53bc8d1-adbf-42c3-9bdc-27d4d2b68588":["0","1","2","3"],"f7d25e04-bb51-41df-ba72-c452c270d3fb":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31","32","33","34","35","36","37"],"32608709-bcb5-4c22-82f1-0b5ac1739be0":[],"915b317b-63a4-4c37-8362-9a35870cbe7c":[],"9e0cc72b-cce0-4555-8c60-9928baea3faa":[],"41689d80-6f1a-478b-ad5a-826ce578b4af":[],"ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8":["0","1","2"],"00e3d6c2-f801-4d91-ad4d-237bada773bb":["0","1","2"],"1c19cc90-e27a-4c31-a566-dce6d12cc7bd":["0","1"],"8b4859a0-119b-4d24-8c3e-f008f1af2f35":[],"eb1dbc1c-94ee-4954-b264-2ba5f2bb6c04":[],"060f78c2-f7c5-4b91-a54e-26722a6a6eb1":["0","1","2","3"],"c483e859-dbe3-40ab-ad85-fdb0e9726a1e":["0","1","2","3"],"d7e83964-79f2-4e6f-ab07-dee67fd9dff8":["0","1","2","3","4","5","6"],"6bde5401-8877-4618-b129-167654a129ea":["0","1","2","3","4","5","6"],"786922c4-3cc4-4e2e-a1af-6f582a726cc5":[],"c6b89f01-cd33-4f53-a410-bd8ce0a19726":[],"028c5ed6-a9ce-4916-bd5a-20a0af91ff53":[],"d8ee4efe-302f-41eb-a87d-4235620299ce":[],"8c415f8f-024b-42a7-9906-fa5d9103b190":[],"f0886e27-8ec0-43da-a659-1cbab4912d9c":[],"9b271475-bebe-41b8-aded-20e21ef4734b":["0","1","2","3"],"fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351":["0","1","2","3","4","5","6","7","8","9"],"60b47335-97ed-4e17-861d-700ea31fb823":[],"1d273ddc-00fe-4e0d-abfe-19b515681189":[],"ff8b35db-2369-4252-b747-2b8feb913443":[],"5830f988-bcfc-482c-9025-2453ea0e5d91":[],"27a36091-2d09-4701-aaa6-228dbe3a2a98":[],"14cfe2b5-1a7f-43d4-89f6-507c0f51956e":[],"f69e8dbc-a536-4df8-89be-06aad4cf7eb6":[]},"uid_to_net":{"_":[],"0000000000000001":["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_1"],"0000000000000000":["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_0"],"0000000000000004":["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"],"0000000000000005":["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"],"0000000000000010":["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"],"0000000000000011":["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"],"0000000000000012":["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_5","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2"],"0000000000000013":["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_5","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2"],"0000000000000016":["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_6","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_6"],"0000000000000017":["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_6","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_8"],"0000000000000020":["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28"],"0000000000000021":["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29"],"0000000000000022":["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_2"],"0000000000000002":["pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_31"],"0000000000000003":["pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_30"],"0000000000000006":["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_4"],"0000000000000007":["pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_7","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4"],"0000000000000008":["pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_9","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4"],"0000000000000009":["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_5"]},"uid_to_text_label":{"0000000000000001":"Net 1","0000000000000000":"Net 0","0000000000000004":"Net 4","0000000000000005":"Net 5","0000000000000010":"Net 10","0000000000000011":"Net 11","0000000000000012":"Net 12","0000000000000013":"Net 13","0000000000000016":"Net 16","0000000000000017":"Net 17","0000000000000020":"Net 20","0000000000000021":"Net 21","0000000000000022":"Net 22","0000000000000002":"Net 2","0000000000000003":"Net 3","0000000000000006":"Net 6","0000000000000007":"Net 7","0000000000000008":"Net 8","0000000000000009":"Net 9"},"all_breadboard_info_list":[],"breadboard_info_list":[],"componentsData":[{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"GND","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[3499.592122094968,381.2251000087314],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"32608709-bcb5-4c22-82f1-0b5ac1739be0","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"VCC +5V","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[3366.1168313046355,378.8059167969202],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"915b317b-63a4-4c37-8362-9a35870cbe7c","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[816.5526985000006,-114.18805750000007],"typeId":"b975acdd-73e3-4b18-a5a5-9b66f369afa0","componentVersion":2,"instanceId":"f7d25e04-bb51-41df-ba72-c452c270d3fb","orientation":"up","circleData":[[947.5,-340.00000000000006],[948.1030000000001,-312.73920549999985],[948.1231135000003,-286.7030244999998],[947.5,-258.2146149999999],[948.7261135000003,-232.17843399999987],[947.5,-206.1221394999999],[948.7261135000003,-178.25684499999983],[948.7261135000003,-152.22066399999994],[948.7261135000003,-124.95986949999983],[948.1030000000001,-99.55068849999985],[949.3291135000004,-71.68539399999995],[949.3291135000004,-44.42309949999995],[949.3291135000004,-16.561691499999938],[949.9306135000002,9.472989500000153],[949.3291135000004,35.48905700000002],[950.5552270000003,64.60058],[949.9306135000002,90.63676099999971],[949.9306135000002,118.52216899999956],[951.7813405000002,146.98896349999978],[678.5382805000002,148.19346349999984],[677.312167,120.32966899999968],[678.5382805000002,94.29348799999975],[677.9352805000001,66.42969349999983],[677.9352805000001,39.16739899999983],[679.1613940000002,12.528216500000212],[678.5382805000002,-14.131078000000002],[679.1613940000002,-43.24259950000001],[677.9352805000001,-70.48328049999995],[677.9352805000001,-95.9164614999999],[677.3322805000003,-121.95264249999988],[677.3322805000003,-149.81793699999986],[677.312167,-176.45323149999984],[678.5583940000001,-203.71402599999982],[677.3322805000003,-229.73009349999984],[675.4824745000001,-258.842026],[677.3322805000003,-284.294911],[677.9349745000002,-310.9130259999999],[677.3322805000003,-338.77388650000006]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"LOAD 1 AC Circuit\n(behind a breaker)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[2521.1223679499117,1492.667604045154],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"9e0cc72b-cce0-4555-8c60-9928baea3faa","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"LOAD 2 AC Circuit\n(behind a breaker)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[2767.5835720784066,1691.9991453659359],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"41689d80-6f1a-478b-ad5a-826ce578b4af","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1576.6917940000021,2672.799167000001],"typeId":"fa95e5d1-b92a-410f-a873-a71d0089e7ad","componentVersion":1,"instanceId":"ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8","orientation":"left","circleData":[[3782.5,-850],[1592.5000000000014,2405.000000000001],[1622.5000000000014,2405.000000000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1126.6917939999953,2687.799166999998],"typeId":"fa95e5d1-b92a-410f-a873-a71d0089e7ad","componentVersion":1,"instanceId":"00e3d6c2-f801-4d91-ad4d-237bada773bb","orientation":"left","circleData":[[3332.5,-835],[1142.499999999994,2419.999999999997],[1172.4999999999932,2419.999999999997]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[3123.2036904999995,1157.474882],"typeId":"5ac8a9e5-bb24-45ef-9b03-1161364522fb","componentVersion":1,"instanceId":"1c19cc90-e27a-4c31-a566-dce6d12cc7bd","orientation":"up","circleData":[[2987.5,1145],[3259.5265,1145]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Main line\n(phase) - L\n(Enedis in France)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[3292.519774875356,1084.5794073453549],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"8b4859a0-119b-4d24-8c3e-f008f1af2f35","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Main neutral - N\n(Enedis in France)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[2953.4352836968415,1091.5820712351226],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"eb1dbc1c-94ee-4954-b264-2ba5f2bb6c04","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[2528.8436755,1583.142836],"typeId":"a64016c8-4d9c-491e-ba46-f626b2aeb38c","componentVersion":1,"instanceId":"060f78c2-f7c5-4b91-a54e-26722a6a6eb1","orientation":"up","circleData":[[2507.5,1430],[2544.3571255,1429.1428745],[2545.6428145,1755.2857490000001],[2509.6428145,1753.1428744999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[2768.8436755000002,1778.142836],"typeId":"a64016c8-4d9c-491e-ba46-f626b2aeb38c","componentVersion":1,"instanceId":"c483e859-dbe3-40ab-ad85-fdb0e9726a1e","orientation":"up","circleData":[[2747.5,1625],[2784.3571255000006,1624.1428745],[2785.6428145,1950.2857490000008],[2749.6428145,1948.1428745000005]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1217.8757440000006,806.7131704999999],"typeId":"21a0a3b7-bfd8-4958-92f9-fb21adb71ce0","componentVersion":1,"instanceId":"d7e83964-79f2-4e6f-ab07-dee67fd9dff8","orientation":"right","circleData":[[1247.5,650],[1228.2216325000002,649.5517129999998],[1207.5982270000002,649.5517129999998],[1187.4231685,648.6550204999999],[1292.7818110000003,925.7259259999998],[1216.5649210000001,924.3808864999999],[1141.2446650000002,923.0359054999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1667.8757440000002,806.7131704999999],"typeId":"21a0a3b7-bfd8-4958-92f9-fb21adb71ce0","componentVersion":1,"instanceId":"6bde5401-8877-4618-b129-167654a129ea","orientation":"right","circleData":[[1697.5,650],[1678.2216325000002,649.5517129999998],[1657.5982270000002,649.5517129999998],[1637.4231685,648.6550204999999],[1742.7818110000003,925.7259259999998],[1666.5649210000001,924.3808864999999],[1591.2446650000002,923.0359055000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"N","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[3393.359241444308,610.2637795986323],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"786922c4-3cc4-4e2e-a1af-6f582a726cc5","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"L","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[3497.068721174747,610.9967802938991],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"c6b89f01-cd33-4f53-a410-bd8ce0a19726","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"LOAD 1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[1517.1631976795416,2554.4111373325836],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"028c5ed6-a9ce-4916-bd5a-20a0af91ff53","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"LOAD 2","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[1050.1295299873186,2562.8970818848297],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"d8ee4efe-302f-41eb-a87d-4235620299ce","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Dimmer\nOutput 2","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[1023.8439203020007,795.1529920546972],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"8c415f8f-024b-42a7-9906-fa5d9103b190","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Dimmer\nOutput 1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[1483.0932434380895,794.8020298127515],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"f0886e27-8ec0-43da-a659-1cbab4912d9c","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[3006.71431,2014.5000244999999],"typeId":"5ce5e9a0-0484-4e7a-b171-46d0c4edfd48","componentVersion":2,"instanceId":"9b271475-bebe-41b8-aded-20e21ef4734b","orientation":"up","circleData":[[2987.5,1850],[3029.499982,1850.8571344999998],[2986.6428895,2182.999983499998],[3030.7857474999996,2183.8571599999987]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[285.6014590000002,751.6867490000006],"typeId":"babbe5d2-1338-4c89-b876-1df438752dc0","componentVersion":1,"instanceId":"fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351","orientation":"down","circleData":[[347.5,545],[313.61446750000005,544.5481685000004],[279.7289364999997,544.0963970000003],[246.29517699999997,544.0963970000003],[460,927.2289364999999],[254.4277165000001,923.6144689999999],[383.64456700000005,922.2590345000001],[323.5542114999996,922.2590345000001],[191.17472349999997,922.2590345000001],[130.1807079999997,923.1626374999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"YaSolR AC Circuit\n(behind a breaker)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[3012.4637827603738,1911.511553397949],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"60b47335-97ed-4e17-861d-700ea31fb823","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[3442.3552975000002,484.8953134999997],"typeId":"c2a09f2b-df40-42a6-8e0c-c519ba38e9d5","componentVersion":1,"instanceId":"d53bc8d1-adbf-42c3-9bdc-27d4d2b68588","orientation":"up","circleData":[[3437.5,350],[3453.0759055000003,351.3743885],[3453.9921460000005,604.2539555000001],[3440.706811,605.6282870000002]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"L1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[459.35242794409623,850.1271975814917],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"1d273ddc-00fe-4e0d-abfe-19b515681189","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"LOAD1\n(NO)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[395.811935358053,841.8286595350996],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"ff8b35db-2369-4252-b747-2b8feb913443","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"DIM1\n(NC)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[321.27957508862346,842.3526361219355],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"5830f988-bcfc-482c-9025-2453ea0e5d91","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"L2","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[249.8597377121365,834.0709109984225],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"27a36091-2d09-4701-aaa6-228dbe3a2a98","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"LOAD2\n(NO)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[191.8459995160615,836.825881731967],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"14cfe2b5-1a7f-43d4-89f6-507c0f51956e","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"DIM2\n(NC)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[124.68264509992309,837.349858318803],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"f69e8dbc-a536-4df8-89be-06aad4cf7eb6","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"-864.00000","left":"68.90851","width":"3727.59149","height":"3857.07477","x":"68.90851","y":"-864.00000"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1\",\"endPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24\",\"rawStartPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1\",\"rawEndPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"3453.0759055000_351.3743885000\\\",\\\"3453.0759055000_260.0000000000\\\",\\\"640.0000000000_260.0000000000\\\",\\\"640.0000000000_12.5282165000\\\",\\\"679.1613940000_12.5282165000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1\",\"endPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_1\",\"rawStartPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1\",\"rawEndPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"3453.0759055000_351.3743885000\\\",\\\"3453.0759055000_260.0000000000\\\",\\\"1228.2216325000_260.0000000000\\\",\\\"1228.2216325000_649.5517130000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_1\",\"endPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1\",\"rawStartPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_1\",\"rawEndPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1678.2216325000_649.5517130000\\\",\\\"1678.2216325000_260.0000000000\\\",\\\"3453.0759055000_260.0000000000\\\",\\\"3453.0759055000_351.3743885000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1\",\"endPinId\":\"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_1\",\"rawStartPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1\",\"rawEndPinId\":\"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"3453.0759055000_351.3743885000\\\",\\\"3452.5000000000_351.3743885000\\\",\\\"3452.5000000000_260.0000000000\\\",\\\"317.5000000000_260.0000000000\\\",\\\"317.5000000000_537.5000000000\\\",\\\"313.6144675000_537.5000000000\\\",\\\"313.6144675000_544.5481685000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0\",\"endPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19\",\"rawStartPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0\",\"rawEndPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"3437.5000000000_350.0000000000\\\",\\\"3437.5000000000_282.5000000000\\\",\\\"617.5000000000_282.5000000000\\\",\\\"617.5000000000_148.1934635000\\\",\\\"678.5382805000_148.1934635000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0\",\"endPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_0\",\"rawStartPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0\",\"rawEndPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"3437.5000000000_350.0000000000\\\",\\\"3437.5000000000_282.5000000000\\\",\\\"1247.5000000000_282.5000000000\\\",\\\"1247.5000000000_650.0000000000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_0\",\"endPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0\",\"rawStartPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_0\",\"rawEndPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1697.5000000000_650.0000000000\\\",\\\"1697.5000000000_282.5000000000\\\",\\\"3437.5000000000_282.5000000000\\\",\\\"3437.5000000000_350.0000000000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0\",\"endPinId\":\"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_0\",\"rawStartPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0\",\"rawEndPinId\":\"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"3437.5000000000_350.0000000000\\\",\\\"3437.5000000000_282.5000000000\\\",\\\"347.5000000000_282.5000000000\\\",\\\"347.5000000000_545.0000000000\\\"]}\"}","{\"color\":\"#0076FF\",\"startPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0\",\"endPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0\",\"rawStartPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0\",\"rawEndPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2987.5000000000_1145.0000000000\\\",\\\"2747.5000000000_1145.0000000000\\\",\\\"2747.5000000000_1625.0000000000\\\"]}\"}","{\"color\":\"#0076FF\",\"startPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0\",\"endPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0\",\"rawStartPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0\",\"rawEndPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2507.5000000000_1430.0000000000\\\",\\\"2507.5000000000_1145.0000000000\\\",\\\"2987.5000000000_1145.0000000000\\\"]}\"}","{\"color\":\"#0076FF\",\"startPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0\",\"endPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0\",\"rawStartPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0\",\"rawEndPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2987.5000000000_1145.0000000000\\\",\\\"2987.5000000000_1850.0000000000\\\"]}\"}","{\"color\":\"#85A900\",\"startPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1\",\"endPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1\",\"rawStartPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1\",\"rawEndPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2544.3571255000_1429.1428745000\\\",\\\"2544.3571255000_1310.0000000000\\\",\\\"3317.5000000000_1310.0000000000\\\",\\\"3317.5000000000_1145.0000000000\\\",\\\"3259.5265000000_1145.0000000000\\\"]}\"}","{\"color\":\"#85A900\",\"startPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1\",\"endPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1\",\"rawStartPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1\",\"rawEndPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"3259.5265000000_1145.0000000000\\\",\\\"3317.5000000000_1145.0000000000\\\",\\\"3317.5000000000_1310.0000000000\\\",\\\"2784.3571255000_1310.0000000000\\\",\\\"2784.3571255000_1624.1428745000\\\"]}\"}","{\"color\":\"#85A900\",\"startPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1\",\"endPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1\",\"rawStartPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1\",\"rawEndPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"3259.5265000000_1145.0000000000\\\",\\\"3317.5000000000_1145.0000000000\\\",\\\"3317.5000000000_1310.0000000000\\\",\\\"3032.5000000000_1310.0000000000\\\",\\\"3032.5000000000_1850.8571345000\\\",\\\"3029.4999820000_1850.8571345000\\\"]}\"}","{\"color\":\"#00FFC6\",\"startPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2\",\"endPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3\",\"rawStartPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2\",\"rawEndPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2986.6428895000_2182.9999835000\\\",\\\"2986.6428895000_2262.5000000000\\\",\\\"3437.5000000000_2262.5000000000\\\",\\\"3437.5000000000_605.6282870000\\\",\\\"3440.7068110000_605.6282870000\\\"]}\"}","{\"color\":\"#FF6E41\",\"startPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3\",\"endPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2\",\"rawStartPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3\",\"rawEndPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"3030.7857475000_2183.8571600000\\\",\\\"3032.5000000000_2183.8571600000\\\",\\\"3032.5000000000_2277.5000000000\\\",\\\"3453.9921460000_2277.5000000000\\\",\\\"3453.9921460000_604.2539555000\\\"]}\"}","{\"color\":\"#E85EBE\",\"startPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3\",\"endPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_5\",\"rawStartPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3\",\"rawEndPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2509.6428145000_1753.1428745000\\\",\\\"2509.6428145000_1895.0000000000\\\",\\\"1622.5000000000_1895.0000000000\\\",\\\"1622.5000000000_1010.0000000000\\\",\\\"1666.5649210000_1010.0000000000\\\",\\\"1666.5649210000_924.3808865000\\\"]}\"}","{\"color\":\"#E85EBE\",\"startPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3\",\"endPinId\":\"pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2\",\"rawStartPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3\",\"rawEndPinId\":\"pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2509.6428145000_1753.1428745000\\\",\\\"2509.6428145000_1895.0000000000\\\",\\\"1622.5000000000_1895.0000000000\\\",\\\"1622.5000000000_2405.0000000000\\\"]}\"}","{\"color\":\"#010067\",\"startPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3\",\"endPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_5\",\"rawStartPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3\",\"rawEndPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2749.6428145000_1948.1428745000\\\",\\\"2749.6428145000_2165.0000000000\\\",\\\"1172.5000000000_2165.0000000000\\\",\\\"1172.5000000000_1010.0000000000\\\",\\\"1216.5649210000_1010.0000000000\\\",\\\"1216.5649210000_924.3808865000\\\"]}\"}","{\"color\":\"#010067\",\"startPinId\":\"pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2\",\"endPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3\",\"rawStartPinId\":\"pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2\",\"rawEndPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1172.5000000000_2420.0000000000\\\",\\\"1172.5000000000_2165.0000000000\\\",\\\"2749.6428145000_2165.0000000000\\\",\\\"2749.6428145000_1948.1428745000\\\"]}\"}","{\"color\":\"#FFE502\",\"startPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_6\",\"endPinId\":\"pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1\",\"rawStartPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_6\",\"rawEndPinId\":\"pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1591.2446650000_923.0359055000\\\",\\\"1591.2446650000_2405.0000000000\\\",\\\"1592.5000000000_2405.0000000000\\\"]}\"}","{\"color\":\"#FFE502\",\"startPinId\":\"pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1\",\"endPinId\":\"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_6\",\"rawStartPinId\":\"pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1\",\"rawEndPinId\":\"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_6\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1592.5000000000_2405.0000000000\\\",\\\"1592.5000000000_1895.0000000000\\\",\\\"383.6445670000_1895.0000000000\\\",\\\"383.6445670000_922.2590345000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1\",\"endPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_6\",\"rawStartPinId\":\"pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1\",\"rawEndPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_6\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1142.5000000000_2420.0000000000\\\",\\\"1141.2446650000_2420.0000000000\\\",\\\"1141.2446650000_923.0359055000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1\",\"endPinId\":\"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_8\",\"rawStartPinId\":\"pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1\",\"rawEndPinId\":\"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_8\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1142.5000000000_2420.0000000000\\\",\\\"1142.5000000000_2165.0000000000\\\",\\\"191.1747235000_2165.0000000000\\\",\\\"191.1747235000_922.2590345000\\\"]}\"}","{\"color\":\"#001544\",\"startPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_3\",\"endPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28\",\"rawStartPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_3\",\"rawEndPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1187.4231685000_648.6550205000\\\",\\\"1187.4231685000_-467.5000000000\\\",\\\"550.0000000000_-467.5000000000\\\",\\\"550.0000000000_-95.9164615000\\\",\\\"677.9352805000_-95.9164615000\\\"]}\"}","{\"color\":\"#91D0CB\",\"startPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_3\",\"endPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29\",\"rawStartPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_3\",\"rawEndPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1637.4231685000_648.6550205000\\\",\\\"1637.4231685000_-497.5000000000\\\",\\\"587.5000000000_-497.5000000000\\\",\\\"587.5000000000_-121.9526425000\\\",\\\"677.3322805000_-121.9526425000\\\"]}\"}","{\"color\":\"#007DB5\",\"startPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_2\",\"endPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32\",\"rawStartPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_2\",\"rawEndPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1207.5982270000_649.5517130000\\\",\\\"1207.5982270000_-527.5000000000\\\",\\\"617.5000000000_-527.5000000000\\\",\\\"617.5000000000_-203.7140260000\\\",\\\"678.5583940000_-203.7140260000\\\"]}\"}","{\"color\":\"#007DB5\",\"startPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_2\",\"endPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32\",\"rawStartPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_2\",\"rawEndPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1657.5982270000_649.5517130000\\\",\\\"1657.5982270000_-527.5000000000\\\",\\\"617.5000000000_-527.5000000000\\\",\\\"617.5000000000_-203.7140260000\\\",\\\"678.5583940000_-203.7140260000\\\"]}\"}","{\"color\":\"#5FAD4E\",\"startPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_31\",\"endPinId\":\"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_2\",\"rawStartPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_31\",\"rawEndPinId\":\"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"677.3121670000_-176.4532315000\\\",\\\"280.0000000000_-176.4532315000\\\",\\\"280.0000000000_537.5000000000\\\",\\\"279.7289365000_537.5000000000\\\",\\\"279.7289365000_544.0963970000\\\"]}\"}","{\"color\":\"#FF029D\",\"startPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_30\",\"endPinId\":\"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_3\",\"rawStartPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_30\",\"rawEndPinId\":\"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"677.3322805000_-149.8179370000\\\",\\\"242.5000000000_-149.8179370000\\\",\\\"242.5000000000_545.0000000000\\\",\\\"246.2951770000_545.0000000000\\\",\\\"246.2951770000_544.0963970000\\\"]}\"}","{\"color\":\"#683D3B\",\"startPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2\",\"endPinId\":\"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_4\",\"rawStartPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2\",\"rawEndPinId\":\"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2545.6428145000_1755.2857490000\\\",\\\"2552.5000000000_1755.2857490000\\\",\\\"2552.5000000000_1842.5000000000\\\",\\\"452.5000000000_1842.5000000000\\\",\\\"452.5000000000_927.2289365000\\\",\\\"460.0000000000_927.2289365000\\\"]}\"}","{\"color\":\"#FF74A3\",\"startPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4\",\"endPinId\":\"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_7\",\"rawStartPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4\",\"rawEndPinId\":\"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_7\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1742.7818110000_925.7259260000\\\",\\\"1742.5000000000_925.7259260000\\\",\\\"1742.5000000000_1955.0000000000\\\",\\\"323.5542115000_1955.0000000000\\\",\\\"323.5542115000_922.2590345000\\\"]}\"}","{\"color\":\"#968AE8\",\"startPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4\",\"endPinId\":\"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_9\",\"rawStartPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4\",\"rawEndPinId\":\"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_9\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1292.7818110000_925.7259260000\\\",\\\"1292.5000000000_925.7259260000\\\",\\\"1292.5000000000_2232.5000000000\\\",\\\"130.0000000000_2232.5000000000\\\",\\\"130.0000000000_923.1626375000\\\",\\\"130.1807080000_923.1626375000\\\"]}\"}","{\"color\":\"#98FF52\",\"startPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2\",\"endPinId\":\"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_5\",\"rawStartPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2\",\"rawEndPinId\":\"pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2785.6428145000_1950.2857490000\\\",\\\"2785.0000000000_1950.2857490000\\\",\\\"2785.0000000000_2112.5000000000\\\",\\\"254.4277165000_2112.5000000000\\\",\\\"254.4277165000_923.6144690000\\\"]}\"}"],"projectDescription":""}PK
     mdZ               jsons/PK
     mdZAT?{  ?{     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"ESP32 Devkit V4","category":["User Defined"],"id":"b975acdd-73e3-4b18-a5a5-9b66f369afa0","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"ae82c023-d9d4-4942-aa8d-ab2ae3c53d73.png","iconPic":"cbf7ad0e-0f08-44f8-98a9-dcbe92af212f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"48.00864","numDisplayRows":"48.00864","pins":[{"uniquePinIdString":"0","positionMil":"3273.41401,3905.84495","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"3277.43401,3724.10632","isAnchorPin":false,"label":"23"},{"uniquePinIdString":"2","positionMil":"3277.56810,3550.53178","isAnchorPin":false,"label":"22"},{"uniquePinIdString":"3","positionMil":"3273.41401,3360.60905","isAnchorPin":false,"label":"TX"},{"uniquePinIdString":"4","positionMil":"3281.58810,3187.03451","isAnchorPin":false,"label":"RX"},{"uniquePinIdString":"5","positionMil":"3273.41401,3013.32588","isAnchorPin":false,"label":"21"},{"uniquePinIdString":"6","positionMil":"3281.58810,2827.55725","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"7","positionMil":"3281.58810,2653.98271","isAnchorPin":false,"label":"19"},{"uniquePinIdString":"8","positionMil":"3281.58810,2472.24408","isAnchorPin":false,"label":"18"},{"uniquePinIdString":"9","positionMil":"3277.43401,2302.84954","isAnchorPin":false,"label":"5"},{"uniquePinIdString":"10","positionMil":"3285.60810,2117.08091","isAnchorPin":false,"label":"17"},{"uniquePinIdString":"11","positionMil":"3285.60810,1935.33228","isAnchorPin":false,"label":"16"},{"uniquePinIdString":"12","positionMil":"3285.60810,1749.58956","isAnchorPin":false,"label":"4"},{"uniquePinIdString":"13","positionMil":"3289.61810,1576.02502","isAnchorPin":false,"label":"0"},{"uniquePinIdString":"14","positionMil":"3285.60810,1402.58457","isAnchorPin":false,"label":"2"},{"uniquePinIdString":"15","positionMil":"3293.78219,1208.50775","isAnchorPin":false,"label":"15"},{"uniquePinIdString":"16","positionMil":"3289.61810,1034.93321","isAnchorPin":false,"label":"D1"},{"uniquePinIdString":"17","positionMil":"3289.61810,849.03049","isAnchorPin":false,"label":"D0"},{"uniquePinIdString":"18","positionMil":"3301.95628,659.25186","isAnchorPin":false,"label":"CLK"},{"uniquePinIdString":"19","positionMil":"1480.33588,651.22186","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"20","positionMil":"1472.16179,836.98049","isAnchorPin":false,"label":"CMD"},{"uniquePinIdString":"21","positionMil":"1480.33588,1010.55503","isAnchorPin":false,"label":"D3"},{"uniquePinIdString":"22","positionMil":"1476.31588,1196.31366","isAnchorPin":false,"label":"D2"},{"uniquePinIdString":"23","positionMil":"1476.31588,1378.06229","isAnchorPin":false,"label":"13"},{"uniquePinIdString":"24","positionMil":"1484.48997,1555.65684","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"25","positionMil":"1480.33588,1733.38547","isAnchorPin":false,"label":"12"},{"uniquePinIdString":"26","positionMil":"1484.48997,1927.46228","isAnchorPin":false,"label":"14"},{"uniquePinIdString":"27","positionMil":"1476.31588,2109.06682","isAnchorPin":false,"label":"27"},{"uniquePinIdString":"28","positionMil":"1476.31588,2278.62136","isAnchorPin":false,"label":"26"},{"uniquePinIdString":"29","positionMil":"1472.29588,2452.19590","isAnchorPin":false,"label":"25"},{"uniquePinIdString":"30","positionMil":"1472.29588,2637.96453","isAnchorPin":false,"label":"33"},{"uniquePinIdString":"31","positionMil":"1472.16179,2815.53316","isAnchorPin":false,"label":"32"},{"uniquePinIdString":"32","positionMil":"1480.46997,2997.27179","isAnchorPin":false,"label":"35"},{"uniquePinIdString":"33","positionMil":"1472.29588,3170.71224","isAnchorPin":false,"label":"34"},{"uniquePinIdString":"34","positionMil":"1459.96384,3364.79179","isAnchorPin":false,"label":"VIN"},{"uniquePinIdString":"35","positionMil":"1472.29588,3534.47769","isAnchorPin":false,"label":"VP"},{"uniquePinIdString":"36","positionMil":"1476.31384,3711.93179","isAnchorPin":false,"label":"EN"},{"uniquePinIdString":"37","positionMil":"1472.29588,3897.67086","isAnchorPin":false,"label":"3V3"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Water Heater","category":["User Defined"],"id":"fa95e5d1-b92a-410f-a873-a71d0089e7ad","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"85e66502-362d-4a26-afcd-97fbc4859675.png","iconPic":"b13518ba-21c5-4f60-a735-1d8041d11d7b.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"39.37008","numDisplayRows":"39.37008","pins":[{"uniquePinIdString":"0","positionMil":"25453.83178,-12736.88404","isAnchorPin":true,"label":""},{"uniquePinIdString":"1","positionMil":"3753.83178,1863.11596","isAnchorPin":false,"label":"V+"},{"uniquePinIdString":"2","positionMil":"3753.83178,1663.11596","isAnchorPin":false,"label":"V-"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Water Heater","category":["User Defined"],"id":"fa95e5d1-b92a-410f-a873-a71d0089e7ad","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"85e66502-362d-4a26-afcd-97fbc4859675.png","iconPic":"b13518ba-21c5-4f60-a735-1d8041d11d7b.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"39.37008","numDisplayRows":"39.37008","pins":[{"uniquePinIdString":"0","positionMil":"25453.83178,-12736.88404","isAnchorPin":true,"label":""},{"uniquePinIdString":"1","positionMil":"3753.83178,1863.11596","isAnchorPin":false,"label":"V+"},{"uniquePinIdString":"2","positionMil":"3753.83178,1663.11596","isAnchorPin":false,"label":"V-"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Alternative Current (AC) - Large","category":["User Defined"],"id":"5ac8a9e5-bb24-45ef-9b03-1161364522fb","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"8a1d81a5-79d4-450c-9f72-108cd2673013.png","iconPic":"aacc0029-e57d-4614-a443-d9bee65b5175.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"23.63677","numDisplayRows":"22.90067","pins":[{"uniquePinIdString":"0","positionMil":"277.14723,1228.19938","isAnchorPin":true,"label":"Neutral"},{"uniquePinIdString":"1","positionMil":"2090.65723,1228.19938","isAnchorPin":false,"label":"Line"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Breaker 20A","category":["User Defined"],"id":"a64016c8-4d9c-491e-ba46-f626b2aeb38c","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1d90a712-93d7-4555-ae10-1782f839eba3.png","iconPic":"e5551f5a-2fb7-4493-9527-57db21faeaae.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.69291","numDisplayRows":"28.74016","pins":[{"uniquePinIdString":"0","positionMil":"192.35433,2457.96024","isAnchorPin":true,"label":"N"},{"uniquePinIdString":"1","positionMil":"438.06850,2463.67441","isAnchorPin":false,"label":"L"},{"uniquePinIdString":"2","positionMil":"446.63976,289.38858","isAnchorPin":false,"label":"L"},{"uniquePinIdString":"3","positionMil":"206.63976,303.67441","isAnchorPin":false,"label":"N"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Breaker 20A","category":["User Defined"],"id":"a64016c8-4d9c-491e-ba46-f626b2aeb38c","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1d90a712-93d7-4555-ae10-1782f839eba3.png","iconPic":"e5551f5a-2fb7-4493-9527-57db21faeaae.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.69291","numDisplayRows":"28.74016","pins":[{"uniquePinIdString":"0","positionMil":"192.35433,2457.96024","isAnchorPin":true,"label":"N"},{"uniquePinIdString":"1","positionMil":"438.06850,2463.67441","isAnchorPin":false,"label":"L"},{"uniquePinIdString":"2","positionMil":"446.63976,289.38858","isAnchorPin":false,"label":"L"},{"uniquePinIdString":"3","positionMil":"206.63976,303.67441","isAnchorPin":false,"label":"N"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Robodyn 16/24A","category":["User Defined"],"id":"21a0a3b7-bfd8-4958-92f9-fb21adb71ce0","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"ae036c7f-e258-4627-a75d-99715ec815e7.png","iconPic":"69c28b0d-a0ad-46f0-a190-03e6ecfe42fd.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"23.62205","numDisplayRows":"16.53543","pins":[{"uniquePinIdString":"0","positionMil":"136.34803,1024.26654","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"133.35945,895.74409","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"2","positionMil":"133.35945,758.25472","isAnchorPin":false,"label":"ZC"},{"uniquePinIdString":"3","positionMil":"127.38150,623.75433","isAnchorPin":false,"label":"PSM"},{"uniquePinIdString":"4","positionMil":"1974.52087,1326.14528","isAnchorPin":false,"label":"L"},{"uniquePinIdString":"5","positionMil":"1965.55394,818.03268","isAnchorPin":false,"label":"N"},{"uniquePinIdString":"6","positionMil":"1956.58740,315.89764","isAnchorPin":false,"label":"LOAD"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Robodyn 16/24A","category":["User Defined"],"id":"21a0a3b7-bfd8-4958-92f9-fb21adb71ce0","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"ae036c7f-e258-4627-a75d-99715ec815e7.png","iconPic":"69c28b0d-a0ad-46f0-a190-03e6ecfe42fd.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"23.62205","numDisplayRows":"16.53543","pins":[{"uniquePinIdString":"0","positionMil":"136.34803,1024.26654","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"133.35945,895.74409","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"2","positionMil":"133.35945,758.25472","isAnchorPin":false,"label":"ZC"},{"uniquePinIdString":"3","positionMil":"127.38150,623.75433","isAnchorPin":false,"label":"PSM"},{"uniquePinIdString":"4","positionMil":"1974.52087,1326.14528","isAnchorPin":false,"label":"L"},{"uniquePinIdString":"5","positionMil":"1965.55394,818.03268","isAnchorPin":false,"label":"N"},{"uniquePinIdString":"6","positionMil":"1956.58740,315.89764","isAnchorPin":false,"label":"LOAD"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Breaker 2A","category":["User Defined"],"id":"5ce5e9a0-0484-4e7a-b171-46d0c4edfd48","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"a038ca8d-f9eb-4e93-ad0b-b831193aa106.png","iconPic":"3e0a96b2-ef1c-4fb2-8b57-d71cbe1f3744.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"28.33333","pins":[{"uniquePinIdString":"0","positionMil":"205.23810,2513.33333","isAnchorPin":true,"label":"N"},{"uniquePinIdString":"1","positionMil":"485.23798,2507.61910","isAnchorPin":false,"label":"L"},{"uniquePinIdString":"2","positionMil":"199.52403,293.33344","isAnchorPin":false,"label":"N"},{"uniquePinIdString":"3","positionMil":"493.80975,287.61893","isAnchorPin":false,"label":"L"}],"pinType":"wired"},"properties":[]},{"subtypeName":"2 Channel 30A AC Relay 5V DC Control","category":["User Defined"],"id":"babbe5d2-1338-4c89-b876-1df438752dc0","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"ac27922a-fd15-40ea-8551-3be3f9cd5316.png","iconPic":"49e5ee10-9185-4279-8a25-10889e7bb4ef.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"27.55906","numDisplayRows":"31.49606","pins":[{"uniquePinIdString":"0","positionMil":"965.29606,196.89134","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"1191.19961,193.87913","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"2","positionMil":"1417.10315,190.86732","isAnchorPin":false,"label":"CH1"},{"uniquePinIdString":"3","positionMil":"1639.99488,190.86732","isAnchorPin":false,"label":"CH2"},{"uniquePinIdString":"4","positionMil":"215.29606,2745.08425","isAnchorPin":false,"label":"L1"},{"uniquePinIdString":"5","positionMil":"1585.77795,2720.98780","isAnchorPin":false,"label":"L2"},{"uniquePinIdString":"6","positionMil":"724.33228,2711.95157","isAnchorPin":false,"label":"NO1"},{"uniquePinIdString":"7","positionMil":"1124.93465,2711.95157","isAnchorPin":false,"label":"NC1"},{"uniquePinIdString":"8","positionMil":"2007.46457,2711.95157","isAnchorPin":false,"label":"NO2"},{"uniquePinIdString":"9","positionMil":"2414.09134,2717.97559","isAnchorPin":false,"label":"NC2"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"HDR-15-5 5V 2.4A","category":["User Defined"],"id":"c2a09f2b-df40-42a6-8e0c-c519ba38e9d5","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"cff7cff8-0125-49f3-ae91-9e6ccc0a4cc7.png","iconPic":"7b19d218-2217-455d-9a43-b73a208c2c5c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.54331","numDisplayRows":"21.25984","pins":[{"uniquePinIdString":"0","positionMil":"144.79685,1962.29409","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"248.63622,1953.13150","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"2","positionMil":"254.74449,267.26772","isAnchorPin":false,"label":"L"},{"uniquePinIdString":"3","positionMil":"166.17559,258.10551","isAnchorPin":false,"label":"N"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"}]}PK
     mdZ               images/PK
     mdZ�&�y`  y`  /   images/8c2f1315-cf23-4ba8-a920-becb97f13280.png�PNG

   IHDR  �  �   ��ߊ  NiCCPicc  (�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D�0գ ����d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c�%��V��h���ʢ��G`(�*x�%��(�30����s 8,�� Ě�30������n���~��@�\;b��'v$%�����)-����r�H�@=��i�F`yF'�{��Vc``����w�������w1P��y !e��?C    cHRM  z&  ��  �   ��  u0  �`  :�  p��Q<   bKGD      �C�   	pHYs  %  %IR$�   tIME�WxG  �zTXtRaw profile type icc  8��S[n�0��)z^�8~$R��b;^eWݪ��HQb�0$|�>�� D�h`�dZ@�&F�Ąb�9��m��P=Eec������O8��`��Й�f�
�Q�A:���{�xt�k��7�����������-eP/���\!�����jS�u�mۃ��Qa;��B�["�,FدCl֤�	�����/�&�S�T�c��\���~�y�_���D6:J&�D�z����f5u�R�����Ye:�010�����?1:9�����{��5nH����^υZ�w�R��WU(5G�Ӫu2j�fo�-���)�:&c*+q�y&�"J��G��|/��d�c?&s&]����VG��^q���@����줁/0�   orNTϢw�  [5IDATx���w|e���3[�����!�XQ�	6�g׻��;�ӟ�SO�]�Slxީ��)6Գ��^C��m7����cӳ��؅|ޯ����y����S�y """"""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""�P �t뎇yX��s*�+��������L����>����<�r�ݵ/�ϯj>��ߌ�	�\51�;Z�w�e[�L�>��( ��R�	�NUo��W{��v��	댍
�_�f�|����Io[����7�9	s� W�>����&A����@��H��t@U���"^ n@U���^}z/[�j�[�*)9����n͚?VTV����� �*�, 4 ��{!��yLDDtX2�I�+�|���5]�dݸy����S�NMX�˯����^!"Z�SNDDDው�]8|�+LUU�S�
�n�u=&҉"""�����]bc�L������H'����ZND��fK�<�M��DDD p�ݚf���*(w��CDDD��%�$ϷX��'0���������p��a���ʓ<���#������	E��Qn������iӶ/[�lBaaAV�`�Դ48��vX�6�-fh�	�R�4J)(�L�O""":t��r�];���T�r:��'O�����z��:<7<O�����F�ۍ��*����v����"�_A��jf"��r�|��������Z�����=v�m����X5z4LZx�Ͱ�����QCrTAii)~[�+¹1k���e�E���;���^�&���� ""��:Z،m�tV��r�}^_��✕Nx�^�m�H�Q�6�5�_�6���At�z�^{�7].��#�WDDD������[u�ޤ�r9�q{"�F"""j����"b�-��t:]p{8�Q��JJK��x��.��o�\.x<,�E9�

�i*^=x@w��NDD��VPX �������}U�z<p�\�N'5C++)���r��~S�7}>*++#�F"""j� n��&"M����|��`@'""�f
�����D����>�,�E5AM	��������r��t:���(4��r� Ȉx>�N�3҉$""�������3ƌm��.�x��N%�������/ �y9�9Q���M������NDD�4 PJٍ�������(��@([�6t �z}0z������h 4��^�����(�i�ee����h�����(�iK�-W*D@�1�E=m����R�b� �Љ�����_�� t�"A��#""����+ �ϡ�ʝ��(�VZV��H�*w/D�H'����B�*�˕@LFx}>��NDD��VQY�D�Y�NDD����
��q@���;Q��*]N��!��%t�t""�h%М��J�u�h_u�8>�FDD��9�����_g/w""�h�UU���S�����G:�DDDdD��j5���~?K�DDDQK ��p�tݯCg�;Q4�b��b�W]t�)���(�i�����]��:QT�L���]ס�|
���(�i��LP�0��܉������2�fJ�r'""�j�)(���ua�;Q��bR
!:�܉���� �DD���ʝ��(�iգ�i0�OM�r'""�v͖�u]X�NDD��u*��^]B��܉����V=u��-�p`""��&uݸ�΁e������h~����*w""�����z���*w""��%���u%Ͷ���NDD�4�߯A� �+�C�)���(�i�߯��ϡE9i��5v�#""�~���J`\�.�NqDDD�N��	�)NNDD��l6[�����DDDQ�l65�`@oW�3[j^���&��Q ""#f��dX�~0�d������%سgv�؅��TTT������PJ�n�!11�������dt���D��@��!"�:��i!K�pr�V��"((,Ěu��ӏ?a�����ۊ����^�'��P�Q�4M�f��EJj*�w�#�c���5j��2a�4v":�(���fM�̡2N �ro!���b�ڵ���O���o�v�Z@��hI��� �z������ck�f,��������ӦM������b6��'�#�P\Z
�łX�#��9|Ĭ�BV�C�ϡ�I��x�d�R�=�m|�ɧض5��Q��V����TT�c�o��t����o�����_���{�]-��O7���������Wa�QG��f���x�� ��ZM�mݶ/�y�y��صk'�5�촭ܚ��-�7���Ǘ�č�wfL����/ 6j���m؀_|	�����xp�e�F:i�10�\�˄� ��n|��x�����Ͽ���"�U�&-��]��ۢ_񧫯��͛q�5� 1>�A����PXT�w�{���?�r�
��Gjj:T���d�B�*w�U����r�~�<��S((؏�L�Z���jVb��d�ɤA�4�������!�/�fK!��PX���gݏ��"�|�M蔖ƠNDQ������3�������rV�u!�a���|�8������x����sꝌ0�@n�� 33]�vEnn.�v���D���#&&�*������ �6m�m�6��
?Ȫ�ବ��g�����w/:��3�Q�Q �-[���x6oڈ��/��̀�B����F�}��nǿ��:�^�O�@�edfb�ر�:u
Ǝ���,$$$�j6n�p��(..ƪի��O�����c���5&������ks�"�S:��v8�vu"�:%�%ؿ?����p�Y X�6��҉G}���u��g��Ĥd�:}:���J�1	qq��6�|o�n�!+#Y�p�	���+0g��{�-��0�{=x���w�޸䒋�)~Y�(�(@)��ۋ �D��*wv������չs1�9�s��Q�����s�>��;	qquü����e�&3��G~�>�,r��G]{c
�Ņx���p�B��u ���B��.|l����7��ByY	�s�f2a���x��p��� !>�EA܈ ���p��31���2tx��jؼi#�{�y�UTD:눈�Q  ����]�*w���������];���t9M3��s��3�>��C��K ��f]O���z]�u�qI��g��o�e)�����.��8"�����ޚ��.@m$�q�L��Y�݋�99�3� �8�d���<1P(.*�K/����Bu"�#�D�5����EX�n^|�%���^��c�!�u�,������,7i.��bL�6-d������H��!!DBv3L�ڱK����[�0��<66�˵1l�!{LL $'&��+�D��0*�������?���9�te�:��}8��)R��ys$���~P`��f����+ ;v��']��(�O�<g�uVD��;f��8��S���/5M�����? /o+���m��������z�v���z f�6�V�f��v���G��4x?����|�=p{�����X,�Z��Y�0�L����zo��v��vCD`��`�X`�Xj�o��
��p������v�����������
Ku��6���������vC=��f��6��+_�Q�ן9p����z���`2�`�Xa�Ya�X`�~\���,=F�S�3: ������]�����f�ߚydMi��7"�^@��U�_�V�Z�S+1)_r1R����& 118k�x���QR\��H.5Kh8p� V�\�n�f��}{�b��X�n6oڄ�{������j�"..�ѣ����!''16[�>����rTVV6���dBJr2̍���/,Ě5k�d�lX��w�Fee%|>lV���е[W���#F�@�~����Т������k�d��[�{���鄈��p >>9�9:|��>�{#.6���T^Q�����u��vj����dX-���+*.����d�R�[�;w�Dee%�^o���ƢKv6r��b�0` R��[�6���k׮��ŋ�n�:�ڵ�������|��CVV6C�A߾}���|iN�M� (-+�֭[�v�Z�[�۷oGA~>\UU�z�0�͈�ۑ����]����4p z�쁄��v�ٯ��BIii��RHLH�#&&h^Wy<عs'V�\�իVa˖-�?�W�~�V�������Fnn.�����#==�6/Z���N���w�Ʉ��"��_]�QPX�������M�w8HHH`MBCR�C�r�ϡ+ e��OPU�Q�|���8��qM�Q�0t�|��(�!.>���ӷ/��!C�b�ر�r�]\R�_~]�O?�?��3�mۆ��2��kf�b��%;cǎ��iSq��ǣszzuN���:^y�U��ƛ��PA�Ν�ēO�wϞJ8�v��ǟ|�w�}�V�DaaQ��P0���ԩF�9
^x!N9eb��pj��{�|��gx�w�b�
VO��SV��;w±��/��=��9�Σw�}s^x���"���D<���Z�DFM��8����s���;X�t)
��k���43R��0b�\p��6m*R���-��������罍%K��� ��x;�iiiw�Ѹ���a' 1!�uU�G[�m���_�/���e�q����\}�j��l�Թ3����S�`ҤSЭk�6��*����#f�{����T�Z����o���hpL�UU���_���a���c�8++�)�dAJr2�)S�bƌ��ۧL��>��~̞�>��chZu�Q@iI	����$)�����nGBBB���u]�̙3q���T�� 6�M3�y)���7����DDV�Z%�{��~��i��Vy⩧#�?~]�9/�,g�s������g�Ɇ�����\��{Ӷ��p:�O>���8S��S덑�Ο��T����䤓O���������9�~�����������EV�ZU�Ϊ*y���O�-���XgBb�\vŕ�a㦠i�r{��O?�'�$�Vn'5-]���u�c��V��?�4_�R�����+���RN�<Ebbb[��������s�=_��\ix.y|>���2����kU�$&%˥�_!6mn���{��ǟ��#F��jk��^w�[m12�����?�)

DD�_�jm��x�z�.���9/6ȓ�k��5��t�Y/]-���"�ǞxR��燝��W.�����_8�9���Z<^o�cġ��������W�$&&�Đaß�L����y#�+R���_��ax�euɑ��GE���n�t��oi�t���߸Q�t�%%-�A<�">1I.��R� ~@��_��[��A�dw���V��H~a��q�ݒ�֩Z�~e�&�,�W�j��""%ee���K猬�������-r��dͺu�:���w�(ej���4��O?զ��G�̬�6c%���c�ʏ���$_*�Ny��$�k�6oGi&9a�I�h�v;�}~�|�ͷ2q�d�Z�m<v�C{L��v�Y���E��5�|s޼ꛮ���ify�ŗD�����s5zL�s�m�`���9�] �6l+�=^�\z��횏W]�'��}��|������?Q������UW�)DfBN>e�E]���b�����o����
���ߖ� �9J>��3���%��^�F��W]]�d�%��N�m;vH������n�#��n~�9���d߁�KG���Y�����n�Y���z��q�v���|)���{�%	���S&O����IgU��0�E�V�V.� ��<΁�,���x}�V�Y$t@����""��[�k���u��)S��漼f�π~hzBb��'���) ���X�|E��4�5
I���3\8�o+]�	���j����h�2�>�'PJ�j��j�C�����߭²%���k����~��#L{�R
%�������˯�����뽤�>5�9�K�����|�p&�y��g�tVɳ�o磏>ċ/�����������O<�gf?ge�i�k�O_Kҫ���O=�J�n��=�O<��#(+-#���?�v���k<��l���V���³�<�[n�۷�ե�����Vs�����f��>��Ar���5����Ǜo��nǲ�O?���|vl�Z�/�Ϥ���`�5T�����<���t����ԍe�7z�����c��
�Z.ս�Us1��d^}���طo���v���T����	۟17�p#�6oBM�4���cࠁ9r��� %%�����{����e˰r�J�߿��3X�sN��my����a��q�駵S/V�߇���:�x����n>�c��ХK6z��.�]�*W�����u�VT��:F*�~/��70}�t�\�
�̞�*���vLGl<r��W�^HOOG||<\.v�؉u��a���՝Ϥ�qW������8���o{GB����x�w�rU6�?&�YY��ݻr�� !!n�شi�l1�	@M�2����8��3P\\�G~�����=Ɓ��������HLH�����]��~�z�ܱ>��4źߋyo��̙31n�Q-��χ�^~�f݇Ғ"��:�q�ӧ/F��A�!5-q��p�\(,,D^^.\�u�֡���^fԧa��������O?��G�^�+��+V��9/4� p��!;�z�쉴�t$&&����@����!o�����=�7?�}�]L�>S&�2=�z���Q��i��z�oټ~_��ٌ�}� !>�i�8�ѣG�ꎀTK <d�ˡ�ܭ�yu�kQW�|�_""��J�R�� ��]��E�qy#"�l�
>rt3U=��N��?]#��^�
���Kc~]���b��_�o7��dee7S=	�?`����/-�[�*wM�[u�w���b���㏑'gϖ�+WIqI��=��|��z���R6m�,�ϙ#Æ�Y�e2Yd��iҳw�F���O��N?S�xk�lشY�+*l���T/]&��q���t�?&�U~��v�r�+P��0_Lf��5Z|�Y�t�KU��V�\��m�����2n�1�4S��*M�Lr�Ie����|Qu�㈓I������%kׯ�����RZ^.+V��Y�= �z�}�(��|�m���Z|ο�����_�?q����k�u��r�%��'���?�DN;��z�����������q��R&INN���uHjZ'9��d������������|�t�d�Ν��G˹�/�	I�^�:�).-5L�_MP����{���={e���7ߒ��� �TIrr�����o���g�����҈_'U��_­rOHZ��C��2�[��ʫs����楗_��fx"6\v��uD午HQq��w��m<�����O?�J���bj�""UOu��)�e����8M���v��
����j����Y��n�^�{<�>Էd�r9���͗���ӷ����\)*.iv;^�O���2h�Аy3ᤓ���(�1
���%1)E���FٴeK���˺d��[��$�kwyj�3�?���|��|���d̸�C�ˈQ�e���a狈���;��ԴN��{�!���m�\�����By��g�i�V2��0��)bЛSM4�E�?a�|��gRVQ��^RV&/��buڍ:�)霑)?���;��_~)���Azjj�|���I(��VFe@4x����^y��d`mF����;���I��������W_{Mb�/�J3ɔi�ʪ�k[��""�����s����Dd�G{\���N��E(K^z�U��x������V��s�ꐡ�F�7�~>��|�駒��E�j��v�!�W�{��z]�$����O>U{�nz��Xz����Ss���ǟ��脻��� =z�6؎�������~{��*�\w��B��Kv��2�5qU��[r�麼�����|�8y�ŗZ�
��,\��?ʖ�[�F���뺼��[ҩ�q����Ly��k�9�u>~u������8�����C-�˴��T]�;ŉ�����:nt��	�6�m��{�⥗^FeE�&��0�$<���n� �z����>���f���
��}6nl�����o���a�X��p���>}zXKgfu�=��N8����:e�D�v�ü)(����[�-W �l�⪫��UW���E�2b�p�}��P���>�)�����1c���Z0@� 8��8�����PRR�6��>�ſ�ݷ߁H��i�Ĥ�~���a�Z[tk�z1)�3�8<� :gd��5E���ܹs�s׮��Li�y�L�ݤQ�^����:�L\r�%PZ�c�������QYY����tPi����,p�W����LJr2,Cf����,]�zZ������v+���ݦ�5;��~+����k׮Ň~�E('�|.��RX�ՊI�&!>>�B���p�e�a�)���ՊSN����S�*T���eK{tcǍ��W�16[���I�p�ĉHMKCs=��=�\�}��V.��a�ē���t;^��7o�?���U�|�-�޽��wM3���/�%_sn<�	�g�v���
��֠��t�̟�em�ӑ��7�x:��55�%i�Z,8��sеk�n�桰��]RM��iF�]�H������^�Fb�#��eYE>��C��A߷Xm�����;���_#G��u�]�#�.c�ߋO>����k��� .>]t�SS[�@VV�/�:�v놙3ς�ln�vrs�"-=x��u?���ۜ#5�b����.@���V��O�>�޽[�|t��s�;���k �ٳ'��2�#(..��o�͛7�/�2X�����_	GLL���V��^z	�`�tw��~�	J��ڥ��4Κ9�n�q�>}0d�P��K��Q^V����@4MӚ-��,�+ >�����餶�>o޼K/1XBG߾}q�9g7���-���N��#G���5�VW����_�~?��6�%=-�YY!�9���ѿ�6m'%9ii��RQQVI4�|�ޣ;&L8�MkINJBN׮!�3f���)�@bB:w�l�LEE�z�!�����m��tn2Yp���!77�ݚ�@�=0��i�M���8�&��֩SgL�2fMk�Ͱ �����`�[e����+���n�t́et�������v�M�h�"�ݻ���5�<q"zT�õ�ѹ3N�~�aUdYY~���v	^�G�F�N��Plv;:g�يѣG���>�ݎ��$�������|�0�aÆ!��s`�X���a���0rԨ�Y�ZC!0�_rrJ�|q���1�� 2?��#��`������ĉk�@m/&MÄ	�����7������Ö�����>�+jJ�k׮0����|>����5���DS��b��9}��d��zz�`D�6�Jm�>�-[fp�$��`ʔɭjwn�0q����%���t,Y�eeem*i��V4���`2�[=�i��JHH@�v���b� 6�a����m��3�L8hP��6[B�4����h�a�Á�i�@����.��y�73���}��r�*���>}z�)�F��h���<X��o��xڼ�A�!11��n�SRS`���	H?����%���xU��HE�{ȥ������
@iY6n�h��]�tA�~�Z�w��}���m�6��o�1z����j�����$''#�Kv۷c���tٶ2��j��w�^mi�v�a����ѭ[ז��`;m팚��{��Q�����Ў��� �d�\ߴiS�o^�2�W�ۯ1..��fXD���F��@��r�4MCL��4�i��RXX��;w�߳WO����l����ܾF���cZ;w�j�V���;����iƗ۸��fn��N��:m�v:��m�-�)���X8���(_��~õ%/�e���f�w�.��c��{�n0��ٻg/���߆���vdfd�9��X���ۤ@��TbVJi!�H��J)$��#T�����6�5�G�����W��Ē����؃�̽�d�`2Yj'f���҉��m�F|\<�����q8���9 �)�@�MHH8��c�=D3V������m[�3���Lطw��vA�� JKK���ڪPR\��6m�j�"9%�]�n6��B��v�8m��T�w��)�.���Lf�����t�x��hTPPgee��Lf3����Ih�tɂ�b����$
~���-�;b�i�bs����j|��������l�Z�'���<��~ط��MK�^�O<�8fϞ��-Q�݆�U�ۍ�¶t����G����6��A%f���n ''6�.��N���p:�H	��pQVVVݩ��~
L��z ����d[Uմ)C�u������j6[`1�@��:%��c2���RZ��mP <^o�APD�(5M����P\ܶAZ4�`��5��2�B���9�+ ddd">DUdQQ
�x'-�n�a�f2��#�Q݋�)A��m�Ř�&�ڱ�Б�d2�|�^�V^OscL ����+8]U����J)��C7k��nGm��f�~�m� ������xRTT���o�]�K�1w�*@����]v����9�`>��M碦��E�p�iLGؘ
���>x=��E�"At�vxl�:i��;�q��;���O߾�FGZ�fmTݙn����+QT\]��(Tk���_�W����Y��Pe{�T�����zЎ���@�����G��e�h~������.���?�Ƞ���ʕ+�t���=�����SO>�?���r1l�0�9@NN`2��f����_�QYQ����r��	>8��4�cbjg�"j��M���x���;�<s�O6�f2�K�.�%:�����r��G:��� �>qqq�(����+�}�h���ښ�����_�k�v�ڵ�|���t��@��}0b��u֙8jԨ&�)���i@��������"�t�������QS�z���1��!+���s_������f�s�7� $�znC���#'�+֭]��]Î۱h�t X�~=���P����ʅ���}[�[���郣F�j�ل��m6Tx=h�Ș�������������mSi�Z?8P=�Պ�x�N�U.bc�پ��&�D-��U�!���`����wW�������rE�u֯��n�w().F「�1�2220|����OMI5|F���b���}�m;vT�����l6dtj��̨c3��HO7��N���E����$�/��f[:n@ v��'MBl\��f�-X�e˗G,�
��m��駟AĨ3�`��a�ݫW�w�;�W�����P�t���ׇ���A׃����S�N=/��g�n�6S���;w�t2�ZLucu,��ƌ9
��r��$�iؽk7��{��ko��9֭]���M�7[l�x�)HLH�SSS��c<�Hޖ-(*j�`F�Ôb��͆�$%%��8�D�޽z�f��������o���\�լ1��҉�&��Ն�1�_��.]0i�$(ͨ׫�?��.\tȿ�
���7�xOU]���G�8���1!!}g�Rؽk76���v۶m���[`ti�ѣRSSbNRGҳW/���� ��%%%��}�Y_޶mX�b�nۆ��b������ܩMj&
���a�4�}�L������ְs�v<��c؟�Ⱦ�
�����9/b�0�7�0u�T���ǰm�j6c��Q�XlA�TTT�/�����m��W_c�޽~:j>b���ٶH�{�n�e8߹���k�j��v�n�Tŷ�z�N��3N�g���/�7��x��G�漷QTT��N-"�hh�U�w�*w0h�@�y֙P���_|�^xa\n�!�2~��Wx��W��U������9g�k3�{�1�32��E�W_}��۶��) �������/t�}���aԨ����$
� HMI��1c�&X�����7o�m�/���|�}{�`������x��yx��'q��7�GCE���!Ҵc�:v��b"�Й���z���O���SO>��^zn���u���q���`�>��- e�̙ga��ͮ�o�>}�h�w5l\���|�8� ���ϰl�2�}���aÆ�ܤ�Ƥi8�	HI1�Y�g�~�%K����X��t����7
���!��W`KcƎAff��L&4��XE�9�zˉ&�t�:�s�u�(�_����fw x9�������栢��u��E���K/��=�����/���)^@B\�O�{L�q�=�*<������e����Vᩧ�Fee��{�2aڴi���>�/pth�5
�F�B���a�x��Ǳw��6������W_ᓏ?6\2>!	'Nl�6�H��Ï��5d��i�pJ�S �Ʉ�.��N��C��� ?���|˭؜��n]m�n���G��O�`ѯ��X� 6.��_0hР���ĉ'W_��ض5�� �mk�>) ���C=�իV!xէ��ݻaƌ�T��UM��y�Gl�:�}��'x�٨t�~������u������� F�Q����C�{q$�ڬ0�-���'����9�L��@zj*n����ۯ?�= �P^V���'.��b�2�5�;�ߪ�^���<�}�?p�����K~�6�L8��p޹���, ���p饗��Y澜?7�p#6l�ܪ���k��r�mx��wO0�ɂ/�C�a��iӦ�㏇ѹ��z�ܳ����BQ+{�+z��q�X��Q�UABb2.��rtJK��{�#6[�!x<-Z���΁-��7�_¶�z�����u'2�d�8�+躎_�	�^s-.�݅x~΋X�n=���-�����+1��q��s��#�"����8�N��[n����P�8�t̘1��}]��>�5�_/X �����Ѷj������E���ÿ_��M����
Ǝ�+.�V���$ux�SZ���/��2�.+����ч�M7݌�k�A�0�58�u]���~ß��>��Ð���S&c�ē#�-�L\|b�1�
�}�̛7e�+~]���g���>_�8?3�M)�}��pV:q�m�#��>�zd��t⛯��?���ݻ㨣�°�Cѯ_dee������NTVVb��}X�b%�/[��K�b��mգ�5׏Q0v�8<���գG��� HIN7ހ�k�b�eA�MAD��W_a��u8��p�93�۷/����҉-y[�чa�k�a떼�u5��[�����н{�QZ�șp≸��k0��Y�r9���T��rᕗ_������/�ӦMC�n]g0\���
y[����c�ܹؼqS��<t����IhR������aÆ`�*�ٳ��z����0` ���PU�B~~�?����Zx�_C 1�|�fo6}>�9��!��_|�Ep{<���b��=]j���x�i�zlڸo�a���@bR�6t�\.8�NT�������P�a��`�1������#Z}����1�Y����my0z�g��]x��G��o`���}�hdee!55&MCaQ��ۇ�K�b���عc'�~o�}ё��	����4q�8�ԁ	 �ł���
�v��K/�T�hӠ.��5�W��nǜ9s0|�p�1�3����Ʉ��r�ܹ+W��o�-�֭���y�|�;�#G�0�Y��=z��g�T���G���>� Ji���ǟp".���%%u�<�����}3j�\���
t��	��+VT�*�_l]�QQQ���2��j*��i�-VL;�T�{�=<p`���S�L���p�-�`[�u���;�g�N|�駰X,�X-PJ�������DGVv�����.�I��e��N �$%���^��z�MA�^/�lڈ-�6��wޅ�j��b�����v�ü��93w�uN�1#�W&ҙq��l;v,�5>�a�� O[ri��(,,DrRR�w#z����yUs����eO� j��̳��+�����<�����	��^��=	w������sϴ[0 M�0s�Y�={6F��y>�h�u.��ge%*+*��x�*ԅ-��!C��SO��/�����ړ �����܇��+���{\s><n*+*QYQ��*Wu�i�|��={��G��W\���!��I�N��aC�5 
�����H'?�h��;����Ç���O>�����b�"p��|\�q�2�T���+���;�����[Ӕ©S���W_��.��	�a�W��*���HLJ�e�_��_g�y&,&Z��[�P�+�j:��}�]x��'0t�(MC�`��@5�K�|���<�T�y�E��y��ͭ;އ��.L�s󭷠KvW�$�WTT`ǎ�ޅhn:zs@��4�����)���{������5kQ\T���Z�խ���̒�����1c������ɓjs9XGH <�<3�'O�+���E�����%ψ��GRr
�=�X\tх�4i��ڶ�n<�t�i��� ����4���vj�_�01�N��K]�������X�����¬�z��rI��o�V@lL.��b�;��}|��6o����=?Z�y��5�����_r1.��|dt�Ԧ�]D�=��ů��~=	<�l{��ߪ���f̀���+W���>_+ۨ�ra˖�����ݙux]g@oV�i�='���:\x��X�r%���{���ö��P\T��e0�w0
���I�ջƍ;�L:�F�DjJ2���
s�p��c�ē��w���>ǢE�k�.8t�N�̈��C�^�0��q�2e
�9f<��{���S
�9�2tX�1�u���ܾ0�ZYj����l2��HW�_G��}`j�H_�@�G��1x�Ph����޽{u	�y�6|x�s]ב��[��v���:lx��뺎~���j��b��(���9��_�ѫWO�Z]�S�f@n.f��\x���������`��U(�/���Fs%Jbbc��)Ç����N�	'��ݻäT����d6UUU. "���T8z�V||���Ғ��/8b㐐�ت�6�L�y֙0` ޚ����%��塬��6�( J�`�48bc�������sЩ:�2��w�ݳ;+��_r)^x�y�m6��@M��"(,,Į]��c�l޼�7oF~~>�N'\�@�v��M�`�ِ��Դ4dgg#77����ӻR��`�>�#u,j����Ǝ;�n�:�^�[�n���P^V��
����@\\,233�77���b�����̄�:��~�ʊ
8�Π�[,$&%Ak�ޝ��p��o�j�"!!�p���G���vv����\�W�t���"�{f�III��p�Dee%*&1�-HJJl�픗���r}/��I+_�Q����Rlٲ�ׯ�ڵ�k׮�w��n���!6.q��HLLD�޽1`�@���=�wG|\��;߫�n����=�4�II�߱���xQVVt\�a����M!P�p�@>��m�Ν�p����N@)���!11	����YY����n{}D�_�7<�ԓh�&4&&f����ڳo���P���]��^z1v;z+��]A���x<�z��z���|��|Д����
{LlVk��F��g���������J�l6�b�"�no�6~����/w{m�p����hَ�6u ^�.�^�70��R�X,�Z��Z�������<8X�>(��ߏd-�fa�! ��o�4���p���~���9�4>#�&���b�u����3�Ѳ�m* V�VKBȠ}0��<8�ېF?��z���ЯlCoo��k?�N^�)ԑ�|?��kᡦ��|	��:Q4-�����p�""��$ 4�ërg	���(J�Hӧ2�E9	���e�8""�(&�.͏3�6t""�������Q4-�����:�E�:�5_B�u�����(-�)�D�˝���;���0¿�h�DDD�>�.��V��0�E%DCm�::QTif��z2�E-�$�6tv�#""�Zv/wщ���VJ��DDDQIDD����Љ����ha������(���;#:Q4����3�E)��{�����(j�7�+{�E��&g�s�DDD�K­rg	���(��`�5��E��̶�Q0"��Љ��� ����ֈ���Z�Я�U���;Q��yl��`�XNDD�D��|l���(���Y�NDD�D���NDDtؓ�Oe('""�ja��V�E�0��Y�NDD���ǡ_����[���8�+Q���H�����Ba�;��#�8Rё ���,�E�p��YB'""�b��rg	����c,�j-X�����Vؽ�Չ���V���Y�NDD�X�NDDt`Fu""��ő∈���2s""�(��ʝ����NqDDD�?ζFDDt�p,w""�#B�m��DDD�,��eX�NDD�Z0�E+�GDDt��ќ��(J���;�Љ���Xx%t�r""��֒��։���T�c�3�E%�!"":"�߆.�r'""�V�V�3�E��*�棵��E��c��Z�)�����Yx%t�C'""�R�oF��Z5�ADDD�R-��>s8K�u���()-�����C�D:J!���h]ס (��4�]���������*�]�+@s�	���jE������U�HD�Q�y����>x<(M�b��d6!PFm�밴�����ػ{ws�U���J ��W�1J�DDD�C!�[�* W�߆v�'""�B���Eo""�Ù���G:%DDD�j���tJ�����t@y5�ie�N	�� ���v��H�����ZGӴ����2-%%�q�Ų������#�aK)����φ��F@Ff�q���wy<�" ���j�U�{N�p0:�%@��iͶ�����pD�g?��������9ETM)��R�V��}gm\�a�:����F�~�w��ի��2"V f��b���1&�ɪ�4��4��4�R�T��`B৪��R5WE�T��k�U�f�.�PX�v����RhxW����x9.����R�<\(T�]�R��ԀR����u�V���o5�k���^�=�:Z���Y�~Ԧ���������j��d}J��u�������4��Z��p�	��ʂޠ��^��u��c�o�5��b�x��/=��WD�H�����9��:{�~���������nHBi�{ͪ��R�4����k?���F��w���'��f�!��`geI��5�|M^�~�������4�	��t�cP��V�p��Vw\��n�f�'�z}���`����~i�'|�P������e��e��FK׻�68�W� ۯ9$���dݵ��p����u?t����������K�Y_��]�j�GR/���\�dX �5ikt\��*e�R�p��I�ɋz���ͯ?��ڹ};�~x�W��]��E��O�����FGT},�4��o
 �t]����߯ ݯ+]~�_��D �_W��t%"�~��s��oP՗]��^W�i� ՜ "�7H"XMŊ��>���]���>k��כ����}{��m�9��g���_y�7���4������]�78�J)���x���q�I'��^O���_��5oIݽj��O ��V��b��Ҡ���"5�RR�����R��$5W��;_���U_���BW_]�҅�r��ȁ?���M��r��7�R����d����/U�=}��Li��i
J��MдڿiJA�(/nKE�c}+M� Д��Ai�mk�Mi  ���;�ݨ�j�,��Q{JNIE~�<�쫇q1� ��)[�fʼ^�}>8u14��4��~�AY4(� ~?4ѠC�I5z�_�h�P ���\����k�R
���5��=�j���5�^[k�ª��5�)S��/uWߠ�cG��ɧLz������-���+��s�|6��0٘PRZ��n�/��r�������#F�87--}魷��ߏ�1���d�l����&��-W�ƥd�hT�Qu�T����7��n+�ꭣ�i�h=5�u ́�Oլ\I��������R��ڂQuU��K����[����_�D�N�	�ʹ�p`E���Hmy]�4����P��nOS
�i]��L�u@��lF �X`����*������t�	�v#..J)j|����Kv6X/�y	&�����D|B��v�G�7p9�� Æ��m;v���."�Ꟈ�����?"1�Xi����*���?�㳟�[��E�05�ک���L8�$�������M�Pغu֮] Hk�a꣏?�?���`��������'���Y看��6�sύtr����w��w��[o뒙���a���Lr�=�8"J�""�,\$	tMh��q�ۏ=q¸�YY�>,DD�XB��23�0c�i11��A?.\��Ҳút� l۱w�u֬^��_	������~�o����[o�S�<�$ŀNA���`��1n�ñ�d2]f͚�ض}[���j
@IY|�!|��Wh�p�RSS�>��c^�~��k�N\w�5�N6Q����[t꜉�cƞc�����ݭ�ye��ڎq������#�=.��xi��O�ظ���=�8�#.҇���Y,�SP����٫���7[,֢`�x�.��˯p{�	�>��3<��cpV��q��d6{323������7�Ήtr��Bb@���:�����:u�e�Z����l�2���V��
��U�qｳ�o�n4�(�����G5�I���6nğ��C��MDD�:�>����k猬7��t����N���?6��""���Η���ILL���#G���8"}���ڮ� ��={�]��A���d�'��}��*�G�w��l1A��M&�;;��"���.�sϽ�>DDaa�;��q���d6W[���b��%�r��j�O?��>�,�n����aC_7�Xٳg���H'��(,�d���>Đ��Щs�-��Ш}���8����T�n~߬�p`�^;��11�srr������G�?yB��MDD�>f�s..�������_�UQJRR���oDm���ȁ����f��٭[ϫ����/��F�����EXB��F�����,��>0�}c
%%%X�|y��j�������G|�}�)$%'�w������S&cǎ���D:�DDD�G����?`Ѝ&�E^�����rE])]D��>�N�A�i4��KX5���t���&"":8���[d�tØqGO���F}��a�u���	���`�|�J>r�a0�X�e}r�] ��}���NpDDt�:u��8�̳�&$&m1z=)9U��u������!�͕f����go����s��_o�!�YMD�jlC�f%�$#77woLL���K(���bٲe�Njuj �׋�_��?�F���0��~�j���x��"�t""���G���={?��I����9�|�p:#^Jy��s�vs��Q0hȰ �~c,X�l&"":�j:�6��f��g�"[�n�h@�����#Gs��������w?��r���]wϊt|_|���O�p��Wh�<zbb������v��ϛ����u�ge�?�x�4qR������й�Kq�Eg''��
�5Q�$�=�`Ăys���8�v�=�x(3���"�Ý9�	��CRb"����6
���˖.���D�ÁC*?��x���vW!�8�f�ٓ�����E��p�ݳP�*�R���DD�c/w
Kf�,\q٥����U�f|ڬ]���8�iS V�]������A�`��BrJ��G;��S�L����x��q.E�� �KF�;�j����GOLJ���y���ED
���/(�v󸸄���3<�s& ��>�t�z_|�N�p��:}P|B��P��<��#�$���x�^y��G�k�nn������� j6Q#�#��),�'O�裎����8�-'�K�.���:$����xꩧQ�D��vMӐ����i�Ϙw���`���8��#��DDD�ܜ� "Z�^}�`f�a������^3N���e���>o�IbRʢ�&��k��!����,$":hXB����J���V��f=�R
�v�Ė͛Z:4 %eex��G��/���4���]�u���W_nY�|n��o��B""���>j,N�xʉ�ظ�6kM3�#�=~�J�^�_�|z�8b���M&��[���������\�;�~O������s����GϞ���o����묬L��^ݎB��ޮϣ+ �}�=�x�	8+��txD��Qc�z殿�����>�L�����(z<�������]�u��xxUȰ�#dێ�ZJ�ۺUN8�$�vsh��m��㏱�c  o��v�����(��߸ 0pА�4�,Fϣ����7�k��."RVQ!�\�g1ޮ&��շ_������{���#�eDD�;�Q��ر		IHNN^n�Z���R(--��+�m�~��ƛ�׿^����oUӐ�)��S&M�{�Y3e�M����t�E��3N�̳�����ۨS ��K�UU��R���?�$��䆬jOLJYq�)����,"":�XB���������p�n�ܚ�kPPXئm) ;w��}�fa�0|D�n/�޽�_9͇}�����HgQt{� "澹�_2`FIZz'��ZUB�W��t����ILf�a�\3Y�n�{>�ҫsmW��Z<=��HgQ��UU �3�:�ŦZ��*��}��U�~y��Krr�W�k�����3g��3���0y�4�qNDD����
#G�i�Θ�P���+/UO�K�""�M�����=c�>�d �DDD-u�5��ڿ\ףS�����Qc�ɞ���.�׌Ӿg�>�q�!K��͓�o�-"��v�x���"�-DD�Nq�*��;��O��!�U۾}�n��z�*��>�>����S
��>�0�9g�9S߱s'�v�u��""���[�[3���&�%T)Z��R����󎤥wY:OLJ�8q�Q�9�  �/�t�~D=z���i��pĹC{՟�������V����G�l7����G��= |2�K����HgQ�qrj�-[�`��G#..n���(v:+;U��^���%蜞f8Q��_X��+�-�Qk��i�ҥ�[����7F��5�V�9-*Q�=��l�~{���[��qY]rdђ%!����̺���cBV�wꜱ����;�����@���������7ބ��G�>�ߡ&j��b���n�ED>������jW���P|܉���7��>�t����{ ��S��d�;ĸ]�u��M�>_�`�f�:9j̸����M<t�c?.��z�?f��g8�9Q��vƙ��UW����^���ēN�����t�������J偗R&�ֽ���xc��睏��^�]'"":r�����Y���G��ޣ׶P=�kwY�|E�������ǟ�G\�vs%)�i�Κy�$ p�uk�ϵQ��v~[�,��1�~0�r��~�?�Ou����_~%9]���jWb���{�	w��魷����|�]&"":򔔕AD���N�b��hG�t��]���{ٴe�{�	!{�k&�<􋧞y���7܈y$һKDDtd��変�\i��xC��%3N?CV�['��j1�X6;���k�������W����G��Y����}��l��\@��8d����h��<!1�s����$"�_~����#��DDDG�5k� �Sgddgǚ��OB�������Ymr�	'~4��S�}�y�:�_��M""�#ߥ� ���z�����u�׀���=����:�\ �眈��8q�46�;>#>!��s%�]���DD��nl޶-һGDD�q|�� ���g���[��f�L�>��=���~��7X�zu�w����c���7��~������̬�ו2�8��cbw�vƙ�fv���v""�����G{܈ظ��-
�J�9b���õ֦�:>�/һBDD�1=?w.�="��=z]g2[��	��"i靾0hp����b��a��""��������N8��8-)!1�悹R&;n�޻��Ǥc�;"ªv""�H[�`  ����{7[�뫫ԃt�-��w]|��h�N'�{��H���o��S�L �쎋�L%]w8�^�<uZ����GT:��N:���@$%�"%5�j����i�FU��j?5�Sv�,t��k6l�t�����1�dA�Ι8pprFf������Ė����LIM�ӳOߞv� p��wG:�DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDG���Nþ�C   xeXIfMM *                  J       R(       �i       Z       �      �    �      o�           ����   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��    IEND�B`�PK
     mdZ�����  �  /   images/6fc4b800-efc3-4a5d-827d-9566cfd108b3.png�PNG

   IHDR   d   d   p�T   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  cIDATx��]	xLW~��d�(%�J"��}�%(�Z���B��_[y~R�R[u�E[[����J����ҿZ��j��B)��'s��;��Ĉ����>���=��s�s��-�37:�PTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��AW÷&��z\I���7�)I*�Ev�Z�:d;iJ�3mtRɲ�������V�$IY6��"a[�d��$}/����~�l���99��t.��$u0Z��d�M��(��5D��a�}0�*�
��?���h��dY~�`ȫq+��L��yY���@���[���������ƍ����0��`�Aк�C��"�|<B&�������r����t�PQ:�;w'N�{˧����a)y���3�t>���ʂ
E@fB\yyP� �f�3b�1�(p�3!�<ÃY=��䫄(�d���?0��&1A3vH�JIi�	�YCd��c,�p?��0���g�Ж���lqtws���%b�G��ɒ�2d'jaxR�v�Zl߈s��S�����_C���2Js;�i���8�f�ɒM>�Q.]�����С�x�g/�5J<����зO̚=�g����f6.:6lX�t]������B��5�D��;ѽ[7���s�p�0g�,�n�=_x��(���E��~/���u{���F�m�6�2�h��!����v����;����dX�i5�7�}�����ٿ�2~޳?��#n������1p�@xV�$��u˖�Ѳe��H�zi��|��u��,�Ν'�����ԩ3�/�5PP��7o���,�_���C�޽ѵK���ǚ5k�t�:>�,^|q 4�XȺ����7!&&�+{�_�~��d��ǎ	SԥkW�o؀������A��n��B�p2�7n����Na��>$3��ARLN�G��&����~�� �����QQ��wq�������Тe+xU�ºu_ lQ������͐�լ�K�.����ԙK�.��9����(�QN4|���X�p&M|�����5�OLLDu��x�"�.Y�9o��&�l7ww7�b�rD�c�)��?��޽E��jO����[���a�0�?B��ۿr6n����o�Y�}��E�E�:uh@lAZZ*�i`5]�ر�u�9Ǻ��<s�4�V���ի۽��1�Q�n�:AƢ����D�?O�F�g:b����a� i4puuÑ�#������W��u� ̜�iL8^<H�Ȏ��ʕ+Bui������®�v�u�zS����u>l�ФΝ�P�U�@.��+��������^M�5c�L�L��S��nW",�Y��e��'""#�|���'B�B�FMТœ8���	�R��ӓC��w��t�b�_G�R׿ƛG߭~=L�6U��?���קў��ݻ[��Z���\�rLd0�q�	��o@Ey.D<kI��
2^U��~�zB�!C^65V�E�6m�W���$!-^�j� ��溃��������͂�٤������m׮j׮����{��l"��e����G�fg�AQ�%{ΫbM�6��F�흚6m"�.\@�ƍD���]P��	��g�ΕG���e?h�V��\��ӊ�����ٳq"m���`1i.�[8c:fd��Y����<P��6���׻�2�sq�{dDG2kd'j	h�͛��)2;U�jW��%�=z|j���)�b~b����!JcӁ�L��+$3�i��ߪ[�Fc�8����2�F����~~���dG��?��%\�9���ɡ���3lw[wGDD���Ç�6�V�Z8AQ?��6U_"���YԢq�0��$��_M�i������W[P��@�nns+�F*Z��@'����!����ǤI��`�<a�CI�>��p������<*T�[�Cɩ�1K�,>�>}�/�h�M�vhD�*��89�-�aq�֭�M0m�t�jQt������5k?C��M�ۻ�Mk5���Z�e����ZSVY'�����L���������'����F����g(4�Ŷ��P�^G�>|<(��p������_�R�VUDK</`9rr��WhI�6��E^��9��~��΁�ʧ(��K�c��K�^���}Ѭis<���b�s���J�efp �e
���,���5��<�5o۶oD��h���%.�sab��F��%a�ȑ4I܍��u�Ȗ-�!00�==̤?�9@���������A��"���K�T����J��2
�������r�̋h���C�Шn+���\�t	�i~`�'t�dA�����Ӄ|�'���GEDCQ��z�5{zP�gA`�@��?�h����\�h*��5���]�r^^^pbb(��1��[ޒbo�ػ^8�s4�叽|�4�@����4}�#0(h�my
?A�#����Mg�<��7��?�il���_ �2Eto�����"����j�37-N^��4g��)�8����&��'�*JBCLQ�JH�C���=d��,���}X5D�2`�����0��g窆(&Q#,���!�.o���e�TF��[���9ʲIQ�[�<l�M�V��|/="D�xOR���vG�_G�3˚��7��aj�gE��s�6��ˋk�Q'I����܊�GBEiB���j���QCG�h4Z�D�$ݢY�-R��By%�V+i�T���I|3����4����ĉؙ}���2r����)���Om�fk\]�zH�|�R�iO�l�Mۗ�I6_dْϜf4G��Fk-匷�ݥe�k�\𛍶���V���_�3���X:�-�b(ڴ#ݾ���KĤ����h$�v!VI~}��+s�^����xg��p�h4"�E@�Ӈ$^N������1���	�����ǁ=j��������o��qbZW�?��i�1��wI�t�G��v��e��^3�x޹���k+�t�w��`-;q<3��rJ�r�##���Κr$55G��޶;�a�±c_�ٿΜ�V�{J9�Ԕd��=�(B���}�\�.1�7����׭w�^v�.\�[��"{x<����̣������{�"o���]�|ҵ�"#��[v��n�ٻoޚ>�Mۢ�̛;[�A���(Ks�#�����@�V�s��I������׸��������gn�fV��8\��@�*e	%F��#�n�����8v� �2�Ǎƙ3�2+yV{<6���ܜ����#d9�¡��ȏ ""�z�ז-_�M���^nzjJ�QNk��i�܇��#��~_�Z(_��?���&��2�G9��ɡ�=�gge|�yx�fY$�Q�/R~�'������ll���<����� ~�N�z�����t
s�PVQ��<^�q�s��mOrrJ@�=�t-���K		粲24x6�;�;�%JHJJ
*�|D��-KKMN!p5�olI�x��ݺ�Ge�F��kǏ�H�"A�ռ!i\�xzz�/_�<�R�u�7�u�����U�F��K0��N�rx����̬L�(B���^b���x:y9��}���E������k��%u����QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB����Blg���    IEND�B`�PK
     mdZ�?���� �� /   images/ae82c023-d9d4-4942-aa8d-ab2ae3c53d73.png�PNG

   IHDR  �  �   ��ߊ   	pHYs  �  ��+  ��IDATx��w�$�u�2�|����n�����`a���!R�/��D]('��E�#���H(�(�D��5�`�ߝ�ٙٱ;����._���~/�U}�S(n0���hTU���2�&ϿYXXXXXX�7K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�}��/��l�v���O���A��'tB�\
(p�s�?{��N�p��z����@^��MA��1V��'���My�Y�����8��j��<&�㺉u����~ �`�tڥf3h���)�3tpX#���V�w�������y�`��%z߃ �j�T��kwe�A��styN|����݉�v���!֕J��h=������8�t:�}��y�`����{גc3���k���ͦ?P�Q(l9�N|�3�Xv��X�~�-�}�{ΐ�E���E_����ݯ�����L&��t6��[�W&c~�w�V���D,��K`	��0ީ�`;����@D �@��}����4�a��Q��@������d|�}�����u�=� yb��~�s������aǇ�}�}+�����t�{�;����W!~ܿ���qpp_!�x t�έ����ƣ{�q���sC0��N���{���sXB��+�ر�Ɋ�d�<�ө�<�O�*Vb�n��~�6��e"�|����@�J 1�vz6��y��#�o6�r>ޛD�����3���c�$��'ק��g=G�S	V�ѱ�Y�b�W��y��Γ�\�:�o�X#@��z��Žp�b�ɤ�5����Ϲl�Z<��G��\3)sV���$�� ��-�
۶mss����~
���8�V�D�z��w�9"���k��MM�$Js?�h4ۄ����B@����u�sd����.��&	]I_5^S 0��q8W��4�� :6��V��"n7�ɴ�)D��FLa��_I�������&�
)�c�vR�͑�X�h�B��T��5�Mx/�8�v�i��󱞬ݡ�\�	�,�S%�� ��-�
o��&�C�Z~D 6�/^�ط�ti�
%'�����$��J�&���l}��0�S24�V��x�]M��yH�O�7�I�:o���ti�IWaC��s�u�e�Qo��Ѽ��~y��uB���x���������1��e�^�S��w͇���-���
`	ݢ�0::�� (���5&8'6�2)D�Y���T��ik���8��k��X��0R��빬����Jrј�:������.~r����y}��>GHԧ��.Z~�!�B7�ϸ�k��&m��)/Zy�Ga��FkRb��I�X��E�r:�mh�B�L�<kL�:��̕����͠i���\�.���{��~���O��*x��L$XP(|��K��q�8�¢�a	ݢ� �j~�תն&R�g��uM���2��d���$}��qj6WM�Ԣ�sA�
S�U7�� 9=�Ԅ��;����K��浘~�fm�aj��8�$t 1x�d�ڴ�Ztz�i����{�{���W׉�ˉ�A���,,�XB��;d�������֌L�Jp�*��	�U4T~��(�XaM��EJ�I0��P�1��Z:2��%I��.C�j���h̖ߠk�A�̱��륅����J��@1���A XZ�5N;b>����&�V	0�~fO�Ұ��}�y��DZp&��{��V�ږ���=���Ծ���N��!��y�S�U����hPL�_GZ���B��e����5����3l�w���ϸ>.+���{��إ����4�[�⪀%t�>D(>r<�W�Ҏ�:��_I�Lj��|o�=y��y�ڮ�2f�EAgݩe��=�6��z�fZ2*���͠>SCO�����ܷR$��ϜS}牴�����c����T"�s�t�Nxdaq��E_a������6a�@�I"6�I�W:�~6��z�%�L�O�e��㨙�\�I��y�L庆�~]�����AS�1�ｮ�m�0R�z]���M�n&R��cZ5�u&3�׫�0�\�a�O:��>�%t����ÇQ4�5I�$�K��K�{�ٮ���ģ�lS36���)p I2�yH^��kF�����^�WMZ5x �O�y����f,A�8S0��G��Ma���k�)0�����j�W,�[�6n�2�0I�!*�I-7i�N�}����2כ&m3�m���fn7䒚t�s��z�4/i��
o�z�� �^�	S��%8�{s���	�1�L���b���2���=d!8N�}
K�}�R�BwL�Wp��!��րI���f
S�6�Q(�h���'��L�:�J&~��^�JHj�J��y�cA���$f���L�ݯs'�G���b��'�!zY:�L'f%e���*�%t��B>�g2ܤ��4���\B��gi����ܟԐMa!�}��'�H��)D��s暓dk�g�Ԏ�yMS}/S�y��l�mf0[����^�Y^5sL�\� %�@���[���K�}30ʉ5P� "߬���E�� �K��Tq3�p%�{R�OoF����ڬ�)�����f~��vS�W�5�0�#)�$�����:�Y�=�i�=�c�����h4$}O��g3'�g�Vp�Xha�ϰ�nяp�����iJǫ?A�P�ВZ�I\fڕ�J�G�HS�S�2���L��s�(�����d�m����fJ�kZ)�H�~}ՊU�u�)�hs���rYۦ�z��I���k��ΡתB��-�ߝ�>�Z��/�z[�/��u�����E?"lkn+�]ajW�XI�dPC�7��^ڥ�&�v�wl�ӕ�A@͘�L�9v2 .�='���O��z��n�=�\�i�WB6]�
�Z�k5����}��5��Ke�sGd߹�����b���XB��Ctjw'	3������g��+O�i���/IȪu+)���{	���oc�isIj�*�$��^s{w�P4h��(y�\K�{��Wб�?s,�C�Y���oaq5��E�!�i�A)�DD�f�K��MB�yAq�`��&��m�@B#Nj��f�c��^��伽�_�q�(v���An��k�e�0��}/��y0��o6o��<�4�;�9��UK�}�j�
2��9+H2�L2O�%M�I�wR[7�bj�J�@2�,y��ħ�oݧ�'���|���kKV�K�;H�j���n��\�`j���n���4oS�#�|�q�8�|���XX�,�[�%��\��Y���)Tz�y��8?�d�v�;ԏ�����s���\��;7��L[3Mٺ�x�3�����\}S�6�4�`��{U��1�
uZ �߼�$�'�yL���ߟ��p�;G���j�%t��C��<]j��e���� -E����׶�f���nf���d���)ᙑ�Ir6߯t=�޼�=�Ǜ�j��u��B��\�@�K�Q�]����H�O^�)����sӱ=���W��-,���-�
(,Cq�Z2.�W���"Ϥ_���m��U`0	�<i\���}f��Ntv�NT	]I����c J�f�[2�[��t\S�7���Ӽ��J�I��YF�߼��4:�ό�7��4��u�U�0���ёV�-�Ě�kX��Mw,,���-�
�����0�\�$ɋ��ME�饻�+�K�(�@Rm�ok�8?ʝ^\^�"�v�yLr+}���X��?OZL���RM�T!�R��s�V�>L�{&�Cy��a���z�?1[��?�����V��1�C|�" �Ѱ\8�hΔr��dE|�h�H��x�qw廤�^��'),ɼ��NL��r�>����֪i�2��UK�}�\.'O��/<i~�m��)Ԣ�͂+���L�I�:��0��^��Nj15V=�Ft��ڦk��t���do��u�͆ߥ�'�Vi����3mM��$������$)��i1�������RX����=��]��*`	ݢ� ������h��7i��Y����Nw������y�߂�$�D	���$�^�ufZ]�y�f�2h��E�����YtP7��7��4�'�l�>'���O�$o��H�73������X3���NW,�[����=ÚM�҂&��nՄ�c����=y�JQ��D����D���'5i3���k+A�f�l"c��z�W���U_?�^��u-����o
-�y�ޘ�R�sMa-���}�nkaq5��E_ap��e[�E��p���&LS�y���)��dzi�I�Z5P9��+�� ����k�R��f]w��nf�q�\�+խW��^C����j����˥�k�e���?�Yά��$yS�����K7�u��>�,���E_��f{��;�&�&I&	阝 3���M�p�Ji�:D�6���箔{�$N�)��J��N���Z�׹Yo=�G�g�t����7�L�[i��i�H
1fj�f�g�}[�r;��yOL���YX\��n�wH������yI��Ip�q�W-qڝW����Z��r;fh���ڹ��S�@PZ��L��p�.�����J�*0���L����'s���d��%s����o]�8'9�y�3e�����a��Rַ��CXB��K���gS�"m�&��0Ћ�ԗ��i6�˽	lS�79�,P��K�V��[��XL�5�j�}i2�MM����qfN{���v�����Z��I��n=7i�75�.�>�mz{����U�C��;�����q`��Fdpip[ˈ87����X:ik�N�фI�KK�2�w��U@�ք?佇�>㈤��=��|f����d�`���_��U�@Q�rǫ(�L�Kj�j��͸o9�S>��9_���9�g�W(⌂t� #.�T���O�V�x�>���w��kXB��+,//;�\&�n��������`1=���WҲ���^�q�c�ڭ��s���I��&י4�'�K�Sm�;���Z�j�7I�k֏7ה����BLK��;3��,W���8������/�¢`	ݢ��ʝ	$	D����I�O���Ju�M�p/B7}�&��2�'}��b z���[�%�s��W,Ar���a^W2ݭ����KV�3K�&�h�A�_޼~�;�Z	!I	�+0α�e,�XB��+d2!��4�$a�)S�����@���v�}���I����<W�LRF�դ��l�b�W�k�uӥ`oF��z�e�W2N�%y?LkC2��,V
������Z��g9���'XB��+��eX��!{��M-�$nӴ�̱z��u�����"�䚺���� f��&�^Z{b�����f��b$z�zz�]�馀b�t�T��ۮ���t���2�4��w��=^i��K�}h��j�d���1�;� /}�$mF��>[=�q���t���s�}�ꘫ���8VR�0���T*�E潄��9&4�ݴ"`��iu9��M���^Z30����t�V"uK�W,�[���ti��P�r��I�+������i��`��_/�r� ����6��X��\��d�x��J���$�꘽�{լW�H
�1Ɍ��1�T��a��dݖ�-�XB��?J���q��<�L��N!�d�\�z�k��u���I֦��js��CۖV�2�+�!`��6o��t�N�J������aV"� lI!ڣ����en(�N[~��S�H	���"f\Z��qh���V��+������f��g�U��|NJ�������u�J�-ʈ���S$/�Jl[t��k���c�(`�q��?�O��ZG��UK�}�t:%�sdm�I�h�	�t��"�Zq�Y�I! '�O+�u�x����)Z�f���^�����lt�Wa�3���m||}֝8}N�	�s෰TE�W�O�֠~�Z��Պ�-;·����l���0s�3�N�i��抇QP����n��F�V�5�=�J�B�?�P�B�T/��P�V�B!UKU�R}уHi�j�I{����U��)2}����E�-��R�
A���>��������|^ڍםY \Yz�cl�,�e��XX�+,�[�2�l�Je���)��K���V�&Ȕ��n����-�f���^���d"��L�J�}���z č�i�5u����MEm��af6��������Io����8|"-^k£xKT`^.�)�I����*	9�J%*�Ã���@��Dk׌���{�J��o�W_}�^x�-:p|�Za��l�R|]A|ߵ�k�Ր�X1gy�D���Ѓ���D���:z
f�4�B:����D�����E��ܨC�r�l	�⪀%t��B�\��Z����U��cvbӺ���B�j�u�v�6 f�<#͜��nD�EQL�ql��q���
��N5�P��Hg�5\���P�O�6F�D��"y����J����4�� �c�Gb� Y��:�-���ȴ����NJ�\*S._�|�z��c6h�5�������ߣ|�.��0��`�@�c�#\�,x��W�b�_�i5=���ߜ�5#c���_�1��[4<R�K�T�\�[+�.�)h�`�`���,,�XB��+3��Z����^C�p��>�	�r2M�$#ֻ�źs�M����������
�Z��]]�!(ཎ���^�\��n�%�D�a��f���t_L�Yָ;�p�O�:��ځ������ƨ֨�u4��m|�R�JK�
��hv�D˵���g
��]&��3,8��\s�V���C�Y/���T�A�p%�^�
E
�)��X��P�f�zT�=���������mh�E���E_Q�Z�K�*P�)��D$�|����р�(����G��u7�͎��˂�(]l�Ƌ�EWG� W�{"C����FW�N���f�K�����Q�������T�\k+luڸR�޹#�	���@��t���0��!l�����Hí�ᫎ���^�U��ȧa�Vå}���y����i�oҁ�g��=*�D�g�L�͆��QCn|���c��0E����n��~�����4::Fs�x% ����ɨ�熱��F�� ��Ld����sXB��"@.8Q;I�ڥӍC;���N����vF�X����ir�2��'��j�3�'���h*��ł�ܡ�5�f(�j&2QÇ�iEѪY+�&+�%���p*�
�t��f��ٱ�Q�Q�xM"���ic�<p%zm�\GD�:,푲�lϏWD�gXcF�X
AcL� T�����h�"�Ʃf�:�>4F�=�w���iZ^�g��јCLʭ����Wޒ�JerÔ����\��C�R���礩R�Q&�s�Y���_��S���Sgg(�_�c7��"�Ǔ����n$lx�}���D���5[��S.�p���J��,���w�K5��[g����\��������fɩ�h���9�5��?H,��X	�t:8��pj�#�����Vgf&�;wR�q+LX��K��0����ݻy���������|advv6�{Y�ó6�l�����PK�-U�ײL�^~�X�	wa~>�R�L&�+�l�^O�Ŵ�h��a3�O�S-V�s-r!kh.�@֓��s���2?�'��`
�2�����(�y�n@F�j������ips5�- �(�L�C;�K�v��E�eQiV���=Z2h�ȝD����mȐ|R�S��%-4C�����{PEǴ�hӑ����|��U�4���Uن�8```@�aqq^�g�)>�M���L���]/G��\wD{wιB�ѽE*_4���0��/0��dm33s��!Uj.�8���3O�C�X8qe칅<�G�֮�E>BY��N�I��v�����^}�����˭R��e��=�
�T�Qw�0pW�s����ń�.//�f3�T+Ԫ���e�l:I0l�e���7�h�Z�l�a��[�u˖����<�o�㖟�?}���7Α���%t�_�DR_��W?���/gg�o*����`���<�V:l�j��j3�fD�*0I�X\51^s�5t�ܔ35s֩T*��/:͖�A�R?-ϑ������@�F�F��o4kN�Q�/�N19��Q��Q7ަ���du�dP�%�zR��Z����Ȫ��W[V=Ό�שּׂ=Cl�oɵi#�N�t���N{b.���(��IQ�h}�l�5��D�C3�g�EU�"|*]���q~C�%��Z-S:���%r�1�W�5�K��-&v����han�i�.��;����04�������|�D�BN���y��)�gs���S��S�8 [��N��=i�`�aÆ���ݻ~�;{�ԩ����D�O粴��D�LZ~K.\!�-��$� ��B*��w������8i1�|?��gY(��-�n�k�mEv>�[�N���ۻ�9�C����>����{�}�j�W��-.�J�����_�����o7m^�%�Ĳ���޻����˃�Vk��Ç��7ަsS(�C؊���hhp�>��Oҷ��=�8;G���/��Ç�<�����ݷ���=x���?���q�ںu����QYfBt�/
����5/*��o6�`��NLL�g>�iڴa�U�Z��]��뻄��������5��{U�&
.��4�]�4�j�u
�t���q-�q�U�U�?44$D�F�x��Tg��TH0��}]p%���ۣX&f���^K9�A���+�^�㮑�Qt4nl� Yz�=Ք�sI�k�9-:�,QA��!t\�8Co��=�܋b����L�% ��q]�ˋ4�����͛��:S,�s&�Eڽ�M*��Ԭ7dm��ħ������w��G���y�ۿ�=��s|^��[5F��y�q�t�M�Ҫ������7Y�*��~�T)��_�����|�����
���e���������'�x��䲙�L���u'�����h=(R��r���M�������h=!knkdЌ�]s��`��y�c�c�.:x� ���˃��B�A:��r+�uW$0,�Ͳ�U&�Ə?�]>�B�9�0�TE���C}��m�F�'��n�i'��_��K2܌x凌���j{��O(�+��Jј��۩t����Jh���D{Ǖ��C����I�yt�qp žy�\(��Q�$�u�S� ���(y�D��$�>{S�ǝ���^�!���2��B9;���v*��G�����ٟ��-�*�**��Pe��$��[n�����ru�,7D-�q�`�;�w;���,|�ŗ��ޓ�>�K�L~�C�g�^:{�<�v�&V��;n��>��O�\���Q�Q���>�ڵk=�ܳk�;�|��?8s���ƿ�Y�����nqY8y��-_���y�s6��ڝ��M���g��x?TG��ZPah�Z��z�-4:2D����^}}��0Cc<z��<<?���S�\eMr����@;v�$��3�����<�����ӧ�+_�
;v��l�@�K�L�e~���􅳔�2��K�3���C��(�S��n�k�X|��QE.Y����&���
��Dn�µЋ�bf����+���U�� b��I���j��~�+h��#�x�D�~�|�v��|\��k�s6^u^���D@�5@�5�k�fs7R�d<�7@�a��zT/.�C�����8��h�>�9��������o�[L�c��#��)��_�_�JR����!�n~v���[ߤY���B9ֺ�h���q�]�];I>k���~���o�����|?�bá�z�F��|x��b�|rr�F�
�?7z�������뮻Nι8u��1A��Y���V�O��o�C�?��/�ȗ�"YX\XB�����?���W�U6��n���GŔ��ˬ���k6��Ke�"���8�{�t��?qQ��a����!�r�z���l�fm�:�����C3~�=tp�>~̷(�"�j���}�O��H�ť}��ߣ%�Ρ��� !d��� &�������!�]N��.^R>���;Z��sz���i$}L�N\n�UK���H�zܰ�#Iq��s㠳N�}5�������\�5棂4��;7��S�}*�SZʮƝ�P�i��y��H?G�X�HQ����]���@J�j�_*T�A�O,��_`���v��X�r�5��C�}��ͤ�BX6%���2�o��*�*U^kF=�A����{$�vn�FG�i�I�|��w9�2z���k���S�������i��8U��|�g������-�h�����j�Ž�e�ڳg�Щ��7�%t�+K��w~a~�5�T�Y��۶�y<oϞ9Os�%��k��)��-P�	iͺ49���ZXb�g! ��_z�&&����,����>�0]�փ�������O���'�_�":�.��?�ڼa���Fu���{�~�W?K3����=.F�ZgͿ��K�+K��&@d��L��mT��T+��Z�s����(֢eH]-��&�N~{;-�h�jZ�m�N��Nnz`��ŏtJ��K�2���t��9�ɵ��VJ�cAC2��H�v�ֳ6�H�	�4���AT//Z�A} �����?=��E�OE5[���}\wމ��E�zq�G��v�S!��5k&Ă��ذ��7nZO����X8ˊV��Ǟ��Y��>��Gi����_�2����������{���a!a`�Ν4}a�^~�Uq��Y�\3N�6��B�s���*��
y!�j���c�bt���;�����N�<}-YX\!XB��,d�A�p�V49�Z�_M۽g/�izf��߸�Xk�h�+��ã��)�3��r�
�"���Y/���گ�>�OБ#G�'O��.^�(5$�UJK44X��w�Z�2�>q����x��5�5I-C�q��`F���
�g2XM� ��t��>C�Er����/���+���۝h���&}�S��oF�'�# N3p��n
,�@�s�~|V�]4�0�J���"_|�.vH'#�W {?N���	5\^|���#�#�-pR���;Q���b7�fw���[�{^B1���
��D@��w,8����#�<Ĥ��V�^M��������&�Q�C>���5����+L�ȴ��ߪ���wA��8���0/YUG���M��c�{�Mڰi3i���q!���XK����'>��o��;ＳI�`XB��8L�^ݯ�p~����4����H^����j:q�I�e������(�?}�ff�X;_�i��(&����ߣ]�n�����ǿ�=���t���={���̌P�ǆ�}qq1�o�|ʤ������b����<���ùV�R��#�G����j��ٺS�M���� &K�M�H<*�ڹAȏ6{|���9�c:R�NsӐv%��n��Ea�c�y�hpD�k��(�k����t��.Ĺ�@*�}��*�Ǯ�hR^�]��5��ڰG��q���^ؔ���[AJ����5E���@�X�`���T��,���}.����]w�6���� _�"a�#��S�@���D�j�����o�a�b.u�)7��N�?�<MOO�w��g��jV����m�x������歛�ο��𨔞��F����X(��b,�[��a	��r��H*�ɤ��a�\\\�%kRn]����o���h��u�����Kn��)B�ޏh�]7G�p���i!�\.Kֶ�Q�Y�.��\�.��
�*�9-:�,�49���_��s���������Y&��Z���;�hJ��a��p����'��JQ'�V�a���U�5S�L��m�6����tk�:>`j�浙Z}Tƶ�ϸyMf�^�|������y�%�,1��TA�7ڙzq�3���FCo��iA���q��
�BC���r�"h�ș�}�X?N$Dէ�v9�.@xy�j0�Zx����������f�I)�@���Ay�Z�*�T�[^*��=I/�D��̧D �����'��O��x��yI��K���z��H�#E	�k����_����ΑQ��AD�#���n*5��]����������VKLLn�����Ҧ�[�Y��'
�H@?�.^��B2p��:s�^۽�j�
���K�� �k��=�Z�n=���!?����+/��}O�x����KD<L��st�軴qӇhna�G�i��[�!;L�|��(D�q����\�j����!���:��N�Q�? �̀2�L����bQ���A�J�~���6���l �  �&k�n[����x��<"�V�%�ZjǤ�ׄ��K�hPՋk�C���+`օW�@�-�����t,�(`N4�x�������(�)���X��m+���R���6�F�~"H��ި�b�H-M�	9�u�y��Gr$�Eoh��B��p���%*�x�t�}GKL���7R��=��T����c���� �ѱ!j��;t� :�.-�i`x��Yh=r�(��{�n޹�ҙ�r�Mt��ד�ɓ���t6*���tgN�����4<>�F|[\������ }�̅��� �����EZ�Zs�0?؊��5X�L����G�й�)��":Ҏ��\�����/��بhF�3������%-�ԅ�%�����OĜ�;"φX���2�+t�u���Ҳ �6�f���ԕ�l�\��U�k73q�+ZG�6���u*���Y��v����њ������L����;C��v���|���k���\�Kݯ0-m~#Q�q�^wg�-�E�s���y�8XωL�QZ]��RD�5�q�h{�`a�Z�ڨ�'��/./���b/�Tw��qZ3����RL�Y&�\#2&J�������|\U/-�Ňze��@N�U�� �w����7ߤ?��?����!=���i������c4W������|9�<_W�K�`���oұc'����䚍�b6둅��%t�ˁ�Tj�o� �Ӌ��K/��r���:�$����iqa��ܳ��.�H5�lf��&?�Y�	tp4Gy��,E��3���o�IkV���jZZ*��e֐�D�?�O�^GY~����8B��~����\~@�Eg�>eͺ�KS�8��9��_�7�BSr35֨tjK�H㾴�j�&�'��a��@�8�^� z��o�~U?=���f���J�/�'o��5�O] ���ܟ��L�ױM�4�I�����y�%��M.�rw�.�v�~�f�)"S-��`V�B.G9�N;J����4><A�����iav����_b����>Agϝ�7��w�yGb3�x�	Z�jU�KT*-��ci�7�z���P�{n~����O鞻o����(M��S.�%e����O?K_�җh�5�K����ykn��b��nqY(�S�Ԑ|m�.�����w%O;@����ť
k�5~��)�
J���$�/��昨���O�{�?AϿ��<�gYs�,���G%b��AP��͛7�>�j������{��s���j~��x��u(3�E~�CQ��!�9�qw
����Y�!�n��ܮ��ĪdMv�oj�Jت�*�����?S�0k�����rş
"��c�<�w�����v�w���5�N�����։��<�fԒO���Q�zJ��-f)��2"/�`����L����T,��ԉ����O���sHS�s�GUC�*���ɓ"��_����.),��kX���p͠ ,;��!`�����[X��ﾃ����^{�mB����oӳO?%��쀜;2<�6j5��[\XB��,�M/�*g)��d�e�D{�6Y.W��K6�c�J>0JgJ%�zI��a�_D:D�������}�8@��� k���*��U���v�9�����4>4F��������>A7�x��� ���s~��	�n��T^�*k  Dg7�N�SC�?M���XK�cU�N��e�A7S�T��t^ՔM�TI�$^@ק�����?�j�f�_����յ@�2�Y��ټ~��c�V����JۓA�f|�nBפ�)k(�vʦ"w���0kη3����|U*�yg�MASoI&,<�y҅e��۷�Ν;��k��4��[�I���7閛o��o��^x�%:��ij�>��I�{s����[��>��������>*�	���3��7_M�����\�����nq9pʵ����tAc-�^�֋6�.--.	A��Y,���d��$�P�֨H�mDIW�ZbM禛n�����=�Kj9s��L��}o%��^���w���Z*f|)f��I�g#2x�7�����w�:d��%Q��"nq��^}o���ҝ��h3�]�G%t3^��$�9?W(��:��c��Uc7���@�K[�y��9�x]�I��i�4y�>��M�B��k\>f�8=6ſ�g��Gz���ׇp�V�J�����7�=�8�Nж5�d�w�c������4;v^��y�ݴc�.z���rƄ`�9a~G�·�~��G�h-�ޖ��Z��*�\�m�M!P�w��K:ύ�,̣]+���S��F�f	������ ��f��M�F��%��Ղ���|.�J�Z���>{�5�j�$>�@����T�'�|���o��hHo��:?~�6m�D����<T׭�������t��Yj�pL#������n��.ҩS�����t��m��d�噶��1h���'|�(�ˌk�t��L�6I��6S���J�R�<&�������@&:�j�*$$S�ig��6�h�H�dCRy\-b���/���q��՜K	zK��D��ս�׉�@�Ѽ�5�;�j:iu���tM$c�(���I��D�T�tu��(��rs��/�G>�(��y*U�S��W�H��Eɜ���.����򒔃E5B�֟~�iz����W��Ⱥ�=h�R�h��$-.�Q>���4�;�Q�_ST��PXf���i��i�P�����K���r���f��?�
�<!��Zm�$�F��(0�7#?6?�)��j��ޥ�j�F�/�?���?���\��ڨ�m�R�0N���:M��H�^���MN��\���A!{�ߕ�83	y=h�)I���X�M�֓�x@�H��S;6���sӇ׈W+�F�d��e��a�+�w6�&�(H�ى���4JQ� /lG��K�Լ��c���v�w �A�Z��5XOץ�xd.`.�R��@@P��N:���8��M�o�{���
�܍�Gz"\n:N���b��$�:���A&f�{���c�������~�Q���3�o|C*���� �w�&2)�kKT��k؊�ԛ���7C|�Աu�p``�,,�,�[\�t�s�ߜ�����/�F�N��9��J���P�8 Z�~QTU�2�䙤�9L�z���!�:�u&X͛(\���%k~y~@S�lzf��� 06:�дDʧ2i��Y����H3OE�A�ބL6�A�Z� ���I� �B4�.�	���y��ZA�J� �7J��4�q��	!E�����:��<����"�A�v�F�ϝ;'D��@4�V#pD���U�5������/�q�et�=66&���־�~s#�{�ڵm�u����h�؎�D;[��d�ǅ� �m�و
������̸��d�A;�I�ZC��!j�[b�q(*��Nli����ђ������-��Q�M�@Θ5	�z�����J����\+� ���K���:��XM�c#�,�����a�rr�e���@��*��UT͑�A���?jǚ�-�,�[\�V���C1ۦ��*���L ~`��B����9y�#��4hphH���Yj^A[���S��pP$��Q?�=�V6:s�>e>�J��L��ǩ�l	��P�̉�n��D]�🙶%ד����0���)aj�N�x�	Z��	�*�$-O�zzZ�� Q*]���2D�si=55%�A ��8-ca����T����ܸ�07��5a�J��hq� b�T��c��:u�|iÊ��>����Y>k���z�F��ɀC5�'�Z;L�)�]��޸����a���~�xO�/y���D����o5
D�C�y&�3g�IC*�u�t�
�'Ȣ�h}�kb|�D�#���io@R��>��2��|���NU(��r�a��~��W#ԪלFʳ�nqE`	����='�af̗��&��TC�(�_+ʬ-�g��͖�ة��c3�ѡq��Qʨ���gL��:�hA
hԂҚ p����L�\���OKO�ŅY�[UZX���N��w]��ב��x��U|�N�J����,f���)A�I��krE��� a��2�k��3�L����眅v;P��Ql���=^�ԥ�InkA*n��?�a>�h�<>��PFB��&˿�X�d�&v@��T�Q��A�P��0�G��p�0?����l�f e��@�Pī����c���[9;Qe:���j���9Z3���p7�� ��*�6�d�������ȉ@�, ]*�a>M^�y���f<����s5J�4�j-�_��V���:��Ei�[a�gق����|�5��nqE`	���X�E�O�����kV���~ ���^�6hfv�*���F4<��.ʀBkG��t���T�7��s�hQ�ҍ�m�`.���Ξ��'�={߈}�q�r��Nd�ad�w"���|�hC����L�e�`s)�i7Hfp��uJ�І�E���8l�x 5]�O��j׾���\�,������A@J�.�8؇��t��bN���|-�P��=qC��~# ���5��>�|����{�-0���A]Q���fLI�us�̵����0�[o�A�Px�&��'��,���O��@�
����
W����Y�� 7@Y�m[�R>�e��<mݲI�ɞ;{��:�{�=416B��N�!��I��R�AS���w�����+�Hi�L��|�ZB��"��nq��a�dL-�C���m��o�Nk׮���k����1Gg�]��}��x�mr򞔇-H-�r���ڲek[+s��[�J� ��w�#-]��ffifz���g�'��cߣ�'�������[��v�����r�)�r������2�$u]��_a��i����A�0���N����Y&΋g�T-��`����6�����p�q�@dW�Uv�1j��l��x/�&��T0��pm 
�b��64{�?�y\�~xh�H�i��a+�\%�F�@] �R��9
��v����W�y�5n������6�K��,��R�����4u�<]<�B>w�,=��3K����ܢ��M�
,X6�-�� ���K��)�����k�;��X^Z���c��~ ~�jy��n^ς�(ҺM�%�"��"����i��h��j��^۽O���	�����/��-.(��6��26�_G�����k�F���t��������}���kߢ��T(HC�Rm����v�Z�0�!:s�Ů��襗^�`&�亵�jb5eL��)�������f�y����O=B�Z��8L�N<.9�R|5�Z�Jz}I'�D*��ǭ�ps���G�ڦFʃ�����-U��h4;� ��B ��ASq����G�Ž�`<��#]��J��G��k��\��1>ǂ��'�F�s�.Y��A��g�e���5�j��=��0�[Ҁ4UH���=ւ��K#�;Y�J}�I�s�/��, ��,4�<��������O��o�7���˥�T���	*��Wb�ugffN�;o��~��TZ\����Ī���3��*ּ|�A����|?.�y}��t��Qz�чYx�#Gܸc��AӧM7\O��ۿM'��UX��-�[\1XB��,��ړ6�c���|��%���1�X����J��ŧx'k>��[�A�g�����qǪ�IIW{ꩧi�����O~�^�)D���,~���"�D���?7S���I�|^_g�E���6m��[n�I��O���-I�#R�OjJ�I�F{ϰC&f�RӏnV@��r�|����g�-�F��6h��Î�a;7[���A�J����@z�m�#����T�q��u=��q���! ��p.��8>dh���T��k��-�o[��+�;�\��5��L+�����������{k��;�a����${��e�,HF�wO�Q�@��ч?� e�<�w�,m�ϨP�֮R��0�m!��ý��;����sld5}��_��?�Q��_�R~����/�0B�ëijvA������[��i�P$�5�ֻ�{ﾇ��ē�d����[\)XB��,�~#@��T� f�뮻��P��	f�]�yW�!�?�SL>6��>p?��o?J��6
b9@��v"@�
A�m�-c,J.���j������>�0?�ΈFU(f�_���~ݒ��3��bM@Z
�:A�Љj�JJx����daw59�L���n5��XA� ��; ������&@��Zs]�� lc�
x�ڹ��q�@�8�4j|/�z�{ Q�0�C��ZtM��@7��������CP�!@hl���Ƽ��콶��,/�ף�Lw���	ݗ�Jt]C �7��T)U��/��mظ���/�kHf�\Y��G������Q��ځ{X'~{�j<��gŢ�,h�t��i�p�>��l�W�"=� �a�&Z31��E���y�vA~���(��W���;�S����tϿK�W��-.�ۅO;�j����p�a���;y����8��a���i~(�u���7�l��y���K�=K�s��e��wv�&�?$���#D1>2*�#C�Tbr+�1�j����'z�]�b>C�����\������S������P���u@��X�C�<�5�ڌ�6K���u�C��~5�G)_n;X�
�D>�����|��LJ��&'W�M�����NS��#�t�*U� P+#�e���9���j; �0bR�3H�a���"�]5��S���Z���q�q� n�^��0&���@����v+VM�����oetz��v��YS�\7�T��ϑo4ɑ�y5��j���'U�a�r�]��8ZAnUP�J��9���^3A�֮�����ݽ����>�c�:���������]���֭��k@ϝ��o�E��:�o=�m�|=}�#S�筣�L��]K��"F�EK�W��-.���M?d�7*��o�;IN��~�cZ̈́�<u������r�J�ũ!�|~��e��i��7� �ѣG%5m`t�����.^8O�s����5{����ڠ���;?M�cC�/S˯K[SO��衝��{��}�ș����؜lV�k_���,5W�� m5f�5�fv�ݮUڎ9��gMV�i���,�6@	O�X��j� t)��s?�� [	*�ׅlUyC�W�Z�~���ڵƹ��5� �jAP6֤�5>k����jzZϴ��=�֫Do���:������F8�ʆ
���'L�0����R�X�_�T���Ւ�x��)p��6:q�\?���5kh�����7_�u�ޭ�\E��O���G�Ϝ�\6ł�z��2EI�sR�D�� N$�8����2��nq9�0��>�úh4s3Ӕ�f��i~n�����W�v��H�=.��{���{N����;?po��vz�#QU�� �l�N�<A�����4xߪ�	�������THj��{龻��kT]�r{�R���(&�$ȇ響���*�'��-G��VJ�J�J� *(H�y���Ą�𑛕��͠)s:�Lˁ�X�y�puΤY۬O/y���k���OS��":j	��e��v-���ɼ}�,�+��ldd2�.���G�q(��tM��dHd�iO���j�s3�4;=G�rC�06�+�y���O���&��^x�9jv��N���"��5"�$�mh(GC������X0am��p�dYhh6+b�A/��:�l��ŕ�%t��B%Y����A��C�R�jҵ�ma���C٣ֈ	�a ���4�Q6����T�:�Ľ�����7�1ڪ´>5}A4*͡_�J�������5�Il�|��!�f]W��)I8����x�Bk��m��SWR2���6�dj�i7����?��>-���m�u�p�����M��W�h{\�V�L�V���L.۾^5�kKU��לs��߁��ֺ�f�{uAh�\�oj�0�c�9�ɪrz�B�fTX'��a����rÕJY*��9�=���Ϻ�&f�q�֭_O�B���c�i�:�A�/������<���iB*杓 �y&s�\�����}��>x��ZIA\@t��*);\��(ǯ�������8�?�^�y�W��-.!���-��=�p�"�~�ڤ��"?<S�.�6<X@TuY���/��>!�a�ggh`hLH���)����h��v��Z\��k0��S��|���.��C�i���X�g�@�s�Q�V3�������v�Ͱ��	C5Z��}�g���kf[O���������[�ӂ1J�z������4`ѹ�R��6A*�뼺~�P���qJ��5JT;k�:�j�07��R�M6�QAF��,��^�������"���%����ϝ?E?���Ig��>D���,d�0�T*-{��v1���[XZ��������F�~�3�,�4���
�Kљ������m�l�M[�Q~p��<VynAH��{�ї��Uq	�Z=B~˵ڹ��%t��B.����`N|�G��'����LHn0�����f����Nh���rl�T%�3��v��@w�q����K:}�,}�_�Gy�����~���Lsm"D!2����9:��~*//҉��ӻ�f-~��9�̜X�4R� ��҇�'JBJ(&�i'3���\͈�6��A�2�R�v-{��ƫ��U��:U�4��j%�>��5�P��V�3�T+٩6�&6*��Ĭ�T�f��ݠ�ٙN��o��Bh�>����V��R��1�G��:�n�4�G��ƂD���ر�t���t͍7�Λn��3�,���_�N?E�\A��B�K�B��z�6	�3ʝw��g����e�R����G���Sg���i�Y��3�ghͺM�~�VB~�=����<L7n�L��l�,,�,�[\�t*̡�K&E��(Uʋt�0k��52$���k9>�=3EKK%r�R!Ҋ
Ei��t��{,�&�=��o��vj�:��P$��������@���?��?��2���@7��ɚI��D�ݔ�W�Z�ҭ�:Z��+LӹYM.�+����T�ǘ�]�ES�9�i���ꀮI���J�:��6�s�pH��Û�f�5@����(���>j�[�b1�=�*8��L�[����9ӭ���s��"s7|t:�Ha��^qh�Y;A'O�����j� ��A~��%��J :��ZPX�RZ���Y:r�yL�CC#r/~���s?MK��~/�f�;�����ȱA��cg@���\%?D	ڷi͚��v�F���%8ך�-�,�[\�AC*���$ZD�܉���S347��O�:/��+�:kDc��f�R#Ҭ���i�y(0S*W蕗_�W_y���,�2��V�i~|{���r�e�yRK:���˴cǍ����o�C�N/�������471Ӻ(V�J�VikI�&Uͫ�4[	�]�5y�Шn����怦�Z���k�9�'nV�ӆ)J�j���7���樫`���y���ZLBo�Ꙅ-�E`L��G�m�{���G�7��Y]	����Jz��c,M�S��4�K�b�M��K��w�}7}��XGN��<'��V+�4�����bA�_z��bxp@����-,�.�K	Y�I��D[MH�N]��jm�̖�iN�ފ;�W1�Wh|<z�;;eM�W��-.��v3�Ji$��VA
~��S���d�
��Rn����Ayx�3^�i�5p���Jb19(,S��Y=d�
�먴���(>NM�Z5:H�l�D�X+CT�7��5z����=!����FZ9��T3����oZ��a�V2Өm�L�7"A�ۡYc�kQL�МAjp5�@� :́kX�ł�Ħ&t��!L���	փhl)��k�l?t�́�i@� �k�Z4?��k�mWn���j�܎f�k��B��@l(J��(�1�U*���P��D�z���6$����nk��a�o�!��q�tmS��8��L�?q3 =��ãm���:\wq�(������)����±���ޢt� �3�?��~E���؂T��� �2����x��{4�.�p�,,��	�w��?!���>\�]�q��nq�`	��P���VMM��� �W���7�I�S����LL��z���8
�t�J�=i�(�&J��>kU)j�q9Ҍ�Z���m�y�[�_��I��G��g���ޒ�ѕ-��&1â&����a�w��(��+H�Asz<��ig4G�� ;h� q�F��xt@���^���A�C���65_c-*ས�i�=lG����b2 �믿^�}������8�����W\���=!kT�{g��v�2�6Ղ��o���Ր���!��Q�Ns�a�Fj�j�X/����XG�]P��ZF�"(��U� �7��dh�+ҧ>������Q���Q�D����?��,���Z���i�8 Č@�k��fM�N]8����� 0:A_�S�EZZ���6G�`)I;n�V���2��nq9pJ�E�٪3�c��+AO��e���.�������Zk٥%֦KT���\Y�q�)1a"�=�Ht<:�As,2���}�v����O=��>+���	�@���!rR^L~~T��Sm$�&o�<��S�9A�V�7֏B/hJ"u�y;��Z.���F�s���;w
Qj�t����j*W39̿خ)e �� dmӪ٠c�Y��0���\��� ym�o߾vԻ
X�
50��:!L`-����Z������k�=�ڱ>3E��x��uaM�>��u�b>�W�U���^�(���>�~3 /���S:��X��k�;�q�@긞��X���Y?��5I]k֣�>D薗�J�bz��� �Ш�4p���t�a���؀�Nb���/��-.��8�Y-�JMʬ��y1�%W������Z}�&�ի&����� vRQ1�N��ÜJ{L	6���@����.=��T�B�oP��xH#�	������ԝ��=f��܌�ƫvR3�TۡjG4̩����5�\���?҆6��7HS΀<p<�h���p��õ'���A, S�w��@�IA#��0���b)��p��C�W�-�}�Av�
�q��z�5��}hyX-^a �n-=������=ý��m�*�l�sDeg�m�J�7S[��ie�P,<�]-�jTp��e��G�V|p�T�45=E��%vׅ�������v�tj�r�ynn&"�'�y��+�{T�z�"��"� �2�K�����ϝ���Mkaq`	��rf3� ���ԯ7(�e(�� ��يs�s�e�N�Q�K|�yt[.EiWu&M�	OKe-T`�����b���V��fMxl|"����СF�I��}br�F���%���ȡX�t5�}��ԗ7+�)��Q��eL5{��j��󎘒�l�B�7l2��q�|aI�(�DM	I+!�O#�A�Ђ�>:��8�w�Y�� _�	��1 V ����~Y���1��QA@��U�6۰�� D,�mFq}���\?������!ta��������
0؎���p�l�d���;�[�.�v�K��-|ϑfL:�e������xL�˕�\����]���y����@�L6O�f�*s5�f:�G����-���-Q���k�Ã!�:�[X��%�sb�Z� +V*�8�Ҭ5�[\XB��<�|֩=�,��-��Bl��.Q&���ay�H���<?TYE���&�x����Ai��mq�F�6�˃�R�Iz��ML�w���z|O�{����?BǏ��#��VщS�������ж�ү��7z�fW3=��íU�T[�A{��)O U�����V�ѐA8^���Xq��Kƹ�r��� Z�v��{=����\4- yb=�����5 �hx��CH@y]uC@[׊y*d`N������u�ݻ7n5��8B�^��z1�F΃�!X`��b�;�x��c��N��1�M-*L�i�F�ߝY{�y.W�1�������hb5:�-��h�����ߒҷ舶a�&t���o����JK�|�}�Ek��ťYZ31)�t|�^�uӵ��{"�LL��S'�ҋ/�Lo��UYXE/�ln@\@W
��-.i/�_�ү�A��W�Ѻ��Yc]ÚtdF*ϱ�NҾ�(���R�.~uԿ��3� F�w�����n��&��^{�5:y�x��y7�&���)��_��^}����~`��m��T�2�P��3ڦ��Xة߮~t�N5�J{xk5���OM� 1�!�����YM� U<����4�P3�F�ئ��Ad �(�)�kBۧ����؏��G��o���:@P'N�'�	"�g�a>��B����{F�u]g��r���� f 3�,��g{�3۲G~�=�c�zoyyf����i4��%Y�5%���H1@�ȡ�:wu�������/h�������]U��{���m�7��p����1~0>��x�
�yC��a>��1����x=���<�_[���؏���
����WߐB�!���5r��{F������{$��Y�~�u.�t��
@ٛ��r��1����6g��Ћ{6v�O6oZ/7ݼJzz���d�9Y�f��F�����ߨ�^�����x(�Ē@Y 	 =��}��6�\&%����Z�T����5�e���j�$�vJ�0,�8n�>/����8yZ�z-�n�L�,�i�,W  a���k2|��Z�M�-�d�҈m�ss�����%��?��n�enZ�@7��iɤ���w�QL{>kIT�J���O�B���-x ��HaQ��� �q<,b?:c�8�mT���qt��`�ê�2^�Lp\k�� �� �x3�`Ȓ.$�a��F���kIx�7]�q�q�9"k׮��t@�A���((��c�V����3��7 󇲀yc>�s�3y�Ix,q�' c:w|��t�໭꺀�?d~d���ZU�o �ݿH����}��N���Ke��Z�i��`=O�:&��.�����e߃U�-Y��7�~ʵ�����&}�yY����Mal�L�D�c|ܚ����ӑͥ#�n��  z 7"���c�!�bHDK+`-��W7ָ�Q�-��ͷ�*����;����c#j�'�@?Rm6䓟���~�!k��M������铧�i��;���j��Ւ�N������wQ>���䳿��5f���Q�/��H]��G�s�6�P�%���pOs�S�����t,`�2��x �� 4 {�8�:���}�k�=W�6�d��1q�J�o�}��	[x2��q.Y��j�y�`,($��� ~�-�� �
l59��{6v����=�n�]�9p�P���g��kbܸ7�5�T�j�wIE��x(�����'�W�$�u�|�-�$F��3T/�$�M���-j9o��n��Cr��ai5U�ץ�Dc]�I�}�z����m��f�������/��ݻ���9L�]��>7s�Y��ee��AY��_�z:�83�ٴq@��تKT�t߮j���u.�I �܈��h�bc[������%C�A��$��k�����+�m�WR-�n��&���'��ذϟ�`�NLM˥+W�.��
v.��X��1���VT�����m9�ǫ�t��(0p�����%.��F�r��g&�o���d�lȊ �;�����LI�1���>�����u`�B�ą9aL�;�.g΁ӵ���̝D,�����b�Z� [ 9�Ͼ���91�৪�S�����-R��������<�~�<R�r,�^��� !OD�1U8�^5B�Q3R��n�*�rSj���w�]�<Yn�������i�ve�`ӫ��:��x���b	���>����MOMH�<'�|F+�o�}��\o4��Lܼ�&�*X���l�B�}��e�&yg�>I�s��TK	d$ �@nHԊj[[�Hȸ�S��Y��v�:��<kVؑ#�$��I:�77������v;$_���dz�h	I���ߖ�}�s�A�g��w��׍��ʞz�r��I��ްf���o��*!�xaX^~����;��V�r��%�)��BT;�i4e�Gbr��]�~��N�����y��OK�#�@����Ke-�?���8��e&�Y�g	�=�1vk�X�����R�F�rB��{����f]=�_��gC�X�Z ���[��dcQ�y��k��1�����ll]o�����r
g?�*� JW�=K��-˷���Y������I�'N���B�fJ�{a�U���ܼVR��?����MYkU|���\�T�ɤ#�N�F:s����eb� �p\z�ݺ>I��j�/�g������@dA$ �@nHb��'�1�eŦ�z�J�hԞp#6����� �b�ڡ&�$�K� 6�3u����~����,f�?{N��OI<��.���{g����EK��=��#�X�2�K�)�F�$ �V��Ao4��}�a��u���Bv@c{M��!(�rn�k��3��{�{E�P�k
C�f'ر�8A�.�LK�O��gR㘘k�	��f�cl 8��������@���Z��7���M��̇2曼0�nt��r֫3��z?s��T$�� %��fے%��tF�i��rIx��a,}��{�op��L.o���vx2�9n �w��=�>�x�_�IG�oH<��M�2c�j�WGep�r��u=��(����:��YK���,��ȍ�1 ���c�`j�\R�>uB-�W;�֗/_�%�VJ_�"�\�R�+;r���e��2�]��G>"1��''��z\w��^2U�2�a�:(a��{h�
7�����+�!��1W�\�u��>PDM�Y�`�� ��d8Z�tZ�x�aV53�	��o�����-�Ы��gĉi�����N�8���<���L�|q9��9�dXF淎	�t�3>��+̪��2C��n-����{+��p]�\�:���ߐ�)J�k���XƼ&0�rP �#����H�(�kj���9 >���)�#�ױ�M���qDF�4�8x#�� n���+��A����>|D^~�e���;e��-�ç�r�}��?=|R�/��3�N�[��Z�h&�0 ��[�D`,��u =�� ��!i6��rI-�j�a�uɉ'��Zg�Р%�V���&��-��sH��}8�$ m�m������#H��hK�9l	_ ���|O��%����\�s��4��p�6붏��\tk��Ɇt�G��m$5����/����mk
�;���4��\j@f:c�l@��76���c���8��0��3�� �� ��M�y$͑U�$4L@ñ�Nz���D)��A�;��?�JIg�S��;����:בY�%�|\���;�1��/��w[���3Ш����|�N�
[.��RѶ�� �QW�N��qIe�v}xmp�'N����[>(��ה�}��V�0::"��w�����ټ*ӳ�t�m�t��ZWn�*<Q�_W�����w�~c��f2��` z 7$�x�����hN7躹`���Ro�d�-[�"X$K��^�S0k+����l�Y���>�������-[�X��p�
Ӎ�1ʫP��|I��W�l�`�ks��e��$:�d7�Qʺ���9W�|�pƐ��q������;��߅?�F@Cf9����Ը����\�.q =>�Ŏ�  �>$�A	]�T2�99�i�C��@�"�5f�c|�nn��ٞ��q?����c���y���8A�>C
�0n�����\����� ���"�M�{%cW��t�2I���F�*�j]�كb�g	J' ��	�&��߿h�w�_�x�	+���e�0s.�Hw�¨��Cv}$š���
�f۔�}�|�w�����س�@=�� ��i�&��F��lr�`1}�y��2vuʁ_;b�@~jz�]��Ue�c=��o�T�}��5�ڹk���~���G���~���p�������G�J���՗���~X"��D�I��B���xC�q\��<��T� ]&k�"��&�ӥ>11f`�dt%�w��~�qҳ���ZHR�83�r ��f�o�����w\c:��O_˄/(:P&��F�<2�� Б��'�aKV���(=�>��^�U�)[�g�3�pe���a�����~�3-u6��_5��0K^�r��q���^��G��D�m"t<+�u�<t�Ø�0&B9Pn�xg�S09*��+�"w�q��A��K$e�P����c���-rX��|wV6nܬk�Te2,���S�"�/���~����#4Mc���@D@�%���m$.�V-��2Z�V�!S����Ε,�<��r<���F�o*�5���]����1�W�25>�m���'�w��]i7ʖ���d4�.Q��m�v2��*�u���0g��ē��mvs��-.�����@�Ns؁�<0�n���}^�2����ܯX��g}�K�,u�ϡ,@8_�3,K(2$g���|�;�	�������yr��2G<cB� �+�0��{�"��-��Y�w��>���<�)>_���̥jqg(p�Ƈ�B�7&X���f�SI�wc
���V�,�B��C ;jȹ�g�L�"�W��3g���}�h�z7�Z�%�d�˭I;�I����կ|�~�a������ܹӔ34���܁��9yg�!���%K�t����V�����,@����i)(�������P�a��//�rC+��H(j���*hI�27S�M|�I)V\��H4nq�t������h����*@��7�f�M�,)	5��mboZs&~�ܯ�뺙7䞻�Ƀ>(��#�j�d��K|�t��5����puG:q\��b&&�@�% ӵ6~`J6=k��C�=d��e�밾��n��Ų�=��q���,Py�+�1~(� ���)j���*+�L0M���"U->��
�u�s;s挍��*�}*��:!.���.�����L�u�]az5�h�K�h�`����2*0_�W*���b,������e�ݯ��J�e��e�ۗ��+6�?��tqN���)�֌��{�]w�}N�]��c��SO�Z�;ԕ4Z����5̤Ҧ�@у��ʌ�O�șs#�R�$��Y�v���{{��Ϋ2��	��Z�Պ'�{ "�r#�N$�usѪ��?��u�n
Ec��D�`��?��mVzċM�JE�z�M�l^"��T�������Ę���*	U�(�R�������Z�N���ruΔ�_��_V�	ɾ��ɏ~���n��w��KtC{W�x�ǵ����~��>�W��T B�^ԫ�F 2����pX��i� ��=X�lU�>��&�>���L�3B=��t�x1�6�{f6==�Y��B	��NkCQ@> ���Oy�^�����r�0������ �Cс�Ƀp�j�`��ݿq�FU欋M����׌+aH��6�����ܶm�ʣ��P%�c]��eK��E��w	��;����K��F*�����F�}�ګF"��'��Q�R-��,����^`�.�ٌ~�j�GR,U��j��"��  z 7"�ݡ&-��Y+�A�1)K��ܒ����H��;V/���u�ι�bu �(w��"H�R�R�X�cPn��;�Ⱥ�vE�򕿑��iqUk�j%i���=weW�N����3#,@��nn���x.��:3:oX����܆� �{ƹ 
(%d�㸴�	���c�lU��������X A�ɘ5���|�L���39�1_$�qc=�1m۶m��p��rW��}�L��~�^+T֔����{G ����� ��q߬�'3�{p��x�3��y�)��U��2)�e�T���&"���Ay��J�A> ���:gxQ�!�r���Gh�!.�3,Ux���ǭ��,����7�(�I�Y�^�_���ju&h�ȂH �܈�ڭf���jy��F�2�K�<zOXU��M,>��>��,؄��0�F�q�S)�f��U�Y�< �;sХ��~�������P�|�%�P(ֹ���[:NS7��3��]�b��@��0�nm��
�T*�bf�O)X����0hwR�B*��5O���nu�����0���2�O��̰|͟�NN|�� �iUc^p��2߲e��+z׮]�����{g���sz"0&ѰU+����w�m�u���<P ����~B�s�:�����c^���FA�zUb�9AC6�%��~!!K2��q�6z�SO='��3
�.\���!��s�e��%օ���9b��Gd�����m�L��G��q͚Ԑ�����Gm�Y�������&��=�� ��!���nj ?P�:��%B��w���b���־��^]7�e2�? �.M`n�ľx1-�P2b�VK������\�l�s+Ќ\�h;J߆���:�%2?g��,%�H�X��1sl�$���i��}  ���K�E`��L�c���K�3���V��q���� ��x��O����
�6�,7�1Xg���F&�: ׄR��qx�Y��2`~��֠�)W���a%�����G��p
��>�ϵ��]?ֲ��}o�z6��(q��H�B�	)�N�2�x�hX�W�,���rU^R�w�{�'����L�x�]y��1'��9.�X$���g�	oB��G�s�êςXG/�����O׫o�@dA$ �@nHP���,�����z>w�PXM��X2e �%�B�5��Ջ7-�)�Hw Y�`�{�jV&�{!  ��,�a��*��ry�6f9v������<d1t�p����� a�.,QX|���6��Z	��W/��E�Y��'\i{ �D5 ,E���i��|��� 4�B�>���f�6@nn?�K�pM2����5��I�2�kǬ{��������`��&s ��qP"�tH%����p���?k�}�y<��4��yT�:�x²��N�d��K�;�����XN�"�mR�.��;l�!b�/�����ׯ]k��{�3x��)8{�`5�΃ԒJ��VwK���)!ɤ8�d���e�G$�Ey�[m�ld����H �܈�"�1H
����zvnF�
3V�R�V�����4tS��֗ؤ#)�����aZ��j˭��*"ⵦ���{�ڐ�&�zuī��X./��\�����n�Q$l���ߪ���d;b@l|�!�&7oYH lY�	�Z���m�9D:n^d�3+��bdCR�2V!�� Fp��#��	`$�A�5�� $8����j����!P$�����3���@@b�=���������w�m�I�,X1���i�צ�zN{�~�ܫ?�MJXZ�lC��x����j��N 4*#ȋ(��V�<X�A��i��E�I)*�cL��o�v�d�z��v���RG�s^�ŋ�����$�k<��xĞ��*��ƿ�v�Ʉd��JyF-���������g �ʤ�[S�G�}&W%�$�le�ʁ -.�� ��1	�"q�v�V,�dnZ�c��Q$����vX6��d�'����%�8�j�q9y���1�4�Ɠ�!���U�+�!�-�M)�;Ћ���;�+�\Z��5����A������%9�?��p�����4C� ��
Y�,^u/��;��V{	�8X�Q��=F��W����p�Z�^�ޞ�Y^ ) +Y�HL���^č#Q׻�e�Í��t���2nt  �M.�cǎ��ڡ0�4�"�ΘX���u��q|��� OX�P*��^���v{�ӝ�7eF���<��{�^|Φ.��*�M]�Nh8��L��,tT�<��<·��-x�6G#i"L�b����Qɥ�妍i]ǜY�]�܁����bU���굫������ҿh��úB�K�҉����%ƕНW+�ՖjqZ��d��[eǎ{<NF���R-�e�Ҩ<���r��1��G�:<A���C`��  z 7"!݌�a���z|¬�M7�$�<��mr�W,���dSS3rn���>uF���2%s����RP��j�X����W6/^�
�}������eI��M��qyG�Z�=o﵍��Z����$#M��@�(�˚]h�k�
�����k�3����ns��G�@��[�۫2� �5�c��zV��[�2��T�<�Z�#�ֲ���
���`�^� ����l�0�`�kAA�g�6�L07��+wc�>)OI��BC �^��gB��\��}!��N76���e�+�@ؕϽ�w����,S������{g\�b*j
f���Pq<!Ըߴ�f�7���d�Z���.����7�/��/JR���菌ܨ:;'+W,�����g5m�n�V�z,�3��߬�˖�~�c9q��>�)*��3� �=�� ��!A�˄��@���ˮ�Joo�%S�O�˲��-k�;�+5Ś'N9װ�b�Ē��%��_�n�&۷o�\&kn��G�S0��ʫ�)�M�☉�N˟����Jڣ��W*�	c���V���7��k��,;����E����'A���҄D���Mm4�
L�����ݘ��R/��4����IX��c�&�k&�Y�;�T��y�|2�AQ`,�}���N>Ƿ�k����|k�P�w���'���I�k��֕�̮kTh\��\�T�8f�������@`�q���@��җ�Ƶ�M��kEdr�(�m1b����[�����L��M���o}KJ�9UP����|�F�8�O�G��0Z��c���t&-K��e�ΝR,�dbrZʵZ{62 z "�r#J(�����,��v�27;\�o����X��6�7��)�޷��^�z�%_�ˋ���-�O~�礻��Z��ٳGf�&m�5zX� �l%��X+�⬺�_�<*�ZQ~ᗞ����G�<;.Ǐ�������%W��5�罝a5���l�J��\�,iMCX~:Y[X jZ�T���^Z�y�%�b��N'�cM� �{B���l���M�5�&��X?P�Z̔�y8��{8�|�O^�k��h����MNvZ���w�˼B���Ƶ��`en�������+�HR��f�sn�����{V�0?l���$��V'~�ƺ�>|L~��v�	�CV�^��CN/^�
D�*W$��Qp�����Mټ�V�|e\�{�'�yP����	�_P@䆤���!w�H@ʁͮ��L.��M����\�s��m�h.�^�D�Z�f���MĥZ���!=�K&�&��r8l���WezzYnF:>ɒ�˥V-�~��1��M���,O�,����Z��� �������?x�~t/��Y�����.c�N�1s���鍀n$%��I%p�}Ҥ�u�e���s��K_����޹o�ܜ'�J���W����:P��{6��*����خmϊ��E���v�:�_���ӧ�c=$����jed����쳯�L�"S��23W�R7�)�NUkW>/gΞ�����lݺU��r����}J��_������+�}�23]�u�6HF-ytxCr��+�B$jc�m0�H�U =�� ��!i�Z�L2%]9P\v  )����$��F�]�r�!g�]47(2��ݎ�� ���O���d͆u�s�n��޻,�{f��|����Ȩ���8nKϫ�*���5�W_���t�d��=��/ɢ>��b�y����{:�4�QZ��en�Z�v���K�4�q���`�r'�o{pL�c�9�[[���9-{ �fX�αI�J��9@,ݳ��!���5�������&8mO��+5�h��)������? �v�����\�|�T
�s���X��zP<b �����+Wʊ՛���J(ڒ.�sϽ�Q��2�%��G���ey�'��������o����XR#捱9'�5�iB�,}<S�Tښ���KT����lC���9K "�rC�I$[a	u6������C�Y����SO_6�r��1g����|ONƧ�e�P��n��
�g�]��֮���~H��g�IY�d�ter�� �dF��� ���!�j�`ԯ�z�q�(���f�w_����G���x63ȩ �-)��a�G�
�k�Ę�m��c�cӺ���� <�ms��x��d��ǚ���_^fY�
���B�bֵ̚����+���!�]����$7R�
k��Y�9
�'����NǇ
I&Ҧ0!1͟�N$�	/Fԍa��J�z�ócme��ԂK�Z1&Cx��;j�~��IX�HzO�?n4��JQ����UI$ch~.SS��<m����>!�\�)8����Zy�\�~�ȑ �=�� ��1э�ZS+��8�]}q�6I��!��slt��g�Gy�!��mF�l��;v�{w�h��)��%Ṑ����W���d;0w!��d<e.�Ҝc ���R�e��C�Z�.�5�;��	�>8��	��l��E`' ���=xz[�0�qg$��	^t�C`Aܘ��O�[�$�����Gv�����ieS��F��)pq=��2~N.v��~�<=��>��D{Ν�Dyd,�0=Ҙw���mU�V��k����|���ԅ�G�o��O��rd�r��QS���VW�d�R;����y�*Cc
�a9y�\�4*��K�d�a@�d�xQ��� ��H(T�'=�� ��	UJ���hQ`GF�a�n���{O���Z��*R*��
y�q=vb�'7ܓ錁4ܝZl��l�"K<��^x�UZu�����KV�w=z��m+�~-쑣GN�~jnY4�Al?�t�qK��qG3��O�J!(S 0HDù /�yY�F+�Ie��v&��"z�����!L�q�>�����O% �\��	�d��x�� �	[~���}�u�x=�m֯��~πt�[k�j��Oy�������Ð�?��c��2��|��tA�n������jX�h'�u�'��<���P�M���۶�鑳z?I��r��)yg�^�:!�xҔ�|~�LM^�����m�����Ľ�y�w�B�Z��ͮ\�
���@D@�E7�h<͖Jsw3, Q�Sӟ�ZБZ[ʥ�̖x�U�_��]R�%X�T)X�n�ܼy��<qBΫ%�������:26\4y�wd����~,�����lp��墠�0�c��-s��=����TU)w��B : $�x�4�Ԧ��F��&���% �]স�\Ҵr;�\=뗠B�9 �-u��<	� P�=��L~�R���úy�۟R�1�>o�d�#�,�3��U(����?��*2�eg};�
��;D�����i�ܑ	B���$RU��],��B8"�\��
�U����:�:�\��2Ni�Y6o�f	�}�������^�{�q�g_��G�������k��hCu�*�G��o�;�%n�B��H $�rݢuJ����~�6WfN&���𑣶9�&�V�J`Uk�1E+*�͕�ZrXͳs�d�Gy�J�V�[c���/�,o��g�06�F�f�K�Б#�b�,]l�h���?+��)�oK2��Ř��<dt�訆�%4׀�*b��F���'�	�c�l������U'���vfB{����Bi���O:�1�mM���t���	!���]�֝�	dh����E���0����b��+WL����(�S2��J
y�I{�W�Y� Q�ÄJ�?	x�y����p���n����'.I.�+�>�aXak���[�f]�=�~���9I�X!}=������K/�D2�ݒ��<f欳x�3�2j�Wt�Uٳg��^�T�H��XF;�.�<g��r��q��׾.}�P.K�v�|���H �,���u���pR7����/����x�X�s�.8���X�P��R�ძM4�6W`Ŋ���d��ҕ�Ys�tcQ��7����1˵���c�'��/|�jWe�p�Y��sR��Z��F��^�x�m�(p��K�s�ò��FL�uQs�v��&�A����B���G}�w�7����L����aZ���[��]ی�CY0�#����fn��毯qM�G���G5k ��lK�,�����{����LuT,����qY����X��{>컃��^_=;���^�(gϝ�e+V��U���'`�͖���J���� �V7���蕗_�W^yU���%�]85l<+V��z�j�	��r�ʌ�d�^�V�cQE�-Zb-W���g���Ĕ�X�R�,[V�����$�@H@�e`��vq�B=��.������Y��y+;��v�w$�%����ų���w��I�~,�C�)�ŋ獄���'O9�pl��ܺE���o�q���?&�HM��q�|���ܤې��ۧu�W�PK\ˬ: �mZ��g�p��%Z������2'�]�ן�g�&&$��!��v��)~	W(?Ph�J< q�[�҂gR�f$~�dͲ�Zu4��B�F8T:���F��\J ��ֆ�w�7���|'�<�6|���1q��S@�xԭg3��X��G�|H��e����e��we���>��'de�%=?b��P/��������>�=�n��W,l�Օ7v���]����T�!9y���:="=}�z��3W�nqb���Y�S��j��rOO.h�ȂI �\�lܸ��z��c��������n�`����-j��ikl���a\X芮�!�: ���h2j@4=S0p/��u`f��e�֔�\�%5�u���X{z�2;}�6�}胲f��<xD���3R��N\�uز~렁e�5~���G�LFR� A�����g�ӍN��ߘ���R/&~1I׶v�^"]��d4ƞI��o��X7掵#�2���j��L�w�e29�9�Z�ʬp��M7�dǃK>�3���@~���.�9�#�cx؁���0g��h[������N��ݮǾGO�x�>U���fd׮]v��K����a}.ڲt�?�i%�h7��"�͸v���Ti@��fOy$����z#d������i������_�'R��ߡ���WM	d�$ �@n@��=�|�Ѭ���%us$1��ql�
B���m۲Neјsz[yW�%�՛`ө��L�yW6��W cc�d� rY�U����o��@�?}H����N>��}�Ld,���R���0�m���.Ѹ��B����b>P �	����uZ�.A*g��3�����{u�dkc�PaM�� ��8����� <b��.�50w @��q/`:�yȴ��m��==v�^������J�1O$b|��#�w�^���;��Iu p]/��{�O���DB4�Pc�'���1(l�:6v��m_����c�0G�t �֬ ��<Y?z/Y0ߝ�9v������<W�U[��~���)�Vi�8$����)wͺ��LI2�-]��۬�Z˱��Ui�e,�3�sJ�rj��Ԋ�gA����q�-�Ta�E3����I �\�\�x"}�ԩX7�x�k.�=P�F8g��1�!o5:�*:b��
�H	K����d�d,n�¨!��s4b�C��A�Z�VU6�ʢZ.��{�n�RmV&�/v��},��M �b��ə���p? R�(���5�g�8 �p�{<��3�� ��d�10/��a��� �p��@ɸ4:�a���( %������xw�y���dp�Dǡc���+W��� �x���߶y�g߾}66�w����5"�����o�`=ùf,�}a�p>k�Q�����1�kb9>��%���Z���DG{�Z������A8�n��  ��\E.�\�w���� �2W*���fC��<.5뉎�'�~���#�
YXTp�==U�$>pėJe�/!����A��*��p���u5�,���u˹s#Y�l2 ߸nn%l���Y$!�xf����ǣ�)�!ȩ�B\��'�B��Z�n���M-��s� Ĵ5�X�l�\<F��q�DI�8{�%���L�޲,w@��rw��P(fqZ�R��۾V���h�1==i�4��`���?��Y�u�P8`�www)8��2&ē��:�$�J]���]��Ӯ`�/͕���F�cd'�u��x���R��1�(��)�;�j(� ���~��	ٹs����o��в�r4��7l���O�ִ>�X 8���u�"��-��v-r��.�����IqH"`�\(ǎ픎�U�yb|(P`�t�s�}����/(�G�@���r1�sg.I>�չ;�ZW�60��Rv��0ȁ!U���ͪwt��k#4���x�c��dUq��+�l�Ue�����+juW����{hV�(%���
lY�S˧@�#rt�{�{�yX�k���WoRc$�� ��nQk)��S�66��Y$	��8˹m�rc+W%�-3��+�r�p���}m$���d��v�U��m�.!���:}���X�j �eKMQ�4rN⺹'uXm�Zs^����A��7q|�r����X�e�~/q+�e�E��`8�1&6u��I�q R,cc��J�� x R|���pGC�����a����D;\���P$p_PDz�! 
@����`��q����N�~�r�x�2�y<K�`�3s�sa|���pX� �T&ic�f�a�f�X�g|�!�$ r]�t�ul���hl�Q�e�O�?���[z~�8273� �3k:Wqyx2����̸Ta��u��yG�
�mbbJuw<�S^|�Y���仩�+��k�T�;�8}s��*F��H�q�Q��@Y 	 =���t��T*^lVebr\&��S9����ݭ�
�	#p!{�lqN�j� F:11��j)I�%��SI뺆%pk'�	�� �;���C�3��X>�����X�~��2��[�X|��cACB��xv�u)	A
�y�f�T?Ʃa�> �� �$)!��7�h9.����_�Z���c����)��q�bZ���]�ܗ����:�*�5yq�73�-�R�^��*Ir����9�ea|����"��(\���~�F��5���t��nq 7 �c]`��PlȜ�o��z�B��9��"�+��,�0��ón>���P��ʰ.�r�T�J��)]��P��{ǽ��[�n��yɀ��s-�=	fh�'s�Λ7�bkQ)��̙�239!w�u�>t�'��������5+l��#W����d�MuV���v�2���` z �-�����mg��
O{=��d���V�ˀ�kZ6��EX<�l��Nh��n���MNy�t%��m7��Z^���%Y���u@�8�\�g����ޑd�%�xK���k��XU�z͖%�E<�`Cf��.h�6� �c�ԅ���� ]�:~MkPX� w�FM{�kx �l<����������j Tzp,�hc=!�Ƨb���⺸R���h]c\�O��#��`�����(:d����~X� %�ω����!,��l���X�渞��<����e��s��iP��7��|��W���G?�
A��9��X[���@��np�.���6d��p�8u��n�LZ>��O[ܾ=���s�R�L���7��;v��@�*~��8�NϠ��M˳Ͻ"g�/Z餮m���SY0	 =��[n�>^�9v����a��3��:Y�n���eK�e���S���g��+����j�a/]�B7Ҷ�� +VW<��V�N)x�<R2������ZZ��%�:�t%�����l"�kzp�C�-aCG� 9|���]����@��L�93�]ɕHWW�8�!T\Mu�C�j�ݨ�`��9횜 @���!�d0XǬ��ۜ$4<�sc���bﱔ®m,�㹬��u���tHa/��`�2� �����?�n��;���+��{���V��j�s�Oz��:�?�j�zM&�+���8 o����Z�V6n�"{�~F:��6|朼��ٱ�~ٺ�V�Pa�_,��W��~Y��6���|��Ƈ�כ����Z�Ǣ�����}V�_8-s3�2пL���Fi�jGdp(/���j��O_���x섍p8 z &�r�244T�8}**�LRڡ^ku�b�2Y�a�.R@_n�f(}�����:�K���i�h��Oʡ�G�^P�x�$����ǭ�ŗ~bV;Z]|�ֆ�����D�Y�f�1ε�3f�ێ��˵���b�ՎՈ� ` k��ᮆ[`�"; 	1s����醕뱆���wT�F\�V,^g��N�;�h�����5�x�����`��Ď׆�=��ٹ�j�$7~֡��]�7��*��&�a����� T��ٌ��z�]�x	o��\���R,V�dɈ[�V��sK��9J������|G�茗�IA�\YH��?�яX~ �5��^}>��>����zT*e9t쐼������Y�EC���6�O_zQz�{��|H��)�pnR���d	�PT��;�ܮ��1}�.��x�rd�$ �@�[t�O��L��N���Euc\���-2�x����K|����ɶl�jq���.Z=1b�5/�	<6td�ߴq��ڽS����RR�����e�u,9�FaŧR	�+8]�<*����?�a�4Jr�¨��o�G��Y��<��%�K�q���N�{@Ʋ4v#�)�\�~O$B�)�q���=+�Խ�[�ڮ���KNc�0�KzW '�A����1G(��م)��5������7�����0>���V8���&t�s\�'������
����r��mx�3&&=�:�p�[�P����DZW�v(T��s��}�vi5u�H�rFu�0.������� ����<����>=�۔Zܡ�E=?,������lU-�?���`�#�y�Ǥ��C�A9e[�K�Y��^����.�u�Mr��H4$��p z �-cc#='N��FP@���U˥+�gnb�V��$��� {d3���=]��cǏ���JR7dl�=�}��������>�8���;f�3>���|Dz{�2S��g�yF>����cPRD~ts��[>�m�� AluҘ'{w3k�y�� #h�Ӗ�wW#w8��G�4�g?u(  k^��2�*$~^t��A	�O�=	���f|Bk��8~c^8���h��}��G�6�-��S��������f�k��hv�	��P@�̀�

�
�p	�;��xM�\2�%��w����Z('�����W����/-�r�����q�l���<����:tH>��#���~V~�3��?�O�I�x�e٢
'J��w�t���jO��Ы����W%�EW7]�\Jڍ��(��33���I �\����%k�Zʲ���4���O�W�j�ܾ�N�8э-�����e���/yQ )�D�[����^��g�e�-�e��=r��!��c�4rnXĔ�wW����G�|_�{�{G�+p�תu��%�p]�ב������SB$�ML��K<�k�Z*K"3k2�θ�����������wgR�sfF=A�nhr��}M���@`'�,���H�B�X�m��n�M�T6�A<��%(B"����=�A���ϰ���n�Ƽh�۽�g��#�c1���JG������WJH�=~�\(��t�,�G$��J�&ɌKP̴Br�w��F_�4Zu	�5�P����7���lܗ_zA{�ay�]����4��hJ�7�$�����㦀.�M�6��1����K,��[�z &�r݂��l��n�q#�@�o��icJF.]��j��1L˰n;�2� 0�}iw����O~�Iټ�9|�e]��֛�yP��2	��@lC+%f����@k6iY�X�ŎA͉x��V�Y	�ȋ��k~+� `b�V�T�u,V6�|�+��s�<��MR ̂'�+���"f�~H�J+��Qix�9c�8�B'C1"H�����L���6X�ZP����?a͟���#��A�c��s�r`����~W{��/(�Oy�{k�,yS
J:�T���V��ho�C�dL(b�<���w\�;v쐷�z����/#�=�ݼW�P�$�ٙ�]�w�ޣ�="��=��7��:���27[oU*� �ȂI �\���]չ�R5	YF���+2vuB��u������ʩ����o�&���g`4v媵1-Ѭ���s��=���e݆�FGZ�+X�t�k��d6f���.u��u���Pp�[Ʊ�wܵufX��y������N� x�jua3�;x�J�ܨ��� P�G��\��َ��@��V4���.i�t����v{u�a��"&�q�0���	�ժƔj��lLMMwJ��f�	�<��B�z�֟�tf�3��@��Ѝ�D>�,=���,�q}79f�3���<U���N�׋�"F�~n��bE�}I��4����9@���I�n��x'D�I�e�=w˧~�gT�k�3���U�;��.#gϪBАt&+c�S�W%���˺H��*�O�G��+�8��	)L�HN����\C�L �,���u˚��S�l�z�ȑ���e�d���	9y�e��|��ec3{��'����r�d@V�7a#������/�(����EX� ������	@/�Z�hw�w���L1E�ɒv��$�1���86�pM�@IU (��N:�3��qM6���H ���x�T����,�d-��u��uZ��|���
X;����Er�f�20���M�6��@B�>K� ^8kˤ�ŋ�ll��u���Ӂs0 7k�Y��$rSy�9���b�_���i���#T��~e��#d4��{���\.R���$Pâa
B?�r�*��!D>##-�������w�� =)�:�	!��<~X��-�l��~샦��&%K�|�	���M��j�b� �Y0	 =����`���oT��m�HWk]A�nh%��M\ڰT��k�(��$��[W��Z�i1T ʇ :p�c������Ԅ,ZX�,�Z�e�d�9y晧;�@�^����N��*����u˴��女'^�_��\� p s������@?k�{�36 ���Sp]d8��(�x�{h|�A�j�s��Y� ga�c� U$e���h�.bf��ݍ��lx:�l�b��1�Q��ZC��w��Ļ�k����/�y@9@i���3���߽���zsZ�,9�1%����+rMN ��5��w`ߴ�7� 2��?�V���)$l�6vRj͒�'����S�WFj���I�K֟ ���*��~~�ay���ezr�>ǳ���{���q�r��������f��1���U����K9=|D�d�X������/ �rR�MM��"�0tg��X<)g�8�w8�,`X� K�g�Z�T�u�+�Z�ZE���a�Fs�Y�H��80�A��ܳ�C
�5ːA��^p�|o�����t�i�� B��7��ޞ'jq<���MA�-� o 1��Lq�I�Z�����j����4�P�`f9�C( ɫW/v�d &;�AQ��ǚ����ze�>�0��˖�i����X3zC��H�:ָC�H���*�����=�����5![�����z��A���w�L����^�Kj�˝?�/Q����7B�Y������y��	Y4�\r�^>s���l��j^y��Չq`x|z�����D�)4ᱜ�\���g�b�9U��?�g'"�ʬ>tJn۶Y�j��ߒ���;T)������ޓ_|Ir]ݺ�N�C �,���u�ٳ9�ޢ���K�D��ȥ+
 �$�rɎ([?�pL2�Y�)��J���*���믿.1��j}>���f5V+e;r"��:�m���B���F��f\�zL؀���%sybo�"�R�yв3+��\��L� i0��@���ذ|���c�8�IW����zZ�H�B9�z?p�33O���u*� �ġP�=0��p��v�ڇ�vw>�k�u�8������ȅ��PV ���AY�8*ޢ zP�c<\nv�-�`sܫ?��9�ԧۛ?t�3߀.w��X�^��>�f<_C:���BjE�M�[?r^��M}ޒ���jbvvN���LN���ԬT�g
s�~�=2g�e=�;��v��c'Ny5����>iá�
li�)�gd��>U�e��9z䄌^�Q�?0:zY-��=���Ҵ�Ѡ}j '�r�2>>��|�R²���q[\�V�Ѡbs���9 �\,�1�DJ]A ����?3+�����82�!�i��hHbu�^�3]ΰh��Ǐ����{v�!���W����o��C�27]� "��2N0Ľ��(�`IP;v�X���&^�QXڈ�C�ׄ�N:�U`��C�v��h��x���%llH~��W�s���J� ����}�(^X���qk�q���d�o��a��P��	ڬ]g;��[���h�Ӻ��h�Ǳ�˵�m]g�����8���m�!:H���7�r��ҕ햁�k`��+��Ɏ�hd=P�9Em�׿�5=~���|V�^��Z3����N�g9��K�ҔH<'�G&�̅Q	GZ��X�;A�}J"Ś>�����{ &�r݂ͩ\��Dcm���k-�[�����Xn�m���M?�0�W�$+O�N�z�aQ
rI��XK�[w���]ͱ����ҕ�KW�d߻�����B�,_��6�������+��YT�C,!O�	o��찣!�,���JΊ���`	CG�9��َ�aL�j�Ξ$1"q����A�!�;���;��(�C��f�,��Y�%�tw��5\Ӑ�)��񃃋�7��/��@�,U?˚����X5�蘝N�4��1�� ��i�3s�ʀ�h�!�d����sn�!��)s�ԴܵB�%nc�t�c��0z���<8��q���ǑL�䓟�Y��(H42�з��s�^��Q��T�m����e�e��,s<;|N����ӕ�+�t.u�����j�l��U��0�8��	��Rm5�<[�L_�D�Qi���r��@Y 	 =��T*�T˹�2�����BqI�Q*��ȓ�z�;�G/ti��s�[HDa��C�T����P"f%YjT��0����䴬_��xCr
��!K���/�H����J�����6�Utq�$V���������i�iX�pSC�@�z�0kq}��a�Ê��
��t�\� =X���C1������8�)y�q����6w7 �F� ���K������1y��G\|�H�ù�"�ݏk��s��O���a��v��o,Qc�8Z�.3�	��k���5�:y���%��(��9���AE�ʂ��V��!��N[�A���XStSK$��GV*|���W%��ސ������4ȍUP�xn�&��ң�ԣ?(o��WFF/˹3�e��e�d�bWb����O ��[A�O����)v�.W@�e�A=��� ��n�+dә�3�ې�%���[���0���A�R�V��!�]A�"�qs�[Fb$(	�Y�l�UK�Æ�k��%�)�~��������j�}d(�v�H` "�.k���u�<��F< ��qmX��֭7����5���NgtN��-
f9$
��jj����˗�0P�XP$�~��s��0Zl.v(���!Ο���zK>�я�� "ң��`�u�8d�� �˚arĳ8�m��p�N%�d5]*M$�a3�����ą��p!�qI���ԍy^�h'ގ�J̑�X�D:�&��>�m�x�1�9"����w���qryV-�[o���}zF������fe�@�*F�V�V/�t̂ıf�\�T��d3��Ǥ�ϾuDS�xJ�d�4]
\�,���u˪U�CCo�[۳t(��֒�J���`fk4�
�a#4�4A�Ym8K=���Ujã:���:g�����j����`���йb��X��gE��ڵKe��9sQ�ˎR��%M���p͆�ݑ� ����> a�l�v Q�	b(Cb^�a3����X�, �7�E�Y��mYq��v��A���	nP�m�fc�w�%��~��z~��Ap> ��8�F`I�3�[�BW7�#�,^�~�Z���O��԰�^c\*��%�,��pϜ7߷�'^���Um�{���)}�F���|Ýf�8󅇌P�5�NX�j�B��ǽ�U��~��P�,��[/�}��M�+���┈����Դ=U��jW�^��r�(�TZ>.}�CU�4W�T"ֹ.�@L@�F���\�Y7�J]-K�x�Y��N�PS��Z�V1f�E��9��`F7�dJ&\?��iG��wX^��ŦH7�e[7�yV�ɢ&1�Q"eԜ�p¨_C���9��n�F�ա^P� � DXd �T2�VڔY��B'���3g->����%-YԌǣV�����$�5pA�9;��X�M���d��|0Ƃ۟V0��p})�  �7�� � 7�ZБ�0f��p,�	/��Q���b�T�འ��·K�|�(�üp,� ��b�,a� �qM�ƽ��V�tz�3�Ŋ����z�K �Y]�����&պ�7(�/
J����z�����;%$@�jAff�d��.Y�t��]E*��SɈ�]5d�OM�u�2��Ų����A� T2 �@L@�e���̙3�7��x5\��rU�8aV9�t�	E�1-��率 ��ug]�3sŶ���$�T�c=ڹ"-3�ŵg�OZ��-
H|�ǒ��2��B�$��� Z�֙܅���HԕL�oқ21�L�0�ﱏ�e;{.j2��"�B��v&ޱ-*y�8��3� p�{�����hU�=&��7��:�o��1&N��QX�TzX����!�����(c����p�
���sp_�t����4�?G3���\���ʁp,n��=g>��17kL�J"�0�"��vr0z���亐����KT�k��E]���Ւ��-��/R�7/��.U W�m[7�E��l.-�RM��s@�y�e9�����n�z�jU*��` z �-�/g���tetS�d�R���[VPK%����mgmSW96p�� ���v#[�Y� �Jq�ڎ�zn#1N��z��)��x�3Ê�cl�}O��W~"1�?km˺w]RCF�	q����V7�d�g�QK`�`l�=��I�g��f�!9������~ǹ�r�^&=�pd�
/{�\ ���G�}f��� �X4���)�Y\�Dx=RŒ˝�e�/ۭ���4��qm�� i�㇄289t��x@Z�$B��u��bIjz߈W3D@>u��P�@����x|4�x
�~�f����b֫w��.�ԩaU.�w�݊�ő��Ziʺk;�s~6�1e+����*�1�&1������>�W�~�M)*r���w���e��2W�����+����G�=w�+?����/�O�xʊ�kC�H+ �@L@亥X,ER�T�O-�3�����Us��]�F/Yj�EK̚8�J�zu\���!���`�%y����*��D)�,n$v<<���+_1淙�q�t�*3֣��j4Z�N��t-��v��ؼ����� ׂbB>�|w���� p��e�Cخ���z�� l���I (A��`��2���{ B ��+����x n�nn��`=ΰ���lr·�K���'I�θ.�N��f��i��H�q{(P �*���k���/( ��c0�c1���rd�����7���μ+>܉�SP!p��)k���?xV
�eY�t�)��0i��-��&�W��;��j��'�Mo�_��_�W^���Z��ͽ�,��{�ҫ5d�8#7o�lI����<�l�֭����s��/�O��[1� �=�� ��n�����C!���+����e���f�z��7޼I��Y���g�����W_W�*Z��R�V�~�ӿ(?��Oe��jo�e
d�=���s�}G�5+�5���P���;V6�f�r�V��rAP�;6;�5f�')�y��ě�t��ʾ}���u��H�;o`�>W�b�l�t��i+/���! �!��X��'u,�������J���� jK�	 ����1�:��б�8K��v��gxc( �q=~���^8s4?/	k��r8Ix���S{�1�=�����{B9����k�ho:,�E�҅�����{��{���JM\�%����j�3`�[���c'U����qU̦�
O�<�29�$���y��`Ǯ��k��3�0y��q�o��Mij4aɗ������uڳo�l��Vy����#�dj|Bn�i�}��JQ�]	]��Ѓ;��3iߝ�@Y 	 =��d2Wi5�eP��*���ˊ��t3]-�LZAzE�ɉ��k�����c��o�����+[�_�.�jv��9y��~Av���3XT 0��hd5���XԬpl�O��GeŢ^9q|X~�w�oa/?5�<��s=c��$����LciΧeɱ�4-r ��`�� �8�bp/�غ�]��� �c�N[ ���*
��c�Q',s����p���>�_����c�s1uf�3V�1�;3��:������gd�cf>��4�9`ݙ��>�s� Y�2��<P�`i����K�<��t�������"U��\�=Kg�^T ��ҥ�e�h`�dHׯ�p�fl̰Kĵ�z��җ�$�/]U��s����'+���ŪX�����T�|/��$��o1V\��0nH5�Y�����[oEB�pL	d�$ �@�[6o^_z����sgOo���;���H���8��
�u�6��c�N�Z��N?%W���˳f���[2W(ɺ�N�=#���f�<�v��L���|�R����e���e߁��{��y�c�d)W��r�6��wm6��0�u��cΈk �\9�W�̚m��K�kرN)q	j̜F�z�r��-�^"[��o���s�#�@�Чk�����Z:\X� if��}�����z�{t�t�3[>�ՅC���Ħ,C��叐 �
P! �����A�2���Rgm|�����kal�&h���7�+w5��R��F�$��d^��?��P�^���?��*UѺ��vmr��Y9��Ay��7�g~$]����_��#W��g��w�yۈ�Ο9��MFVߴ�y �1����a�V>%��yX�'�,K��tue�:ל�I �\�tw�j,Z6u��C2>6�I�\�i�袑���~��t3����N6�\WFƧƍ;�Jv�@Ak
�`�X+�����P�cA�S;�r��x@֬^&c�#2v��Z��L^l�5� ���5-8)���5Ҙ��0f�ڷ��ڴ��=Ƒ�p |Yo�D9r��5�Ef=�ǵ��ǲ3�Ł�l��q��Y�նz�T�o���k��O��oMJ7<=M�Z��`,̃.��G��$��K���X�[�n�����
gy�sp?h$���]�䈂'c�䋷�i�\�l@X�Fk��[��H�?��6<���T)��� ���GZ�N�/xA���$4<�����/�?����o�������쏟U@�#�Z�ƭ�j&����{q���v/��Y�|H"H����rrj��g�=�츮3�]7�{;7�F	�"	0��)*��$K�xl�=~���qX�Z~kٖ���g��ئdi$R��D��)f� H� rn4�������>�oZ�������Ս{�N�:U<ߎߞ^L�xr��tO޳���;;2� Wv�Ҥ��>t����z���j�&�	��x4F��,��E���KƄ8Fˡf�9ڵ�-*�X�����&;�a���>'n�-��ժ� @�7��p��kf��5��,��[��+���غ��5�]�n]#�V�&S��F-w�8���!�Na8O���A|�st^R>�x`�i)�
����Ph�M٪��~��l��]!�d��k�1�th闞��1w!�a�Ԅ5\��y��/O= VX���h�^��F�5��Њ�_�@�A%�G�?��XV�4b��Xh��Y;�UuZ�B)�V��ޭX�����]TA�!�'�ꪫ��믧����I�Γ	jT����(��q,�)���mx�1(��ȱ��E]���ӳ�2�<��<�螼wA��l�59�cp��d��Ό
�$3tz�-[��������ر�6m�(�Y�^�T:ƖS��������MW���f#��z�$e�z����k�5����~_@�t$dcF����kif:'@�ۇ�S���T sӭ�-C�lD]�ڍL�M��n���vkC	���5��s��,�Q Q*U�i�jǾUI��y0��q����j�.-�R �)�q Xmo���>t�B��X���#[�����$:@�#_�.���0 =� ��ڹ��|��&XGx*�4��ֺ��£
�oB!�v�d<j���RIV���?WXټ�A+,�[�>�rQr>���K��'��z�z����r�f���L�N=Fo��:m����|/Y�J@�2��H"dn���0�y!�ȱ�۟|�I��s�'�Y<@��=K�5�D����ѩ[㱔�d4�$�1z��+��zg���ٙ�+�QWo��GOS���NjT7�'p���޷hF�.Z�����e����[ǥSm�I��t�ƍ�qf��:i͸a��X�����pw���u���n@�� U7�r�kM7,=��q�:{��v\�
��$�l���d�MO��E�x-'S�VU�c�ծ��ʃ���[�qf�B�� SF�T%[Qw�\&yK�T�?P� �x��
�%8� x���Pv�P�����<�E��"���j�� u�����ܺ���y�dZ�<B�}��s~���������K����QZ�fmy�%���G��W_I�V�.�H8�VRR�$�LM��i+�O W��b�Y�X<,��
����8LKV���l���42)=@�伋�,D�W����i��	?,�]���ͽC������a�F��蠴�P���o�Ca˔�'$IQ:;��]��x�����}�Du��mtv�t<����"KHL�3��fز{c����IQ�Wo���4mc����a�]��Uk���[mF4�q�P���PD�:Pjr���od5yc�gJ�b�^jg��+]��&V_m+[V�ܝ��K0w�mc���(]�ޏ��+Q��� ��)��! �€{("��Aܿ��	�-_. �,~��q.J�&�)�-,p(�k�����u���1.>�:+e�&���/Q���
`�A�>���k�40�^z�+E�D�b���a�S��٩i�^N��9@�|�)Z�|%�[��~��Z��"~{Bt���T<N��<e:;�����/�h���E>44H�:�9[����I���w$�p��O�B��'D<@�d!Ҋ%c9�g7+(�1qXbl�����[4;��x+ܬ�#g�M�P0�MN C<H�J�^|���������geC~��?���'h,����^�Ϲ��	 j��{�9�@��o�[tf�-6�V�l��Z�l�g䓤�&Z�������f�e]
2�"�����pS���䬹�5Z���n��/Y+D�R����r�2�i
 ��ĈkN	��-��ӆT��j�k.����a9�k7�,X #\���t��i|[�S/�z ��z@vІh�@�>��Hr�o�I[�n��"Ԯ33Yڽ��v��6�z($I�JA������4��C ��de�Z�����h��7���ҽ�vҎg_�Q~�P�����9~��i�+qGIMHHj^x�9*�<~��������4Y�SB�]�G�N��s��;����:z��؂������/�Y>��o�!Q
E�V�+]�䂈�,Hlˮ7햍R,��R�"�α9��%j�pHX�J����߅]c�Ȥ� (�z�7yX|C�Oѣ?z��A?=��W��I1O����*��
������G᱊�IF�j4:=C�X\2�� o3j�Hn"�4��k�c���Y��vѫ%��[c��Lp��ͯ��w�����q�Wk[����������V�ޏ֨+@]-_X�8O���ư���Ni1�[��^����HT������0��(q(k�J�It��@V:�͆w7o	�s�����~�~�Z�L=]��g�J�)��u���r����o��:����K#?>x��<,�h8&�yA�P�?$���ό����b _��O�Y~M�b3t�,{������K�K46q̪�k[�'D<@�dAbY���Ƃȏ�RF��8o�	ʱ���2o�
GRizjV6LI c���;ʖ|!�5��Ѱ��Z�:k7��8���]�k�� �t���M���S�?��M�>��*z��f�s7hB�S��e>a���!
p����!�!9��^��d���y`^Μ|.�»]�M��[��;�Õ�`�86��-g<\.r���:�^��G�:��c����_`㹼�����V��NXI�c@����O�<)nz-8#6����4�@��Q�B���k��-�/�s����+Vс��Ҟ�T]�A�'r�x�0gi��V�-��L�'�1'Ϣ�xhX��wn�R�N�3�دP�g��A��D_ B�/[*5ff�v`<���螼gA��/~����mi~b�-9��-�I���?�{<������H���2��EbQ
��4�5L]�`��b�,/Kf:\�J�����;�ŋz(7�ы7n�[Kb�ھs@�����{j�����Yz�������3��Z���luek��]ƥ%m�d8���s��Z��r��J�GRO���i�*	���1r *�l������ x���U���QW>��x� ���: NT9���2^���G�xd�����B ��B�%sZ[��z�6u�7`��z�������?��?��ق�,`n_���4xzHH~�s�;�7��L)%y�-}�l<�=BRԒ��܍ [�>��F�+�_����a�!2
	�l��l�=ݓ"�{� ፶:6lX��|�_~ИmT�yJ�['B�).d��`������~�wM,� Xy�Գ3S�J�*._�j'��st����@oZG�?����uwt
��.8��nQ�Sw�[��nP��A}�����D�7|t�oU��k,{�K^�кru��ziݺ��v��w CmO�� ����u���#�.e���z 0��q�ޝ��+^s"�M��pM�Nk�,?~T\��RJ��_\�Q����?<d��q���^
!�-���%p��hzf����@���H( rC!%Bu��	�f]�#]Y�q<�B�W
[�Q��a�kٖ��ū	���-�ϳ�=�0��'�&�ܦ9��Z`l�؜5+���U���ё�p$H�l��XWc�^;sIu�����~�H�*yc�J2[(d�˰�k�@.����ѹejnZ�SAq~�����2?��nV����3-�k�����:�f�k�7Ɋ�����w�����z}����4��@��
����RB��9�1�0��%p��X�;�k\������T��`�P���V���)u��tp �Ѩ͔;��j�Ůk����IƩ�@�q5!�P:-a�<#h{MR�L�/ �O�z�zMMN��1>Gk���8��y�@TC����-�鲓��)����L�=�+x��!+4�1�'�E<@�dA��x�j�Z$ �}��qq7e�E�v<�z��Q��VZj��~q�bS�K����F&2>K8�Ô�E�Ȥ�x� #�/��4�a�9Ǫ~��67Xji����;�>�>Lw�N�s��ݞw�:�Q�cw����Z��DE����2h)��(�d*nf6X� `XŚ������+ ~����������67;��/LD/|?Hr�g8n`�b��>�n��]�L�|�>�9���3�N5D�3a��$��;<�+����b��]�e\�e��Յ�j�,���{B�sߴy��v��)�͉҂k�w�(&�`@�Ϧ�<"I1*9"͆�tH2�C+@�|'�r���'D<@�dAm��l��cy��j6�9rzf3hԪmr�c���GM�n��ʹS2ѕ�L,S>�$&�%{@$|�v�V��*��d�(⿆�~��u�k�����M�+�1��&��=��ֺ��T�r��|ݱw�@�w�\��tl��ݵ��r3 $DK�4�� 8���b$ʽ��K2�V9�&���ذ�U����׬�]o�!�1g 5@<8��;���Lr7o��{�����6TF�:������Np���j�Iwp��Os*�
4���._-�P&�4������(q��N���[��[t�]wR'�KȘ/�����~�|����ZB���V-K�a*����ӆu�������4x�9q���G�(y
M+$�=� ��'��y<�%3؆����Rl��$���I��fK�� `	p$��	�RkH-6��B!GQ��P�c�2�V@S0М:y\6ydc��6��YA2��n��r�[M\�(c�O��p���D(J��kFy\q��mk�MI�d/'v�����9 ;����PK�ݓ\Ig܊��(��x
�����@�1w<'X� k��{d��up,q�1B�Tq=|�s����vxX�������2ڡM.����=39!c�^�R���������؈d�/Z�D�0$�A)@U���k�TE#]s��ŵ���@�z�n�kMK/���>Ip�|f��2��4�D��x>���r��������M�λ��GJ�!��3�Ӗ���K���L�T[88J�|�Wx�(��h���O<� ��'�x<ҪV�v��vG����/���EdږZ���e�	�g���|����3�L�PD����C(�u� �F�"���x��Q{�J�u� {�n  Rt���O���*��3���4��<u�]���0&�Jk�!p-�g�P+\-}=���v����w��ݮx��^7'{�E6�&�q�H�q4Y���`4+])d�Zԭ��mM���,�Q����X��K.�ca��z�߰�q�s��0�C�,s���,���܋6�Ar*5�O��m����)��ߚ����N:68$���/�g],�N:�t�ڴ�`�s�E~��>���mt��J~ ]�)���w�F�_�~�v���9�����������	:|�(����{O<� ��'�V �A�l�[�n�-b�_|�&���h��,�7��E;w�2&�.}�����������䯞�n���s����˷����/��\*�������ϔ�N	�⨠���۵�מ�vS�*�*��Xn��/�tl�j"j��ֵ�������J@�>��J�5�n���#.ۚS8 2g�uN�����-��9α�J��`	67�"���r��v e<C��1Z��↫���_�9IJs����o �_�b�(�j��rP�?)�w��W&:��4)�x"��mO
�i5�BC|��з��99��;ߕ���B�V��lV�PF�g�c���/�?)�	%<P���h�Y��A�S���#�r6U)�/:��a>�t��7�Z�����Z��/��1�ē �{� ��X����I�36c�C��� �%l� ᨻ�G6jl��b��K��n��B����u{�>-IQ?���骫�!X�����(�RQJܔM�:59J~_�V-_��\M�|�ʼQ���$9���Ic��uus+�i���M��jV�Nͺ�Y�r��AQ�h'v���^4�O���G)W�w�<����qw�^�^���(�ntSm�a��9����S�U�]?�KZy�amk�9La�C������5���$9���c�Q�ߩ����e֫�l��0xV�X":<Dp��r���������L����	������kBu�5�=�q� ��tQ��Y�m��&�������r�*
�T�w5��Wl����'r�A�/B�xr�tO$ͦe�b	�R.�E�%�/��2'�da����u9ot}}��>�����}T��2�Z�)� !��-��n�Q�E�ʧw��7�Dbh��I��)I�
��}�#��tvс�G蝽"��R�}AL�9"c���N�s���+k{U��1�]�U��i�� :�WEb~�qxMzS����$3w��\�v?ʥs���;���h��=�#��(pko۶M�e��4�������n�:)/�� /��R�;�'�������hֳ��2.,}m�J��xW�$b-�J���A��R�t�8���(^�`4A��;��f
&���x�9K�K�R�-� �C�a���-^�'J2ܡd��<x^}}'Ba�����ݬ��V���'� #$3!$��;o���o�m�*�Y�\� ݓ	��͛��t�-,�^��a���e&u��A��z�7]l��v~��IL�e����'>NI���zX	8xX����yz�՝�jE�o���:-lt�X������^�����c�l���6���o͹���l2F�u��O 6rX�Ƞךw|p�Cm�v�6ĝ� �n��s%X:77hk�u�˵�V�gp���G=�?��U 0k�U�'�ns(L \�  5~c������3��� ��3�)�T2���o$���E��Z����7@��\�Ƅ ����޴
\����AA�u�9���D�>���l�\)IIٙS�ZX샧OJ5F.g*��PRP��1��q�]�?@,JS㔈�BE�jI����(egr�l�z�?�!����磍ǨQmy�'D<@�dA ݒ>�h���l�+V����O(��.��X:j�cRZ���# 6_�j�h�ǿ7l�DO>�K:p`o�1��C�S���K�J����C��`�U�jՔ�a�6Y�a�r'�0l���]˭������p��dV+@��.+#��.?S0~7:wBZ���e�����q���6?��NxS׽*&�k�RWo����# ��Lq 4X�8 �yxV�w�3r3�c �\?�0W�<{X� JɌwZ�$�Y�#V����0��W����q8�y��F.��9���v�
�s�r笯v��:�_���-]B;_��՚��E������ɽ}���{�����۴%�~����-�z+~��)����Y�H�{��4��;�7B������=Y�0����_HH��dGB�>���E���$e9��>�~���Q�3��Ɇ��w���oڐ����@��<4|F�F� 0*f��lg��+���c��=*;��sx�� A�V(
�JR㶘�-��o~���&�[t��	)���/����C���'�q'ٹ���V��Ν,�Ob���;��Ϸ��U�����{`��!+��c�8��aA+'��7���N@�A�T(_�4�P��o\����@��q�FQ��:'\�Rg���5����j�q2�a���T��wJ -���z՛���AJ���z��<�W_}5����>�)�õ�$u���e�tl�v�x��n��?No��K��T"I3��R*�Q��sKRY1<:&1�tG'=q��oHP�<W�7��*U���'D<@��=����ַ:*�b nXXgEPGG�e������,��3/��-��"�Z.[�Ǐ���s�Y�[o��n��6����/~���j�9���������H���xR�����iJc�a�H0AccTak��V6q+�.wX�)_k�w�`���m���l�ŝ/������Wi��Ẹ�d*����8=���R�T���lɼ���Q,HG�3=�s�7L�O����δ����c��?'�u���f��U�	rj�l�|��`��'$ʊr���k�;���l������Z�6�s�kY�]�6���z���=59�&��b��z��s�d�c��3]�2晑�4�ϵ=��*N�ĖB;h����,���N�]k
c�(<�k������f��낎����f�S��ﯽ�F��?�S��x�f�F'&���G���?I��_��������3;��8_��K��\�c[�"���y,��^_�B<gԫ�2Ѓ'��s�W���ݓ"�{��f���>l�ب<"�;�������UKG�C���ܹS\����e��� C9�2�"Xr`��x-8Ņ=�/�b���N	(tvfd\d8���BI����]��t���B��*Ę�3�l6+��HrxnP,�޻W,vMDS�h�;�)��͚�zu���Ǹ��̍!���N��n:��R����Ķ��6�:�r���C�\��C����s�=�V� �>�G�߰v5�ڈ��Zh���%#��W����R
����;��d�>�t[k�����D9Ͳ��&@�\������������ ��$v�g����o�SgF�+�?@�~�v��Ř��]o�G}�.ٺ�&�'�P� D�b��<�Wӓ��||�G��7e� �A�`Gg�(��H�\A}��_�R���gG1GϏ��޽�'��G� ݓ�e�P(b�"
�l�a��U��&��ϻ�{��ɢ�����J`�g�D��[o�I������*>s�֭]#���7wQ0`��9����Ա�ϖ���7CG���I�U������~w_���&a�EpF��ƤZꎗ�o����BW�v��g�S W��5�Z�q'����1�S��h�ݝ��m�����
� ��ƪ����	�)�@p�����T2���	<mc���&��<m���h8�F��.z�'�h���'�	<W�����p��s�q�6+n���r�oL��1�����￁�%�Ʀf@u$�?����K�xTB'?{���l�*�� ����?i��-�;A��鬸��	�dg��g�;T�6)M���+�c�N$)��*6���������V@���o�"G�xr�tO"v0i��M�X��P���J�{��x;q���o�#��H(��
8�׾}t-o����K�=�B!�o���ǎP"�R���F�$�g�B���Q�Zb��$[�l�U˒��r�� ��N*Ζe,M��֮kJn�=Å7�����2 �`�%S�x�����-[]�u���u�縭}�g�پ�{\�[]��c�Z��r�Zu�+�� ��p�� \�P ��|6���9�=~�x�BV;�m޲E��:��0���u�:B��kz��0����dh}9�7�X�x�|-$�5�)1����_�?���%�/KW����1���:�U���������\�x�&90F��s]q�V��?�"�o�%t��7S�X��_w=����_�Eb)�6ge1��Uc˽L�`���j�:��⧞z�^}�5!�i�[t��W���:���k����'��G� ݓ
[���w�ɜ6]��?����;l� ?l�)���^@�7d���L��2iz��')�����7H�,7l��4\��o��=�3�<C�b�.�h@���<�L�K,8 �Of� ��)�&c��z( ���Ԓ(��0���/�;vP�A��c�,��>�-_�����_"7�N�v��K���%�?i'ƹ��t7������n�����:��������L�|���<q�>t��9��Kd=�}��π��w�b�gi��J���?�u �"ܢ�t�K���H��+h�[u*B��ׅo9O�O����>Mo��� z�����ޖ��Ԭ����-_�\2�7�_/�ƽ����ᓧ�c��7$����~O޻P8�xl��41:I/����h�R.�p��#�u�կ~E�7mB\�s�{r��tO$V˶��(~�٨; ���� [ݰ��Qc���62�Tҭ�R�$3$�Nl��S�[��gw�n���-i����$:9nrX����Xt������tl���^�~bÎ7�,ӄD����X?���~��d���z��;����?}�c�R�}��]�Jc��vw:D�q��ݖ�|�w��A4���L�`�Tu'�Iy��.��Ѷܱ M�����o<?� �(A^+ܫz/����7b舍cU���c,e����rWo�"�GV<�,t��5����{(!���h�H2#+l�~�M��;S�LW�d���Ft�� �yZ�d@�_�z]w�5������Oҥ�7�~��;���w�}�������M��>6[�u$��R
oD_w������1`M���Aj���.�'/�~94,/�ݓ�.�{�a#�e�A����l��jW5�����l�(�1IP���C������*�+Eʠ�4��ykՊ$$������F�#�
%����Z�b	e�����j�R�z�!��\�o2i ��/nx���PwV�%6�v�3�䭿����|P,�0�Vڧ?�i|(%���ص�<L[[�*�i\!�.��� ?��:�Lg��۞�ߖ-k)����f��ۖ�Rq��XWԃ�r&̀�{��d�#+����4��F��C�#I�({`�[�IF��P��>��Z����YMr#�d8|v��W���~IT��嶲��FQ�T�v���>G�2�� ���K���ҫ��q�ѐ�5�9���
}��	��S�I.ބ��x���3�Ҙ����(��,�Z�D	���-j��
��{��U���B��O�ɯZ�<ݓ �{� �D����S�K]�C�����.�o� |&�)�ۖl�l� Dl���5c�a�Hl.�2�=�|����S?�A`\ʫ*ee�Uo N����F�v�/u�Ţ)��,�KΔ����4q;�,��n:��nw��OUw:������t���w���Z��&��z�@�TM��Ys�ו}͝,��r�%����7ԝ\��! }�v��$�����2G���� ���t 2��Ф��]�ַP�R����#�9p�c^X��}`�}��E1)ԫ���ڤ:~W~Vh��7lZ��V��0�Cq��{�r퇎��bb��w�d�c,$���1��g>C�R��}�Yz�?��G�����VX���5^*5$�29���\lr-�����V�.z$y��y�=Y�؍�r@�Pwz<a���@��mAqC�ŝ��	J���w����Ӽ�"��zP�j[s�������~�tU2�W6�v'1�,�f�Wʕ�;�1�6�: �2�^�������Lk�Q6��lY��\����6;��jw���q�c\w���V��x���t�%w��1n>?����owM�����8E�Bwz�O��ɘ(_�k�~�u�ёC�h|dT���*W��x��wg:C'k��%��(?��-����`�Ń ���1� ��l��I����v�x*I$�2��I�3~o�H&'@��}����
��PpM_�F��޷����R�T�c��l��{�K�Yr(�x�����w�BRoD��� K��>���d�C��ɞ'�\ � ݓIö�z�f�B1�q��ٲ7+�έ6Ũ6:P`��'�)c��'��xv�7C�F��z�ħ�}A�Y
���P�a,v���0�6aY~c֚��nKh��EC�ܥ�$������h|^u�c���/w��ɚ�,l��|��Pv4���v����ݠ���d4=G�Y��k�_���7֫ƭ+_�g�����q�����1��{N���`��$�L��n��fn$"�Dr#�ݠ�������Q���`A@�Z,��^!�`��À[.�bRo:�n�1@:�a�xwR��ķ��XI���L7�Q��4=5f%�ԑI�.oՒ��kl�wuw�8p��=����Xq w{�\�$�|u�L��
A^r=0O<9���'���R���!7����}���)IkG:��T.P8�8�f�Z`Ǣ�.�Kq��5���y,��r״�%�cQܨ�G{�E��SY)MC\ܝX& 8��sk�۱m$X1h[Ow[S�����?pNL���ow-9D�j�B�s}~�2=F]��v'չ3��u�:�^s�<4y�+�%Y�<'D*�vނ����{�@�|�*��G�]��hkV -�"x��u����g����g�wDC+��&�i�U�P��Mm{��+x��)��w�F##�hyR� 
�W�_^�-e�C6:�N')_�:V|YB2�J�R�.fK;�'i!��h�����u$S��%,��oR~�D�8����C��[�x(��ݓ�.�{� A��0���,blܚHnll������]�VG�26�D2&�1�_o�+�����mh8I�Z���[�%�4�
yJ�z��^�����g�_Jq��Ξ��s#l�UP��v{��eMP""�X�}��:o�w���[જ &�2���݀�]zq'��q�ou��O�S�WEi~���bא�(.�D-m�<~k�=�c��Ki�w�u ��xR��-־�ϋ���r��qܕ�\C���Nvp�#����qڔ�����]8q�(���AS������0�ې��jh����u�˚
�R�I�����u�n��,Z�]U,jX�#M���Lͻ�ՠ5�.���Yi�����$��g�彃�������@�n���.�(�Yow+�&����^���+T��( *�:�������=Y���j7�u�L:�l�Lŏ0�9�݈m�h6d >�ovufL�3\؍:�QK8���M�>��\V � q\��?�E�z9{��|�gRs�ƅ��m�T66h�)%F��FX@�m>��l��p��~��,��:��M��]�� ���&�q'ɹ����Njj�+ kL��%N��j����YTA�,y��U+~c�5�A�m�Jp���P� ʰ�q���Ic.Hz����n 6��0&���y��a�לX�x���@֬]+�¿Q�ny��I��¬��	~��љ�'��L�m��I���+p��I�v�����h9b 1��L��/��/i�����=gF'�<HO>����}VK�v>��ϋE��O����~��Lx棿q7�Z�����������E/����=Y�X��]��_�he�R��5҄1Ul����X&�]�H��X(�� �e����0[Y-z�G?7l|��N�_q������	���G����a�x��ys���U��*V""U�[��ni��¬,ԃ���Y�M-^\O�˾_�&�n��0�e� =��|>K�f»]����It���	wj}k�\����
�x�3j��ŭ� ���M�W@�0�SY ɋ�R�M��od��,kX���f+XG�ˡ�ֿ���e�u�ȫ�q�\��� �7=�k�:&���X��r�\?��^���[��饗^��)�R��J�$ʀ��Q�����5�;{��1�S��]^���>��O���I:�o?+�Q���nv(*��C�v������^���d�o�d3��g�3}�o��Yy��J�<� ��'��ZMq�wuu�ҥ�9�28����O�GP��n�ի/�x�׿�u'��  %ݑa+g5jѥ�]N�_�Ԁ/_eڥ*�Z��f?[k1�R�$�P(G��x��m�$�����
kS�61�)�Rb���Z��AèH���%��rܼ�87�B����qwaS�\c��:7n/J�Ŗ�o�)���*�ZNC��q� W�� 8(Q�O�igػ�mt>�q�wƅ��5X� rĎq<,n ,�vHhp�*J�_ K^�-o�lz�
��"�e�[s\��`Wap��;��6�cĥ�Ư���ސ� x�Bb�X��h�ʕ��?o�?����?J�����{ĭ~�ݿA��즙�I�ꪫ(NPWw'���� M��Pb�.�zzx�B|��p==���;	��O<9���'��
�K�6nX] ���96cp[')��'>A���/�bG�2� �����K���M��J����J&���k�	�U�R&\���͛����=;��?��MP�aʻ*�9�32���[��ycGs<l,�p4�ve��F0�o��	L�Un;Ip�RQkZ��N-mu㪥�q�|��o�r�-�%>�g��R��)��
���s}`���0����n;JK�햇=k8 �R������R�Rn�:S$�� c�Q���$1�2��ʆ&Ժ	nP�Qg��B \-��IRc<�9��:�g�2nh���i�@�l��2<�D��[ͺ�c�R� ߑi�g�[�Z�d3� ޢl�H��v]y�մd��z������wR*�A=]�T���d���k��B�n����o�L�TLhi���)��^)V��(5ZU�VJ�5�>�9Q� )��}�֒�O,u��!�p�̰59=�Wh���'�U<@�d!b7m�lJ$���VTOO�l��6]�H(L��چ���su�!�Ѭ
{\�Ae�[o�U��O}�S�@��UT�M��瞕����V����F�����3����	 ��9�hN�~�`�R�ʀp���E?u%�y_�bԢ>� GK<�  ��IDAT=��qmP�F�l�RS<�S,�$9�$uHJ�ڞ�l���0����ĸ���>H���A(Xw��İG�8���2�^sb�e�Ȏ �-�jK�ꍒā}� ^�@3�Z] �r2��ՠ!��{�"�oD�&e}k�x�r�+�_:�Sp��W���M�X�~�~�l�Y����}vv��;@�|V�E���Z��A'�?����}�u̕�%�� G�p��Z��`L����9��B���CM��*+_>>���n���xԄ �x}��s7��9���UkR��
�w�������_A��=��WT�������1~���M��]���gE5b4���NӞ���K6Q�.)��sA�"(dA�l͓"�{��;�t*��W�6�U������a�
�L�/ܬ�ûڐ���7����=���{����젩�1� �R	��ݜ� ��kW��y��!���W,���P�"� ���Q���u&�,(�����~��1'�q�[�p�la�"˹R-�\� A\^Cڒ�=���9�����UMZ���9��4$`!9�_�SW���v�d��$R�K��"�����
�6*$��b�5kR'-�5����5����+�A�B��Ut�����}o��e�&$�BX�B&�ܬ�R���xOغ.UK��ĲG�"��%Ȓ*���*�k��2��uv�H"%�~�gg��093+��Cg%N[�H��;	�OZ�"�.��3�~nEz�'?�G�x�*��*�Mf�?��(d����~@�it�����*�����$�y�(e2ݴn�E4xj��ŢT:!����x��M�w�<�����,H�ʵ$93I�O�hP_�Lw����;�r�jZ�~��l�Y�o@n�P�_̠T��G��c�8~`�2�TK�|��8��� [�*�Xr=����٪l:|�!4�i��\
�vOO7%���Ǹ�m۶� n��7�`�~�t$%�Yb��S��u��p��w� E�a��L�����9�<�v���9�da����`$((M��ϭ�El]�~[��xHx��I.(���c+�I:�Yl��9�Eċ ��xxÀ/I�x؀5�J�k3虘|C,eH�Aߕj�O ��L+?�eu$�՜�@�Ȁ]��M��o��Cҡ�(o��IB	q�}N" bߨV0��d:#އw�?��c�o��ü�P��X�9���4���
+OexP���C�Z�y-]��:{R4:|�zR��G?B#�G��@�F����τ}��{������%:x���_�c���Z5
x�y�c'�K�?�` d� O<9���'�?dtәEm�nl�(K�bcE���kN�2꒑�5���5�V��J�ҩ����V��>����Ӳ��ࡇH��'��?��;^k��}��w__�x���tR.?� �-V�C?|���#t��a�o�<��G�1iǪ�+���!�p��b�E���$e��0�X���>�E �@[��)9+�ȴӴA�R��� ��O�Ib�;�qM*�y���* ��%#;(�{0�\�&�P�xL�G��4,��gD�
�p��B�놵О���.b�l�SJV���(Y�����A�
��Ʉ�7��nHKS�������2?o�+��C�}hfrBX٠�4$ҐrDQ�n~�Y(�ihx�����I�<*"P��OIr�����b���Ӱ"V�	@A���������+E-�&�|N8ar,��+��Y^s��;��5�5�]Օ7�fV@����d���J�^y�5�F���(�	^�'D<@�dA�MK��X�;)�h%2A�9���.δ ywO�d����nk�?σ��g� ��������/e�D����:,4dH��;z�.�h-��2�\�H�S�vE��?��?����H�WwO�l� �:�Кe��{���2�#Ng6�ڵ� �|�AS:x�3�W�-Na2�5_.V[Ў2p%ө�u����Ը0��c�Í/���MX$���b����(�k��
�d��{�x|��_��&י�^�ZE�%��
K�������a��x�I��1`a>� ,�BY,f 2~GCAq�7��E�8�Qϖ�l���Y��QP�*�nQQ��(.�PX��|�,?�'�������2"���`m��(�����@q�� ��{��G�y��"�k-MT�)���$�X�8q��a��I�P�n��6ck?ϊ[,��w���*��xm���-���*+;}�������ӿ?�4=����QX��-z���nk��� ݓ���l�M��!�`*%�E������JĿ�= �}_�:tċa9��ba�ݷ�m�����/�"���K��.���S�pj�k���G�!��0`L��ҙ���A���*��)s��7���q��7�.c�F�k�lP��<��	�v��-_7ܶRBf��/�����8,��5�P�p�K/�v�Ԁ�s�L���6>��U���dѷ,�&G�Y[��2T��J�ɢ�
p#d�j�%���+<��o���@K̀��X�-#�)����ߠX�p��u�6*��Kh4[Rڅ<dv�
 ^�BMc�W���M���d,.��OGKѺ��\Wa0���OA���s��̦=BH«�����ˠY!�@P��vc�)�;q�f��@�@[�5�!���7��Ò�8�~���9ާ�T7�����/��l�w���S�*�"rEI�C�_��1���6�4�	���[�#�߷D�(�����N���5���X�N�'��� ݓ���o$��b����]W6XÎ��͠=}fHb���S�nW���1��}��ߧ���tzp�z�A��<����s8�1&��d:DA9}F�P�[E]�Xuh��RWWMLOI��d@�V�����+�7k�u-��ף�.��Rⱶ��Cn�fk�&u�dW��X�H ֶ֬�5�9 #����:j�9&�f ���^Ӛ̥��t'�qh!Fl<�U�$Ð h�֭]N�|^,aű�I����|>Z����,[�߇�8�-�φ.�89(u�蒷z�
Q ��J�V���c�T�NH���U�i�����0e	I��H\��N;NO�x�,^��o��V�x �0 V�п��?!����w�y���A6����ij6Oo��G��Y�D�4��]�D!��5r�x|&��xX'������饗�W^��nZ�%�w���}+!VLg���o}��������0� �CJ� ��4�5�x�%�8��%K$qtl�N1�OL���c��OӒ�U�۳�ϯ���T$:�u\�����,D�[��T����HxJ"��V����X�϶K�P�������$�	a�N� Ha�D���AGeQ�"�D���6ܯ�XR��~
 �a6�wl�dhLSņ4��`���-0Ŏ����g���{�b���7�-7_�N΂�^è�f�lߡ#��C?�d�+V��̧idd����L-wgG7��w�~�Q*�%{�7�e�o���6�QlS��y>��������]�{��R�=������N:p��d��d�����~��l�'��X*�w�B|��]����|�v�m45��l!Oݝ��]2�A��/�Bg��h��e����1w�	�����~��z�@=[�o`�t���%�ɢEKx]2��_���x�q�)�|�et�%[�][�V��s�O�)U�MZy���'����.
�T��T���������z����+[��R&/���
�m�7%��4��M����/
D�P�(ItH������h2B1�������]R7/��HlTyν�cS�{�a)ml�ZR��X�5�m��XN#g�����y1tOοx���BD�Q�d�ޗMd ��q��NX���%�$�	Ԭ��E^��H�\K6�m:���J��o�V��E�M��X�am#�J&EQHD#�M`�=�a?���띛���6��T�7)��I����Ufe�%G��MMy��2P�tvI����>i����D���ʒ�'s�{D,���E��:;��l���'����mI�~5�@H����.�Ơ]�y�x8�mX/�6|v�v�B���<��������u[.Ƴ�t���s�Je[��*U��k�;��o�*Y3����� �����7⽛6m�~�p+'i��ި\ ��
�5��:���{�_V�QQ�&tf������GB���7wʽ���(4�z�-��L����h���W(W��~��Q��l�PQ �	�@#	��5���D(B>o5�	}�x��
ڰa�x�6�o����_��dJ��9 �F˰�S���ߑJK������JE���n�5Y/S����s�����K�"������oyIq�\ � ݓI��-�am!m�i ���A��On�m��4o���2ꏑM&2����}�h4�@��Z�Ir�naQ!3:������t���il�,=���t��i�z�վn��4з����ĂW�Y)�e�>���a�6UbЍ
[�h�a��7v�v{�-<+|]�	�|ߥ�腗_�Lk�S''s�n�f޸g���Sgi`�R,��Hi\���(g�8#Ih�P�V��d�5$���H�ҩ+=���9� ���._��g3�h��u�b�~��/I���-��7����X� �����ٻTz���b��`���Q�Ҡ��%t�M7Pg�b�_�L�)-X�"4:q�v��K�}�q�����Q �`�KQ�a�B�4�;xB�������M���| 3(|S�;�y����J�x�:�h�"Z�j����"�Q̗��^��IRgG�^����t�C�9��t������+.���I���� r(s(M�W ���V�0���n�X�G������v�C��͐�P�C~~���NG�p���Q� �`���+|r<@0�t�� �唒��x Ȫô螜� ݓ�4�j��ʆ�������ĔNUHUZs-D�Q
,\��*IWp���X`��r ^r�܋�[�s�Q`�(R�(�Y�Z��W,C���$^?:>&1r�b�$YIY�.�������3b�(1Ďa�J�)>�932� �mۯ���)��9�������GJ3�2:<�c��d�pI�:���Y&�O��L�Ū���c6K��6b�]�X�P��q.Z���G��Y���]D��S��|�I��|+m�t�(E�b-����AɮwP���^B7�q��<f\ұXT���&fi�P�m۶�o���Q��� @!�V(AC�9I:�x�t�o~J���a,⎾Juw��	]{���{?-�hQ� ��*���xv�b3��˷���={�h��RZ��W��ý���hl|�b���*+=C��;�g��7���x��{���zy��\��M�>Bq�;��=|-tM#?�fg����/ì���f��=_�R�#e�<%���v��(�UC�d[u�vG"$\�i�6n~[і��2�vx5��Oηx���BDʩ�������}׶P�":ݒ��vS�BMwS\�`��;��b�lZb��
A���?3�"nZ���
՛����* ���q�W�m @�4q<�8&�,�����5[b�5��&e�@���|f8���#l���;�u�}�EZ�b-��{@�}��	ڲe�Wud�,[q��l.O-u�i�ԉ��,���R�-R��c�gF��Xe��A9[�Ӂ��r��C���&�&h���⎶�0�s�(Y�M����^�����*e*7��R��h���.�s����jVxjG��3�K�P��{�շ��]��$-_���}��5J<��?8<E���k499.�y���4t�5^���6m��m?:v\�+3S��� ��L6G����LO?���C�����*%>n�	ڻ�8�H<+��Kv�B��.	q��!��"pP�9�=j:�����W�����m��D��M�-p�Zo�I"%�:�@AM��0����	�
S�\�$Z�N�Q<ȊYW��;+�@� �f�&<QB��D0�NZ���'��o� ݓ��g��Δ�n����:,r����o$}و�Z��Q��>Ir��!96r�p�"!���b�(7�����,�T`++� Q>'�B�a�Ih��oI$�ʀ �+��P{��]��v;�jސQC���&}�[ߧo~��R�� p SY�&[�/�~���F{o��CE���I�<�����[c+k���aV ����M* ؎��dgs|�M�d-��=��E\8P��w�ƍ45��&"�&�RZ��赝oK���̔t��fe=���M˓�������$�	 9��`��c��� ��/��=��<߂d�/XD����?"��X	�Ύ�_�՗Yiu�(cKf:��@���V��s�Q��.J�%��X_(���3�TG���ɱ$��P@�c�N�:.JO�&�汖�7������G�֏�r9 Xk���^�΂�/B�8�;�4�U�9)}û��H8 ��+H���ˬd��=6x�0��~	Ws��G<N|���n_����,tOοx���{ް����?�B~ِK� �r��q@m��n	%(���GW.Բ��j&;k��1��K�M_�٬ś;���9J ��IM�Q��C|����m��_Z~�$�:��Ki���g�Rt\�A�W�Y���o�C���a�ǣf�n��ub��)[�9Ðǿ�d0� ��)a���m]�P�5*�*_.2�aE�������<F��TKb�I[XP�JO񀔕��	}��DCq�r�3X�ed$�	���M�V�������oG/om�j� �¶�Jf�P�>����cJ�Y!㼯�O�p;zB����4+E�V�����h4Ӵx� e�]tj�c�j�-�[�/�[C��"�e.��&�{���X���(n~��-�0x�a�<�O/�m:Xxe���>?Ŗs�-� ���P��� [ՠ�Y���GP�`2;A�**�]Р���F�m�T"Tx����9r��7�J[M�� ���y���=Y�����e#V]��*b��>@ +4�.�.Pd��	9��d%��A �q!$95�í�,p��[�$���rڜ����04� |K���E�u��v81	�8;���e%V���f�bC	Iwt�Uh�ƀ
614A�	_�[ZH����q�g��cB��x;��Z�����f�:"E,6Kñ��'�4 �������=B��kBꂸ|�^��fx�P�7>>%J�]/P,hQ�3-JN�R�{I�|C��w�-�nV��T�{$ �d�4幦I��;���k�/:�<��% ^����Л�� 7tzX��e�Iq/�k��xԴ�55�
fB43��ǎSO_/�-�b���6k@yj͂�e��P��Kaq�L����c4f7e]/꣭[�ʸR����w���X��R��� 㽒,}V�p�a�+S[�P
5����˚uk�ڛn��E�t��!�?�]��|M���O���		�ds���4�3�~�n���҇�=�߷�y�FώЩ�hz���v�Z��xr��tO$��ecsGb�:�2��c�Yp?k����l����'ܲ���!i'z�-��%�]N�>���曒T�:k0|�s۾�(�����=�w	� P�[ ��+��:�u6)
\�����S!��c����â`���B 1��N�ak�?�!������͖(@����&w:�I:�q�Mt�e��q�uJ��70���7hY�Zg4֦�d9��-	[�=E�*��p=�i�=�3$�	9N,-n�D,$D=�Y�Ig��T"��ǖe�ǃ�˿T4�x�^��lљkQ�/ ���$e=�`����#^C�1�����Icl5�T�g�So��$���u��2�t����g�}V����NnE��J�k	Ӟӊ9�rA����'����k�<C�$������ eY���[d>��iZ��'L{������Ŭxy������_#��fJ�P
���#s����ipp�~�� �ށ��tO.�x��ɂ6w��$���]+\�(W�����A���+�ӏB,�Z�.1(k��&���mt�w��eK�o���t��
D��[��=��|k�~i��@Y��ua}C�ݏ����(;���  ��/��V�	�ڭWI�b��_�fǣNU���E�fM���F]2���k���,��w8�Bְ��LM��@B�I���gB�Z�6�R�\(�6����.|�!���4�A��>�O�� H�H��ff�R�NFTD6`��S�dZ���a~���ʸu^d�Ǔ&�)`�$���5זi�L9"r�����fg(�Vw��)K�qAUx����e���Nw�4���@��M9W��F�(�I��4��H�zbt���;�g�jt�{����R3��`�RM��6�ox�pj͡���g��N�:a\󁠄�χ�<������zϿ�,�~���gO=M��w��\4�h�Ӣ��V�uW]I��<�,���~��.ɵ�A�kECԝ��y;}��oS��Eq�<����螼ga��|�A��?���������f�Iw�����/���/����/�Y��K�A��;b����D�:{���+�o�r�^�p�r9q�6���Y@|���j�[׀��Wu]>W�O�L�o�#�*=�� W��!Ӎ�n+��$�_��S�־�`��ҟ�ghf�	��� $�"�|�9�8`]k������0�|�
AI�d3�s /@�j���(,>IPl:�{�X樕����kbj�]5���us�c�l�2Y;X�Rg�{�g `�����J�ibr��#L��E2Z�J�Vt����.��l��&-�5Se
 �/I�ȑ�2���ER^���u����yxo��!� ��+n�싵	QFFƄ(k����!���r�B�H7�r;���������]�����A!�e��L��ヴa�
�9OA����K��י��Bގy���=yς����߸Q٪�w@@nw���o���_��-^F۷o�{ｗ���-V$ -������k��C?|�>񛟢���ߦ�L���ڵK@ɸӧ����Xx� ƄW�l�#�x�b��Jk�tZ H�\�#���k'���i��.h��ڊ�[�*���N�U!и�f�kl߰�ڮy <�	ֳV �&��7� zb=�
.��S+pZ��x0S�0�ឧf�t���3z}�
A�259.k�~|��C�����N���4}�Z 8*,ħ�-[�o:ΓX�H!׵��F�(�P�O��));V�ʕ+����xA�M0��N���������������G��s�o�xh����ҾE����>����˶m�C��Ν;�}E�/�k�v4�)I�˖,�5@�}2��	4��Aa-��7��}��ݓ �{��C���V6����a#�k4���X��+<ѭ��J��կ��Ĵ��ٳg;5(�/���/�w�A}=������.�x*���: 5��t�M��#����5�3����eLP4P�t��	z��]���j���Q�&�X��}�ڏ9�:�7�]�:F��8��5Oc����
�5�e�X�o��gpC�yX��N���R�  �g�tq/��(��k�R %��Đ�L;�UxFXWxF$��
@k��c� ����7:��k�-gg=��M���J�wY)sD�A4�����hy*�#G���W��k�,���IRc�6��?;�ա��3�s�h }�}�Q:��2A+hюgw���9+����q�g�ht�,m~�v��L�00��ė/a�P{i�eЛ=��Y�\� ݓ�,�п��6�� $|a��\� �K���.
��ђqOԉ?���Էh� 	2����[�}��t�B�����{�ivUg��|9�W��CuUwW�V��d���A����g�xl<`{�ƾw��0�x�����aB"��$�Z�
չ�+���|���O}�g����;�Q=]��s���h�+��]R��b���z�Fk��9`.(m��>H���c�y��	�6e�mن��2��@n���S�!h�3�!e �	a�5��&����aޘ�%��|1es�������vC�z}�d@�+�<^F���r�K�`����35R)�p.Ȁ1n�lg��NiK�d�T&˝���w�H�z� ��N�����:j�1xہUc�h;�_��╷����������Ӳ����d�k�����g���υ][��	���ɤ)|�0?�P�ݪ�^⽈�����߰a=o4g����%;=#���}2?�(�V��@��sIF�+�����{����::�et�vt|��%���eZ��Wn���5����3��X���p��>08�1@=��0�8!3
E������{�Z�܅�c�N���?�0=���}����#��!�sutu!�l��!P�Ϲ�\[k̜8d]m�R_����+X��c���y]� $�P'd�c�=ݖ~��vX��Ƅ}s��3�l
s�������;�0��E�Qd�8&T�}��m�b�0n��;��^�{�DR�mi�k�W1���G�.y���3���zB�&�o�?�0x���"�Z]P�=����aj#�
R�xsoz +b#�� -rq��
�q֭�x	��X<�xa���0jTa�]gg�g$��"�N�<!}}x�y����l\�ޤ+IP�`���ɟ<dJ��g�׶��?^*G.�M(��Я��j���r��.�Q�?v�8'
;���?~�t���	�5��%��|�+�xq�����f9t�|��?����}�a`�{��ˮ��
p�micNql��G����l�>,��ηRdz�l	=6�J�� ����mw3 ���-	?H	 ��}�х�3�,���?5�0�+�������jߵ��\pM�M�I�0�Ӝ~���'Z��$�">��Qv���y'��</�4��<���`XT� �׍V�����ǽ� �ix�s3���z��'�FMؼQ� �f������<@��F8d��T4^���M�ٲ6��x.\p�4x�h�{��E#X3|]�rz~*�5@ ,�x��G$�c�=�o(�e��#$��ڱ��@����*��!yp��p|te[\\����r��)��Жa����y�W�����u���(4�;{q������9������߬�fʦ� ���n����	�۽m����5�e�/6�/~���i�"�:� v��Q��-�$�~���o|��:��|�ӟ�������$���E6b/uI�%�9bs�!cJ���h�g87�k�殓�6��>6�%W��W��nگ�{���}ZAk���\`� x��7>g۬�
t��9-�����6��|{���V��FL,٭��a
�==}�t�1�u ��Jh�Ӝ�=�MO`�@8! [����(pA��À�����Z)	�k��8��{��[R�]/�;ɖa�����rǵY���À�����} y\�];�4���ݻ�u�S[]�	�)&|W�Y9��)�4r��0����(�HXz�����^#N���	���%5lv��'��_���iӠ���g"u�3��K/ȗ��^S�TV��t�>����������/�+蚃�t^7A F�T��L2�Qo0ɲ3l����w�#��{��06G�\�HＫ!��n��>�����g�zZFGG	L�b���`hГts������f�]Xs�z� 8z�(�� �0l���uR7��X̓�\;��ܻl%��<���[eJIs����es���|0b0OC��������kU�Tf� ���Bu��R��x� x#`�׍@�j���V�M\p���1��C׸y����>iZ��L޼R,N���iң�E��$	".�r)��F 캶�ز@�C��z���1��߃glט|�� �S,���<��јǎrm����Ǜ���p�x���#�BE�Q�6��ܴ��Zu^KM��ر��x2��3�����|��ߦ�8h�/�|0���e���5�	7L���At-�w� �|E&&��3'�� joh���b�g�Q6���:�!ǆ�p��܂LOM�ۇ�9�VG] C�2�������tx���<�-ke��:��>�|ȓzD8iɁ������쿭 o��\����zs��{k9�@ �3��}����i>�q�YG?xi1FZH}����P2��m^����6�����QA��C�Z� =v���n߹CN�8A�#"%D�50�E��y�X�0�.f*\�W� p<�"����n>�2�b?s�1$�5�r�:cȔ�mܰ�9���E�a�mw�����E%=���>�y��R�4_Q�(����_:z\�(�wttR)�H0�9@�#�m߹�]����S|���?����k�I5�R2���]"_]f^wllB^|������P4���
.;;ȿ�����*�G�IR��W�ZB�r�����!O%Mr���l��Jb#��m� ����7�R��9ZP�h�� �?U��Z_ޚ;�<$�
�֋��1�\�<o��wO���sm��[ ��Pxw��5<��WFH$��)��a}�����Ĕ��&vfχ(�A>���W6��مE�o�r˭o�?��)��Xo4���T?�VhZ�=@!�@0��놐<E]rYz֔qEY��M��Ƴa�+�l5�6E`(�����~�tQ�\({5�5Gn�|
{ �!; ybc~xs�v>��ǮSt'F�F�(���S�z�_��:�BI�l��p(�ү��y���Ɓ��ö�͆�u�Ú� OKr�zD �:���拍5�R8^�8r�)��q�&u�-�Hm]��F�gpp�:��S,��9 �5�iyJ���8������& �	�r�[s��m��
q����t6��V������� ��+�c��Y{Ŝ�b�	b�1s0�qХ�������n]�^�nT��L�z�p�NQN�>%�
�{��ǎH�jJ���6�5�|��JL4���������1xp/m�����8��]��;v�/��<�4��Wܦ#0�\��+Ȁo���)����@���oH�-7�D9Ԣ3�є��
� o���[B�~2�LQ��V����wn��sj���@�{WO/#�B����?����k!'�0�� s�dY�W��h6�.�/��ޘ�U���\��+��tK���18$9	vj8@j�J �8�$�D"*���-oy��f ���m�6��qL+ b���:}V���P��g]e�=v��َs%�]뫱�_�	�j�3�����|��[V�5k|���h%��i��"���w|�z���6�fЄ��=@�8���� �h�
�7>���)�֯���Wy����������iI�Z^u�����%N��i>h�kk82��{?�W�,Z�_�!Sv@x�~Ȫ��%���/��U	�׆띛ZKn����U�3Vp��iOp�G�����]��Vi��mV��!��n�,���@��n�^`×x*��D6_��06�����������Woe��J6S/<�S@2�%Xh�j��:7W��ꮧ4^Y4��K�� ��Lp1yjS�ddP�(�߿� m;o�5l�8� /�5���Ы�Q��;K�_-�����o�{�1l��z��k�߷[`�u��}���w�!�f+�{s[tx��l� =�%Z!`��M�=�<�{�� ��������]�D����3�r���y�69��1����<y�J�x�0L=��7�:�����չ�_Y)��j��Xl�2��
%�ݻw�z��5pıQ�������f�ƨyHנ��,|]K���:s�1� h�V1q(�z��x�L5�*���0\+jk<����m,�l�z�g�ډ���>��cMC7gݭ�£D9@�u��3�Q���Cx����dK���C� =��2���ʫͲ�uu� �`�W�0��?�yp��L�>�.����f���JM�א��̓Qo����/���][��6
a�gA܂j븜�g�G/��Uw޶<�R�_����u�w��t��G�&5�!�b�l` a��7ld�uY�ԕ쒜�x�Z �������D���IG@��Ȉ��,�T)@2V��t2�&�AKT0�	kzOY�\�~�6��½Fh��V �ad��?7`�g� ��#S*�=��#* �:��q��,�Q `1p[��k�0ܚ-y��d���xbX��qVv�\c�wt�K��KO_�	��S�C�����t�i�h�٨6M[O�#6�8��	B�W��]IR+���l,�`]o��0V,M����L̇�z�Qg��I=�ɕڍ`i�U/�j7mK��@ F1}�����l[[���0E�R5,h�G���^8F+��z���j��-�֠�����A͋(X�=�����A턬Gj<CޓP�A
��Q�hHtpTx�t:�y�K�=P���vD)���X�K��dh`�l��KR耇y���L�X�ujAO0�Q��[�'����Л����ܚ�<K� :oysH�bݠ�?48`*�\�i���U.Ŀ����b^网�̡gB����������1xL�]�|�n����V�9�ZC��
<;���A��B~^�=�k��>�lA��xȏ����1|@�ǚF �4�ɄQ�S)�ь�b!���b#��GISڰڳy�o�ES3B[Q��H4.����yE�˦[�-v��Q#���	�k��~�.=2�{��{��
���?��8���;����jq�~�VUaf��~mKU*��0�5� ���[�q^.�	z^�G~s^#z�����j�����D�Zq˿ԃt빥`t�f" 5��@����͕�C�RH����\՟w\�:!�eOB>1ak]ܛ�z�}�zyO� W�mfc\�]���-�s�Q���ԉ?<b����`}�j�\��5���B�q526����̜�-,Ɇ�Q�9kz�"�jl�a{�:�R���%Ϋ����Z�+:�tR����D�R ǳ�g�?}�T+�܌aA�dIH5x*%}�t�Q��.���ݿS�_�K6oޤ������3���_8)S#g$V#�Ts��Z ����s>��cM#��y0h���y���(��p������;�M���F7�����4D���_�u�����W��U��׿n�����������O�g�y�D,[�mۋ�C�Q�����o ;@�^l����f�0����䲰�;^7�R,����^QO�aIq���a�p�;���g�W�Wx���[���|ù�=["�Ӥ�!۽5�/-��@YԫC(�
�~�.1ԨL�ƚ"%1�i���*9z�;��V��^DUCI�4�W����+����E��C�K�(���֩
�0h��k������A1H����z��(W�sn�,]S���Y��H�d�8����C�F���TP
��L%ش��0�pm�@C6�둷���nC��_����i���~���}���H��?�+�5^w0�rR��r��>��cM#��	5v�d�!͛o�Y2�mfSv�}b�7x��y��g�ȑcܘ.M+���	���������n���У37��׾�� 
]��G� �06�����9�R��gIT���Qǎ�;�+�-�aZ|�q�z�y��y�A 7Xj��xy�&r�n����elm7�l^k�^|�-Ys\�<~��ф�i���[
�0�u£{\�0�Wn�1�v7���Z�����G�{��mrס�ð3�g`�z������@�.;��`�u��o �ϭyv;_��x��������$H+!d�;�u��/c����)׈p���V`�9lr�7n O�P*�ё���LMLJEA������L�kt4� ��q�M�9!E��2�gG����&���zi��ezfN��l�]ۮ���v�A�+�w�-�r]�z�yY��v���?~�t�i�B �����፾������6n�$�d�\��������>�zw�c�8C�P�;~����~@���:��c�tS�d&��������?N-�M�9",<5=aj˗W��i�x�9|o��-��mA�P��ح�������|��J#�vyk��Jt6��J�kU#�{�[�|���i�h�?q�ٮ����}�،7MϠA�Y0"��C��:�A27�[���˖-ò���r��Y�:C�`���P�s`�m�'J��.���nkV����`���6u�˙�V�"hz�AY��)5y��@�Q�L����RA��#b���z{Q;T���U#k��B��k�uިFNJ�����h�����^��ލ�g���Y��I{w��~�����2��FB�-��9�?�q���XӨ�kRU��-�bY��ݢ������m�2�A��B����t�b77�?������%�zs���	����Q������W
� �'�x�" a�{ʪ��j�PR��6��4*a��~����K�����5�L.N�<L�"73=I0@�S,���^���P�*��Pu�-J]vÐ��ϴ`;AeOػM=�)hx?�����������7j�W�7]�Ԧ4\�3��n:��n� ����3/�m-����e��	i]�#��W;>!A=č7� �>KP���֭[e�SgϞ�rY��|�5��F��l�A���|,Siz�n74��ѿ<$��ݿ����x���nx�(���=����W���СC$G6�$��'@�=��hRv��*��.9v�%�d��yۡ����)i��������28�U��y�#�n��m�d|bYzz@�t��a�:�MΜEd���,�{�?���*�i�YZZ�k�����u���76X4��|��%W�����[o�E�/O>��ttu�{���?���4ù�f���~&��47_��` �v��0(OPT�Æ�o�>���[��36�q��͍�B�8�?��?�0���)�3^#��@�͛Ӌl^V6vY}:�e�l[�e�f���*��Ps�d���r&��i�_��1,n5��HC��Q�4�d����!!�c[[�s�[�~��q���kj�D���/���{�����c4�Ф�(�x��s'��19����G	�b�6*�9�o��=���a�<��u����?ał�G��Q��s�ѐ������f��O����L�1l��F�͸>����vٹc�������7dvz\����ר��K>�G�B�!CD����v�^��u���������XR	Rc�V��m�*z��?�qŇ��X��<�фzT��é7O�	��m�)��P���
�䱟=idV�Q�Q/�����Z��M��}�ѻϴ���\N�]B�W-W��3#o����K��l���m[=��Wu˓l.�O��T���H� ����I��`��h��J�Z����D�4���nU?�^3�I�a�2��y�4�m��j�5����i���+U� ���e.h�a@H�Gd�9q���V�ݜ�R,Q�ϰ�������F����ر#Kܣ��vr(��.I,l���&_�	���ȱ7A'��8��ޖdffNv��ӝ'�[O$LDP���E�[(`��T�&Ԧ�N
p���Wըsy�cM�+G����|����Ї>${wl�'��̙3��kT�C�~��i�O�T�����s�d��k����z��e�����%ԈH![FEA3oT#��+E��+0|@�ǚ�eq7ݖ�`�:u�`�\66��۷��8�4v��Լf#�l���U�|�m���N���۽[������mn� l��cQSS�? >�����\<�v�qwYAɖC�Z�2�Ǧ�6�PC�w�kY�_2��՚'�r9�[��V��)Y�-k�ܽ�W�L`w��cY��\.��lNٜ��*��W��nj�];��!��
�Ș ���f��A6�]ط��^+��_|���ad��7���.z� �h��h/�ʔ[EC�9֤TA�yUBј�f���z�Z�/j���| !l���ٹs'C� ��8}}��F��&����g==���ɋ��X�Q�(��u��۽{��+E��C������NF�%]���y�'���C���^�,�[����r%/�Z�O��d2-�@��,^�}�?�����?�4���(���2�6-����	��D591-�z���w�U��G� �4\�`C^sÍ�u�������%~��������^��o=��fmw2x���m�/-,�[��}i$G@�.-3o�a�8o z{{� ]��Mb%쎕JJ�\"�"��d�bg�l�6��k ���uh��fϚlg�u˔� b �{8��F�5�V|�|�=����eu�	�SBTA�ꖙ����/5(��M��K6�g̞��XHz�*���0�^g�<�&5���뱣w:J����G~bjR��h�����hY�4�P��t0`*�X�X^Z��~*e5j���:�+2>>���߿��b0̬qo{A�- ��O>��fg�=C	�ǵ�^-�Ϟ��+�}Aԃ�	��J��{�����>" f��c��@U����YC���%��Y�����ַ�%i��%��:������y�z�U�4˲}ې�בpD�U�)Sc�r��qpN(�V*���:���?c���5تn��Ŧ51����/���'HX#�;veD����􅍶��\,���9i�2`�:�B>'���7��e����bk�0���'+~G� �f ���>� �s/^"�b��RO0�{4���<���q�QR��g/��Q.;�z�Lڀ=��^����[�4 c$�`�Cݭ�̴6di���a=�ְ�%��0~���0���|<kݝ�[Oo�������_z�`��ॻ5�
�T�����W�i"��Aq�Z]�X$J�iE��p���>����4,t����[���5��&��6���^��H�E�d��FX҈9A��;�6���3��Q��x�0��F,�|Au^�1��hg��;?}�a�Q�:	HBAǕ�I	�ejrF��ѹ�lz���}{�Q�Mm2�Ve�sU�����^�ׁ��
>��W|���5�f3�膉�8�^��Jy�$��t��;︋-9��x� �?���N3�y���|�m���m�߆G�[\��y����҂�)B�O��S�oW�KGw+�P�T��f�)�T�b!1���n����nV�4A��tIC䉋���aj�Zo7�Z[m���j����5Ք8%O�����g[��Ȑ��mLm|Е���$��rͭe�w*��]mTV��� ��b��D��-,����NO����Q�,+s� c�ܨ�,B���S�-`t�BbY�UH0�p�q5��~A�!� wWW���N0�uvu2T��	��!.�HH{g�YI�c}�Wx?a H�h�-C�������{CC�^t����/�Vs���D�=��ޣ?9��s���_j�1�E����>��Fd���n��ߏ����3r�u��dzvJ.����Ã���6s������>����������?���?�4�ߐh8ބwo{~~Q^z�l�&/�|Z������������x@^>u�~iR4�����g�������u�6��|�	��*r�7�FO�Q4���Z $�1S���=wA���0o�>�cs��q��V,�x0�OY>��z�+�᭛s �1�o��G)H}x=d��(�A:���0*�M�S6��a�ݩ#�J�yP���V_j[ƅ�wȕg5LzSgA;R� .s��1�7�=_w�ǫ�0����QO�p� 8��W�O����.�W��*��Y�g:�y�{ט��C4em:��Z�D]x�������4�:4�����=������-2�e:��KGx�\�ɜ>W�r�Ү�x��z��½2�@
c�뮣�����3�=�J��h���:�����j��Ǳ�:����"��a-��ߦ��3��]ݡ�ۙӣ�˖dpk�l�H ?r�y�_�#�5��=��lX�E�iR&g&�S�=�����k���u�o h�	�g:ɬ>y��I�p~T7�i�h��^^ʚf0��I�݅�~�(�?+�>L��h˨Wm�� ��vd�l������Q��ق|���'�m
�������Axmذ�ǄW_(�G����e1=^�^<�B�@�,p��ԃ�!�����6<�&<s��m)
�n�æD-�^(s�M�öyy��r�g��I�O���:��,���o�w$cd@��%ṃ���m���0=�Æ�1 �Ss[�6ٳ\�?�� <�'�=t�ۉ!̭d��Z*r�;�h�[Tp���}�i+�ݻ��gfv���ɗOH�����Ay�-�@����Q�6���I{DȡɟlKJ�z� �Af^=�EgDe�۵g?�?�{ ���s��2�Sn��mN��> +���`�ےQ���k/�L'7��ժ56�!���Iy�N����%i?}RbI��'�ʲ�}@6nآ����25��J��T����?����k�H�V�V ���7e�4�Q���Ar��	��B��+�B$/�8
 ��0�I�8�*ä�2O	d<|ozӛ�����f:��z�h�^��Rf�D؁9���@��V�6dfnV7�(ôd�Cs�bZ��s��xn��>@ǲ�추̦�n�u�6�nAyi���0��$2�P��W���@�|B����.<o�q�6o;�!2`Z�<� �iy���Ca��r��]��&��{i�	b>�J!���}�5L���65A�$���7��55��248�X;��6�z_��h������EN�>+�7�~��\�(%]�;�Cv��%����(�204�u���&�g�ѨŔ>�Q��s4� �8��A�\+��>�N(�C��FF�"%�۰�k5#��`ra}¼w5�*��
��-�|���{�4�D����%Y��Q�!ېD<%�|I��e��I��$[\���E?��+>|@�ǚ�n�
�&6��zO����+����I�� �rC��;'ы�%���	`Bn�eL
d�j�9g�<!�[��� ��52��������p�zR/��^w���h�ɼy�j��MI���<?�<�9e���a#XLE<�ƿ	�֗����K>�#+�
8+�
�5�h�c�{-P]�a�۴M_���껣�1="^�@������_�9ã��gaLDlq=�e�h��LM;^�@��Ԯ~��g�%[�aqK�(K��D�U_��u���� �d<f�T�}�(�r��E��a�᜷�y� ,���=�Q ���^�����E�٣�>*�Ϝ��}����,�4�A��1^������+�ë��Few���xݬtp��&2�;Gξ���Q��쐅��������Uc�rÅ��W�@_BN�HG�����d��������FS��P5D�[^
:�]�{�PY���:����r��>��cMC����n�u	Q �1X��FMA�D�V6dL7C.�K�)�~66Qq�w�b�|'ʶ�j^z��zd�����?�b�摡��O>�6(A��.�yF�ۄ�Q�D)PP���*����֬q��EbQz���V+,�2�j���^��@x^����~|�q�.�° �?�k�4Iu��\P��`�	����i|�R�!S:�V&+�ea!G\*�z�!o*.x�u;�]���C!��0��L��Fʼ�o��]��������4U�@���q�=�5�u�����z��>+��U�0�əI�bB��@�%r���|�vf���l������O��=������g%,h!k�:�!���F�L�&�4X���0�kBA7҄�EU���K�Pgi�4 �8�魞HDP
,�~��W|���5�$��(�{c�ݪ bRwI[
&�D��;p9��ۄ�����֧c#N�gX+�<���n��|��� ��|�Ŭ~G=l΀0�u�B�Jd.���YP�;�y�P.	��-��$�������²�/x�M��o���qYZ���6|�g�H�P5 �H~T�Â�6y�eUM��n�ۂA/� �+�(��L1�\�2�v@�4O�6���������"��p�נ��s2�D)W�v��������^��B.pc����S	ӏ|zfJ�%AC$m�(���S�zQ�%
~A���k�=N���s�@ܛ]�To�&ۆ����	��}�w�C�^dU���r���n���H�jD�pȤ��r���F6u����OkL����FZ>O��{,��%�? �`\�����`�F$��xlouMU��q���2�{iy^��9��I�hV)C[,Ȧ#?��K`AD�����t�i�&٬Tk�tZAP7E���� �V�C����5� P��3mo�.9`B�,!�b#	L�j��
9��Mk��$��<����:���)}%k�Y�lg,�W�y@�T�~zbV=�	�t!��+����S+��Iӫ��'6�3р�фQ������饋�^'74������$.<>(�a�ߵ}�z�������C��Q����'��rY9~�C�����wk�U�wh��tu��>��	���m͍^ ��$�����#R~��@$�9�φ�r��K����o�󇟣�Q��쬦�_��M+نa��-1�)� �l`�.pI$�TP�WKq�gz�ۥ��]N�,�^�	@��_f��uF�.�6�	����c!�Za#���w5���F�@ӕ��y��Z���ť�٠�I�>GjW�hj��}�� x�nG�!�H��"�XX��y�����~>��~T2m=��-������_J������qŇ��X�P�ht��*��KC/�\n��^ �T�I������M�d7x�ꉖ�C��j�F�g�H.��s���3,�4�j<��1��!�;'� d+ �[��V���?$�sFV�:�A��G��Q6����S�AH!蠔�j�4�w�K>����Y�Ruu��W��y��#���}���#��=��#���*k��^s����~�<���tD8�M�T�f	]�tB�6\�ŵ��`�
C�6z�l �v� )x���[���R���`yi^����y4�5+Ive��@�������b��z��0��.��gH����w�y��A�!�
��:�0�q�A�Ȣ'�ta��Bc����0�<Po4��m̰Z��|�3�D'��13��k�W|�k)��:xn�+y�5�y¬$�[\�Z�b��\����#1MF$���w��,[�o�s��?vF�.N�����3R.d��y�$��D�����>��c��̰-r���.,��ع���zol��J��[6@Q��w^��=��ϡ�	r�d��X2�\r�\MC�B^�%���ͼf�9MO'��F�V���}��������0��8B� ���{<�&S�m�vu󭢆H'�:(/�:*�3�d9G�	F)F'-��w��C�do�����/��x��S#类e��낡���`=�͛[�y�����@iҚ�<�aU���q,|Ɗ�@�J}�*�q~�����|�����ٵ}�!���`4F� QJ�Θ�ó���	�4�X�.]�����aF<0�H% �9S��j�Ģ�2�՟�U�z�(�]�������V�{�d�����&nK]Dq6o�*]ݝ��Ϟbi���_�2RDG=��T���ַ�Cn��ZIgT��h��5��K�O����,�g�G��B2������>��cͣQ�9��J�y�ݻ�V0�C�W�͐�������[\���,7�d2BV2 
�* 0�ᑣGe)��M����!��g�s] �
1�t�ؿ�Q�b��A�Y�z�;�)5>�?M���f�B0�Z.��+ez��.sK3�O}������o�>��?a���'C�Z.g$m��cO(����G	��؟�ѣ��G��s�����^�7\Cђ4�,�f2 r�x��`G"�'-����W�8E<@%�i�z!W���'��t���d,�5�-�{MI�9F�F/�5��xX�[����������駟���%��w>�~��~�9FRz�yxǕkֳa0�i��F��`�8zI�7�����0;�_;;���3�7��u��,4���Yo��W��xD^!����w��(��+�K�z���c�|�4���+���QCi
%Ӳ��5r�w��]~�]�?�C9t� ס�/�tO��Pj�Er�{�*{��A
Q�n�N�@�	y��o���я�B�CV��p���^\��?T�XӠ�c 	��[���@�*C�[	�h&�����ʃ>(ǎ'�ՋɤۙK~�-7˯��oɳ�������JF��dS�|�#�ǎ˗��պPn�o�	F�ǹ�X@ ^9:�m��y,����^�����u�����������l	�P�sW��A�B]4��G�`�7��w����FдE�X��C�=9wa�����C�<L��-�~�_Tb�*jL������e`[їŅ9z���?��gE]C�%�
(
���Bj(u�8�=�tMC��&U0���L� t&�Ȕ_a������յ޾}��3?*���mD����
%8����;��v���Q���*�K:ʨ�5;;O��B�mɗ����T4(|F0Z��[�8��nۜ�����:^)!����r^% z uO?av��'�z`-�I�馛Y��>�|X~�C��~H��>'gϞ�p��,7��ZA�
啛7m�L�S�&*��Q����!��?��W��?��_g��_��+?|@�ǚF5�C
���$�l��P$�7^����h�w�L�|���x�[�y@y�Q�NwЛA.��F�1�Q��ߗ���ߙc������}���,�y.�f.n�}7��
�
" �q�׫��w�Ni�J��N'B��W�E���<-[\��dQ�htbC�򣅼l�Mzxh��ղ��B^&����]"��ʳ@.����
�ǔ����qΨ��p���:���wnf��@��I��0�57G^3�gXw��k�f!~�R+��S	�>�29�Tb�� �jE^��e��C񦇼έ�`ڤ\�J0&���^��M�F�ɗ`]�!jD�at�PF�Ȉ�q({[��!�e���O,"���� t�<F�4�g��ӯ�5����0��Cl4-ܛ��d¹��_o:F�'5� J|~$H"������c/!�mo}yP���'�OY��Q~H�:;efzN6o�#���,/��5�*� ��B���|�����/ȷ��	��D*>����������)M�|f�	V Q�۷����g���, 
!����]
zq9{��,N�yݲ <_���S��3��������-s�=}���s�*1��5����4��Q�de=��GH5�6�m�,�596&��u���?:��m���Ș6Wq �3H~ �b~YN�|\A��^v�:��j(H_o�[�m�V�8w�0�K�z�;Y=r�i�	�k[�]A-��蔅�Y�o��N���u� �.��tU
9�Pȳ�dm������߬�/�=պ���py�1�}BD'nr;��i�K�|l* QF�n[V7�`���#2`��j���r�t/t�
ޔ��B?W�A����.u��ra���z��5�x�F&�D)���՛�w�Z"H��}'H��v/ n��(��ϝ����>����c�ʁ����	\$S0���C�%dzrN�}���]�7��&炁��P�988�H����M/p�\���?�4b�Z�Tk�Me�"B���W�9ܼ�(�˞���1K�@�Z�Y�fj{�C����C|�a��[���{L��կ�.�N �nIV��!����D' ؤgg�)���8+[6�JL7߶d̐��3����*b`e�T	� ���%��^8wV��M�a+X����q�dȘv5�u�G�p�.�fX� �z�������>5b(��h*�6����iv�jWC�7~�ר���=�k.�)t���z^�P�jJ��J��%�:���̚�q$�f*���� �(��$Q���Y��:�ޫT��wo� On�X��^wc�-l:�������g� �e�с.�P�P6�G'9����B:7�Z��9�a�(�=jK�IN��D��J�F�h��	p�HTpՇ��K>���p��"�2#�����g+K�j ��E��qGf���dWJ��}]�v�87Gc���G��v��H�d�\.�f�O��Ǖ>��c�����-`X`��GfeH6�1���h��|��?���M�3�����4Jb��������27;#�(7c9P�4�MX7Y�|	X��	�<��&=ƺ�+2>rNA�(��+��T�Nk�� >���)�---�-l]�Y+d~nZ7�H�ʇV�Y��rY����M�7̋m_�ˬ�ZQ��z�󞷜Vp�$iBA�9��[� ���8�jJ�:�u+X�1�Tg=r�;�e�g�n�Oۗ ��zq��R�|��v=z\�]w�E�8��Bd�х`v�z` X��%�Mc���h)���B��� ����[x_ׯ_�[7"P�T�Z���{��7�eF����G=;����A����o?�MF�z����M�:�)P*$�HBд��<�U�OU.���� KK�r�vIb;�����]bJ��^x�9�ȲGI��4�32b����W~���5�����W������U�Kg�R��٧���m;to7�)ȑV�B��zT �)+'�̵�u��jb|\��mRW�|졇xl��$K�T�F�|Eo����e]q����ղ,.�JD

���b$wU��u�գ��4�F�@���AxBkMGj�<?#�BD�ɼi�45�Ã-m�m����/��{I=u�I������xT&�'$��T�dhd���<KW$ƂY�1��֟dh�z�)��J�P���J��l"��,�������[<`;���y�)�}��} 9���Gt)��Q�0]q�,wH���������:��%���u�_/��v��;{Vv��Ő6�~%#�J�Q&�0�b5�"��`H��^q5�md{Z�BFx������/�'�5O��P�F{�*CC�d���|F��eٱm����;���#������aUc��1����H70�Q���j�ƑZ�,���^d�������k�i7t�l ��f'�т�]*V�ĉ�����������o&X �N�:ɐ9@*iw��fy�;}D������(�f���w���<����L����:IQ���Gp�Ў;�˭��9t��g%*K[<(����R��3��lF�6���1�!,�]��ݸca�N
Z]�e(����
�mD��-� ��ԄMsA���\��#���5�rhd�u!�aj�a �c	�*@���]ު��6������V��l � �W]u��>��[n!9�閜�gV10�k0 ����<��K4f>���< x�]��9J���p	h��+r��5�H�����fm7�;�SuE� �4x�ֽc>�|��kt�q��G�:;���V���D��ܫq��%9h�5Fkt.[��G>�����yV�0hy4�����y���^FN2�i#��S�fi9+�{evnZ:{���BC���2���j�]8��<��Is8���D|�8\���?�4t#ut3��=�ϟ��'H^V3ܶ��P.�ȨkF�^#  Lq���=�y����wȗ��W��KGHx�aU�<[lбxd��u�b��0jv��k��k$�A� 뜓:�D$H���"�d��Q E��[�����ʖ.�O�m��J9� 4���T ήh�0,��S5����o�z�祷����uB��Z��!x!�P>L>����w�n}���_8K���x.���+܉�1y��ë�5�����3���2���ؤ��؈�����k%e���M���=�1���>�nc~������M��\<���ʼέ��O��LMN�����s���x�M�Y���hg�?^�"�>7;e��z]/^"Y�\�$/���P�һ8/�$��)�k`y<�V6�~�NP�@�z �.��}��RC�&�TM�yW�gd����;dxx����mˤeQ��~���)D����?�q����X��� 6D��'�ƌ�Y���d��A�]�9�`�%��͸=�EA�H,,�N�����O���y�ͷȯ��W���wI��>��4�<�����hl8��0u�M�v[3�n��*K�����J�Vd[�t��
�(�p4�8%��$ �As��Q�Ԣ�=��Ky���%J�
)�	��=�Րn��8���cc�= �Q��k�;>�P5�Z.�����Ly	�@���_'t�����ko���R܇^��7 Q���I:��W��s(dڮ���Ju�2��)+ ��-�)�;�|�z�{9?#�[f���Q�&P�3�~[6��=w��q6_��P9����fe4�b:��"D�D2�vRC�#LO�\J��['o�ݲm�V���ޞ<yJ��'?)+�շ�wP�5� n�*z����x��0��H4�D���K�R���_�*�\��Yu�k�n���{;�drbZ�uͶl�ȶ�'O��tm�	9u������G�R �T��Ҭ�ү����t�i4��F�Z�c�d]�z6'O�bh���+w$�-$ �z��Y�s���|�BO'�J�8��;����;��vپ}��7c�G~�f<a�t뵚+⊎8׫ss��9R�
e!(�U�:G��y/��W0Y^����V�H!`G-8�u`�c��}���G�ǅ�]c^��p���Z�9�ߵs��O������t�����:�D������K]����+�N�� =�Hؑٙ)J�"b��ɩq2��m#4��
`�]�X�U5�r �
�H�W��5������ ���7�5�;;۽f/5�,�Q���lgu�!:Mz�8�q��;(9="4�KY��-�d��-�Hld���|V����&@ ƎH��s�ۆuM�4��ظn����M���?�jԔC3�z%t���b��#A�e����t�{��AӠ�^?��Q Vm��Ke}����� ڵg�Ԛy���O�a0-#�r�ܸ���mvhd$R�ME��\���?�4B�jM7�jQ=�T2E{U7��G	f��F'�%X��ErU"#���fB҆U�T/�4�h��˩��R�B�
B��U��[���NZaT8	���J` *�r�z�ѰD�;uСR��?����;}�W*��`^<2��I��?��8������0q<s�����i6��U�>x�흒i���A����\��5��nV7W�&u�a�[� өU��s��#��e�fF?.�^4�YP��*p<�t��Y�Ww�P�)"�qY�h<�na����|�l�
p���Q���ѰC5=���H��Ԅ	������6X��tgR-��f�(��J7��!Du������"�kK� Η�<�GF��c t1`��p��֢����RL����?��qIt��E[�-r5�QVW#�[�:�8�*ӳr��9�iF$�4R���t��C�P����pߛN��s�����t�i4��&��lU���zW�*��e��"��ըkV���b�$+%�IÓwL�<�&��պd�&Ϲ4;iJ�j&�l�=�wǭ5���%fa�&Z���ї�pP��f�f8����ˎ�W.������z���^-��.y�Ǐ�7���v�!1-/����D�0��lRwtO�����<?)[�l�TG� ��O�����}B	�,Ǫ�<�����j����Fo�i�#�n�N��W�u�ᔔ�
: o;v�ӧO3V�v������y��S�`���J�H���;w���ٴ~#K�PB�֞1yjq��r����:�x"4Eɥ�za	���,� �0k���/-/�+;��*�DX�o�Dc,�߁�W�TɾG� ���bY.���Y�V�(O0	�{]�UH��229�޻@=�?�������b6+=@���7��0)�l�w�x6ݲ@�F��t,B�LF*��|!�ƕz�ͤ�䭒�AFo��ˬ��ձ[bm!ܧ@U
~�W|���5�H�� ������ag�A0���7O0��E! t[���qB�:�ꜣ��<�*�Q��-����5�Mh��^¼�xD;��X'm�w9��G�n]ꥢ�WФ��1���M"���iCz'����S&�9���J� �K�g�g���X��Nm�~Zj��C�������6��Wox�>���Fl�¦�5�Hm ���"F6@�ꫯV��J����Ȩ���2�~�5��Kޱc�s���qZ����E󛠓��������\���# ��^;�[T��� �
!���Ȥ��wW��:#$乙c+��5  ������$P����T,�.{�\,X�����%�6՘Hv���#r�M���g/�� hC� ������O�<"cS�rn䒫�J�S��+D�cP��G�w����%�< !$&#��Y���UP��ep2b�I��6��tvwɥK#�z��{�����t�i`����GA)
����1����Y�i�U��$CA*C�5�ްYb�E*4H�T*��r�h��+����)S5�&w�r 5��p�zu������|��>�M�z�[*�td:hl��Fn w��A
�X(A[(醭��ut�����':��^+�gQ=V4�V� �\%�I��w���F����u��-Dqۻ6]�q�Z�k�
`� � Y�|�@�%��J�����MCU��s�=�p4@9x��QB�k�5���#
�(jS����F��2��<뮤+�*�x:�L{(�Zq+�cewm�[�m���=oaaY�zz�q�	y<�~|>m�z�l	 �~��ep`�t�AӖLH~eI�;f�b�ոskҋ�[����	U�g{̰�+f>�s�x���z͓�]V�Xt��«p.�lh��'����>�������ҷn���-��|���^H:�p"����Wx���+0�&A�Qb��Qjs7HV�i���6妘͛���s���C �B�S=A���`
��гf�<A�rɭq��f��#<� ���e<`=�Ԇ�p]�_��CE�2��j�l�(��^�{{��H�4�[7�Ύ=W�ٙEI�z<�F	�����D����/2"�����'Xg��Qo�ZB:������E�Y��|�-[1*��N2���a����?��"1F�oPs��
���%b���K�ZZ�9�����VkޜZ��و�a�7��z��V����[>�����_��Ӱ����aG#ʒ4��!�������/:,���;�-�Fq�<>���q�&���Q�'{h�t}@l�46.��;�Ƀϫ!�Q���r��g�۷b�P�Z�����hB�`tp�s����EYX��X�j�Me��Ek��gG::2�4���U�/[�Ǖ>��c�CA�ـ���/�F�G���Je�QsHÎY��遡|���ێ2�is���!8S�DkM7R�]�+=FD�Qz�����	�E��u7���y6FYkldLNC���T�]\�ÄI�2� �ĨS�j�PΥK�$ԡw:j���JN��G\�6��+պ���V�a���K�^��-�4���bv��5�aU\]ץ�z�f������3JxV��j[�^w�u\G���Y�LO��5� B�����G��O���WS��g8YV��Y�>~�!�^�4\ϼ�}������g)#��� �J<%�|��	>�> ���}^1B�US+��I�S�|tL.\���4=s\���3S�$�E�<���{�9
�U��r-�Ȫ��֬�`zJx0�@z���`�W\wE���H�1}fhH���5�@`T�X��J��tv����˒J��R/�ՖK�\���?�<���+XBp���P&r�|݄Y���yt,q
��   `����� �h�V�ȯ:�XG�8A/��� �p�R�*��8۔* cSooK�U��ܼ$�	ܺE6o��/?@R�$>�<tȈ���Y�~�,Qݤ�If� PO=�.C[w�%�XJ�9������J!��f���$��6�B�"��s#���	Y[0g��Y���e���OJ��@m?�nD ֶ[B� S�C�B��>s��돂�`�M���0��M�$���;^��J�ڹZ�����o��L�\�~׉�x_��繆ۇ�Q%�2��w���|{@����g)�+j'"!J�ί���_��du�hX4k�� l�����/�ᾰ"A=tk(�l蘴�s<s�^�-����D,N]x��M%��yY��!�w��۷s���)y��ef��5[�|N�DH��+����t�y4�=�:HF�F9P"i�LQ�l���¢,-�P��b֫C��P<��':o��sG��? �!?�+�B ���!�f�5�ho���*�Y��_ݽ%�^%�bڻ�S�dp�f�g�����\������zva=Ζ�����m$�ojfR�ф�u��i�y�=���Ϊ�0��I��}���BW40����]���a��''�[���58&&�x���?�
�Ü����m u�M7��j "�mɂ o��<�Մ�qX����%�����Y��bH��T[�hq=������|k�`�w\�_��<�&`^����q�u�(�C�8  |wj�]�pA����F�%�鑕|I�(��pj�u]	ئ�[�l�����v�f�H�M��y&K����yí7˥���}N&���{�<s9ٱ}��z�r��z�	��x�����y�����{5�����IN�������?����kIݠ��Ն#���G�8 ����:sV�=��.���b<�-[��3:�@X���mf���$a�E��;�����F1��)��V�����[��f0,>�S��L�f�cW2u��.�NJD7���.zWTwS����Y?�3��` ����p����z�g�^�&<z^��\���n]����;Fu��X�MC�C4� C��j�~P���37nd�^�a`~֣��Ȇ����>����a5W|ǒ��:�`�8�P	i�+o����l�%<o{����Y�Co�����o# 6��,�0��S�#�x����%6��f�eQ5�`�A�R3lw��g�=H&�2~q�M]�MS�\�l<k��-�ɺ�xl���mI�Ӡ�~����P,�e��l�ݿ_>��2��o�n���O����܌tw$�#���x��/<���ڳS��}Cy�?�Ͽ��?���/'?y�Q*�e�#��Y�����t�i���$N�!C���k�b��SA"��2l���c��?~�sR��f�.1ݐ������ o��w�'��������=��Gn~�M�я~T�yɐ�Љ�a����-/(��Ԡ���_��~���_���u��Sϱ�ȴ�9�%?���g@ъ�P�ʱ�'d����ꖗ�gX�^�~R��!*�^�z��<�>|�ൾ�W�� ��wu���#/����$S���:{�< ��L+ЊG�<� �AOT���ȁq�g���)� ߃�~��E�Fc'�r�x����,�Ö�^���Ld3�=&G^w�:�RF�*v�z}�-�cbq�n,�� W�]� ������>�@�i�Z��9�~� ���ٕ�qd�޽29�,�?��z�!2��w$J�8֜C�:�
�xf����ױ����}�g�;���9x�9�������]�?�W�J�z�1�ʗ�����dqvE.���o}���}���p̾XSx��e�Ҽ;qZ�$}�>���������\	��2��#;vl�M�6�溏^�m�NeR)��;\������l�2�(���� 7���	}��W��x:!��v������p�;��`����{v;�5�s}��!�45#���_�׾�f�� T��g��JY�($293-��{/�Ȇ�cy¿�ύ7�ք��+��j�����6*_��W���z\k�]@�=s����S'���۶�~z}�:�r��r�������42���ϛ^�\� �u�B8^����� @p��[P�� /��X�]�x*u0�,Cݖ����՜z�#陜�+E},�φ��ZY���0��"��ɴ��A�@(���,t@F˲jCRi��(�C��-x�:$m]�no��SPc45�t}]aK]7*ck�5A����/�2���|G�G��GDׅ�6mɌ\�7�q�������d߁�dyi�kybD16m�,��^:��Rsr�jP��+<|@�ǚF6;ӯtJ� T��=�j��<2rQ�h^�y����v�ǎ��������<�M�$����}C���������~�dey�� Vaݐ��&<�/h{����^�Zv�ؚ��� ��c?���2=�@��w!W��[�z3A����譣dm@�iH�B�^�@��W���xV�ׯ��	FL���;v� Α_��m	Ҷq���]h*� P�EQ�ؿ�*���5�GGFd9�c{�-%����!qD P2��Q���<�� �����c=~8?B��dg=t�c/UM��j��b_�%��l9���:��U��.5[RՊ!�<�=���A	����z�ջ�Y-�zz��+�l���a!:�v�!�Zض}�[[��D P��H	�6�UAi#:�Y	ڢ)}�|�����������w������Q��յ�:9�ʹCuW��Z���P( �����{���3�べ	�@		ԭ�J�V�:�s�]U]9�:9�����>j�O�޿�1��:a�o{�+�5�|D=�uk�Ȇ+��W^~Q6o�Lo����������I9?xQ/6,�����*���{�t�
	c:��8��НqYcll*����ֶF�%<ԡ��ښ+��;9u�,��0�?��wl��� � 8`a�T���<+�vl7�@���(��D0XGE1���)�+��XT�
Ţ�9�&��O�@��n<�ܦ����n��4�"r���u����c}��_�mjX��ߜ��sTEsY,�b�� <@�9|������e�f�v� vzb\��� ^�p�t�w�;=j(\��_�0��X7x�F#�41���V_�7�|�s��v����3���3R�5�zC�#�����X�����K�p6 �:���)�Ҩ�^�:7���^�����I��ҘA$!p(��ܵ����脇�p_ax �a�#S*W�p��<�/�a,�r�&�����;,�_��]��{��ӀPC ����~��r��)���7Q;?��_HZ׷�i���OMZ=�k�J����U��S2��ܞn�T��IZ�+XwW�RuB�Θ�� �3.k�xV@xִ�ds���WvYŰ�#�����P�s�H����D��O*Un��-07mڤ�[c�6}�g��9۝'M�M��B�<r0�8!Z�h�bJ�nz�9zt �PR3I	�&;9>.c���.�u=��D+���3�5_L�=z��u�]�?��e6=� ��ad�?0�q����O?��y��2GS�NyT ����)������֮�H(�{�V�`5CܺF�`@.��$����MӖ��Ӽ�Nf#E��m�Ҳ3����hY�e76����\*�qi)ץu�e˓f�|�e�{�����|Xa{�;�j��H�"u����?b�׈H��7��U�H��z����p�xdbZA_�s��*!�&z���s�^�n�A::�L���K�Xa>�TO>��454Ȓ�Er�]w�����]���c|zTrE��A��PX��X��	:�e���
�A���8�2Θ�� �3.k���z�5�mz�ؼ�����IY��JpdAB�{�a)�eE��ÓKdR���-���祹�U�X�F~���dth�a�t�sySӮ7B��F��T�w<C�5���R�ݻwʖW_fi�q���ej|��%���b�*>OozӁ=������ܟ�w��ߙ�g�v������}�>Q�_
���ޱ�Y7�!���A��}�*�p��jx�(��u	q���a �`�|�����G�Ҫ�Cyd�M�38�~�f��Vێ^�%f�������ڶ��2y���=rۥb2����VJ��m�-�8�|��l[�j#���{���,K� .T4��(G�b�ӓ�j�i�����yr\�` B�9b�e�u��N�A?��]�.��r�g�ZH�X����i����Y��Z�� �u�Z�B*�<���� ����ݿ_"��4(V������z����gǩS'��e��^O4w ��>@w�e�?�G�L�M�����Jfe�����F�]8�*l�ȡ#L���'Z��.XgΞ�{�����<������7��/eK�
�F�kxRؐ�� ���ߵ�9�l6-˗,�?y��2��K�ϝ��۫/�(gO����s�9iQ����M��c��G,�JQ��V��<�����l߾���/�	\ ���+�6��+V��z\ ��dԻ}&���k���*�ͤ�좆^�F��4�@_�r%{��9}V�F��񇂨U��yp|D�y���6�@E#��9���^�SS�8P�}�-/�.=��ؠn<k&��#H[�x�����X� �K��MD��p�hXS����|&��a}�X����W�pC���-��7���E6�]'>oP��I>�ཎF�l����O�;Z���I���j���I��c.v����} 7����(#%=���6Bt���?r�dΛc��s���f������h��U��챣�w�^R�P����-wg��p ��5
���r��1�K�`��B�Bp�禨����;;�
>=�a幹�ر�D7�ǧ^�z{��p��Ҩ��}�2��g�'����N�#��=�<�Ub#%i�=��d/���1x�`7C'��Y=^���tn�����9�E�2���1�PW�l���i��uk֒$0D7r�P��ȇ�'�u�-��~�sy�/P�{�{d�;;d�+d��w�k4��Z\0�E���'��/+-�2����x} ��������z'ዝ��ġ
�����9x��C@C 9a�_G�(�ŭ>�`����TX����޷����P�~ ��ʥ_�G
�x����4^7�0w���5�A6�Y���Mgj�*�6�z��uk���|��x����M\���z�<zi)dg��9ǝw�)�]{���]������ؿO�ۺ��A�^>��o��sʥSr��1��#?�!# 3�i��;䆍��pE%RA���Q��(�[y�Y4�[��頑V�<7���~�3��?�}t*%q�3fy8���W���]���O�F%iROnB7��,�l�egk{��+yٶe���G?f/�x�ɐ�h��f��y�-Ң@t��7�Lk�sϲƺ���!X�����,b����Y&&�� pS4�`|X���;�HcS������;��ϔ�216IFu1S�B����\���dSY6F�E[,|2�?,[^MƧF��{n!�
a�B�Dm��x�Mb�:�TÔz���6پg����9q��/��<
>.	��;�o�Q\9�����D��U�^ü�9�C�D.�+��i�Vfw6S�]���9|�%�b�j��-����\�������P��:��@Oy]�2��2�׋v�Xs�o�7�� ��^�!��I҈bo�J�t�ӋDm?�=�� [����e�o�M�rQ �W�(�굫e��>��G?�4K1�џ�Q�λoD���1��������hD�#~�h�=�I���THJ,쑞��j�P!��b6%����٭�y��h�c�à�>�L�s�<+o��l��6W^���ݹ��p�)5\��O�u�m�D��{���/C1�?e�_������_G?�����Z{s����Y�;�C�
3�P��/�RMΜ>/�M���fj�SS�C�8uJ^��f��Y�[)��⛂ʾ~���F��_|i3ۀ��o�Ma��z�Vn����:Z�(���5 H0=�b4`���2=:"K�6*!w[��&�wO6��6<4��[�0��_��[_��]�5=="3�	��,�/驊�u~-�M��q |8c������%�ַ�Ź�MN��Y�X���X�IZ�i�C��A��!�kEJ���m&9�PLǹ�Q�	��04��;�8�MrkV#i���r��	��.��Q��F�q����}���(���9jz�%5�J�f��"4�6Kߝ���N5��Va�_w�q�<��R�y�L(���C`�K�b J��P���V�G^Zں�����j��)�J-�p�^���ѭ�n�ͩ�Q���;��<N��?VN˩矕9�]l�z��Y����l��!	�B�o�]Ϙ,��M�]��QkLFǓ29���'@	��ߤ�r��ϩCwƬНqYC�I�M�ԫ`�k�"GƸ��J99v�a +���@��F�
�1���f���c/n�,�v풡���,؜yX������^{���Y��r�8� ��w�̙��w�1�IN��]��^}EΝ:i�=�����ٓrap@�� S�iK65��Ç���U�#G�Gй��+��ڀ�-�\ ��.�0��|�JI�OJC�I�3�~�ٚ�
���|��:|V�z�t��@X��~��)b�y�!j�A�CFQ$c��	!ax�X+��1�پ�y0�qoи��1�Z~eOku1�c�rSs��R�C��"�A�AG	!S	b����N!��=�g���	ߠ�O�]���Ք�ԁ� a�������`�OLIGW�t��U��D:��x�ص�<���.j�g�Iz����:;�$�:()K������|6cڴ�T�ei(�r�����p@�ا��d� ��$s���u�񬍎����D�hK��G����@�|��U2��/V���b�g��p ��5j5O����*LZ��E�;�^eB���+�Ƹ���d!'�S�H���������jx����zex��=��#���oYܐ��,y���?8d�Lj.n��Ĕ~��@,�\Ȳ}�ӧ�5�0(+8�����'��\(IG���c��'?�II��d�O������YE���42|������V����y��Q��\�TM_v�r�$4p���m�Q�ӗ?k���b�3G�m��]D�^z�N>����ф�6IfPB<�c]���=G�+\��+<j����YW�ϫ5��E����cP��T6Z����C�%���
�Q,�:��e0��:�ވL��\B�B�!qz&�:}h@`�_�aD^���Xy}��d&ůbE� ��ћZ;$m�g/��B�J�G����
!-�g�|��(��NA����4Xc��YJyx~kV����LS��Eio�g�\���\�������Exs�ϕx*-�3����Θ��<Tθ�ᮺ�!�m?0�pB��R�>�J����.���mP@-���z(��K�gx���Vj���6eEy�g�C�fdD���� \!�
���C�m�jHLz\tR�&g���7�BZ�S����K���N�2_���z�Jy�������"z���0�|���k�r�� ����?{��� ��P��J�f���������{�Vm@a,!�mj.z���M+S#/�28?*>�߱6��QP���AH�|���9�s�iߚ��z�~����'h�F�t����UTjYS�&k�%r�v;R��i�B�9tIC2����V��hب�r4Dp/��g�$���8Ӊ$���J$��s�xP*��J�>��у����||bFZZ3$G˺�#�J���ΆpI����m�55�������8��"44 hP����T^�ѸLM�p^���Ѩ ��A�m�R@�a&�����g��p ��5���ڞ�-P/ �d�{:�e@�0�y _�z���T���?ۊf�l/ g�4S�@5�ӼUO��y�W�\Z��-���[�����d߅7mlb8��z�J�E;�z�7�ɫ[����
y�������$����麼r��1����Y�a���eV	Y�bt�1pM�9C^ZǺ-�t��+�z/q�cX||��ҵj�3�Y�:A$��(�-�
�������wWM�x /�z�1��\�m]i��'M�R)U���I"j� ]�8����_Q��#;�����^��Co��!2��bN N"�12R���h�À��h�� ?����EA����*qK����{&{F6����Z�B?����ʾ����ǳc���Ĕ^O��-�cײ�
{x��sc^�D��#��s�Z���8��7_=��nV��Z]�(/Ԋ��8��=@w�e��ˋ�$���f#tk�a^2o6P}��<5������P��eB솽��lR=/�ϼ���@���	F���Yb�x�-�':<���o�����-<� ����W^�w��utʃ~�y�ޅ}ra`T^{�m����������W�#.+���ٙ��c�!��a�*C�0���+�j$�O|G[��^��Y��E�<�~��a+��J%��u����k���=���t}$ǎ�0�Ǭ�1r� ��� %mCÃT�[�r����q{������C� W̩�����^�~�ZA@��.���tnj��t2Ź�x�A~Q�����G���AF���H�s�(��/����? �O�����Fr۞w�Ikk;�56g�����t!����U�>��8x萬_���I�c�������*ql�����Fԥ���n�i1��B�ҽ����O�Ղ�]�P#D��g�tJ��\�7�Τ��F�I$��Q�Egf���
��#��Y�;��%&�R!��݆BȺb��Z;'�2��PU%� CO0�fHPs�;6�A�JZ��b�O/
L�h��r[���Vq\��R�`���O�00h��rE2�AV:~��O��:���yw�N�{�B$ �b)Os~�z��}�^���8�%=���,/�?#˗/�?��g$�����u���.�~�z]V�:��)�MY^}�U6��F;$�@��I&Mj� �	qv�3����������z�Q���e	X�h���3g��c�=&����}�s��ŀי�Mz��#��d�T|�8K ���ǖ�h�SP���t�,�PeCi��|�75r��1�|���� ��5:rX��A�� ۋu
�x؏�b�S8c��VԐ;�^=Z�"J3��CS���op*֮�B�9��> ͭ-�>��z�X�˻=�Hͥҵ6���HsS��� �[���=_�P��̈�lѨ%���(�w�3fy8�������"���<)6\ts����z�PR� ���s��T/�����{x���PSl@�l��G���)�d,Ƽb�����FY�`�l~�wK;�<CQ7 s n��m3���u��h8���_�~v�Q4`c����c�v�b=z�^[����^OKs�tv�K.�d�Y�/�e.6idnD�ɩq�ó�I&f�y��a���nz�<��0y�򞸌���<���C�Xc��7���Y���'��������J��ax̙;�k�χ��4�W*��VȨ�65�������?7=]�̤�d��\�qN8am=<w\_D019%?�����½�dSF����I���l���O��܂��4Z��nnl�y�L�N�-��"�T�����Iޫ�I]��ٳK�y��k����ha�L[����x+W%������yz+�z
��O����Ӹ|���d��>��N����\83$'��1��djbL�݀+��3�1��tg\�p�Vjހ��I8�W�H�¾$�asY!wxX3�=�@�O7�h�B&M	���O�я�sU�r�W^y�l߶� �Ps �{ݾ0lmv �ݤ@���l__	g� �A�aB�ؠ�z�)�) 7�t�}|�}�3���˦�Ix��\��nqy�y��P��:u���ŗ_V�4]�i|�_�x1%I���N���(��5aH>���ay[(Ŀ�Τ,���p�|��wf����j�y���[����G�w}^�F��?s��&&��7[���W^�����N�߸�s��b�2��-��� �L���V�c�؆�6"*z2�����G�;�k fCe%c�A�����TD�����ͳ�6? �!���C���z�)�a�w��>19&6\-Ξ�4pS�A�ZL���v��L�����S#���=����0�	׈u,dff��-����4��C�Ի�zd��+dٲ��s�.�pJ�VTTj�C�sƬНqY��������b���Ke��^n��희Î�ǌ�����uG�0�7����h�2���;r�7�|�<�����A��׿�Z�������X����l/^5�8������6�<�zG�Ǥ
�r0��3 ��ƙ�-U\?�ؔM>:_'H�}�����Fz�6����jJ�u�M������a���XБI����Ҩ@���f���"˗-����Ĥ]�@�5�z��eͪ��m�v�g�D�� p#��G��O�9a�Ǜ��Rqk���Xߓ�����˰)�	����KMX_�[��_�ͣ+1�W	�j�)��øh��k��V���zc8�M:)6xa��<K�P���~�S5_�[BM� Ϋ��W��R���%���}9�RQZ�%�����!)B�U�������!����QJ�b�Xa`Eh�.��
�R�\�ׅ���O<����F�n�:IL�3��=�WZ��ok�KwG'9P̧�WO>��[Q�U+���g��p ��=��ZW�o,� k֮�W��=W��E,Q��������g��_��I	�ƌ�Y B�h`�S���X�Ȇ�U��ޕ#��u��i�b�U��bsF}5<���i���?�@���" ���F��y��[.&�T�G��[2�׹/����bȭ���R�a�o!�[�ȥ$��0������祩��Q�4H����k�1��L��QH46�d`pH���]�Z�z,r��Y�!>��1@�o�.pm �h1\�����A���]	��5����Qo?�B!�u��n�ugn��7�w\�y���A��)��>?�C�4Zۚ���
v @��f�����
~��`����4���6��.[İ�a�=.��LN&H�ǔ���?�3�=$������[Z���MNN�: B<c�VN=�{;>9�{A	��#��n+�M�9��g�� �hX׼���$�p�A�M��"PO!��("����}���}���Je��>@w�e��[�-@�</^A�r�Ku����6�� "�
,k�.^Ȑ��mS��x�Q��FV�gZ����+$�����ɓW|T\cx����EӮ4�75�.0t|�n�SgN�=��fY�h����+����i�([�X.�)�X�A��;��zz����!��!{Օ��1�=����;v`:���Eϱ��p`z#� w������tx�1>��ѣ��p�T��#�n���r2 >�<6;�QXŴ�@����T� }塺��& 34@Q�A�@=p��!}����bۣ���nT���=�A��Ax��l���m�4^j�t�Lb�������o�-�S��X� �
�Hp<_��:r��A� ���c�� ����G��D�P����Ul�g����HVDy�)5����: ��&,z-A=/�	�Wt�1����-YL����C4��o~�r��!�5D��I8r�,\��u�'Ύ��%�d�|?�b.�ӯJHL��v��g�Ru ��>@w�eݜ��pDA݈� �A�6���V�Y!ﾻ���m��N��<Tض����;r �a�DX��/��6ѫı�Ի��I4$�#�^��%S��wSc �/*�u���?OC���M>�˕�V��]�V7 q:��k��F6n�J=�݈�V��׾�m@�rɆcq	��A�F8 �ӗ*F�n*�Uc��G����-�ǰ`���nv%��
�)�HF����q�hz��cE��D$\U��o�,0@0_C��a<�4�K�c7J�`< c
`
�������jx��Mc�
z�p�霑{i�l��B�$3�ƒE�h�����w�ex�i����l�5�5�7Q��4�0$v�e8Px����w�X�]��cg��a���Bc�o-�x�HU ��*�BIz���|�K�z�j��?��<��/䪫��_��_���ݗe|t����II�
��Ц��?|\�z����h�o��t�z�xY�Nٚ3f}8��� t��k�4����D "xq+W�R��j��#��N�ܪ�I�Q=#��'Ƨ��}���M���J'���qCf4���Q���¥ 'x�^��fL��
K�Իs{�?�:��+lk���w���ݗ���.C��.�o�\}��*A���	�Za����ѣǥ��C����$�.R�ή���Ъ�8�k�8B��<�bހ4ś���'��;-�t��(P��hmc�z&�p~R��!BcZ���i �!����T���sF��Ng x��&8g[.�ܹRRO������$�麝<y\�8ɰ���Ar���a  ߝ��Xߤ�a���S�%�f2��c�#�FA$d�\�_��6�~�g�
�yMN��#��,s��{܌d ׍�?"3�z�(��1�c�E�� u�tV��GY?��;���QZY"I��J�͐���E���q�,���R*�׾�5ӗ>2�m�5}��9[����7�J�V��N2�������8��������8��<@w�e���S�l&$J�\�^C�����9󥣳EQC<���,
�#C���ƍ������#^����>�Yٶm+�Λ+��x��h[��O�v�2B�G�!pa`c�j ���pCj(x|a�g�y/Y����� ���d篹j���g��FQ<���r���w�PTV�^+��P4����"�\?���1�<�q y�d�U��8F�-۶���� �� �u��yF�� =��ّ�\����z~УG�4:��\�����$������\7�K���|o:����c�� ���:�5��0��ZR�@��`�p9��B����N�Y��WW�#	B9�����>�f:��W�(�~��"8�ĭO��k�
�R�~l��Vm�K�1�I���;֮Wj���"����!��7�E��'>x��ş��Ϲ3��w���FR���j��L����|Q��w�j<554sݪE	�erb��Q���*����Y�C���j�]�V]�\���M���QC]t�ԥ��>�
�Q�
���<==��R��kЯ�5ҡ^zR�h��������뮕��?�e\����.6g��dF���M2���l:�Z%���M��w���9))p�J5	E��sK���I�"���D�U�0� �t�2i�鐪�n�S/_N��6�bq��e�V)@>/���ꥡugH�=��ib�������z�:O��\�: u�w�!
�cht��bnoP���%�w�d�].��`I����	J�S%���:o�����^(KC�`���\�Meh �cX��Wl~�;*J���'����3B�%*�!ڂyn��WB�|��=z��/W�:k��P�C�����W�:z��]�
�^�\�ϥ�Qq�%�����
�>��$�k�&zm>o��P�I%f�U��$�t��5�Y#7��J�Z��t=������|�������� 2`�]�&dIo�L���gd:]��3%��-����	�����4�\O�{��>�wP7t�.g�uƬ�r�e����&]45��8
KҮ)2��Pegws�h�q��9�3��0K�ʬ����?/7�t����.ϰgË7*byؼa,����O���Nom
J������x�T{뭷$����+����GY'�����E��w�/-�m2>5�s�0���><�	ݘ��n�	��JE�j��˟�#�O˻���t��ԩ��ͦ�l�Y`H7�^sE�y�@�lw���� �I����
G���(�F9T�`���`�S��{��:P�C(dE��ff:������X����� ��$�)2��9��]'��C�(�7o3�a�� �z�р�Ü���#�.��5���*����(��e�2��d��ˆ��T��*#�z�{<�<:�s{~�$�Jyv�Ct����@%QB}:� ���'������[}a�D>�	Eb�[���ko�"}KW�ј�u����ys��!ʒE��&Ϟ��[������+��3�1��tg\��U��]C^����X�d1�~e.��{ɒ������1��7�i¶��� Ȫg<|qP����ˇ>�a�����{�Uo�,�����i��Ƹ䭾�v��T����  ���ǎq�G�Њջ�[Ǐ�Q����ѻ#�d믾J:�c���%�<�$�b��4Q���$��ꁖ*e��3w�;~����/X���\�rH�f��`��
���p,h��E����c� F��N��2r�YS	��EA�EI�F�Tҧ^�b���4�IΤI"��� ��� �5�~`�27� Xd����]���װ���.mv��Я�|,��4�m��
Yۚ�l��M�)W�/~����kl���ԥW�0�ۊd�g�M_s�9�s����;R��"~L;W��-�y#����a����0�mT�00ix�QB���:z}g�Lʊ����&5���[7�ƍW�!�2��ӢF]Z���{���Q����1��tg\����%��P�#?	� Z��5�Pr����N>zw�>����O�{�~��������ٴy���{�����m!�%\�3Gn����h��kW���3�:���/������-}�����d����<���{�r#O�\)We��

��M�����#�׮��n�M�~�m�5� �X�A��V�����>���K%�]�v�"���[dx�";o�����	��3���2?�%��5�����<]��?Dxة.�c�d�ɩ��* �	 ~��En�r8��X'�z���܆z�^��U+�����'k\�(���H2x�L �:�B�`��!���Σ^��ظ	��B��j�?�!���f!��j�j1���v��j���k0�pm���w;�O��%�m8��.I����ހ}n�k�����i�n�+r��7��U���O�a�G���i���5���[280.�-���2w�G���>@w�e��[��C�Uÿ�|QF�'�#I�3M(�T` �p��Q���b�A7K°9�ܹ����0�`����V X�7T�%�fL	�D�!O<�HF>�xIo@=s�S���g�����!Vȳ��f)i��l�P'S�06�������3�.��}˂�>�8�>���6�w�X��㨿���wv(0o ���F��z�'^(f��s�.+̍kR��9O��_�����8�U7�1�$�)m�d�2�1r�,زek�)�DbjX-�Aq��'�i��6b48~l#4 P�=X?��Y�N1W	#z�b�r�dHd�M[Ey�HoV#�_���g�F�ǘ��1aT��7��F��Vo�4Tnk��J5��m�� <�[����o{ܶ�o�6"D�\�r�M��U����zw;t	��������V�����_�������TcpP�zk�^_B&Ʋz�sd���F�O���S'�:O�8��<@w�e�j��Η�UR��6Y�/�"�1�3��t�p�_xu N��St�B�0X�]m��Wc��K뱃l1Z��� j4q�����p�q ������ϙ���e5��1&���a��m�t��e�8�	���~���6[��0J(b��B���ak�毠����O<�24�@<f)��x$Jp�d����:v��jh���e�>�}��-v5�b���d>�w�^��� ׎c@�^;�dP���B�_��Zy\������cتr8�i��#��{+
��;�]��ikm�@"h܂h�k֒<�셳�p�f�ղg�Nٰa�t�wpN~5�@8�:@�@PY�Oۺϕ�a��!�Ӹ���k�@��+60��z�� �F[]<�U�N����#'�q`��M��}N�E����^Lȡ�G-�9�tu.�p�QΫѵf�:)�^ĳ�
G����Y�C���	ּo���7�j�k�`���t��;��

¨͞�������6@l��4��2�ө�E��ՠ������qk�ѲQ�����E�BH�D;��3��y���y(��@�.�E��	�Z�(�e �B��p8HOӉ��/��.�{�"�����W���9'T[�҉#�:��������5֟�����%#$�ɦ9�ֆ�L��%VŴ�9�.4QN���ĲjU]UI��;��0b*=�R�e`h��Ćf2��^���0Akk��m���y��M{\v��q~z�(��䡇����I!����Foz5rzΓt��<4�+ղ�}��������Ǐ=J��m0�Xyz���w�2��C>��!�C��n����˙α������������A�J�Ҵv(^�����/�� +Z{��F�F��IiR㳩є�-�c���,i��|<.�W"����Ę��:cև�P9㲆��/z��*9Z�b}3�=%�xF�eF�D�L����f�s4"��R"�VY?���wv�R�D������ɏ�7��[���4�]l���/�H���&��(�I�G=|ݵpdH)F�V�Ur��sVϮV%���H��r��iy���h��C��QS������!�d:#7�|�D�����>*{v�2�`:%!5�ȵj~���<�q�_�1K�9������ԣ���1z�K�>F���PBC=:��m�\ ˶����i��7�e�M����H�K���T������#����6�-��wv�!Y�l�s�eR�3w�,[�B~�O�C`�\�"D��!��N��y�5�kG���-/�K�#���0�M��C�&Oo���/@���]�Z��c��ư�8�M3��������Ź��VYлPj^��5S��\���ɡ;cև�θ�Q�T+�`��e��e�6]T�{H,]���5z�~��jV��*�i��E��<�e�,zl�d��o����#��&�����>Bڨ�P!�ja�y�{�lo	�	cr��B)�fL����B��wn���un!�W��m��{�;�3�ʙS�����r��Aӵ�S��s:���S�+ɲ=x�W]�^N?Be8�E/�ڙ7��
������Rބ��U���M{Q�qW�*�r��>��an�C��DbF�� �� ՠ�	���V��s��JpwAaMLA��~�'�K��wY�A�������s��R)�0T�a��9�cr\߃����w�p��^��O�'s���<!sj7�{0 U��`��g"Fji��b��b��mF>�cs�����s���G�1N�8I��ھ�-9]�I��ʢ��e�6�
Uz�e�4>jz���7�LHCK��kB� N#
Fk tX�Θ�� �3.k�Þ�z�U4a���0��Xfki��52���Xm(���P.=3��X,W)���5�GGFXN�M�56nl�)�[��޴B�x�l{m�mϚ6��i��u0�&�}M�Y��z��}=�qr*!}����>)�<��__�=_�5�jL��2tq@̟�y��W^u�T�>��5�����r�y�ͭ�iW,o��j�3���0�67ĥ%e�8��C��R���5M�$�z�h �F-ȹ���Y�F����y��/���L�\'`�#�B"�r�6������έnh����+$�k����X4,������{4G�y�o~�_���}�Ш ^q�����@�z�86�WK�:���(=�߶��c�+�|�[� ��,#�J!�M��K�l�����鹙*����Ƅ�0�c� �Wb��>gtv<l�Jp�$������?��_��5��LG��`JB��Y�;㲆n��b)_�����eX~Wp��������p��7c���%�+>��O�}�c�°��V�y��ʮ];M����k�GM^=�Z~V�)����;c}  O���O
�T��K���d\���{�֌��z�P�V��(��6m�$ǎ���(>�A8����t�����E� �h��|���1G��m��>*�ny]V�\.�����[��6F
��*�6z�{Exa_[����Sr��YY�j���_���ܱ]^z�%���e��>��߽{���_�9Y�[��̒�/~�"x�<p��q�m�ax=��Gu�?#��.�/}�o����?�������&�Biki%B�'�MS���>�!�3<������Oפ!����0�>$�x��F�t��Y1i)��q;��W��.�iG77<x �����{"2R���9�>���}�����r�R�ÇL.�(ĳSRC4�b1�צϻ�"-m~�W�)�̵LO�HM={�'@�hmm��3�1��tg\�Ѝ����k�LIR��|.���y"��W���wx\%��%B��x�O���{eמ}d��ܸq���_A��{F~��sRIE�4y�p�['j������m�������x=~�˖��0$��nɌ�Λ���o�믿Nֺݛ�z0����~*3��`w�v���rZ�/�e����b�\��!���p��iiX�TV)��)@���wG���jS�c=:�4˧>�)Y��m���򋛙{�xݵ
��Ɂ��exlTV�XF��/�KXo����P2���<p���|�Jg,\��=�m���z�0�Э����Z�[��j������ � w��9xh��]}���j��0�^<�v::ۨ>7�w���G%A(������zo�jƸ��6H{�G����3U�3iЊ~`\Z�v���燞�Ǌ�gHA���M�{����̥�
�3�Ȼ��䆛6Ȝ�m�S����d߾29�������.*�TN����;㲆n���n�C�<���|�ᐴ�w�KC.`��Kl���a}3��[�IO��(,�ƿ|��<<����o��%�����_�Zrټ���YU 24�AL�����Gk&��2�U ,� ěP��n9��X��" rl���sH���I�,Q_��������^xAF�%����1��̨/(���ˆ�{<�2��=��_ɉS��z�U�~/�N*~2!�Bt�C�B�v�.)J� �?~�19r𐴨{���~*o��]���,[�\�y�Yٳ�]���
�y��4eh�����~�3�(+����}^��47�����S`Nw��u�+����nr֍$�<r��o+��5��aL��_yg2)��ڍ���?�w����{���M�|�R�Qo�o�4رіz��H��/=�v4;�D��Sϓ���1���d8��n�j�����<��J����/B�_�z�H} ���y�5�Γ�߲Q"!F*�Z��OP��W�����d�oȡç�]S��T��i����;�F*Uf���y��x�sϽw @.�$/��ի)^�<���
<��c�Y��ںuW�=���\�Z�����KOwER*d5� �1��H�^� x��������O����3)c��Ӎ%f��F�yao���d*9i��f)��)��������:Ϥ\8wJ���v6��X�� ������L���G��Em�{�
�\&C� ��fG�!�W�K�у�u�#F�U�����9TCc��oIT����E��*��k���a����Y5�^���x�0�ʛ� ^=�~C��h��O ���lJ㬼3�$�M�z�Ly�p����u�"�䔰�y�ݻ��^ܷP��d��^r�,�3�ِ��k�;�>M �q]�sf{����V�n�cwC���y��Y����-�������,t.Q�����Ck?��Q��K$�u�WȠ�e�\A���F�/}4�pKE�Ʌ�;o�{5"S1
���I�9��4@w�e�_�z@�&	�խ��*7�t#7`�����G�SU���/�;'O������}���y�����W%o�7�|S��:-��q��K�7<-���"��V�f����e{f��H
{a�f*��n�d��1,
F}(@�w_�b(��,�Պ��aX����/?��Od��iY0�KƖ,���]�l�P�D*+C�3����r��=�Ikx��-P+s�q��9��@�V�v���C^W/���^�[_G'�� �p�@��G�4��w�gr�h�S��'L8��B^�PG�oQ
 �K
F/�7;��ܱ�TxSo�̀ȿ�;˜6^�Q1��=�@<��W�{n�����@���[�&]���k,-u;��zצD��{��6��w�(h�a\��\��`M���X�xS��.\�F�J��}{��=`Ń>C�<2_���5��'+֮�e�7�=�Kjʆ�	4��@"�Fٰ~�<��k�͋K���Y�;㲆_w�x,��ʮ����޻��ȑ��S��\������&����n�W_�b��k���#k��@�ح
s�tˁ�����������v6�v��&���D����ٟ�M7�O~��'B�_��$� ����QA���}������BA��Rc9�|�V����v�����r��~��4 GELj!�`��$s%5z����HC� ��Ks<F �)xN+�������m�s\Kj��k�$@��U�`A�e^�L��k�Yy=V;�
��C$b� p�{��I��ŏ<��g�QCo�U�Y�gSs�t(�
"죞ҹ!��Ⱦ/87�-0n�f��0�(w��M�2x���������{�T�!�����O�(��.{��*T��\��۞4�v�C��Z�ҹ�zVc�,B���V�U��@�#	�J���,���'eѢ^9y�ϵ�ͭr�m���7_����'�Ҹ�6�$W��Z�~�$�)��C�����>��"��� �m�H�Rg8c���θ���֯Y��xV::��ƛ6�&�I21-�(�.���m�0���.6 9w�<ʯeيE�}Db���P�mX�<1:y}�_�%�>���<�Fy��ڼ��u��b���,�\.�� �|�f2���V�x#���Ш"W�Y!?��I�cA����s�9�f�Ź��Fjڹ9��._�ܘ���gN��b�h��Q�n�O>�aI�����o%��P궢��w�N����s�S��������ab�C� ��ym�� ���I��xh�y����Ĩ��J�b�+�,Uc!F �p�<P��ܠV�~�b"�(+0����9o|�����y?��!�{��A�<zo=�ˤ�����X�r�dR3�7�#�2��h��׀05����u�a@��aɦ����ȧ��0Mc"�Ͱd�
����#�߇dp�T0޲����f�����4���6��q#��<�^������R�{�h����$���l$s�ܠ����ge��9�W��|�e�+/�H�H����I|�ؖϱnjj��Ũ���(�z�b�2~�=��&�?��8��=@w�e�����������^��t��IbfJ�ᘑ����	o�Q�e$��4O��"�0�W���/Js{��\�Z��>2��ы\AmA�؆�v�Bĳ����t��m2��@��C��)�R
�n�[E�,o�<5�Q��l�a xtn ǡ�L&W � 4���ʊU�e�w��[��'�T�K1�����>�~�[��L�wv�Թ������N�W�k�N�X�z&\��W�k5!g��b�z� �a� �⑃l�&(+�W���&�����#۷�u�֑�p��Q�����`H)���5V ص��9�������g� �g���O��C��Ģq�������A�� Z�*#�p׽d:&ށ�ё�_��g�����7��*Sj��TC	�����=PC'�1�����G)m��g�R���q�`�Xf���:�1�a��1\ ,T)������ b�[ ���8.����u������oB�B�X2�%�`�/o
����[n��'ϐG�l��L�X�sjX�K�W��)<g8c�������=on�Mw:��cS�T��4��xز�v[Kx����
fy���%�V��w�-�ջ<z���w�_9w���d��FF�5�v�n�Pݵ:� ������3Tߨ�����u%��0y۠����@�`s����ǈ�$SP�cI�#�<"��1Y0�[���Z���eNW+��ăz=SE</7^'7^�����k�ʲ�YK��ȡ=�$=5� �gLo�*�	�lR)2�M��Z=dl���M�H�g�x� ����X}ק���C��6�e�t������ �-�]�X�f�c����Ő<���\��{��["�����)������	�s�.9p@�ٹ��AG�'�C�<��I�5�XN�05���{�C��T����ǚ�؀PPY�n�/@�D �eS���#��#��J⭺� ��Q.,�|��Ft5�RΔ�!o_(����C34�����}�3ʴ�ٿo����ԼR*�dF�Ά������=�T� ���i��|�@����Θ�� �3.k�s96[l�`\C�-GM�*7��d޼yl��:�r�"n���t�iǈ�l|���7�%����K���?�q)��֛o�K�~+i�[2�5j^h�R���y����Q�<22"�#��9���s�yZv����Jz�K���5�0��G�"%���4<����*�4��d��H�gY�C��OJ�+���ѧ3yʯ��;���+8�ڿ�e��259�P9J�pL�����Any���o~��R1��($��a����R��F�M\����=���1D<�%g��y���kX������Yϸ����C}�!qpVyױ'�n����\-#��U*�t�����Ŵ���w��E�L3}��w��_H�ټ�L- ��^��JI$g��N��`H�iF:������`7���n����G �_Z����^���^S(��x�} �ُ'�\��}D�wӍ�r�
�eSlV362D=����=������z���ǖ7���i�W_-mme\���^��{�� U�kf&g8c�������n������|��J~࢜:}L:$��t����L� �ʎ���[���?s�]� �N�>-�?���ww1	ŭp�4� �&;\�!�����
�+�R��!^�O|��-o��ߒH0 s��]ާ�)O�+s�/�����h���0�}�����!�\�|�3˖�7IWO7��Ȑf0�$���̤�6=�������;��Y�&�(po yW�5/ds�˟�B��ͼ6���m�~�ht���p��{ǎ�A����W��3N��11>���s���w�
+�v�U=�Tvܰ��������>����dǎw� {��)������Y�=,{��}�XQ���%�^9T ��e�P�;:i���1�l�Z�Y���g��|��7�{X�4i��&�`������/�� SO����j_�H�V�$�h��4���|xI� ��n��&��׿��6 �|	Z�Ui�k:���8y\�u�X��`�A<'�׃�Ap	p߻�:؏Ǉ�_ϜN�����Q��y=��d��ݲg�.rR��+5�v�֜1��tg\�ЍХ��ʠ��n�F��O�_���Uoo5�2 �0:�)h@�t`p��Ml�� q	�P �����Y�U��)z���2Z�rSL�p$fB�"�%��u��w�QcC�p�45Fd��U�J���6���X=�B�K/����!�b��m����n�������
����%u>)�T 1^)�;������o2��S��"aK���w�)�c+��{۶m��c�T��z&�� p��=�JXq- nD$�<�6miޏ��կ��8G� ��K���в[��0��x�<�-��50
 �E_t|���ԎG���`��ut\{��g���S�6��u��7�,+W.gy�w�&/��U��|��E�ʡ�G(:d7T�yC��������%�M�s��l"�y�:w�������ܸ��D����Jkg���_��\�f��ՠ7��#8L��y��F��ׯ�F���8� i`Sx��dD�A̵�o��9{Zn��6����YP�U����Z��g���F���d�����g��p ���M޳�k��yA�9���%}��X-5��g���lS���	z����k�0�O|�S�G.udl�x�
�k��G�������R�W��J�!*T#�{���!�=��S��sϨ�:.{׫�TU�uX���;�9oeۙS'�?�����.�7J���<�� L������Бc
,
~!�	�Jd�����H��Eɪg_ �/ ���R��eٚu��k[���%ndsA^����уE�n���@�OܖsE����ҧv����Z�Z�ה�.}(�G��l5�
>0����G��� .v��Č��'>)���y��W�駟2�
p�hL:;�����$�L$/�u�]�HK�0qm��VAGwk�C��lg�mOQmp��QiWP}��-FI�X�����=8���̛�D�+��f���+�9�
L*�S ���q9!W��F��5B
��z�\�B�B�`���T�X�*�"P�tRc�!q"܎��M��ٯVae�jAr���R��c����C|�Ϟ?����T�Xɻ�����:cև�P9�2�Dx��wn�ݏ�#<�b�B��g�k]�t��u�]r��A�;q�@����=s�'t ����`�o��d��(������)����R���8'<�r�L�yaS�l��(�
U�̋��zޭ-MrH����=(��88u��^D��,�h��� ���!�� �J�۠_�=CO�����D�j���Y5��iw�\
輽}'��J�4�)"iK��{�[n����O�d��>�;���p(���k�;�Z!m��h5�l�u�v��Y����(�\�]	�0(�b.��H�5����:�5�'z��P��_�<��+���&��IvE�cG��7���/�~�̙3��3�ú��\,��� �x��u��m-2��[����q�d�5���|��߰�J!'F�h,�,.��2���޹�c�����/�� ���O�q�~�����rT,mF� ���&I����ѮUǽƺ�9���_�����F<Ͽ�I�ီ�\2���:�F"�gq_�듸^���&&��g��p ��>9�������W 
�t�Z!uy��y��7į�,<�Qݼ1���/���瘫���kY.�M|NOK��~k�{�1l 8����b���u��r�i �z����=��fHb�� W�X7��~���կ���՛��6ƃ��� :��D�!&]��r�1��Qҩ ����/��sd��j���@y����/��oB�`����?�R3���=�̽��P/� (D D��6���-a�;u�aDẰN��Gc�iDJp,|��ۃ� O�̔ J��\g��5�&C���G�S�%�$z�.�/�Kj�m��������:��PB�uY�;_�X�JΝ>Ŋ�^������3
.EB����d��"���q�s0���u���޾^����$��[m��]5I}�y��	�:��'��M͊���+�TϫTK�w�z�(�@*���ıc\+�� �	^$��{b�iv��5�:��OI�ܪ��>��\��7*�p�,Н��D�����"F��jaZ���gw��t����5`�zM	6���O�k
B~��r��w���0ˆFG��ȡCd�{����v��U$LX���7CѮ��'vKA7gl�02�/곛c��,_>� �2%�zy�lδNU�Ĭ�xc�='��b�������Zs����?v���ٽ[bQ�e��}�A��'>I��_<��Və)����g˥�a��P`�����na6���g�l��;<o���>�W̍����q+ꁿ�/Z�"k׮eH �(
r�۷o����T�E�+ZZ�EFp�s��rM�F`������Rմ#u���񐆩+���<>�u���+�-��O�8�m��-:�$�l~����>b�)��2��=��IY?;2ԯ���czF�&�$�7�sE�{.��j�r�暫��ֲ_�_�L�p$���b����L����µ㳈�@����5�$�������[��lI�nD��eB���#a�֕��8��<@w�<���m������ۅ>�U�k\�y?EI\�n�eZ�����L�8�U@`B��������{��uUYûr��I�n�eɒe�9`l���`Hü�`0����<�,g[�eY��d+�V�s������k�{K�������u��#��ֽ��{}�k�}�]w�S��k�Z�'g�yw?��%y=�@4�O���ܠE
�2Ӝ%R��n�Q�c�A�L��2:�G}T�%�޷�>�f5���B�.�gf��'���6�0�m'����eL�THI��$�}ۖM�{(4��{�	z)	��n"a��i��o�s��S����2j1�0��Q�x�~�/�6���ODJ��tʮ�;�ְ;XǴ6љ$�!ώdv�T\ V��O|���~B����S�`v�g�2E�<ET
А�/�,��<�><���Voˠ{_!�nvM���y=$��Q���pe����*"5z?�O����^3������ �JU�-nOI�[t��!���T���ԲP�t���Z��-"&� b��ky��GG�u^+�(�gKL�p�����싞/@� �vY�'p�-��8���Eb��5�z��*��]�f6HT�-F�����	�,-�j�����L(6Px�Ua􉞐'{\�l��R�t2��l°����𧪛�l5R����+�"֯�X��je�QO=GO3�HK":������N���Rp�#ǎ����us���)��l�Z�b���q�Lim�l)�S�D�eQ����"A��@�Թ�i�Ȝ!-䬲1c� x� ux�X�@�S��k7uA�>|�A^;��o#_�� �Q�kȚ�a�>r� ~<x�o���epȧ�K�1 �R)�ﰥ�^����w0
�`���O�]М�r�r�n��=�K�`E"a�	sC�F��D'���G��V>�I�	�Ct�+�L{�ۅ�.ϙnm�DG�$�>����j����+7nA:%���ͤ(	�7�ms�p����~p̐��ŏbC�LaP�AZT���˦i�D"!�l�ю�~L6�~�BB(�#�:��8��q.#?{�̑l>�VhpB���1�R�d$>tcv�鈅�ᙣ3��� 
�7���kEh=�`�P���t�6.ʋ��B��i���/\OX,X��0��Eo�+��� ���	|�Rѡ�T����G]���Oʴ�3��e���M����9��T�z�%݌�0B�{ۤ�]�vI���g����m��+�G�c��n�')F�Mp@�޳]���Z��m�����$��8 z�`��| $�y>�n$����  H�O?�s �p ��t�ʕ+	�&�>*_��ef=�}e�+�O��a� R��C"#״Y�XS����F�����M� ������>0���%S��H�9V��'��������KVn��J�٫��(�D|��p�`�$&s�;�F��髧k�LC�(��z���Ri��~�����4�����I[��cj���>A����\އ�A�������>}�NJ��|H?��Wy�Ϭ��$�qA��d�.���8ϣ�q.�s�T�4����b=N��8�%�#��^ج��+7�B� A�V��}�$|� C��"l����[ ���xM�9��_�e]��ZV��[�!����������������Y+�p|k�T�G�)�R/�k�e(�s���Co����M�T(tB���eos����|�?'t���K��T��;�BUR�^֥Zω\=��Cx��=����+���f���g��rH�34T���n�aD@�w��۷G�,Y��8tŃk���rm�-����&�_K�"r�0 X�U(�ۑ�����ҙ��&��!R��b�Zu�`�O&R������i��9*sg_ǢDx��kU�w�p�,]vǞ3ݒ�Ee|dX6oݬ���/�Y�UX��c�>��9Sϳy�f�2:���0fUT ���w}7��[[��3�c�]���WK!����TC�|�Bd�E5*Bj���h�@�ʨ��<*�^oLNV�ٷo�n�N[V�X9����cμdm��h9��(�ۆ���p�d&k�OvEcW0s<�|�E6��4y���EP�3?Fƴ*����AX��XW�^?��m�ن��ͯI:>���
Ѣ)��_M��Bո7 ��v��4�H��P��4�g����'���́�9�7�c]rΡ��Ǥ��2��������k�����&�d��L�P0�Q1��ZBM�^��'Ήc�����ڭMqN�<�9s���0�m�}46�C����%��}�&9t��x������5�MY�;�і)����:TE̚���
�Q�&������-�W|�薭�@԰:��ͦ'h'��N[��r��1MV�]�p��Y�إ���7�@둅��)��V�G<z?�̤��g��iҫy���ǧ�^8�Fޤd�x���XF��^ ����yM��Ӵ��zC <�G�_�X]�9��e���<�d����#r��Iٽ��?tR��\L�8K��TFe��Q��x�c,����j�EmYV��OV9��)�m��DdJK+7�޾n�z�)��F=0ژf���K��<���w��V��@BH�f��dZ�z� C�6�\;dlx�z�5��r��tv�SZ�*(��!�x��1w����ߣk*���,MO��}~xm>�ݩ̐�.�`�$���2ۮ���ק9���wC
�bz{��_������Ќ-Z������ �gI\�<�{~��Zr\è�9�}#���� ���cMlз�v���D	���/�'�=�r���r�r��y׹@�ǫ�E��K/�,�^����~�i5z|�r_r|FDI���	��b�ye\$@����7z�j@��,��%6l�������&�^zY���=uj���\+�r�h�[� ����Koo7ea���
5�� �(�+��@������6<}����ݱfx >Q�xg�e����ZJ�!�5m�lX��鎞<��_-E�G\���^}5�7>��lڲ]<N5r}lؒ�ʨ��<*�^o{D�1.��!q��z.N�{����3d�zY+W����f��R���y`������9(�9��둯���r�k宻�%q��)�ҥK���Y��N9������
y��<������Y@�������$S�?� ^/�p���!	��exBdނ��)G$�DH�Z�EӼ�@�s�e̾���u�8+�-g�6wDМ��(A!Z��%�\¶��z��`�d��;Ը�+��!٢�P@�&�l�����e�Vss���d˒�y������Kz��j,?k�*K�.'@!l�Ndl�r�0�m��a<~�fwo��3�����vz�0 �����lY��a�(�/�(?��${5���U���y@=pT,�C�z�
jN��gr� �@��OA-��ۡk�:��!�U���ɓ���{�G�����z#�F>�C��葃l����)M��;Ŝtu��k[_�|�jȅX��~�E�J1[����@�yu��S�Q�t�!3�,d
c<:�B���4�P�Mǥ��$�f���C���������ך��t�y	���뮕��ny��	��Y���+㼏
�W��!�3�s�����5�6ˌ�3�+��5k�ғnh�/�q�_�N�_DM�|а��\��V�^#+� �;���r�W˲e������Ш���)�;!�
�u¶�i���^k �If%py�����oH=�t�"zsc�e��d`pD[ڍ 
��|^����7��(?���Pl�ʥ�݂5~�U�
 �`�������F�^��[n��\�zТ��2¸ �S��#�����Az�N���6Y�F���&���������p<��烬*�u� $ԝ777Rm�����Ϟ=[�=N@O*ȡ*���,O�s��R��z��g����`U���"�덜�~�н��i�]^�}$DR܎ �Dqzz���-������ȡ7c��3����(�<��AĀ*�j��hH��� ��<I�q?4|L��O�aw�����M�9�f�@�U-5u�j��r������d��޳K��	�;q��(�����g�c����6O�E/Y-�f/U��/u�Z5`��N䤘���X�x����{�!�Ta�W�y@���=���D��X�98�7K���
�  &�(�NƢR_�hHm�ID�g޳g�;v�ʩ��ҳ��G>"۶�&7�t�z�U��|�]6�d=0B�۽¡�eJ���w���j�p�ۧ���M;_��c[���ӹ��V���H�0%U��� cB�t\�پ�52�� ��� ���V����e����u���@G8J�z<�tfy�8-T������{��ʤ4�X�"(G�V�h7�6�VY�������P�MT�g=o۶M�C-�� �Rt�21�EGS�s�x�a2���6��#V��<��R�ϴ�t�D����g �@Dbp0�G���ř� "��F%d�c�!0��5�����*9u��p��n����{#��Dȝ'O��x>��ϧ��1�L���X�`M`0���6��	�R��=q�ǃ0��Cn�ʗ���M:H��)Su{YV�w#���;R'=]Q�U��¥%������֭a�{Z���6i�eK���W)�OH*�(�U�y@��s��%��v>���|6������f���n���V`�p�2I�����?r����L�a��
��ؐ�����!�@յ5$��졳�ʪ{vXyxlش!�2:<"����#�����@��3�Ĥ��C�(��2���r���O�[�[���<��3��y�ׅ������hH�s������f�&@���R ���nK��aI�@��~��d�*��sV�T����t�];��~�����,��	�ܵwL�� 0�ڤ80�O(h�Ο˰=���t��!7[��a����Dk��|��s�N��j8%3,|��!���BT���IN�:y�R^�r z~_�G�Nf�(硐M��
���b��ã���X�h;�̙�Ƞ�O��C�+"aj�]��A4"��ү���T�RF�FA���)�rJ�2��xX�+.�L���\�/�G��AP�(Uᠩ��Bς����	�#�����{<��ǔ�-�ؤ��9�C$�H��FE.���O���>*�^�2���d@��a���2U7g���m�S(\��(C�K��<[Xb�̦?(C���M/"/�O�R�8Aю4������;���qXlx�\w�x�hՊ�(�>�Nm��i���T� |YEک����+ܻ�b����}��Kk�}J��m���������a��<��5��<٩�i�����!�����2/��!\*�ɘ8��15b��5�L.����`B�T"��y��l��F�լ@��a&��Q��!�����îvmSejk3�$�3�j���YMm��G���8�RQ���3Ϙ��
lj5)6�z�`1/��(����1]�<zm��� -m�h���L���Ei ؚ�o��ed�d�.��ƶ�,�����޻h,f��腡�� ��hi����t��?3c>@$E��֭[Ձ��Kj�@`�}�\����5F�j$�5���L��~o�:M"��w�A�\�Q�E��z|FƆiP:Q�Q�q�G奪��=�ɑ�����@7J�1kJΰiN$RM��ߡ�6k���A�2��(��x�]� ϊ��8��R]f;O�dP��(����H���
��d &�����d�9>�;=��N��{���ﯪ�
���ή��K&�!��ss���jڇ�ۏ�;�t�z��<g+�!�˲:�&�Ȁ�!KLz��E���/}�K1��  �!IDAT���׿&0�h�2��a�za`��~��,h��R:����z��"���� �O?��\�a=�� ن�&�{jp�Pps�M����qY�j��}睲q�S�[�Dv:�t�~`G11Q��?X����w��l<7�tSvXt�h��#5��kT�[#F㤲�E��!��󗉋8��%"B�`-}0@�$�"ԙ��N��a�5��lP�Y�x	�h���_���6��ܒv˖M����Y�uu��������sF�/�@H�&	E���'��H>C��W�xtlH%����o�o*�2�� ze��1��Su��������acSD������,<����I0`�b2\��3��pVt�E���������R[WCO�NV]x�\}��r�]wJ_o��¥T΍�r2摗��;�ƹ��Ep ��L�"������K�&��.Zg��I���^��R��fP�s�I.��D	}a������m`��=��rި��@H�Bt�VI�PM(��,h&�#��01R���@$@#�����Ѝ(J� o{��a��k�Ex��`)�D��9|��_0O��yG�5@����F_��������֖&�!q0Αc�5c�-M͍��C����kd���V���u�~
�45�赂4���oji�0����9Ͱ�X녇��-����ݱ��X[��i��ǀ�?�q�:��=t|�0��#1�}����ܧ�ᕗ�R�� �'��qih�ȩ�#�6s����^5����
iiE}���d|Xv��.yɨ���W�����ʨ��4*�^o{L��N��\i�IN��{y����>MF�GY�@���ӭoh����G}��9f��A��Ƿb�r���?)?��e���r����� ����!a��cz��?vX
q�����u�־	0G��۾������~��5���VS�	0�%� ���r7���&�KMD=�(����aF'`$`�_9�à����(A �{}C�����܇n^_��Wy}��'i�wۍB ^6�ap[5�s��n���ƽ����g�k����@�W�FJYg�XR�N�>�����{﹋�������r�dxxHZ�"Yvҩ�ն5+�6m�\ W��0��LLf��뮓�~�+z�P�[�`�x���������Q
,�eb��d��ݖ�7����9'&S7��eD(���z37��р�B[��cɼ�R�H��:�2Lm����~��ҵ�J��p��{�̘�B�/�!SZj�}�f9߾]d��[����S&ғ�ze��Q��x�Ý���b%6@ 
��(j��۔)meB� �����;��9˟����ӳ����?J���3嫷�ƺg�q
/kn[�[���oſm☝K�f�ɔ���G�����z��\42��W {�PԪ�/�=��F��e�����S9�u�M7������7�=KІ�x��Ο�K/l�)�-�O}R6l�� ����xP��Teۻ��O�x�{^����k�M A��$�����j1��`y@*��nw��U�0��)��w,΂��K%3̯S2�(�M[ؑ��mx-^���n5>� �y}2]=S\��ǇM#�зo�*�#� �1?�SG����dhdT�M>p㇥E�,x�����$֯_��eΗ3�O�0u�:��˺u��~ "��s�I_� ����y	�H�`�h�R��$�!�)mS���~70�<;u�a,�A(�9��0���$OHC(,;v�k�y���x�O�_�J��#E���{O�=w�F�g���0�|����W�y@���=�Z&�j�O�823�|0ڡr�L�z�iz��fB^�p��������۾cG���7	ooP�������� �ʶ��cCE���<O�p!�j{�����xF�������>�[7�I���b�� Fv�M�u)>hD�GX�/��NKK��C����HQ���A5b��w\s�<��C4CF��-�KK�U~��_���2k�,���W� �Y�t[�� s�f�s�vT��1R���;{��vZ�{˱4�L!���O~�����3����a	�)ȓN����#�u�$����}����Ƨ�U�z?��z���q���d���g?����5���7������_v٥l|SWW�����R���1ft�w���/�� �m{e;#h��:���u6W ���뮻�x��l�o�y2�@>D����q�w�jL�}Z05c�q��C��W_&3�̤���7��'�]����}R����F�5F��4�ފ�^�uT �2��hj�1��⋶t�>q�����&%7s� B����O08~�$��h#�)�5n¹CnSn��_��@/t>�e>��yݔ�D^�ͦ/�r(��?ȱ�Qr�Ժ��ˇw�4 =V="	ӦM��� Wr����轝�G^���Y{����>ٷ�i�
�k�G�Ǣ���[61 �Gi������Db�^%�b4��A�~yf�$,�+B�&�P*G"�:�H����z�J�$���6�y�T.�h�����4�f��)Z��:�9|���Q��a�ȇ�/�c#d�����?}�������NM���J����n���[���������m�5��:�!j���x�B�.����_��e�X4��{B��ITB��A�^=Ͼ={�]�'N������[ϲ�����7��!.X5��:�C�hu�3��ў�Cg�TZ�EOP
��<����~?6��-��]"�Ɍ^�J�j�20�����x�Q�mT �2�e�͝ohj,��Ƈfx��\���86C��p ��*Pf^���5=��jlݼ�̂
z
����+5��r�9^1mZ��Ur���6�5��A�Mw��/�,��>�Զʜ��e2��]=*�׀��d�^�?�A���b.:�>f��y���>q<�q����_(d�S�A8�����[ ���k�ԱV)�4�D/;�,
l�;0�"3Ɛ(�Uӕ��[A��A�������|r�[����^`h���g��SO�SFI\R���tN�U`N�w]�5�WABG�Μ!�_�^^����t������@�\s������
l[��9	oޜY2>2��p<w@(�5c����u{�5�����e��	骼!J��P��Z�*]{���Z�2�m)��:�0m#ѼV� �3{�L�!���_����R]g�ytM�6��J���p��/T�?�pȕ���ȿV�y@��s���ǎ��j����3wY���D7ׂÄ��_�ݼt�N��V��C��H�=��L=OB�Nʪ�L�����cQ�rC��_X���d�sރV4� w�q`T�����x<����*����z�N�!�P�V�h����(G&3�W�pmM�:���䥻ׄ֡�V�Po��\2c�,�S���n=�g ٩^h�Y�]{n6�H�:o�u��@oe���'n�ߝr6⮟!|�ܰ�a��<E�N������h�R����X7�L$��N������Ω��I�5�C&�Q�:�E<nlNR ��.���͞-;��`�,=}�S0� �%(�=�=��`���f{W�L���/^�0����{˥ihۇ�+�L������������5zKF⯆!��)�a������1}w�$�%,��3M$�����hL��Z]c��y����b��_�T���F�+�m���td۶m�qD�%�O7F�<�2Y�H���G�Mݴm�Q���&�;]K�)a��R�I����`%1:� C[� p�9hĂ�-)�F	b�)ꪱ��	6z�5��m�U��q�x���V���ʰ8���Woq���2�}��68��lx۰p��Ǳ�'��jI�^7���@�u�/�Q7�F�5���gXK�}K}�=�{�r�ˬ�w�=y���ӰA��#�ys�C
�_�P � @�ܒH�:�~Q?�¯��@_��2�l�j�����Q?���ǭ�cBBUKM-j��j�/\-����7�������@���~�I�
���u�XWKAT�1�B<X����,��a��|���e��s6�s�2�0��V~�l�t��W׳��*\�w�.�&4�����u�z_^��UҦ��ht���*���8����G:�q�����6��D��ɿ�V����dr�E+t
F	�O7Wt��3����`������ջ����4>G�4:2,5�uE����w�o:�1c��m��[�n��pHl��d8)��wA�Pr����7�X2h۩��%:�g	E�0|��#�>{�\�����+M�8вn;W��AJ®7�`M����e�Q�<W,��=/{�vn㬗.�(CN���Q,���/@k���z�u�
��C�?�t�s�m�T�[��^�=ֈ��l_�¿����X2+��L��nYtՕRLg�ﺚZr|#i0��V�Cy��)�#^���+����X5���|���I���
�`:Zb@o%�� k#��(�ߡ��2�0s�%�Ǩ�(jpT;$���ѱ��_��+�����1]�[��R�q�G�+�m�X,Wz�Lr�*^6� 찑�i��AY�4<;l�`�c�X	�g�w�I	����tJR�\��>�P���'J�|��0kk�8o7�XI�31�uFq��i�00�Zt<���	r�ɉI�M}�OA��B����7��3]��j�Z��1��B�zA�%:���S���B=��U�u?_=Ť�7F�k��u6MR�QF��Wj�a�7���9W�߶��������ڠN�v8���dK�Z��2�^�z�%��7�ְ��TZ=�0?Og3� q���ed�N�L�s��H�C?��E:k�%��?���/!S�ġ#��8�����B
�z�dR�_�N�z�u4�z��0t�D"/�w�|ɤ�A�nIn�D���fv�>���N0_��^B���a-Dk� 쟷�{�����"t��J���Z��������dE����3n	��R��������>c�VFe��Q��xۣ��:��L&s�"=S�}��5jγ�"�N��l`�{�F6@5�TdC�YQ�E
^Yx���[7�n�Ep�C�#˰��6�8͞�w���K�l��7邩A�(B���\$�p���%�H0R#����
ֱ�|s�����)��<D�����Ƌ�W-��߾ �I����8tN�xKG�|�3���'T�����9�h�«����DG��Uo{�(�@�ո�1�l.k���F��3��e�%��.B%Y���Ψ����X{6_,����j �P<k���>���ԖV���e/z<_c0�P��U���*�)���Ճ�j����T/|
5���R[]/�h\�F�28�w��߭b�����q��dB�eR����H��h�,�炪��4u��]�����a��A���9�"�Z�P)np�_��kR�"( x6W✲E�?���]����z#�����Dl�Qg�!��[|ά�L��5J"L;�u�����{��6I��k��k�O����� �)Y���8O���G[[�dG��O<��Z���F���i�ܠ��U +��Vl��b��S6� H����G�t�k��d2��wU�PK�s#r���&\���^:� �s�����Zt��<KC��M80
nU�5�v��Qz� ���!i���9�f��'��Mv��@X6UG�=�>yc������g�q��)����
����ڵK-\luO�X	�F ����Y��y�7mZ�`�T-@�0B�l��5DB�	?�}c��"4�}����v�+J�0g��'�����i���Q j��S��ĩ��`kkkd������XL:::�����;|�0C�RC# ��ʰ�]G[�E>+�*DW���x�)"
~ |��y}�*�O��涙R
�q=/쥗n�U�Vr.C��2�Ɋ���|q�����}��:�&��K�1-�f��F���������D�(��j���X:E���^�yF߯ںF-j \uŕ��X'�?�(#4����)j|U\�z�"��p�4����z��"a}��"/���?�]�m���`(y\��Jze��Q��8��[�pa�#�<���cn��Q�3����07�z ��v�0�F.�Gт�������7� �-1y�|�R~��+[^�f�JdX�\n�bm�vh�&��$/���aD4˴�3����v�':O��L�˶�[���ȡ��G�u��[&�,�T�@��oY ��w�sց��y����{r"�9��-������p����=d�תQ��?>/�����eyz�?�0=l����׌�n��~����-�?�-]����=��#������_n��6����o ��>�1~�{��.%X����(��~]~������/���!��ԧ�������Y�9��/��"���!�����X��`�*�*��{��n��ɟ��g$�-S䦛>*a[)g������������t�p��j^��%By���^qS���p��r�����~9|�0���>#<�J��5�&5��zlZ�G&��G�:���F����v�P_�����}�V;�;��{�{�$�,A�w��:���p�|��|���b)'�aٰ�Jik�h4+]]�R�V����T#��Oڦwȯ����a���œ��*�oe��Qy�*�\�3�H���eX^��!]�t�!��ysd�u�����x�����D�=���W�X��M2�� ڛ�.du���"�|Z7z�=�2?NF7�ܳٿ�n�M�w�����	v�G���=r��X�����{��r��7ʶ�q�>���=X�CGʝ��-�#�'7>� @j����w��a��}r�t�<��sl�ZRGq^t�$S@@:_�fs��7.tIK�s4ka��AI�e^o�OU9D`x<���<�a�����.���{��1Q㋿ñY?�������΀� �^. ����7�7�Z�zڱ�;�����hl2�B�h�jV��k6g�F``�(��8�Ii׾�.Fl��)ٍF-�	�1m�z�9��b/�6ly�q�ԣ�;26*�%,.+��eE���fٯ���ۤ,�(���3Hm47��154%f��0�\��\q�e|nXCD_6>��=zX����W])���o��Mʔym��� GO��r\�z�S�Ζ�sfJ]}�d�	z���\ �Ϝ�9��ޔ�i(ɬԡW�y@���=t��n޴un|2�vXm*�Oko��s稧x�����*FEΡ�d�Pl��������x,*O<�Q���K,>�R��|����5<��;)fR 2��j���1ӯuZ�<��Tp��RC�Z�F�YW�t	�{�A)HA{�	��
����K 4��_8O�,[���V�cE�u��ռ�k@� �H���NɆ���UoP�e��I��$�$��е)�� �L�wmPE���/��;����G�����������w��g�F�w����������P���{�5��uu|4���V�V����g�[� ���غ�e��/Z��!�.iD`��~6mٹk�d�����
T�C%��������~�I����+�g���xB7���g:	��,���и����G}$F�i������,�c��>���D��2�9r4��w*���R�U�.l6=�KLrN�]w�\p�
������l�b��f�?SD�w�V0/�E�6�eW�����S�����ٔ�����%����I��2*�F�+�m�l'N�t���p��f�t���
��?�Q���wѻ��7B��I��?�����{L3�����q���b�Jy�ŗt�N��9SfϚK��i����Z���.�j��Ҕ%H��f��O��{�>���+e���
�9�Q72_�^�|6�x���r6l�B�8@��z��\{����?����r)S�b?���hu˙��׹�"�r9���?/����<v@�["7��������� �4�)חKv� N��0��� rl*Rc�����px�v<B���h��n��v�^0���(�u�Ñ*�6"�g�`����}��ځ(�ɓ�jmd�����癜���j6a��p�Ե4��������LN��"�4h���^%��� ��;��g�bVoi�|w@Dd���T��7٥��·`�B���M/q����y�K���!��D-^)��f��XTF�b����Ғ�LK0�c��w���0C������؍KeT�y@���=Z[[s�-�z���-M^?ac_8��:qLڦ����L�ou��_��1<ޕ�.��w��Gum��G���vʻ��7��u�� >�����~o�9n��O#Њ�-˯��~/�j��T��w�)?�(A*�V�Z�*zy�O�MK��#�^��jÉ�V�f�4?���H��v�<OH.mr� A�Ćk�y��T)p��Y�r%�g�+&G��y�ү�^X�o��q� 5�F�A���C�H��y�Zem6p��s��ݑ�6@˃����|���g�?̃9rH�	���+�n{�;��r���gh�?����?�I���x<Hv]���=H�<��w��P�J=��x)]�H�Z=�,k�!�LH[�t����HMJ��`��;z 8��hH	�/�c��A~�B�z��kO���g'݂z���Ө�Y�o4|���AQpBP90:��B� �6�[0��iB���ys�3���d"I��O��R���%�3��󝆱��xG�����8���q.��p��~�ח/�^�n�`�c�۾��%O(�����%���OA,˰�nh x�;v�e�W��W\Cp���g$�l~�(��]��jwP��6��ޤ�3K�!��K�)����̙8�	Wɐ%����N�OfҬ��B�8�D,�\lM8"��w��VOMI�Vm��2frU�������b~��組drPԳ �t�������Y4C�s��9�K�ێ����{��ӫΛ�=X�8$T�f`���|��q>����t����w�����o|������\}��4>����(�z뭼����^�W�9�{B9߲eKe떗�6'9-o�|��S��bw�n?A���C�)S0]ѐ�/du�]
�x�rE��^���a}c�z}�ԇ��%�<�ɤY��֓j� z��0���ߝa緋/����ӝ�I�e����]��`��y����)k֮V��t�z�}^�`�����'#�Q�yT �2�e��U��z��x|��46dx4���K����̔�e�e`����k�`d_�N�}��/��Ɠ��w��1
��wv[�|΄I)|��vMu���ظE� ��!_z�|�+���{C��[n�K֯�O}�S�;��q�r��>ʰ�Wn�����H��l�E�6j��
���q���H�x8dT�p���H�^�_�����>���7����b�9�`+���$)�}�o��mذ�-@���I��,C淟�G� x�����=2��=� mם��`�q0�x����	p���?�a�P�4��ڧ��@���׫[_���w�����[G:���hiJ=F<��T'O>�y�Ǥ�O��fr��/�嫗��[%?��L�7K>t�$��뱏+H��s��y�d���� ��g̜ɵ>y��:rX��KMk����73�s��qy����(b�gS�b���ܲe+]�i<�R�P+.^G���ǎq=��8'��H�$R}�[)p��&�,� >z=�ʛ{���+!mZ*�2�� ze�큐�O>�-9�% H�X2����.�|R�@7�h4.C#'eՅk	v㓮�3d�.cI��r���ɷ��=��o���e�{d��r�UW��Ȱl|�19tp?�Q���R���z�^5�̃'�uk�����A��+VPS��w�K��أ,k�>�eRS#/1�Wx�k׮%0UG"jd���g��7�浩
��E��!�c�e�<4�|�۷��4�C���Q~�� g竩�����z���#�s됐��̰9�����_�E��ܹs�@ �,�cl� �ED^x�j<��@�%��]h�)����	�A�?���;�x!�Dn��~��r���a�%�mX�|�t�:&c�잆����d��E4�}ة`������_��+��T}f��|��o��/�R:�������?"����\y����}�ލ��c������N�w���+��52ej��{�]$��]��>��쥗^ʴ
R��#�� ���{��#ᵫBq�O@)��]��v�RC!%S;�$��r�HN�8�sm�r^��^�}T �2�u�NW	^�GA,��Wt��U���a��.M�w;�c��u�F����L�U���w����uy��G$:6.�m�
H,>n���<&L��o�Ac� Bκ���)�b� lb���#�������~��,:�A�ddxX���os��wN����y�/����K����,v�;7���U����{���,%X!ߺc�+��w��f��4��V� p@6��,��X'��W#z?lA� ���]��/�`H�������@x�8�9������Gdyp����.m��n c�l���*Ќe�����.�L�'��a��3�<˹X���"P�����'%�T`��������_��Ng����뮗��u���i�>x�5�����ȣ?"�\��!u�ȇ�/��|����;���7J��w|�A�:uJ�c�<���x?�Fx�=�(����73ʀ\�����ګ��a5D�L��"_�kw��A��`��y��]I��ZԸ��T4��zQ^۾W�	5j"2�H�2*�<�
�W�9�;X���Ka�yII��{	I���Ț�6�Kͨ�54D���� �6qR���M��{%�W��/~�����?�/�:�&��ς�~��[�%l��V3<�O����&�����oHl<�\�S'���,�?�r� �D,�F�G7n��TE�<q�j�,Y�D}B=�	(q�(D� �9"/�d�B�E�x�Ϛ>MZ�UArphPB���.���A�kb�r
��;���߰�y&�*�nx	<`_�^���F���[⚸K��R��{��k�/��r�@�I��1;o��~Д��wX{Դ��G�׵���S��W&��hÿa��cG�\��PȩϿZ���;���d��t&bI��V��.��xB��n�>�+�֬��3g�z\�.}���ky����� �{��d��r��A}W��Ç幧�f�;��u�� 0T�n`����~��7oz��	�F����M��%Ԟ��ǥM��d�		E<r����n�8�^�?�3 ��Sv�ث�_�^���R�q�G�+㜆n���pU)WȲ,�`ש^�B�ٵ{��������߬^�@x� I��M' ��ƍO�c�="�Ǐ2g�m�Ay橍,7C���3)vZ9W� ���=�V@��b# !䋰0���<�Q����A�ē�6�y�U"��9�y�7<6�{D������=���d^�#5$����g%><����H�㓆p��wz�t�˔�����6��!w��+0l��#�`�§M�N�5���z�y���Y<c(��댬_����.]o/$QsF�=]ៈ`�-X���nGxv>��9A�aD���Gc����U����@��5��O��
z��t����c��Le~=�H�G
K���}j@������>�9�Ŀ���Ȼ�q�$&bR�}�kx�D\�CE5���U�*}��ɠ�>��{�K*���}j�>uBЇ�����(�(��
���j �������Ts�!�N�*)|�0ŉ��e�+�_�&�V���QN�R��N��8#��t�ڋ�ʡ����/!�Q�yT �2�i8���nҥH����pʒ�Nw�&y�+�d��X�mk�c�Ǩ�
3���P��+����a|rB~����p\Aʴa�S5�ނE�@B�_7i=��Z�~��Ϝ9-���*���
�����z��˛����ydlx��XlC�k��F�=�y�D+̡��O=K5`-�z#�#�^�hm
o#�^�m��Ǟ��ߔy��5�m�܎8`�)\�n�s!�a�PALs�9O���d����� + 1�7ae�f��� p� ��ڹc�Ug_*���1`4���Юk�<Z�Y�.k�r���)H.o���=����u/^(�N�f	���(������!��׾ʨG@�sh�>z���:��-_�t!'�g� ?���K6��}���{d��9����r��!^���#�/�������S���6J�m�`��=sv���D2ٔU�P���zQȱ�Ȏ'�.5B����cR�����.I�2��%��]��r��K2��ѢTFe��Q��8��(8
U�@��5X��1B���X�R?s����ꭍ���db�3Sl7A}8J�N+���FP�P�'@����^��EP�2�|_��רQ>��Wn�� �I&dHAr��e����Z�������"����Bi#�OŲ@HN��y@`$�W��Q�Zc�\R�\/�PS�^5�ﺰ�ڿG��#T�{�٧M#�Y"��Ҩ��끐��v���nwO������~9����� ���)΃|;����]�Ʀ&��Ǝr����>�bx���o����7��^����:�#�u"hI���	��y���c���Le���)D4��Aܮ"��@h@��ӧ�ʮ]��r)f&����!/>���S	��w�Apt�����d�O�p�)�鏾C��J�?��K�բC��e��I��3�}��!a��h@��H�s������D(�y��F�t�Q��8.oI�./U�R���<6$�J#|�!py�?0�-��OIu]�d����8���qN���no��6�nʦ��9+$nJ�|^S�+�u#�r����!;�͖����	�ֶ�S/�.���M&&��ߡ�K��z��x�4-Zw�W��;�2{�<� �\� ?��_�m����=&������fMѐ�X��mjn6�b
Dcј\���z��;5�Yu�&u��Q���D
����i�n�`{C��u�ֱq
��dє���:s;m`�����Ϲ��������M�X���Ɵ�������
T q��e��x2�,��- kww��T�ӵ�9G��X���q^�Q�'85�hЃTD\����4JvY}��H����b4�2�s�Ёߴ�Eٽk'��{�G�(�Z������3�?CO:�NP2;{w�.�_���;g= ��/�G�����	Av7�����:u��]so�أjat|��@S�H��k�XM�y��#AGX<��#���k#|�q��������	�q5bgϝ-C�c���2����T�qN����
�*����
óF8�^ Ox�B�aq��&P�Vw��
���}A���1l�̱;��e�ӂ����T�\�����Y���=���mV�wu�f�0��0�=^����IP �����MM<�k�3�A� 	Y�ދϫ����pL��ihi�l:���^�ð��$O*�{�^�~�"u�SP�g7>�����~Mz�tXح�h,ǑCG�F)�uURWS��ٺe��1�N�:eB��W+����:u .8 �����a���!�ŁB�]O߀�VA�����Aą����
���!�:�ƁC�:�(�;�n.5�z����`
����pt�hc�_AzP����KC�a��y�}F� `
T��q���(�>�����\S��c�F�z��iG�5��ޏֲV�^tҼ�2<h�F)#�}�x�;��Q�3a�A6����[ �Wr@���C#��n�D�h���g���u�VY~�J�#�S�q�G�+�<䯍��!��0���]^�	�'
IO��T�r:��TK�fyt��wˢ&�`�N�"�mT٠cr��Po�vR7^ 8r�v�4����y�u�v9��.uKe��Ùv=2A2o:G�N+��䩓���1C>x㇌�i�l��\��b�}�ꝁܕ��x\~���ȸ�3��U��T¨�Y�l �݌�n�b{�8[�T�f����		����S�8�����$1��Q�ෛ���������L2MC������ϱS�[��L��&����7]<t-3y�-���j��q@�[�"?�pX�I<�b��-_����~HF�Ǩ��~x�h�:(�ć�M
�v��f
��#��}��w�V���0l�����=h�bB�����GD<��u�>FSH�y��)���cH�(�C�����e:����;���낮�n4*�(I� ��M����*9��8��qNá;g&�*a/E	{�뮏�+ ���P'm뀧Ha7K�!�nt^�F�4��,��S�9�Gۻ�$Py�!bMNNЋB]06^�b��O�DF=��H �
�u�uR���ʇG���u�6��ୣS6yD֬Y�?�y/��靎���7�<��߽s�n�.��}B#�aC�O�V^#��^ѽLs�?úb^�,k�̡T����b���u���ڧ�~�v��`����1���#ɉ8l]7K	��'��U�@μ1DUt��N7+ `��~�(�̜%�(Ӱ.0&�Dr�LΩk����o�1�<u�i��Y=�'�2S����V���_HldL���;�)�hl����%�d�S_����9vڅ�%�"fg�)پ�5��z/(,��\<������a��%+@
u�#xo't��<\�2��H8(Y50����@�٪���Dc#$��pҌӤ��Z&��aoU%�^�}T �2�i�|��n�dj��^��%��ƘZ��� #4� �9�*�ON�x<̑;�� �b�4B-KT�(fV��F��v��y^�7��o����!S�?#�/��BZ�zmPT�wjÐ5�3�xy��z�����%�F����=�
���K�a ��>���%����Az�H #�Ȇ4а�!%�<+<:��]e��mL 쑓�����z������7����*Lcׇc�@C^��a�l�ܘ;�Ɏ�&Y0�蟞R���� ):��v}��.�<��� � ��.p���x|&��R4��o����/�ۿ�npjd�Ͻ�wѓF{Q�s��:%����R��R��F+Hà<np�_��\q�r�5W�e���X��A�|ꩧ�5�t�t���<�?G�[p.�" _^8	��|�d�z}/ۼ"
6Sc�$'�RCI=������U�b�2�>p�W�mWcb�<te����,_vA��2��� ze���M��K)� ��-芻��\��d9K<%��0̉&Qv�2���6��P6T+�^e�c����µ���cV���<�3�� ��R���w^r27n`��t���И<���z�4��ཛ�9A��x�)SZ��7HmuD�͛��k�@A��;vJ_��ׯ��B5�)I�n2I�V4h�����<��C�����5�w�e�\���v�O��\!���#a���Yo�H0�q�|�;ɂ���?,##C$��E��V��P{~��W �n�*�<��Qq:���p.'���Y��ϮI�P��t	�"��n4�ry}+Jzl@:,�j�L�"ߺ���^�������i��{t�y�M<�enJ���(��)���g��CZ�J=�^B 9O���A��xh��|�5�]E���2sTo)��>��)2g�,Y}�
�={&���^�B���?��N5t��	����Z���Z�1s����%�:�]�_�NG�����t�K<���S��JJeT�y@��s��;��1��
��Α��l$N�a̪p5���=N �&�P`+2�ij��7���8eH��H�� 	����S�Г7���>�����l�lPώ�;F6c� 9@%n�q����v;o��z�*��x\�z[�������z�	���Ua���R��x�(���QFV���(=�6P+�Ovr��
t�\����Y�x����[���׍�@��dg��_�9�R���+6�	O�%o����]G���'���X޵�g�i�8��sZ��wpxHR���!=���˴3��5�ՀH��:9��بz��I$��e
Egҹ	i4l��FI��(�z,;�Y�yA��Z���9�Wa��9ϒ�+�G�cr�ĉ��=�p��D`�y��>��>v�sy���Z>��O�qYE�fb2��b�!",�� [(ɂ�sdZ[+K,s9}GC~iW�*61�?q�7w��~������|��W�{z��2*�<�
�W�9IW6�t�����Ml��Y�{Fg��s�)�6��9�َG�}�v���<�65��u��r���\��}��YR�P/�bU0��i�	o���$�
�)�}�\uܬ=�qMim�טͨ�����!e��O/.�𱛜0��zp�_�PAtǹ�PF5�}R��/��^$�-2���ǏQ#F<;�."({`��z"�*{ո;]`x.˻4=�kk���GdӦM�� ��b1��9n��F�^9}��Qf�5�2����`��c,&�>��!���
���Z3�]��ᱳ{X����!֖������a�Ľ��@���t����"C��{T����������=�,ǆ>P��g �`�n���K�y�yH�xg��������}��3��:�IFIJ�3  7�6/u�N�4�k�e��7������tK(�����,����~5��̚�������e���a}W�f���E���q���Rэ�G���D���9*�^�4��#\]Ŝ9�a�E�0��eXx�����W�^)N�S��W˚��h�H�"��ӟ���?�u��,7��nz�(�Bx���Aw�b�{� ��۵�بq.l���Px�ؐ�)�;������gJ��3`���vK��_���(�z��W���/c�}�F}��ԩW��|`�OH��`L�Ũ�=�B���k�j07��@�A�4 y�; �z����T�!���CKK3���s�4:��bq����J
�t5�z��G��24<�P��}��]TO��3�2b��Q0�HQ��a���5�:���,k��i (� �&[�R �K뻁���zy�R��T:cU:LH�J�%g�P6�gmK�ڑ4��c����ߓ�4S)N��T�;������u�XpJ"��-������#��)��l����9�tH��q��T__k�%�r�UWHuM��IFr�	���J��.l��S.��y�Oˑ�G�3�
�W��@��s��ǡ��^*���#�v�*je77����n4a��z,�p�G��;���-<6X���%�d�?����1c�n�Ez��O!ת��*��ɶ7j�\04"7���N0�ˎm>��|���!�"�@/�z��ЎՍ2-�>�o��-�}2w�
)�|�+C��F-K�����a���d<F���t�5h������$���6�3X�g[��-涇B)㡎x�lx�$l�r������u�I3!��[[�ȡ�G��� 2�h��g�NHUu��}�F���/��1���p�H#,_C��[�X�t�M�w��ߚ���:eϞ=�O*�f$��������uAR�n��e��|AFF�e񲥲h�Ry}�>�%�H�$����|�h�w0�p> ?J#C5U�Ԁ_�����AV���(��c�l�#��r&�7�#�]wݥ�Q��^}����ʈL�|�Vq��A�B]}�����i���&]�2m��3�E�9Cv̢ٞ�P�[q�R6��vJeT�y@��s U�'<B�E�[�p^~y��x}/	\��;d��7c���v������m�y��C��=o쓛o�Y��Yq��?�����I����9~�(+{��{�f�]^���6���nɒl�r�lp��n�MK�InnnH!@�IB�(	�H��ĕcw�"[��Q�hz=����w�����?�3����~���9gw~�k��%�;@��T�e��O҈��� C�< �R�QZQ��(���icE�T<�2�dϮ��w갸Q�X�Z>(s,�T2MvC�1��(��]Ft_���"��ֿ|[~������>K���&�W�1m��Q���F3� U)�1�k��^c�1ӌ�Nv��n����}g����0���"�0�˞V�?��  ±�y�ܹ�t����ٲ�*��_���/��;�����fd`pX�� q\���<��ȩc�lIus���EN��!Ȧ�cӡ�@��K�}�(f�;fϒ
f�]��LJ����H${ʵފŋ�����I���k8���p�y��/T�ӄ��[��3��w�&o���X/%u �����o�o��5&�ᄓY��d벥dD)e玽z=B�v���<cA�i�̞�)�y���p���y� ���%�Ѫ.�^�d��	]�P/�	f�W�X�1���!����Hg����P�p�<*���g	LX�1Z��楛�dp`�$1O<��<����ls�tg'b1FQ�F�,�H��tՀ����Op�Xt�Nh�|	�f.�Q�:���#�f#�'�o�
�.u���@fh[K�v̯�XR��j+j''���9���g"� hQ,������/�G���g��@.pQD��;ƺ������a���'>��)��q�=y�)���F��,���;���!�Pmd������w����;��F������}r��o���w��~`��׼�g�(G#�`\�F5J��E-���9�';v�欶�rIL�/�=D?J!x.�͛C��i�|`kCV�\�0�9�a������s�.��sX*$!�S�͍R����䝷�.�#Cr��t�>%+�.������R���'��,N*�$�0�!s�.�#y��af>��I�y��019!Cz��L�&b��λ�،L��Z.U=��]wJT���e�t��MH֡��-,��
��+h �C`��E`�h��'Oq�F�۳:g��3ݜs�xQNh �l,�b�P�c�R�ZE0�<���+�a~��5B"Mmr��q���#�pԤ��9�@c8F��ZJ�����j�d��Μ�%x 
D�5�����/���d�5�vq����-����=�|�r��w�#��k��NN�� K�jS�#x�ǽiTcFP>@������)�h�l�>�<R�h$�8 ��}GHނsQ0��MO��kkk�|�C����wHqrP��~��'6]|�l\���g���G�H��@y[��;fu�r��'�Ͳj���$���`��z�i��Iw�)}^\Υ�Z5�ש��3�R��Mfk�/<���WG �I���������z�<��G�'�ʭ.^�@��I��L�NW��d떫����òb�J�sDc)�& ��R�	(��څ��۵}���9��%�=1���ԂLՠ�y� ���E�9����뢚#���ji���QY�d�Oh�b
:�]]�LS]�yy��(����_}�e�Νr��k�N��V��o�^>�������������
E6�!U���Q-�ϧӣ�M���ӊ� �;����N�^�n�ē)C�}t+��0�d�"�N�Mi`��mDA �FUNd��yT{�p�juT�ə�dc0�����o�Q?_����OH^�)w���r�Iֽtx!��c�ǟ|��e-�-������~�C�y�,Y��Mz�;��x\�/��/���fy�Ձ9"��ڢޏc b��^~Q�>&	u(�u�Q��y�0DB
lW_%o��f)�)U�E�ɏ���ޓ�J'��+.�+��T��:"��qM�<����[n�����t8.ڴI>�7#��x�Q�;Z�|]z�&ߊ%K��_��|��T�;�۽�-��e
�;�T�!��nx������>c��mo��(�앧�~R���HҰM��OL#dF��Β��v�:|�NԜY�����%y_P"@�&�I3ˁ����4�������A�a�,	�_8�~�"5�ŉq��w =�Y(�b��Q�mLCZu��%\'5b蓪FX�7��Ex�4*�  �HfY�r>w9��,����+=���[�[e��9r��I���2�B*�)�֭#���?.���gYƼ��7�\�F��t2�D�1a�b�ۚ��o��Ψ�嗷�O�Sը�l�P>|X�{�oˢ9�����{HFsy�i�ɴ/uZRG�Zٰ�B=�a�;#�(0�E�B����G�f2�!��q�R�@�{8
h��KLuh���Q@����&��zdΜ���
޻������.�T��O?,��ֿȳ�>ˈ{Ӧ��7���O�3��W�{��=﹓]�]IƓ��ϗ舁;=�2t�}��l$��@u�ת��Ǡ��l�H��h6��^�QF�W^y���'���Шދ��eP�wǬv�ù@f���tZ�ڷo��3�k��2ݒ��t��3��}G\u,P�)��G̔����(`�WOc�"*M-�
�	鈵ˢ%�J2��}�ꬡ���B�_2������o{�:	o���1D���u�F��1���-Ȇ̟�rRkK�F���hLv����@���j��;� z`3�����z��XZ�D�����v���@zߩ{���Y�FF9��g�NΖcj\H!$��u�]t���\sYΞ~�iC��������i4s��7����x�a��?���LoZձl6_s�{���5�b꾜'hΟ��)nl�h A}�ca��F&iu|��{�M֮X��\Z�.\L5�R�0��p� h���Fd���0���HԑD2BSS��_0��k�g����`1�$J8ac�H��;jq��})��s�a���b!F̔��e��R�̙��}й��3�ŵ�l��T8����)t��#`\�b>G^}|�\D�C��ǏvɂE�%��܋�	Y�p�:M1�3:��}���:���������gg��ػ{�l�t�<����of����W�ftxX��G���˖������� �Ͼj�G�Ȣ\}�՜?_�z�̞޳h<KH�'���#q���"X��{�Iu�z�<�[��6���H���� ߩ۪˴��C8�0wN��W���H��>y���e��#z`��(�SF�$*�{`��@l�(�Ԛ�ܪ'�g�ʳ�|��2h�C��������m\ ����ܰQ,bc�ٞy�{����4^*˷��H�t���^6(�7=��<�HE�d��5�f��t�֍��y�$/��]�ek���j���)�jtC������/�$�/X+�M��F��w=k�/���/�U"=;2��l�,���G��+�x GM�#u��-���8���
.+)h���=F��3� ;�*�ؔ=:֑) "zň��`V+�lRko��hl2T��,S��&(�<�0t[c���c��P`^����N	u���AW<��\�� �1�1�>uZo��K��n�Ɋ��HGM$�Q�~ %�2��Č����/��N��?E ���^�:�#Qyeۋr��G�v���X/�dT���Y���vKS[+�o�م��F8_���S����C�ɔLf����3�P�����h�x���c,��*m{�En���`�����ohh��:��x�2�ݺ/��ٝmr��O~�l"�����g���@R��x�������+ ��Λ�،�r!�R�R�t]W��t�8���F�'uq��4�� ,��X����m W&����(]Gh�G|�T0���S�r�`TŐ�N�������o���R�������={X���Q,�ѮF�al�5�iO?��̞5W�{õ�~݅윏+p$��F8G^�	��g�S�dǞ}�J߰�"��O��]����ȏ�޳S),�#�>6�MH�����Y�x��UKK�d�\3�gv{��K�T���G�/4�f��u��w��9l̾�Y�4��HA�VG �Qu{kIt���ǥ0����80�U9
�Q?�_�T�nz�IY�'�idȈN�WxL�x�F�)uf&�`�PkBA3�ǎsU@�;{V��eѢ���ϫc�A�8 7�t���9:�w�D�Ȅ"�T�h���2�ɤ����qlom��:|���D����s �t,%���作'�����hw���Ks]�6ކY{��~dǳ
�f� ���A�D=��!���R2=�ْ>�!���J7���䋸�)��-��$�����3�<)�����X`��@lF����!�C��(G�V�hqb�",n����M�A��8�p��2�nbjML���-AI,j�سɇ	���U=_��B�rPu�icX�.�H�N(����r��A�m�V0h��@F�o��;�ˈ-�J�a�7[����G�~vpD����Y���b��͌�!*S��n�����	���)�����PA�����`�42H?�,��J�rd �����T2���Q�f*�\�r���(C�u_d���Ld&К�v1��������x�N≌O}k�=R���!����1Т�,����z�Ca���H��4'�9�4�+���/��o���w�/���D:��N/�ߢ��?����@^���?G>j�(W�,�雜dv�����E��욦8�;��%�#��
(�5)�q��1���f�h�ٔ�3=<�L�0�����J��ƱD������3��>��;."���v<��8�"�-TX��lsk;���2�>}+	,��d�6#S��WJ尥´�� ���X ���ъ�.�0�-=�ioD���f'�.�!�����oh��<F�%/8��@�	Mp�yc��\9�9<8D�EC����B\��Ƽ�^&f�*�J2RΫ��ՅuiS{�2�M* �wt��<���f��6�����'`oٲ�s��
���jt��#c8p4�Ɔ�-�SG5µ:�pF&'rr�W�]p���wP~��g-`0��s$�T��C��c��)�#�����g�=h���,��U���m��W�(wͺ�(��XT]�r�@�F��F�h�{ߝ�+/�,g�X��nb�]8rW��;{�Bɏ��|}P*���{ꩧ�ȱ��ַ�C��[`������]G��x����b(|��ᬠ[-�秊Y��,w�^�&��9р2�>@pH8g_(֚���+�k�i���}�x��O
<w+k��*x�"pL4���>���${��(�Ye��+K2����TM�d:�X��o�(�v�, ��fdCC��
�q�+�P[�LfX�h �I�`���"l(�!�I�vGC-���[q2��J���� ۙ�"����Ξ�ś����t��ڌ�щ�"��S��g"��R7*o���2�C�skG;���5b�(��ϥ�t����avm#���F�C���P��B4�f�J�#�Gz}���,)`� =��������/{õ�ʃ=$�3�^�n<i@���-x���y����=^��-X�Q�$�/��X}���)un
����)�'�7\'M����[���N��z��-$Zٻg�i���qL�ΐ'�S؄�>�N�m&�>3�:�����_�lꨞ7���ٍ��&=����%x�9�� u
Ǥ�.]��ԁ����ۿ�}t���^ukǃ��=l*̚�U�|G�R[ *��GĤ�j���ngt�5���:.��xNI�k<,����v��(�d��<��n�6#IV*n�\�0��t�0�ѴƨiPr��1�����uJ]���M1>|Lf'��I"�t�ˆf��c.ӹX4Ѱd8�#,ܖub�2�h<#;S��jHas�M#�R�8!HU��w��Ȱ�-W�g�Y���m/�Ky�ؿgwM4)al��l�ȃ>�q ��W ��k6g�K��/��'���y�3}��ժ�Y�z4��I{��2��"����a���K+,T+�b@].$�C&B�藠�0��qT�|��Br\J�b���7�ճ� �Q7:����2�S�-#C^]c��]���CC#r�=�2������0Rfo�kt{�0Y��9?�7���c����̀�T��D��e"�i䃳X�j��mæ-�ཋ/�X����L�O�R�9/_f�$ �B�sd�@h�T�!�q$��@�i{/Z�s��4p��I��7D����%��� �;� z`32]��p����d�B��� �KɊ�
ծ.�N��Ya_Y,�Q:@!�Q9��W�Z��cǎ0{��A�@�>�@ي��� Q4l� X{���l��`!��E�Z&��E��j�k�<<2���)z��F�Jc'9꼈��	5]���S'��g?{��ph�CP	B���~���|��G�n�� �����6>c"ư�@*�?��qޘ��3w6�p`PC��Z�[�&�n����v=N��"c_*Uǌ�پ�7���`��`�|V{��Fx̨���U��� I�7v�}��_�'ٽ{�̞3�]���P� '>�讟cm�p0p����@F�8�+��L�9B���˧�kg�f[�S����ŀ�����)X��)���A�)P�gY�l��L��w<a���P��FB�?��ې�&	��*�%�lh��uB���F�#_��FB!=N)`�y� ������"����>v֡���夢�$u���ʦǙ��u贂ʻ��n֣1W<11.+V������ޟ�޽{#F�\�m����<^r�&9}���BHD�8�Ijr��F�ji�*S��.�K�[A#ׁ�>ٸi�W��(v���|�{X��t b����u��O��]	J��3��������[�4� D� Iht�v�yp&p>P2kЈ
h(?��%��hif��sĈ��8��Q��9�s�(�R'L0��:L(`��k06�K���t�4���'?�)�#T����e��E|���ַhT=���{���*]4���D��O|���3OS�i���
��V�<�c�RIa"!F� KL- TAT�h `���=��1a��U����8w��H������F?[ú��F>��,?�q��*���/�k�
���e��&�xt��@��vuD\�~��I7$d��%�~�ξ��q��|�}��<Jj�T�EܭBAZ�=1s�v�, ��ffUÂi�h(�8�"M-���x&B4���Z�X�E7�9b���N�x�F]w��CFTH���> W]��ihHt�s�h��&�}``�@�(z*�77�5noF�јQ�#0�3R��6I���.��-;F�,5*��l�
��z��F��@���wH����ui���{@^x���C��n|��K���u���Lm�� kP�^vŕ��1�#���?�q*�}���y�+��/�h�8���+]]]r�eW0�],�(��	�����E6����@��ɧ���'N�m����/|�w��&L�669��W�D�z�GDv"��ǰg�F�8p��F�?F�j�|��g������|Ե8>�;�<ܲ^ע��1N �3<:h�>�
�I+�cAc$@d4�/t�{b������խ s��J|���]0k��q��Ȝ���ڌq�3��c����|���38IF�7���W^*��. QMZ��&S.�喛�s���<�Գ̮�A+�X���;O z`3�H<�4�5u�pu�z��Y��s��ֆ�ܵ�M_!��yaID#��~��y\���A9t�^�)_|q�\����k�5d��Ms��t�",Dҵ�d�s��E, �V��n,�`" @� R����/VB'���b��n�rG1�E�s��
h�bW�;���L����A�u<�`M���n[�|�H}c�d'r�\�I0@�h8�f�əguVp~ ���p��?�����-[��\iZ#���,�L"q���(�|�*��#Z��l�T:��o�f��]%�e��u���Ѩ:_zݲ�㤾����e�~W��PP��j	u��r�	6:���=8f�Sr��έ��K�ٔ��76�U,�~����	��104�����ѣG����@V�^%��M�����Q���^ɛ}�g�զ�A�J��\N�OJ��(�'>x�� hl|X��8%dA����$_��7�iA��"vʊ�K�h���.�,͍ͬ�GÞ,Y<[>������?�}�K8��E0�[ ��Ț��A�AqԸ=]��Q^�|�������PJ������}���~��jݩ�&lQ�C
��!�h�QbwL���Ozщ�1FW�H��Q j�gVC���8��ś�G�,(X7n���jH]b��8�T�Y�.��9�5�c�l8��!n"b��O%R��ҪQn�������؈%F��4�Utq���?L����o�\�ϛ�����p�c.\(����$��7�����%�6˩���ǲ�+�myWD�W_��b.��d_~�ev�#��3g�����Qx):\h�CC�Ui.��靀�y��|����q�Ӣ�k$����s�������1
o�ZF�dULD�s�1C��{�0��;v�`#�W\�y�\!/���+u�[�x-�3<ds0Rȉ���l�3J�9u�����2'(���Y�t)�W׉�����7^w���'?%�7n`drb���p :;gK&ݠ׭�P'3�)�\��g>��w��/ex��Q< ��j`��@lF���G"��F[��"-͍�b�
��+�P#"qȢ%K�����~��ӟ�������7t���۷k��jX)���aini��{�����Z��멄�hż��ƿEfЉ�� "��e�]&-�h�)����{X�;;��jGY�'���NNL�.�&),����s��~�UH�L,#xW#��$'l�'e��Q��x��$	D�}g%��0�1�q�~�6��8��\V�b�̞5� D�k֬a����i���v�7!��kb�JP�X�d�tΞM�ji됵n�,9�߆�F	��f ҆�=F�|�م��av�Á	�c��#�A�E3�`$X#��2�X�k��o�F�l\��{���Z�����H���stv��~v��C5<8hg��z�8A��~�Y��7^�^.X,s�dlb��hQ�=j6H�6��R�Ѩ�����:�[�v���=æ�y�g�Y:~��/�%h�oVǲN2�zO�;;$��#��>�A�K%}B��\�y��^�V�{�e}�J��a	,��h�6#�帊�ꢹ�!G���s�:�Zo[�,�5�i͸�_>[Tp�S*���G^y���.pFV/��`208L�K��$�	x��Gt���u�XPmDgǘ�Dgk�
g�_q�Ul;��+Ԯ | ,��f�/_*�W���k�ʡ��9�擺��Ă�Uy3%F����bDZ�Xƿ���nے� ��-m��1�~`D�VČ�g��� d\d�q�9�t�M�<�ϔ�^���z3�mJ�Z�o�F�n�J��h�x˛o"�;g�Qvn�#}��uj��^,�!���F�$/�DR�dC�/y8�d547q�+�����0��{
p���6*�cy0�+���8G�F � F7����L���絏����<�C��Oɺ5ȩ�]�6͎�`;6��Ʌ��:ijm��;wȏ������[�T��:*���o�����'x��r�lq!�a�-������R#����u2�s�,�?O�Ι�N�^_=���V�cO<�RR0��y� ���%҉�b1�WT#�ʙ�%���.M(�
)���)�<9|p��\IS"x��}���e��92�8ñ8�,��I*S-K�3jW�FG�����;��)xl���� �u]���9r��p :"�|���x�ʉ�,�94�%��it?,q
��pv�Ԙ��?�t��D'��Ҭ�.�E����:1����J�ᣣ�2��Iƣ
������a�H��8���GĈ�}P�r4���?\GP��z��C�)r?r�#���^��78%���}\+��q�t�[�9�밀O�D�N�瓸@�!�>;S�јߠFAF�ǻNr����(�Ȏ�+�s�O��6u�&}�N�͘��2R=�}��ҷo��R2'N�6Y�f\�\k�D� �=�+�?�{��!����&9����#�dr|�R�84 ��&u��&�������L7���P�(�DF�X��5��H*��?%��Σ�،��º�c�)�ʙ���q��KǏo�:iji��0���L��9g��Ѯ�
zI���7�����[~�ིo�.M؋��5�b�̶#�}��eժU\ı�#�j�1����L�U����h���]{���X�O��0��4 Q1�lk6���Ƚ)�9?en#N�\g�O�aCւ�����|@�Mt� ؔK��O*��s�.���q]+
 l+���[�qb�+W��[�+#w�v 0�u�i{��V�e0U �Җ�V�(ͼ<�gѩn���Q3������!S$e����IȚ��F�k-������q3?ڷs�8vԶ�Y�q���ܑ��M�}�������b���;b�����}}��fs�ф����P���O.��b����:O���̓Oȿ|��2:8$�	Å_��I�������#�Y��T���g�_o��ޯ�+��JH�v>- ��fd�C״� �&��E�� ���]:;:�(��94�/���e��)���?:��)����F���rՖ-� t��m��k���G�%IɄ?g�IQ�J\H�����ݡV!��qp*ȴ��@���ܳ[���J�mG'�b>d9�6vz����=�?�]���V�&�c@��;ߦ��;��F�9���Q0;/�� ]^e��d?�4:D-�b ;�Jc�FZX@V2�xz�rc&��:�""Ih�gsct�%iI#~�]�U ��q�r���c�ۙ��.�B���G�C�[�����x�-p)@×�fY�l�Ť�iiie�:���T��Ą:g���d��z\�a��yWMt��Z��q���Эٲ�uĬC�ϣ Uo��6l� ��=�vJG{�\�~��~��T�{�'�J]Z�����i�l{�9�xQi�5W��3��G�h֬&=�F�:v@Nw�D���!	"��Ϋ�،loqĬ����>i�kT����I�?o��s;e,�;�N�9�߼��|��o��_$����P��x�ER�Jj D~�_+�J�kin��E���`xޱH��cIy�2f?��3��*���T6�G��x�G�UC��.���>�N���lԎ�7#t��Y����������L�S)k���k�7:6̨]��=����T�E�H�'ň���Fi�49R��M�{��Hۤ�I،�^ !��k���3�NK�١~7�Gb����Z��#~$TeD�T�+�XF�:ȣ|���:<^864�Q�G�q�ᘠO��Fr=0�Q�M_p�U��8��x$���ɮ�^�����V*���L�>�{�P�5���7�s��/�����Ô䝫�W��%�|�e���?ȴ��c���L�َg�~B2��|�B}�]
݀6��{�g�����u{M�F�A�{`��@lF�'���LV�h���Wf�u����ua{A�����HF�ޓ�9u�[z{ �bɕ�ƸLd��,^�X.�K�E��wJ�H	��tS35�㺐C�
فx,E��2A�
pD�gN�HǬNu8b$q��H=������qv�[����Q����6	KE#ّ�A֏�~'=���n�vm�L���7p�cp�[Ǡd�:!�
p�1�8�w}j\|����ıcSLx��6#p��s �2���>��O�;؎�7�憎����w���Ԩ2��T#��0�v&�����%�/���@�����T�R%c`��g!_�;م3��vg�nF�@�K�w=Hp�G� ��!`K�p��'�ǃF@8^�zߠ����45��:F�=�H��=��K�#����:���I�+7�)]�A�b� ���W��:ҐNq����I���;���$���)xp�LVdpؕ��Cr���'�b%O:ڱ�Y�r�t���}w�{��~�+�L���"�h�̢v^- ��fdH�c��^4���i���֨k��6čhD��?,'Nuˮ���%�8fa�XcM6s��Qmm-�JӺ���9}RJ���ڕR�F=
gs��P��F.[`g4�ЬG�����N�l��j��>n';9�����q��	)\(~a~�z�D�!'d��9?m��ac�F�F�ly��C����{��� %# �(��(��#_˴f��:Q?�?��ƖX��n�|x�~�h_Ɵ���������k=I�� ��z"�s$�o$j�������y���|}v ;+65�3�v�U�̀��QN��b�����V�lN<�H�E�w�pP�COz)쬿�cwL��>��X�`],��<��:&C��㝷��D(��D���!�T>�-9u|�oX+k/\��϶�6I�d��<����O>��?��9�
Mq��_ =��.�n$�J�)��ɢE�dV{�<������ə�I��O�<-ǺN���S�i���WdY�t�����M�g��L1D@@��H��F#���@n�^���m��#��e����9��0"��:
H'�K�t� X�� T�Lq��5:��4���;D���6�f�9\K�㧕s���tN{�3�w<;�dj�7E[����H��?�����9��Ba�)�ӞN1��LՒ���j�Ŀ�M�-3T	�"�B��T&~���;(=W~MӠ�=���7U�0�X�� õsxw�s�{��|(e45�1"��-�XJ��=ʶ���^u(c<a�q L�#o������[�|�#�D�q�LNN��a���:+!
��!L�vFF���/�ɾ�����M���S]�r�|�u�j�Z���>�	'	 =��j�63�d�.ꈌ��yK'���=���9]���;$㓓Lk#
D� �(�����(X�G4:}ꔼ���f�Ȃ�c����h�6	�U����V�Ԑ�Ge#HD[͍����MG�>S�ȟ�rA�X���:��D�$b�>u�ѻ�)E��F�:\6|�Պ�+�U:�=��khF�"M��o[���*?���@�.�*S5{ېW��ᩦ3oZ����v�Ӂږ<�ٯ�x^�y�{�6������)2,x�=��I,E'w�Z�97ix_ͧFh�#�W�f5�؟�F�8:ɻϜ���3��gL�:>��Y6�g/������'��U`� _A���F�r%9t�0���Q�RH�o0�U+�l~,bJ0_��Õ�l��� ��#~��/!��d��&�ʉ�O%�RSSE�<Z ���R��W�H���ȉ"}	 �!uM�L�W��X4�su�L��k+HN0�v�����[��K����n�F��|�:����ҡ��<e�Bm�f7�P<�������.:���E]�Z)I>���ա�7o��k����˦��]�6]N�r�o~c�6@�ejQ&^ ����(3�N�C����S'O���5���R�w}t���Y�LE�qǭ1�M�اt�Q*`��wl-ނ�݇2�u[�R��?O�7�?t�c��a��Kg�4�a�5�j٨��Ke���pl���D�L��@ �a������`��H�����ζ��GZ;ڥ.��x��tw#y� VJE�#G\���H��O"A'׳PD#�:%�D6 ���p�1�������pF��$�T0�)ܫc�ⶠ��wBz��K]S�\q�r���J�ptx8`��Z ���<߰�S�\�3=g%��4�͆�#��<_��HVFa�}54DO`�����x���w�n�S�N��m/I�dR���"
T�RG��Yn9�}������uȩ�Q�0lk��M���g���|� ����Cۦ祝.��̴nؤ����z���87:fu�t�_{�Vy�;�i��:�Z����G�0�aϝ�"Lۿ����3�^�iۭu�O��M�[s<�������ۧjZ���q���5r��1Ϊ�9e�M�4���ANS� ��.���#b�G��wx k8���8hj�k���P�9�r�؜e1D6Q�pol��{�$9 p~x6@�GұC#���!�rG���$�"�-���̠�M��H�4Sz�9���
�"�t�<Z ���tw!R2��$؀�`�m #�Ʉu�2c/�g!JtB��q��K����{X���ҷ��ݜ#�:~\�_��ɸe��==-l�ld�mcp����9�$�W8� I�5���:$PI��+;�gf�c��\բ[ȃ"3�?���Mrv�
�� ��������9����-�/�@��j�=1#j�pV"����&�ZT���i쐿o���o8�3��ͿW�ا�w���mo�řj���1o6fF�ʮ�\�F��	���7������q�11��a{~6mG,d�~��U���i�33���r ���lDVpM1��h��襨�i���L����l���Ƕ����\�Z����Ï>B
ت�k����J��.��O��r,�]q��M��#�{/�_!eHs �������D,�d�yJ�v, ��fd�h��Q�k�(���w4^b���bf.�\��J�0�Y"�&jߧO��S]�j@�H	Mq�G�2�k#-X,e�Li6r�Q+dDY1]lQ@��S��5�8{D�)I&��W#b�À:xq���$�qw��D��#_̯�4r������7\ô�U�u����~��W� ���Fʵr��1��c�՟�ׂ���{�]���n�~�WA�=WD�ֺ]j��O�z���Q���^]2��l�9��L9�l�
ƒJ�dN���y��r<Cy�<�+��fA�d�s���Y�>�'o�Lc�>K����;��3���CfϞ%�����5��=�W\�U�ʜ{�����t�8.�T�T�H����Y��"X�8���X ���(�yX���Ff�b-��B�E�R�0C��4��,��7j�X��Y|��j��[���X@�X�́,�1��v8�QWQ&$���1@g4s�Lƨ�� �e�R�&{j��g�^�;����S���g�P��v4��+6˭7���qP�{\�E�g�KP�{��6�`���� V�����.z{m,`Ow�����������s'&X�b�Z�<f�m���-��8���M�䑟?��r��W�Ow[]u8E�'�1s��ܔ�ƑAv�GQ`�{�J���>hZD��d�ʆH�ϑz�t�hjó���a�����H>R��q�m6�Z��=��}�k_��~���}�WL��;��/r��B0XR�D�
9��~W�P��o���I�2�܌���0���2���I�?����b��Ϋ���,bF�F̑ޞ�(����D�a�?˺C��F� �I�? ���w�ٍ�TqI S� ���
Ivb��l�s�,]_'!�8W{��TZ����`���G-0C���`q�F�(�"�F��&����q<����˯H�0��������\�����{cS=S�P���'k3�V-cs�����,;��f??ޣ6�^/+�j�Ѧ;�N�ۺ�t>zkv���Lu�ێ}#O�˒:q��h�V6�&U�Ow��Z ����,\(�/��3�j8lz
�ZZ\2�M��|����x��?���x�\��*F��:G�N�v�����q'ҖI�u����]\�={�ș޳���{hތ�#��K��gn�����?)O�,�q��� Im>���W�Z��x��G}�5����.���ff��Q�T��1y�ѧ��--{w�bV(�#�ck��W =���a����MB�MD� ֤.h�M�DQ�����$۪A�C=#G]L#�8շ�
 �@���/�u[�����j��(��?~�s���Mr���JE�r�Lǀis�0��n��c�ݭ�"SɆэ��@x���S�k�%s���j�5]n��8�֣�נaw��y�o����PgF����� �~N�js��D��?�O�eW���HG񖜡x�B#5�T���[S��WSѷ=ƨ�%ՒS)}F���8Ʀ�#>[�<��-���L����^u��޽W�|�tP"�u�*P��LyGj�	>�s�<Q�vdا�MRZ+��%���؆F:��H�Ա��9%���&���Y��"���sD��?��t�=� ��ٸ92&;��l�2t싼��l�J��n+�<'Ƈu_�i˺W���dͪ5�O�t�$%����r�ߜ�; z`32��mt�Mj��>%������)�H8&ǎ���zF���j)��u#*M+����|7�L1��}�$`#&��q����,l��X��1*�ܶ��I}�H�p	 �&��j�X#�aw�F�`%��Lj�/�T�d�!��N��ɩ�6��k���uމɱZ�7�q�h�)\�[�|&��`;$k)k�( e�������9�{��a��[��ULu��Kܧ<�H"Ƴ�~�N�E��$q.�가4�f�ׯ�E��ə���Q�	qR R�u8����r�#� ^8O�D���Ԯ���R�.������@����c�rX�y׮]ܯ�5�j� f�恟>D>!dG��<6�wS����J�B���`�
���&�wKʅ
����}� �����_���|���(A9ޯkX,�X ���4��*(zH��{�\-��.��K3m�y�fC�`��4��R����)T���dG.Z"Wn�*�����7�|��t�M��;rT>���J��DP���Mxp�/X�� T_�H� a2mt�q���,^�t�������Ia�gsҤ�A$>y�|w��]�ݴ��u�-�LT�i�3���F�辆�Aj�>����cA:ijl�Fc� f6�G�X�k�~�]����Uj�����5lR���sR���Lב�5ep�#­SP3��v�OP�h��2��!�t��r�7����Wޗ���E ��N4��:8xA^�����5�c�:�)J麔i�s��w8���~F�`)��>�Fm߾��1��wz�p������k�8O�#� Y��~�3��鹦eٲ�r��q�h�%rɦ�8��I7��R��{�F�Ey�{�+O?����mT�z��z`��@lF��R'+>4�͙�)�W.����ˢE(�(h8���}銥r�7�}�= ��=$�E("�뮿A��%9z⤬Z{�l߹��tц%7�R8�|��4�>��s�=��cm	�낌�-�o����NZ�6B����w�G�?�l�&S�c� Tv��!C� &�rv(h�B��$3��lm���}J��:14��5�`���\>��� �s����ݻ�G%@X.��2���ˍ��Lq�s�?�E]~���3ئ��jHhJ
֤��������ʎ�F�����v֜��v]�t��=���i[j��=����s䐲�H��}ý�h�qμ�����y ?�g�
��$�˂��4Rn��'�1�Z: �o�>���ޜ���ر.�(��oP^|�F�ǎw� � F]|G�Α:1P
#�T_Aڿި�G�Ƞ�_kK�r�f�jY�r���Lʬy��Y��g�����i.\���Me�^Ku]�T*��;� z`3��=�!������d����p�*}�"f�|1¸��tQ��[HOH��3~;L���	��7��eނE��?ʮy,�	t�W+����F,#ŋ�$
49!z�0̚5����C$�hB$��M�Y�B0����,]����!��+��+;�a�O��uf�,PV}B�W�M[bHfnٲE�4���!0�F��f;ǭ z�c��vף��}q"��jyx��~�q�߭|����h��'e���Վ���dHǫ�^8�p��#��3)eֿ=�n{�D���:��m/���H&�Se;;oޭV(�b�ma��?�פ���կ~U������O��x�t����:��dW�·���e���Y,Z,���_�f��؋�xC=QP'W���H5=l�Qn{�;d�%�('�♚��!��I�B3s�Β����F�d�>��U��ĉ�)�j˯X�L2uxvK�v�- ��fd���M����~��h��U��[��3�jo�d�|hdT�.[!��-���)7�p�<��S���П9�+<�����K�N7Ȏ]��n{��y,����KϪ�Ar�L}����9G��MN ��"��h�Fw��DZ(�K.����裿`ǵG��#IDr�)��2�'���g�Q| �I��)����=zT.��i�T:Ip4s�.	KzN tS�'���x�l&aFƹb�ǟ�Gk ���������ݝ2�����`K$�&@����tV8;����9��<����^������7�KˆQ��Ϡv���?��4��Ș:j!̅�Mͽ��b8<.��:�3a�>::&����E�vu
�ώ�4� �����t�Ѧ�Q:v܏#jHS���R��ԣ�7����<fu,"ndm ����+8iL�'�`O,���-0�E��>�=$�ioi5Y	�.��T�Ӏ���V��A`���@lF� P)�.�q��Q?�sd���*��HTi�"�w�za�\8҄���S�^^{�Q���t�Q���/]��3��s�ɀFg�J�E����,�UE�|�h_<r��ޓ���V0��L�c��olf�`iol�X]Cc�`���!�huwf�}�x�jv����ǌ=z��|/��jqgz{��G~.��.�(LT�$�.�|����n�i-}�w�8Vb#�CZ���v�8��^/P���l����V�̰�95���{U���O�b� 5�ˤ?��$-8.4Õ*�.�t�l�ݣC��ܤ�^[���B���u�<��I�җ�ĬK8��:'���� �h�9z,�be�B���a��T��y��
�!��#���O�����4z!:�P��r�ӑ���lt��f��68Q�̀sr���́x��p���~���gz����r�80Ep#8���f��NHG�,��3tx�N)�&x_._)^I��B)���C%T�V��z`��@lF�p�&��3 y��aA]�t�FJ��ؐe�Z)����]��*���M�n5��?������� r��-����QX������9qJ��$]�Փ���j�e4�Mcݏ�T���t8�}V�"�88!�� ¶n�.lvpK�6o�O��ͦ7',-�1d$:a�pL����1:�{� ������AQZ��@�:]4�z^ ѩ�T	�8n��Hd��T��L��̠O��ٚ8J�j��?�p{�n��q���]S�/W-�l�_ތ�!c @p��B�p=���r���G��ڥ�&B��Ma���U��;��3��E`� k�8�l�9.eg̍ӑL�`�l��X\��A�/�9z�	���>{�~��]�0�0`T2�ڸ�օK��u�]'��w�4���^�\n�p�$��_ٶ��T(��K7_��{?�>�Of�n�[�^+.�K�q�N�K&�pزz�y	,��h�6#â�А��4������9�۷o���3���{wm��QFg`QC�q��Er���u��y�oQ���'���|JA��QnXLW2c��� ���P��:@?�pL���"�N�|���T�%��C����( ��a��s����d{ӹ�Q9i��������}�s��ё!���7P/�!S/�z���m:��`�mz;g^��l��q��(@Y�s�֧j���n�pdJ}mz��j�}�����&|����9]���8q9���L���ҋ/+X��]�H�3�az��[ء,*�5������{��H&?�{ȕHL��F��(A�f��AD��9����E��p<b1�'��K�L�d�]�p�1��A}}����;�#;w�$MKc��O�2�����#24xV�]�Q�;�����ʬ�=�^PT�nm�%�C#�2��#Ǐt�+/o�����E��̚5+ ��Ϋ�،,�;������߳�]{��e˖��d߾L�R�CM��Iu��#�������� H��Z�J~��?��|H�;*w�+��}F�O��x]*����ڪ��k�:h��Q�:I (�ʒ�� �E��Ns��)w� �����8������6G�2a�:��(�*|�H�[�T���냅�ۼ�k_����r����0�T�q3D�與sA�.�k�L�Ƽ�����_8G�l�}J�|:�@�2�M'���vְW;��p:�B��P����ϙ˿!��+N	�� U���o?Cd�1�|���k�S�QX���m��S�MXډ�����^�:XdAP+GT�U�J�<&&&�TƓ��M�t���������>�%K�pt.71���sTK&S|�~��{���6Ҩ��u�>�2�s�dꥭ����Ւ+������G���棛6m�Wgz�%��΃�،l͚���u�~y⡮744ևuݵs��PPG����l����f�QA}�K/�7�����K2:Z���v΃#E���]w}�MK'O�d��s�v9r�L���9���hC���љd� z��
Rf�����D$-y���-f��x��H������r�ixx���x"�}`�'�jmX�K��L���	ՀRd�k�W*�\#��a��Jfj��%֫�l8��(\3������Ʒ��uЮ{�Tj-�^�I���;�:�Z�ݝb]�����Q-��	�K��ڲM��I,�โ�ݔ L����#�>� ����FTgHn|�v��@����SR�G�(8��ut���ߐUI���2Ci}�6n�H����>X��T�b~Xr���,B!D�h�;p�����;٣o �e�ʉǍ޻����3��9 ]��2}ԏ�%�\"M-m<7�����+_�����>
�3�f��ٲ��$��γ�،Qƃ>�����;�⪺L�yYS,�K/�����$)`A�o�>y���_>��rJ���������.��'?)�4*Z�b�,_�Bn��z�^x����Iʂ�(���!g15UCˊ�6K��Q��&"L�Q���¡*�h������5kY�Mh䅮�ɬFkn��OS%G-���T����:����� �]2���l.��L�|�S˹�������o��!�A_�Md�2���U�	K\&�*�R��h��t�2�o�Ng��/�Zc^�@n��	���)��F8&jQ�H͉�Ӂf��h�.(S�0}Pq�	2��s�=�Mի���S�j2aF]�j������#�[>�ֶ6"���t��}�[JAcu��A��Li��pM��*	v�eӑ�Ϡ!���<������K1���Nt��~��~� �Q�ס��i�n�7g�<��S�h�"f������!�ՙ�3w�w���2o���;� z`3�[n������?���?�D�P���sh����}򔴷w�R]�A���Ȉ�4�"��76�"�Htp�6ٶ��E�@ #7>�E�f0�\��J*��HYţ�&�C�T��qtbPRuW�g�K9��+ ��)@546QU,���UA�Mc�#R���㧍��_�
�0�aH3*����uQ�sk[�46���
�7v����Ѳ��Z�@3j���㧍*�XƢ�×UJ��,����Kv��;[����&N��H>u�^�Yw�������#��g��D�quB�� �e8MQ����r/���9��`<6�ȯ�GC�ַ���Fz������Ty ϑ���X�>S?��O���g�1��bp#8$���"�N��G��zN�Ž��ȟ|�stB,l�ft�i�����
�MwO��y�O�����#R���Y�m�g��~�������&%���, ��fl��u��.ң?����T��K��a����4�!��ʕH���*
�j�Q�m+W]�����nuu���,��&5�uˬ�"B-�\�˞��)})���)b�����R�3�X�Ou�&�p����(�:�t)R�3��E��[)R�O��K��e�F1�p����k���~�\Ʃ��M� Uv|+xP�w�{ $��O{>�����i�sצ�aI\㹾���;��n����j��m�lg;�JV�Lq	}O�Qv�á��u|4��c�F84�y^I|��i�f3�a�d@F=��c:r��>��8�b΍D���\�~��c�2�u^Y��;�Ig<{&N��=��d>���F�q�6�:NU}��T^�;���v���y�l���x<��E/��wtt���475a���hS>
��Rɑё�lGG{O�.�}饛��~�[_�{?$���d�v^Lޒ.�v��z������?~�]�(h����cq$��
�!��:�������A�~;_`�8YL�1�vn��>��Q�=C�j�H�j��`[�jQ����g�ay���Z[����3�w�́�j���a�T�9�5!-ǧx���[�Ƕ9���Wya���?���<����M��(͋�C����]]]����)p�1c� ǆj�� 4� }����~7�a~
�zn��t��6�ՄT¦l`f�C��z[s�����3�W�� ���ԯ86��ʣn�F4h����U���w/\�hG8� Y��J�JAtB#�I���!��!�*��H��.�{���P��P�sL������̏^�j4�`�>9ǭ��7�V]���\��ש�/��.����B�1�#�w�S �,��;�JU�W��Y��W���¥�>�au��b�\i�F���6����C�|�	�D]}�1�X��x����g��u��*��c�	,��L =��f~��]�?��o|�k����������D�p��l_G.���N$	�C�H#6ԥ���)�;�k]�]lO�h�O@��!1Dzۉ����,	���uĩF$�E4���w4BX����ׅ
U��x�^��1W�
�x*�wl�Ճ��U���rK���w*�P%R�}T*јƈn(��ʕ��g�Rz6����D��.[�d�����*�X�钦 �D�-[A�F#�ʕ�Ys�g�����_��_5#�j�Ws�B��ӿ��.s�B�Ǵa�E�,�*t(��9,���X��{���o~ӟm��g��e��8N@�X`����y7�_5��<�C{�F���ϕJG�F���6V�t;�?6\��*u0hm@�;&ǎ�h(Qc���ӈ��˧�>����7��G��~��U�U�"Nm;�!c|�p��X�0�!�R������J��|�.��L��X`����kf��-͉EB���xn��X%o���Q��}sk��i{F�l||��G]�����'�P�&Qf3�&�ȜLm~ӝ�ȫ�.8�t|q��b0H�C�c]8�x:E�4R������`X`���X`���&'+Ԏ/M3�?������G@�i�CC5��4�f4.�+�j����I�[v������v�R�Nզ��H�X��gz�a��������P*��8$/K ��_b��kk�e�)��L�M�����cP��/�O�dR������CW��bӚ�~]=]���W:�CFqmz�}:#~�1 "��D"��d&!n(�NyL4�r9���5����� ��5��d�T\�V��H�.�!P�9jC�B�hHZ3F��R�Mgεy�r���W7���Qξo#u2�Y�ڪ%�)���`������ݶ�K͗�}�<}��<�t�q�5��{�- ��{����cc׏������;�hLfϝKu/�|A�԰�����z]C��Y�e��E��hH��}�Z�}��	Հؒ���s�U�]�a���	����8�,:�������S0�e�2�^x�#u��O��w�gsX`��f z`��F6�wf˱c�>s������-r��K��N��,��8�����N���X��S�H|���f9+"bA�Ε�q�)��W+�Y�ߦ)�ըk���-�ۨ���'�;`�C�>�dÑp�X��[�������}��7@:$��kb��kd���{�F����6]��K�7B>.�Qw�s����l ��E	�I��n͂m,���4жLu5~w�;yլ���W{u��i�|��m�� �棤y����r��ɑ��^s�X.����,_��^70��kd��kd�憇�\��7�4�Z���������"�����l6[� � ��R��Q�����b`�5������5�1ּiҰ���Ύ�Y	U�U�������ں�;;�_V��K�}��o<�_�m$��{�, ��{����}R��Gbh���8�P�
ʍ����>}z�c��{k*��(x�5:&%����Yـ�U�ZŬ[4�N(�:���z=��7d�u9��\�L?W��Q��/8�Nccc^��1 |^�6��S@�ONN�؎͞={��cE�t����X`����:���	}�U�<��������H(`F����� �|�cBg���g�LU�_#iVm�=��g��~��W�n����`X`�}- ���o`>��Q��X`��_Z �X`��:� �,���u`�X`����@,��,�ׁ�X`�X`� =��,��^ z`�X`��, ��,��{X �X`��:� �,���u`�X`����@,��,�ׁ����W2    �����D 0 t :  � B�����`@� 0 t :  � B�����`@� 0 t :  � B�����`@� 0 t :  � B�����`@� 0 t {uUcrC%%    IEND�B`�PK
     mdZ�S��*  �*  /   images/cbf7ad0e-0f08-44f8-98a9-dcbe92af212f.png�PNG

   IHDR   d   d   p�T   	pHYs  �  ��+  *�IDATx��}	���WU}�=��9��HIH ƀ0�`X�������6���x^k��lq��`#N	�����4�h4�}�t�}�]��W��}�"^���Y-I4��]U����/��?�/>�y%*d�ɇ
�g�B�|��y&*d�ɼQȃ��$ɀL6#%�d*%	�"#��@��,�,�K�e2q�B��	��+��l6����@/#dzo4)Ch^ׂ+7l�|�y��'�=	��8�v'���42<�$&����D����fYK�I�0�l�D�?/ɚr:��:W���bP �d����{{���I�B**+�lU3އɰ� �)g4�Y3*)C�x�C�Ȋ$�U����J"e�#+J����YVT�٬��T��h�Y>H���\.�'�7
I�∄��EbגB62�,W�H:0����,Yrpk�Y��)F���s�ZX�`���}�
aV��<�J�0�d�(� �$h�3j
U4[�.���I���2t�Q(���s��T*Kߥ�;�P�v=}��BU�-UMe�'��4����lN$�4l��m44�p��9�N�������Y��l�>�$0��e��L�I�B�n��5�`+�)O���y��Y�pͅk�s�*� %���s��y�����$c>ɼQc}0�I�ɬE��,�"I�Y�!Y���D"!�a4�D���QUF�O������ ���^YI�|�y��_蘒����z��s�_Ba��C���Bd�����>#��j�)R�5Lz����ItWȳ�=�Á��!D�i��SD)�ww!�;J�=&i��0T�'D	ˠc����lk�� �b�T�N���'>�����`JnwN3��W��p;F�Kp�m��K�ǻo�����i�-�*�_���:�<gO�v�����sh�<�[Tկ�֭���x	�AF*�FZ�Y4�xǃ����0%|EP��]�&8Z��T�Y�p��N\RS��^�,f2��Ukq �A�>����Euu��c>}��z��
�XX���M���S���n�\X�~��+�\q�1��`���`����Գ�CI���r�C�����M~�������,�V��X���sp���^q�Շ���G�����wg����w��p<��������|�n�m#�*����	����U���>fYPӀg_x�&+�$ʊ�q����ƃ}�h�o`*�B�Yi��T��T:%>���l��S�
�-�/��ccî�҂��,k05>�5��lQ<>O�3������z��
	G��;ή�兗���=#��2��I���cA��I$�Q5A���V���U��"��!�cF�-ј����"�;�����cIS"4	�D�8|�~�������C���:�K��誐H\��V��w�K�N�'�PѰp	�v',d% ���VL����'q�qAͱ�C��VF.��L$��Xa��&���$�F�VÖ�ν�Ѕ�X����1�")���W��`�ؤ��� ��Ǡ���I�Y�A~�[.Eg� |3A�-H'b���$��.C���pm&���
��'�}DXGV@:��.��Y��gggdVE����LN���%��� 	���ͨ���[�?�J��T"�EW���aLO�`���X��2�W�a��V4-^��gN�Y_UQ�q_R���1l�(�� ^ӈ�b�����s_ɭ��5��ј�R����BJ�+�7<-��<��d�K�6�7�o ���#�矠�誐L� ��\mkkW'=����H�+��P2�F 5��X��9���am(���_���~ψ�fQ������.+b�\Ϳ�g00؇� �v~�SS��{�<�c~P�z��
q�������K���	��
���6��*Q^^��������l�e�K�3���[���N�?�F"��7��511t� �x\X+���Ʊ����Lk+]c�o"���'�xI���Ϡ���C2bq��Љ�n���0�������qb�cP�>���H�g4�B�gV�z�`���m.�+`-��,V�S@0���\�����L {��0�P�a���_G~d��_������-&��7����.]��)r�	r�L��E�4`
J+�16�!v\���LJ4[�X�%�H$���A�����ő��Y���9{EXE2��{a��E~������3��3t-'1S��r���U�%BY�L��
I�Ė����z�\RY����ӭ`4���]	�UX'�Caa����C�EE�!h��lb�/d{�gccc�3�+f�Y��f�2�����B:;;0�ϐ����~�xP?���X�6�.F+�P���ߠ��\T(�1����0g�L��AqY).l�)��t@���ⵑ(sVL�|+�-'���S'XJR�J�{�ɺ8���Ҙ�0��s�s��ش����#�a�?�B��PE���G?��}�LN�E����o�;��C�~,^�
}�=�������J�j��+`�!�_s��QgA��U����Aq;s�m��PyNY��Z��z��rhp�a$�-7l!�~7n����ص{o���փAo�U!6�j�"+F�"9q]�=4�V�-�F�@?�.�1�C0��$v�1Is!��`e��2X�X����s�:��}��4?����5
O��,6L�M ���`�ӹCO�U!�e�p��#�ۤ��;�v�����K����^*�¹D���2+C�eW��VCn�	b���`1�g���gr��{0\Y,��0�Mz&��J��T9t�,׃m/�Wށ͑7�G���������C�s�ݤ�b4ȱhP�(+�YA�f$GK�ee(�(�!AȖ��I��ҙ��Fn�Z�&��l�Ă.ʄ������(RN�,DXJ2!����٬�jl6;
���~�K��/v�PS]�@0�*+p��׿"EW��;�[�r	����㥗_���A�/\���L���؞��CXN$r�9A
���b̕�h�o+O�PWs��c�\F�_lA�VT^���>��7$2�`���8{l�\}.��#8�v˖-#�6�EW�Ȋ�gh��_}~�����-������D�&`��')2b2h%���H[��Ա3�c�"�.�)-����/������Ur�w�g��r�X�r���?^>vR:�֍U�k��誐��H�������3��L�7���wv�UP�a}��*�#/����<����r
%�+�s�Ba��ȅZߴ��ʐ/�.�qJE���;�E		���m��N�d�㍷�b����S'�E��[�e��ѐ��3������&�0�lg"�G�΢�4Fb�F���^���%������+��U^^.����+� .b�<dE����I�y1W��X�T�����3�ԗn�ӦE��
aX����*��O�=^m7>8r��k���%����HZBFղ�i^���`�m������ʂ8T�����H9x+��O��\���`�F�18�O�t3���PWW�k>q,��*�z���?�	�]28Lxm���z㞩��>������q@�����P^�΃j�Z4�d2� � �3�|�bQs�sk ��@���f2��H�S��=������]o�Bxfm��1>�G��h�Ǯ�M���zq'c���ci_�YQ�@
��3�|���%pY
E�GEe�R�\>*W� 2���[��K�dr��?� �8(�e���e6sQv�7al*��a�ۦirRH�g�S��ȣ��k��V�,�1��.�)��t�'��?���@Ii"� F�F�S#�k\*P���N$)2^XdB��D��J��a.dH��bk&��VH0�����bQC��3m��!�E��z�-ho;��k�㲍��܋;����;�Խ[�%\��3�3Jmm�ܲ�k[6�d['�+��CeE
��������w۶aÆ��k.�� �(�f��	YIKHr֖��CZ����D9?�Z�X�b%+yx�Oo L�[e:���i����(v�Swf�o�=������y�Oy���)"���)1serУ�d!��~��,4�=�I-_��!JG��
V����33WI�N�>���Ĵ�Zv�lNli�\����)�B?	�c0(f���O��S��}��o{V��ޢ�B�����d���	'n���y�
Jʱj�:T���	fDI9��}��"e�Yܹ�h9�Y%��ҙ\բ�s��֬���d0jۼ��S�e��wq)Y�g*�Ν{0�ۍ)�!.�Ѡ�|�G�f�^�-�9d#�����k��/߃w�݋��D�%K��� k��ġ��tٕpXͨ�����ag�"�V��WA��G�q6�W!�b��&@�&�F1��t��1���_(�1�_�	=�ڰn�������J�����n�z��
a���A��H8�<b�<�Ņ��񡴢c.?ފw��K3�N�Z�Q�
kQ�(Z���ɞ$KR�l\N�V��'` ��V6����E��'֭���W��m�8|�0.^�H4%5-�(���[tU���D]m�z������-JK���L�<**`t܃���	�W���7�Z���E�n,$��[�V��0k�����:�k?�eK������l�&��jCS�%8q�V�\�}b;��|�\��uu��&�~c'YU
�z���a������v�0�]�L�s��Y�AV�N+)$#�δϋ��Jb��f��7����,����sx)
��h!E�g�A�Zڻ&����C�4�GØ�	axz/)/��=^
���o�lv���[�߂��b"�c���y�Ld滍���c#����#��&���ܰ�@?��������q�\���2�Z��|f�O�1&�����s\^�(��u"��&�s�k�RS��U�c&r���)�2�hi`Hcc��qa���;�^��-��7>��n��V;|��z/���g����ن��
��Rϴ��4EY\�`�dGlu;i���'���h�[�� *f�H!��ϩEc�4K<�Q*}����"�"������ٳV�O��=� J˪���&�Z�ZJ�/�*N�-�.Ϟ>yJ}����A���^y�T�]�إems���s�k��$�!用j�(#��l�|-��w�X���G�SbFQQ!��+�p���*���{�"II��_ǒk�5k[$N��-�FY4C}�I5�mWW�]�ށ�
�
��bT��D,��K� ��v�koΕ_��(f���S�YY�b�<��DB����B�6��R���,�z{PXP�(�F��S,(t������ÁCm��ýRC�E��L�044����R��NDbi��_`Ś58t`���ZP]E��b�X��kڪ,Jzĺ����dr]��Ė�"N�g��O'㈑��-f�"ڟ�U�f �SK�,'h*�����Q\�������j�ͪ��?I����ޢ�B$��5����!����'��,1��' ��;08<B0f��bCm������H��K��}V�u؊�Cz��3�3����ӗ��X(z+*v�h�t�pf����y_	�F�s��3��[n��	z��Q��Ƞ+��e_}����HS��Eό���EQVY�<��(W>��]my��/�n���oa��{�0��V���������JI�.��e"�I�D �px��]"�M>\��!�`d,������n����Y���Xo�ׇ�����%�y�m��g)��:߃�j�=y���(*-C��U(��k�1Q��lq#��v��FSm%�6+<�#G��514�DB�j�����p�c��$.�Pa&�&���k�Dج�ϊ��M���-8s�����z�V����WwHK7@o�U!	��C�j]ݥ��ի�|�|��?��] ��ru����}9�������$X�U�2�]���uxg�[I��>.�&��B�]�E���"��;;��\*��8Q�#�J��{_4�VV�c�@��+ω��>�'y�D��Z�z���;���?&��X������c1�N��o�q����!�>Wp��]m����)Z
��)ֲ��^�#ַ�D˺��U���������"��z� ����0��/�����Z{ǹ3���I��O ��k�����Š��ˢA�s;T�ק�Rh0Y��!�Ոĺ-���х��6[P�e�U��>L�"0���wZ�5�/H$�p:�[n�
�k��sQD|WLT�4-Y��L�ߎ"�I�}|��MAN4�$kQ4�O��r&���4�.�ҫ��Oi��P��.��#��څ�pd�^��3�$*�ax�BX��P�'��������[a2�p��Y<���zյ�tU�oe�@������@Y���f�H,Kpv�ͷ�p���^E�4������Cx�w�<�o�������bH�X�Tc:�2� ��T#�M���H�&� ���եy�&�vY�=A�`�y�sW��*��A���VBza� �B1���N���>+������v��P�oބ��a�,�艏GBŹ�!�Ҭ���uR͂j�-�󐆦z��|?����D9g:#���v F�"2�ĬO=�ȴ��Z��
�za9�f�h0;�sG7���㉨h -/�j�Y�;r�(�sb����N65aղE�A7[�q��8t���z<���ff�������+���6���S�[��!4��ĺC~���� d&"lFQ&�
��<��O�D~!3>���I��\�����a$�x��a�{?fg���I�Ϋ����E,_�\� ݟ�MRt������qW.@�+���&��'�A����^�b�1<�GOO��Z����c�`� .�R��0Y���_�F�]T���TޤQZ�B��������1���P�[\R��#G��n[6,V�ݙ��l��;�"*M81�ʦ�Ŵ="*��� �܎�*%\��z�ƆQSjŵ�n�ٶ���G��y%���Գ�/�W=Sb0���"�`s�5�F3���҅�p:���m���L���0F~�<>��%豹�f�Mљ�"�]XB>AFO�y�aŖcu�(���T�W�(���E
��֣d!�Q�^��J�5��b��-�l���4?{��-��_?%��7�X��pth�c�)�M�"p��c�����@�߇rʳS>
��t?��7���&����gd��,V�l��K%�()-���^'gE���� m�^�*��+]������e��eJ,�.���@e$����y���0C��׏k?~#���S�MzE%�������Ս�q�XPP�鄑�f��K�!��2�nb�I��s�.�u ��@
�6�ESi-m�����{���ʐ �rin��M8z���ct�z��
i^^��������>�F�����_R"v��%Y�ق��2�T�#��)DFg�{av�!����C��s�<�r���eee��skCw� 9�$��JK�yJ��s����ˤ133�[n��:!G�PRԀ�U���;X��	z��]�&�˖�O���_|�E��`�lU3IX�_��S�Lx��xQ1ƆzE����a�K��;�q�>�İe1�M�m6}g%��b��ň���o=��e=Y�⥍��酛,����#��ލ��?+�j�����?�=�R~^��AoѹrQ!Rl|c��{?��H&��c������D-)J>C���clM��v&�2 �@L4��j`�;Ol
�~��������|�X�5MX��������z	�����)��B$'&F���<���&g��WRb�FgїJY�!��|�|�g��$s��u8`!��H���
ь]C��]�Qb�ee��s �>��x���O�[��d%f����Lb�#���s�OV[VE))����E��L$���gPV݈�`������؀����<��-, ��[tUW�3����H�ml!��©��(,-�e���Y�;.���b�S��������0=�\O7�t	�8r_!�"	��,�g�߲9�(�iD$���(��
x�Xl�������v9ɏL!U�%(�d6�IE�@wѽغ�� =�ko�����j�K����ZAs��5S'�AeY���2a��9�Q��*�ML�.*���h�<�@P�%h& 2��He�h^��+���&DW���kP^Q���ދ��>�uww��+)�s�>C���d�׈�
	�m��d%G[O�Z�G䣵�����}H8��b�N�1Idp��UB�e�(�Y��q���!���p5J�L������0���4�r8�P��$��-,)�bAV�"�9fHF�_��������]�qn ��PLV��#�Ȑ�*x���q͍�»o����d2�����ɒ���R4-]�������F����t���L��]z��Ѱx	�.AQq9�ɲ��Ӕ��a��{��q�q�팀Ы�������C~'���'����z��
��#�H'�R�D�Z��f���Ǥ�z��:-c��C�ɡ��;�׃��j,ij@w�X�����ɓ��n]�8^��2�mk,<8;����s�g��Cl��w܁��^d���j��ڍ$L��op#���^�()5iR/��$��J
2�:ڲ�k۳"�$���ϋRN�x�GS�	L�n�C>�OlL3C���!��7R ��1FS�)���TTV�v���X��NؒLf+)�����E�����w���Ь����5������}��ܡ(4��,�儢IѺ�=$-*��`ݪe�����A1Y�a�2�M����4pє�ID�4D��EY���xR�_�w����.]��6]*��"���3�� ��Q
m�zZ,!��7�u��0>r�����3=�u
�E�M0���<���b�k_���b|��G÷�wvR$4 ���z��h�G��K/!�RaLGQ� X#�w��-8��&��1T���p����=�Fi�캵�4�!G=�yY���]m]-��b3BD����P�h9��]&�u�V�����#r}C��ۢ�-F5��}���;&Db�"*�ɽ��MX�t�	��B�o܄�1�)4�?�w���n�/��&�m{_��]h;�&�	��ƆKp��	�����wcjj�y����i
����!@��C�O��8|�R��3?8<�]���]grZ��^��!�T�[����Y<A>��_��|�۳KXΕWl�G?�]���V�o��;^����0���Ά�~�J��a?��������:o*S��]�TU� ����12�CP(��a�pۭ8r�0�,������}x���E3����~�,E`�R}�%2G�-:W�H�g	�����b6�U�MK	�:��F轃|	��(Y��#	���_w�Up�c��}�!���$[T���Ξŕ�ՕU0Hx㭷p�L;zz�(���n��F 3q��,|o}��y(�"e����;����h=u^r��[���x��!�غ�����Y�u�})���I"t!:�L(-viU$̘���:D�j��f���p�R�	�<���OR�v

�=��S�3�"!is$`(7
�i�F�,2YZ�*��r㺏~�v�Oљ	z��Q�B�Vái�����$9v7ʫK�.r����]��6�.��Z-.�`尲�n'zη�F���sD?1��{<��r�=�Jlq�	��&e~�W,P��Ef
��k�k����J�t�"/��MJ]n�L�_������)%�9u��S\�XT����G��GB�bwn7 9�˖���b�f9祤�vV�UN۝�s#����D"���U���ʒrr���W~�h���G���	�lR0� z�8��"���V�F.������a7����b�~8x\_(zC��4���2Q�;a£�
&�_���]	z:�	�|(+)��\x���LL���XpMϣ{`L�{=z���Z��?�5�r��U+��
��e��7�wI�=��\T�ޢoE2�]���6��?}�0Z\��u�31���^:z_����=���w���#2�q
m�;���e���x�����s�k��+�����W^���E����������5�c�uå����P��gX��l�`��&�,�X�b��>�4[/r��6,h��?8|~���~#���$a���e��L�11�%˘��$���J#�D�^y7l�^�i���IB�[�9O�	[l@<���ᳳ�t"������Y=êb0������	�ӥ��,������Yu{fz6�N����Ɔ��[tU�wr�f���"o��?5Ks���:�u;R^A!F'<���1��J5�,��BcZ�����i������_���l��;� r[s{h���/�����nj�l��_�}���P�%��$�ɧ^��u��3j�T�ɬ:x K֛M�����یw�~Gl%��誐{�r���o��{�L�r����h){�d3�Q���C�wj: Be��j���פ���X_/� x�xl��\PQ��}꼟/��V�%��Ǿ;�܋/Sx�x5*Ii�����l�5�b�zIDEwomen���oJ��Cc��W�"}rח�(����޽S'����~��_�O>�\w�w�TY�M&N�KiY��V�*?�S<�-�t������{�݊�Kq�UW�?���]v��#����IJ�u+)C���Z��#�dI�?knc3��ͳ���9��]��(�+���/���.�B�|��y&*d�ɇ
�g�B�|��y&�(��5�N�    IEND�B`�PK
     mdZF�i~�  �  /   images/85e66502-362d-4a26-afcd-97fbc4859675.png�PNG

   IHDR  �  �   �lC   sRGB ���    IDATx^�y�o�U߹�������$��$YÓml����ӡCU�ؖ��bl�iL7Ch��!@H��ҡ����Օ�*����ƃl��,����7�������]l� ���٪�{~g�:{��k�9^�   @ h0���m�i�   @ p^� �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   <TU��tYE����^��}�w!�   @��J�����s�Ҵ�1˒��䞝��_�t)��(���EQ��8veY�eEeU��M��$��yQ����CKK��6�%?�}���v?����|���   �<����}�K���f?�mw����˭V+���]�v��p�i��s��%x%|��4s���E���(��^��q����o<}�ռ����o��+� �W 2@ ��_��[���r��p4��<��N�'q�z�~�eY����n\u���E��(rE��5�k��*��*w.*�8n��[U�$���<�'���Ao����>�W��}K�����K@ �  p@���_�-��o�Uu�sѠ(�YQT�4I�0��W9�+W����]7����v�-�y�$�Ue����$)�$��0.�"^XXpG�������?�.��	 x�|F��   |I��_�g4�LQV��Ey�fi⽲R���\�f��v{.��������q���E��o�����)�Aq�ī������������ر����7��!��K@�b!�   @�/H����O�]W��8]��&ij�Zye�[bZ�\�W1���ή��]9WV�%����%ᬟ��z)���j�+��?�}��C?F5�_Є�s@ �  �	������sQ�3�V۵���b_yA"�G+D
Sp*<�BcUY���=7�\QN��*�g�6x|��g���������������/��g�   <�~�g��ue���v'U%	^��Z)^	� �+W���Gn�?t���%��*��ƉD���UY������i������O,-.��7��۞zN��8!/����! @ x�D�ϟO666������8_�Y��>���O�x>��\��\��-�4���]�WB$�$b%x�vw]�Ԥ�]Y.IcWv�ݨ�q��eY�i��ǎ͏�-��Mo���=g4^�F��;�ۇ   @�Y#���oM��]�g�������J++�[�9�F�ϟW2��t:�{����?�c���'��:�v��z�8��,��r����4sY��7��w��ļ�u�1_���t+��^��Kb7����Ve�����r��v�E�o�c���]�۰�9�   |�Ο?��Z{�E�B�f��|���v#�W�|>���N9���۝͕7r������,͞|������yy��j�ť�:q������ͦ���c��N�m7�繉_��*�-ސ�vX�:M�s�,M��`��xÉ���~�~G�~��@ �@���mok/,LW�i��ҕ���������#��d�L糹sլ��~`^Y[;�@��w�4��iֺt���.J�?�y~c�j�+++i\{x}H��\
e������W�{������!
m�	l���u]�!xzu�.S�n�[�r�/z���G�-�Zs��J.@ �������[�&Y�����;����,�LƓ��S7�F�ao6����Y�n��w���7�tz+��kUU]lg�Ս͍WW.:[�r��vkG����g�4�{+�Z�+��=�ԓ&�����t:���N�c���^>�k�@b�9�����۝��go>��7��/T���}� ��wv�KY�2n�Y̋WN���E�����^\\\*�����gY�&�I����\�����x4�~o�$�t�8�tUV����v��\�ӽ<dۛ�������!��u'p}@ � ��D��ߛ-�^tn<y�x<���h��py\��W]���p4����|��4s�O����;n<�Q�$�����y��Y֊WVV�����ʻ;�͝�f��Ӂ���=��&t�VW��+W���UkPȮޗ�������u4q"�����G��P���O�'O�x���w��k_�ڃ��4���~A^��q{����׍��o~�'��������f����jd|
ש%���-t�uUI��p��I�<����ʭ�rqi!�J�,�r0X�vB��v�p4,v:��u��^w���t��j}���>2��W�vze>ɟ^YY}2I��<o���gS���������@l^�   <	�{�ə���O�:�����[���O�E���4����b����իW-�LUN�V��&әtC)�!�mY�q�jۿWWVܑ��\UQ
AHL���g��w���-,�x<v�V�b|���v:9P$    IDAT� �,�G*[潻����W�D��=s��ͭ�������*yra���ӹZ���v��x�b�WY�<o���'d}<��{�wskkmoo��Ҭ5���Z�&I�U�p8r�N'�9�Y+�]�rcGiQ�&���[\Z,u\_�ݎ�����ڪ���,��,���1#�Q����m�M���T��f��oQ�J������l:�������M/}�ՙ^+++&���tʅ�������Ǐ�g��~���=L[�F����WVv���S��������r��v���ne����Y��?��y>LӢ�nz�����"�����S8o_�`?`n	� �{�ϟ�wv�3���;z�h�e�c�?�x��z$����M�3w��I��[ZZr�/_��]��������q)A<s�<�.q�O��y�&TC��Y�0w�.^t[��nqa�zݎ˲�'��J^e�� �l�
˵+.�Jl�����dmm��G�9��N����s�X���Ӂ^���t �4�İ~oν$.uh�����H�n��EY�Y[}j>�(�>��葅�ړ�Ї�/�����|珟�p��?�r��=�����MA�k;�'�ټ����Ι�i�R�v�]�}�����6�����b)����d:���=7��}��JFVJܪn�l>7a[�2&��d�Y�SQ��N�k���iZ������knuu�mnn�����j����ZeY��.�:u*�Wݓ<�Z�i����c���h����`�O&�X'&��p�ot�`�߳�$z��,�*.}���z d�>�=.{ݞ	q�S�Ntɋܼκv��c݋^�^�T����^Y�f��dF������q��[��tsyiy���+I�&i�'}˹h���o��t#���V+ݟN'�s��R�jR��EQ,�ǎ�>��.T���է?��ꮻ�:��x�y-������'@ �+I���#�N���J����`�8����v'��/ݰ�?t+�+��j��d	��dj�Q�P�C�+W����b)���[_d����|,׬�E+K����{衇,�aia�v��CJ�0��z���Xh��Z����y>��������[��x��)�,��y�/�()#W�
�H�Ԏ;�.�.��\�Ib�9˲T�7L�����uUmggǴױcG.�v�m����~�o��7>o�x^^�����t��zW����p����mi�eY��u�ťXbLVb͋��)�a�H�*�@B�o��ޣՏ��p�9��� ��ܒ�˵u�؛/������$�f���î���rww�l�[n>�cms�b�����>[;��������ŋ�3E��F�$A<�ڶ�|��m����4-�BטO�q�nǭV�&�=h��4I��`�����d<��ՙ�E)�E��_���q^�Y^j=���3l��������ի� ��q�^��N�]����:�{0��u�45�����X���E��w�� b���G���&��/�L�3�3����ask�?v,�\�u_�~�V¹:3�S}?�ά����5�8P�&q,���VҠ"Q����'��L���8��ι�(�v�4fY�RG��h��neq_���v%{eYΒ���&�YUӪ��ը*�$)��h�P��~�·��jg�_--mU�����_�����B�! <D��{o����Ϝ>��˗�������z����z��:�Lb���敥�E��ZN�1�淽=w��	7�L�Q������l�Ξ��u{}?�ƾ�B��n��]�$6��G?j!K��n<�V��U���+��%�� �噕Ksߣ�>�>�яh��G��[�P�2���\�H,�l^��j��+	N�ҿ�$��컍����M���������}����^�����:��ox�w|����ϼ���[�ο�|t�䅤��^�ۍ^2�L���y�W�A��i�;*�x��1w���|}}=�`�v�3�닲��8)KW�Q�>�QF�3�*a&���ֶ��4m�BQ�����ڪ��ԋ+]C/}F-P��RBp4�'TF(&����г#*���ʵ5Ź;��㏧G�������1x��5���WU�T�T�������b�V����G4���s{ �7��Ua�RK�ʴٶB���ʕ+q0p㑭������ʲ�}H��M���<y¶d���IH�c��Z&����3��*P�P��J��mmm;�b��tڱ>�(�r0Xt��[��G��>��������7
�7�?���l�8�@u���o�k�>���@�ϴ(�W}�ղ^~%��{1�5'�q)��i��$I�V�m�{8�b#AL
�`W?�z�� ك^��E��;-�n�e��f�ҖP�Ӗ�N-���R���T�����.ky��#'�Γ$��I:K��*��b�JG�r[�N�ZU�[�Ngc>��D�w{�'ՓD�^���YM�v:�|ҞTyޟo���[����?��-���ב��� �U��c��ϴ_z�ԍ?�����{{��c��</�K�/��hT�:uC|���k��ֵ�aG֎�G}�bs�ɕ�G����op����m��`��;q�;v�w��[���o���3<��g�ǎ��jrE�$�(���L�8�����9y~'#9�z�x�����"�S�i���j��	��<���8���)���x�}��h4.
�P���W��y.�q��W�*}ӽ���[����|V;�Y��W\�J��������t�k⸽v�ʕ�<���9�;����<�&_���M��nG�EbdT�;-#P@��R���a��y*Q���WJ�J�9�f�.�L}/cԿ�ʑ�V������[X�l�*��L�x���Ϋ�q�J˪���"�2F������g�'�\�����^�V� 1���'�k����� �%�������t:��H��</�Y��(��(��|�Y���]C�Q�~�@Mxű	u��ޞR�-��*�Y֭�Mc"�<�z�$�CL����l1	Z_3=h�	2O�^z`k��X����~��?\bN�	��Hp*�ٲS���ړeY��Jh�aO��G��b��s�(k����C1W��_���`b���n�+�mca.Ea���A<��e�g�I<�LM���m���8��j�!,�� <�v<��Q�*�g�@Vxz�_,X�N�mJ:e�ZhJ���N;�X0���]n<m���n��'IR��z�,}<Y��6��T�N��}��B˶�|\�����z�(�~ͦ���w�\�W��a�n�&Y֚��^U�$��dY{;˲Kq�\���b��,'q+�fU<rU9q�V���s�<Ϧs��ؼ��/�D�����f�w������,N_�4����s�>�%�{ݽ�ޫ1���r��g��[����h��o;v��w//���ڵ��3goi%iZ��?�_z�u��	w��E����*���s��Y��Oژ�9L���S�np�z�8y���nqq��r�6����2~֘�'Zv���K���nr����D'��#��o�:dSC�vU(O(�Ue�����p�������[���e���c�^������ǡ�	M���Nq�ߧ��.�(��2�����C�;������������/{��O�Վz/�������|�D���t�<[K����=��mnn��j�o˲4Ue��gϖ/�˕x���(��mw�w�~���cy׹s���R�j���Tq���}��]��v���f�Ф.�'�p��U˪��g�O<n��.Zy>%����4��������n0X�Ѕ#G��	�bd,�ǂ�͓�U���塔���SV�`�`���p_�&�e@P>��o%h��{�Kصfa��T�~�C�qQU�,�$yu��{-�����VJj���DĪ�Al$̵h����HyFm���
f��ĸ݃��:8\qOzpB����c����Z��(�Oq��u�j����ġ�E}�~���g�<�A$�����-�������B ����>$����ޣ>�Ng�]\\��]��P�Oy��¶��}�]�`P�Z��]}m��X��7�`��a���[������	b߄�y�g� 
B����ص�5��xњ�G`>��Q�Ċc���R5HB���w�w�b(I�c6�u�{~��\}�lc�\�O��^���L��u�waQw�(R=�:^�`1P{������󂰮���Y�{t�����Tv�ݓ,K-c:����d�¦{�#��e�x�4M��E�4汋�.r�8���$ُ�h/��^�ZmM����*�QU�q�W�عj��8je��s���y�-�E�ϊ,˪��A�yUe{ډ��I5�v4��c������*M-77��8]�<y�ZY�*�~�����~xn��|�����'/��/�G����y�`���')�x�j%����N@�e�V�B��l�E�l^鼩Y:�#v���,?������z~llͳjEek6�f����:�v5m������|�1.�k�M&݃{o�'Q��~�錿@D�8�g��c��=��iԚ��Yke����i�<�R�·j�X5!���������[U�5�Z���Im���޷v�I�R�w�q����+��;���R�����(��s�>]��U>���"��O�������ޥ���}��_\�����0���[��l�����ܑ#G˳g�Ə?��m�klO����[M�nnm���������ܹ;�r?,ϯsG���J��]w��Į�Q�V�Ú�m�w>s�V�}�c��;n�����7g�O%��خq̋l��k~����ˢ,��͍�7~�7,o��U9�v)��[اnL�'Kg;d�6Ԏ�0k�K;̃镩����Nݍ7���[�'���?�귾�>����W��_1�{����d2�vV;�ѵ��8N_q���{����$�B���q��m��f�2�������-w�q�����*��N�(vS�T�˵~���9���P���x��q++��ĉ��Ť��j]���/_�l���_���K��K�/�Օ�R������|�ķ���N�nu�J�^{u���V?&�%:��[�Cj�=;�!Ճ��]	3�W�^�I��ջ恬's��lIgϰ��m
���o�V['���-.zqP����gW��z���G�j�Y��D���e�=�M��o]O��5�Щ��{}�Aܒb�l[Ư���Z9︾\��8`�;KP��ыm[�>#Y\$���������@��{�9xsCY�0�����^�\�O��h�h4��}j�S�/!����(a��� �O�6(�&x�vc��z#a*���lץ��y�5��Ff#zA*{V?*VZ�݉�^���>FK�J�hů���P�Z��}ɓ��B3����W5��^�o{�칲�K ����ņ��[5��mmm����g1pIl�9O�&�_��oj!8I���Bb��kaKݟ�]��w <_%�j���p�/��6�\������a1��e[��EL�_��'+��Tj��}�cгE�_p��O���Z��a0;�b#��L�DY�}B�j�\����Q���;��p��v�T�bk�S�0�:�Oת&�i^�y�β|6���N[�e^z�}���X6yQv�=ݺN��z��W��'I<�YY�8N���W�m��2/s��)�ٝV��Y��iEQ�ɪ��4ɪ�|j�5�Nm����J|�ԒoK��~'OY�dU�đ��(ɋ<+�"��?�1P*�Q�Ω�S�F�%U���W��_h9��/�Y�¶؝i��/�K9`�|>��H�V��,J��2b�<��yYUc�dY:�NgC�[Wj�5�Og�B;�v1�N�Y�M#�&�y1��,�#7��|��'�M�v[;�U���·z�n�]>�fUU�V�vUN�]Ͷ��Z���u����nlT�kk�����������(�����ҝ[[����;�\���?��C"^�(6~�����v�l��*���ޮ%liӘ)�A�Z|�Ue�sy��qKZ;z�yv5�v�}w׋_l�Y�l���	�v�l���~��x�V�A��:tя���_ph�_V[*U��P���z׻��K�]n�~^x������o���wm�o�՜�-
�|��_�x�	�q�j>��oz�7��{���?��|���
^��� ����%�I�:�:�.m�YYy�'_���q_+k�yɋ_�:y�Dz뭷�흝R��&MGj�g�%Eɨ�=�ʋ�.I��ڲ�!���r8�Wɶ��c�T�,T��f�<��4W��_�'k�D����i�[�u�%��cǎY����j*������7�x{s˟�����߿��d8&�wv��U�����20����`���i6��}� ��B-�}�\n���0�G��n��~���3�;��*[�eR��8���ݛD�ڥ6�-v����7ݣ<�>�IIj�u���g(�3}F��8H��is��{R�G��Y�ф��&�Z-�Z�r-�B��/���9t�~|=n�D`�	����WՁ<�p�1�����&s��b��$]j?����D�v�YɄ
	M	b��a��~���e�j~��*_��B�{BK��b���bD��gDqc�~�@1�ynI�O��Z|�m�+Ժz�7Q�P�C��r(��=�~�d5%k����=3�=���B�>^9,n�s�4qFaa�(�a��O%�la�nY��`#6I$�-$�u����F��]���v��vdG�NH\Rey�N'�΍���ښ���l�]��P!3z��;]�۠�,���*,�$��@��ؑ�m��@-�F/y����A��g4��ł�F���P�y��Z��,w���Y������Z��=��6�S��z��[+ܬ�yf��~K�'�J�q�s��K�kl�c���|Ȕc�M��g�:���F\|R��r��d@��q��󂗫��河��cٵ�#I�E�Ï�4K�{9 t�zqe����um�H�W�D^��|6׎�A������(�?�N&�Y�a��R�9�N�$�4ǖJ~�L�~gS�d�����vi�g�i�)YK�Zy��U��gu�^,��t:1��������9��J��J���*�~�j�QX^]��4=�6��ŕ��Mr@��Y����ͭ�B���Hĩ�L'6��eY�'�����f�r����</�QU���t6�t:��l6.�bE�$��8�6����h8��,i�:Y<��I�����D�@t�n��St��ߚN�?t����n��E�Gܤ�+^����c�{��^w���R��Vn���ډ������S����#��$�._��n:}�yx��N���n��X��q�9�ͭǇ�{Y�ƒ�=����[-���V��a��9*���>�H6v���/��S娢P������'Vh>�g�.v�~�ؿ�Nfx�un��H�$��ċ�;~ꧾ�;X�������k~���
�_��_�>��ϦKKK�s{�<�W��u���x4������0��VN����KV22��K���"/�*!��5���K�M�u{�-�����hT�J��<y����N��iG�N^��e+��c6m������(h ��B�Y� �H���e��zo��;ku:-y}�;�t_J\�
H�OM��M7���8���V|��&MF*q&Q�kx�n�A59�^,����%�D�y�Fc[�x��� &t:����'i��������=�A Jh�E}�{�0�6.~ҲrjÑ�z�R��)�L���D����*��� �T>E�v�s�G�c�uj�x8�IT"�DW��ja�'d�S�A��jF��%�)��(W��@<_`A�{��K�x!`q�
��g���l���-��V��]ha�#�*�d6	\]C�ӄaq0���������U��M�g���t?����'4h�$��=�~�֓���0n\�n<��^�kBTv'&�d�ŗ�/�Rۃ���p�P��4�Wx�~g���Z��N>��8f�~qbBV���~�� �k�P'o(�Cu(}�H�B�BF�ۈ�x�{��_���O�p|��-O��I�+a<�aW%������a��g�o�w�W?��{v*��V�~���|�^��>��/��4x���Vq��{_�ӿ�;����[���� �-��(��*�}��d��^�܅�	�-}i$%�&u�?���^�_����E�����?�j��Yy����yĪ���u�P��{���P���;��Õ\�;��kB�����eu��o�d�agF�ճ&�	�pz���摐��2��v�mI���)+�:q
�    IDAT����Y��z��W=O�N�Sja�C��c&,p%���aGF�=~A�j�&ZN�w���7>�� ��~��>1J�� ���\����V^�r�Ǳ��5����Va&��v����;kA���S�N���-s�h���!ۓ��!J�ʗ�;)�Jz��*��vR�zE9��}v���4����I��2/˲�&���ӓ�d�����V|��[�����;v��{�k^S./-ǿ������cv�k��B��ɓ����Vk���f��h�ꩧܙ�g��ή;v⸅4Y;j����oq����������OBQ� <�����w��ͦ��9�<WoW�}�zhṵ�e�h+T�*��/��/���.�s�.a;;�^>�Z�Z�_�@��x�FXP�vy�k���{��SU��������������7��q�ϩ�}���M��^�S����֢,�-=�ą�������������a�N���$�bN4�����D�]m�?��S*� �mm� ����z-�q���d237�ԗŲ��YH4@���Q�s�����Ah����Y�vJ��g��ì��O?�t|��q���W,NW_͛�Y�����+p7��(��2��	sm�j{[�;?H��M7�d"[<�:��f�'O�D	m�	���4��B��o��ګ��ݑ�O�l٠���'�6�מUMn��U��~�^^���Ԏ�&�ڳj����:T!�����i��U�&L4����щN���$�x&�U��ϼV��ZE���յڛ�aZ$�dGj��>����(Kk�a��[[�N��ˤ{��).K}�'3- �	-1����O�Q���D����q�^o�=�v�L�:��EJ��'�N׽�>m�V"��	�d��V�u���G6MZ�2�{��	���݀|n:
ێ�y��Z�*�#����l��*�����8� ��=�0�á3j�1��5���:$�� �,|C���	���>R_h�!��d�SH��5+5���	�S�|�1��pr�eJ��|ȅy�����v4�{���[����N�_���eĞ���h�@m�݅�L��+���/T{u������Ņyլԟ<��4c�,�<�/��������3Ʊ��L���El��:���Ś���K^T/���v��ߛw���K�Mg>!5xHâ���!�%xyU�%��aW(0��;"&tK+8X��z͹1��'[(QY_�k�Ì�B(�v]W���˗/�Yc�8����cA�	�^xK��yAs���b��
[�XZ�{	�4�T�<�د�Xc����;����x��ֳv_jvtM�lX�����}~'G�-�k�)O�2�g�JI�*�?A�����gX���C���ة1G���X��իW܊��,1+ɕ�"�8�Z���Q��i���D�M/�23vU�Z(�[�}�-KKK3��j\�t;�B�&��U����s7�xS)�����;݋^t�����L4��\<��Wd��SO?es�^�B�ҷ�rf���:9a���ٛM�j����v@E��y�t���k׮����W����ܧ�>#�>X�C�hüb��`W���z�v�~���=�ȣf�g}�=��{] �:$�����P,�5��-�9��gϤ���!�?�O��~����;�ę���`U%}���ϗ�)�S�����篏��ߺ�����)}������%3i%��U{ȴ���>g+)J��	�?H��I.CN�$�V��gӀ������L���(,�O�B$��+w���vwwsy�%x�W��͍�:)Ǘ��Jy!�3LD�xJմ��
�taKO�S��&ۦLӃ�^�/-Kwd��m�ol��+T����ow�.]2���J��r(;��VĵU���ζ=L���[lҳ�ʺh��*��cڠ�Й�^���:x�o��%�����Sf�AK����,�����R1����@����1�A�g��C<��,����%{���?�~"H�7m��*���`[Mcl�EV�� ��PIh�y�b][�C����<��{�h��P��A?�#�~j��@U�Bp�n��X��~>���7[��4��w����-O��c�v�b���Z=��}/��A?��M"Iό�B�>�0��޳n�
e�v�dbq��;�B<��U��S�E���=E�'��:�Z�n��A�t�-7Y��{˽w��o���DK�|���$̐8�I�����{|���[��x������>��L
����gܷ< ����`������ɮ�����/�� d���:d���{Y�7��u���/���b^�_�%b8|�]Z{�$��,���z�+g�>a�ě����}�R�����z%ԭ�h&��%�h��Wي-0�0"�OϺ��: İ�!o���%�󃒑֤�;���(bK,��� sbԡ�U������^{�C|y�M|�bB�l�{��d/�b���5,D��Z�ڡ@��BK,�B�d�I9�l�\Ϟ����|L�2�C��Ⱦ������Ʊ-f�i��k�{��3�{ް���B��V�Ǣ��0�Td��[B�G��6�~����#�X!/�|8N_��>�ּ�
]p�^�m\�p�k�n6��If
���׳��������h�Q����B��Z��L���C�|�����A�$�l8�4g�z����bg:��
)[_?��O�~؝8��������?���VsW�3g��m�/v����'��+��M�	^�5��O��PL{njի늙�;	�GyĽ�k_i�Q���^���L,��r�n���,��������D��x���^]����=�P9P���a^��E�9�*y�˳7�U���SO�Ν����u��|�7h!2�#���v�&D���n��҉�_���~i��uC��}E�*4��O���._��޻���O���&v?�яzO��оjPTb��?aF����m�۵�&��A^��M-�g2)��q�j�q���O>�d);��FK������@��'6���ñy�?� t����ȑ#��1ඍ<�"�J~[Y]�%�����GH����uْ�5c�˙�|���cs�V�a�NBW[�2\m�ϡb@%h��J��o4������&�u��䁓a�_6�E����U�	$}� ��������y�*�V�I:��%0��+�V{/���D��K����\��O�yh�~����v^`��ĵ<@��~����=�uHB�h� ��lb0qh����:	}a�ǻ�W�P�,5�(���O��!�A��{��V�ru&��!�q���r�?��>F+�;�\�pѼ���b���Ja7:NZ	�����먅����F��lL���^�5�t���'ݹs�,3X"M�y��	[T|��pǏ��lYM��{̾��J}�c�?�^w����>�s
T�DL�uY1�Iμhӳ�����?N>L�{�CB�8Y�ϡ�-]���S���>�W��X��ｧ?�0��PB,�y�,9�{4�ת=�A�A޶syX��K�:���{���[�_(�v
j���g8�ə�X��xe=!��J~�P��~�8����x3C�v}�p��}�u�"�\^z����m[_���P'�p8�~/�u�{��Q虰�x�"���������4O���q`�Z*t_�����R�E��q0a�g�3��� (C�Ex��(=bX������{}^]�Ǉ��~{�5O�:�]Wv��7����ٝo�	Lg��U�C�tȑJ��H�w!�"��汷�z2��K���£�5��>��':��%�`U홗�A�����M��V�Sdi<���Nz���C�B>,<��N)��3�ɤ.��żBq,��Լe�6�� &�ލSm��ص�)m�o	�v�]��/�X(���}��ti��$��*g�d2��:"������{�|����㛿������>����,�W�^�m\;�U��F}�X]h�����X���7���7�t�U[q��/������~���_�2i�[�<���۰z�`�o-)ܞo�{#;�Ї>�~�߾ׄ�6�j�Y���K=�>�~�-�Ü)[Ҏ�W�WYy�K�.���U9�W���e�ݶg"�)�nA<�O�#G��+��O�r���������}�3�������9�umƕ��?}�K_�-o�ѷ/�G������Y^�:�V{JVS����2�+W.[�ݰ�J�@�z�݌\�x���gY���w��]�%�]�pa��'��x�қ�$���y~tssS"֎��jz8Z��:�,��z���g�ɤUO�*7��	��`�K�	m#�D	��%��[�a�P��젆�'BH(I�I���Q�v�A��_�X�G�'ݿVg�:��]uf�	��}���b�>�&�:s]"��V�y���P�A�Q��W����4��j�ı�C�_��g��#�����?4X�3�U�2���mnnF]'l����8�Y������^�x(G��B̪<���t���AI"L�f��2�s�}�ٕ�<��Ӗ�xmc�^D�ٽ�:�O��"L��<���9�V	����j�dC��hP����:�m�{�%����}i7Dm�HW|�&�n�5� y/����c���>C����c��� ��#���؋�����v�Z��=�.zo�����a:~B����@��P�j��'zI���e�!FU�B}�Ŕ��W��{O]�:x������۝��A��a+7� vW
	W�'�{>�Vs��>Z�;2E]ø�&�V�]�2�����>�&������Xz�v4��D� �LI�݋0Ä�yur��s+��4��r�>a3��p�R�0 M�����-�\^�:V\ai�CLX։MV�^������8n��8��]{0}ȄّF�"[��"�	ֳb��"(̹��i��{aK[������"&�b����	�ד
���l�j��]?\���y5�(�T��؂E|½(����y�1�:�w��g���%��b��*(��i���f�ĲU��Y�hŪKR:�u��V��|�,_������l!�z�v�Be�R#ǂl_s�v�R�6�h�Q�v�4~*LO}l㴅:ڂ�	1ǡ�;���J����٭vv5H�8��}�Q;h�[����}؜E��j�x$����I���/%*Q��~�aw��Y����n��vw�����׼���D�e�0N�/������~�m���*=�q�r`��-�x�=�!�浢t�=����_��<�
��s������Wi~������S'�������ߖw���x�Z�j���㥅E��`�MyXu5��̦/}�P���������{_p���~�m��͵�s{-�A�w]�|�o�����s��N�k�?�'2{��[a��^W�^�%�|�5��t�n�����|6�t�8��v{���������?���ċ�;�����t�TU������f�7����^4��u�8�M���E�����z�`�*3����A����Ǣ����m� j�nirz�
M<�� �B �8��S1�*�&C� ��!`�=�}�Q;eM�C̪���VW��:���I�<��=��^M+k�7�z��~��hҐX���nw���Į�lR�>�O�w��V~в�k��Q
=xv��%`���0����Y��z�V���c�g��e��M}�Ŋ����y�ud����i��`{�δ����I�[����������I�\�SB�&��Hu}��{����'9L
a�>q�Z���ާ�k�6�S�	L|e?��:��W�~�[��~��WF��
�I�y��(�'~���u�و8��$J}�}��ڢ�+�T�m�r��bA��[�V.��6[���n���o��be���Bu���-��Wu�{8�1�>��Y�v��������o�9�'���q$�VO�Y�CW�]����L�#�h���u_��2u���xӻڙ_`�e^��`������O�����S	�̨M���)��3�m����K`"ӄ��5Aja^h�f[���F(QX߷��m���01�1�!8�9����=�S��	��&�r}R�����;�q>\���5���WL�O��]�L<�Ƕ�1(�"��ɍ�$�:�ل���P.J�5����B��a{c�A�G��x�=q-\+�j����#T��p�:�Zs�v�B��ƌP?��-KK$�)��V�u�;�o"�s���*{O�r_$Z}_�C�B�����>B������IY�܃0[8�B����ϗٹ]}-YUX*��\UL���iU�E�ƨ�W��Y��zs��c�Y����7���-������p�b�yV	��!&;�����I��m�m��n�ɓn2��յ5����k�í�`%��
 A��m��c>�w����`P/f�ck!Hv����.x5��I�-
O���w��-�|%�~e���
�/���e!����w�����ʝ?����?��}����p����1d��0ֆ�����p�/{�ݿ�W��M�u�ó��}��ߝ<��7�y~�|>����;�$�s<���vm��m��򖷸����v��g{{[A�*�*~����o��gΞ)O�8?��c��ŋ�nͲ4�?y���x�����?﫡?^j��K�������v����l�X��EQ�M�7�ey�,������"/��"��y�)��2L�U�X+��v��C�a���i�mKiwo�\Z\�A4��CB�hH:��D׬=F�B��-�C��X�~n�o"$L��]H��u�t�zr���ղAP�e�֓�ek��3��$�=*=3�M���b2UZh{g;V�j�X�O�Q	9y��`���W;8�N���E��vS�r4Y&t'vh���U�Y\$�4X��tm�l0���>�Ė���� |������/1?|`G*o��uyֻv���)i�S2�&U]��>�5ē^�����MVqDO�)q�W�PuA}��ש������u��~��{�������~'���kK��vj����$�c��y@���rnIo�F8�D���xl�Fؒ<��jQd���'l�}�~����Raj:�N��A�!(����Hq�:�Ӌ6ُ���[�WI��vG��Y��$%�~N��Wo��Br_����ra�~nq�
��L���l�m�y�$��*�;��hѣ�$}o��u�q�>�Ӯ�
�[t�� ���'a��L�䅟/�e�H��ض{
��2����I=��8� ��sۉ�$iz�.�-�/T��$Ϻ$�a!*n�zM����PBc�� �C�Cr���-*�m�N%FB؅��ק� ���uBN�<���M�-����� ��m�R/���z�^�g>P�[�����`���y}5���vT}�B/,`��aa�� tCIɰ���,��-���Ƌ� q�*E�C�܏Ma�/�؄E���ױֲ%�ݺ�Gإs��{�1�w8Bl�?�����0���b��m�3%��l:�-X��>Y�v]W>x;u�V6.���RK�Yj�<��z�!�0P"�5+'�q�ۿ�;lN��?��n4�q_�9ݗ�=������U̶Xh��SM��yr}���=z����X(���w���'���ͻ��='�ˇ?�Aw��;�j�Bj&:l��N�rԵ��\Z��s?�c?f���w,��6������p|�-�?C�V�Sc����?�G6�������t�����:��q_�u_����5;t������Znye�<}����[���B~�W~������'��}yQ���r9/�Ţ(�W�\�
�sébſ,,.)���0(F����[�F����+���X��{~+���_�ۭͥ��O��.}oQ��>_���k�]�]*�Fky�w8^j����n�+�j0�'K�8Y呢(��l1���i��̦�SyY���|1/򥲬:q)%��v�ݲ��|��n�b��(N���IT��lނynɚƓq)qy�,�������E�|4ZT�V��Z�R��G{L��v*��7��y~�[Ž�����i�qQ���h�/.,��N�D�&)/��@����Bb�2L@u��	a�VP�.[d��:�p��yO5�k^k�ߟ�Uonn	���>}U����H�V������5��3��    IDAT�'q)�Q��r����Wv�&����PX���������C���Dq�ڵ����kfξ�ުM���jwz���A��h�0��T�<�E���u(4�q\{�ԗ�_[�{{�୦�� �<��3}]��`啔=X-�y�7�v�<�q	Y��2yu��B���O������N���_�
[�����(��{SMt���bM����]ً��*J�a�G_1#71��>dM�W�i�V��uBdJ��RR����	� �\�����v$~��
�
e��!��x*�e"N�]��>�6�	�i��za��p�������DT�(�B�%�ڢ��A��8��5��mϺǐ�瓖�(�t/���0�@�Fa���0����Wտ�3�1�۲�P�-�<�V�d��|��Õ!4.�8n	Ͱ�o�_��D�-@+�~�?G����U����S%�+xB%����X�m��_B%To�/NB2�Ć~�qG��}�̓;�}�{<Ǯ�Q6�*a����-���*�s_&R	����R�������&������~�����
B��c�M�-��sѱ�Z{���}թ�
���1t�`��
�FJQ��$��h4����ߍ&&/׈�Q�DAЈ��RTC�u�N��w���^�1��gC���H��O�n5c�5�?���?�^sɱ�l6߁<����ٽ��z��&�=��#�o{��s�w�� �f<�p��N�ѱQ:15mA�ˎ�S{�ҩ[��xF��������իג�����hFU�s�)'��������dcp�@�ə�m6�PnUGf�H���BQ�e2w�Z�dC�.��2f�?�	x�5dKQ���_�4�;��A��O=Ų�ۮ��� _��ivv�9�X[q��}���d|��ѥW�� ��W}M�Z{_�Kc�K9�$��J��7=3����պ�kQ�C	��Ɨ/W�o=�'xS_�����j��-�c�:2qe����՞��뺻�����^��n�6@���'��|��5?�.tw��F�U��뚓��.�N�w�$���4YM��Q�t]JiX��Wk�M�>�,g�h4�l6��Y�@K�`R���9�#@�D��X���P��q�����bҾˑ�H��._�w㔟D�%��}q�j��"�ʫ&&T�=b&��_��3��9ڶ�`�
*��2�t��LX��� b�1�N~��Ȕ� �
�
��e(�4㈇�l@i4N�^��b2D�m,� 2 �Ť�4�$� �RRF�ͳ�u�ܸ��cLm����:�&��-�[E��j(8!��UI�B��4a��bF��`��ƙ ��d�)I�?�ĵE�`����4�x-�/C���hA��s�[@��m�C�T��H��3)��{�^0�1�7�j�Uin���4A>��eH�� (��2���t�v�@�
�@j#�(|��Sݔ�4~�����B[�c|�H9�`]:��<m��(��s�����y�9�ŏ���}pT�d3��1� ��	I�c|��h�D�qS�a�(��~,����t	��8�+QV�RiFcZ"�X����J�D�ؘBd��.� �
p�9�om����l�:�	�9�S������z�(6�z��i���'JC�?㬆S6A��q~�5��p�q�Ԙ�?4�a��v����u�i��6�1�$À� L�8�(ж\��0� H �A;�e쬢���l+<X��h�s;g�F~�,�_�CqLZ����qM� �q^Y���	��ctw�V�t�e�q0㡇�#G��=ŵ��##��Yͩ��"+��t�t��={h���F��h��M����bz��J�����K)O����t򺵆&�m�m��"�#߳4P�{z��=�^�Bi���KH�g~����xqN�tw����_y=z�G8z��fh��1z|�ڼi3-[B7������b�r���[N�r�Uk޴m�6S��m���c���7��߈�dU�ă�r�� �N������l�ru�֭*_(�X��+�i�����$��>u��r[`L��уC����8���d�߼ꪫ������{������f��k���������\=z�YN��QRq<�墿=T� dP��=��W(��$I���f�\G'�II��q2�l6� X�CݵZ�����g�z�-d2�����r�V�N��,b�@���ӎE���l�hGʹ����� �X@D:�X꤈Ns7*ȳҢ\e�C��p��3�Wn�X��-}�%��w���>𹙼��j�|!��i"j�c�57`G��׆�E�Z\��ڂf#�:��ϒ|%�(���B�, &4\�N�E�Wu<ϒ9�ET��q���ǿa��ŝ�`Ҩ�@e6����-+������]�\���(T1ϝ�,��Dlq_�-�	w���g"����\��GD8�iS���Z��+Y�!����=Fď�
��(Ѹe�
�)�8��c�D��9�Fc�a���d$3"����i�(p*���%׾��t�i�!� h��J$Nl�4���a	(��J�u C�7��l���9�XXę����� [�k��� ��gqQ/�4W����~�,��q�Fi�4[ިP&�`�o��I��D��Kj#���H8��]Ÿ��K� xI&ׂ{��5�^�wzj�����8O��=6�=njp��Þ����(:E�1�97�g��A5@\ L� r��Z�A#������Y�j~+ �-�F�nV �s�B��]R���1Q��5�y�E��!ٯ���	K�2��v�c% Pn�9v,Aej~����gG*8۷og�P�(� M���3u� w�t�z�V�Ɲw�[�M��o�Hh�f|ڸq3)H�q��E����}���E�֭����tp�`�B��(.x6ca�!#C��7@���P�M��rn5�ez�H�ϲ·��|`���_�?[p
 ��4148@_���<O�q�t�_7L#'�Eψ#�522��_�������2ww��/��u�֫�8�K�����SSp= ���1��B��.��M��P�
`�Tv��]]��T*N���-ǡ/._��;۶m[���;���/�P�8::����"ʋ(�R�LV�� J
Q��@�p\��]�rǂFcyWO�x����LO�J��oƥ��2J -\��I�Y7�7VC@Q^�� T�v�(k��9�f&Il8�
�#)d𘮀�]@/k�FaZk�X�#�ŋ��n@V�۬�:�[C�(0@8�"%���V��j-��s����� `�c� �X �hS
-Q�d�l�BA�jsw-���=�.JU�����p3ޙ2!<nȈ�!��H��\��ɴ((����51(��b9��/�Z�,�	E;�P6��1�e"ͦ9�|�d�h�<�����Xd�0~�I�ֵ-�"�(��9c����I�8.RD�>���+i|�!H�����(����������=�,WfWY��&d l�� �6�� ����� o���Ie�c�l�	J�d���pі{#���Lx��"P�ӮX8��[�U� qA;R�o�L���Vj_�����>E%� fӍϯ��G��Ǎj5�@Yʃda�L�v�9v8���R�䜰�Y8�ss�,�%t(�|N�8��3�+�W �P`	3vlL������N�c��F��Q����T*\��U��7�g�mb���B7��8�.F2�.]'��	+�&���@޶m7�	�1�8!��a`{y��?y�A�=�u�Y���*R.\{�K΢rw�ܹ�9��>8ppl�F�ڽ����~��d$:��q��=̩�O��Rd))�r�Vn����m����ˈ﷾y�]������"��Q�_^i$��Ҷ��4hAMD}�#�Ҙ�������$��Ȯ|�6L�t�?���"��CC\�=2<Dw�yk��t����u4�b^4�a&��}�}���q�Ҁ��A0w�B��$�."rr�N�ayy^X��
�B�b�
�e��w���U��v:�x���������=<�HaB�!��֪�Î�>_,���7��xa������	JT�����=�W͹'N$�^�h��T�����@e]W��f�,U��hl��HGCI�i�9��F�!6;
��A�aA�6E#���ʂ)IP,�E�)����@���)�d8�*)]pC����6c��l���V��*�qQb�j2��pÂF��q%�U,�~�"#rjd����>�V��*_[&��
^h |&j~(����8.2���!�q[�-Q��h/�%�!I����av�%�`9G���2iRP%Qi -5���}����	�ߓ�$w�s��Y!dx����f��qlt�;;�R\����I,� 7 �5 �E��w��!�g,� 6bo��.B'B
�p<����,w�4z��g��p>�7�C����lIQ����(�dQ-ʐ�NH�؇���".��8?�A�3���a�n��G
Y4�Q� \h&�2c��X��}�1��QN��@Q-٭�0�Ծ�Z�����Z 9KC�2�UDI���
���9�:� �2�!6��
�%��.6��YD�%c�6��4�`�̩�L�g�E�h.$�yD8,RH	�e�z�y�Y�L�ų�j����1.N���t\3�
Md����p��8@���m�-7��E+���[���-�m�Pi�����B��؆Zţ�-[N5M���ݻw���]Pl��:��s8�g��I�~��'�������v�߰��(�=u��-*gU�PgZx�9��wҚU+�l/׮������Ym�<ԑ ���j]�����]GO��e;��A_��[�?��C{��}6ҎFK|tt�~��d�\ֹ�M�Sf\����0:�a�ݰ�pw��Y�H�qS����W���|��۶m32P/���4|���홙����l�a�����3HR�����ڲ�T����s�qN���Too/��喯����%K�T�X�K��]�F���)um.W���o}��p��]v,��B#��R�=�玌Ī��7�f�K�j��u2I=ȇaҕ���j���h*9�"j\)��Ѩ�SJCQ��fɀK�<��5�x�Ş��6�	�.B0�ZL`[�WC��].R+2�zl�ִҙ��� �� dtr�+$�2��t��&H�!J&�a���/�I��  ���J�� �T�s��m�"�6���cQ��#�.86"���p'�(�yƈ$��(q@���/�R,�(�Ĺ�8�B�aY�/�J��D@ �� ��jժ��2"|L�`�R��I�d'�b�k�"��ַzٰ�I�ǭB3�8Hq �Q"k(�d��3�upF� �*ԘΉVZM"���}ʽ��6�� c|�o-� �{dZٶ��)�2ET��)�b��Y����Փ���L{z��J�ml��1��8l� j�41��F+d�Fb�����@�����2�H{�Z�q] �8�D��N`
#��d$��x��~�(�:�n�� �A������q� hp?3���p4}�q��W�_�0���$�viKmlcim��L�z.�a ���F��?CxN}Vw������y�F��Ғ �?��r�ѱڷ?��g��̰�U+��nQl޲���>�%���ldd�Ќ.�)^��كw��H8�b9��5�WQ>zGJLW�)� S
,M14�-Ow|�Nz��YK:�IwG�;�L���,2e�K�Dq��O���5�\��433E����l�Y�����N���@��?>u��8ԥr	u's�֟�t�蛶m{��/Ԣ���Pg�T���&"Q�N� a����}���������	��k_��ڻw�i(�G�g�f�Z��]�v�=�o�b>�1�r����o5nng�X�c�����t��ܩ�(���W
i&�t �t>��b�2��
��Q�YiECav+W�DQԭ�����(sss^�\V�>�2B��dy(�0i\�,8³��2�Y�GS�g�!I!�r�'NS�h�%������i��E�������sM�� ��\ +�OI4`D�-�}n�NX�ܷ�_��q��U� ��yJ���F�`�s�x��Q��c���x�ϋ���������E�
�m�/��[I�\�iD`:�=m�е���hc?���*X�*�����t7$`-o��N(�_|�.,�?���1c���Rpi�Ϙv��.�4��5�[�_�"L��k�����P_D��&Jk�D��k�'n��%8��4���j
�&&(�H�[��]��4���mw�l/�Pc+l�A��ka�j�j�Dl�����7��}��ڗ8r<���&]�n;\�	� c������Md eB�0��#�I-�A��f�c��9�ڰi�}�1�s �����K+W��@G����G�+���}���QM
na��k���?�7�m����a�y
��/�⢺��:mKg ^pxW�\���Q[n!l�w�7���B�������w�G���o�k�f���v����j�?ae��k�m�1�P������M9��j?~�Q:p`?m`����/�2=�ē�y�YNA��S�[صq�7��uo��B-p��~����v�|l������8*�Zz�zzzZ!�r�S�ի��G��-o�C�2�Su�}�� h*�	�^ !ɒ�͑��g��ɹ���������r/��;��X�c��� �?��O{�n�����; ��b�����x٬�9.:,��sc{A�\�\/St2�@	���>�SCNJK�T�8F[�|���4M{�8�@_'���G+X�Ez�6�E[�B��P�"b���z�j#ij:�IT�F��i͙�3��ߦ([�#Bq&�(IT�6lT���,`�st��h?(9,�,������3��H[�֒:�-����"@��ٔ��n���DG���RR���k�[K��k�g���g�0 �c3���yxo~a��m\�_�ؗ\� �g�����ب78��,���)�^�߳6mp� C]��m�L =h{�$(��wbS�hfl�5�5)�o�J%Π�8��#VUD(5p��G=6y� ��d��+�3�\4����F�d/��7@��b^�D�\�t��5�p��}��,\�p��]�S(�՘�n���X�N���B��m4��طs���@KPC����=s��e�p���~�X��r�͠c��N>)���{= _�s��@^|��t�w�Ӻb�Jڽk7��/����Ɨ�s�x�}�z�Z��ҫV�a��p���-Y����yp���d̶�CD����{�T,���U'�)�o�Ŝ^��YѦG-�b�� ��#�0�͍t�%���� ��{��}Z�b5�un�t�k^M߿���8:��O���e�^���P����N�z[W��˶m;�B������Tp����]�f�r���GC����vz+��ԛ6n�ӳ3�E��b��:��}A
ixx8DǛ���(�����<����f���ڵ��/���u�;��X�c���#��<K(��=D�w����g�755���\�U���T� �=�O���A�G���8�Z��(*&��Nt<D)��qܣ�.%Z��Q��Q1
#�+f�|	�h�R{�-WR@$�yH�-��s#� ;����q����J9VN��=є6;�X|��X!t�F�� AC�k�9�à���*�%Ϥ�m�N|�����l�8N�CY�)��7	������~�Y93\8;0q��J�v�,�5���p  0o���Y�BX��42]tX�"B|���-_�����ՑF�WtŲ�,;>0�� ��&��s��x	g��0l��e���kQ�,Ks���#tM3v�0-��_�K�j7���+���Z�.���Ǳ�C�d�5W("�8��7�@��R�B}Fmڴ	:��������e�����w���vÆ�t��ws��W^I��w�	P~���� ���o}�;��_
=��NZ:���8aJê�k����:ۂ<�v�C�����G ���u)�DS    IDAT)Xù�����>�Y��,3	Z��=Oэ7}�9��
-�Kk,�D2�ٿ|_���|�Y��Y
���^u�JVg���_�+�/��O�qjg7��x�>�e,�-�#���uۙ�Nz�+�����s����gsa8s����Q��p��A�~�RQC�#�y�fDmibb�=թ�i�����⊕+�|>�jqh����D�Xxd����f3�ޡ3Ȕ��۱@��ǰ @��w��˻��{{�R��LNN:��7P�9i�f
�DU*�!j@��#
�7�Bܤ�
Ji���&ITNSg�qh��8K4�t=�I!���8U&�!�V� �FҤ}�U��"�)&�k��1�$	��G �C�ܵ�-q%Gl"��:X:�I�k�Z�	V�F��-K*�e�L�֤�h�h�0f
,v�2��Dy��2
��{n���h�k@?� f ɼ\�� ����6S>�\���h�f8�F�(�e��'�VQ`��X�l���"�U��­�يV�s�Y�]�[�'�08��]�/ 7
4��g"`.��Ç��A$���/((���x�RQ]�2^kÁ�����-�n�M7��^�*����D�W^�Jo��}��g�I7�f��������_��8j~�9����w���n������z#�$%n<�gQ<j
5yP	������qt�Tȷ�hL�����xl�e�F���� ����t���7h�n��rP�����Dt��+��o�S2�}�O9Ҽ07G�~��p��. u�v��I33��8�����Ü�B ��p���㴗����,�u�]�_�N�j����x�[��/I!;�a����i�ӸB�5XT����{�n]�ꢾ�^�A���zn\.i��?66��\ד�^z�!u��:�X�c��~x6~��' ��MW�\ũ�Bov6U==�E�g|�O��a&� ��E�<_봜*���@F�Z'�9�l��a6���0���N}Ju6b���Z�$ ���m��������B�0E��`D��t�4%0��#��{�U��qc��.hh!XY�����R���B8�`�B#��~V!]my4�x�2JN��v):Et�z�oF7J۵u�3w�h[�h$��r�����#�x� C��4th&�^&�!���C��C$i���Y.B;~b
tJ=42�N�z��׮����Ϡ���raa�n_��ӧ?�i.�:�sSC������g>��֎L�l�@�s�}ͭ�`Oњ5�(��wP��v�	K�f|��xbGw����)��"�����raG�5��TjT*wӾ����چ��q���ӚD��N�X�b������ p�*x~O?m+����w�#S�_���1Rx�n�}���d��o��������e��ٿv]�/<8 ޅ���u�r�w� �{zj���{�r�����484����#:�#<<�����5%7��}����c9�����9D�t,б�z��"4����7���Nw�s~݋"���mz��4]��������n�*����䂉�U9��0��g
n�Y˸����~1�υQ�#'�d2��8��:N�J9����ϓD�w�DY�y��h���Q�j��d}��G�<��Q��6��Z-��a����8�>Q�t���i��u'I�$l4���?����.;iԛ�|!�L-��xs����޾�l�pх�L�K���'v�B�� �ڻo/�4׭[G��'��:��x�I�g��/у<�Ō7n�Nk���z���MR*�^ ^r�A�q����R�C{�즮R��"�� ��B�¶���V����nŊ̥�(��hph�����1�5�FŃ�ö���q����۷r��hX�4��;��;\pרU����FG�i�[hnn����hvf�c� Ƞ�p�j>��]e�?8x���z����x��''������(ʙց �kxOU"~.�^4#<���0�|���s�kpp0���R�uNPJ���|1�����^�tW�郲�:�X�c��:��-�\r�%~�1������w�K�8t萪իt���>�����˖-�cG�ѓ;w1W-tQ̶dl��NLpdzݺ�h�S{ό������L��E�+WQ6��/���H�E���}��RW�D9p�S���a�F�W	�2�_C���s|�j�A������̖�cѭ)
��X�	�Vi6������^8�8i����uk�Ү'�����Z�n-_(I�̴�5�p ��_�HM>�G�n����B��Z=�+����f#2GDs�פ76n�DK��ӑC\�
PD�!@����Р�`�RJ9sD�wV�X~�R�[���������;�X�c��:�X�g��ygo�rpd��s�9w]� =��cMPW.��B�'�[�j5<p�*�ˎ!`�Dr!�5;3K+W��Ch����Rf��OP3@S L�e+Vrњh�t���?����Y�`ux�(l������h�_���2>���v�~����[��+^执�Kb���y��㼆�`��I�j�ϱ�߿��}��J�֮����;�q���Q�����<c?t8Gt|o�Ÿ�
��������޲m۶�g�o��{Ϲh���?�~ff�=����C��bQ�*�h힘��7�󱣓4�t��$���/hӦ���ΝL�.�(l�gs�=��7
ݟ|!�n<�u~ӱ@�t,б@��9,��׽�ӳ3���.\;<<J;v<�*S�|�+�>�Аb��-��G~đ�+V2g���+WҡC����b�
zj�S��h�4==�T��"�;�l9��zZE���� ��8`��o����(��Pk��*<�Fi b�n>�z=��+W���Uֹ)wT�����O�t�!���\>�z�+V��O��'Y��𡃬Q���`����d��&����B�h�z6_���w��m����������W�f/�I�3=�M5+�@��\�<�
�W�a�8>�vD�ќ�W��5H����uk�B�-v�Z�AW������(ow��:�X�c��:�X�y���/9�-)9��7��g~�J��6m�{�<�@Q[���ffgi͚5r���㓓x�FG��ѣ\�p�l���@�^d��]��I�hB�,��h:vl��8����/N5��LdW�9DiA�(��8��Q^J]��E�����0��t42x½5Ňk7�>�z��^�:�"�VْFCT�X*��� ]p������!Z�g}�ۙ�EtB~��A�0rlF�$	�l&�5�q�\jA�ֹ��;^�~�9�{��-���zsm��z��u����^��x�ez~a�/��!�a��("�`�ׄ��Ç>x55M���➞noph(�������|�|޶m��Ǳ��U�t,б@�t,���׾�m�j�����wu=��N�P�@70���?�>1=�����L���	����[����P��r�*:z�e�9.2����.[F�b���"Œp ��`�!:|� �8���A��ǠwQ
�ʋ	tXſ9\ʭ�xk�]��e�˝ۚߴGk9H��f&x�#����q��B��󐑧��~ں�T�ȇ�;����:1�l~���8���<k��f5,7�ynFa���\���n9~|�7_Ā�Fwvvr}�2wea�FJu�i���5����j:�ܗ���I�,,�ѣ�X��Z��͸��K����>���΢;d��4Տ�Z��׾��h��:�X�c��:�X�c����^|��/��?���V>��Cܵ����tOO�B��U�z���!��՝�v�I�Nb�U�92D���8�T��Ӭ���+"�˖-���"��"͏�C�2��]�x�t��e�l���L�4�3��/(SS3�����)N��\���!m�ٴ�6�MG?uTO��9l���*ZF�Li@�������t��E�]M�8Nc�#l#l8���~��i8}}��T,~����_�^�����_��V��,,� ���U��� 4guu��.��e����Ao��'Og�徾�����w����7��Z��C�=���\܉�>��vggt,б@�t,`-�K.��T*���+�t���q��8��GG���!�{�}���hϞ=�!2��p���Gi�I'���,Dȑ����z����4+@$V,]:N��L��!~-�)x�)9r��8���~����	 �^Sdւ����:3�	`I2�̀���.=zl���������"x��k���Ip7�!̞�m�r��Vڟ�uu���.��`?�W����A�she7�]��q�С�����NDw�F���G��o;es��s�7���7������=���.�V�n��(�=H�5�MZ�~�\�����Gs�s4;7G�&'��뱐�e�]����52:�,
*��]CCŗ���؉�v���:�X�c��:x�-���ι�����\r��AWػw�[�Dm��8�����]w}�^v��ȣ�p����4�t��t�u��׼�5tםw��ի����c۷ӎǟ��O9�v��E#cc�X#�be/�y�)7���"iBG'�0ow����pV��sx-45=���u��p4x�l��8��ǧ�o��[x�7��F�1P3��y0�,����MͶo�/���E�T�e˗�`� =���T�����jFW�D���d���0">���F#��}� �7�j�^Ԁ��??459���V��a�>�}�Zoi���ņ��;�Оr s�B#�a�W��J����}�����n�JK�.����ۺ�����7�y�y�v,б@�t,б�/�.y��o����7���C�so�0�w�������y�]t�%�Г;��s�9�u�f^����W/��v��I�~ի8Bz�7����}ڸi37�cJ@������lk�$ǔq=��k/��� �W@o{���e�4pw�]�<�ڡj�A_���|M=��� n]� ����jQ�L�/�D�$�D�YxtϽ��+9����n#�!.���M�:>�:�Y��gx�5���^6��]
���o�-�7�<?�xq�[o��w��£�ssK�MP�����	A���ϸ����@����	��"R_��u__���W/��E���������5��e���w����Od��;�X�c��:�X�y��+~�����������W^y�ɬ��c�կ~�~�w~�@�D��J�J]]%V^@��(*�� �*$������G�j�z�z��~G	�X��~��F��6��J�đ�~�8���Ѿ]��J�UT���5������o�����?�
	 � ˠ1@< ��<VhX��J�`���eI� ��l�˿�1AM E���}/�n����TUDo��`�f��z�Y?K�j���YN9������Z���M_��m��9��^{m���[?s|�}33ӿ�Fq'��Tƥf�(�ъ�/z˩[X:x��/,�./��A�D�5��������?��O~�\n���|�X�������Nǵ��Y��c��:�X�c�_X\�ҳ~wpx���7����RB���_�J�����733���l6�tl�47S@����`)2l?|�A����X����^P$h~v�V�]K��܄� �̀)F_7�#�1ww���#�&(�o˒�L��������\
D{ҭ�~�~��G���tȖ9sp��ܘ˟�R�1 .su��͘��j�#� ��ۻ�������G>�a�H4u�6M3��wV��Y� ����3>�)ͺ~����t钛�,Y���o�����ߛ���h�V/�H����I�F#�(Lȵ��1�]�����cG9- /inn�2~�&''������}����_�%�} ��}wp`����w��_�y�s�t,б@�<�8��3~������|�o.��Bu�豸Z�y_�ڭ������RWw72�t޹g�$U~�aZ�|�ؾ�^��8z{�ofY�C��Be��L�z{�h~n����|�#�Bi ��tx�l��"�ۮ��x���B�����(�P3^���۾~;M9�Q_�Mњ髶���@j� ��f��
:�sx�>��������W�����Y�"_����,y�����Ӕje�����)�=@�vhp �S���w��׽��_�y`����>⮿������WU���A���i��г�W�
^x�"N?�tb��;�#>??�r ��"\~�gқ��&ڻoo��_����Ǳ�%_���}��W����گ-MS禛nR���*533�tuu9N�Xu���L#��O�Ɖ��|a��m[,�I���߶��&���Z�Ժ�b1�{�I�V�W}��ժ3���$�T*9�|�I�57�.�Q�8��f� �l6��� �r���D���D��?lA.h���*��
Z:�F5\Q��)���2��1U��ņ��J8�a6�n;v6�L����������������I�5�hNe�9}J����J7u�<���{���6��y?���tV�ɻ4Ǡ��~+�v� ������k�1z�јH�����8'���۳TZH���ڟ��{־��p?�����t�n��Z"�����MOO�����g���^�w�Qq�o���7]N���_l��Ӊ�!����ްasǎ�M7�d���s��W�gj���S���3>�;v<�&��fgl��o��3�km�oέ?��_���t�M �ɽx�>��W\�p�m�����:��X��g����ĥ�^�C��#G&��������~���g>�Y��e/cU��/����X?u�q���op�ђ�KX��?��
�>r�������t-_��x�'k��Xk���ː���*<�����O�'���J Z��a�����~�V��_`�+���{_қ��\�Vpl��Cm�8���� ��K/~�$�G��@n�
:GD�z�J�n�#G��׿~[86:��F�z՛����C�y�8������N-,�Uk�Dk_;�B;���
X"� ������-[���E3�3t��16�� A��\�����Y}�i�х]�����}�ݕ�=��R������C�Ї��� �^s�5��<::�lߞU�穱1Wek%�����y���*�Ӛz�8���@��n��r�v�$MpS*�IWW7t�u3lROW�`���T�V%RJ�<1P��
��@t_6�u�A��j�f�k�z���C��`6�71NC�2��͐�Q�I�(W�^#hdr�\6
r�L�l��q"����3:�b��L6u\G�@g<��~�[�R�������(vc�F�����92I���AS�������0RH�tuw����j�%��=W��ϟ�ku��2(8�z�����So4�B>}C'�"?N%��y��d2*�b�/���7��X!�����2�r��(L�z{���
H�2<?b���Tx��AS�ge���N�֍F#�}?�V"��
yt�I
�B��J�$�i�FhONi�Xk�7����8n��e'MS�����\�Y(7͸���D�4��0
��J\�&�Oy��� [,���^��J)��V�Q�vK� ���7�͸P�QGn�Ď�p�f��l6i4Q.WH���8*�bS�I��^�ѩ��>D�1_�$��^)כ���q�Ui�T�B��n��ƈ����-]�����̶<c,9��\�j7Ց�S�M�ȅ 7~��
%!�㩔��s����K#/B~\���$�x�`�*�B'ՔSrh� 91��u�$r<����x&�lj�HD�x��b�9�G1��D�r�a��e�Y�Z.��2~�fq�4�x�(�x|a�<�G�����2��8��0�>[=��0�Q�����H�4B
�J\��Un����x�^�g=?Ci��b��ԫ���0Iu��|^�bc��Iy�
�X&�~�i:�������|>
�(I�8q]7�=RJaHi3�4�q�8�I.�m�1��u�</�y:D��	��DI��J{��?v]�T'�#�s5��U*m����A*4���O[���p�$q��*G"Q�	"S�����:ѩ	RyG�_yY    IDAT1R���qL�Ps�i���K=�`����T��Џ�J2Ik?�M��|�� ��"l��l�O��Z��eSE|����X�Mgg�i�\�{��XJ6h�,=����������y���,�8�%[�����_t�E���aOo���S��[���m��LLжm�8+�r�
�����yƙ��#�pQ��@?=�k'}�;ߡUkVӉ�i���e��(���Dx� �*\D��С�n �J�c�-�0kpL��!`�`n ��u3v��d����n�� �f��N<״`���em�p��h���P+z�������e�v���@]@qZOw7U��yM�9���SS
�����]����Ë.��je�w�w��G?�����o�������s�s�A�C�������N�֭[ǭ���╯$��R��fff�/^c����l� �7n̝}��4>>^߻�����S�?���[�Թ_�x�r~v��5�L&Ӻ�l��D��l��r�y ��֔Uq��X.m����j���\.��0�fg#���F��]|�X�q�a��@1bΚ'Wh��uY�8Z��j�h���2$פ  �\N�Y_�����wvvF{^FA����G�K��(8��А���c� �I�BŤpt1AZ�D���Z���ˉ�X+������/&&"�k�}B��[�������f��`(p��?F!������rڴ8�`�G�/~#������,lR���$���/�4 %���n~~^�㞛�S�&#���V�� X��86�cBDS�\�`c�؟|�{ �{����wao��|&x�'t������u>�W�8u86�L�&W)]�U)h�v�d����Ts�uh"&1����mp�`\'������a�P,h��;Ʊ�A��1�1�(��I���	���-'ͤ	�&�W��9fi\'�>�3�����m&pI�{�a&_�V�o�(e|
F��$ &
*�X��F
萟�4�}�u'��y��p,D5\קuևN�p��㷉r=7FL�]tH�ٶ�<�0�	�P�+|f��0�1`[&m3/b���O��<'�B����PJ��"/F9�݊�Ɨ�V�q�T� �_���Z���DkTO[Qy�2�1gAMp)Ld�0�����>��+���1�kP�V�k|B��,���Sȵ:)� ;��|�pjI���Y������)��B�)�k�/��8!k�z�BU;�m��|H!E��'G�p>S 0;�M��8~����(�v=�n�WEe����	�P�DǾ�����DgQ?�G��Lv%I{'��A0&��h&�uS�N�&iC5�r�:��䪦Gn��;I�LRUW��<'��V1 y�P���0���i��@��M|�Q�����F#��siVt����رR��ۛ"��� ,«�����T���K/9`L�A�'����_�r�韾D�r�&'��W\A�B��
��Ɨ��đ#�i�&��룹�yھc;7d@���D1sz��-23�7M4Gr1v�ϑ�ё!�A��0�����Y��kR\�v�=���w�N�ٻH�0��v^j��_<���6YG�״�!��Sb
�e�]��ׅ��c<g�o��
P������驩x``��N'��>�Ğ�^���x���o{����<��Z��v�Nܨ7�Z�Ω���q	�$[�T����16������=:1���D�a�Mؿx��1�^������=�:E��r����~%M	�o�$ �]�.'%]��|7����ӛ���.�s��(���cjvf1�Pk�cp䴧�'�Vk>�En:� �Y��a@�S8o����yH�R7[#����A�ׅjN��B�@a1�����10aca�uXb���\c�(�  I= �b��2����3$SG�@
��:q��z��TIl��� n������>����>r�g����Q�i���q. �A"b�Q3 S\�ѣGi�ʕ|. �x@�8R �x pM��j����T�9�罰P���0p<�1��ax� R�;�'�/:���{�X�`W��{�,^�"B�}�5��8�o^��q�����)C� �s�9Z�>h|?�!�n��Q��g������ ֑�-M�����#�+.�2l3�d%ep\X�-%�3�c���up��
�]���[�W1����=���&ZT"���{���7D*��k�fjR�a�l�g��g�r �Rw�Zx��\�_��M�L�y��l�$�ϠOY,9j �r]�qj����{CV  �ύ�h���8:�+��U��&�\� �1΃�S�9Ž�����:�N��-pfEB��u����E!� E<a�u]��u+���'�2S���-x�xqƪR�Y|az�'�)χ���ր���(����4���
qAsN,~�hvg����MA-mPܛ���u�����0o�;>�D��	ǘ���|����1pM���g�JF��i�H�i���XX��H����Q�^E���|>�	�?w�=W��\��<�C�qJ�~r���N�8���")Ju���G�JE)"�C��D�$ҩn(r���T�(�%i������8Z���$qY��٬��l-��r�J%��d2Ŧ�9�_U������ew�u^}��'h�m��C��
"���'m��8L޸d�R=;;��G]{�����#~q�m�1��Z�K_�RZ�d�׽;n�ˀa�`�Y�|9
�鶯�Ɲ��qm��R:����U �\`�5��WC��������`�Q�`
��x��L濖J�)qd�\�b�m9��-_���wP3�����Dy�)f.��(`k��(r�?�v�"#�-�4�t���N���Ut���;�Q������6p��R���P�(�es\�P�˗��4=�"��l��ڿ���U��w7�pyF����C�v���.��:��3���.�s�=�M��{w���ƀ���zsa~!�ROLLx� ������!ꈭ^oh 'Dp\�Q�����I�D̿�A7xfz�#f�yv���!Z�h4�v��M�p#��a��[�Th`p�$&3�#�!n>^�:� �Xx�� Z�Y�!@�  ��7@"?�k������:G��m&o��y#�h�F���@�����+B�����Qg��I����(��<!b;�} 86b�?�M$7��X�(@���x�s�B'dx�: ��a�Z����ʈ΂��4~�- �b�,� v"�D���7��Qk�e��Qk{�X�%v��
:�3Z� �����"���`rCd�͘�t�ᨑ7�3�|\�7QM�"���Y�)���G�6�@ �A��<y��k�aq���d����&Ƴ���\@��=5�Qx[8^&��� M���OaC��#g�1��s;���@���%�3�� ���X|��j�v�bW�[~���CZb�/�0� �p��1>d1n �˜�~⶛jd~$R��$�v>1�d9� m{�0�����Z�3��`��-��B!�?���3
C[�#�A�C��:"�fnr[c��?s/���p=�^!� ����DtΤ�J�����c�b��=���NII$�S��Ea|ǟ�>�XA�}O̀iRr,� ��8&[rη�n�)�vc�\������pk�|x���F&+�`��e�`�x�A�Ü[�Umƥ�Y��Z����3�6s��x�1k�#g�Z�_���e���6���=�S1��ԅR�4�r�US]]]�V�*JAڈC�z�X8�����|N7�D;�Hx�Nk*'��0���zEu�uq'Q��䲹j5��F�V�sٺ��CGU,�&ݦD	�MW9L@�Zk�?��Q�1�U�J3���0H����UiQ������I�D�S.�I&`�T*E�%^&��bɇs�IR?L0���Qty�$��r�
�"8�����􇆆y]��;�eN/��g��Gx��K7���N��c�	��u'����iz�ǏҺu'�S��r
4�����]�H��^�k��ݻok�/c�)��e�켉5�H�Y]]dM��!��%�혊�2����:��4�[�1�]�Z����Et�8c�4_��$�'�8ñ�S4��N�y`��6�Hg�c�9p`?gI��������n�˥�����֭=��/���6Po�ᓽ�Jp�\��j�ޥc�!%��y���*���)���e�_N?��}��餓O��[Oc0e#�J  �u�Vo�~&^d�ZC��J�0���p� �k�׌)��8�� ਏD������J��f`fE>���(�@�pG-�e�gB�&����)]���	nnn6P<DXP�%�� =bDD�9������T<���"��Q���QE�Ϥ6L*Z"yv�jE���_|�S���We� 6�"��#��1��F|Z�g���<pD4��"�!�G�# E8w�i�#׆�`�/S�Ώ�q5�R��Ga��op�v&�ց���q]x���A�rL ؖcpKö�R؜��&����^��/Q�Z��)S�	 @����G���Y���"`�Hv=�l�S@��l���:;�n�k���׀q
�ՠ=ʅs���	�b�c�&�3�]a�f�'��Ǒ���s�#���#�^���xA �R���3#Nn&Y���$�+��+�hk��b"�ߓ}��D([��ǒ�n߷L��o~�G *�,ƥ<O�D�1��x-��a8��z�ڑo*2�g�����d�-O~'`��ff��xk%��~�G�ni�H[�O��=m�^��aGc>��yv��4��g��e2|���sC	2�R��,��xN�csD��5)�Q.,��L��`˽�h�DO��Y0QM��V�S�~8��~qdUz��Ⱦ|�s�(m�z��L�9�Uh#��k �F��g�eC���K���xʹ	��Q`�/F��$�/�L�I�fƺ�k��u9Z���PC�!dXN
Ͻu� ��,�0;�1��e'������p��j:k�r���l?M������#�)i�-7�'&5P������`��u`_x�ڝ5�Q �{�4�a�5�y�L6C
���?��b͓��������3����L�4��$MsP*�g�F"����M[�����]�����]�d	ϝ���?Ӧ��	��U�V�w�^�^�@�����N?��.�	E�������"e`���S{����e�\�"l[�2�M�Lp�k�8��F���{�����4q��薵�X��v�3��k���$�]��81&�������^.t[�j�����,نc��.�,�����Sp���qw��ozݶm��Ǽ`��Fih?C�y��f>177�J�qLf���GyD��p�)���3����ן1�ݴq�/�8� 6��̴j6���hÄ�h4b��x�\nh6�
A.�Eڇ9���3��J���L� 8�W� %ȼK���r��O���D�o��5x�.G�lAJ��	���nY�\��h�/��-�R��SƜ�C�� I~Rm:���^���P�S�QD+ ��"� E� I�pUmO��x��p����
�pē&Hh�4��V�v������x-�@"�8WL�f�4(��JTGƎ'-��0>�lp�+�PNÀ�������i����j�ٴbl=Ԟ�22؏���/�͢�ץ�-`�� �x��8�k�3�k�M�{��X�5cc�A��r4�'<<lP�Hg|ԏ�D�'m�^`�=�����0�#v�')V�vP�}D(DBj� ̀���<F��o��D�e�2�C�Q0���#��ޤ�o���4��b�t9���sԓ��R{�K;9�͸�n�QW.�8��Y
�r�s ��A���Y�J��3<l��4R� ^ĕ����|��Q�W8>���S#mڈ;-[�=���ϗBy����&Y~&��R%r�V�OT�!���3;�XF�8���iv��rx���07ro�8aG�5� 6D,�c�T3���T+�l��P<��|��&cc����aZ�(�1S�%������1��v�q&Y��SC�O�3�!i�g��e� �<W�a���# ��2ob54* p��tXz�����`=0��3�U�'��uq��
�ǜ��sЈ�
�\��533e��c�|��|�Fb����	����5%v�6��ƸGƖ�a��8(l� �KH�	�9W����5܀��8ˆ��q�p��Pr�ɼg��mI�~�^3�Z|�e���d�l�2g�,w�t3N��`����!T���1@������	�q1����"������Pxbjʇ����XX.w�?K��w��UA��T�Hm�X�=�0w��#M���M߻�ڴi� ���:������]���@6��D�D���=��ъ��Z������)�hkO|�������r�w``������&�Ʈ�n���Z(��2c�k�:H�c��~�L� 6lhQ&�?��zz�[����P#�,	Е����\6o��������,��Ol۶�S�zA /��O-�����'�f^�*Յ" ��^ea>��8�w���-[�z�7m�`����zU.�tOO�BԴ��wZ!b�IX��� ��ˍ�dc��M�� ��*�yR�d�������HE!O��� a��1�0�W ��m���Z��6(aDCp�"�� P �.<���H��2�0�u�5&_��?�\�VL&�CHD�D7[��2�.G���v��#E(_�Vc/U"	�� E	D\m�!��,�uM�!�"O�(�G��ky�dBC-��/�t~-��+[p�#�-�2��H.���-;��5��O���"	���`��`
[��L4 @�/�v�04���"���f���� ��-)H���,� Y�`#�_*q��D��Z�Ţ����ȍ \�`���ļ]K��}�"�i�'��� r�X�%�K�>gM�T :"�<����8yѱEY�d|�u�)���:~�J�b���f��@���������0-N������G 	�*�-ֹ�g����m�D��B���8���م�ŒC�y�yq�P�}��m<C�{0��K\djsݚwL���T(T��[,�g�����)<3Zl�[�qq.����#����0N�M��{�t)��g����1C��g6�e�)�1��8Ѽ�[�,�n�<�� �/��gF��b"��$��(�E-@�g�(�1(�4.��费>����������ɺcǵ\/� Aqh��Fˉ�G{��y���2�8�:V�Q�)x�H����1�����4�uDB8�L��0u�=Cd�D�����1=5ej&x�4��m��α�� ��
��}~�(�����^�]��i{�#�E=��F+��G�:��f�5<��Χ��ź����(���� cj||;�w<��0(�}���� �������h�L/
%��m=u+8x��ȶ�z*�������AI��dp�h�;�����r�:^���(q��ӷ�����l�Moo?}�#JP)��mE�-M��mm#T��.��-�+�
۞�
�$�O�[�����vev�<����K:15E�J2���e�=�z�%�.w߲m�6+���K~^� ������̆���7Q��(�ʾ���4�''������s=�."� ���l�������
*<�x� �	
�.Q^�Zٺ}1���bB�F>Q��h���T�D!�1 i��ǖ�?&�V��V��,�g�|Z�"��V�E�T��4�]89�b�D���k��X� f
f��*@�6���n�C�*�:�#6f�d���V�(Y"�]���t�Pc����Ij�������MմQw�M��ߘ4%2�E�B<S3��V���U,J� (�s��5`R����H	v�	q?$j�c�|�V����ʌ�;�K�'������s��7&L�����B������VH%=�O"r1�{�N�����Xf�    IDATB,��(>�B�g�h�g@�����.(����Lt�<�o{om�u�w�sΝ�\�j��Je��ɒ,��ellc���lpҋ��:��������0���Â`��4s�n�-![�JCI5��7�������w%�4�ut$�wת���w�����9�����!Z�\��%��,�ƚ]��_ǵu�ְ��3��b��l�!>�}��:*�x����v�k�8=m���?�u%�z�_�gL���ř��ƚ����B�(ˆ�AV�Xh��x�htp��[�2�ɭ[��UH��b4n���݅r��2��V�g��r�B�u\�DQ��[�J�xǄ�4-2��&�v��VKs���wu�
�*�hz_�ww��(�3q�+ޗ���~]�L^b��Rӊ�tm�@��/��/�X}��_�C1���9]#~ݖ�;�q]:c����s�����6-�qAnBRYl���ן8$�^seu��]����\�(�ğWj�牸���\���r1w7�=�Ŭ DO����O����Ҹ��N�t|��GA�>n�g5V�G,vEF�Q|��ƍ;xq->W�8��\z����wB&��̜�g�1���I�'��>�P�U���;\q+����~��*��:b�J�˦1�9xi)�|����㧭�Þ�{�̸q�}����y�P�%n�B";|vl�n�i�{�X���J4}�+����K.�������̣�M����Y�#Wm3P�9Pׂ��vm�ύ(95_�<W�Ţ�m��?������>S�]��)���4�}h��Arr'����c�l�Q,S�������c�?���֞|z�<����"��Mo��ܵkwPZ2�{H������ڵs��+.�^y���s��;�y΋�yx�2�[
��W��=}v��?w�uE�_"q�]8w�%�p���̊���J����T�&W0өS�L�3~Sh�d�TJ)��#˃6M�fEP`8�V��bj(P�IG��C/�rsj~Y�ˇ�����rŜ6�h�Y	R�0=Z�y5�Oi��#զ�D��}�.r��۴v�:N	f����(��V�.d�y��sT/#3��XNPv(���P����ɧe�ln�k��E��h6fu�*=V,s�IȬ楕5�dŭ���]��x���A9�r�1����������[\���[�YTu<.�􀈮)]˧�mk�^�	��B��z�^�~��9L4+\|`YPX9��"I)��m�8�]�?D��Bښ�-���~��J��/
�!��8[�8�U�o��[��<��-h�a][|K��J��͢�nA��syϏS�x]uYr|1�~u���a:-��D���/�������E¢̞1�ϺHt�eT1�b�����K���/0���,���R��a�VH]G���HG1눻�L��޾O��^��}���P��]'���-s�:���<������%���� ����2��[\ ��Pב_#Q��	���[���5�1���-�����[p�~�.����N4x
9�>���B���7��s������]�;W��4g��S�E�ZL��7(,��(Ztyl�_�f�/.�bI����#=��nH\tLΕ�ciTs����vw���W1S����;�:�F�v�Q�<�s��S?m��<ϡ*�mGf��ֵ�{A�V�	gϝ���'xb o<n�����PZ��1�4Nhg��p�j�Z���yRsd������g��}�tұ��&$eT��-���W������V�l��=��˯0�{��m�S-�&C�������y��A_��<����n�)?~�D�b�$�/��rOYh!)��m������4��ʠ���y��m�z�w�����0ޙ�����l�����y�tD�9�M�o���w���/��̀�h����-����ѣ�ʩŃ��׿���W����,��e�3��{�}�鲱�iX�2�?z���t{��w�y�_=�\�|�W�����_���ܹ'o_]]}O�߿!I��|�w��ևgΜn��1Bzue%��-Z� ׄ*����:�)��y�t-��DdLe-�0��y(ߪ_(�W9I�wܺ�?'���V��V$JH�ߛ���u��ض�����$z��r_4��օc��~�Y@]���r6�SZo4Q�z���*�ӑX�m��d�*�*��L�T�;�(ʭd�J�����+A���z��>�>yF�.?�-�LX�[��>��K����e�s�GD?�迬IK�ī^�O���=�5�㼸m���'M���)Mރ*KȆ�\r�%��A���8y���*�r��I;V�ww�q*��ϭ�jC���C�����u-�t���-��z��t�J}��c�����H��E|00��]w�e�P�G�����o���ͳ-G�^ѻ%�-�n�T?e��XYO��˭7�a�<wC$�~��ȥˏ>#��ŋKVvS�0	�����t���N���D��5�Ā����lg��tK�k"ָ�z9w�\�=Pu#qZ��,״G-��,iхE���?l�j�]Y[�q�������[e�"��P�ndSq�}���1�{~�1�{�_�.$}^���fv#&"� )�?.�ݲ�g
���c3��VMw)����j{��8WO���0�Ϸ��Z\f�`tK�ϑjӯcbޯ�����/'���5�~���&�]!�Ϫ/����ͤ��B?,�]��n*�%I�q�DڄU>�=,}xK7;�-e��s�廇�bj"&#���e,c�Tt�YW-0ls��2շTBV�w��k�\�.L�j��w��5^22�F�M�E4 h<d4�	07E���-p��Ȼ{r��i�F/�ɬ]�nx������lP��_��_�ڟs���oxc8�ȱ��s����%��n�a�,���9�H��W�'��_~��$���+C�XD�x�8ȝi��=vL!���^e���?;V/�]�$�}2�ٝ�
{^[\�(��6�{���?��ٳ�L���-P
�I�.|��3�Cl�nV�P���8��-���n��3da���f����h�"�gΜ�D�gϮ�������F��?�S?��χ�}�6^�[N��'?�sמz������H��������I���0I���5-�Dɱ���/>\{8�.8��{7��5a���a�]q[����Ed���ߊ5���mY&�m'�m�̳��k�����!l+J�\ʠY^<�I}LB�D���Y�K_M�ԕ��v�[	b�-}��X\�U�_՟�]��ͭ�:Y}'�#��[���J�z����D4�O�V���$��#p�d���rks2l��E�ڗ���Jɧ}�1�zɟ�3]hB��dM�-��Z�����6q��r�>��ֶĨ&p�����+M֞{W��{��J�K J(>|�xk��
\Ǡ�H�Q��OA=����A�M����ک����];�,ؤ/��������Շ��رc��k����74����W_m����u-������>�*�z@�I"Y�ݷp��-V�Pb���������ĉ��z���UjG�� �-}��-����xL��U�S��D����4�%@�b�_���zU �c�=n�-�g,ǭ�D����8�=�����gu�zi,_s�k�g?��h�EƔ�w�6�g3�yh��3$f���x�G��9x������*�#x�q��е5kSׅ��z�)w��O�K��S���+���Y�kUף[������a��/��@�"��ח���+wAr�>+����9�~�ˈ��8�A�,�b�J�T��9_$�x��r˦��ntA�F�p��Q�Zs�)���lkm�v�&��n������v�h���d�,�\�eY�\�Zƞ�R�����wOI-�1?�^&fʬ.�'^ގ���y��l�Me%�������J�/
�w�ww�p��s�,��h��f�w-���\F�De�Q���������3%��+n�ǌ,�J2�R`�L��l(c!�~���E}|h�V�ŏ�TϬ����D��?C< ��[t݈s>�ls܉rk�� LҢAh[([<I���ؖ�Wm���s�ȑ+�G>�1[�J��������ݻ$�����P����s� K{���"Ӝ�*k�t꙯y���C=������4�[Y���C��tW�,Gץ�UG���E��i	N�'��>�q�6!!<�򅖿�\��'??@<���w��Y܁���rUd�ܹ��H�c�V~�QΝ?o��Z��ۖ9ix�K�_��oz��]�z��_J�g��s��	^��`���w����{�ћ���5!)�O�9=����ȟz�D�܄�V3_]Yk�"w˜Z�����s����mq[سw�=0v��m=D�ä_���utA��~��٘Gtl+�t���0��ߴ���EAY�l<BU�	ãFu�e����)�ᴽ�U����շ4�F�mD�4������?o�kb���Z��ru�Ь[�����/��>K���IQ�cYQ*�L��Ԕ	d��S0�Y�إ m���+z�[@[�e�B�2�`��'M�B��C��A��i��,�:w	<Mb�c��$:�Fc���$��a�F�-k����\L<�T������Xu7�Ճ��-gsm�F���Rol�*}�t.zp��ڲ���6ӹ�U_��ﾵ���B�>�1����B���ks�(���{'��t,v}��r=���d�}I�~���]�-��&tg���-Ϻ�}�X�j�}=Pe�ѢD����>��1���g�9eX)-�vߔ���`Ό����o�~Կ�[�����~���c��Ų�G�)�Zch����:�.��~�]/>��^׻�CYc|��=	C-F��,��eT?-�vi�w�d�/�Bom���*5-]���ţ����t?s�kQ��_w��_k����_OT���Vh�ъ]����]�.-~n�0��2�_��_Ǥy���S�Oٱk����RbR�Ʈ�=#�"�s�J�y�ͫ�[g���X������b�|�����x���Q��8u����xf�4�,�ʲ����,c������k���8Ǩe�m��e��vsA-~��t��Q^_:�]�:O��L��j'Kb.�~*;O�����y4BlY�yQ��>6�-�_Z�=@��CY
ܷT"L�������߹��]
�O��_��an��E�풕eԶ��w�,[GL%g���4`z�]����oy��m?򑏆V�T9�{���������l.���v�cc(n*;�����8h�Sc1��={���n������<��I4�)h9�Ceឿ�;,�φ�ϪX�eA��J6u���+�r�x���䘃~hk���o�x��&x'-�.v��f>�#���������ʵ�N���fS~�������y�a��WVqe�Ю�ⱔ��'Ӽ��d�׾�+��[n��g���o�����u�EQ$?��?����tsw���N�h>�/[^^V-k�:4N�<m��*��A�o߾T�.�h5h6�ۖ~Zf3��Z}�0�OexX�[ܾ��)����+�X�ȷl��oc�\�2?;M��ߖ,��o2P̬����m���m:^��%�c4!�L���3�U�y���/.E���M�p�ҍ�	��#�tg�����JKC�V�M�zx�LP�Rtt�ɳ�^HL��w��Y���=$��rV�D��G�}�p�t~�6��N��[=�f�MaY%�eD?5���W�b���hb� ��b�Wgm���r+�=��C��=mY<�\�>^�iV���1S߲@�
]�v����tO!�~�Y����b.��#�V6q�?�'V�[Y��>�#����,	:F�'4�x5=O��[�n��1�!/�ǭg�[�����-�-s|z�.���\zJ�L���U�������l���w����d��>���2�w�P�:o/� ������l��(la��Ec��I�.M�:o-�t�8{}F��u�Jz_�k��0;���zW�bm�O��$77���5BN�ܭJ�V�������HzO�D����t�� � >�7]�z�o��ѱ���ެ,w��ir�����J���u�רm�x�0W�zk��9T;z-.n7��}kS���:�/���b,u��()c���ÕZ�w/?����<�?�,���{n,��4��v��RV�3~kn�sG}�p���v1�~-��J���w���_ϲ���]e>�HǦs�N���̌��Ug0P�$���W�,,鿮)7.�*�1Y�Y�g��OB�}��[�=�(Q��P�����:��������zF%]�����rn;�V�3�����������t|���|r�t��n�U�ٹ��P����Y[�Yi��9��O�3KZ���2�>�S��{��{�/��/�˚+b�c��M��o����S���ǎ=jnO�8a.�_w�vm�ܙ�<(;pLK�3?��q��w�������J)X���\�]��?;7?�����'�`SY��m��o�wLp+��|�uW��ƶ/&v�}w���V�=�o���H�շ�j�
��~�~(��_����>��%v�X���m�w���ݘ"�>��c�#G�h�|�+�����>����c�R���Zx�� ?��C����{�-/�\�5�W�{��z���|T̮�������R��������0�RS�&���U�}�4��u��2_�X�(�[Q��)�*�`](^>�� �"�*5I�e�Ge�������v��*>�!��h�T=YK��W)���IB���Mě�d 0�[�q��+E��]�eZqp!f[��V�nz�cY|9������ĩJx��}�qUQ�Zݕ�n���kR�O{0�����������z."eM�skD���#�݇N�:���\}O���w�"L�S�׶m�zl�Q��]�W?��ǥv$�\���19}����Xsk�D�Y��̬�����=h˅��)����o.Z4��X�����#e$�]+ed��׮����������MO��aV��,��6��d]�z�Sx��q�_ҷ�}�-cb�������������x?DN޿[�l��}��g��v~�]�:�()=����`�N�[�c��6����u�t�Y}�m��,8�O�m��_�>���/�|�s۾m�xLtf�*ŋ3�w=����פ/6&���ʷ�}��"B��x�r�"��5�1�5�������{T}�nZ�E���ݶ��1K�����H,v���v}1��k����Ԏ׽��"��*2�Y�4O���c��zdA�]9�ta,k��]q��|>r�]۶p*s��X���L1�9[�-г&����Js�Q,���E�Q�y���r'Fj+Ι�O�ˊt1B_���ǭ�z��e���ЖAȪX%��A��h�p��]v�+IgJ�[�p���p�ˌ���UHA߿�Х6��H�+͛�o�>;��ra��[����>gצx��L��o���Í~���1��M;���E������X��ҁ�zq�c-�*^�by��U�+�#ǂM+�}����oyk���Q ۹kwx�{�>��o�Rw��Kh+�	^ϝ�u�b8�WX��Rp���*��`8��J�R�=���&S��X)���=�n	����޳�Q-�6���z�ŹK��qn�"V9q�=5;��z�d8s��Y����f��I�k�T�3�0����[�Q���������}��i��M�d����3���1���:v�t]�-�ma><z���;�x�/\v����]�x������>������D�����|���y>ؚ$�ֵ��-�V{g��q��j_s�̙}�Q>��f�$�|Q�������j_��&�D�~BJ���U��:[�M1�0�c�v<���fi�Jː�f�e@�D���z�J�p6n�mr�"&Ib�T�S��`�2��o��o���I[	ŵ�V���^�%<��^>==ee;� ��2&~�1��8!7-3��Le�¦�$Z�R�����=`���|�����ҫ��*����"l0����.�Ԧ/ZJ_QY���D�T�u�\ ��ܢ��Ē�������N�*׹�N?]�4������_�
��Rȥ%`�I�
@��׫q�7���?X9j%��5W�+i���I��ܚ�|;�?kQ�V.W�TM-V>ڜ��"fr�N�?��2�22t�q���%��JZ�<��U��7`    IDATTn���Ϯ�mj�Yב/�4��t����
�o��W����%|�`�����-�.8M$�/Ll�\���LG߲T	m���Բ�j��s��Z+�Q
G_x�;	{��uح�~-y�=-���;*x����˒�c�M�/����r��Z�!�uݮ�B;W^f���Js��LT��r��S�^�g�p�W���'��Ɉ�v�"��>-�yOx��q����[��=U�,}V��JQ@NZ��Zf��M�g��-v����8~�E�Ħ���� ������[s�[�\H{NaϦ1�H��c�JVef��R��4s_���](c;���}>>1��3S��+Ziշ�b�.In�йĒ�Q��q_q�\�T��*�s����x��C�?_�y�js��w�*�[n��3���g_�ճ��Z��.���~�2팜8q���(F�=�Y���xl1�h���_��E�D�}{�~�z�)5�D�������jO�%1�]I�᧟>m�
e�P���Xڴ�R����<^�ʫ�G?�1����C�,����D�3NCtG��TL���������v��@m��{���u�]oB^�x�F���ʬ�ʼ��6Y��ϚK��OYNc��ʲ-���R |S�zLA:Sڦ���.��������X [\�yp�3Ӓ��}R���c�.�ߋ��;v�P�"+r�{p~~���dY6����R�v_�Cs�v%4����͵�Si��m����?���ɽ�����JR��n���0K�E�|�C�����g�N���v�V���ۣf��o%���l,v{����b�_3^��vw�����P�TuMUsL�Z�r�h�[��r�V�+U���*=����l�҅�A2�k�U="�Ys���A%s�o6���v��EI�{�)�`�(t�0J�T�]G���<��N��rJ����~���ٙ�p��G��pmu�7;7�k�Z�S����z�z��F���;�3K����W�͢9hLgâP��~6B��!�.�%�(���Mͦ]�tVdYZ���os�Y�=�7���!��hk�Z��Z�D?C����T���d��L6���,�K}���$n�m�E�^S��Z�_;6��+.^�1@���r7MG�Q��3i�\���v�Y�	!\ظ�m�/q���e�;�N:��H�iVdô�]+���x���'�����NTF9曵ҟ�\�������e�$mE�ɽ/I�F�!A;lE�%�Dk�Qk�'ma�T.�)��B2�b*a:	IgT�Z�4�������C3Q)�����*�1����ǅJ(ҤH�������E:�U9���H�z��f:*���]�!��D�I��yG��H��DU�:���*��Q��jTѐ	%^�#+u�hC�CR��onnvf��J~�o�[k%�Wyo��%DTe�R絚��?̛�F*�[�4�����t��d���_[���1m���T�d�XZ^����Q�������^�A����/ŢU���8s�-�T��,`���x�w$�=��]E<��d���[��n#z/�����ʨ�q�R{�W9>6/a=�F�B�|����YbU��h�����Z��E�[�Է/R|����g��"�틴r!���H� /���
�%t�kf�S��Ō�a�(S������S�r�
@��/�|QMT�ڂ�$��(��՘��|2�2���1��lĩ�]��2��U� ��g�Jx㦅l���L�4'n�3�ڥ(w�<���[\	k����)$H�}��+�+r��w#��}^�O�$f�P���0a�;T�R{��X�/w��r�K��K������I�ƝΘ�ͅ�D��(�+�/|�N���bi�o���[_p��?�Z�-���k��淄}�C�{���G~4|�_~��r?�9ou�ˊ���<ށPW}��w�ɧ�UW�+�&�o���4כ�W1�����r�kn1��0�w�L�>��C���,#����z�^��\f]g�[\�)fE��&��j��:�(x�i�k�4h�������'�?)���S���U��V����t�33�U���}�7!o{�m��ɓ6�g�>m.�^_s����W_���#������A|!ޏ����g�2�E/ˏ=�Qb~��wz&��;��~=z�ɽ��29q�D�w��bω㏝ܻ���x��<�m[����,,,$3�����l��a}}6�gݹ�͛�p1mw;��^�gA�f;Z)��Zì(�Z04�Qa���ۑ!�F���lT���QZ�2���,ϳ�ʾi����?��,I�N��I�I���`��nt{��Զ�,l��}7K$��bX$�0
i�$Y�5�Ծ���wҐ֗�i�e�D��̋Q#M2��V��h8H��<i��m���n��4EF��K�d�b�z�Pw&E2i>e���1�HeW�[���lŔy�3��|���X�!�Z���&�^o����N��.B��w{Y�lHh%덙X�:�LO�.\�E"J��4Z�d4� ��{�-[��p(�?HF&�m����,���2X�!���E�,�ZtiG��!����p*
��l�3*
mq����Fh�[���t�h�������ŋ:[�Xv�Xj��D��d���G�53-r:�{f�-w�L��~�h�t�ϺQ�����/�Q[��KHsq*��t�jӫ=����dnn>/���̒�U������S��-��/��|�-Զ��<���|�`�e�RX�]��[V(�z}��R�iG��ve��B�!6�ev�}.�eE�^�LX����"�\t���--����:K��3K��<������3q7/�|XI�T"5����u^�.ow��~b�����*�)�YY�c��8M��l���]8	0����|Q�EF�1�).'��o�����w��ѱ���+���nw�b�\4���Y�]f��T��/���B���}�Yxc�t��{�'��O}<,��ąg�I�!Z~�2-f�3e�u�F�����*\��d��7����d����e�XU:���I���?l�2>�=�}+G�{Z���G/���KOܭgѵc�)���~����z6�g?l����G�ѳ_����y�������r���j�r˚����ͥ���B�$�����w������G��ӧ��33z���ַ����v�{������y��x�[x����J@���>u{*!=y {���O�<��b)��o�������W�������g��$�7_SS���D�~v�SI��Nd����嶗4��DBϿ���As�w�~S���%��	�ì1j$��K�a��v�pJ�R�Qxˏ M��m��Qn�)L4�R�i���6�JJK3���a���(��`;4څ�Ң�F��I�&�`�Hv�T��|=M^�I^���F�ݖ�F�r��e͞�Di��eIQ��F�H��aV$i֐?��xQH|g�^��j�[�Ѱ����I��y��,It���&m=o��A�!SY��`�i{O"��ng�~���(&��N�Lq�
�]���	]�l��eh�A�tY�A?&����Z�WC������V���Q�{�Vk+��?�ti�|8F���r��q>k)�C"Z�����+++���֬��ڜ��MW�Wr	�&h�|ii����&Syي���\�Vo���P���2L@��g���F�,��@cZ�����m����t&"Ʈ3��	��kA�
$m7lZ�7���X���GAJr����&�jv�-�L^�e����n��y�]�������n���De0�������ܜ��ښY'�Bx����ŃvBe��L�)�9%V� �b����D�V���������K�zr]+V�bM��%#���mneNbY�u�X��b��X-S�(�ۑg�e���윶m���7������-($���{�7������D�ЅeB�G1�R���׭p��m�f.b��#�̟��'��+�:j�_���C1�����^�A���p�����}��,��g��M�T{�V�����v)��d#�A�ԯ�F+�&�g<���q��������}�ex�s�r4��ۭ�hϞ=���Р���/��Ū{�ϟ�%����o
������	;2]��w�z�u�{�����o��o9��~A�>�0i
/f�z�m���=��{ｉ��x.�5�p�	����h�>>��_J\�KlOMM%SS��qv��DB[�~�%�h����������]3L���R6��|C]�e��Q�XR�����,�����2c��~+�VZ��YMi(9g$1��Y?�5�ͩV�8BY�sY�cE�tFi���F��9Z��@���N�Ք!\�7d5MBtm�ﷳ,I�a��2�����3�)Kvik4�Gj<iHi#+�Q��p%��6��U�\"4E�oL#�jn4̟<kFf�`�W���oj)�M �#��l���M�h�-�!���Ĳ���#%]n4ZM���5[9�#�Czmu��$>��/qZ�L��F��^��W,��&(�b86ܧ������eY�Z���ж��q����%��2P
��>��J�
6�3��,����Se��q�]�$
c��,�+�N/�^�		�I7���S��A��A�SFf�{'O��u��� �M�"���I�k�ko�+wԎ��]�E�d>	%�w��ږ��9գXnM�q���b�2��Rc�ٴ����Y[hH�*+���'X�Q���Y���K�:4X[Z��=�~̖��B,�b��2���.3T�[���K�T�1Ӊ^^���sS�+�Cش.�VQ��y;�Yrԯ~���·}�Ï�؏[�	��w�w�O~����>:��g�ڷt���6X �,�s���'�G^qUx�G��W_c�ִ����W����+`ӊN(Vd���ea.�>u2��;?�� ���Z��8F2g��C���[�&���?�n�d����?�X=�_��"x�w⽤��fc�m۶�.�]�w�~i�ݻ��c玖,�1�b���T�~-d}_[]��[ػ{����u_�����}qϳ���"�4|qrK(��	)�[��LN���znn.�p��ff&Y^^���ED"��^O��e�Y"{�7�(�,�E�P�z�DZGb�ݞ�PK6�ҫ�\cؐ��|*�a�)����5���a��I�2њv�4���$n˟!M$^����iV�O���L�vai@���I2�Y<.=��,��D+w1,�"-����FSA��6����E֐WI�$�|F�Q�h��� �L�O���?=J�$#�:OFr�)�&Fy���F��,�xC=�KE��Fy��;-�6�C�Hd4O%�ͣ]���TO.��6
wh�xW�g��N�L��9�m��Zn�V;�wM�6��^U4�?׬�E!��R[��+K~�~G�o6��jhA�m�~LAְ �F�w{=�<�z�*��,m��ޏA}QM�W��/��"._Om�JJ��Z�P��xͩ�k�K�xK���#��U������1wo3*�y�cY�c ��P
U/�`ŌJ��R�����=~&0G�qN^sk1��\
T<����`bq����������yY���AVͅ�9�ұ� �����[Au�O},u\����ĜҪv��m��B��ԗ�M+�Q�����L�hbw���L�h�W[1�_L��W�Vۮ	D��=��7���_��ό�`|�?���+��+�yے��S�fyy��S)O�*�������^z�p���a���K/��W��e��
��Y�𷴆�����fg���b�rլ�e�������Z^]1V���K��⢴d����v����=iݵk~�b��5�}f�e�9��i(@[����-[t����ez����[�ϟO=�����ss�z0ݹsWسw��{o�{��t�M�Ợ��"�4@�� `��o^_�r�� ���cǽɃFWY�gf.$�����YI��Q:̥��F���J��n"a.WQY���F����y�dyޒC�D{c4��4key!���Y֐ی�HՎ���yt�ɂ���3-d��"���h�����9��N���.Ƚ�(�NQm	a�3Yċ����V�6�E1jgY#S�Y#k���Ei-�YCޝqA1*F΍"	�"�a��n��._�X������E����n4tN�"�(�߬,�E���F.%�C��E_�I�GA���-�Y��g4*�L*!�6<�hH,G?v3s)��m
�Y.i��Ǣ�%����3k����L:?��JL�}1P�yL�!Dw���K��*�y�]���mk�,:F}ʟY/	fw���}��&�=��D�e�?O��J@�ݚ���,-�(������ܪM��ĸ��������g�tt,�빞/\��>��qc���yc���,����Y��O���`;	Z�^HT�8y�����2!��X��Ñ����F+8x0�Y3\q�	^�:"���t�`P��O<Z�,,]���U��ҫc���U,5F�ې�����I���/�R����Ltm�T�.zM�>+z�����Ȧ0Vi�4���T�;vl...��~?]���6����v-e�������/y��ʵS�{da~��w���ۺ�����߁�}!�@ /m�sp뭷�>�`�u��dv�T���;����\�0���C�-���ES�M٪��Q����������Nw:�N�f�kk+E����F�ΨH�`4T�4[�a�ʲ��e�N������ز|�!i'IҒp�F�BgMY��C�@˙W��a���(�I�����N��6_k}R��{U�L�6���~�f�E_[����huZ�zɵF��̈�V�/��F���ʉ*���ʤ��%��\Z䴚��F���7)����c��C�����;��\37���͚܌n'�!A���e6s�T���(�t�0��h%DJm1��MJ��6�r�_;
��<��.�������]H�>s�����p�}X壿��o��oYnc��J�+��'O��z ;vl7Qy����کhay|�*��Z�W	�+��*�˜�7�� �"?�D�hm� ;73mVj�%7/�|(�E��7f�.˖�b-k��T%�_�w�]e�(+�>C�*���}.�;Yh�fw�����O�puu%]__;s��e�^z�%�>==�SSS���(��Ԃ��E0  @��"0�2dM�u_����ѣG�S�N%r�{r�ېķ��h���5�66�(E�OYȓv�K�B��4Y���a�-���[BG�|a4�
�Y���e����9�*_���&ic�����z�n5���.Q�1�%�+Ko����7�l�|aG�F鋮L2J{���l�j���Q>ZN��B��<�&�p��G������������;[��u_}�QГ ����g?k����[͂}��-��|�e�ܾm����b
1�?���v�5W)�:�3V|�K)Hqx&�hZ��?y��p��y�V�ܻ�k���EA�Y�cA������T��?���T�Ĭ��hi�15��<���Yܦ/x�rb)�
�0�g_���F���K��^wM#I�����+�\�o��g���w���u-?�� x�O��@ ��s���ߞnݺ5ݻ�Br����R@ʃ��;��h�,e��ߞ��yb�ư�]����������O>�R��9|�p���YY���˂`E,�"M�^�CE���!�l�p߶}G���=�|�[���/�ܻ������=���',�,/��ki�$h�2��r%��,�^@GbYrUA�n�5_��(l߶#|�S�����%
�ͬqh<cų2�����<Gt��Y;�y��;�<�///M�޵{Y[?����_�����_�� ���8*  @ ��������{���n��Щӧ�%ac}��w�ގ|vϝ?�n�m�kz����S��b~c�;���۶{b���;w����[P����Z@J��������}����\�"�NO�v��D�W�p[���W�KKLO&嘮O%{�����%�'K[��]׳��@:�&}}�~���.�=S�|����p���e��=�u^��[���~��i���܋������   �$	��������_�8r����_��U�ۻg�e8}���H�_	�X0�JG&_��S�l����հeqф�`X�F��4�ڳ��Y\-G��y���~��)�E�J�zF�f�ҠT~�[g��*�    IDATj��dM�o����\*���������p��3e��{.nc��zvj�I���p�`�W�a~a�iQ�n����?�����w���/�ہ��   @��H������W]��z�C׭����ΝS�B� �VW��U1�H���U��zؽg���]^]5�l	������7�(!W�Ç���W�]��Z^�R����φ�U��lԡ�̻R�Y�X����{�*KJ��Є�$x�_��J%������r��!V'tW��Z��gա��i�V_/PQ�1K���U����|zz:�ۍյ���}�g?�����Cޗ���9A �  �$������o���o����OR�������ť�&t���Ξ=g��JC�������׭8�\c��-[�����0=�<�i��W����L +�Ī���*A���_>fg�Cwc�,m�f��Byn�+K��TS���&d��bK</n�~��;�;.�٫�X��ڜ�/��O�ޤ�߽�]l#�B"*��\�y�7ff���­��z�[���?��[��'_�./�Q�  @ ���n}�?�����oݺ�Q����|J��;�7..-����}��s�,{�
+(���ʊ��X��gf�ov}m�R��:��ewP��ѫ���7}N>���h�Vda-����ga떅���b�˗W�T��$xU2\i┗Y�n�Πlk��EB�_+7=ZŷO�w컱����1K�_�^g� JK�hq�J3��g� �o�2�ڠ��,���)Z�:�N������}�9������xѽ�/�!�  @ x!|��o��[o}��R��;u꤉ə�١�J��W��ٳVnqq�	_���+a����l8�B���&�UiM��
�������*�m~�f5�-`M���O�$�ܱ]%��w�I+c83�kn-C����"�ʠ\�r��O�U�)����󰺺fyx%�%f�Y��[>�`gkW~�zy%>�_���w����V��f�|�����s�������������_�q�R�@�~)��  @ /yoy�W|�[������]�p�� �����K�_�Ғ�W��KKK��V�rO�~ڄ���\.�;��}{������lu���j�ʯz]Pel�hdV�ق�Ҥkk+�����V�|s�`&��>a���� [n��(�3��>�)��h4T�m۷������lY���7T-p�}��n�
v�G�T�^�D"W��d����1����9s͐E��(+m[����H�
ߡK/��k_{�7���/����   @�eE�n�q�Uo����?��|fkž�]�v+�lz��/�*�� �������رc��,ʰc�sc8q�tX��l���|qێ��뇯��׆�ьAl*���1KC�ŋ���T�N��}��y���	W//\ZY�X$Eѐ����t����LMO��K˩�_�,lyu��V�6�[�����^~�,����:���,�Ibnr���~*��Rw���y|ǎ�ǁ=���-��������b��   ��	�y��c�u��~m�H���l�v����,��t�;����ì�L����Ç+����C�n�ݳgw8t���c���ի���!m���7�l���DLG&���'±G6�;�����z�^黛�2��,��(7��<�����ư�pvv������Eq����͚�{��-��t�z���T�����\KץJ	<5�����F����m�ۑ#G��?��O�D�Ab�����4�   �痀������6��_�m����o9w�l��
���E����7�w�u״ґ)PMY��p�5ׄ�����f�ݻ���j��۝�p��W�$m�?�	LY[�/K£�	O=y��|lc���j3�"�,K��n�͏V�W)���ݓ�z����RC�U���W]����;���}���15��;b�}�!x��x�i@ � ^��������־+�^<��n�}!�+���z^�o��q��?/1��Z���뙛��e�5����m
b���a��u�
O�$3WY|'�<Ν=ڭ�X��rk��@�C��m�:V|B�w��zP���Q>�*�U׿����[��|�ϗ~f�/�߄   @�eH@n_��Ow:s;��͡(�>���I��nwv˖��F�ۘ��O�a�ܽrT�L�4�0;;�GE�k���c�nZ�~5�[��<��p�������Rò��,�2�ʏ�)a[�3��6��lҿWAnY�>t�-��ķ��[���pH��SB�~�i �   ��+�:�pfjaa~feem�Ә:�5�WdIv�����<��4�23;�j���VVV:�Q�P���������5Zf��J�5�����1�[䣘w7SڱAh�ZV4BAn�\n��|�%�Ub��[�"�h��y����W>��w����r�/��_=�@ ���H��o�=}��Ls}��f�/O-,l���jLu��Ő���$y����W�$�)w�v{�̿��X&X��f#_��=�"
Z��U*2�+��!��exdo^xB?%��A���)�B8x��Ƕ����}�{�������z�޿+)>@ � �E�(����Dcjj����ص�����<==s��tzf&��VtBb��A?��E��3�m��e1�������������d�xD���[��J_w�u�`˖���w,1H� ����   |���{������ݛ.,-�`��y����r�Z��3(��4����҅��qA>��Ao\B���U�wg0���hI�b����*�ɏ8\w�������<�����/ۡ��  @ x!	|��?7����Ϟ>�}����NMO���ZtI0��,p-���Z�V�W�Wi��%_�~�?.8!��\dٕ�D�����v:����_y蛿������R���R-��   �-�����ei����K�0˲#�vG&�4W��4�;���I�6�4���X����+Q,Q+믂�$j%��RК`�b�=���{�^���ݻ�<p���|�C/Z85����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@���� ��E   IDAT�u@ �   ��	�go^J�a�    IEND�B`�PK
     mdZ�  ��  /   images/b13518ba-21c5-4f60-a735-1d8041d11d7b.png�PNG

   IHDR  �  �   �lC   	pHYs  �  ��+  �MIDATx���	�m�}��}��g��{�M|��$Se;�58��Īb;M�D�#"���v�N�&�ӊr`'�؉I��h�6���7�[���R"QI��||��<�i���k�s/i.,:���Q�;���k��^��   �#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   om�����^��f�m#�  �I�z���'�X+���~����������޼u+�0��mc�6��<�~���~���7~�����_ϊ"�ײ�gk���ol���٬��'�|���[B�  �
��_���֭�'��_o���t>����Ai�6O��㬪�&��\�W�7R���e?kB��7򪪎���h�յ�?��ß���?��z3|Y^  ����3��÷n��=G��?d!�鵽��ˬ,�UQ��~��/��d��8��:�ě�Mo�x�����<o۶ʲ^����,��(&����x���������7ڿ?���"�  |����?Z��;����U������*�z�q��ZM�/�(��i=��Y��]�[P�BUՙ�ۙ}��{=���Q�������e��%^  �ߦ����_<<����B��Ъ(���An��Q�BS/�'c%�\�������g����Z�/ϋ,﩮7􊢲/���~���e��!���oVWV������4���?��K"�  �6����g�I��Bm�����r��i�[�m���c����d��,����&+�V]��U[�i������Mn�lgw�/)���+fs���   �M�鬧����l�x�f^P-��=���IUƐ��zv��k�)��~�Z�f��z���|6��,/  �o��yV7US4e�_��N�k�xo�f_h��w����(­�H���ח�*$K(}8y�V��������?����w~�w��W3|A^  �߬��SO[[[Źs��~��Z�_�{��j�r^ͳ�*��,s���WB^U�n���+vn���7�W��!�?{���Л��vM]��.�f�wX�^��Ex  ���~���W�d�lw688�Q�$7��}�/6O=�6�[��/��h���'�_|Zӈ�f��jl������ܞຩ�����tBl����\�?TM������}�������i4�o5���<�g���  ૞��2�qcp��-6k�hi���7KK�j2���٬͛���;�o=�}�lv�eg���O��;*bț�ݫ�z�כe����ŵ�W��GI�-�N&��l4���J9�g���Tڛ��I���4'���ݪ��S!�/  ���҅���F9m�ނ��ۺ~��ҷ��m�մ�-�֓��e�����6ͥg�����Q1)�v0�NV,�Κ�n4W��djwSIC���r���x�A�7y V�}cϰ���r�DB�zz�5F����+��mz���	^  �U����h��=ɧ���7V���l6����b�r�͎����?8�c+�;�yu����a�w2�~�Eэ�n��ӯ��e�gYӕ��aV��{Ku��泬Q�-GY^�ƶ���e���nz�}��ƃpS���|���/�?���a������~����ֻ�y���t�Ak]������o�u�|p����}4���Ν;���J~|tT-�,[+j����ٶi�)��O���G��۫�������������� ��zO=���p�����������Yx=g_XrU���fVգ��g�����h)+������;��㦗�%�|���R�n>>>��,{(D(��g��d�z�S�͛�߰�:��h�ݽs'[__˪6��ka;+����`=�ا0����j�ťKK�d2��~问}���2�&�Q^�����������������?���]���d*���������|X@A����V!7;::�,���Y;h�4�hgw�Y�X���[ߡ!���5'��KK���Q��<�=�ю��μ��t���qc0|�v���yu��w�굳g7�E�]U��+�i�=���eo2  ����|$?�^yxm��3�#��Ł�a���8Wa�J���PU(�1�KK�����zV5[B�ܡ���d�[8��1ΖF�L�������y�Ӫ^[������R������WYD%3�^ӫ���-om���g7S�qv����|ns���������7��n�������|4���5��᰹y�f�՜I޲�Ww=������ǳ�<�̿���;;��~�e���U=����0{lavTE�_�rn�B��<�u�x����o�7�픃�0����7�m��;�ͼ����{zt�է���}t|��{���+n�f�Zb�֒{B;�Zj֚S�nf�i�!
�O������w>�?{���,�fmu����W�.]��F���2���=*��~Y�>s���t2}՚�;�^{+���v������?�Co���G���|Ŏ������-�׍s��(p׿y������ �Uɮ����K��z��n�X]]����Umn����a~<g��;�p0���72��f�o���e�̮���77�fw������t��-#e���m����3�̠̠���x�^��/�ij\.b@+B[x�p�����:W��`0X�498<x��>���[h�S�ᰜy]�L/��n�����ן�f���W��=�y��f(�+p�c�Gu��?����_�/~%+zW���گ���?����
���_��}����Ɲ;w>�5�K��G� �l������Z;�3gΔ�q&�
h�.--��յ��T�«����V�d2����t_�gZ��s��l'k�ժ��$�Cm��N��d�^�\E�����~�M�w��W��oŶ��lln4v���Z�y���奕\j�TV�uo�w���R���}�\][Y�Lf�kCA^�~ǖ�YYY�4)I���>j�{u|���vs; ���+���|}^ǉ�u �k~��U��wfٷ|�F��o��������r��g�Ｕ�8� h4$s||�����sc[/;��t۶ǡ�B��|�(�;�|;���֠_nU��`0(�Ӊ���F���͢>:ڷͳ�\��yW�T7n�h�\��~���m���w/�G?�TK  �Y���w�,���eQ�X�X�'��ں]iu9-<SL&�ll�T�Ӫ@����׽�=��욮lyw�N����=����:��gh�#��J�_��g[��5���RM�{���@��!4�5����$�-�F��|f�?���eZ^�"������^�>V���������G���+������~��o�r�Fѿ�����ǰ���S��~������=�ؿ���W������/��W5��'h4�;[����S?rtx��1��
�]--/����}����m��6��VWV^UF����ª6�?�ZS�h�hXB�p�Zm�����ڛ7ox�T�nU�=���j�PJ_k��k�hH#WX�ίC��󐫲��`�߼y�_K���F?�@�{ܾ}�T��}���p���̛�4���>G?����M�[��,[8��ݾ>�5$b�QP��������8�?��t����W�ּ�9ф�^�W�W����U�3��|���,��6�Ѱ|��K���K��Ȟ�yĥ�b��`��]����l2�����F����ʹ]��a}V
��x����^���\˥u�����}�Y���
���+�-�Ϧ3��j8�5�8���:i�Ț8a�ƙ3�5`*�3k�Nl�ۊ�����ʲ��n�g�O�����R�{�r�k'�{�Y1����,��vЯ�㶱�^O���Z�\����hu���[i76v��͵v{��OP �����|d�����G~��۷�N���e���{[�w�据�*��u֯+���]��:�+�Z����]��>�E���;�߱���?OZSX�(U��/��<罯*wPi�����j��2�84���k��B���v�]V]��}/�pup�k
嚦�~����C�����V�]}]��������Q�E��X��4gp�k���v��C���ã��3��J���<}�����\���O����y��?���S��o?�C�+�C�n2i����|����F�@͙�3�ŋ�K�.U�Ԛ�3u׫��6�m�VϓVYCi[9����L��;;���ʒG��\;H�`����]�T@�Nt��h����Y�����zB*s0���gtwwW=���;;;�B�\�v��p��x�k���
h����C����*���Y;0tz�܂�����F��i,
�^/��@��kGU�����`�֚'H���k}�Ν|�B��>[G�Ϝ=�ˡ`�K=��/ߧ!�|پ�ϧ �kk�������Sdt#���¿
�=��z��6Z��g�u�v���z�ɵ<
졆����=�s��]k%?`���sv����j.U��L�c}�R��`�@�7j�2��<=���.ʰKס��N8�\�g�`�l]'�<����`0��e�G���@R�I�!�o��m���������>_9��`��U������s�e������F"b+=<QGډ����!�g>yx�����NB3[�֖�f9(��ر��=;�G���|��k��5�����e1<��I3,g��R5NڪZ�ٲzy��S/�G�q�������j{ܠ	��SO}[���_l<a�,��S---��AL��޽��2A����E�f���k�%&���� g�����<�ݹ}ǯ���|d״��N��K��9ш���ƙuz�wKu�Z�!�4qF�N�3��[U���m�>���`>�t-*u��=�N=����da�v]�N{�e��"�&�e������&��=�vͶ$��/�K�o��'�}�G�ҳD��^����??x�\��eǫܾt�^u�?���?=�Gkk����zr$�o��o�X �l8�2���zGU��e ��-���V�a�S��A��]�����*�Τk���_~��L��
R����B�Zg�A�a����0�]�ND߳X�֭��0�H�'}O;�>�!����I���r'a'�eP�;�?Ph*�8�^z�=������X_W�To��n;z��R��}?$�,[��(��k���^%���F��}��K�E3��o�;��Z`��n����u�C7���f�jh
��E=�
�)@��˗}�=�&�{�%�@[��D�i��R��Myhi�g��^��w���ݬ�y� l�:M��tOu|�����˯�@�F���Nj
�
�z?��n�����C;��$�Z^� l���9�󕕕j6�ض��ZFՖ�a4��}��z����~Zμ��^��*G�5�����f`�W�Jhp�g���h�{��m����=��^[-p�R��o/ڄ�L���_���g,������}v�zٿ��wf�K5;�~���	N-
�e@^*����Vi��7F��c�KCv�f����9��a�m~�6�~�k�{�5w�^{�~u�a���~�[�o&֒�l#�hTU��ܚ�ڰ���a]j�<�loo���Gk[&�@ڭ?���zO<��/q���nj�V��ƍ�����u��n���3�@�åAs����u��n���Z�S�O!uem-�X��D]�Bn��묮g77��x����]쭏f��A뽬z��ŋ��۷ny�,�گE����5�����zO�O�m�kr����놏~߻{����/�>#yu���K].�Ƕ��pWGX�#©��Թ�^���,u)�������{~V&Q����fŲ�'��w��?�goa�c�7<z������]�z�+��ї�������>d[j��C����=���{��^�x��֑zG�m�S�_��Q�廟x�Y���jc�Li�sptx��d��F'�tjV� ��"s������]�
C��rM���7|Y��^[{]L=|+ .�F]]]�҅���Ǟ�\|����{Ҵs(��z�L���<��*kM���li�d�i��v PY��·|��>{yjv	m�M����ܢ�[�u�U�hZD�յ��a�k�c8Uֲ�T����g��k�(��u���~'�zC]o��4��;	xT��J6��p�<��f˰���TC��Zh�ȧ^S��������I#O!6,˒�Nx]T]�<��'>�P��O���V^����(�$��캣6���u!��R�]om��t潣��k��^ʢ�W/�zx�84塾V�x}����C�I㦊�a;.���^�]���>0�����s��A��N�<՘�9�xJ'E�(`����5=[1�K���ė�i�x/��[�;�1dǓ���dg�N?~z=���!Z��A����9􂍖�ΝG*=��X��h��sȢQ��|ړe?�>��n.=�/�uh,�2"���_���7~��Q�n�O4z��1�ʇ�>ի�QjD�+���5�T�f�����S0W-�혽#;0���C���-ˁm�[����+k;�Gv��7yy�ֵ]Aډ��qoП�2u ���Zi�~V��Ю��6j���NG��p�N�#}�fi��V^c��jk�Y[�/�9�\�5�/�hϞ�i�Od�<��/<�{=������+��ͭſ��m�[+C�>��p2Q�'�A�l��(;����l�7�G�����Vϛ���k�<����ʪ~�X&�7�~�o{�:7>��������Ǜ�l����ύf�v:��G����ht���~��X��pҋ�-��h���p6��ً?�u��N��`6��{����?[���Sf�|� }��>��n�\�ˑ}�}�A;��b��I�ŗ�d���������x��Zí�z����hmۨ$���~mڶ����rQ.���ӷs���Å���j6��&���Q~�Ν�������U��6�p7�s�nJ��;�~�[_���^}]�eG�@������B�v���]�����|��9s6{���|�j�������ݺIDm�vm�lvəL��S�׫/h�s����ڮ�S�R��������>��x��"L8����c/��K��E#���d:�k|虾sw+{���s�������}zx�c���{޾tns4<>�ٰ����_�C���;,��-�>����c�|,;�|~�����^���4̬�������{��M!:5�E6�����A���w_So�BV������ܹ���x�h'�x��B��4��;/����[���u�V~���|��f�;2��~��������W_������e��m�.8���
��S�������=�+��@��]�5��z��c�a��\=��bn�Ƣ�>Q��Ϫl���S!H�A�⁨��X⯧��%�ݖE� �4�љQ��/˼5�P�����5T���3)+P�US��H���=���4���e�<-��q�׿��O�iOX��
�)��=X��逬Ю�S5Tt�����i�S`����i��ZFՆ�v��P=�gϞ�bi�Fr�?!ؗ^+��p���S�J�6�u�co!�~3�����Z�:�����"LK�]�^ �稆��2��y��We
�ڟ�?��F�C�Z�J�!�嫞�ڷ�\w�wz�PH��^S�[ˣ�t����Ν[�?Z�0�I�ˢ��5�-U���w��i����8P��֥:����M�N�~����'��¾����kT>��z�QZOZz���ԃ?����qR�+������,)��i<ݐҺM_�>�I���t��Ok|g�����wSǹ���⢥�'�R���p���7��gZ���(��k
��?�T8g|��S%Q^w��֫�le�f�sϏ�&\<_k��4�G��8<��Tk�㣱̮2+���C���lZ�hZ;i�u��m�FC���X�J��X��f�5\������E�����Vu�m��]4��� ��7+zŴ�TX��	4o���IQՅ-�h0��~����m�ׅ�O��DY��U~��l�h������lP���t�����>泽�-��R��
{�fسw��jM�YQ���O{sk�i�򺢢�E��X��W��04����h�Q6�-�,��iE�0U6�-��zM3�UYU̧����Ӄ��W�Zc��G���p�{VG�dz<:��e���j�.�k3=�`e8��{��[�ɏ}�G���U��ٱ1��u��'[�v���hǃ5��z2k�̦7��q�Z��Rê��6���6�O֨�k��Փ���onY�>w��M���n$֟q��N짞���������_k����^�u�kUϩ�q��V�����Pݨ��o��M?oZv��aP��t�޶�c�Zh�{�nv��,��
������<��*?��`�e
�:����xٮ�:g��E_ޢ���Mm�x�E�z���}��z\7Ξ�nߺ�Y���x�UU�!�|3�΁�,�|�M;�Z��;��5][ԃ��8{�Wl]ݭ����[؛x5݇������+�����[�ް����ի�߱���M�����������wd�{{����ZX~�v�#�����ga�|e�/��[�HK��:���Tb~���1}��,�>`�R��h��T���Y�'�.6?�?�kR镕����������677K]ptq��������vqU�TX�0H�M7j����S����Р���̃��o
M�����Gٚ-�BT�I.L`��TI���g?�Y�W�/^�ϧr�Tޡ�l��B�&<�PaU?S�d�u�����{�z�=oZF��omoś��x�����3-�NZ
�
���!7M����&-��kZ���4��'I=�
�!��_W7;�eW����b�ƻi�$�ƞY}O�@a��'?���z�0%]�_ײ�w��Z/��C��ֳnrX���~�����k4����������P>��׋�/��AK��Z�z_��<��%۞��b�y�D��7x/���?��;K��!�R���*_'MzPx�Ի�&AW �6PcR�e<����Zư���XU�ƕ�᳅�ƍ����.i�FL��"9�7s�O����ÁOѣJ�~1Q�@���s}�.6�Imw,[񩆴�n(��z�t�֍��M$a��d��QjP�z��ު/��'�6�dFǺ7�bX�bϏ���+)dO|_������Ko��Q�آϛ�#�2���S/`i�0,�2z�U��������N�q&[�����u2_K:6��X��r���~F����#D�0к�s\܆���:7��L�Pu��F��ױ�-��3m�,�M�S��7\�9)��d/�-��tПv������>�dYx�)T����y�r;���Ըj�6T)���C����׫����M�&S�J߮{����as�������(�y8����U�3�FeQ�m�͛��p4·j��m}��W��GiT��.�Ւ]!�H�땦Z�W����h6(f����}֨��<p.��T~6�k?��+?77����%��R�u*��x�-Ν~ޝ�f��Tg�:�����sQ���S������Jĩ��t���ʶ��>�ܶ��ř�a�Y�)W�M3�Mgc;O�'��ض˼�+&���^�e�l�_���z�/�ǣ�5(ʢ���{��Y�������ѽ��?��O���e{�Q]����w�����.zCUYD��>��Ғ��};g�!��\���S.\��y����^��5��k�^����ϛ��s�ƞc�{�pX��g����Fo���y$^=���o�G�y3���^�L޳����ɾ�unq_��o�-�[�����7*���5��|ue��r�w|�������OngoAoj�|�r��ϖv�>��s/<q�?���w?p������)Xz��s�=��d�Чq��i��6��mٙ���ÃR?��N�
mv�kbU�`��;MLG� �a؞����d�Q�a��]���	�NB�:
�*�Po�B�vv�"hH[?�״ךF��J.�Ë�K�`j���Ԕ"^�z��������=�-����(������P��=�}�%�:�ؓ��)���7̾�B���O�vN�y�M�EP�8�R�n
�
C�����S�{��K�hi[�$�C�v�N��Zn]L��T��?u1�����n�e$C[�TG
@Z}ch�xAN��0uJX~}�<����Sϥߐfj�*�{*O�.볅p£�h��!M��7��xE3Fh�J����z+���*�IR�E�JU!P�YW���S��^�>�k_��r�n�X#�ϥ}Oˣ��'>�Ҷ���G����}ݶ���Xʱ�lZ�cR�zZ��� ����x��:}b�:LA.�:���C����ɔ�:٧}�P�<�}�R��|�>=N\Z.�ꩌ���v�´�8�[�z�f*9]Ýz����}(�ظX&���y�k�}R=4�N���X��+K
���I7���9��,��./��xcdK==�KqtF�S*��c!��7.�K��^�D����s���-6�I�%Yz�:��X^�b�o�f�^D��,����Ư��zzuG�F���ì)�b�$s%���^˩�;�}�º������b��m�v��Ξ�����֫�R��w� o,��[��*��B�.b�Ow�k�N����t.��~�T�Mׂ,��~Vewڷ�N|�2�1��l�:bA�K�4�����`����:ɨ�>���j�������u���f�I3�����a*�C*J��d�=U������c�k�����,Ko��q��U��a��x`�U������Mq5���;��^��]�x!�Y��ͫ^�wo{�;kf��I8�z�Y�O*k�WN��F�:����Ѡ���M��,�_g�č���`8���P _]9�8ZZ���Uu�W>\�����ny���gׯ��]�t�υZ���\��G���%+���צ8���F�λ>JcǺ��Օ5o��u^ZU�({��>b�O��l:	�A�á���h�%\�EG���(�k�2�*�;;�'-���k��H�����~Ly�U�V��LI���|�C����õ��?e>���/ފu�oj�={�_7�?�����~��X-��W^�[��+WF�����I;س�=��b���������^}�U�@���Z,־������v TK�`k�jԍ7
ӈ����
m:�h����NT^{p��'Le�9�d����ð�@�)mj��F��ի�� �_��_�/�wIAp����on߾�ꤳ���l��<�
,�f��p���^�u���{T��.��,$[8V/oO"�㐲z�ԛ���iBv,��$�n���t���l}^����B��G������^�rٗMR�j(�X
u���+�� R���3g������X�����&�=(:3���P��4oy�3�G'f
�j��B^����Z�\�ԯ�z�x������FL�M�O4ڏ���룿� ������w�?�������Б���O�Q��C�V�b������GK�<�k��'�T^����E�~Fvq'l&���z�N�k�nݺ���Cxn����~��/o�Xd�E����^�12�]id$� �3MMW��8,��o�0�=*S	ʪי��>��O���X��آ|�,A�?g���m�!�67N��_����;�&�Tc�?���-4����,�t�JB ���I'j/�-zHO.��B��h0��JJ���F����:�<.w��zī���˗z�㴈Y
{��)���n�u��E� �2W��y<���������a��b1�H��K%L~��p���4��k�}|6��)��eѺ�q���T���ŹK�����0b���c���˴��频2����/\�ؤR��˫�]�p���:I���oW�#PM8g�͘޹1�&�w�Ӻ	�V�aw�O´�E#�v��U�S��Q���Sǂ~���<�@���.��E��okk����M�/4��?R��W�d�̦�ڰs���/\���l{�:Q��^O����ԍ���;NoiT�,�Y��̏���}�d<�o��g%��j�	K��O��_�z�l�-Νj�k�L������fב�xcVQ�#�;l�u��u���z�y�JSs�/a_׺����Y��GZ��Ml����"�~�4��api���i2����ꩴk�N25�l����gWy��Q��&3?G�q���0����p�ѳ�׿w�xo��0��s��ѵ�	�65켬�U몪C��v�����������c6fH�����5�pi�/J�|�N!�z�eo�4H��^��zx��.t�y��c#,���s�=?�iƲ�虧���7��~�/��_����h���>��3ӷʃ)����䓟���ő�����|���M���ֿ����y��K٧?���I����e��~��ϫ��o��ڥP�Y^8w^;V�D�"�^�Z� ��cvrZդ�
=vQ�4��.�z�ّ��y��FAHñꎿq��~+_�Bq�����P�·n�Ց���5�t�bx^ʃz�;==������A�N�]x��<$y}�}���yo���*��^z�j��w��B�-k�=p*�*d|�3�Y\���w�ν������|���}����2��L��؂��Q�Z=�['f���-2.��^/��Y�լ^�F� ꤥe�t+��b8�O�#��7��sj��� �gv4�3]�p��r�pL�'�xh�r1�ً3>�Z�";o�]aL'B�z����t�J!��g�3:��*F�?�s/��.��t�K��ԷeхFu��	9Wl�$�Y.�K����RxJ�o��ç����׼�A�������!�pTOp�e3<h�`ɾ��g>��VￖA_W��BR
���F�P�P_�q���<��t1�{�����m��c-C(�Q���_Lg��n����~�>�,4'=�����l��3�Ts߯�p���4�3-�.�jx�ѕ0u��{���=�E�C׋��`��K@�����|��=?��m��c3��bq:��^BzG}��8cI*Yx�>$�~����I�j*�H=�u� �=���i���Ϟҏ�w�X����R�tSlz�r}�E���
q^��=Qy~�?����S$*X�a��T��4����Ǜ{�h�s�=��T���|
}�~��Ҕ��g��pt����w�Zibi�OU�כ{-c��=�&�fִ��I�V�M���Z���k<�s�]�
f�Hh��-�f؎t2�ci���j�_ͨ��kD�=��o�/����E��⥋�vwv�5uD�>O���J�q����l:��Ԩ�yR��m˘�ȕy��`uQ���d7.{��ꈽV(��4�̭x]�����!���5�u}Ӄ�,�g��G^�����+޸�y߽�UǛ��>K�ܷ�,\�.}��롞�����SE�횽`4�ٹ��������7G:w���F#���/���r���k{gVJ��f8��`׆�����ً3	���06d{�8�T��A�Щ��R�F*����m;Cb	�ɱ~rJ�
���rx�p�_�z��{VD��p�iHei���ק�e_���ܧt�3�}��;:U����-Cͮ_�~fk�����~Ys�?������ޮ]o��S��-���c�Go~�����a�#7�ي��ȏ��o�����|�{�����~�����r����	Uh�<������?����}eeէ��2\�'v ���,-[эB�]��l�W�����g��qc�ñz��*��_{�5�F3.�e<�)�gO��	���l�+u����������K4w�nXe��'�L�a�U��"��vB�3l���VQнs��7����D��"p������&����ʕ+ޣ��jY=p�ƺ����P���~�EH���u�ࠡ���ʕ�f~!TN7�h��6R]�JO��/�^�>K�Գ�^j���>������	7ˇz���.���^��[��Q,IH�d�*gi���$݀wzhT�A�vP`T�������FF�6&�&�����Zq�:秧��z߲��^�k���C7���}��M�}W�j�ÂZw�X������������v=�j�脪m������?�r���'�𰩐���ը��_�{��|t�(C��5�vo�K���k�w|�wf��ԧ|��τ*���|U�<��:�ҷǁ-����X&���򗁇�����׋"�i��,�b���i'��*,��������2z��wn�2hY}z��Q�-b��A1����.zX�8$�����4|���p�Hurm,MHe�ϰ_Ws�	��o��A
ۗ��O�/��7��S?�z@��Y���`�u7n��r�´��!4��+�����kR�a���e���4�P
ӄ׉=�gR(^T@�龃8CJ8O�Q�S��xc_��s��M=�>:�@��ZE�(5H�݃��h�F����'.f�y��hAZ���L���=�鳝�?R������Ϝz�&���|��\S�h�3��59��O�a(�����5�n;�>w�\������������^X�[�}-�X��q��~7��xՊ}�p�I��q��Z�"�J���z�z�LGz���G@|��ҬG�S����z�0R5H�:���uGjB�sii�ܵk���Y����4�Nh���;/j���P��_�p1��qM*�Pǆz��������zGr�P����a��뭪j�����凉5P��>^V]�j����S�p�mm�񹺺�S�.����,N�Y�V�Zeuޤ�����554�c9R�ao�ޢ� ��P/�OE\g:/dm�q�"���{:�∠OY��|����ݿ����>�n�/n�tՁ���'�I���,�L�*�X��,����ܡi5Ká��h����:���7������?Q)w�=s���������G��}�7��Doz�m}nƏ�}�W���~���!��������T��=Ԇo4�9�0�؅m�\�@��ӆ�?�`�mۑ|m���O�����?���_nYtݍ76�j����o�1[�o�s�ӟ��B�O�a���`��RM���6�,����*�ܠ�����3)��K��K#�D�p*�A��f�~
G�~�L�a�j�����`w7���Uk/����x���ih�[�
H
��_{�C��O?���"�}��E��իW��vҁ���2�J{�$���e�^�س���V�~fgw'�\�'b��zb�5���B�.n�q&�4��!�4���~#K��N��>���u���ށӼ��Y�C��j�o�����x��dšv��?��gRo�/_�����c�z35|�ى/����Uk0�f�{[۱qΗU�&��u��K�M)k��'΅Ϫ@�j��Y�l�xhR�Nd���>ָ~<�춳��
�j�h���mg}F�tՇ���Ϸ���������~�Cpy�ԍ�M(�2��.�v�[��������l�{����	�a�C���,5:���Lge�Sc�Kl�j?W�O�A�]�z���q�muˀ�}Ɗ�E�b�/zC�,	U�����J_K�P?��rS�9�3����5>�|����tꦴ�,3�4"�P��YM(og�p\�a.C��h}{�y�/.,��gQ����c8�}���X����4A
Ⱦn�U޷sk*7й������Zg��4�C�}/�Cݡ�����9�{qyb@nJ@Ky����|5�Z�x�T��9γP����ң���K�TF�3��ЋJP�y*�ᓐ{�(Ќ�G_�Gקra[N��Z�
�i"��$�4�����W���9�O-K�<i$���ף�<��4�}Ҳ�O���у�⾘k=����NN��^���WG�-�p4����`�e�-�g��<=�Yy�*N�XW��k���j����+xC|3O��׍83�bV#}v����h�^K���E�S�c]'t��2�U�����qM�fi��u��Z�\YZUO�ȇ�/��Ӎ�>\7��w�F��5��7Z�䲋�/�yH�#���R�'�x����C�fo��:m�E�z������]�[��R��A��A��2�"��)�z�/�Eqj��GC���5+ܯoN�ſi�*n����=
~3o�d
N9i*�C�_�5��]޻w��lZC�o�.G��e�E��j�R�ؚ�W���ε�v����Gٛ�+x��������s�,;�������}���?����{����6w�wsk}����
a�5�B����co�?�ܳ�|i��5�5�c����v6Z=c;�߱�',����0֑ܳ�~!����[����(ֶ���ۆ~�.�8:8z������Ajg�l���@7����Oeѝ����'�t'��Q�eRo�����&�p�V�p�=��$���n�X�Z���}�{��:9�"�C�
7�9�ހ���z��\:j�_e$zʚN��fUua�,��߱���I�xN-�B�[�8N����G7��	���Ah�ۅQ!k�J1K��i�R���xײk}�b���,����~|�Z�D=�a�ǞA]$��6�LH:�O�g5$���f�:�?�֝�N�YR�`?>�yb'���O�##�;�y���t���UϹ_��w4#���W����?�����y�k׮�6���_�p��n�)h�E�X�Z�:�Ʃ��������K//jm�}��>��؋��*�Ϸ�h���𶎴}`�yE�OAZ_�y��"��k:��=��P�H�[�8N���R{�d�7��{�E��rORR@��>�������_|�?tv�Y���,(��~{33�%](�$o���z�:��=��n6I�e��Lә� �z���)���>N�A���\K{�5c(ܲ��+B�.O����S�ԥeN�M?5�N��Ƀa3rě�⍘�7@�ϖ~�V�4L�T|��7��M#X�҂<�P7�S֧fr�O�Զ��K�4Yq�C��������>O�/ͪ#xT���,_��'��T[��C��5�?�����e~��{����>_�nu�}?N�φ�ºN�Bi*¸��?_o:��=���p��#�c)Zӆ^>�Vp<^�ӝ��mo˿��ɍk�Ҩ���_��ë��ڷ����~|죊a��8c��w��i�K/�^l�?�dȽ��_.�}P"M'Z���F;��7͢�(��сT�i��;��>��:DO��9�gc�Ǘ��y�]3,5*yШl]Hӈ���z�h����/�����|({��+a۝*�K7��c;���i(c��ڥ�@�y��W�˛t�kR�R�q���ٺ/��TB���E�|c��j�ziQ�U����<Ue���6���+���"�T��#z�mg0ibGђ�����*Ubf׿fue�{Օ�V�W�V�J��k�����7�ƙ3��.ՙq����or��ޏ��ŋ/>���^�����m�ǋ����x��t6_y�w�~��G�o㓺x��kʦ?6?r�T9�.�ڡ~��{s������^�oݼ�Cۡ�/��/=x��?������M�8�w��������>��[�������n��d,�fG�M3�P����d�����v�<6���Ps�.ښ=}t��]��T�g��q���"�y�t(�̠Q��h���4����ׯg�iX������0�n:Jw�~zY2��.�:�]����$�rx�}O@���v)��O\�w=��+�t=M�[�k��O����Y�LS�LgS�S}������'�&�/�v�j�8���T{�S���9#�g��Q��eA�M��3�%~�p5����lt�F��EXW���*9� mM��j��6�Xc�;j[g:�鳫�F����ۗe>���#�� ��w��i��i�ܯ�k��y8<0���c]����=�y��w)ܕ����'̉��I��q��t��͍z��0�����я����O��=�xͨ�m�7S�k��.L������y��G�%�	�7�~zXI�?��N�8��=z^FT��S}M=����iĬ���@U�i��>ǵE�~��:�����=����pmxl�����&4:�z���
�!�����|رi7�itf%ֶ���cT�S=���{�^��x�b�:N�;֠���)H���ѣm�3,�^��ӽih5�ϼ������E��Eu��A]�4�v
G^�Tᩄ�t"�w��".��J_�<_�y���5�>�2�(k��IH��P�J���T!=-�d�����5�8O���+��Ѣ�$�<��W�MC����z�oh?Uc6�]��[,ch���NǺע�0�|qæ���m^/�A���&3��5��\���m�q���� ��X���Fc�Z6�W��C�چ�75�2<;��Ž)�<��G1 �M��.� v2�LQ��ԙ�$��r���X�s���<�h�)�)0i]�b�Yz�����G#gi&���5&�z�����T�WqE�K��e<��X{�������T�f0	3�.�K�(�+��G��]��ty�z��Nu��k��
]>�X��J8�S=��>����9�#�?�i�w�t�ZwGǇ>z��a�L��8O�(����f�qX��X��s����<ͦq���]t�f��ͼZ������0�r�6�ꉍ��$<��/V���c6��//�(boq/K�C�s?��|9Z��ry��m��M�]}���=�?��зյ��iT2<�`���|d������7}߯H��{�'�_���?`;�v��g�LU����l�޽m�iF#�^�������T�r�����_�������������p�m���g>�3
��p8ؾx��g677�l]�/���5��K�|�I]������W�u�褅��[[[�wxttk��[�W��~��j�1o��֒:?W�u[��Dtv6��_5��u;���oG�f֎Sv�|�.TM�]�K����-�X�(U��'�褭�����of���N��¥f��k�U�_������^�S����u;����/����&����`�T릇�4��y^���i��b���x\��G���4_f�}��{��������X��3u����p"�g'���:��p�+��]��G~a]ZY��>�oo��i7�ז�~,޼h����Lei(=�(�Z�<x��-�I�5��4Zjz�����BO8���}�s=���T?���O���2��u���ڜ=s&WӉKӔ��['�]�z��ᑇ�6>�lo��C4M�Bp��M���M;�o�Os�څ�. �d��4�K�����z��N� ji����q:�0r2YLI��LAV�5a���������
�?��0�F�Z�i��zKfވI� u|��8�z���>����v�0s����Z�aj�P��!i����� za=��Ƃ��nj�ǯ��c9�Ɩ9�$�@?�!?I�G��i��R-������x(�Q'=�1>v[�'�N��W)�����H�L�������n�Ұy����j�/�ZOa֚c�)<�z���	��r��R/a�=5�Ҕw�O�i��<�_U�Ǜh�0k�b�t�����Yf��<�Sk:.�?+h��~�È��Ã\TG굚�}������}�Nx�Of�9BC���������4��0�@��F��p�r,'�73k6��;6��z�4B5�fa�����"L���W�x܄2�����l���\�;�1͋PJ��~SW�1�z8}�U��*uO�}JSօ0\���|݌,���^w��H�lј\^.c����W�Q#n��řw¬0����E�|
���J'���1�*��qs��㾌��fu��7���8E���7�@Ϯ�[���p�\����9{��}����p�"�i],��4�G{��7���ł��{��L���N��i�[����ec;�i���{���Y�㩝W���wըn��w�W$�N��7O����[��*��:ǫ~R]�z5�76*��~������S�h]]�
 ?��~2�ƫ��s���/��ľ}�~࣭��AܟxS�e�?�{�f�_���3�.��������N�v���R�4˳^�ԫ�%���|�-�����;F4�rɂ�Y;�k=^��|:#;I��gRǓ��(8ߤ�n�y(�b�!r�7��ԓ�z|��Z�:ع�PQ�H�S��YMOǉ�!>�z��O?�XA^�_�~N_��B�=�i�m=�U�r��Z����h��YY[���4g���X�^X`,tr�3a����·>R��*��kě2�8�Yx2X��-�"ΙY�i��~a�J�c��TU�Qp��$D�gni��fP�k*&��$���AM�wY7E�gS��w��w����u]� �O�K-�z�Ğ��?��\ܬ�j��v�T�&H
����B�����wa��T�aL(5>��PW'Sť'���>O?d!�P�BT�6,]�ROc�b,M�������M=��җ�����O���0�9iz�4[F�S;�����S��y���,�\��
��{ol�u�	�Ϲ�o����T�R�ed�m�8�1�M1V��h���p��A��?:��#��+���S`A��*
n(O�O��Yʔrz���;�a�^�Z{�{^�6`)�vq��~������[k}�[Pq�c3V����j@�ʼU��)�}����~�6����U�	g99�¡M����<i8���2{�q|�Ț7^ x5�TC�]1�J�Z��J��Q�ٲ�b�`X��F�~_�)������)7@Pˁk!����W�f���֊�/�}�~U�7���0P�Ds�ה9�[�f-..p 	X<����R|�ڞ*q4s��pf�	1�:x�G� 4�xv��]&��!����mܧޯ��80�5� �h�U�g��'́��y���e;O�Q[���*��yJ)�R|!Q��R%8�34�N�h��	�؋�T�-�xn����&"O���%SiN�89Wrڕ�Z}��Ca���8.�\�����V�&T�G���=H�2fRWZ���"1�%�%P��W(ϗ$�c_t�!�ײ�,���I<8��'f�ֈ�����s��Q�.��K^����9������׆�7I�=�w&_����y��uF���L)@~��Qs�˿�y��_�ܳ�xP}�?ŋ��ܜ[Y]�w'K�^��U]��k�"}@F�+m ��z׻�y�q�T.._��n��[��X��o'�h���آ��Y����;�^_���M�y�봉���:GR��Y��~# +Z	L6��bm��@�c/;�@�W{�L�#
δ�P���mӵ�;�ori\�p�*[*-լ_�O�sJ�u�zI8�}�ɨW��p='�Ђ�j>�%��%�[���$S�
&|�z�V ���>��"*lkvs���f�͘����1J2�3,/-��+,ZK��t�\ ",��q8��v4����B#Z�W=����lxNP�7�c�kA�/�V�҂8���)WM�	�0�l���ޮQ��PN����E�*U���Rx9����I
����$!iF2��y����z�-��qQo���c�
_)�7N��w/^�Xr�q�zp�<��S=�
\5��EK�Q���^�7����=P��h��*�@�� ��Ӱ��2�z��>O@����ڔ_�Y�xx6U�k}f6�cƱVyse�7�<sMfU�]U��rQ�QC�")7�V��R&�����PVVy�{{ݒ6���}5�f�(��V3I.1<YH^��oD��ŋ����{���~�O?uV�\�'���H2>뵰1��D{\��dH�E����H:E�1 t�6�g���~i��!N�uK1'��H�e�~����$&{~�xMlDӪ�p����J
*�x���.��3K�M���ø�{�`��Z6�d fHN��8�X��aH�(���;5��'N��H �ن\��/<��P_"�=�0���4[IA�4�W/릆0{��W1UϬx��F����5\Z�Z� 	�(�?��=��P�]��RM�?�� y�)�o�M7'�6��3�����K�X� E����>��瀤gx������S��U+7<z��/sw�=�ȱq�:(cZ�{i��D;/�M9�䄍�̙3 �0�����ş�&�a�fD`��4���N��z�w���A�UX�cڞ��s�>��D��\Q�6�0>pdm�Vwas��4/:�w�Y�������px����8���6�$�F��]�E�C�+@�hH�����h`�D����n����]C�܋(P7�e̘��Qšm�*N"�����3�"�b����ӵBV���A�t;�!mqin����k��H{67?9k�� �ܺƋm��yjX��e�
�W�.���no�y�,��ڹ����>�hU
��Z�,j��i	�xS����hcɳ	O3��V:A� �S��z�8�륅XU�M��G��X��V[�=�5M�2h4^�K�
�|H���~?�<R�0/����qQ�׌M{qe��r��Z�s�9�
x5��@T�'�'�K}�Oi U`�T6Q��@�ЄD}��1��Q8)$����+h��Ӫ�A�

J�p\���{vRr�(�CP�����\�v[��Ā��}K�G<|�m��u��e�(rB8�D �/�T��}"�1��+c�G(�������<��~��kA�/�zww��8 � ��c�vm�s�����m���R&�i�$4��5/�F _x�1O�|B�ի���D����]dp	�ױ��q�x�ɲ��5m ��$j8I��0����A��y��x���uդR�A,����zr�l�������3A]������b�&�ӧO��	����F��u@��U�ڒ�¼w_H?�5S�����M��,�_$����_��z��Z"�@���}!�\�N��{�����|�ڿ_�^���R�W��R6~yV����؀���*s��V���Κ�H���ws�w��ǡ�UN���-����Q�U��}�{�S��8{/M�������&�]��h@�a���Ewms�';����>��rg��A�n�:
�I�ץԞk��fڦ��|"��P]?4x��S�������	� ��׮��^�����L=������ţQvSa�L���(IeY���9������~M��A�D>7Q:b���O?����d:t�l3mj���O@�����yD�r2�C�UȢ�\g~ց���ȱQ�H�q�Z�v�[�+���,�'��m.0��A=�hL��Jf��A����U�1�����G�d�xʂl��#��� R
��C�� A7P�8��*g��݃@|Պ[b�*jx�)(>���Q�)�
�4/��$ԹTR���z&��(���q��^��3x�po����7���V2� �;xmk��Yl�x߃GN�pm��l����S�����m���C�&G�$&ڀ�I�{fwo���(�V��~w����`��-W�	-���RP���1�?�+�O��G%�E��mP�$?���:<G_i&\�+ҨB�״�����)�� 9\�ܫ�TC�Zښ�9�m�"��ɒ�۾�w~ 밖�N��R(��Q�'�\TP�k�6���q�kԾ�A�C1�v�Ǌxnc.*����JZ��Ӓd�R°�`�5��̫�.}��3�T(c��$�:I�D�5�V(㟍e�O#?�r�c|ćK��Y���b,
,5)K�4���F�^#�>��{���o�u�O�n�D׃��~����ί� �v�ZZk�z�>�$��q���c:�Я5`���=_*��ǣ5�A����[�O��T�|B�*������f����>V�B��]>�:�ޭ�k�)��? 0G�F#6����#�0��'Yr�ԉ����|������^ॉѦ��L�҃_���2P	mtA277k!����F�?����g>���CG�"@\KWo6B{���%�6m��U�*����������F�����C��C���- �hԊ��W��=��Z>7�$����Vo؟#�ݡ�F+�1��M�����*mlmZ�;^��Ԯ!0����?��Jy	$�j����ı�ʍ	�3u�����̳�`ۋʋ�&#��j�2� �>{\A''��r@�^��Yz!u/�B���׶Z��$Ud�����q��+��A���1�@Ze�'87x�
j"�9��X�,W:hv:�86~,�ic��Ƴx;E
��y "�AW�
�X".�$$���|��7��4
�@F�u�W.�A���M|�������^��d�W��5�L=˚��*�(��Ew"]0�*�&X���Ox�h��c���6M\Ԍ}���"'ꥮ��YEI��2�ArU�P��(�
^5ζ�%����a�!��Y|��5vz�lRJ��T���T������'���0D���;��@�4�T�t�hw��\�П�:�=���t|Gx��q�M�-d<f�8:>���^o���S�c,`���	E$�����z{{YɑքG Z}��)����no��9X>n��fN%A1�ʲ��7��zI��ƀ7���z��W�0Hh&26N�9�x���2�Z�t�*h����O�ד�ÇLg� ��,Giؘ"���7��8���駍BY`n<���+��V��͐��Jz����x~��/�$aR]Q��C������f'�-�޹�����/8��W�+�R/z�ɖu��%����M��c��x$C�s�a��������P��|c7NF�;9��G���#�?L��ܠ�� o�lE44�Ӟ��4�z��<���j$H>������?�y~�>�gX�-d� ��(`1���{�'�x|���g�ɂ�h`�O۴Mۗl�?l��v=_{ee%
77�B`{�ZE-M]���a�k�i��27C#C�h:�V�z|�6:T㙣E{�֐9�z���(���QgfF4]=���e�j�Є����K�߱���{RLtq]��|4�c勢i$.6����0t�g��$���^ˇK���PY�;３�� `u�G�z������W�{���G\+{��6��^$�b��r{O�r���hm5�7.��Ǐ�=����޴ܭ~7��ZXє~���E�i�ޛ"�n�i&|ܘ���E��M��5�T%��r��U{���%�Z)n���eR_G"����ꨣe�Fy.�R����'�D����d-|�:Ԟ��Rm���V�D�e߈W��/ޣ��%+����.��0��=*��8v�'����%Ƌ&l+e���&�<�LY���c_$+��|vf�-����}I`��d����Zjzݤ�__/'?i��Ѡ}ǥ֋��4=���c\�Ӧ2��$���]��&HE�Y���@=����k�C��1��)dp�_��G1���9���] 	*�-�Js���s�uVr�J�n�V<'K2�im�vH'+�:�T���~�+F�P�X	$ �q���@�̮�|~+Ip_���`{ߗ��
$�W5�	ߙ;n��<���lH�y�|����%���G�Diw岔��1�#ǎ�PZ�Wx?��G�?�Б<�F�}����RR�b�8A���h��v3�:�"��h{{�^�|�B�Q"�i�DI`�����Z�S��K�]��3��N۴}�/��F�aj"W �{�#������4��v;�ȣ�jQ��jP�D���4��f�x�4BW�¨�j�e���w�Ȯ�]�
�B[+M�f��y:�����8ɤ8N���f"�6JD��\���L�&R�̒:�E��R�(!�y:4I�	�0i����c�^q��bS� �?��<��D�#O	�d�J�aɳ�u�� �i�a�z�������Ϩd���{��r5T�K��a��߃r�a�)�W9�J����þ�ɹzg������&C��vv�����G��֝���p���k�����xDcӺb_�9�H�
�7c�"_]�DP{��T���o���(�o �N��">���e�� To\�`4������jVc������SC��B��;���l�#t4o(�3p\�C�'@wDt0��Ƽu�-�-ơ�|��ﯠW���oL�p�+�c�_ ҌK�3J�wv{{t,{�葬3Ӊ��q��NExƬF��=n�|�I���#<��#e%�mI�f�*ԫ�^��pv}��$�8����"g��<^-�˰fxO4',B]��`�8�>2!�B�Ъs��%FUA�z{5�
;*s
*K(���w�h <��n;c>��O0=f{k�����c�s\�7���=}��gb�hҮ_�}ŀc��&�p�E�1�������l7*��L$��\�����h�9L"��h����g�=�E��q���p�] kk
x�mڦ��l���%�n����)���s���kbǱc��mnn�,����l�vhi��qL�?�#?�����dY�L�L���<ws��Vi�] �8O�w@I�5{�'��'LYa��(zߊ���+��M;&���I�V�d��N���95N� ��z�y�mUjO5���t�Da �� ��=p.�vW ����*l8��MTu�o+F_��y��H?��F)�����.���@r2D,��d+�M��ـ�����������_�@X�/�j�T"�S_;�;\)K�i!_�/�<i?�,Ss� I%8ǔO�d5�$���p�cP����CN���@nk��*��Gu.��uy<$��R�$I�'�
sR,���,xԹO���'rĪ:�h:�g,U�f���T R�U9D4��10;$��x�Rڷ�-���B?�m���������due=�x�"VgΜ�P*�D��p/@��C��Jǁ���U)emY�4"����e�Ī�U@�$�~�M��RH\ ��}?)=�q�y��Z������ �˹T�u�]�����zn�F�4�ZÉ�7�W��fr���:d�~"���z��;;7��+A��o���RTL�Wx%��ׄH��x�@����y�,�ŅE^8�Ñ�ag���Y�ow�gqJ�O�T�q�^�l�v����{>iڦmڦ���%<�����'��� �?򑏄33O�<�t:��ʕ+���af��F@���Z9�n!IH{R�y�&���h����y���!Whk9B�u�1Hw�`Z���'8��h��K�}6_l��}[��dpH�0i���z2��s��q�{�/���忭��
}V��R�Jd�M
>c�������GQH�L����򯪅�U��M���{�Y	���+y�*� �E�G ���&���b
MH�e)3\g�<;��z��ӱp��Vm�jiaX�_^�D�ܹ�mH�E;�e-ẻ��+��:p��.�]2f*�pFCn x�b�G�\ˮm^��33�S�.]Ƶ����ozӷ�'�|J0��܌}�+��9�H����� �r�[�������fsk���x�����%#��^��_��m�C?�GQ)A��O��g^��������FB�<�|r!��]&���)T�_�M����*k�?��sЭ�-��:$`�9dp��`<���l��"BR����=�(
�f��ǎ���+�4i�4!���T~qE� u��Mv��ǂb������-����n�^/.1k�ӦY�6ɂKɚ�J�M۴M۴}�5�_2>��ݾ?�@P�����~��v~>
�4��ZŹ��ER� �I��(&�8SX��$�r��+Ж8���6%u���%iڦ�/v�����5�����*��, �V�%t�R��UU�jR8N���B}h4��}��ta�I��]��C���(9�LJ�Z/?��u�����r�	p5W��v���k4�����8 p�/$Y/	\ P�;��LiD�sYq᪳����B.�[y���,s`�2'W�D� �tc��ӄr��Ѭ��!۳�Ι��6����ٶ���� js�s��5�j�.���Y��Ck�'�4;r�HY��Lx���kR.�*ka	d��Ɋ����k�+��o�)O���{��� �K�4�'�uf�|֊,[�ȨL�/;l��E���4h�Z���t��,A=�E�g��;�Q�y��*`(���Xƞ���uC�HZ�V�-�	�dRW=��;�w�ANj'VI�����K3�>ml��nw��e���sڦmڦmھ6��U7�Q�G�]����{{+��x��B��a�!(:����0�� ���$�5�¬!�S�a�v�՛��~-I��h<��d�HҬA��V�5�]��:�Z�?' 
�IH�[G��p ��� �qq��#�:"aL�w�����zc���I�$K�9�m���:�"P5-���yJW1���q����}�v>�z�VcD�������C��ĕ+-�?�я2��e�v�������+)<d�o}�160����Rh�Ɇ�ï7=��Vp�Aj�)UP4
PJ�>��suE�,�0����0�zj�p���������O<�Ε�U~/��wp+Z �~�'��v��zю&��� hϟ?��4K �
�f�y��F��P0���Y�����6��`�=�������^�VnV�6� � �gZ,�9�g�2��ymɺ����|��������mڦmڦm�^�T8���1+ ��m��[���V�ٺvm������U����lnn�����q���Xcn�+�1���ϡ�ҵL3@8x��,�뙹��/��k}�aMe$��+�&,i���'(^^�_K}�y��Y_%��+@��p9v�^#�_F�W��ޛ��z4�wg��,����K�
	G��((+��8.�2���vv����@����%0-�b���/ԍ����ڤ�r�r��d�CyYS4+�9�^X�w��:�D�2�|�R�^[3�c�mڦmڦmڦm�^�V|���}�<����$g��V���G��%�c��I�a��*�@:� l(����Kc�&K!�`��{gsWېs��8�(�@` 1a�aa]�0)�	�@��U%�PD���TCp- pV�`LJ?��Ja��"E)��t�'O��'��R��oy����x�ݽ=���3'�L ΁�-��iѿ�k�Z�N<��[i�V��S��-.�(ٺ����Y?xZ�\ ��i ����I���S�H5ʮF�F��h4:�jՓ`ZNxڦmڦmڦm�n@;r�p������ՠ[���EA���!R/�'�T���W���k sx�9�V��-�0gF��X3)��vK:�j�2���ag�T�)�$5H�q�9k|��yի_m����C�7�3�`R�������۝�&�K v�S>q�����5��λ^��i�z������4WT,��y����FvPo�����z;�%��P�IM�P��l����^w_*���������:�5s��id�gΞ�gn�ńdU�;E��z��^3m�6m�6m�6m�vZ�ߍ�q�r��q���3����C��7QP����iϰ�W=�3 ��5I3
�/�+%�A%Ș��:ۢ1�A�_So)� F�U<03mT�t�V��6����a+�	�mY7;4�N�\�x�)�9=�W�q����DD��\���e�˄;��Ue�F�in��V~��q��A(�xt��"6d]d�c�:�0�뵬?e�vg4��Ur�F� Kf/�a���p�g�&x(�?g���ft�1�}k#��Ԓ��<�B ���c�w~�w2TT������(�C�gnx�޴M۴M۴M۴��l�F#��fan�m\�
��m��,vqa��wQU����"C���l.]��U�\c�E�<�a��`u:���/'jI$<1��B�!��VM��c]a_�"��1 $�U��:�&�8��zmlVʢ�w�e�3�A�l,�� j��
Y��V�̄��^:�p?�_Pp��´Z3�zb�����3�N�@!��^��4��KK1�d6��KQP�xx�a�)�������c���`GG�X��^��9��)��P<���滿�{���
�q�
?������o8⟶i��i��i���m8k����<��"�v	{[�^��VWW��_��+9����0/���20Mg��1Ph8��`6���J���[���'����\a�e�G `G���?c���Wo�W-�r�}��<��7W �*oq�YH��Z����2��f���d����E�y�9�~�����%p��'�z
E:p�ؼ�+������ݯoxB�c׺ɬ���8�qݍ�#������������g>��;��;���/�������of-����1}o�ߝ�i��i��i�����^j5[�oo�DR��~׭��;;�%�y�Qs��q����j��a�ᔪ���yU�(mE��V�o�E�,��T�ջ��2�CA*ə�M|�߭��5��P�Kx;.F"��	5EPD}��ad4+���*�*�N���\ ?x��/]6���O���~��x`�;���������=#��j����Z1?��?nG�8|)����V\��"T���A�!�q�hL}����q��� ]�x6<�2ommE���������r��?�Q�]����f#�zx�mڦmڦmڦ�4�a�ު]���%��{=�v� �6Sڭᗛ��������[o��<�ȣ��;�2��>dN����~��桇6�[�,www͡��r�|�<˼׵�$�PU|il�Ĭ/}]U_�&�F��L* ��m�\b����J�}��e�H�"|9�R8��L�%��@�:#z���w��W|�����{}�s!�,5�����h����Be8N�ݲ=���ަ~^YyI�/�FQ���$��A?�D�ԙ��"2�.]�dn>y�Y?�n���Xn��6xp����d�������W�q�=���ɡ�`�����}�#?�#�fڦmڦmڦmڦ�ElQN��������7~��̩ӷ�q����>ko��Ns��%s�=�`Ł׼�5�1�|yì>D�������ҧ�~ƈ�C�^՜=���d������h�=���M�r����(,�@T)FzN.˿��x��^���9_������	`A�P��J5��nW|:��h�^툽���]���~����e\�2ʋ��M޼z��@���6 kp�����8�z~~�����7&�����8�F�1�F������?f.L������Q�� T+�e �]q�������������.�?��ٯ���"zoynn�7{��������i��i��i��i{[�v�e�QT��3�щf&l��4s��?�v3�0o��n�B�C�~������l���w@@����0�6���{˙[,"yҬ\��0R8�sЦ 3g%�;���.{�����	J�E�7
"�B��,//���Cfkk�A���q��V���Ѣ�V�[�n乺�`�^k@ �Ԩf������������+��#�T^����"�H@�t���pr]-��t�.�ƣ]��ŋ���\��a7��d��w)=Y��Y� g�z�x�	���d,rgbp�,;��q�b_�������A�ַ�5��w�L�G�QLV���o��_���y��߾9�䝶i��i��i���e�4#���.�3���/��G���UfgQ4K��By
�՟�V�=�o|���É�'�'>�I��3g���>Ips��&K�ɃI���B��eު,��D��J|�a bz^e��V���HS�]��.���P<�"����D��{�C�>���R���;z�$�=�,V@ w0L�����.�Q����C��0��Ȥ�c3���l�%Yz�̙����ho{�ۀ�?�ۿ�o?5j���?����e�}Q�Ui�~�Ϯ�[N��j�I� 8����"H���o������T��w�ü���ݠ��g�~�Ի������uu
z�mڦmڦmڦ��hY�Y�'�h<�!�z��F������-��̃~��梦�7��>VC'c����?~����_ ������g��z�����g��0��X�m��ƃI�"��<}tO �<�ʫWg�Z��t��Xa�˅q�czXkskSj#�^�l�k�����4�{�ሿ/5 +@/J#2�������X"*��vw�\/.̳Q�vh������fL#��:���p�G�`g��6[u��//�d�+��ԙ[~������Ǘ۽ �[�9����`;M��v��t���3�td����x�	3ә1�k���ORG��pk�
�E�N~�{�c���������y��3k��^����O��/���;��$�K�K����hwvv Ob����΀������h\�/fg��a�o�����ϱy�n�������J��u��N��o�w
��������^������}�_P�vw7��d�u��Ís@�^�O>VL���h_��V�=�m��������t�	l��Y��~��S8�jfLo㪸t ^GYh:���z�U9w�>*���>O��E��{��0[��K��iѵ��z����њ�a�9�����hHj��ꅼ^/�z����r�2_���Ö�����2Q��y��KE�y��w��sh�;��bo��E'��܎�������U<���r��^Z���"��[�������yΙŭ�/noO�s��%��^��i��kw�w�q���/4�qo�<�y�7��͋����>�h��ާ6�����/h�E�]\=���Η;'�W����`�g!�����-o����w+�qڦmھLK�6�666�G>�s��haq���O?m����o�&� \xi���������k�N���g�⅋���#�i>���ʹ�s��Es��1�i�>/� ��@C�^ XN&&�t��{0�K����+ڰOnom�1�-u|� �k��s{}u4`5���gt�R}.g@�k�1�x�m:�U�7�Q��D@:�Cf������C���
>�ŋ���������zO�T���"��}��������F�c�kA�'�lX謧�z�+o��EI��������Ц�A�����$�x�+^�������W�^�i������������t��/��/�_IGľ�]���v�뗂��[���������ǵ0L�͠�|���׋t�i����<Ӯ�� m,̴¼��84����1d�Q�b�g�� �3�f��:2v�AZD�*���=��� z�~�zH����d4v���|a}�Y�n���M0��lgm1HF}�3��[[��"&qmi�QO�Im.k���PM�0��64��$M��Y/�"qE֠��k�G�h�X5�9$�FY��i-���!B:�a�h�l��(�p?���z����[2��۬����A��2�2d�f͠�����Z��}���m���`�G�fv;��㒃�m�5�$ٲ4��^o�7�)�-�&����'����3W���Dt���bqa!�wM��8L�4c#��(�<��	}�F�a������\�������KÂΗ��+���lw�b���Wy-�>,�tدS_���y\U��O�-ƃ�1Y"E�0Ɲgɂ�6W�Q�4�,��F����$��|�
I��.���$B��<�Ie(@��0}˟��x0�G�Vkv|����-�[��(g��|8���|6恭����`� CӞ:�������Ռ3��|��t?��1��i2�h85�[a��H��cu�l,�������|�
m�,��5����0]R���K�gR��V!-u[�[B@3yȖu.rA���l�(4p㽝K�G����R�4����3�]2�ji��(��]A�R����-�{���b3�$�t^��@7��F��:om�Cyuz��hp�,����c�^�qR��i��sp�`C���U�M�&޵��p?��S���O�?���`<l)蚨�AP���B�6nϴ�Ao��?�I^�~ż>f���i�]
��4�\�d�cW��9ͅ�����&��&��wRG/Ҙ
��"�\� ���h�c$�$G"���m;�R�2?��r�����:��r\��y�Pk�X������/sIÁ�@h�D�+�Zq��	�V�|J�����p�4��"*"����z����ѧ�s>�9ײpdsפ��
�F��>��A�_4�u�)?��f�h�w���v133��bic� ��yc�����"3m/I��6 ��7�԰��K���ѥ����ի�����x钹��/g��ɓ'���ڥ˗�˿��8Y�}�ɧ�ͧOq��׳�s��8�/#\}��ߥuE��)��M\SE`��+J�6�Af��^ڪ�n������V�_����S �I2.ύ�`�E!<�g�>���׾����r��ss�K��v���m�ms�lҿs�q��̧���y�����K�^����d�4{6%.M"�HK ������{�=�gΜaj���a���o6k��L��v�xx�� w:x�<�N�!�뮻:��w_�~����g���^�|��-�?���F�b�V�!�`�Ή͙:����BN��I���w��Gx���)���Υ��=������3��:�F�6�$�6dK�Iy�i�KA��O�1�@n(^k����6>C��8��[I�� ��cIdU�{���l���k��$����^pv�a�:	 26 )e�~-��I4�9�n��I�-����_��A�pyD:ρo�����W�`�ࡢEa�&��������������v��V��,~b��:�/�N+`с�4�3�����軝]!��wlv{�{7-B����� �D�?����D�A����KKK������8���EP*�$����s繿ѧ��K�'�=6]<[�M�h�~�|n;X�gX�9����С���@��
�^J�!!*p�,^�E�������p}�v�?�Cc���z��
��A]�����y�=S0$�ȩظ.� ��;��˚��紌!ԝO1������u�Ι�./?���s��S>�XQ 3
EK2�}D����,�E�R�ف����#��z�c\3�(�ņQH6	�t����v!C�!VW XR��*�^���H�	�UƮU�o%!��w"�Kx����M�;��>�V���q����=��{��Z����0�����>^��P�%�@=nX}���� O���N&�X�0n$4�ҧ9z'�ЗQE:�E6b���v||�k?��%�^�cر�h!���qGh*G.���2n�Xs��A�K�z��f�̍���,a�a[l�X{�����H���"�_��L��I�R�8?�!���.L)ػY��;�Lc�*�<Ip�YlȺ����lX$6��p�$�l��c���8��5���`��]�A<�o�F�x��yt0ۉF��}*�Ρs�#:�����A�5%�!�Q��g4TpIl0�������"��MC&�U�y�`Ȱm��K�l���4y�mlt
Z{Du��JCX?���;��$��E<'�kfgyo:{����?Kkl�5g��C��z�!�O���������sV1���rv}�{<}��we��jf�}����H��M���礼F^��*p��ʹ&^��oz ������+#<e�a~����e�?��.���u�����7 iMxь{,>{����#��-��{�W�~����o>��Su�#�/�]Y9�I �>���ُ�<m64c $�ر!��k��O��y�7��^?��8`I�Q�a��e����.�!4�|���c�XDǏh�^\YY�{aq�n��|� -��nw��A�-�'jHN�y@���M:�k�jt�N�1O<:��Š�7���s�a��������F��; P�z�I
@Ӱ�� � �0�p�Cyk�3	��?�+&,��L�΅�gee��'�X�>��>y�$@�
���@�gP�@ ���W|����Bf$���2�Zw4!-��y 7	$�t"4&��è�,R�w��'C�~��b�v}�0WUYX�S�N������<ȶ�2s�,a�
x*a�Є1M�l���NCGZ�@ߣ~fapȝ`cv�'��~��C����q%D#��
��� �j�s�^<��~�s��ˆ
�o3�����<O9��
��
``(d�;��k��܏�V�y諘� :�I� !��@����HYF G�%B�5q��G������xt��y�-Ƌd�f_k��X���ɞ���Ɵ��s�8kXN^�}��Zr_U�QMn��13-IƮx�C������M(��F �Ȁ����.5�5A���!B���윜�Z��\�!�I��}��?@�|m#VP���c�6+e@�Z�� ˎw��<Ɇ.�x}9�ת��2S��n�28B�1����u��0�� 0TbN
a(����uG ����^���/F_b.��B�T�r�x�����I��(��U@3r�)V��D�C���H-{�`
��"5f�$c[�n�����@�0?�G��r�$�8����7��| ���c#O >ݧe�Y�2�)�TΊbS��?K#}$s�ף<�S�z�^��z͑����5���;x�# YA���a"ศ�E+%=
2��B2v��h@ڤa��qV�XV�l7�g;�GA/�h�؏~Ϧ&����7�����EA����ԏ[u2�>k��x�[��Gt1Yܳ�6�t4/�o����<�;�w������]���n�^K�`77�9P�ɘ��{���ٳ�>]�z�����H@;rD���?�c�c|ƍ�@�s��ڤ,���}(�T;SO-�:�/7&��M�qTUR���6�և\���j&���<�+�ت�X)r,N�G�-ɯ�<�!�׉�4�Z�] ZM��sϞ�O<���]Z� vaXb�.��
J�����8f�o=~�Xc}}��Mi,ߘ���7��0.������i&�%�qZ�"�Q�i� (Y��_��כ7��������'>i^����[&�`�7lԨ~��'�@K�@�ho�q�wZ�JZ���<����(j�4�����Z�bW����x8�mr4 ٓ�Ѐ���bp�+��4�
b��O?�#��l52�I�/�\U�@�%H^�vw�|�x�����.o\f�,D�l˱2��!  ,�R��ǃ�6X�^[��f��|_�`{05�w:l^ j��ƕ���x�с��x�f�yx�|���7�Z,U[�r�p��=*�y��Zl� ���޴��ҭ���4��5`BC��@߁7
�Bǰ��3��Zx�A�{�H���4aPXCA� q� �N�� B=Z
0�k��W�Qo7�	_MP2���ߘ�z��ClL�s�8�x&X��'aM��Z�Fϋ���,��zb��W3�pX�^w���M��H�x�방J��ȏ�L��% ���G#X�7�	�ɆC��F��k=}A��ê�彼�P��_k�Ðs�ʐ�)������B
Ð_�5W�1�3A����s���/#>Y���To�c�)�E�az�(�<oU\��R�G�aFɲ.�3KZ�q�uB��-���p���ƞ����� �:k\*�q���|������@]������E�Șlh�!�?B�Ք�J����1ck����иM`��Ӌ������g}R�<�&8�r{��a�����Y?��5i.hߋ�RCFrؓ�O:�=�5`	�{ų��Ղ#PG2�\�7����C_k�8퇎D�I�9j� p�g�s�&q��EF�D7�)�v��X'5Z��Ԏ��1����� �����F�����(�8�zX���#��Gq0�PuT��x��1��*f�D@������_�)JV�%���8d�kd�ө ֋� ��̎�#^oi�,.-Z�*���egI�ތx����>�{t����6�9��w��|��YJ�)D�`t�!�L[G
�޸Qo��ɸ�b0��q�>�j1��=8.M��w�٘V��mJ�	9���VhTErUb�Z::=MZ[$�-�4	 ����w� y�3m�^m�u�mxi	��(��}��q�'�In^�d�~7m~߸��K��u �5޿���$��!��U�<���� �mgn3W6�r���ŋ2�i<#B�v�PyO�w`P�92?6y��+Q4o0J_`U��5��>``�j�#���g�t�~까cꭅ�������LQ�<l����}z��	c��GX�(��HU]ȗẰ�<K�����#�nnn43�i\�|�s��̍n/���Yh�{�����4�gi�@�9rđ�d|�A^�������
���ln��6vnx��3������B�xq�!6�~��^?b�# ̅F �(a�#c��ᖧ�J�V�>����Kvd�a@�99وxP���,Z\\b�&!c�lA��޽q�m���k��l,p��{{2��m: ���z� B��]�x�ݼ������� �9"�@��_zW�yx�`�U/��~`�!�f�n�l�t
�	�QO&�N�Ä	�ǧ\<�ܕ���a1PBHQ��B¿	_�xO��>mBBQ�˔���{��K�6�{{6)|G3Y� �ց�x_(9G-K� ���Y.i����7��A2���1�7���+�?�G`��0���X� &A�~�sQ0
@�F��͚=@�!�y�o\k�h�{��!r>�W6�r.��פm8�/�p���GáU{�&�,�F1Z�#���+Eס�RZ��?� �zo�W�&���=K�����t�\��	�W��x��d��9�)��?3��p=�dM��ܩw�@�>���>Y[�9�E	>s��n��AC�'8���E
d�Z���:'����C�xpX�=x�x�1j��'p���@|�1kdf��gãBk��]��~�0�}+�^(J ����2�z�qǳ<���"��r�aʚ7p�� �X�}�=���v�: U5݄�[��O�+U�5ӑ����y0�	8Z	������5?�4,\3��ǥU1��<�l�����U��k}> ������_^�+^�!���꽩��k�衆��8��gI��Ep˱��蜥~���1� ]"vBݡ�v�9��H*Ŧ��Q�D�z_M��q�s����BV�5�#f��}���|�DP��j+�Vi�������P�8r#³~�I4C�����؇��]�s�2ٺ}I ce�^9Fd�Q�N�eH�h�E`�u6Lx����.�"�X�9l�y�is�@��#G���,��+tz�J��"oQ�A�}��L��b��Q��t���me-�2�4��P�Pl����[[Li �	�*�ߣ����xʹ��r�z~�ە��hT��!`�3��}>u�����c��s�Xlx8�1�}ǜ�_���Ml�--.�940�~��U�����������'wx���p�܇i�|�����ٞ>}�}�s����Ϙ��1?񶷙������ʯ����|��쮗�c7�P,�P;rԬ,����M�l{g'"K:�B�A�٤ͮ���g, ,��st���e���C�[Q��������:���V�わf�)��R�J�8��&�� Ā�Z��n*�N������)_�D��M�=R}8��^�!{�ěpd�p	�T ��'T�}�C�9���u�U��N�8��U�=�0@�Z|���CP���N��
�AA�C��Ӽ�c1@bX<x>mx�=o	��>�G@��i�\q��
0����<�lL�YP�+6"zQ�e����1'�~��/���+��fv~�&�"�% S��5�]#�S��s6X�K��x�I6V˝��xh?ʑ���=� T�YZr�b�x��\-��C�ǧ�TDe�5�[� 5�DF�|��T-=�������)�}M�!����k���2J}X��y�EZ<���RYH�A�Cך=�`ת����yO�P%*\N~�;jlc���-R# ��f�N0���Q��r������1`� ��t��}���Q�W>������O��}(�B��N�Ay�j�gؠ#����Q>���3q�QH@&Vk_�;|F �$t�8D2�`Pσ���X��6rm{zf0�aXc���K�~�^/���ue�5R�)I�x~�~]ӱ�g�(��3�^0"u�$j��x��Oq�1��%���3�R�F�g�x~�D���7��� '��B�
=/���4�&�r]�����k��+��S�Z���1��` �b�3�C����W��=��7D�E {�#Xs�{c�-�(�xZ�^1�ZFف���X��l�C��QF�Ұ�x����n�Aǘ/��"#�Gu����Tg��k��<�k7��α�s)��}����0Y���JTC�kV��!���vK��З�%�9?F|B/�K=��2(G�3�\��NO`�>�è�v�v$^��5/^Hh>А�h�y��yL>�䓼?��n?��Cf<�X�;z���'>��-H|%Ɍ�����u,-��s�8��(�	�xM����7���0���.�	0�����x���uLuΔ%�%�!k�_�5AN4���Kd8It{
8B�����w�����55Z��1���M?��^��E��l��ߋN�rj���3<������S�z�/��i��uҿ����4_g�Po��wޚ\��?�أ�����Dw��e�m��'N0�����s����`���Ǐ=�E8:q�x���\c�@-�À�{.'l������̌�8D��3i:���@�
k>6�Q�U#�r��<b�-����}]A_X]o �����]A�Q��L����3JdC���%`�Ԍȇ�q|,���<���p�jL��z:*��S�	�����҆0��a�e��z�>{�Փ���+x\}2Ρ?u�d�k���IڃWB7,L�[[	<���/' ׬�E�sQ��*/��Uk��3Α eY����?ހ�My�F?a���3�{�~��Q�[�L�%VpB�I����C8Tiy��A�y�Q:���r֠���ە���q�{�MC�U�n@,ZJ�*�Aiz# �H~Sn`y|6i1�Ǎ�c5��`I�k�O!Fx���X<��x��%�����&���_/2��)H#4��Ŵ�o�7[oXӚ��%W�t�x壟|l�:�7�}��h��f��Q��_���3l�G�N�Z�|�fʹ/�&�h2SDt��$I�C�m�!�=X�VW+��C�����B�� �
��1��o<Vh��b�]^�z?��s^����C����{�����Hx�<Z3-�v4�������Y�}>��Ng��[�D;�D!3�0Wz���*��x�E�En����p�
��1���Ft�(�K�z��y�k4�����՜	MRE�9�jV�4�9jk��.�D\Y�؋�Q�����ku���dQ���/�*	˨C�F�Q���eJ.�+je�dh�1����(%Ʊ(WtJ����j���N��砋�{O(-��b����5Y���f��G�L�Oi��lfy.��zG�א�Z�U;b�W_� <!r~�⳸V|7�E�@��Z��R#�hA��$�ܿRh}���F�R� .��!u� �9];�?{�9�#ĝΌ�P�Y���@a%uc���,����>�����A��p)��d����j$��K<p܃$��xԗO���E��(%�d�1m&ί�T6�[B���ɹO��}J��x�D�c�̻�}�<D�80���i�w��R�����}��5�T*�;���>t�Y^Ye��N�ZpXw��ř�_~�ˍ�v~m^�y�f��������&�yZ~���f��f7�n�����1���� ���^�:������sL���p�<�i1�v��1CG�)'����Mu3d/2�"�V�n|m��c�k�
 h����:4,�h��W7/����?��c㳊��4a�ƛ�,�)���)���ɒ��\����1Ǘ���7*H�����@M<)��K��� ��}���I�+�EiJ�П�L>������.�[*�L2���J�j��� ����'�N��s(h�ϋ��RfjF�^��5��ϊ���U��hD��R>,�UA�$�L6'L\�D���$�XǇ&n)�C��Ӿ�kF���@��#G��������c�?��$�u�|�O��=�z�)&��¸pc��/j��L����:�X�9����[q�V�A5�X��(��+������c^��p�Gd��g��|���l򘇡H�
�\���e>�`��~U�㓓g�<�}��ϱQ�X�s���B�����D�C���?U��q�י
Aߟ������g�G`�ycO����^��>,��<�ћ���+��B��y�LE�[][+6�I?Z>�F;rO�H�V�Xc��U%�V�(�R~V�������L���]3�؀R�q��,�7 tS^~�Z�B����T�u�u|��\S
S�^x���f�{�J��1��G^��.9	?���:��֘G�+��tL�8f�	���~�<k<���%�����\�� ��Ɛ�[���N����t�@_I?����O$�!�T��>7��9��N�0qXS�����5�?�cpm	Q�5 1���?/U�i��$WxjH%��ΧhB1�O�e�_gf��*L�����h���N|�-��i���n��SH"�dnѳ���Xx���G�!@˞[�̧�/H}�-G-DՄQa��uV���'ޓp,�ه��D:�G�r]+�a�%���Ս`�)`x�só���%?�=�D������B84%���&�����#!n�؆sB I�5�)EM�J �ɧ�6ozӷ�X�؂:����������j���S7���:�g��C��xѨ��o�/����������������Nh�,�DQ� �C�ڼ��bc�����m�ݦ`2Z�����o>��d��9!Yլ�Z�^	�ҁ���x�W��j*�P���E���ˇ˞�
 �b��h�X6Sސ� -����w �� b�a��|�[��*i���h�A�y˽/.�����bZZ�h�縩gS75I\�L6�yo{�ht]^.(�_�ԛ��`�Ӊ�g�D���
{�G�r��f��M�?��[|\��h�ե���5�\�g�,����V7�j�_(i	J�����`<�*��SS���]d�P�00"�]�*�k	u�O�k��E%��E��@�s0�0�k>k}��	7h;;ԫ6���{:q�w��5��\��A?a�`!.AwMh]r�m60����f�Ú���iҕ���X�[�/	oT�虋�g1	�M�!D�̈U'Z���8d��D�]�i�&�2ܻR=0�E�r���d�~P��c���������14J�$,7ә+���1L�3<�S�l�}�P����:?G���\k�w˝�HOǉ���x�l�<�crf���!���S�kb$���ض}x�(ý��f�����))ʓ��f��Z5d��H>c<���������U��YC�r�	�-Y۴�uz��'B��iUri�s��K2�����ӥ&;�^u��á�|1�R��8C�u	kV�g^�N(�`�kQ/���ѵ��^�+��p�tY��d��m�$S�+��j�hc���ń�5'amo��8˫+޸_+4�ǥqt��i��j�,GI����*�P�-}�<�d�>����^K��e?�g�QE���Â0(��wN 2��P���?�Ix�e�ܧ��z�=�Ja���P��S��Z��^���>�{�4�����dRjX<��tF�sS�0�,󟛌cyv�S������92 z��]�rT���:I�V(Fܐ��fJg��t,���G�N9K�n��%�B�9�P�=Ĩ���c/��;�=����{^A{�.+2��;;7�����5�NϮ��O14ni՛7T���^�@�B<���l-����~��+� ��>/%w�ڕ�:���׮]�P3P�mR��B�N�&����3�������ҍ#N��.9��L=092�
�e){#6���۶����>\��5QB�a8��������ذs��%`��\V����E7dp�^$� h*�~}�����$�P�fݣ�1��a"ϫ�P����#�aJ�P"�����.XlPJ�蠖�(�E��e�3I �>dY�$����W��zPԋ��|i(�������6r<�8�"V��	��'�{�Ƀ�r,��OgE����5�ᩱ7�
����.�5�+�Ǉ��-��8 ��4��sĸ�|yC�l�!����:�=�<~��9w�\Y��p�"��{�5����x�D��-B%�K$�ʍ�z���`C=�:��ӈ��1\Y�
�]7_�!��瓟מ;Ϟk=�
����������צ>Ήs��Qy:�5���9�1cR�'�\�R~O�O�����B�Rt���7\q��.���<�xi��+ր7�1����))�O�i���av��5G.W�7�0�����oJɸ_�/+:x�~��$)P7Q��0�)��1����t��f����s��.4}��*�iJ���dMd��dK�>���R�jH�r]�� Y5|�Z����s�9j��a��E~=P��2}:�4�M@��$HM��1�&,U�ᵮ�-W:�C<n5Z�k��T���gS�o���k>��J�$���Gc�V�ʋ|��I��a��s,�h�Q�z)15��Z���1X1��4J���G�2���
O�icO�K� B�8����9
�u}WN���(�DS��Tv�:@upy�4��J�W/v�@R���/�A�i�N<��_w�d"j���l�v��DI�݀�_ĪB����9��*7V%>�nE�xK�40���f2��B��D��Ct��S�?v�8�s��^�� ��D�^���-�� �~>�خ _�6�7������a�� ���G>⣉M^�M ��=�_�`9$���I���k���.ƧN�4���KV�|1�������n���{�{ݸ���t��M7�Po�gghb��Ď��2O����X���$3�\��Δ�#���ox�Y���;l`���|��&u���,<*:���3b�0�ϳ~��\�!��'|����6Nd|���u��o�t�K �7���A�~����'b������*�׷j���\,��� �I�@��b"���<�Ǽ����-@	7�u�^�t�����k�b��Ϟ=Ǜ�t[�,,,��e'PjX�3& 
��>sXݘLh�pے'ڨM��h���`���ƘH �d< +���>��~�S�2�~��͓O>���M����`b��c�F���~��864��) �b� _��� T�}���7g%�q{���뮻�k���.�5�q��O0�����X$J������@�Te��TYU�� 偉'�i�D�*?R7=���������_zȱ0"ԅ^����fD��c��c�Y+H�5+��gq���g��W��|�3�0�FF���E�y��]f�O��>���rB胛����R���z�M� ׀cb\����csC�I�x�T�t��I����xV�*�}5ք'�������/��"��I4��Q
U�P�����@�ȅ�����N��Q��Z�
&{�=�I��jx*�Q���J��MT���R�f�D2�W��0>�9U���AW�7H��h�?/��pDΕQ0�G�S^UH)�:X��,�j��I���j s�>ӨIDA�gB�R�ҫ���k��Aׁ*����^uQ�)�3��y�_�}��P�I8 Y9`q�4��?q2�kyY4G�����&�Z��~��&�iu�PiTT0K��ͽ���س
-J3�=D�ulk���&��L�Y"QՄT��1	�S+�Q��Ј�zu��[�~B5 �j51`����o����W�L������NB3j �'ޟa����զ���"M�D0P���;����8��.�%1D�2��=#
����sV^��g<������/�Y��a��C@�셽'�(ϩ9?L� p����QN���?���E�O������߿�?��7���Kx�p�����@��_P'�H��o�W_���Z�z�
���Y�/\�����9G$?ilL�O�&����^���������u�0�{��8L�_�1��p8Tﳀ��6EGT+$t�Kle�p#��x�`� ě�J���������ڻ�`K����}۽/�6sf�H3#����1`;T*��+q9e��xpbʮJ�R~�S�J"�S�cRv9T��<$�)I�Jv\+8�.$@�F3Bs=��w���Y��Z�ϞAرAF^�~TS3:�}�������_6I���{��F�(s&���a��8���0���a+l���۱ٞ��> 6��{b��n�歛Y&Yi��QV�s+J�������]�^���V|o��n���T(�HY����w18�f5�����H���B�M	u���B��+.:w�j�a�&qYE��vP	��=��(,��7L�񫻩W�.Ӎ��@��O��O�'q�z�u|�FO�es	�X7�9i0����A%\ڌ�����P��o�-H�X�]�+	�NQ����׾��/�(qQ|��P�CRzO=��=�X����Q�c���ey�m��}�x�Q��H�h�A�[��q���N��ޕ�¥:=.��l���}*|j��I��������r�d�4���b5��kW�^��y��V�U�ǟ��!D�6�szm㈼ʫ���D�Wx��%n��8��mc:�(d���_���q�msz}b]r�/�#��������o�@��P����'��N¤P��D���Q�8���_ۚ���Jʰ8��Q�`�?;Au�q����a�/D�>��(k|�zo�������^�j�����9�5R��5Ρ�"|f<cȉ=l���mD?�Bw��".��18��:�~w��W��ܨ�����'.����Ha�k��	��A^Y��Ik,�ҮD#s�b1t'�)��� ��0���y��hn���u|�lp��Շ	ҧW���Y����~�ɔ�՘�m��>�醚v?a�&aZ���~̶�1HǳQ8a�.=����.�ק�d���=�'�q��:����8��w|��iK�xf�7,(3	5��o�b���+<Q׵v�S��,L��,�!��X�fl7hϡ��B�M����~X�ھo��|��]A	Wa�N,g�0�����﫧�B�,~u��
��ڏ�*@�}�>U?'�Nm4uj������7�_�,��,�������C��i��/���KBs{��YX�9e1�����+��>����h��6��>��o]���	y���[������W�_X���8�U�B��o��o������E;�������v;��#o|xr||R]}�Z�w��=��#v&G7�b_�v-,p3{�ʷ��%b;o�!T0�x�'�&?ѭ����M��ߋg���$��V�M$N4�a��͉by���#:���pIW;��$�+��w]V���έ۾,!�f�w��f�k~�i4�U�6R>����?S�#E~2@�[���8
����&�u�|�c�'
q������ڵ�����O���Ʊ^2^Ҋ��C��?�}��&�(pi$*��h���0��u�.����t�)N��t[z�*S�k��/�W���v	ͷZ��م�f���;����U�����kqYbݯՈ�ѹX��Y�`#�a������̿��/���)����$�K�V��m�a�G��Jxz�1��ѳ8j����s'�m���;��f�F����\u�1��筧t�K6�c���I}�׊�NP��jT&~_�P{z��x������QJ}_'
���Y�'�'^j$^:�����#n��)GC�X��B���z������kmW�J?�~�V!j�l�ĭ�Iۗ­�����uЕ	_�1^s��rt��~L�5� �I|�[��QX^;�6��a��Q�8���*�T���g��/��q�7��h���w|�t�_��Wm��VWr����~\����
U�K�ǺY=��J�\���|A�m+�YP�?^jå߻�Ą�C,X�ϧ���KM\�;n�qR��3�S��׿���	�^�0�2^�������,��k��ɨ���6'��	A[�$E+�Q(����]�D�ޚ��:SmwC����N�Õ_?� �K�
&:A����:)��{�	����}����NmUѹ����k��ܷ�������&��F8I��궟�����g�e�����o���Va4�*|m�V���߾���K�H��⹍�V6jj�5;GvuQ?��e5��ˍ��Q��+���_�v9~>Զ[��>��_>{��đa����o#���J�J??gik	�٧?�i�9�֚s�z�q4^����H���Di)M�k/~{舢��W5�����?I���p�|��qYg?���J�]��?��٧��Ӷ/}�+_����C V)���}�{~[�Iq��}�o|���c�=Z��G������k������(<����}�Cϲ�M�|�۸��ov;��x��Kn��v.5�.nܼ٩�W�0��g��;l�èH�T�pcQ{�:��㊣(~���/����T�ee�8���K���j� ���Ku:��;���D��h����m�`�	_����F؁i'/čtZ���:��%B�lv�uџ̓@�W�]l5S����~��jQ9\>�߷��!�fd����HΨ�AO�.�Q:�OU8��L��񠬃�nK�~��^7L����G>��=���
q�u��ӈk���;aM�����G?��ȪɊ#)�Y��`CMX���C<p�v��%�z�N$�c�Y��б"�-���]uP?�p���&�EK�Xbhю-�%���A9v���+����򸽈B`�ֿ�����˄�g%��������Q?�+^���}�k�����'�~U<t�n��)������so'�s�:k����/�(�������]W(�}��k��H�^/���>�w<Q�s����r�F�%v�3��t���~7Lڌۛu/	�~/�hœX=7�S�{���[Q���_�x�������p�>>�8�_�xrq��G����:��Y�"g��1�m-�7�vs��i�镝X��T������5��2���.�dJ�� �ݷ�J�0u�N"l�B�Ȫj^��V�~����X��pU.�N��+�8���u���f���8��&��_lۧ}�_gmW���ye>���C�z,�?�~͎e(��K�k�FI5w����G�?��e�N���z���s��z�|G�����.��D,m�}��_J2��-\ݸq�����:k���[��	F7�~��/?�;�}��7����|O�n[�����0�\�K�}/~M�C�O����ZP�銭x�3�;�3b��xB`'����u�d�	�~���tl�����#����o�ۇϮ���Z���m���-���(\a��sm��F?������>c}v�Ä��H'V�Gw�u���J���Ս����apeN�t;�o�d�����^�GO��a��N��_��N���|W��� �9�>|?�K"��ŉ�z��O{����{��瞳<��.�T
��zx�K��l7��W���X��O�a��7<���#�l����R�4|7�����=ӳ�	~����GݎlV懻�z��u��{g�κ���_pgT=��oy��߾�Π�n��v;��ѱɰ~��`��A�ѥ�tR���Ck�X��3����3���+���bH�*���āp	�VG5bV���Iq�-J| �NM�a�/�]8�*����~)?��
���(�}=��=j���X����tg�����C�o��\<��ã�"�ek#�Z
�7��y��%�FY�vq<sWA�0��wa�ð���~k�
5���QH� �}tae�*�[�!.˻�ڹ@T�	|��G*�}MJ��f�5~�KV�?f7���g����X��YvZ�z��O?CK��;:��>d'���<(b��٪U���W��ͅp��mS�������ݦ�k'��o;-����2�-����t���3���tYX�l�^���u@�I�'��뱆 ��|Zo@��e8?0a;�_�m��9�Fu������?s��q=�6�#�q$9�X���_�X�<փ;c��ڡ���=j��Ȩ.���&��x����c���'�|I����5�Ш66^Yp��mxX��/ �;��+Q:Pk�����o{nqd1Qm�z���"����x99��oN����҆Ǥ�s�7n�qW�M[�N�89H��ަx_��V΋0ڼb�S�~���B�����9���W^�e�E��.�s�+8ƓG-媰鶞�?�='���kX���JWشA�^��*�JR�y�C	�ܼ}[�MO�$t		ǉ.|N��3߯=��awY\)��xa�+w��k�����,�j������-d侖U���������9ƓC?9��P£���s��Bk�5`'���_���'���"�����l�����>��1ǽ�O=���o~�y{\���d(�&i��,,�_�eN/�t#�r���1t�p��3g���g�f�:�\�j<�3��XC�f�_�|<�5��~���x���u����l��n��N*�1B-$�ՀuׅQ��N�����awhWW$O���ҥ���8�� �/��
��~~O�Gc5�&��	��Є�xU)t\^e�{�h���b46!�z���%���v�q�6sk ��"�^�ڦCP��������89�������=���g_N���Ν?�}򓟴En�\y���ߺb�ݸm��u�z�۱_a^�F]��{��x����|~�Z���5;Ij���'�=��������?��r�t�ҽp�����rY6��h�h�|UN����b9������[��Mpr|\�xPk�5�������؊�]��S&Tq=��J�.���<�a���$��Ƨbw�f�ee�W}�{�C����ۻ�~^��X�=2����ޯ�v1CK���V��[��_���Sj�ո�i�d�2@�vҭ��K\^���d:�6G�g��j9o���6�����j�엫Q?ZU���{������=0w<��g��s}8g�V�P�»m���]��]������G������g6٥۫�^��#��)��Y���Ёw���u��ns��r�}s�Qȴأ]ޛgC�t����\t�tv��[M��P�z��/�`�ˢ(��:/��֤�Z�ݸ/W���.���fv��
����n��Z��s���sl�~�/:_=�Ka����&{�2�a:�A8���+w7��ڮz�1�ܗ��������{�
�m��e^��^ݷ�Qv�XW�Ct��{�{���O��4u�����d�w�y3r�o�Q˺n_���7���˄
�]_�l1���myy��.�iF�۶��Z�-��c�%i�M�s[�)��ځ�����)�8~�p���\�B]�t���k�{
ݩm�.���ʦ��6��f�U���sҷ�~z��}u[�|e�I�r�6�Rn����D�4�֭���U��8���V�
�%ZN�\��ں�lӑ���2!�z�N؊�PF�󋹖���2L6�|۳"��"N6s�"�Մi�2T�:!����:��J��þ�SA�t�Hc<8꽉�G�P�џdn+��&;'Y�iX.9�WOV2�\C�+b��w߷�XcYJ<AQPW@��k'���khue�ãN��Xb;�n�����N�4qٿ��R�_~��otZ.z�GӴ�)�E&Vǫ.N�����9�6�P��x�g��#�;��m[�+�,�k�E����Ix��]t�`�p�/��WQ�N����&G٢z��u(�1,
�A��F��<�Y����h����5����2�Ez��߼��m����zrզ��)&��Pc��������v.��cc�>}�ʕ�CYAZp�5��|���mW��1hB����j� ���
��o��久\D�fX��������bw�x�J��uk�廑�uS�S<y8�p��H^|��v5S��:�~��k�yVΕ�?��/�Q�mԵ�Օ�7om�ǉ�9��A�=kߠA+���wV��P��N��>���bv݆]�s��bH}v�J��mđ�XZ{����޻Tq?����~�-}�����N�on\�Q�Y��u�{�*-��>
]]|y�*����3��^Љ�v���t�^���h�X5��W�ޯ�������p��i���}�z|W���~������A#�ָc�O>�����>��ޜ/�W�݃���+��F��.ٿ��_��o�;���b�L�ut�oo����v�۹*�O�2��ڭb����,'Kk�1����n�Xխʹi�0T�O�m��Ա�I��k���}�_w-]�^��o�ѹ�k�7}�[����I����̒;{s7���;8T�Dd�������h|���R�������G��������]�����"�W*��65��K���������;(�y�.��a/i��L�[t�c�Ř����g��#��t_��v�.��q����NW�|T���lk�P�/lDi\�ŉI.�P��'�z����	^�Nd�.����_t���G�ښڨ]>��4���b(}�U�ʝĭW�n�pa����:.��k�~9r[VZ�>�M˾Q���'j��.]QY̗E,;p��N��	�;ؓX����aU�ǵ��YQ����n��c�bY�j�O�����Z�O�����k6�{����ޫ]l�'��R"-u�ޜ���wM
s���׸ڣ� ��wvv�PW�祫C��s!��'���_z.��~2�p���=��ea(��$D�,O�����O�w�"��զ��uA���ɷn��B@/6��ʙ��:�������η��}p�ݢs�>�o-K�M5����RW<�Η�0m��F�����u{�x2�δC)�MDW����=�7�����t�UG��h|zX�dT���bH��]��?������tuz���8<����h�]�!;��,C��pE�}>����@,w��g�TB��c�4_�s|1�Rl�ڇR����U�£�s�����O�։�檌tR�=r}K�q=
W�2�\���N��6��*��	���n%���S'$��7����+a�ɲ��m�K(i���aۉ��"LH/6>���#�����EE�G��<��<X?��ڹYy����v�����Z�?����5	���wf��_Ȟ��3ٿ���NN����ٽ�'��O4��;ww���٫>�~?��ת{��~�z�3 x7~�#����s����t�����.���=�^x���~�7�}�����������Q�r�~����0���==���������r���Q:wy���{�
z��F�:_��!����5��纄��3�&�۲ZW�;$�j�e�rUI��=Q�;�c�]���ծ,4L��
{>.+��]2T�'��k��a���i�B��Jwpw�л�cK�V.���$W�X�}��z�[]����d�k[Ml��\���
�{�;�B��+��t�����$/J��h ZA�DJw@q�w\��P��]�-���Vwi_OQ3`�:ުdF��F�ҥB��:���w�Jg����ۧ�L��#�K�\���� ��
������+�J�'��w����ʍ{�j��G��V��B��=����ۋK��m�y�1b���ྈ��6l=x�E�鎳�7j{;�]�*B��fY��������vqt�ӥ^]
W�רj�y�H�ڧ��x�x_�碑$M��"6�_jԺ���G���iif�V�f����l�����E�ԥR{*�Pē_.��H�a��OG�����+���<􁮺�ٷ��*l��z�G嬃�m㪈sA6�6�m����|~lK��whX$f��b��%o?ү�6?��U�K�|���(p\�&���q��>�k�N�ز�_����݆l��b}��&!�ْՍ_�T��q�3V��(�J�b�����$��ĞĪu�I�-�au��P��+u�%���*�IY��^��
ܾ�&p�a�K�Ha�
ue#������t���m�UO�'n�EuTR3�9��f���m�.�]����¯��j�0��t�pdeV�WX�m�k�s�X�������O��F>,��rN���dT��tqq�̓�w/m#˝_a�Ug����C�{>�����PN�%7n\�>���eozӣ��>�1[����jm���߷]x���+��^A������R�����A����S����~���	���N�>�x��/|!w;����S�Ϗ�����s�C���n�w���[[���x�O�i>��s��A*WP�g��|� �j5ܮF���}誒kex��ܞ�.����&|�`����c�o�������}�`]��Ua�γQQOTR�~��i1,V�z��Tg�ue��p�V�p������d<�pR/�l���Φ#�k��>湝w����Z��.�Rٍ'Ũ�U�ʔ�d\k�߅��p��KK]����G���0��0p�L��²;�k�l�Bh����T�֥򢛸�ȿf�/�� �#-�H�Ze8��ؿna���a4�;�����h��.��z}U�#գ�hv��UY���Q�r����e�.,S���J�p]���H�ޛ���"��ӑ�׶�m�Ӡ���0z�j�Z�=�<�g7ڇ9���+cYHh5���Ia~b�:���F�5�Q�؛��g�C=��6Z�m�FC5ҥ������?9��nv'�����>P�=�����gvm�{<ֈ�&�N�d��Zy�r�� �s���R��Z�.P���.$��F��YgW����Y(Q}�͏9��c'z�v����=����O/ok�͕�V��̴*�,*�k͵�:�(/WK?)�Y����9.���vm�r7�t��W5�U�����3,m���}���;*�aҵ��j�׭T�°/KhZ����	����׼uQR����lXX(U���;�"����FWU�b{Q���~~gw��#[-�J0��:���~�C*E�W��[�I��`gM�+?~y�k���RT�T��*�6?�GV��'��K��g���� �{n�A��o/�dW-NN���#�>��3����Z'�O�:]��|�w~�^���V��<��4��>�����+���F���
~�Bm�,��c�>{�����}��
�͛7��.��}'�>��(T��'yY����'�]��O���F���F�<�����y�k5um���R5E;���ג�������U��u��v��R���^jb+�R
�e��[�B��Ë>w���+{������Ǻ�?�uV��V������
T]�)'e5ҤH�6��f�ە�J�U���ͺ��u�6�r�3˭��;`6���ד���J�^� ƅ6ݗ;@ꅪ��r�kH�R@�{?���!��r<�-gt�`��6���dU�����v=+	���mA_W��
�Z6���v1ua���/TۨI='��b�,l�˼
���^O�`p�L�Z�B�W�%���Z�ki.��T�e�HR��.7�Ye\_,������)
kU�z�[�B�0��9,�k�]��vto|�;ռǉs.�BI�}r���[\���j[��}�ф1?�V�x�!�BW���-�$��;wl�1��j�"I���bxNH��]W�ߋ�=���ua�طe�ʥ��h$�VԴ��:X赳mJ?�����Qͽ�*}ow�����8ʯ�U���F�7�j����0*j���6:���etUN1�Y+��Nq�`���2���g�6t[���okͭ����~Jj�m�X�3v�Ѯ�z���MV�
u񾋎o�=��T5Y�z����DfdԜj�˰*_:����ኇ�C�'���'�d/|{�/����2�*���0ʝYK6��2�v�����U����ݣ����v��:. 3L��	m7z�vw����fy���m+X~��+'�&����6l�m�阌g��sV\�t)�x�~-M�d�0/��p�6�C�{b���'�_�Ǎ����w@��;8�B�����˭���bq��L�Y��NQ�swBP�����U*�즩������U!R���o����k����z��%�Je3*;����|�����Ε.�V\�Y6�|���D�9G��x�\�)���=ϱ��U���_��>�Z���򱆖G�������wO�P�Ne�/�.�+�Vlt`;��*Ս�V�w騮���8��Ġ�:k��w;�;zL�	m��7z�Ʈ@
�Zz��?��4qb�O�6z\�8?�
���n]��l:���?r���e%%K��X��2o�1����/�>��2��5�b����r�T��B���Cªk��J�����:Z���/�+�k�g^��䶹$��ȺE��c��hq���d�Z��t�l[jw����ͱ�a''�]�¸B��&�gu���_:�N6t�7o�*���7�������m�����wAN�.�w0t�Љ��}��J�G�_-a� ���1.��R��[?�����Z�����6�#��M@��ˡ�%֥�:p?2�Kh2�JKT������e�c�m�Fb��]���;G��´�O��}yS][�DkZu��bi��z���5�k�����+jwם9���n<�;��w:��N'�;9:�"H�4/ �%�����3r�����?U<��ӹC��������b:��߼9�U����٬)��	�:7���:�t�|��M&�������Éf�������-���jݪ�{ѭ�z�v����M\�i�]][#�E���{U+���~�Ye䂷�na��*�f����42�:���Z�C��W	mm"Ug+�V]V �]*/�T��jՏ4�%eM�k]�rq\�>�I �݉���g��Y��[��
M�T9L����dT��B��y�W���ڿ��/6K��|����ȯ/m��*���b9�e'֍dVN-�kVd�꤭�⭕�_�S��M|�|���Z�t��4��N��ltZe
�S���*����M3ȭz<�mVوB�F'U�������DA~ݿ«~N����	)�k_�*i���9=�z�P�Y��k��@�b>��=޾�C���Z"�zl_�۬�䶢/3_z����muӮ���ӎwX�_/W��r�o�^\-n{g+{�{�Ӻ�^��p�����^���4�m���>o����E'��Yx I�ʁ�Q2d�����[��:���-�իWs��k*Rِ·��u2P�՚�.�۔@%�X�Y��g˝i��c ���j�m�s.g��F�3���w���~AŮcfGu/���S��e��KW�ɸR�t�q=j]��J�Q�
�#tv�_���Mf��h�����j�jJ��ʅ5���e��W�h|�n��%�;�7���%��U�}�%�G�ܾsх����ڭ�;w�&詎G^��e��ٞ٤?mZ������I��A#�]X��Y�}���������g�J�U�۵��_����_���bP���В1tɇ�PUrR�~��F��R�f�-������s��I=*��/���1��{����q췽�Ym�vN6FV�� ��}����=ԣU�^����}�}�{���U�� @B6�����'�xBu�ťK7�+W���ҥKZN�����=�_�q�G�o\t��ֻ;�`ݮf���/�NQnXU�ޅ���h����u��뾿�:,Ha�.�� ����y���f���}��u��E����r��[8���W}˳���ѱ���F��a�X+a��de����ۡ�����Y�^|����P�j�52}��K�����N�ܹ�}�}�w�����o{��܏}<{"� �W����|D�j�����8��S���?�ښ�vaq_��Z����Y�����^�Z�Vd��tb�RT2bەZ�S���>�h���CDVՓXFP�J}ٰ���n�{o�f��X����5[��:;�g�=Y5o�~nj��C�a���k�v���i����'�O����1��6iN^z������l>����N�'�щ���Wj����  �&UU9���z�ﻇ���r�:��ՉJ��^-^�C����EGf��X?�.��q�Wן�ާ���U���7C�Tm����O��u`P���ʸ[}�:RX?�vm�42ۆ��OCl~��q�f��G��ʆ���5^�p�կ}5{��Kٵk�*u�p' '�����٫�  �&��}u�����J7�U^�eЭx�,m$�:A�e�.��DFg�5��j����2�( WUjg�0��;�����uU��)��j����\�=88��Z�������B�V�S�՟�<��a��F�r�~���k��_��ް��ݵdu�͸�y�{��s�}�v����M������:���U[?O�  �I�zy�ח�syk6-�_�2����=����UX�x2��+�b��jzm���:�e�l[}�߁A�q헶�ä0��R���؊���6�*�H�:GĖj�E]4��N��E���ܲjy�1��:e��yb=�Cp�#���6�¹�����*[eP���uϻ�N'ŭ�7�w���w\�~��X� ^  �T�e=�͔L��]1��u�ڱ�""5��0*�ynm1����-�����*�5�©"�:,�!~�<���6�,�u�����\��K����[���w�G�m�؅j�_�<(�n.�z�XJ�Gg��|�/��������Ϊ��\X��������5��*��k�e�n�{ӛ����UNX/  xMra���W�+��В�.���ɤZN�6«�`
��ԯ��[�#�e
��@}qmB۪�~�}a�׺�s��yc��_Y*[�պ?g�l��kCɄ��(����0q���8<��ϙ�]�ޠ�_�dݯ-c�ZY�������%�7jt�J|���Vh�ʾoK~ےӵ��w��������n��ˏ��-_�߻�^��  �5i4?����ߛU��k�^(��>غ�W-]hti�q�֤���[��j���(����hh+���U-5�;;��Ivxtd+��!HV�-�l��C���о�86C��l�e�Ȧ�6j?Z����Z�p�.t_kwZ�d�5+�]>{�Lwr2/6WZ���N���;Ē�\�~��S���1��G���w���B�V�[,���b��"[�J�r<�74��({5#� �פэ�n�x�_���_��|օ��;;��X�E^�p�J���j��{���P��~�+OW_��-�?�U��=��}����p��jaU6�+G��C�-Y�YX���*��Bo�0�M��"m;�W��teղ���[���!cF/�?Ѳ�UuG��Ԏ�]$4k�V5�[��j'V( �0^�r	�f+��'��mݯ-�<���VMS(�7��m���s�����j�*F�  �I}꩓����o���'�5��v^?{�֝w�{��ᡋ��I�jڲ�o\����hl�4M����|a�pU��nm��&���I���8�,vP���;�uZЂ�������CnKǮ��᝻�����+�����qպ����z��o�p����7=U��Ϻ����ϯeYw�e�Z���h��������t��۬o��UUu
���c�=6�~�����?}�Uۅ�OC�  �YO>i!��O<��ŵ߫�˟�;{��~������mU��Jn޸�����y晙r�xRg/�t=��̭NV�7ͪ�h����Z�ί̦%����*��a��H�3��ժlBAX�x�GV\[�n��K>�-�������j�TZ�򥋿��{���/��ɫ�[�
�  �����~����o����?qt|��.�~�}�Ѿ�Oܟ�������'몢����c������\X�U[lmo�m�~�
�y�}V���eEy�㰺]-={�j�7�]4b�FtZp��ߡ[�Bs�vvv���>p��d��  ���w����'������mko�߯�w�}��.y��駟�w�t{gw�p!W+�������Z��N�[�:�3�(�Vck���:,����wJ�����b̀~_u��z4d�u���md8��\ݎ��WF��<��"�  leG���O|#˿����ݭ��㽝��]2}t{k�m[[����x]Y�g����z<�N�˦�jc-Ȳ*�4�ۏ+�u]������R���&��|A]�}�v��ڲY6j�[�6c���ޗ�u�t��E�  �.B��Q���Ͼy���'F]wg��w~k:����j?��������_w���z�jh�]5�Cז��Jf����%���ٺ�¥-Q����E#*-a����V>Q���Y5M�T�bk6{v�/^���   �z��d�B�Y8��>���?\]�p�>:��ݹ�X6f��}���s��Z�u����e��y6�N�f��J�ٵb����K��:�땅\?��N��_<�]Y�����lo��l���gxY^  �?��a��O�z����z�֢i�Z�L��>�v�FE�/gp!�V9ú͖��|���z����4q�~W+���$6��+{(;���C����~�����/��  �=R��G?�o�m_�ON��x<.��R�V�$h�Zۭ��A_�hnݏ�f���P�n�ZݸR�-F�g����#��V�Oo�^w����u���  �}жu]�#���B�vb.׶k�f���]��[(�6
��l�}��P�տ5QM����il4Woom���Z,��s�ۑ�9�"�  |��=�r����^E�   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   ��� ���=ׅA    IEND�B`�PK
     mdZ�+s`(  `(  /   images/8a1d81a5-79d4-450c-9f72-108cd2673013.png�PNG

   IHDR  !     h@~   	pHYs  �  ��+  (IDATx��	�U��Ow�Iw��C��" ��!�@AP��EDAYUa�W�A	� 
*02��8,�2�b�ٓ������K���;I�[����w���[U�T��޳�gp2Ƙ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!�[:	�9%��f����Bw2f1X��D�KhI=¡�5�~ww�{�<˵X�D�lii� %$B[��tϙ7o�d���/�����̙�ؐ!C�5k�S��H�A��y�X,B&X�0���c;�d��3g���������D^�����
�::���,����={��6��k6?�zD���s�PX�.���"���ں+°�ܹs[�O�^��6	GmY;����_/B��-��Q9rd�4i�6�<x�xhw���5�7?�B���3��Eh�1
a�18���DxS\J3f̨	�СC"��V۶0a�gAR�+,��5j�:��!>�6����u���X�7��6����/%�',B�V'�������,��Gb!���LS�N��!��tꑀ��z�Ҷ#F�)S��DM����-[Z���ؿ˯p?�r�����٩���z�&�"ԼDe��q���F V����]lK]]]	a�	����Ӵi�j��ՋA��7�,d˙�l�rk��`��r�~#���B��V[��E?]���m4x�r�x���g/'ӴX���yd�� _&��$a���Y?�_� �zX(ai��^b�#���r�?�J�D��v�ʛ��l�H�FV'�Cp6`�!�!�ۢ� �G��=�$�Q�v�h��Gr�'8�Y�������d�
�P���քo��7���($KD�_V�,�h� Hx�6�c�������}q�����n����
�>oMX����y�b��,����v���5_���D�L�@�u�~�LSaj.��3������F\E-Y>Qg#q"c��v�ob�
��ۙ����g�A��`��չ��ҖQa�b�,$ݧ�[������[Ա��d��P����q�QS�,	�ňe�ԩ�c�Of��C�I=���\�ųΥ,/EX6ClGh��:�N*��a�I�!F[�<0߻�8������~0�B2�0e`խH�dU�U@kI��s5��������+ �����ܯ��B;A�F��$Ha�q�Z����7�[�*�E��a�Ex�Qf���bPFU�2o]?�Y���		R��L���������������F�I�<����kl߀�O��b�Q�RS�5dȏ����Z��o����l;��?M/v5:�p��<�8\�%�����Bd���*���D��"T=$@ji�H�d��D�Y
�(�P�KA���z�y�>��X=_$^'+���B�57���q�$|��d*�E�Z��Y�L�c�[�g��㓋`���@�ݖ�_LQ-���x~N�E�զO�����ܲ�����d!��꠺�6��7�I[V@X@Q-Ȉ�a�?�<���]\7�*���=Ԫ�g����zs+AM���`�R��m��8��y���8�c)5]%m��x�x�D��@pц !�hʔ)�O��R5���P5@{ڮ@d>���h~��^�Df�q:2��o%�U�)�9�&�ZqTB��	Y�6g��Nթ��X��}^�@1���5,��yd8����V�~�19?:'wb�?�M�Ѱ�T$;�pR�54��gW�����/��1ad�����Y{-X�_c����y�Ơ�h��,5PV�"��N�a�56����_I1�U���dI��M�v5Ǩ6�(�8�1u�T�����DVbt�l���H=^ Lbj\T��M�b0������Xj�?4%{ ��Ն�_��S:�*"�F�^�Q�}����"Ը�ճW�(g`�������T� ݈�!����/�H�eɳcWW�ֈЉwZ2�E�1�C�S����8j��.��ԣN��'b�?j��-����'"N�&�PX���g`�M�1#;����{�Y������Q�����j�G�wc��������c���\q䖟��Ν{Q2����I��)�n�kh����d�Pc��/g��	��1F
4��Fûru1tvv3u��I�U�.W��ܳ��OR��~� X��	C�}��Ř(UDg�����K ��9N�r�*�Mc�4e�{����d�P��J9��uKtHԗ;�#�J���d�K�Ո�]]]۩nMC[T���ɢ���3}�)�E�qؖL�M�W";&��H��az�`,Ig�.|UG�s�r�?����"T��x8ń���T��4�L�>�[�����G,�1c�v�(��@k�"}'��1ޮ���Gf�aÆ}PM���K�ئfe7)��s���(�$D1��ڑ}�&ww(�E� ��M����ch_jUDO\Ɨ���7Ѭ�5k}�-�CX���X&�W][�q �-B��������DgԨQi�����G��Ͼe혫VT!�W�Ƞ��y�k��ה��R���ٳ� -7�n#G�L�[��m�0´d�a*V�Fd�%BjJ������.�Kh�G�{h��8�?�)7�<e�w����灲��5k�f渄 QjIկ7�1q=�x�Q\%@*���ٮ��?N��� @�"<-1џ*�s�|E�a\B���Ɯ��ٹ���Q+\�Ov=��y=�p��r�P�D�ArN�./���Dl�V߫�{v��[���z�BX��2�1:$�w�<�����{9��E'�b�Hۢ�R�9��l:��#F���)��^���1U��ފo]ˣ�oE���}����	V�>}�{�eV�PqL"@&ш��\�؂����$4 -��(SemL��1k���x�Kszi2�[Ru�;�A|_E�WԊ�6p}7q^��'S�PA���/��y�C4~�4�V�?�z��ItBlDv�U�
b���B:w�eT�u��F~/FW��UZ+���;�Ϊ��;�6a�E��rhx��$Q�.U�"w!��q��F`vG�&��ڢ_L����%!��?�Aמ�5�I1p3�dg�,�qQDT�����s���T-jiH��&�B�֪�o�䎋%���q�X�Det��`�h�cY��A<6ͭjr _+�I@$$��r�ȟs�)�/�`V�����7GK|�2���-��R���kܙ�C-r��.,¹�{M�g:�Y�eլ��А��J��*6��,�9+�/Ǔ,�zL�fg(��j�A1,,�9��b_*�Ǒ���*~�05+{���|�c�FL��/�s�;�Ly��:��H�Y���s�>Ǿ/UkT�޷?#�S��F��{ǵY�!���=��|�v����#G��ݛ�󼷫�K��%n�����?/����A��2�02�~�	r����?��Լ�%ֈ)jԃ7�|�}}�����j�#���ٲ ����r�;���:J�q�a�-Bv�3^EF��PT��6���,�M�^�>��=OxN���ke�,Q�ZjnE���{��D��b�7Dh%�ݑJ���|��o��E����B&?�����5�����9�|����Y�D�DX���C�o��by�峤Ooz��U^N�w�D_������v�Z�-���^䏼���V'?	��M���i#�Ѽ_����l�MF{�x��1 ��Ѓ�	!�j��g���ɓ?�hy%��3f��o��ƥ��޼�r�;���?EH#��䡫�fe֕C,�j��"}a?G�h����&��X5�]�$D��ɟR�*H%@[s���v	��~�/"�W����Go����?YF�u�Q��-h��uCUr��(��@��d����oGt�{�7-�~�s���]�'�\S&M��z��q�m<���x}d�ŋg������ROeh|�D��e����ya~Hg]e��v��Cc#f�b��;6�ڎ!C��z�d-z~��4eg]5+((W6N�=ߗ�{�{��>Z�t���X.1.d]����* �Y+r)��#�[��
����:«� �}�������q;S���:�E�엻�����r(�M%@���*r���n^��Y�E��D�hި!��������,�����k�8j����d1z�ךC&:�߭�:%���T����	]���n2�����<:�/QY�K>�k^L�O�V�gb�������L�1bĚS�L	�S��}�V�eq=x�k�L�7�c��-�H���>�ǻ�!��i9�/"Dd!�h��p���������1��d�.���"���Xw�@ϴ��c�m�7�߆4���2���1^,;ڊJ�ތ��GD@��k���F�<���J�.��y�%�7R�սK�����p���f���O��Rz)�n���2aK>Ӓ-̆k֮'|Oq��������Z���X�H,qQ��?�����~�զ�d;�/�ٻ����v^u�_?z��`˘w��� ���"�$�5'm�S;k��q%-"�1#�2�"b���l'H��;����u����G ;�W<Ԫ�
�'��!��k��JS��R�3#�E���>�������Q�]u�E���^�h����x��#�ҮW�x�@;>��"BS�NUѣ�#�_W �W�	��	/��K�Ҿ$K����<wX���z�&}��'�[�`_�+�8��^�ճ%%��Z�ukZ���E2�7�����<-�h��"�eBZ>ŲZ��;�[B�YB����n ��0ߧwl�gE巼�y��f[���8[��,DUi�s��*qS��u��?�:3���}�?Dh�1X���!^�ړ��5\���4�Ǘ*��zѵ��cR����z�<^��X��o��|*�uq�S��9�4ە�Nშ�(��*���&h\�ѭA³e�v�}�"��}�^���R�2o<��f�8khq��Ҿ��#�#��Ļq�7���u_.��>.�A��	�`'�r��ǟ�@Y}�^�0�뚞+�'�k�(Z�k��I����,�7k&	�Ϧ�G+/�2����)�*nZ�/������Ӳ&�s�G�OV�`\hs���|�rboNE�z�n1<%����E�gI�l˓z�	��V|���u���VeJ�����"��E݅�9'���1l�;�r��t�"v�آ@B������é�K�9[Xf��Nc��Bs-5��.e������Ձ1��?��?�B��1©<���d���ٜ��o�Ӳ��T��k�b�k��ݽ�8 ����L_��F�j��Q�]���UK��?fi-%Y;�܋���yd:�ng��9�����3~�;ᷩ�ⅼ���S�׾�Ғ!۰�N���DU%�::v�s�1�i��{�����|� �ePŪz8�݌�!���ZgRjxw����=�Qct���E��ԛ��ep��Ѥ��
��B\�Y����߅�5�������$T���(m	���ʴ��4{�x�D|�����K|�<�q�&Mz?˝S?�"�y����}/�fi�lp*�|�/�|0�zZ�*=`F��������԰jj|¼?�L��V��u	�����l�@�ETk�D؞pvi�5Q�v��pd�n��u���s�u�"�'��,� 58�<��xG��k�	[�G���}��}��T藊i�����r���m�E�o/��$�ЇROSs��%�f��^���r9~��K��+��E~VSW�<����� �͎�.�yF���P�ի�ZDmP}}Y]�p������^���G���E�^X\ѫb�M'�|����^yh��h��א[�A�'�C�$}�"܍9��sH�q۱ ����/��z���y�2�3���x�[�F�+S�#�=�=����ٌgv���Q�T��C�I|n�Y3O��[7�"�.V�<*j�7'��--�~ȾK{{Üs�h��� �ٝ���9�ۍ��S��#<#8^�po�3��25�m��ѣ@���a/��XO�%����2/�*9��f/��l7��e[_=7S����<��z�wD�U&�Eyi�ު̅���q<�M�-�4��h��<'��I��j̠��M��F������2���ėZs��K�U^4x:E�^�T@��U��<��ݺJ�����<�ߓ�����<�����r�����N��s k��Q>���D_��W��H��HYH`��V�R� �q�����d�,oO=3dT�a�T^��4�g8.O_=�*b�Z<�;ؿO�i����n)�k��H�5c��h:�� �b�!����>���G�Rt�Рa�Ϥ��ɓ'��Lb�;�d�p-�����l�թwr�Z��BIϊ2���a���@_���"���?�r�$OU!Yx(��dP�Ft�$�����l;�m*F�ú�����qٳ����<C����z���vWnQ]��=�-bu��3u���<���XYH��w/%E��-��P����?,�U�%���B�׫8+��}+�����,��ʗ���iӦ�N����gf�`K��C)����$�����d��5�N��*����X~�l��*�ݗ�%�{�tG��0e�\T�6�J��~/%.È��e�De�P������ů�]7�`~Ká^"�e�}����"��!;���K��ӈ�|���wS`*��x��<�M!3��*��Y6$��S�X�,�B\�c)�l�����i�e�Hl$@��$f�H��_i����s�^��ա�~�q�e��0u!h�y��"T}u�%�=�1Pa(s�lO=��(B!���U-q�
�Y;�aŠQ��n��8� q��R=Ӳ�3�-E��1��
{��'P1,B��>�7״<��Y_�<�^-I���b�b�݄��iX; *m�.b�t�~i[�\+�!���y�|K��t�%/�W��<Ѥz)V���X�
�%t+Bt�(|��H�m������oM�QS��X"8G�f{X��i�,"�`�����&�QO�e%
c�$&�����/�ŧ(�� @�!���z�r4���n�?+Ue����d9���>"�. �e��H�%��:e9\O�u�DHT7����,��X��#_�j�_/\���!�h߮��f�z42��8pd."-���A��H�?U��Ρ�!��6��Y8���;d��S���}o2ʍ�9��㾥a{��m��Q�=iN��3g~'�(V�Pc�G2ƭd�D/���V�ݚ��G����45�
�9^VP�K	H_�+��X����J3�����]���ނ��ԙ�Lo�noo�V��c�}x���L�!�5d�[X��g�p�/1�n,Nd]�FUl�/�~bt�5T'@�o�"n�5z*n}��n���gmc�i"�K�YR��x���b������YLJ��X��p�5����XnT7��֛k��iӦ��s�D�/���L��w������W�c-@�E���_e���_�u"�c�l��Of��tZ'�˝_�&t�����P�1��	�f7���<��c����dފ	��g�ϕ�HUL����t]2�E�!��b�����{�p�J��mpY�����TRm�c%@yN7�prB�����"Ԙ<"^d�3�e'f�D�FR��1�!�az�&��r5�:j���DP�Wt��L�ajL��4g#DXn��y����˭L%7n�O���gΚ5k��-�$�y����/%ӐX��yy�_�U�/{]?��'(n����4�Qk�&a<6�p;�AnaT�K��2{ɀ�"��<L�:���ZQqL�,�ȓَ����o��[�q�<	N�

?ҹ2Z�k�N�a�5>� >�"S� �J������.E��хi�(�œ49�������ȑ#kn:�`�k	_M���U ���X>����}����t%#v�!����¨�r֌���Ū�QŽ�b�|$@�q���b�ip,B�@E������׿6Gx�N-@Йr����Ss#+����h�*���2�il����
`����Fc/D�V��T�Or�2�QXkS4�G�f��՜A�]k�'>Se	�_�\���]���T�P5�1N��}'D�7�ѣ:�)ڍ�G��p샩9�f�^q���F14f����veߓ�T�P��O���p`yb�~��!�E�5X�!:�㾑�],�x�r6q���
�8��:��IDiO���jϤZ!,B�"2�F�O@�n�SF�|ﵺA�B�<��F�c��RuP�Rf�:�ͥ��6�	(��zd��\m���QP�Lb������OF�.���ڠ�E��\P�����%_��\v����b�A�N!�=S��Hb>�$@���m/��&SI,B�f��4K�U0jԨ���z����H�/������������mν~���gm���F]P�B��'�ǧ��T�P��H�SRO��K&O��NeV՗D3�2���iWD�N�$�d�k)�\�o/p��%@����P���b�W�zP�|jf��믬j"ś��<��V��%[.#���欛bYV�*,O �ű�s����ăC����	`,�!,�?y@?@�c[B�gKU\n��Ϥ��B�gm,B�'2��5��BT�c�����5eEV�Jd�<�D;a�hD�E2����V2�*��J�8�wtt��z�r�}��hm�!(�֛�%B�#�{�ߝ�%wI�}Y�� �P����z�ȼ��<�.k(��š��>U�a�{���O��i�osx����߫���\��� �V�Z���r�w��!���T��:_`��=*����=i]��u�".��J2M�E��1Rߠ�W��O'c��b��%��%@Q�-d�H ���,�U�sS��F�ʶ	�Xc���]0��9:��ƾU�M��""2Z�sJ�t.U��ꧢ�=H�=Iu<�����S������,�P�3xȢ�GM�h�g�<�kc�,��wɳ�F���P�h��fyu�<#������N�&tL�S�]��G�#	��1q��-�v\\����mrO�A��&�"40P����,Ւ�/��d��"�KLd�h]bT�,�y��J�N�rS��b�����#�c��%�Q�\�i�7�5�=�\�3`�,���&�If���m���RvB(�i0���N��:����]�_�"��џ'�$XQ��!b�/��W�흈�D���Smz2���E��?A~��������KDB�oC jC�%
!R��H˘RG��(���߅���uq�GRO��_�#L��f`b2Bn?~�@�<��LXkg,�w�]eWTgG�dt4��$b0�Q�fO�<Y��+��ˈ���{�}������.6Z��X���А���;c,�!8�XvR��4�#YoǺ���B�fp�,H��S�)X8�T^Tݎ�}�E�,�p�!5z5-0PT�/Q'V��
��Yv�a�+!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ�o/�9��l�    IEND�B`�PK
     mdZ��/��  �  /   images/aacc0029-e57d-4614-a443-d9bee65b5175.png�PNG

   IHDR   d   `   �s�B   	pHYs  �  ��+  2IDATx���VU��~�� ;�Nk�}�N&hEa�i�1�)h6�#9���$��A����:�4JEѨ58c�|(��|-���l���yv�;��/��Cs�3�<�������s�sιoq�
�g��8C$�"!�	q�H�3DB�!��g��8C$�"!�	q�H�3DB�!��g��8C$�"!�	q�H�3DB�!��g8��ӧOR__�'---Ikkk���� ��/**zOysssr6�=!rj�~���Ǐ'���I����>����(D�s��}ًlA6A�nd�(-"=�-!���m�t�A�?e����}�����sU'g�:�TY-ׯ#[�^I�:|�ԩ)�Wb\RRR�455eH��%8��3��PΦ���+�&���Zҧ�s�F�c�3
=���ݏ~�B{���D�7�#D72�(~��c����F-�٫�8����7�n�!�*�7q�'H?��S�w444�KdX��w��A���_%���i7��觑#ANM;�&u�l�n;E�I/�}�{t�����Vz�3�^�x�;B��{�Z��p�
��"�G�y�3'�� G������$�嫹�QҚ�����/���!D��0�_���Ƞx������۷/�\����L�"��)�V�����;��@s���E<�0u+D�"8pA�E>8���b��8�1����ݛ�32r�z��>v예�B�7UO�-�6/�I�	1G�a������z$DU��=����?�⫑��]�s��F�[Y㔉8�#��$�bsFOA�4|���N��ȗ����~�rM��D^	�ի�mm�!"�!��zEEEbÕ�ȳ^�K��������O)��A�G��wԕWB̙8f�����/�#�V�!��	��q�ku��wg��dH]���)�"�9�Vg���䕐�#'�,�ְ��z��"�v�nCC�?R5٥{mu�@DJa�t�k��|�I�$$,��V��9RN��2W��R=6�}�~�F��5	ɉ!_�u�P�U�?�_G�+�%#U=�h}R������'J�{f�'N��zVB�6�����9L�z�g���}�s/�]H��2��lޡ�)�?�tϜ���k�q�C�gI��p�u;��O� �	�Q�%�ڙ�S��Z��{�o�7����,k�����'ON�n��`��FZ녆�R]6�=lB��8�/�7(>`=1s��N��Wx�ˡn?�h�s�ǒ^�5�I7v��H�n��γߡw�$]A� ��NsG�eCx��m���vmvG���_Y		��J��а�Q���~[���v״�k��ѡ� �7A����B�{�#2l�뉣��I�Z.�=��9��=)�q�����~Dccu(���Z���t���J;�B�o�g�ڌ��MB>Nن$��!�|�lS"�����+)��5��{��B���%l���9i~U�^�°����܅V�:��5���}�ey�g�˹�a�;��!�詶P=�w���VB��4���
�)ߢ!���		����љ�=0���gl/�QK[S��}y���
io�dǩ�kx�����9eʔk�-[��H�&}^|D�[����r���2k�TP�i.�1��{5���!���1�#ȿ@�v��l.
m隉�m�_-�C�!�V��i�P-z������?1�-4��W�W��/j!�L� ��`g�2�ql�K˗/�f¸��zY�4K�����N��6�!�H/��0`UMMM�,��ty �'����No�����c��
F��!�m��!aVc�y�+0|-eu�&��g��~�Ո��՝u��!�t������i����n�vtq�&��8|�NET3jkk��0 �)cN����QZ�,��?zmYJ;N���!���߮�m���{U{x�[d�cW�Kݱ��0�%UUU�I�H����㰫3}��D��,�l�1| 1���Bh�vz�+d��HjnKl���v�T�ra��<�	����Ӈ��/㐗4u���D|=/yw(T({Q���L�;80QO�n|0���鉕�>��y�:	a�J�u3ΚH~.����PYY��رc=��/`od8����y�@��#G�藫���0�<���1"ټys�/�[��%�)At��H[��)۷o��
}Uer�m�{!}��I�oЎ?��|�!�;�C4l��,$}/i�Z��a�9��q�-��y����{T���y?�JB-�)Sѣ�yJ�<�]�ΐ>?Q��SC��yR��7�Bи�]��HК���{�P�5b���Z�� }�'�ƞ@�	,6��/�moh��z#��-����VGo���U�]�����R�؞�攲��ǉ���-b����c�l~�m�l��?���/Y��	�|�h�.�q�x�8P����xq���e�Y��ZQ�~����	�4�� �d�i�X����lV�s�(��"ذș��u61����ׇ���}mXP&�^c���Շk/�j*6�#����t�g�p�r���n e%�uhmNC&Q���v�.�-h��hX[��\�\�}��a�DkA���~Dz����IpG�`�
:�ӗ!8�	�x���%7�<a=�vSAo�\I�R�&�ۑt��V�$�`�a��'?�S/��bm��� }�\��Q�ꬆ�:�ۀ�[�7;���kB���R�\d�i�������a;�-H(//�,���N��	i96,�2V/R緦��E�ꪫ���	g!B�M�����?��F7W����?#��g��8C$�"!�	q�H�3DB�!��g��8C$�"!�	q�H�3DB�!��g��8C$�"!�	q�H�3DB�!��g��8C$�"!�	q���n*e��B    IEND�B`�PK
     mdZ�1��� �� /   images/1d90a712-93d7-4555-ae10-1782f839eba3.png�PNG

   IHDR  T  p   ৆  0�iCCPICC Profile  x��||eE���Vx�*�g\�$�{�R�f�IvC�]�%�lv7��l��U����E�4��)"ME��   �4AiR��=sg��E?����d�y�3��)�s$���_�`Ψj�̝�h�{���{�U�J2:�T�͒/�,\���Ց�'�~��ǒz}���J��~֝1�p I�W,��K���- �~��g?G?K�0��g9z�J�'�7q<�ݭ�S�d`���>Iƭ�?�ha��������sA/=a`ͻ����;c�I�*$�̚�x��ch̹���A��$c�\�?<+I���g�\�FЭ�m�Ϥ�%�����2���L�Ve)cͩlf���:�����y��C�4MR2M��4�1�5�kʴ\����Ӕغxx�ඝ�{Y��"��t%,I��ݒ*��,iƫĿ,1h�HZ�Ix�:��&��;�%�6I�8S�ׄQ�u ���M��{���K�<@u�ǵ�1c�%m[��&���_��^[�/X:<4k��j4m��>o��Dғ�,�6�~{��ǆ/<�����,��qA��m�b��(I�x0I־<�m��d���䶶H<os
?>Y/�*����������\�\�ܖ<�<���|аJ���a׆}�5��pm�C��Z}T6jڨCF]6�ѕ�;���ţ�����1��yb�cg��b�?��qG�{`�F����J��x��V�b���X�UN���ʌU��j�w�ֲ�-��կZc�5�Zs�5���'k��k/[g�:����7�׽�+����p�m�y�6Zg��7�k�1�\���6���͏��~1��m��~�u�J~��[l��V�m}�6�}y�/���EM��w��W{�+I�ͮc����r��[O7]v�v]_����w�񀝎���-�M����I��y��[���>���w���η�n�պ���K{��6a��ݯ�c�^S�q�7���侳�~c��N���L6����۸�����l��O����[,9���.?x�e�|w�CN>l��O=r���>z�1W�k�=z�~'�;�SZO}��#N��ߞ5����\r^������{~��ŏ_z��G^���Z��p�'�=u�/n��/�~�˭�ܾ�����;���{ο��yp���,�����ɦ�����y~ʋ�_������ޘ��No�w�����?���-�D�X���3�0
�]�ɇ�׍�`�a��='���W�4n�q7���Ru��W��r�*Ǯz�j��~��׼`��׾}����z����kn��F;l��&�7=u��o~����K_�дE˖Ӷ����m����^�ts�ǿ�B�f�o+�5�zzc��m�n�f�o���;v����>���']�v�ΏM~i�w�>v�M:d�nS�N=������~�w�i[M�e��{�����7��+�Zѷ��[�o�ϔ��s�<`�wf3��}/���9��}h޳��\���*7^Դx�%��ׁCK�t��g,��;7}��C�=���W9�z�8j���8z�1��=��?8�ǟw��?���kO���מrթ�/������'��s�g�z�~t��G�sȹ�w�����'����-��܋g^���/���h��+߿꣟���r�:�nv�6��׷��q��7��r�慿Zv�Q��x�Y�_t�տ��o����w>����z��w���������?���{���{��?�������?v��?|��?��§�yzڟ۟��/��m�����?���^�����m�+����߫�h~m�ק�1��ҷN��eo���s�~���><��?��֏�[1Ɲ��ɿvo�a�&������/��5�ͱ���t�����J�\���%��������k���kݼ�=�<���������������	�]���'��֗�M�p��-w�j��{o��ˇn{rӏ�^��+���gϱW���ߪA�7��5�[���o��rǖ��|��-�'�z��]��o'?������Z��b�W��N]�u�n�u���Ҵ1ӷ�}�{�y�^˿q�7��?}�����o�O6�6c�`�̡Y�g9tھ�w����>5����ko��-j[����t�qK�9誃o[��w���|�f��#ڎ�����;�裎9��s��q��	w����>鹓�?�S_]��io�����=�3�?�}x��|p��}t��?^q�xQr�'?}��]�Ko����O���+�ꨟ��S�>����~q�����ȍO���/_���z��nk��r�:���7[�6�s�ߵ��{���u���ܿ�s~?�����8��=鏧>���S�8�O��?=����L�ˮ���\�����~a������}������m�^������.~��7.y󊷮���8�����{o�k�k}8���Ώg|BH�#�Q�Zä�s>����G�ї�i�_{Ӹ�ƽ=�ܕ����ʯV~�ʕ���ڙ�����k^�ֵk߶���>����_��FS6^���Mo����/nո˗fN8|�s��q���~y���]�i�扵ݿ�o�,;���/W�[�=�Q���v�n?f�uv�b'�������:鲶_����o����&����;�N���[���ݳE�iӏ���=~��s{����ߒߞ�7k�C�O�犁�g<8��̧g�0�͡O�[mΦs���8�kA����p����r������J^{ل���~���C�v��q������Ǭ{���Z��<a��8���'|ʲS����ӎ��Q�}�1gsֱ?:���9����;��������p���s�~�����K{��.?��<��~v�Ϗ���kN����~�ˮ����n����~y�����<s��r�w������ѿwW��U�Y��U�w������s����`����������cW?~�����'�}j������g��������=��#^�ދǿt������W��ο?������k���[;����}�9����]��߿�?~��_�譏��ɇ+���,/n�$����]�b�No'�Ӯ<��wW�x���a��R���k�L�R�H`�k��$[�̱j�Ks����#u�l�)y`��������%�Z�Љs���־w�N}'���ڤ��������8-I�w/3������u]�N�������x�ۿ?���x�̞l�����񊜡�!�*n�Ff�����+x�O@����D���W���������M��Fo�����/�����o��*_��'���c��㎡�m�W��#g �N��޷S��a�! �~ ���C�B��9x�-��|K�_��	�v7����x��k>�b�|�x٘.;�LaaB���}�A�U�����߭+Aֱ4�m�'�lP���T�jK�$�����o��ȍ�7"����T>ukjA>����AYƀ[ǀ�	��ݴ��P7�N7W/z� ���!�)U���a��&��u~����X�~��,w�����\Ɠ˰i�
�>w%Mu2hQ�IԞ�m2�N�Q���c���\��ȌdD��q���C�&���Az���>$d����fh�Z�'���t|
�RY�,��b��O�!�/��Mg�5��d�!e�l4�W�1���,��6n������>��m>�b��;��bNV䝽�Z�V*��zZ�ۻz�vW[�g-�3���?gh���EC��U{��g.���^T�7s������2��}r����]g-\0<�?��������6���ӿ��ٿ��L5��I��d�:Ј�������v���T'��tu���X�i�2���oR{g_Oo[�$1��ή���m{m�sZGo{c���jc��}�Í�ޖ��m�}�Szz��u�M�6���=�h�:�U'a�s��v�o��Ο3�s���B3V����wϮ6��sw[�.��)S?�-=m}��o�X����jk��n�ȻuL�Ԧ`�X\_�NVm����̘�jmMp�XZ�R[˔��4V�L��l�h߫mR_�Ծ=��4�6����X��>�mj_Ǵ޾V0L�n�m�:��kjOO�Ď6�T�؆�����胈����Lo{*�K���Ϯ6��T�[���ՁP��U[q��gTZ4;H�Ty��l�W��ͨ�'���Se����͝8�����6eR�ܕ�{ں��A2˳>�4HqbGK��B;�G��6����o����l��Z�X٥��7��x��}_�Wml���tN�ڻ������]�z�v�ֆc�6N��m�{_8a��5u
��}��V�L���݇�����1�����'�����L��[�i���pJA�������u5ɾ=ܿ{��rB�{�=m�=�L�sT2�v����Z&4�#�dk�Sa%�Z�״jT-���U5�Së�ո0�����|��OV���g�"X�E�1+MZQUvSߏՌPR`M5��Q�)SVWtU���/c5�,SUY��pK�	&S!*&J��%3�GGX8��S��ظ��~R�D&9��(-m�*��J��t,�,u�gBXj��GF+�⺒�И�?v4�yVe�k�a�c��d#T��Q�Qe5w��"�i�0��2��T^�b���Yn���2)-��M���(;��1���"���L1[5�$�}d��������יѴ���(Q�T�1�����*V(3E��A�d��8F�4V�Ɍ�c��:�d��wj܎>K@����u^� �h���F,˔��g	�	�&B2�II)�
���DZF����f������D�љ�)��ĖZwdҰ����X��L�-�z6)T�Å[�)�Q��pH���� �ɌT�&d��Y-���:S#�z��!�&�f��c��3���VO` �rͱZ�o�Z�yjmN!�0jR�z�՘4�\b��6�*�ak�����$U�,�*+p��aF�jR��	N��\#�q� �V*���he���5�2)�r#`��=PY����	I�]O��X�m	��b�ؗ�}a	Ο�贄PX2�P9U#�ġk�R�
[�X6�hN;�#�feʉ�ڹcq�O>�s��#��I����N>'��N*h��,�B=��$�!�Ԓ|)�Nji��n�c&ͬ'���(�p�b�Y��*�5o�uDF��Wd��֑��d4#����� mWp�ďȝ
Rc��0h������ؘ�QW3�0PZ���P�
���{������V0v�c���P�GW�4��)X6l�,��.�9X��
�!�
�9�[G����9~��;l�(HѺ�f�S-S�e�)!x p�
6.!j�T����(��?����g�(�����"��U���6U�TBR�
�#�g�k�C�GX�)q�>@9�(^{^G�PEi���p��A3�6��[=� �i�������a��hH��K"�:�+���疤
5�)Ed@%@�f�0�Ԃ��@�pĄ�2�+8#�j�FZF`|!Nj{���6�8Z���7VuA��BpO%N�W�)��J���F��* M(��JI��p\���mf��RZ�@�H�X�V+1�_G��Y/!��R2L�,ڈ
,E���u�$G��¬�z8;�pxX�2�����$M#,�(nY�$����q1����% �T��qdX���i�F(%�:��f@V
SK:@& {��ZJG�CiZB?&9��ٚD�68����#��B���Bt *��U-
K�YOh�m�f�U'U�ۑ�`�F�wrHaL�>��@dX*2-�aF
VO�&a���dH�Ҍt�֎��0Π��a�a�{p+`W�ϑX=��4�גpp��wX�EE���!&: u�"$\�%,��(]�5D�����ı S�c� ��)����W2�>��E$geK2��[��4�I��L�ɠD�ӒL��H~�4�L
���<p0L�_�+Dֈdڥ~��5���e{���*e����8t�đ�U4���u�b2M^�B9%��W-�=:��Q��:H�'���j*��b�����H�#+ ��'C2���U}GA����#�t�^
�uI���(B�(��(��g��z�-�'�X*2�|]8aC���
$\챾#�#<�Qsʩ0�Ó|3b��%eq UC�AHڎ�,EŔ�q�9��!�������{8VSVȉ'�����J���LX*/Q�(.8C�����<�BF�E�!GqQ���cF�f$�.Z芑%E��! ]�<���QM��|ᨒ�#� �t��
�����[�*d�xc=�g >H�E���H�tMZ,Ք�1�����Fy�&B�V1��Y��%�֨\J���nIu'�i=��u D�����Uj5:f%�@�`�P=red.��paι���� eU�:p���:��d��/�� `d��i�@x6+�XZA��?F$Y\80��2b��T���9e��UB�����P=^���c\*��8xPޒY!]� �V��Ǒ
��"�{��b��2:S��& �!�:�hH�(�� V�-q�EGAZ�H�sN
7I�V�Ҳ�S4��"'g�z
"�U�Ҭ�g\,"��J���L��|�
I�GV�Z?�MK�F�\�5�r���K|kT�T��|�����@��%�5�pF�.��\��\GU����\�l8;CU$��'\zH�=���EO���\Ru&���qFs�U���%�=����� ST=�j�EONY���*ydEU ��1Z�-�:~��6p�)%��r�YL�d���b��e������9a�Գ��{6v������M���'+�& 08���34�=y��D	Q��a�������K(=E��B\Flir���irƥ�lG֔�{"IǏ�'�Hwa��o�T%�&@oq��q��ʼ8_M��%3�ۃ�b��V�9��&S�l*+�AظO��lJ�3��L=��9mI��R�|"	@LU"CY)���be
0@CN�ƔH��
��²��b�p����"�p�1V�5�e*` -�s��6N�SF5錕=��� ߗRM2/��:`=\`��g$�p<B9-U�Ud�J��%^3�SQ��rߔjT��D�r�J�f�d�v-�Ne�ڒ1]�5�JPq�lؐl54����֔@ˢ'U2*i#OE?
��dX����k�U02.:OH�Q�N%�IoyiS�l��xIFu[x�n�>H\�����)*�k*�"�PO%��J�Iт�)�r5Fኍ�)�`ٜ�)z!*N�*�@aX)=yL鑘(�&QBS�Pw���fS������ğ��fya3��ss"��<y�����%'8Nk�uC@���� Jz�����?���\����l6��T�'�/����^II��i��lѓ�}�]	XC@N���e./����?9˔�G:Lm1���\A�	T>���y�U�'�,�����9HZB`,�r)I��5	5԰�
���5��ꎰ.W��*�ɍ��e)|�I��)0r I=%�������V�5�
�R9^I��=� uTCr��X0C���2Ms��}Cڢ��R�l�}�O�Ӕ���27�M����C��
[�oG����U�YQ�Ӑ��e�5�Q��<5ݏ �q�!���[f%�6��R�EO�$=p��D��IVҳ �
�vT� �ߑP)�[�K�m�	T�b�S�`gy����S�[��(�
hKF�`��=�Td��~����]ʧI����Jz��39��T_�G����2Y��>i�,/=��J�?�GOS�ocO*`[Jv32q����0�Q��I�  F�ψ9=n��JCB�4u,.Уz"C��j��V�a�L�F����B�\3�S�+�g�%��
�8��È��`�);��)^��O{��y�f��H�4^�%D�J;��pY��H�M�,�a ��E*3����jUYRU�kK�\:w��9���.U�����n``�0���m��}���7R 0x�D����C�C_�!e�BX�	˥{% R���(��2Oغ� �]�/��'�YHH�С��p?Tc��VL*���0����H?�!��j#�I�:�r?�8!������TN�tY�4ܕ�'�7-J�1�r{� �	��T==�AX��7�DQAf�f�,.�U�&��݁�4�dh`�SWa{�/�_����{����IlXn��ɪ��ϭ6/r�a��q{�6ς��6�̈��-��Y�y �K�U���dPt1D4�;`����DO�讑�HXmރ��5{�������?wh��>&��x|�������}F^���*K.I��K�t��������4�:dP����H���H�#T ��{�JIǫ�S~%y������ h�/��\+]��ܓ\�Z�R��x)���"���D��c�����U�hϵ*:u�I���"x#^�������i(�ʽ���v{c:��C�-F��Z�I�����YF����7C�ܓP>'(�6�KK��V���rNbk������(�V	hH�ؙ�� xG���'vҩ'3����>�@J�xuJ��]�ͰObe~9�N<W�M�|6hDrR�r#����f�5�(=i��$N �t�HQ�o���M^�j�#�*_��õc/�A��)����O.(���� H3?��t�x���4�<	8�G���+�$\���f�̌_�R���r�p�9�?BA�7�F�T9^�2g�)��'�Hs��HL���8A�� ��ۚ零,גe䋤��61��taF伂�3g�������ʜ��o�z��V�F�7+�n��.3s���K��]�|�J��Ѝ�8�;��q�/RYDG�QE/�u*�Z5L�g��t�Ϗ ���,7͜���'��Z�x����r�.+`�ĩ�n��Q� !�UH&o<��7'�4�U�+��kԊ���@�T��eF�����^+h5�!�;^���{�X�C��C��� 9�ίݑ���@�4��u��Y�9��+H/�&�nq�2�	�ȯu�d1��+9�M�l=7�)xh�T8��M���>a
E*���b����
�IhWn�E��j$S���o�.�K�+��X�R��
 ��"e4���ר���?�"��I8O��+DՉ�Aa��'�:�zI%d����ݞ�ys��[--���^ؓ�Y�\�D/H�DR������b?~0I�ϓ����C�k%���Q��y)�z^���!E�Γ�%�$t�xYD+oR�@f�P{�y�!?�%��t{*'c��%g�[�t ��n e�������O�I�dA�G�xe~A�Z�~0Lt�H�����ێpL���T��*��y��`B~9V�`�y|b���<�E�k/��כ�je.�y�Yo���qs��j��
I3�I���y������g��z}`)=%�y�������R��/a�[-��� )� S���]�k�>�_/�f�	@f��Y�0T�5�T��@�ԯA���,�K�t�5�<���;o��̸�6��Ht��r��Z�]�Ԇn�3^s(�Z�(Ȭhu�s^�_���w� Y���cO��10	�)�[�)�7r~0�% D ������A-��)��L=��0��n\x���@�5�)>µ$bk �6d��Y0�	r�y8R�\�<bFK�ޜ�U�[`F�@:�8�!����pR{�����GÌ���	�H�<o�a�h8X�d�4>��aA��y���*����!�����F6�*�y�0ٗ�cH���Z���a�n�$O�g1�����P�D�j����Ѓ��7���"��{$a����6b��-0���2�;fȨr����cz��@fao@�1M+��9�[�V+�z#��6��b����O���0ئ��	2�L�4�g���0�KY��GHNI��[�0o/�p��yxeP6La�#$���pł#��@	£�z1��}��ȴ��ĆxН�a8%�~�Ȕñ 'h?n�0nһ�i�:Sx�2��@r;�!R#�a8��c */I�a=o�a����Mʤ�k�ƹ����0�),�f���խ�Kg޽�.����<��X�v�#� o&<o�a�~�
��o=)�q#���r  ����E�"<�'2����rވa�kK�Dz?)�=��@Hʻ
J�6-��T�⁴<�J�x,"�p�Ap
>fa�J�q#�4Ͳ�aCʺ=�ټ|#�����D��*#�F{���2�w
 U87Z�_o�0�|����7S�,�mHD5U<�Z�CNJ���a���y^)����SE�04���
�~�>:�y��a�=�,�l�y��H�b�<����d�tg�������^��0��>���a��� ��ԍ+-�����މ	XH�T ��ވa�+B7��@B�r9Ȉa�o� �ӤB�����g�ܬ�,t���(1t@z�����Ւ
��>Ȉa��ZRp�*S���1�D����o��/��LF��5`p�������`��JŞ�м"��T;��rO���@d�0�����
#�u�[`	�*�*�I+�<VFC�-�@��W�,�Sd{��^s�C9o�a0�I�$G�y��?��a(���i�f� ��a$!.H�2�|<>��H�_A�*0�1�:���'Dw��"�A���R��{�,#���)yH+�a>���H�.���9I�L��"b��0.`uX}�Ï1ZC�����=�����:tCLR��T~àU��
�WF��v1�A5`�q%|R�HJ��,��4-�v�y3r
8���W�o�a��PI�,ر�F��e�I�:S)���Ak���2:�"��-0Z�<�D�g��sSà�����������yC�}_cR��>���|MAE��>H(`�i�k*b���_Ae�O�gY�&�"��O��@���1���BE��)x�R��ރS�������x��OY�:ӾN�"�Q���p�W�l<o�aEw/>D@�;�U��8*bEy��K�t1�x#�Q��^ri�~�=o�a,(���8��vz=�F�~�!�T��G��y��Tg����0
��?'��Ǩ�6#��v��/����/߈aa]0�B���X1�,0hHj�*b���^��@�P�R�`��0h܊���a�~�O��\�n��>1��9��t9�y��(k���7S*6{���е��`�' ���#��pm~o`��`0�sH1�Ί���{Aj�uRGC��Ҥޤ1��8UGC����T�����a4}7U`p1'��up1r���K�ky����g:b�|*��^$�uC~� /1Lx�����g:b�qo�#�q)�;�h�>^5�i�b�3���a�^�Oa)�
$�g�7bL!y �GP�i��-bL�|��y� H���1�PޭhE�<I�sވah
xU��Q��c1C�FS�ɏ��w�1�~R�TC�1KG�)����ݐ�r���a�<��C87#��/t�0T����i±y��#��!�j��?��M�wL�0�>���[�U�L�0hUAa(��Wf�^J��0huO�2Q��U��(B𴆊$���+ӷ�x]7�P�wx����t'�-0�zC7��0��y1�f��>��I+<^7�P��;�$�{�D��"��V$���SP�e1�c�Fp�H��&b�
�4�
�M�P���-b�J_7d��|�Dcx�쀀����j=~�à5�����p ��^'M�0��K����㐉*lP�d��&b�߇�TW�����>U�ݕ�a��W.�u���;��F�1 ���&b0J�@NH��xC���� �I��}��Dc�{����k�����DCu�`8�Ӡ}�a�
*�=�F�c|��D���zhv:�q�0����w����R�ve#�!��^+��QXl�-0dX:�V�[�AFxc�1e�!y T�9[��)|�l҄q��ue1��/��l�O����xa#�J�>�b���EK�Ҭ�-0�ʐgY��#?�Kp���06sϸs�4�4��h#���4l��C�|l������\�#97�y��A$�BH�y��t���җ���s�P?e>^f���}/,�y?��S��>Y��
Q����-0��Jc�P��;��[l�0�A�0�^�2��8��X�ҍ��B��7�I1��YAH#U�Fj#���c���.Hӕ�-0�h��?�q���ECu��7v�����ك�MgA|���6b��p���0N*�-bk�2=�N8Һ�Q�[`K���y+?�Y6��.Z���k��պ�3^�N��� WuQ���   	pHYs  %  %IR$�   �eXIfII*     (           >       F   i�    N       %     %      �    T  �    p  ��    x       ASCII   Screenshot(/��  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:exif="http://ns.adobe.com/exif/1.0/">
         <exif:PixelYDimension>1392</exif:PixelYDimension>
         <exif:PixelXDimension>340</exif:PixelXDimension>
         <exif:UserComment>Screenshot</exif:UserComment>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
����  ��IDATx�콉�۸�%�R.��֝������_��V���$�XND ���t��v�R���+6�0�����e-k��IkY�Zֲ�)+��e-kY��Pײ�����
�kY�Z��BeԵ�e-ky���Z�/����W�E*������+?�Wj������Z�^�#�� )��~�:��^T�#��J�_��m�P�B���kP�? �����S�מ���{������)��⽭����
�ky^9Ÿ�2��S����,�������.�[m-g����k��6�y?Q���������S"�)�h�;�/�����b�<&;���%�+U%�Y`��$��\䬲2������W����b�����m�.�z9Su���dEȿ\Yu-�+-�{�H�8E-�粒�K!���ŵ��.�:�{��r������31���Bos0]�YU�[9y�s�t:O�%��F�tc�����
�kyvy*�����<�g^N�W �"ߺ�9&���H�6z�~�iE��<W���oVV@]˓�S���cs%�/���ߜ�ܮ2V4�-3[P�>��\�g���M��nN�ƧQ���GY��
��
�k9Z�#���T欴����F�RZ]�S���k��Z5�Ci5����=��aHc�:���yb�y�o'x[�[x���UAG��&����*`e�߽���/O��S����#8T`Z�E@52Z�tx�~�����oT�qt�Y�K�}�3u�]� :����^=�����O�-�>}_O���x��Ȫaϫ��y�c^c+�����Zf���R����@[�1�$L�t,�E��@�X����2��~�����z){e0�ۇ�0�Ff�1���
38�
���
��Yg��L ����T����]�������9�+X�sw8Wf�� LNc9���РZ�9�]��-+���*?`���&s���1͆5���6=���"3@tz?iا��F���v>f,�r�d��M}S)���O����|���ӹg�I���#q� :A*P��AX�&m�f�]`�`���I�(�����^��ȼ}�?Rl&��n���m�й	��k%hg��4ь���F�'�"O�W�ݨ��+�~Ӳ�Z�� '�E12Zׅ0f��
	���0��DxگT0H�~�^��A�*��L�DPX�\�^�T����T�RJ}���cLZ���m�S���f#�&��lz=Q2F�c����$i _������jI]@������B���K�Q��u��YV@]���`Nk<b�:� I���4�Y2;$ #�y�,P�03�����o4 �R��@�JA�)	"�� ���=L�c�+(UlGPG�Z���>ȬC��.9 e~|�6�N�7�}N� u 8�#�8Y'��m���L����F�&��
@s�^k�>eԵp?˩f;P��=K�O��e"���l�>*�ƫ���HA� f|���}��q<Ui�����&p�
��z z�*!��&�a�ߎʂ�32��ޕҵ������'?��*e�T�N����Q�i�6�z�L����n {A�f�1|M�+���+�buV�}ղ�Z�D�(�Q��@�%,rd�0���Yԇai PԖ�����W},t��e�S4��#�c��Nu��Ã ��+Z����2Tk�&+Ƨ͸��ઈE5��TL'���v��m�y�z�}/`K���2�����q�ir �zXUf�[V�~�@�T|��h�򊨯ZV@������	L�k��a�zI��P�'�0T#���u>��d�5
��k�^�؞��C TX�s�h��v�J��O�}�ɋ>��Z�[ֻ�(�2c{���i؎Vo��(D�SV�V+�����J��*��ꔉq�;��AuQT~)S���w�%C�f:�6���^ky��Z�D�aQ0�����ab{�P	0Х&��� ��Ea0��jPu@Ы�1�99��~�*�J�g#���=Rd�������d@X�>L��^ݜ.JӺ]���ưN�h��Y��_��+�0S�t�D!��=�kݧ���U �R/��xq���b����
�߮���/e�;ܞL7�M��92 �u�Q�z�J��`��3�b�����	�*�=7�������H&�:�x>��9�>s<ʂ��o$P%�?�������~,�@�R��r�U{��܇�ɹz��E���aL�� �J��6$L,��>V������nY�g.�2B��?�^S�QHSv��#�� Jb=1у�U<UW	�����۲n#+�iw����Y+K݋�lT��t���!y��a��9�>�=��x1X��3�Q�80��MM�_���cF�mb�}�w�/b��c�.]�B�K�����jˬ[_=Id���|;�*��C]�u�
�?k�
�'���Y��Q4�(�򧴟���CuT_Tb�����h>
uU@1��W��(�H�%����>�u����p ���BDwڣ�R�^ҝZ}��:���� M`�ƻ� /��6,5�*'�[8j�PO��%K�e1١W�t"_��I`�%���.��#�����'�^A���
��r&S��	#�3Ճ���M����������\�9�ol|�&nT' �]�;+����'��A��8�ٿ�\��''꣆�	����F��M2��s�SWj&Y}�AY?���<	e� �~�Ć�"Ʋ���82H�w�����E��Sz�≡�9�N+��NY�g-O��njY�	"^N#�\���$�!�8�a0���
|2�Q��x*`nD��X�+e#����4�L�Y�2f���HH��[���Do�^ �aol�a���j ��L@8�> �q�4�Bn��ս�M��^���U�oj/u��Q�F1��'�8�'VWկ++���%?o�,�:̪���h��i�������Sa�c�cnY�k@M����(�@�O���vy������\
pe�:֬���f� FuIvy��0��Ԩ>�x����_[�]@F�B�R�-�/��P����>?���8��ꞥ�4!� �^���h�����n'F�}����hp��ak*���	�&�����>ki�
����Nr��_��}�1�k>�AY'{  >?	 r|� �-ؽ�xS	��p�,�	Os�5kz�4tp���r��r��Дx���*�j&S�&�l̐� ���ɋ�����v�s�S;h��D ��9j�*Wq����̵��j��Wb���21j�~��t?�S{���ty}�����U�fe٥ ��7���Ze��O*+�����c@��g��TFX����Y�`Qgq�#SQ7)=n���}����%"����	Q��X�$K�k�~�Y��3�k}�VZ�
�NPQ�;��X�W���دS3A���\�UJn���FV��%0����	�&�X/˾��`A�N�<�� 5�8�UY>����"�.��X5���f��r�bi����eԵ,���t|�j�q_�=����c��M���&X�ᜯ`ZԪn��z,�j��������+�Q�;��v{�W��>s����f�����q;	�b�g&��7��^�F���aC�6&=h E�̘|a!�w4�l����q������+��zӵ�\Yu-GXf�Q0����}���(!wib�(ْ(��%*�N��Pr��2�Ә��A�� �� �u$*�of�RJ�p�NQ� ��#�c��swY��H�/Ġ��TǤ���t��,s��vX�
��؍�t�R�6u�_��x�+׊�߶������@�O)\��yj��'}Cuf	v�Qu������O�Ы%^�7 V}7�X��w�^����t�=��"�3 �3v�5˾f����@8��~���$�_ �3���@�G5��<����(��Pw�i����n����35��y�q�y[xҘUN�VeԵ�,5���A�;��ߖ	z�h@J�Y������"�����>�q��a!��7��!u�f�,��f�Ϋ+�{Bl�<����p�&ɐO�ˆ�N:\� �����4w�����8Հ6�S\��Shg�6)���`[�ۘ#��0�@uk������Vl}��ZN���q��wџ�����0È�-,�A��PŵI���� 9�rT��.��T`�����ד�4�9���k�j�Pz�$������L�9��R���ަϟ?���/�V׵�TCӨ*�r��c�F-�K�Q�keF����H��c������>��
�C�E}[~�y�+��nYu-��`��>~���nM`c�6���{H���>]^\�w����Ǐ�N��ٌC�ܬ]j��V��U@�u��y9�+�z)Y�9I�Vr�v�(�7�v���.�����?�d`=��T�ڲn���;��(1���"�z&��v��d��&�3hCe MA0��$�	����X.̳ %j��VM���P���v���:�U0��&s��-�3�kj>�K��~�>M`����]@��;u�Z�0��KՔ ��VD,�jb��W��J7[] �Y��ڑ�܎(��/�>ML���*���wϠ��\�b��u��	#0�W���1�� �3��J�b��龓�`��A�c��X?�Z$⦝b�W)+����=*0����I�����9{K����s�!92�1?�?��/�����ҧ	��M ���]�%�ذ��{��kg~��f�A��EO�ܫ����sC�?����U����1��L��	`�'P%VJ@�ɬx��32r��ov�`-� ����D��Gne	� ����b1V�6JFO]�4�
�/ZV@]��3W�A-����F��]��K�5�U;�2}}9��O�" %y=����W���N@K�U��?쒪X�F���X�Պ�Pw���~�ji���1�ը�h��t�� ���2K=�������y��Z���b.]b�ww��N@�W4��^#�,�`VՉ~6^د�X��چ{_�R�^V@]˓J���6%�G0�@@��܌�j����?�g6�)���/����h:
K��Sā\�r��`ѺXڹ�<7���k@��� � @��(BE���r0%����;�����3�U���/_җ�M��QX!�Qb�UG�����7�@L��î���
�k��A�8rɦT��h0�G�cԳx22}x������0�n���-m���C Q�ya�ǳy�j���>�l�	��N�{�Q��='������g5P��E���,����������/�y;�#�z�Yu2�ʪ�D��P��q�Z�aq������������Z--;4�I��;Ď&������_>��������l�����?�;�B߫�ig,ѭ��k�����XfZ�����\c��xG+�X�����y$�|�.�M���[���gw��j�LSYWP:m|*�,�9�IV����
�kyva��A���g����=�ǿ���믿N`�^���Q@ S�z�{�������^������	rmS��a�t���_��c��� �[Rn�Nd��u�r�Ng��VV��eԵ<��(��f��Tt�M���@���w3��>L�)����`
 -&��7ʤr0�����0K ���l��5�p8C'�Y���+�(�7� ��{%�]�T�'uK�ٯbkU���Vd-/TV@]˳
'�`8ʒ�sԤΚI��x�����4��-�6b����"��1��_
�	a���ˉ��g��텄���L�3M��������s#O/˲�/+���YE��� n�zM�D�R�Zԭh��O��r�oލR}#g�3.����_KP�:����ID� 5�!�Ԧ�!Am�EuGPV]��)�Ϊ
���/��|}Yu-g��2��12��>��_\hb�1Sƭ��	'�3��^�z��^�%�Tƺ]�dݒ��MKA��TS�^\�bV���SUk��L��Z^�����g�����8y�c� ��E3�5�Mԗ�ʄ�9��o�N��>~�-����l��3��fw1�Q���3*�b�$�ww�@�Z��g�P������^ˋ�P��ҳ�~ga��E,ۙ�K���q�aj3�Yu�l9���MY82��*�Ю�9 ��VI@�ȗ���nnnd�BՍ"�ku������p���FYu-�*+���6 v�5[u���fqMa������0�#*� �c������^Q��H
���޽���?��$-Q̷����w��	<����lX�ox-�QV@]��:��R,�S����r��5>��Kiu��aJ���~�-���c��|d‵�U	��)k�9 �^� �D��ޞA\R�&0�lu�p����b�.6[[Rf՛�nYu-GJ͛\�T&4J^҃f��]ɡ�ܤ8����)�S��2|d���qx�s|}�L�U�.m��Q��=,�ਫo[^vE2s��4�J��Q�Xue;Lu�w/�W�/�$�'O	��������m?�7QV@�K����ϩ�Zg�w}(ńS�����d|!��t}}/ ��d�j��i�Z�I�\��o������ˀ����/]�pػ�D3E�骪��y�괝���P�O���Zib�K�vͱz�QH8j��1�w/+��e�1�OYP�|�P���.���3��$��G]ET+X��s�֗��&F����R�ѭ-���8�C�錴'N�M�d'@���~8p�n���jU�w��ny�� �U����2�OS�b�rnYu-M)�w�1%���e���ձR'ǧ7��@�]�G��W c��c�[���6[ ��v�J#�S
����EO4�w�
�!�
�k��`��H9nM��q��$�֤� �ܞ~����L2��`�	5�d,W=�Ǵ��_V@]��%lHݗcZ%�AX�D^j�z�%Jx_&*_ƛ�MN!��uԩOk��eԵ�J��z6����<=#�3P6Q� �#�ܲ��b�L���V�f�2ʮP��,��r>�͢']i��)+��EKT�	�*��ſZU����x6��j^���?cy���6�-=������b.Tk��)+���*�rѣ/�=^Ԭ����9�^��.2C�|���D)�>Z�oH;��5���t��Z��/+��%��O�������H�U\AU���y�ρ�W�8������ ��.��ujߢ~��<�N���*����Z�(=�R����{��T]�h����e��K���	e�49q>Y��U/#���QJZ�(+��%��^>�f~�) �g��-a?��	Q8R@@�T.���K���4�q�XF�Qu������7�0sn[!���P�R�*Yq�cb���MD~�������)(?���הe�_3��Q�/I�$$�'���1������Z�E������:�~�Ė�*'�;��,�G@5bK���U��^�J�q*�t���5IbiZ�g���bv�@\�;�+�u��5�
�kI� ��a�#X&Cj��=i��<ߗ�p�O�a��S7����}�"W����Ɇ*I
B٨�d)�W�>�U��k:e�#��e�!�g͉���8MH��?������1�QB�T8
�tӬ�%M�g��sr�1 m�tmVKky���ZB����V\�ޟqJ�&��ђǷ���ߥ���M[��:=H��O�E�+����4��Z�٧���;�.5&a���/��ۻ������U�h6F�҈ﯮ�����C.�Q_�����gЇI5FDl��$�Po��~��1a]O�H>=�E���5�r���?j1��X�Y�e	�����1j�~��'�����n� ^�Rٳ���<�D@�gs��T�Z[�S�mYu-�.4Xm	���j4!@�����/����{U$:�tq�d	 �蔱Q~O[�*�M����
Ƽ����)��a����s�׿����P�,�k�=by��M׫��h���ީ߶����g[;*�`@����"������-:�w,��c���
�?p���at�6̒��
1Qb��O�MH�7���6ݨ���#��3zc�wK���oRV@]˳�XĘ��:.��EJ�~�����	DiI����������΃LJ-kc=k�9
G�M���;1�>�Eh�م�'N�������ϟYM�T�� �IE�d�Pb��K�P[�������'ʏ<�����g�����72If�Q�SY��J�o�>�T*��I�puy�����XE�8�l��?��^�b��6��1�Ll������f$�qoT}2��8q��r;�<�* �Tz]T �!��u�
�kyV���TG��,H�DYұ�����ۋ-9}ާ�>�뉹r����?�طD�p��bL��"���p�`����g�����ݝ���(���RK�W���t�ky��S��$j<�^��X�d��2�n=I��w���~zu��yi�/7�׿��>}�ȫr^\\�Rǅ+z�L��
/���ӷ�[aϊ�N�vj��4��M��?������N��zg�0K�/�Y(G��&6Q�m/�ar���*��ɬU��疷4nj@�i�eU��������/�Nn@����@�6}��O1V]���֞�L��o%]k߉���.R���ŢɆ2�B{Nm�ۿ~K����͠J�I�
�)��e���
�9c9ѭ
�)c�����F;�^V@]�3����Q}(Ch*�N���n����N��ߥ/��ӻ�k��__]����һ����w�����ߜ���-�׹�OJ��� �������a�����F�|�)�3j�~��U0���/9'���=���Q�vY�(�!��7�����T;��YC�x�"�N�F��<"�&۲'{>�yx����<�F��0��IEa���Kf����˧O�Ç��g����Y 0>O��_��O.��0�(�e�:җ����������Lc�>�OV���,xMPȮ�ib�Su�>�����e4v*�W�.D���,��Hk,%m9�d�Y�;fy���7H�_PC��,����vé���J��Ի��W�4���}^���8*�'4u4���T���t�k㿙�N���O��*��mTv�Q>c}b��b�~����8[Rǋ��b_i7���~z�������K���[���;V���)��9�|�������Bg!�C�I�x�ډBI)�>1�/7_�����>�Ko���~��]Y;j��(י�c����v;MBW�ӧ_�I�C���ּ�F�V+Ћ=.�cT��O�鬛����q��p�:wdDپ!թ���2����縢̧�� ��K-������8��b��N<��I��R��|
u�C;��,��FBp�>�vNef�"�m!��Xr��˒pH	�Db��9��}7�GvP'������J/&�~��h���t��p�Ʃ.{�_�~��"� �Xv�xUR�j������S��:��g3��)g���9Kg�"���7�˗/���n(F���q:�����uY� �g6h��=�F	��tu}�>~���׿�=���_9���X?���(�?�����S{S��\jm������ ���I<߈�Wo���L��U��s�"4z@ ��@���ѷ��%z2+0����N-�^�L� p������U���j	��-1t��vKK��d#h���n�<Qo7%W�a�;?ed�8��PDI	C�$ȝ�[/.�	'f��/�;%q.A��'༘@�D���{v#���y�Olubg��_%�Y�5�]���6����g�C�"F>d���{I���w�N&֗�OߧɈ���ECmyr�	���[�]�V@�� 3�T����ԾW8�ي��|Y\��Ѯ=o���_�1JO-���޶ ���A'����tt��x���R;3���U����S�?�+�Y�+W,U��O��č8��7p��[u������7~|��A��l_+B��� ♁��1�K��4�qRp#�Q�ԩi@�tK �����Yw�NR�� �� ������_�6�����ω=�w�yֻjl:��(��2����.�劮7*S��>	"mN=�1��;;؟<0��N�Gq#@� �d�}�u/1��d�Ԏ���u�Id��&��Kn[ *M�^�~��ݥTCv/�F��h�:j:���������J�H����R�9����3ڱ�.�.��N:�N����i�^��I�"R$߹���
���Q��.�1�t
��p��\Y��%KY�@�t>�V�W�� ����X��Y��[�q�3�쳯���xQ{^L���I�><���
T	�4����	U ���}����T���|�T�	Ǡa�\{dT76Ą��! 3��ª9kTVJɶ%���x�R����$Hf����n�����.a)ӣk�$�6X+OgN E��3`�X;�>�'�R�5��Nz�<��Hi�OU����r�?, }`
#��_� o\��9��^�@���Iy@�Yf0P�b����yǏG�5y����+�\�s�\6@� V��ض��x�a}��:����H����ދF�q=���kre�28w?�'��4\��+�h��	H�w��Y����{)��wiV�:a�����[���Uyb�@霱)�I}j���&:]�$�����6��q���[GF�Sb@ꅹwj�g��`�k��K����9I��44�#�N�t�,5���#�DVZ�����5�=��c��GH���,���b"	���Ԍ�ţ�_��D���^j�e�Ҏ�]Y��ce^�q,�9�u��L�����BK�C- ��T�}����uD.N�E�E�TD��E�٨���Tuˤ&[}��<���o�W��30H��:+�'��'����5�p�T-ꐔ�{G�+Y\�Xt�2`O�l� ��f���ML V�3n&Pl��ܱ�	��TA�a�TW��j����̾�*9Y��ҡ��@����y�����̛(/���:�y���Cl`P @<�Ɖ�r:�3ƚW�.A�/~^bKK��F�_��T��C��zܑm%��}Yط�ޞa����8�|����/ׁ�Xerյ�a�c�c���E�/����R����a��R¬o��	<�Ȥ��}%��]ۑ\�R�)[;��ψA��V�� �*�^�7|��P__�'2�#1��r?ZÝOH�$b�lBxrc�|DG]���/X3�س���|V�ey1@E�!��l��'obW��h�o���#_�\�1�c�wv��>�T�m�`/2��Z��1��zC������&�����1�	�_��Q�5H`�ͺj�l���� �-"�Nܳ�����]���!���3��<�tA����F)���0#��1��I@R��z�M���1c�N�Af:�P�y����52Կ���;πG���1ql�G�.��%�J�q�nv��+�����/*�cq�)�d�ŵ.k���\���ŷ�*fb�.7<���Ͱ7E�D��k/t��G�d�'��稾�A�Vo�0�þ��ƄΗ'�z�%uGJ��O�*��{�p���۬KR�b�fpʝ�`(�����~�:�6���0Hv'����u{6��B�V���YH�卬��;{���S0~���z�����j��e��I���+��@=!��1�Wڥ0��������m�<໗�Tk
ի�c�0��Y�s��+߇q>�G�k]��":Μ��R����+��=��&�B��Ĕ\�D�-#������ ��u�ڛ���������Z<.2V����1W�x[(Ě���٩�� ��E�3V�pP=���v�T hT��*��k���%�/��\4+-H�P�Z�ɥa��d}z��:�Q:��"�9���u-#EI�3�d��c�?�y��Q���硄�v���K��Xz������P��j)�Qt�\R�(貦~��GQ	�dl�1t�J��Ԓf@cU�W;8��V�L1�DT',��D�Z��l�GJ��Ei�5���%2��銁�ٰT]mS��i�"J$�)̔\���W��&�7�0YCTY�J����@f�#IAَ�@���JT15�EW��*F"84"|d�&�4�(���ˋ>J�)4{��E���m�>�1�)�O�i����;j��RUÁ�I��f�=��>�0j+�����U��r��E�E�P�ndP1K�^siZg�
�480� �Ć�f����[�x���-͜y@��u,uL�f�#�w��B���o'�՜v�zv�MK:�xYc�%N�\a���6��^�:�QYc������'�ր*��%�'^�u.��Z���Z	�(�J?��L�}"����	�f<�O˽i?���`�� �uס\��6w�>@v�O�'*��� -��ȟZj#W8G�� �-�]��::��N���RyQ@��!sg$�|��"l����e�ΒC�l���f`��yE����g��<Х-%���,c?����q��!�tq��3�~��p��ejev\	2�rr7�VuPлFܿ�J����7~��:a����3�O��������[`�Z�3�d�H��v���I�~��x�ݜ�J���
�biu/�$$-������g�ɟ]Q@���K\
	��&����$E>�q�¾~�%lu���D%�8��*���%šw�A9[��QTꞻ��u��nd"��Ȝ�a$�cy��	b�h�V����-��Y��_�2X'���%t��� �4�`�i�$'M�G�[9ׇ1��e�5tXڿ�~�2�����Ъ����ĦP���xn�s� �ܕV�A��;7�`b��0$�Ʉc�*|+��+*=�J��� 5�~��C��&� �a,8OP�t�3�59�4fێt�v�sT�D��h��N��A�#�J�(k=l���97�U�@�,p�j��)���ⓗ�9C����c�	.�D�6(ĝa�ib��������#��>�B�:e�����*�ޔ��\���A;���E$K��6nu�K�qڧ k�qm�!��ӛ���<�euLa+�	�<��tT8��&b9d������D�B�J2v���ı�:d	X�&�>�?����Ʊ�-�OJu?��Z�v���l#kT���C?̼�(6;�/v6;U�^OX���T��{�E�!<}�|�:밦�1�9��3��0l9��Y$֝*(V���ƅ#EX��$�".��.���^���z�5�3�)Fu�ȥŪGJ��?c��,�Pf����������Y-f��ji���NU����.}�h��9��J% ,�I��R�L1&A����ڤ��z��Vf׋�`'��T��7UEu]�y�J�3�?� x��/��k���UW0NX�x�yS8fh�{�����Z&�(�QQY��M����=؃c�qx~{o���֓b��i���Qvvx�52:#�̐����U؈�z��Pq3�.�rn��.T̠��_�l��e�b@�װ��~z��r�9py#7�R�x-����@q
PS��L��@)�
�RԨ΀��d���`�hñ��ز��Ȯ#&f�h\����m[�K����:ɽE7��ڗz�v�c3~x������Ȧ0!`��Zo�7�5`ܭA/2��>��6�ЊU����aJ�]�[ĵI�����P��<tϷ�/��s�E��0�\���%)�����0�U$&i���Q\)�����2Z���" m-�fU��}cG�iZ ]pW,���\c��Ů��@��Nc�ǧ\u�Ȏ�D�ܴ�P& s�yjo.~�v"C�{�I��<�#,�0B���=W�F�n��ߍ�Z�
/��a�Uv*��U��Ǚ'�7Pm2�ve�����u�^|ib;��i��k%n��	�Ŗ&�F���O�F�ؚ�����CP���!b,ٖݡ��!� έ;@7J:�T{	|��:	��@4��aS�?3�A"�x�$l�b6�Z&���	�������R���9ӏ�"yj0��Sx֔a9'h-���!CՓ'i�z5��S�sZ:�ߓ3:��_��=8��h~ן���Tgt�{k�%�}�q�,J��4�/.@n$$ת�V����NA��݃�mۏ�D�HT��<U�r��~F<��y�7J81�g��Śq�MO�U�f�gL��y&����wl�G�����O�y���@:*�w˾r���f0�8����i����e�P�OI�1��N�I@G��ҩ�;y�����Yg�.���a�`T(VQZ�^���A�=OdKRe�L�x�e��n5�+�Y�k�t���Q�-� Z긕�"f=�gc��ߖ���a�S���`z���	O���8��x�����B��r)��5B8�ee��|YC�0�g_�7��%� L�xfG�<G۽�V2���.�ٺ��.S7¯��@�k��Z�4C8|�2\�E�pb�4!&�F�4��F��g��ߤ|5���):H0Ń�O$�ګC�����T������e�I�x���:( sS�$0�
���n�Y7��8�� zUѱM���Bu�z�,Z��~�����6"֢.t�U=���y��B���k����RW��p��"�*��6�>aǥW���+�v���~z�>3���@��>l�j�(2�@Ҥ1c�s�Y����:�����2Q�%�����CZ@�zKX�lq�ȈӼ}t��m�*w�S�j�>��������ƖT��R^\�g����.�G:jC��^40���K�I�IJ3�V���$'���_2}	K����������� ��ʒG���=G��ZGAbq���L߫m�t��3W��Nv��G�]�CտEXZ����G�/�r�8��B0J�>���>��U��L�;^�	҄��]ib�~â?9�[�Wq�S2Ј5ok�%ֳi��0���W��%��z��\���'c���. ���xȚOKU�l֯:~~�`�Kg��d�����<�*����A�s�{Z��+=&�1��ɹoI��xnէuj}�n�@��i���E�p#`BU#���I��(Ɵ��A�mJG���ޞ`_Ǻ����i�u;y
� �P1�y=�2" =��z�sPe����Iq�G$ 3��A ]C)����~�KP[��rw����`���Ae�Y�k�j�x+0�=h?�/_1�q�\��ЎK�ij��U}V���&|��J��_�������ұJ�X,�֚y1H��R��F|(�!�����o�T�H�����(������ˢ�=(��G~�"�[?W�BkŴR�����ٮ1(��Ϭ�H�����2K�|l�X9s_A�-9�PN�0�8x�}�2�>Z��+=�2������ o��-�@��sn]/9��V��&o�a�QZ��֮���c�0�s�i��*�������=[}XdWi3��H'�t,�p䙟�R��?�f[I6����C�_Gn��c]�r���G����.d��D�0�Uq�:X]�%O�J��Y���+���o���wؗg�yd�̗P � h�� ӂ�#��Ig>���EQ�~�$:�]�����M�����_��߶�6Z�8�Da�nd����E�WUf ^�!������CCsZ�w͘�\����+Ku�V�����H��W��u�z*�:�rݮ������b� ��$U�4���8�glمʏ�V�lr�2�o1|x6����pK0Yg,e�!|l�?Tq�������Íu�b�_5��=ZC�V0�0Ք�M�3�LXT9kNd<)L��#
��<�rՌ�ab���8����L��N��"�P��ZG~	�|�R�F�L)>��Z<9�=����(�(������+u���,`�5$�͹�d�P�ZJ�:�������"R�e�+��Ѵ�}@��:��K$A�am]"B�u� B=0�yN=_�-�1v�"��D�k��Ɩ��6�n/�;���E�h�Q^I�K��k�;H���t�]6 X�O���S�S���Xfl�c�H��n���=�����b�g^F&c�YMP� Q��yT���fnP:eU'-�;ة�.g�L�z���$,!-}[l2d��~L
�Ơ�B�x����:f즶w)�bT���n�y���yZ,����Dm�oZ�����E�N₇N��lܠ�j��4d�T�m�}���[�<8��A�z��q>k��js�|%�������� �4yb� ����+^����f��� ���N2�嶽rʆ$94��;�<zL|V,�&]>�����E�J�W���X�3�W}Xo�<�s��ļ�	B�'��
i`�����1	�����W��OGx0��,�nNf����˞���Lr+�F�L,���]dr�	���+�̉Z�P�& uum0D�! m�e����<g8�[~D�<�,�^Ȫ�)�x���2�^]_ْ��Z�����7Kf��:�(f�9�����[�Η}"_b�KZ�g�܌$om�:C��I?�?�߾�N�0r��ʸ���.�#C��ߵ��+��4�T�'ХY�"\
�u2#���]���M777lp��d�%��Xa�����ѻ����[k&x�)��"���"p�K�F�4|2�J��r�9?�������#/��/z������xz�p߽7���,���ޥ�������X��u;�wf�z�#,�:�\��%�k�}�K��	>�� �4�O���5-�Y���Mw��[/�����L&�ƫ���{(C�Y^P##�34�x�ۗ6���$GxxxH7�`���?T	 �}4Ηz�.�5�@t��@�Y�'��I/���R��>�0�g"ѷ ��QX�#\�V�~L)�a�/|�9�qӛ>���{�C�܏�ՖUn�1����hr��=z/��W+�s=��Z�/+I�,��#z.����s�@ ����5�|ʽǱ��g���x��BWP��4���2nDh� ��R�-�b9]P���/_���F�D~�q��~�u�N���D��3�a�P��D���k���m�����ׅ>��=P�ds�A���S�i5J1A�5@m%�;��I�!0ݫS�K�Kꉐ�E0�ܼ���'o�b���=E��Xl��eM��È��Aк�&S����r�ֶ����W�_-��1�tQL}�lح�oR���o5<wG�F�F��`��]g: ��I@J�h$���!��%�*��P�ak�k��a��#W���"�֚%$�tN�٠�_��Gˏ#�~���	 "[�Ҥzq)z��v���COYo���+H�-��W�s����o)��%��z� ������(sO�B�%��m�`��z�w�}�Ep0���}�]�o'̷^^P��a6G�X�H�4_��4�_י
�X'��I��1X��Aj�7i�b�E�����|��AZ�UK}�ӓ�3:ӷa�g�Ο�i�sp�gO����R�#�i��qTGF�HP���>�LsAy����=���m,���۹m��<b~�K
���ā�V۲��
+�\��Z&�׿������RS�)�7Z^	Pk񽠃B��E>�*Gꇅ�zU��N`J/b&P�\��W�6��uᅙ��o��=ٯ�&kR�cSƷЉ�=��%��>��K5·��D����H4M�S�h� ��/z�V�m�S�n�o�\	��KJ)?������)��d��v��]jGXѳ�v��(��\{;$�H��k��cSj}yQo���6|��Z�]g��>�h@㳦O���Ld��AA:2z���RI�'Cd��+;��-$��`�(�rhڃ͞��( ƙ�"�٘���V�z�{n9���^���j�Ƨ=3S]B9H;��X.p|�Ν��k���L�*�M���������9��9�'0�Zǚ0�*V�����G�63J�ȟ�1=;\̏#��˷u���kP$����;z1��;[e$Ѓ� ��pq�ۋ��$�$�H��<x
������gx��cS����+o&ϴI}�@)���1�_�������U���3����J=Ѿ9���F�9��9=
����]��R|z _4nW��U]��ŝ�R���G�[J����J�������O.��;���t����k򵋺`TBH����~N0M�dz���֙kY���0�	��K%�>u��hb���R�7O,���)3<�~��-�tT�N̔b�1!��G����T�篪�p3a=�C=�)���)�OX1�@�Dz�	W���U����}�3W���=�Q�+P1,��gi����і�3�ŒF#��egO.�/v^9<���z�}��M$���A�8?*Ysa�E.Ƹ�4= 
U%� ~��S	�GY�%��t�
@��}��;�Z�?>�� ��c��{Y�M<N���\���d�l�R��`|���y�`�BES\�CN=D�K���>�6�g''���dv��~-�urX��/��ҋ�/�S\�o���&?LqP��2��5|61g�G�6�~�D	����i�~_(`���0Tnw����Dz�%�:4z��>Z�T�(b�m:5�~V0X��S��F���@#Y�S�c����n���Ae��%'��9�?��4��D9bx���!1=6���H?A� R쁅�*�v�.�(����L�p��zۥ,���+i]�.�>�V�Y����!qK݄:�u}��@z�.n�r܈���= 42�ri3V�-��o�C}�R�r��ܿ����@�Y�F˘%� ���,a�~N m��&��_~/�ԏP^]/'�%��#%1�k�i�G۽������T0��@'���S#eأ�LL��  @�����}!��י��Nc��h��Z��,��R��*\����Bg�Ԓ�]}�5���B�n���l����_������������
�?��⓸55�FX�JN��?����Ӛ����F���gc��?I?b��g�_'�d}���Z�c �?����yY8ƪը�$w��l�G��.��J�����6b�QO�3��bے�������,�P��l�d�ʪ7���
L�/�.�}ʑ� Lt�)��X�1C@��t�K���@�'u�h�,�����[^���{L��%�窶�X���J���U3�㾩��1����:���
�E ����c������i4tp�k`��N5Xx����VE>�d�ҳ�r_Ͱ�e�(��-��HQ�*�G�	:� �w�5�fj��6 K^�no�^������1��*6VEA}ͣ:��?F0爥m�T����@����>>�ϒo�O���(/�P]��6cs�MӳX�gL��b27'������M,u�~����=e7�~S�R�dY`��}5��0�k$�5�����8�ˢܿ>��4>a��������Q{�#"?B�cݾ�,��0������+	�H���g����F�֡�W�������j ���J��e��RZO�BL�Б�l���$�/�������ʱ��O=�����
��翻�*;u��$)N	��Q��|�W��ȿ���Q����8��oE}�3�Ғm�g��S^PӞJy�d���g��K�G�a+��K�`U�p�ol�s&���ĵ���~n �~����=��A-3�����3 ���X��;��
9 X�P����V�:-��H�Ρ(��o����DQ��K��a���!����X��/�	���m50T���z'���� ��1�XT[�l�7;�w�z�~d����"3�`\h��|Yv�[�ZX.����V�z6�>Z�X��4��!�x�t4��2n+�,꣼�c4F5�)��#�\�~�R�M������5��f��&/�"�zf2���b"U+�G~\��^�0�����m��+�\�F�O־b���f&�/a���Y�yb�K��ۋ�U�������iN���͗�(�'����ﳨ�3IC�|�(��y�K����0�^Nb�ks�����$yȒ��꠫�R|>]�3d��~�T	�ru���Z+AKP��"�&�dm��z�B����'����'H��-�WQ��{X��O�\�'���z|����]ߚ���:��-4���j��n��8���j<[IFm���=ӳ���җ½�x;�3֣������לZ5��_�$=���&Ss�֐�f�Rr�lE\#3]f�U�ٱ����m��}X�8�������o�_L�/����K8[�}CF��:�
c�X�����{�Dҳ�~E2�K�j���.%/���fp�����qH�"�x.Id��C.XS5�юY@���Sr��yL�b �����#�j�-��$΄s���b	����+O�Fot�q'� �?귣e�.a�������I	�t{�uIU�������fle���^��Eqd���x�U�.�{X�A9�L,��AG8Ez�@�=	��P�M'�Ғ�wdB�;�S�[�t'��h�:[_�	��z�ԅa�[]���;:A�!����	�DD���96��y�d��<�^$�m���+zfo����C�X��8yHHH!�+�rWEX�vƜ��o�l9-ufOYO��%��ӘI,$p����+�"��̞��	:��v�r~GΚx�I��'�}Z��d�K�r�߳e��DPѶ��js���R����KEX���G� ���8� o�����Pbg�,�(��^�γ=�$��O&�φà˭'I�S�ֱX㩀��,�0wg�9��p����&����G&�����^`� ��C��=}Bѱ�,s �%N�l%���$��vL��M�� ���b���X��o�
��f�Q�I���z�L�~��'��:��̬��9L�9ko�#^;�-���� �۔-�o�77:S��� ���?vj�3]`�2O�I������Q�L��� �g���K�ԽUrX�Wj�)�c���Y�j��~.�;�9+0V����U0��F�y�A���|H�I �� ���6e��\:d������W$�^j)�lfnD��̸�˜�.z��{I><v�8 ҉��ن�X$�(g�8f�r X��6��J�P�bͶ:�U��)����G����0N0��w��J�oP/����K�5�?���m�e)ȡ����GYlG�V��XԩD����ʈ�!qE�ZA=�mu����&��L������̥��N=�
T��8}�����ꏭ�����-����I7���	�E�y(�u��!�:��@��ʬV��tK�R����c7:Wڥ��w���l�!tؔl���X���(fS�+�Ӑ���`I�� Ԩ�3���u��}ϊK�sp�~oI��v����`y���_[0)�� e�����������ig�9�xo�� M��2�ј��H�0�D�%�[��5N�xN�`��7��~�dʈ�<�đ��R,X�5�k����&�/����܈�GChZP�S
v}K��s�����˘QDU��Y�b�_;�f�'��=�$'�#�ǃ|&��W`���D9ee�c?��d�;�nܹH^t͡�l$�O��-���3�AA������td3��^��n︇�Qn�aĤ�8'�!�����p��9�,�z\��xZ�=�,|-���V2C
���оᜦ��dV\Uà]���I�AӫD`�?t�Rע�0J+#��AW��G&}�'w�k����ЖJ$��%���DD�\�X*ʹ^��'�:p��A�Z�KL5��QX����c��a�A'7՝��V`0�����+����� Q]���::��* .(�IE�biV���f3�~�j
8R�?Y)����ti�^\�Pe|��Ҷ!���\�^rg5�gm#�]��`�1��N�&�r,�y��0q��7�7U�ܐ]�?w�x\`�-s��9'$w���"��}��Ṅ�A%Zی�0�g'�
��X��j5��W��x�t�$v'��Qnhޱb�%<��4��e��ζ��#�Z|�F���)�Ⱦ��vVyq@��s��ݵA��G`�+��X0hM��V�}�}wq �8N����o�$��P�O�Y�H`�c����Nv�P�H�����N�R�y8���C�|~UW``��v���"0ڶ��]�q��i9��i���1o �� ��u�_�#\b��._w4i�J��4%kK��Qg^�֐]����D����ƨ<d8�>|�$<����cPQ��k��,X��������T�� ��������(�	���RO�j{n0V�H�g�e���Q?Vy}��ߘ��C_�lR��E��5R�R=����(��5xܨ��˦S-bl�ԧ~�E�Q�Ww����nzN���V_\�
�r��\�X'���z�:�( t�~d6�DM~�T�POf��� �%���6��v��d9�;�3�6Q/BI��Ɓ��W����X@M�u�i5�o���L0fE۩D�_Ä%��w4�C�n�v8�:���#Ť���G�:St�B*�X�����DǓ*�+k���]�Y�8@�$�4�J ͥ����Mn��1P�{�����~{��&O//�����J���W1���/�HU��L�י�t��iz
MX% � �xE����]�h`�a��FW��?-U�|N��j+Ǉ݃ �AfXQ ,@��������[ln�"k�C����B�L���to!���9��^�ʝ���p>Z��@ld�ո��*WRq�$Yjl>9ó�dI�;�����;�2Ք��=k�)�]:�9���
���>�����A7'������)�i��UQ��n7[/*�q����J�tp���B3��K26տby����80;7d�p�/�M��}�+wqzg��U>�<�9Fs[I֑��c�uT���q�T@��-1u��U@UTX�2^�U7+m�L3�y�)ݧ6NQ��Daj��躑Œ�b�Ds��k>Y�ze ����)+�.����������A�����a�𼸽;�B�*q �K���8%Lx��f�L���`��|����u��0�N��L���ܿ������zc�����<�2�d|��h�%Q?=��`�J:T�����
��R�o�`ا�EWh�dƦN}��	G@%v:5� o覊8�c�lƍ�	P0"0ݲHݱG�ݞ3���uPX]�C4d�=�}�LMA�L���I�X��t�Ӣ�qyq�{4��+nQ#^��ۗ���01�VWȤ �bt��`ME�{�Ԗ߉��<��ǼT�1��Z*2�/y��=:�}�$���tw�(t�`�Q��'�A�SX�}��uʌ�Z7V�h�%zI�!��QV�c���ȒY����h��vA�Q�O/ ߹�&*��Bфgb���� Ǜ+/�w�A�.f}c����i	�(l>uuP����W�d�zƤ��yk@�Cnl�/�T.0a�����:X\�A������	��.jBPG�W5Viup��`Ԩ}k��̪��k0��2A�=7�'fS����{խ��?��Km�e���Gz¹���I��J�R�T�TIG�%%O���Jm���X,fM^I����%zA�Mm��c�� �@T����-��)���XS���K�˳��z` E65�74��Y�dU����J��{�������ҍ�-��3�]�dKi�Z��=;�d��A���~H���r��$!�t��DQ2�!��7����e�pR6]PJXT8��lLQq���̌����. �>du|�.�%:$(�!�C�Δ�)��l�b��I�,T�ӕ��S2��:֤�υ���DDG� kXu�H��fu�zw	������ Y:�:�'��vP���<������J���Uc_./ޱ�:B�~�F���C���{)���f��(��bn�ܹ�����ý�"K1`��E��p��&�UuP_є�!)��f 8z���$��V����LGN�C�Az5F�z�z*�E̚�4����$�:\�lb@{��0���@�g�����)�\�b`���=��X��;���˽��}BO��-�0�%��2
�7'�r�Lm��v�# �ؒ��̠g_�'�e�ܛH���W�g��:��6�������aM��i�6 TFZ�XƪR?l/dI�i������G�[Ӆ�d��A-҇}�����խ/�"�2�}���A�͕ 6�qlE���oJ[��|Xw�[34���4�:��X��H��cm�?g�F��t��+C��ɕ@[��N����X��W�©/��db����vȀ?w�ۊaj�{�����OV\��uc �� ��Z*��S��,�{�*+>Y��)"��/�	P��X���4���`��#ú�D��YX�J��elā�-����pD=�m���Y8�� ��0T�s��A"�Lٖa��	 ���=K����PV��] [�BD$c��6���W�u�n&�,&&ºMgК����T��Rq�٭��~?��Ĥ�$̍���EϞ�:90Ҥ�e�Y��u���Iw�/�4�Vtj[�{����.\�,`@�#龻F7� �]Q߈E���RU3��(ZRl��F/�+���Ґ��W�jd��MP%p������p��p-US� �9x~�1�m���PAĊ'���(�=�Y)eq]2N ��	v �e��n5�#����$��$�1�J�X��F!�B	 e&����*�������5q�z�ሀ5x�!����t���_DՙVM�`�ES�mi��1��x�:U�cuw��X �>�%�S4|�� ����D�Jϐ�a�`�M��'Zu�c`T1�c󃻜L�{�������c�Z�B2�����'r�V���t=��"��
@���Fm//��O��&z:߀�d��lL��-����l���(PA�������S�}!�w����l��j7+�|L��#��(�SQ�=D~���8*3X��Š8ͶC�dz+Vpg�퓊��C�H_�|�@�΍D��\����X�R�n�G�8ۈ`���T431��]�"D͢�C�N~�u@b��:s&�1�ؾ�ќY�4�H�%F.�:	�'��@`Á��`��h+� �(��hYL|V_��
�~}^$��?�{�� �����oLO~���v
���P�_���wPo��zw�7v���M'0	�"�;TY-�����,�<iJH4�8..��|�V��t>�汸�*�n�R�B�KrۄD@(�j	l�"$k�L��óH�Т��T_n���S�3��d�@U��e0���3e��avfw��w=)��<�`� ��Mt�� 08�P@��`@Sp�`9
��@����l�R�A���P?F�\��+Wu�	�`��%�,�O�D�p䗊rp�A�eL<�2���@F@?�26��d�io��j���$��&؇�N�
|Ⱥ����QR���
 �)��S����;>��B���-b���Y<@F�Xu�zIdZ+I&f�H��Aԟ9�.Q��)�$����t5�'�F��;�O}v L���Fb�cɑ�B��d»��Xj���P�{3VZ��ox�~r�~�Z�/Y�t.a)Jy���`GN���cD��ˠ���͍��SGﴓ��Pr��Da;Ӎ�c}6���
�������r�tM*"ډyJ�*��K��~�
�b�ss�˔D/#�e�|4���>7��(�zU�A���� 
JZG�W���-Y&g�V �j�%\t��H )��ϋ����Jw�YL�^�0�����d:V�����n;����DB@I�;<bF�D�9Eܦ��l# �wʼ�J7�%�J��f�:��)}���[�<g�"׸`��5u�$X՗u��xŀ���% �&BZ� E ��T?IЫ����7-ߑ���������&�����n�����6H'����E��`���0.:����������0�}������A��-����bp��"��� �ҭxݜ�$vw�B�b�����D��M�f�;ҽ�9h��Fk7Ĭ/����K���|�1��1��%	��;*3*oQU]�	M�ӄ���hR��ѽ,M��5�{��a����u���K��ɑ\��y�O1���ܛ��PwXt#k�j݇�j�j&�2=�)�%"��jHOp]q�HV���t���>��˧���{���	,�b�!TŁgMҝD v�~��|�R����4>17��#G�~'@-�nQ`z��c.}̎�����6،��(8�� 4Y��흊nce�Ȇ�k"��i�-�٘/�f�.�%���-�.2t���	�݃���Z����t�U���3��p�uΖ���t�"�o���IPp�2�W�,��ى�4{�#TқT���*e�Z���Bi�=Sa��à>��S	�T�gD��)?��]���4!��9ݐޝ��C�1ۤ+IvR�ܾ�5Z�ɜ��\T�ߨ�J�e����U�'Vg�!��N��:�ߦ[c�t/>ާ��w��΃P�)�~��s-�&v�NH#y-^A?j�W��+Bt�T}������N}@̌�49�V��6O�^��f�l����YwV�H	1?�a·���)��F�,�����K�=l6˻���	���{'S�K�#�suy��$�_����6�I�򜲉���)TW�Th*fhto+t�������d9�zmL����:[������5�`{{�
�yD�{�RD<�H��˜�?�y>�܀�����_&0�¾��6z���M.%�O)�,� 5E��S�^�����A�Bo��쫨���%{@���@3�3��{�\��?}���%���O!	K�4P��Q�%	�.}W��%��X,�Mk}��˫jyl[`��>M�K��f�5�UAe7=|X<	L?�@�[�'!#t^��72` ���f/b.��v�řKR]�-��|f�kO�u��
N�2̂4``T�d��_��E�c����<��O���|﷢���A�>��ED����u!96R���j�3�7�W�8�:%؂�o��W���T��MY��{�%>�[��%`c�(6vgz��s&W*�R�a�"}�n���  ���	�=S�aU:I*�'P�ܥ�|��D�M�/?�i-�(��h�7]�/�tщ��	��n���d�OWWW���;��������1�C%d^ꂅ�h��PV7X����?��h,��U���YWbl5����苓e�Ec�\�^F,��$����]E�0ѝ�!À��� ����U!Y9#�w�;����V�L�8 ꢌ��h�Fź8��!o�e�/���tkC�	�7��Y�h�\]yj�K(W��ݻk�1�A�j
M� B#�樖澟긕��R�idU�͏�幰e��c欹� Rt�w{�s)�T�jA�oʢ����!���"��Y_��՘Wd0֕�ޛO(:�?�ްh���F��s�s�3�x�ߘ��DX:KXh�Ɂ	��e��u!�	Шm�y>��s��OO�}���[��K�8��f�>�$���n�G�T���G��S0�]9  8�S��ջ�,�� �P�_�i�L�ڇN}�s�1!���L�.�hˁ�IV!E��+5P�y�&=1�ۙ��b��Q��]B��"u\�����;��i"Xl7�`D�z����_��F�,1�+uwb�%��~��j jݫ�%��s�ԉ)1{�Xt����v�	f�{�����qT6L�A�WW���*�M��o��*�29���Z�{5(���~��*>ݖ��n�cƨ�,�_��q2(���D��+�Zn���R\�h��Ơ�	��F����&��ǟ|<;ū��������]��E����������'6J!l�:��
��'DQ��lE_NR��/����X�i�E��	�`��$-M��p��$�h�>�و����Fa���|�����1IMt��3�0�{z�U�/���!�g�۝�X��ؽJr�{�o��W�*_�ڸ6Ɗ	���M��D丠�Cm?1��-b�"�Z?g�^mk���ŵw3% ��*hRq���r*��;%B��<��uF�ل��4m� ����!Ys�E�f�-���o������{�_��#�a,֖#^�������W	���2�V�K���MfF�rP$���;�P������Fگg�:7n��]:�75)�I���S.g��j�g�|����% 5�� �ٻ��S�ygɐ(�樽�։�y�ό�>��?�g��b��/���>O��X)D}�\��o�^%��ͧsnU�b�ʔ}�gz�������L�B��K��8R�����8���ACW�86Ց���������\B�j���$(���A�]�`�W���V���؝�a0~��^)���;�uauUӳ.�_e���Y���-����e�a�� X���Rt��?$�E,��NU�wVZ�誸
�D�h�~��:r������@��ff���#�$�~�z4��x��R��g],tT�gm�
_>��_$w�.ʩ�������;.��+�ƅ2�}H��.Y]�Kc�(MƟG���oI�������!~��ݠ�M�P�,e�d+4X��|hl��'�"Y�0ܝ<� 	�������dH����D�������٦D_Nm��7�jh���BWt���2 U���NP1�Ө*�=�>��&b�f*��x��]� �w�w���܃��MmMR
Y��
R���ܪ�w���w�z�'O����B�lT�a�rޢ��HO[),y���x�jp��]k�.�&ˋj�ϰQĿ���n��c�4 �^C=�ɳݛ��tk�Q��V]��U��7�)1PIr3�6�@:Y����d�%��#r�M��P��)S2�l5���'[��N��T"q� �D�AAO�	Fv�N��".�d�� s̫Qr�)d�\nؗ��:T��,�	����3ǜg�O���:J��I��3�3J��U�Z)����(*��NnH�/
ҁ�{�=�K7�_����������'�	�(S�A��e2ݚ[���M�% #���2��U��QjR׃��ˌ�c�E�!�ԽK�&0%'}z�u�8���z�ޒ~w�����,�c  /�C(2�Q��{�n:��Lз�"�h=�_�_Ӌg�4��3��5[��今��q�Q���*:�����e�v�jd��������%������+�2��4PF���;h���^�FD�ܫ���z�^@��ڙ)����˗"�,�3Q�
��1i��U���ģ�-���AL��2��v��S���U�Ttu���ԉ�߅�
�I#���Y�{Sd�N̆���
D iY�\T�\��xœ�����E���������W�c���i�8�m������)��FA��)�D�����&'cz�mQ�sv_Y�a�4���/6�G��t�>~J_���������4�X�d�^!}�IX�
��/%3ը�|P7:���m'�/�J�4��rY���>�l�<�q.������bS������*�臚>�oϙm '㛇�3G�t�f(b��h�ׄ(�+�Gǐ�D>�IЫލ�'&CL�~���8HV"2!	�_��fы"��P��\���>�e�U_Ń��u�<�ۡ����D@���Y�'�&x+�M����B#h�������V���ʢ�vҮ;h�eo,�CV��O�7]:L�S�A�Q�"LU���Z��� �~��=�ʴ�C���-\�ڂ,����?��Dz��ӳ�B z��l��P!�$�1�;���D�/"����{5�D����B;�3�(d�4H;��&p'6�˧_������?uB�i�>TE� l8٤ϓ�A<UHj���;1�>��\D��yc5,6z����������d<4PU{��ިu���G��Io����2Ҹ�Б�F��5\ܛCs{*`"�V�®�x��9ZDf_X�hPYRh�}�XJ�14�����d��4�9���>}���]���4�T|��˨���{[�^�9�ʕq�ǽZtK�)�ؖ&�N<�H$�	����d�[q��������A\fh�^YQ�:� s���ɢ3�U�������N�>�e0�_���d�H0���
چC�b�ih0M<������I��c�@Y"��QRn5i���~���xn;������ƈ$'��0�':��%��/��p����G��\�������3%�J�:����I���*]7��D�'�&��'ѭ2�>��QU��0��������QX�C�L�pQ�F ����"8:}�����ޛ��m$I� 2��M����ε�ξ������RK)�ue&s7�dդ�R���J��@Dx�����U?�~1w�+��14LCe=&s�Ci8'C�.�"4�ԩ���pO>�D������B@x!w��5�	�f���k�z�j�mGo�+�£I1�j�����R~���45)f��czƖ,C�z�׫�vܱ�Em	��Ò�1	 R�(��2��К�:����P=�c�	�����Q^X��'z���X��3%
Q�3�_�}��x�m0k�#ن#���
x��캨�/�37�h7�*�b�$h���%E���CՇ�<��4�6�mU`��{��5����Źk9����=�Z��P�)����b~b�s��y���.�?K���f�5daJ�(ZU�g/���Μ�`�S)}v�'NJ�k.�:��gx�ue->�C-a��$�d�	(��0��z>�.�W>�̴��M���z�6>c�ׂp�8�.x{�x(�;�V�y��lrm��S7�Z�e+�N!��TjQ��ޑ�<wk��E�1���9�5r��p�B��v��z&X�Yt�`�!M=�ߔ����J5���0��h�mn2�8�l,Ww؏sm�W=EL���D�$g�����F�Ң�g?���>}:{�o���@g�p��lH�ObSR"&]������**�0�d��2���\�ʒCAT7Z���G?��n��E����5��K�,� ��M.��� ���,�?=}����콙���Y�T��a�u�8LZ	M�?s~�'��ĄJ1�3�󴧟���!7�����S;&60&�$�����S&�0���i��;�[;g��s/@r`^`��~FU��9�G(�cK���hG����	W�h�])�j˒H��B8�cT�,��>��3�G��Nc��`�|&�������ݍ.plXJ'[+��qmj�y�8��u�J���7o�ۻJ��A�������4�<2�O+%1:q�aG����L/=cO����~xf�)��'�eW �W
�zL1g)r����Z	w�{,�^��&��STIR�)�v�/]X�IF����u`�7jU\m/eQ�:[�k�9��}ǌ:�ʁ���V��xޏ�\�|��v�B�a�&��'Ǵ@�n�(��_٠:z�s���;�z2�E"*�p@�t^T+N���fˊ���:��|T9��o֌�l���ZU3�� ל�d��e�n;N�c��w�3��v++
 �:`G.Z��I�JL�!	6/`�'��kڱ���V�k1��F��t���������o�T��A�".�aR[�^�Xc8L���C�p)������]1��X�WՏ�8dt�����0$H�a�y��y���熛�9४q�&t ���k�GG�<����Ј����`���t�#y��|�G��J3��G@�c�'���T��2aA.;&U���gaޕ���\k>o�Ã��1šb�<:E�HG��ð�M��{���8T�@mf���?蟧��ǯgPe�~.���Hub��}��Co!���P ��P'�i��s)�����ߧ��L"�p����	���&��pI!��h���S^G�Ϊ���y�:��.��/�D�#|��v�+��S`��~����NՒla�^����<����//�"�ґy0�s�VS$�\���_;��&�g^�W0s�ѻP�

�3���_J�ն�.bx�vo<�8�d��||��4�:9���#F+B,��V�����2�<�Pѿ:Q���vo0g��v�y<�э5L����S�˰�VJ<��65j�n�*C�j5��9��Lg~��16����>Z�:8!SI$5�H�r��>K�������6�
�m���R���vj��	����Ԩ����������]��'�S�5�^�L��o1�'˥vcL)����ud��X���tޱQ2h;���v�ׯ^�gO�R��O���w��Ҍ!�ф�ď�;�=��0N�*[��ZX;%��O����R2��2�0䧧vM�=�Y��[�ؼ���}�~��>��|}n�i۪�J���l6��20e$xd� p>ƷǤ�*�(����sf���Qy�vdab����8a�R̈́�W��K���Rqo�g����{�4�[vBPb&tL/=�?e���g����{�em�Jx�ɜ��L�);eޕ��۰?�s�q��U|(�!OR��.T>���@m��&�`���j�T�� z����$��0D0�mc�R�!*�P�myS�t� �ٛ�>�����Ym��{�+���CJq/
�-ֻi$�b�ɸ�s�0N���NT".�>���Te��E��X�.b���=��ކ{<9<(	Z�g��*	;�Dv�͡W�L}N�\��0P+�c����+3��Ӈ��D�6�3�����M�!D��
2��.�U�ڢd�G<X��/�|�y���l���q�J�NI��|n��7z���������l�ۨ��`��.�K�u�E9)�]b��Ҕr�k1E���B�E\��r���Tjŏh;vdsvn8)6O�_�|i�5>�|����&���Q�*T؀�s���D1Ñ�By��ݠ�@�%���&e�yS��JZ0V�	
���j�h���.�o��������2i�������(�e��
wl�{�9��=�����<l�U����J�JY�!.1J�o�'��֦��p��Q}F��/Q)U�M0|���G���C�&��N��u��;����W���c��K�?i����;���'O���O���p24��o�æ��n�va<M�i�j8��S�B%�0pKer��K�ǂt���l��ؒ��-�J
GSBF��۷o�W��X���Ƶ%�!��z�JzL���2-X���H�x0E+aeN����J�a�ȣ3���雦�z�B4Y7�	������w�x�}r̔�C����eڠ�26������_�+���[���t�a�Dx���1q�J��,V|Q��!xIQQ�"O���@1��s���7�p����`����n�Q��,�n��\%N�~S�m_,�w~�V%`���O&<�6p�e'n��Y�Z�,��g��K���a��2k��wP�C����0�N�1J�4�DŢz=O:xf�Xp+#E�x,�5�f��9�F%
��o~�[��0�/��(�~0�����fg��+9ԫt3����j���"��̽���5q�]k��������zE�A���H��u�d2����]�����Ci�qt��������ϟ�b��a\����h��.��B�.]gN���G��K�Qa�L�N�U�I4����"�MY�@l�*�����%/�����_q�^B瘡W�mChw#+�rW�+��k(f��F
���Q��k�k�[�We�2l��S����d�o�b�r:������zmu��B�M��[$\�)�wGά8����[��OG��F[�͖p�+�IȈ����m������;n���>��c�m&!j�?��lp���A�D���&��%h�I�U$glB�U4x/�M@z ����ij?���{Ǯ�Ϸ;�,����G]@����6B��jM����G%,n1[��yG�O�Jÿ�O���)�0bZ��)x���і��SP������*o� ��؟���F�ڄ�1fK{��j�E{K���s�&���CaT������e��I��<6��[�8�mӳRb������:�M��Y�(P:O^�ѧ��C�iK�2�g~�%�/��!�pKwR8n}��h+���*FN��}f��y��?81<���h+�*>H8bnS-JE.��W8l$����qlJ�;�ލ���HZ2!z�J���d�1{�8��l����3�~�F�=~�,��%�~��خ��A5o�+���;��ޟ��f]�~�+������M��� ��������`4�!��QEk��1{6��"=����X;ULLnmY��C5�E����x�q�T
�l�55����]��J-jX�%	�K���#��"�x	�*�0��p㛰@�xC����\y�kM{Svjc=qq�g�`�?u�%��p%�Xت�""�"��wPd�}��w�{=[y�v�ÁGA�T��"�w4D0�+������w��і�y��o*8��=u��f�{.XC�h��'g0O-ܺ��-sN(I�j-L��N!�#<��!�ҷ�s7�}�7��ȿ:�A�Ӿ�3`m��4P	����$�k�޺ ����u3z՘��B	R̘�ߘ��EC~�s$G��g}��|S]P�XK����" �*�c��~�2ե� S��BL:x8�p���l�Q=�b6:���J��_�F�� g1�1V��%��</hK������<<�c�l11<_nH�IS%m�#췶+��>��{`��c!Y�*��Rk�3:x���y�'po؏������~g�fC\p�f_�d��Mr���.S?�h�
*a^���7e>�RN�B���X-��HoA�b1S��� c���ᓧL,}ʴfq?S�5qH�L��.=3�?�=��)���0 �ss����4h'�$��tol~��|����5�lS�獹k��yW���lH،޺�����l�����6y�ư��_��QJQ1���5������wy���ۑ_��eզ���߳��VȢ�hGl�S��{���f��K��F8���-F�p-*q�.�I}��<={�<}������{��/�L_~��e�Qr�J�2��<�`�S��״e���Zi[�`"<�H��x���:�J|Ԡ��Ʉ��LkNb�޿��b�=U�#'z����P�0{FJHذ��P�Ht�ʛ���'+���C��-��D��:����H�\F��lP��69v*�[u��!����X�H�7�_�`a�N�3kt*uM��U%L
g.�Q�!�8�:*��68.I��B��}w��Dr�Z���]�L�M߹u۸�[��Ċ?�Uw�v�9��s�9gs���d�@=�MUu'Q�a�@�MPR)�el���W�I�6)��2ԟ���j�3Y��3ӽN��-����g�����8g5y����Ώ�Lo^�v���T���C<�UKL��L�ڥ���|T��#��7�̆�^���~�5Р �?8!��S�Y8�Ņ�Ǹ�*����N]�P�3d�ǘQꐚc!�Ÿu}TSŚ��x�%f�w]`zx�%t1غ�Y����$����T�f�A�gIe�S���b~�<�~�,�#��%���Z�%�.���a$,ԦAp�whڄ8��C��rƲK@9#U���_�Oφi��'f��VE쓑����l��(CJ��Z�����9J�'�����Hs��,�A/+����w�]��/�79�N$l�M`M<�2$:6�˄n��g9;��\���75=��E#Մ�p��}h���1m���/����e���<�ﹰ3WEgN�mM��*����
��}/����[ń3��L�g4�a�-CV������]z���׶�pHn`�M"m��-�Co�zXm.���zZ��RqQMNI�@U?��"���F]w����<��C^�x��熐�Ȟ?>;N!�溼�N�Z�F���:V�Wn��<�iZ&��yP�藶2��.aOS
�⒝M�:�+}�+�g*�K���q3 oTmRDi��w,m�dXl�U��d�oʖ�)m	���w-��+kõrYW��"Px��f�^k��^og�w%HLob`9�m0j@y��뺦h���Oo���G�4���@�6�yc���
;w`��A��~��)�L�p�{�r�C���bx��6���
����j�GrA�#�'�ُ��U�B��d��sR�,	�����ca�`�.�aZ���7������E?��	a�d���t�e�~�16�Ǥ�K���/���-Po��T��x�v��Tl&�x��<~��޻g���a�ċ�XT�>,,���q//"���l�6�mL+�܍.�b�5�k=߫2�bQ��qSs���dֿ��ͨ7/�LK��q3H̐!�S<wHn��&j�4?$�c�~6,&[�3�
,��Cc:ۘ؏L�zҋ���a��4V#�E[x.k����16VQ'�~��si�I���j%����^��)a��i�{�f?��mO�{��L#z�j�[;c��F\Z�H�|�t�P��}���GJ�-�������3�5����n�����)��#`���dȌ	��M��$�]aAa'�2�b-�)��b��F\Na��ә'��8�x�lJ*���׾�*^G�Ս���d��)�J�FVJ�ŴS����ՄJ��Uo�U�/��=|�0}��ז8�P������p��O$��͆�hV|���I���e�+Fdk���
�_W�;?ӕ����ޣ��3-�Bz�08 ���ݺp�⽉����5��`�|d�������y���cNV7����o��8�}/��F���6)�A��BXH�>�<f�;�"�G��E0��Nߦs��e�hs���茆��,7������K�׳�X��В�ڰ��Δ$��Mq�~ʫZ�
��yQӿ?3q�g��~2��ɽH���յ#~z�=��0�²F�v� �����a�{�u���z�����I���H(�a)v�1��q�U�"m��~�!a�Dӥ����'���P�U�֬���	�ɫd��%�jEj�	�I�aP�8,��Ϻ����1<���khi�W����{@��̴�-L�d`	�F~c�w������}Ć��m�A��&��w��ϖ����K�{kT�ɛ��Glc��rs�0j�l<70�'�4Z� {zv���UA<%��F)�n��s�}�6&V �G�_�(��	��>#"0hf���86]�Y�?��rp�X%�kz�S��mx���Z�9.�a0�`�vPՅu��0�J_�ݧ�'&��Ffd�����}+,Fə��EV���s�a��K� lKZ:T5��|�O��ĠT&gGIQ�q*ȄOR��	|���&��<Ŝcbc�X�������nG7��9�>���?|�����H�{��f#��nY`dPSr�=lÚ�O�d�]k��Z���֚��ܽL��'�kQ~G��*�y8�_|a���B�?�sN,�6�5���.'n����;rG��)-��ŋ��ts�U!/�����^� `s���>H�MԜ�[;��QqS�@�Z����I�}L��v�Ț(�?:,�ș��%�E<���8�H�޼��r|cq}�ǄQ5��X۱�6��	Ɓ\Ri,�g�3#;FTP&����3�8��ͥ�F�H�lܑ����"�  ��H��~���ڌі�aщ���_�6S8#��bI��܇θ�x<���̛����;4F��KQ�UH�Q��6��a���EK�ԹQ�|P��Im^*D����|�	��n�[�]��L��Pw���<Y=��o��I<+�6�y�0�B���~��O�R���5��Z@;V�H�B�A�Ob�k�u�wo�y�0��b4�S�Dq��O�����We��8�^&R�s�DE�~��v�������F�F�9p^oq}a�<�DU�h��ydJE�� ��<Je�����������Ed�܌�������7L|J�}�I�mYW߳�'V�i���o��席m�U�)���,�]�q�M�;5�fS��׊�l������ʒ�^�aF#���[�vq�2��S&5I����Шs�M$b}�����>l��0��Z�,�LF��T�C`�a���٣=<0��`{������
!c^j��:��������&i>�qc��.�p��k�1yAʾv����h�!�Đ�Blǫ ;�5�I�%k������Z��0ʃ�����4*e��3���c=��D��%�D���r�'�eq��_A�PI-��r��R�\I��w+�fB�����db���L�I��r��f�>K|����%�Mj��Ϣ�	W�Ϗ��
��6ucݸ�[�����{�s�u�)�h�6�e2���S�H�HUg���DbIjRf4���c�0��8���� Ff�֫-j*6�s� ��n����ίt-���ZK���������u���!��`��6�f�/���<�� u��㨆�l�X���r���Ζ�+1�vM�SMTL�D=T%�ںcSB�|i���	"�ף�(��}��S�,�j�]Pث��F[sAS"��*{ڷ��ݴK�%��A���P,��p�R�t��;��2Z�h�->�35�n����o"|vA�:�G|��l����۸���fDL\(V�h4��I%�?���x�F���M����4d�;� �m��S�d��c����"G��d+W(Ai�27Ei���)�"kja�K��$(E׳kTeXI����;%�C�G�r�<P׿E��;��f.�Rg&x��
e1V����j}�Ɋ��|���Q1͎��~���_�9��N6�4�";��%���}���cgo�aLi�B��TOHX����S�	 �IjW�%	v��\pD������<7unդ�k-�k�e��'�E[�s���w�u��<`�HV�/������&pO�;N{Nɶ����V�'��^��?cM�I�l7��#�>�1��Nwb��[~��]�*�9���P�j�v�~[�������rx&Q�h�� �G�N���M�f�䖚;��	!���JY2�"�.�Ehp/P��b�ok 	����j��\�!�h��'�Ql�k�DC��jC��ŕ'���f�cP�W��c��p�.o��G��4��S�D�O^w�0��:f2����2�b"�}�I���.���6��:E�nx��}�Ml�����%"d�,�ua���Zz?�]x�,Aab+i{��X%^'z%��Z�v�`���ޟ�Y�!�Si�7[2cM0��p�"�o�ݭ��ǎ:S�r��s<�ݑ��"A"�Q����H�Dэډ8��O�ef&-lߍ�)g��I��1�x��تr�5�^ƕ6����x9p}�S)R�_F���߹z�b�`��\�*��J.���b΄O�1&�2	x����U\ۮ�M9l
�ﳤkߐ��ʏcPü4�T���	�[�ͷm��R����˙Y��3�j�`I��6��H���R�	V�(k�R�OSP���%.X��~�W��$���<�.f@�3�ro��ӥ�z���)3�{�N��f�0ɮ�cul�0[�����Z���^���k�̍��G�Fڢ�Hwcl�J~�\"�l%�F�ro��$�'�ؕt 6jb߽{���hW�{}���\��<U7�l���q�JM�d��L6�(����I�Y�ɦ��=5.\��+�V�^�����#)_��0̓W�f�ڐ���<�}X�nvU_A2�ߎ=�A��/q'/���!:�gK\5<��ʚ]���������	Ob"�1݄�o�gZrfU�P���M)�s�����4��w�)c$�ρy֢d`�vs��k�@!�Fb��pp1���ޫ���46�5�F�H�G'�{����)�{��#�Ɣ���LT<����f6��*�T���i�G#�p}0�ɍM�m7���ףO6��懇��/�W�m������R�Ri�Ί��9���a��I�vԝԻ�N�m#�x|�Rs��ʾ����YE�FV b~u5�Rm�=5�K\?�M7Ơ��)B��rR��
��[9��-U6ܤ׼T0j�ɛu([�6�IY��YO��/*OrO��ş�Bγ�c�O?]WE�,Y����Y���g���ΎBQ�iT��%��l�Zcb�&��p��%3���3r�wKZ��-ZDm�KP�*�QG�Gq���ӊ�js��x?0����;��'�F�unB'!U/k���vY�F��N񙰼S.��!L�Sl�F���l��rT�9A7�
�-�t��A�q+zc����Ax�8L g�^1>z
W�·�3�|ΎM�j��/�}�<�ԼD��M����fԼ�=p{VulU�pdG�<���ءOԣG�͓� RT���SR��Q����%&V�W��7Q+V":��ZS4����w�g�%��Y�Y}�̨;vO�*��$	a !�"������5,�w�qAn*�-���<FҥMX�9I֭� �"V�5O��%L���)��Ż�2�D��B$I;ϩ5Ƃt��O��
]�L .�
ɯn�U$'\y��x�tFYb�9"��uY�7b�v>�TE�G�F��yOET$!�h�^P��:������4���Xsp�rhGU�QI�ﶵ�L�����7à��$��B��0)��R`xKz��Sp���ɓ'f�`T0y\l�r�,�ML�)�dKD�ת�N	&�YK�4B�i
��p);�NI�LE�e^��9f�:~;�Ϫx6�������X�W�/�x�Q����V[n��U��3������rv)��J�E�Y3���d���6�E������~S���|zQ�y�;�S�!�ƶ^K}�{�{�,IF�&����u.�{�k�><)垟�z�~��V^f�>�)�.��ldQ�4�h?�_���_�S=d{�i�Q��sa�lr�`�n�k�X�*�]�R5�W��o�1U��nL�7�nZ���>�.���9%�uO�|bޝ)P�����Fm��H��hb�/��S�#�,�uAmqJM|��+�&�+��4U��Z��j�ro�O����g@!j��U��*�q�y�6�z�*�0����C�r�b�Z�g���I�W���3�v��R$��(��+Z��
��!�]���3�yoAj��k�P�JYxN�D����B=�&{���$�Kɮ���7�f}Jx����{7F��0���^24�m���9gZr�u��CJQi�Z�8U�b~��%c|kF0~��d6��X�sp(���cjf܅TV��0�p&��]w�
�PǸ�y���4������7��"h{q;q}��h'�Z� �?UAw�g?�e��^��s�%�;<������~&�+�{�q�M�������|Wx���^��bx�f
!��Y�08®�8�����l�'fS3�����	�RR͙����t�J*.D|�Ĉq �����5y��AQm�U���ĠSu�8��|q�cx@UC��Pc*�:���E�Ŭ���"w5M%�kz�<��|?��t�y��0�����7�f�����~{ZOa��P�H ��DsQT�L���h�����E��w9^{tvj��Y��������9�Z0�n�J8j�S�U_�]U��iLn��z��
��`�Eqvސ�m�W��U8����w�,�F��s�p.�b��6���GȀg>��Ԡ.���%�,[�t�+z��T<^�,I(�\��RX9�TmT��7�H�7=��G�P]�'��mR~4��q����v̹�L�HFq�$\ʒr���^�j�ɫ��W'�{��*|2����c�s>��6<���ɼ��Q'nڭv������Pog/�;�:.6�^�����6�E���2ڭx����7�_d��X�M6�<�����po��^�ҳ$s���ĈBި�+��7I������-[�%\f��觋p7`2�I��;�i��1NΦ�S���;��ݻ��j��?eg�E�':�0�{���ꈡVʗWw���:�/�$�D��#[�[���+�:��d�SYI�$�^�:hpb0ޗ�KpZ�-�&��m��Q�_|�=��/{Je�E��a����I��qcB��h�I;a�I�)�r�y�QUwl�J�B�y"�J�YA"$hQ��:�k�V[����Jδ�>�ݫ``V����c�B��D�q>֫�|>�n��uC��X�A��h��0Rx��P��>��;=�����7����sz��T^g���FŐ�,�-���>Ή!{�\�kܑ��]�A8�yŽ6�:O*��7ޚ��w�����a�� �FC��`�M��ʤ5�p���ߔ�:K���G~�e*��v��OE.��v,�M�W�aSI��k�`�\ֲJ��������ϊ=<:��>Q�*�B(������q3jb�Xj|R�����~,6�L� j�'�ư-�CY��LБ��2�l��5�5�)��O�]��'ɪ���?��\He�@JQ��o�,jw�-�����PKS�g�����}h6�n0���5�r<�J��vM
s镻�L5�rSj��������$d��2����\{BE)U����)�S%l`���׍�=B�h��驧��8��\���M/�����
N(SB1��:O@�x9Rɣ����vB`�)UQ��GO�~�����ѓ�셅<*�"W��!�����ۄ����n����hPe�����T�9-��$��Yh�I���_���ƵA�
�w�d0k���
[�bf얆Am	0��X�d�;z$��Ґz�0������wCyq���]`�B/���N�E���!Yq��40��y\���K�w�^�}�v�ꫯ"+�dS��T�`[�ɚoV[��2q��#���*��K���+GH�U���ͬo@U޲Ċ�]V��gR(q�r�,��w� �l9E�ט]�$�/7!0I:��5�Kżҗ/_Q��|!�g��Rz�}OvO�)Z�ob���g�R�������O(�sa�%�U�(_3��V/՝��m?*\��u��ٟ��Ų|<W�zc�aPn�@����i5ySR�jCĠ�L���Ճ�(J
�_�Ʈ��E!�H�6Iw��D�4[{����;I��D�̙-̵��q 78�	o�[OoM�c�'�i��H�����m�e��q�������8u�4+|BO)q)] �lǊ0kA<5UU̜�PØ���N0J���8zQK�p�����������8�2�\�J�HsD�x*u>��xa������~�"�4�9QЄ���}b������<���ׯ�����|``�V�<ЋoA}Я�s�Q��WlC��G~���#�ټ|��	 �G��ΰC?�=�V/���RƱ6��	��L�ub�U��~̸S�Q�)+w��o�8�3?n�Am��r#@�$������~� ��nnI�T��R���r�EYL�S�5��kz[�񬚄��G�s��q�|'���<�ub��/�=x���w[Fxjq5�������읜6�i�x޲���hV�&��V��*��r��"��m�W�U���
���m��Z�sq�e�ɬp�"�]G��lbyd��0�/��Z᯷�� �nB�[g�L�Y���Eo�Du��b>v���nb2�5&�#<5�N�?���g��s �-^�B}%�px���<b�l1��xC���}i�jT���W���j�#��1M�o����^>!>�F
�-m��M7�7Ƞr3�V�!�Dɂb!��aOE��\S
�P�ca���S��j�N�K�x�]#k�E�H$廇:S$���o�CE�N�~����$�U�(���z89	�!��q��4���+]ڽC�q6�[{�a�IMwd.lB����DR���'����D�]Y�w��3-�U-�m=G��楕 m>��	GkсpÚ�����&�=8�
�£�.��"\?�`0�� ��tR�~��Vx��
��q7��6�j�v�	��4�{:��(C}���o��b�Te��_�b�}7�F�{��������A���j�R�7��"�\D�K�qmJ �)ǘ$y�Y^OM�?�O���{� �Z�{�2�="a�k־��RC�-ED*�^I @��"�;��%x��"4��I�a�Q��t��4�\_�y��6�.�P��l����:�j0��5�õo'_4=S��E"�ײ�)1,ł���bl���a��R�ZO��*�RZJ�U��j����z_{�ٟ9d�jS9]�gm�/��~V}�FUa�̂�X��^%����h:��w�@�)��J~��w��4ajl�Ö��CR�~�Y����0�H"���{�"�)�w+]pBO-[��rj���/����\���䰎�:L$,]Ձm��
�w�k-7j�DqH��8��(�O>�?��~�Ǎ2�80	q�~\���x&�<׉�f���s��@l^g��y��Ք���e�)6W�4g#���'��O���2�-)�BJ*�!=7�����R�solV���P+�80���̸�vQ�o���7�� ;
p[ჩ�'&��<��ǆ��*�d$�`���ˆ]*�q�?�hi�}^Y�m/'Oԥ˺@ͫ������C�cf�!��{;�SƩJ�YT�
�R-UV�c)W�)B�\|�V�� ������"c���d�t\����^Q�ˍ�������N��L |��̉yx�JG�Am�G���+���;c/���d�Gl�P5��<Ø��g�7��Q����
�����ɍ�<��ۓZ5�-k���S�#���Z{�gۍK���`[y���̝�����Oz���Ԋ$Ƿ )'_`�āY_U�H��ϑu�&V2�U��W�^�&�70,���J�첉{b^:��ݰ�$�,/k�6�T�R�lO�����q���T38?N�'.8���Ԃ/r^�*]��`��6�BC�+<�k����z�Zo��1_��M��t��/
��Zvo��9W.������U�GPFDPr+s^�TOI^�n��#�`���X4��ꌋ����
W�f����������v�Ҟhܩ�n���b�Dz"�{��hj>����Ơ�$�k�;�����E�P��2�6�����4-�bM�NڥZ���)wH��HUkm��G���!�싁��?e�jng���^�6���8�g�g�}��r��0�Xd/^����B�l�7�9��s�}�����J7�����'�V$/<B�qe2v'FV��ȧ��<�����o�y�ni��?e�U� ҄�#biH��=te���ý��7N��3�>��c:���E1[���j��	��V.���yY�ʀ-�����x@�����y_���޽���7�C���G����9׆�T�[�dZ�$�����@���~b![9�"�+!�뷪�Ġ�6դ���Ę��p�NXxL�s0&%����>{o=�1��jo�������&�g(�c��J��l��� ޳�*�,�C&8J�h�ڍ]�*J�+o�b������������������*] ʘ��a6�yEA��qBx��ਧ;��сe�ONnY�6��0�K���	>��$XmSX.�{�̮�j¹U�Vм����:��5�E�J3���M{�N���l:6�N�iCԐ�lڵ�����%E������}Ud���Ko9��*�x;��;|���m�.�ZG
�v˚�)�Q�R�o��쪫�	���%���yH~���Qlw��V��v�^�6o��Ƞ5��R�sS҄���u��eA},~_u�x�ԁ�&WuS���A.����߇�u�ׂ��ίt|2��������@h�k�%��pG*�S�_���z4"�'!d�7�t��N���+[�3�;�����V�|�>v�}���kv�84,3ۤ<e�{�.#��zY.]O�������ac�g�!��u�ȕ���#���EB=�\R�����9|��m f�֨�>���������?�;�路o������[\kj[b��u��݆2��lx�p}�$�jӌ�Q��\q��I����G��4�!1�VK�r�{"��s��m�i�t��ـ�̞����u��ᣵ����vaK�~�Ѕ""����4�yd[޳�O��MK�i��'Y�<�=U����� Vu)$Eמ$J^m�1���v[��&X� ����Yb�aB�\��,$,M��6�m��w����6�(�x��v޲pV��Ȅ�i��m�\\���:�)���'އp-��1�Lh
}N�'5��/�z,�T���z�\�q��*�{���nU�M�c�v�x���A��]��8(K�v����M:mW�I�X�Ǌ�����$0�8L���P_f��Pkp䪜d���FU}�U�AG	�t�����6�tyv>���Hvdr��m�(��;��'_}�~����"{��-=�MԢ��ʰb�LP��ۗw1�U��l���^~����ٴq��ߋ�T�>�9��V�!��߷6����q��0��b���s��j�Բ՜����?��.��dU��]�䞎��&�j$\���Y�!�%�:�G�חe����*1E �d�Ol��d�	�Jf�N�yc�mjW��[۝C���ڿV�ō˜���U&�����JPO�G�o�ש���q�)�t1*\A�gfHu�Bj�F��}�'��L�,<׼�  x⻐����܋�Rnt�#C�	{vzf�Tޏyl�c+tX�Bd�&�R�d��ie�L4x��@�1&�*N,�J}Ҟ#5%�/'����n�T�K>M�^�J?��4�|��<Kx ��R������K����O���o,y�>TE^^Cm�qښg�t\��S#�Vz�*�<[DC����p�ɥ��!y-$�aPž�/�b��h4�c}P5i��m���F���"N��a���S�G>����-����Q7��2�*ڂ
x�yxC`��V�yj��>.I����ItR��zks`Ù�l=g�O(������{��Sp�������E��j��c��@�`��ڧ&�b���^R�����#�#��3�^']�gO�hp��$=�O.�=H�@H���㣋��]L{�����Ù�R��0�_���m�⦡�3{��/���fǚ\L���p�t�N�;�I!i�z{h�q�����a�mw�X�����w���w�������_��g�LFŴ?��LT�A	qc�Һ0lV�,$���Ђ:8���V�G�����6i�
L�0�g�b,^� �����QH����đ�/~�n�D+��W$�CD��d78M���|�Mu3�w)FDx��\�pA�JP�^��If���<��Uk¼dz��4G�5�\^����1l4�Ϣ��{^�z�D{�!�X��w.p=�ܜ��S���^��(�nj�qe~������M=~��8-]���P�)7�6O����������`5ޅ�^42�P�G�&�('�x�����nha���Yzj����̸�yK�W�"~Xވם��a(!�grl&�\��".L�n��L��z�g�0���wz��괰�3|��Q�߽uX �,����'>�C	�b��X�?4i�)U�!]O�emjF��d�W_��5+1}�Q2*1�]pQs�p��\"1��Bs��Е�z�z�,���n$�Wa���U�Β�ǚB�(M)�ISs�fPX0���NJ�M��Jx�/�-""�#i��-��:�\�R�SJ1��jGov���d�T��$t�/�:�cŽuQ�!�z�Fb��C�L�%6c�r�u5s"lD��}��ޠ�o4{!�<��˾�c�(���İ�XgZ�j�LL�a���`�Ō�;��9$���{�浽��l}kb��A�|"z�"ɣwk߶7��]c�o=��9�w������`ċl5GE�g`���M,<���򦀎��B��������������O�
���p97&U�>IJ����Y��[7����AIoN5���Ej�Z�k�"���"�V<�?��.g�0���K�Q`�)D�E_ʁ
Ґ�8
 �-�و��0sr#�4�J�ʣ��2�*a��Y��QE@V
J
�56tE�
-vP�1�Z��$����U��T7R�ĕ�j;KDn���0�a�����Q�ǰ]�Nt�OؼL�pI���]��-*T�.���-<ӛ���!�1M͍M^ͳ\2�5ljJ�v� �}ZaG��=������/_�1}6��w��0�n�~l���YW� |�}� ɂv8� L74�x���{lpWy��-*�#*&��F}VC�fN4��B�`�l0��JR�I�:�,nMa�U:�� �����>;;M��������OfP�{у�SqN~Z�	�Ө�_�k� �r@^�w?84�KJ���<���e�D2���F&�PW
<�2�B@��y�.���69?�v���$&>6!��qr��k���u3��,4SQwv�b/i���g�2������!�#����f�Sy�%I�jr�=uURt�M������U����z��;�pf��~���sAT��=:�τ�p@�G*�X���@����LM[���}��u�R�8�{��>�kR��\J
T5�v���h1��h�.l �wgI�?���ԫׯͻ�c!H̆x����VO'��w���ᙺ �g�k���h����֌�!'`%@wޞ����P�
�l��% r!����W�d��pC��E��w��� c�"�`���H�{��rE��'Ӽ���Ȩ2Mr��_q�Zi~ޡj�:�|uE>4�"���`�i޽wwތ^]L�!oJ���e�#�Y|�G�1�F�(�T���W�ԝu��ʼۊ��-�h��V�+~�q�κ�}�ٍ;��GAp�wlj��e�L� *��~O6��0_���&윛�#zhs�7��Ƙ���n%SGx^j�~��5XR�h���T'dZ#m�EO���7�BJ�~w�
�꺀��>�����
�-�B7��x/zWFJ��&ХI��
R�_��"�9'J����"�п��{˸������G��-�-�d�s㨢��4??��]wYdK~0#;M0�n�9��8���t/M�����Х*�l�4_�A�<RE	x����8w@)0�,��&ũ���I��}\�B3@j`�>�YUbS�A�y��(�*�a���̘z"o���4�f��$̢OXI�Z\��M��koP	�'+S�؍{�]٠v�(Ł��k�(���x��ݍ���k����<�B<��ܨJU�E��BA��KyB��q)|�e���K��T��B#�	���*!�揩�����W��U�����ͦ��Jl�/�7�s�%6������װ��5��uaaTG� N�g]�՘��Q����x���-@ ���� [�VM����V�������� o��}V�D�T��RPCE��J/ɹ��=�:�G�m�(�޹e�n5�ӎ�B��r��TE�'����&wG\e����Ŋ3�'��*����S�0��Wa����J���0 ����Ҽ��Z���q$������i��0p�&~��膠LD";����^  �T^�����c5�;9,�S���	cЧ��<�`/H*҄s4�F�_E�Hkz��<��6���ZkR1�ڄj����{�.h`� �������<�g��t�(R�j(o�q�c�y��Ġ��E"�,oV�������S��
[�)���JT�& &���{[\�m�Dx<�?�ǭiZ�t��cM9�Y{�J�w���31��Uv͂sNV���,��n-Q\K��HBGwS�v�H��9�:wR����΄5p�(`�|�����tMX ꫪ���:��U�at��8���4U3�P=��&�\����N..4U����c#�Ta�v^�
���U��hao$hJ���zA�B����X��i��a J	̓hs�<чDy�?��]ޅn�`��#A*8�E0ƫu�@ڲ,zK�nr%*��a�(�{��+����#�qqn���@J�M+m�6L�3'eƷ�0��{U�Ǫ���*�Q�%���6�
��__eoʁ���{R(�O�4X����`��S���{b"~��ߤ?�H�~��-�ќn6��ݷ	�C�Y�m�=z
2:����a�ob�
��E��%�+�!9�^B.,9����7��-w��kqm�^�
�Q0���0�)�ζWޣ=�{�ZbjGa���
��	h�	`�x�<A_D5�;h�����ϟ���kO5g�sohA��l�ý*�u��$�+x��Rq�:PU:w
�g�{c�H0����8�S�)T`�t�dŹXj�V,�7�ғ0ql:��C2������|�o-�K���8r��8IגZ�����o��h�6�aeЕ%Ji|�{�^�sP�����<�O���&]����h�fP�#9��Ul`�F"ܳ�o����㓉�h�RG��Z.���S��䕟Xa6a���SY_����.�<2������O��ܻ?=z�(=��K��ަ�O�7�s��]�֧���MS�RB�9Z%�DL��$8y
��`��6��S*/��e]�������2�OYk�Ja�mC�=lt�l50�imF����"���@q����l��C׃��
��6$,$����F�꺡����m՜�R`����o�ۻ�q��O�Q���|g��/�������o�3�N{�Gg��y�6L� 3U�T�I�HH@��3��ZK�ܴ��y���N	�u[y�Pn,xň�i�O�r�AŸY�r'9�Lu���z��դgޚ|�]��;�� �Ź9`@�oz_3~Sx���`H��j*7��YhU���Z��2RJ�qP�G4�?7��(�{�_����4��ӎ%a���k�T^�Ҭ�$�\���[]���3��<1i`���k�L�x�grc����u�I��(U�5�<0�id=�c�;O3���a}^N�IYڑF����Đ���j1c�>����ݹs;}��7V�䘠ӆ�0>�}U���v��P�C4���ra�/X��zw�	su�;oYR�ز�j�f!��u��`{�^LhlQzZ�<i[n����S^��j�։�L�B<Vc>{T8�����h��Թ����0��9+����,��c��i���e���R�=�(�L&Rӆ!GV\z����rVG�DS�bbO|�!	ѱV���í%ܐ�B��\8�!5z��;���X�L�9��*�fj���9�h���r��\��,)�p�%8N0Rn�˹{��U�r����_�A��J���r��
S9��y��v�}�:�x '�7�_�`��9�C�[&���@Qj�-[
]�T%�v}����4�Q��(k��\m���*G�l�m�IE¹ÐY�|�C�νN�c��V���a\Lggo�0�B�<!��<DE��D�����O���u���$$ �d��+M5Y��Ջ�'���r��{D��5쮬���p b�M�L:�� ��|;oB{��֣{|v��Y��Ng���ꍫ�Şj"�綢�.��./����#�DU�UL_{%�bٍqO��tow���:����b>�1e���b��}����+�t��}$����i���U�R���ׇ��L�o?��X>����6O��YӲ8y�x���w.�b{	N��a
B��O��	%����5����P/&/�:����$
�4����2:��%?A�5��{%7�?P���6[Ye��]�<cGS<����/~��� �u�XQs ���<��Q���� �	j�J���;�u��^G4�n�WQ�ޖt6��7Z�&��x�'%˕_��4��T�hYn
5�w���=zDZ
�31��4��������DZ�J	���M�*�)o8�i+;�#��sM^�ހ�Q\�^�	��R�21��D*�yҩ�V��IL/0��W)/7g�<=p�[H�ݚ���Z�}�)�CyL��v�?�gD�f��lg���9����Ժ�hL�����KE؏C���%bk��_�Uz��M������y��9������=KK_br(�3
��a1��^[)T"N���(��B�y�z��Ax��B���6����{5x�Ą����%��y��!�ٗ��'�WyA�U7JT�.�ӷo�ح�wݝ��Ի�A_�~�����$TӀ{���FUE�Ks�j�q��$��,t�a��7�G�2��F�6��ԥ�ئpI.2�s��HҸ;�"��,Ř��I��x���:�PKx����qbL�����&&�-����x^P�,jP?o0�-�q~^J��.����B<}W��6Mk���hH�Qɭ���5�!?<ҵ)M)����ս�Zm�1�����sZX�&�Q��0�!�����!�<�z�l'ˆ{r"yhNEvTI��w����o�����8zN(LT�(B�(8T���7��"&�š/RKt�N�|�T��ABO,}�J��FT��ƁV�b�[ے�U��b���yy�;[�R~�Ƃ2ʍ��&��ц��#�쭫�7���-��"e
M�$`Tjچ�a8�\��c��K�f���uS�A�A?��t�*M�Ŀ�{6_}��e�_�|e�dؐr�R����v���;�ǫ8?*�Zc��;��،0^<��	�xIH
ѓ�鄰H�A�B�(���<���y���&&=�a��aˣu|����?^e�k��YVF�yw��mD�ztˋQ`DYߏ��g:���b��m<����͛�0�z3*���2+̌`��;��&B�7]�?�۟<^�� Y�^��SV���~�B7k/ݹ��Ixqp�ݽ�~C��R��8~0H0T��Ȕ'#O$�4��I,pI��Ay�v�(���f�|��${�����0끥�loa��I�]��S	ݎ�P��eN�̭�QGfХZ��Lەq]�����G.���
X|������2�$$���G�����{�L��yX)�P?�0��?�ɩ
o�#���t|�B0i��m.���r��K����N�=I��zw�E�Bi��M�ɧТΚ�(% ��Ja^(��<�=G&0�w�9��CpO�F�"�*��B�a����E����E�6���b�j���cP�E+��v���i���!Й6����f����?��?X菶O�=��P`���g;f�#cE���+�����r�����5�|��D���L��<��(O��CJ-(�<X[��^n�G�����s����T( �e�7\�Olb#1��e�F
�1�/��#S3����_���4b�5�[�W�[���s��K�7�E��1.v��{u�D𘞟׽�0 G?;��hX���{~�s�_�✒ޮ,:�0 �pː��=]��0Fh?��jx������g��Ma��ig�;c�
��rCq��h��`^㊨��X����Ն��=����߽w�q�c�d��#�h��	�DTq��O���Ï���p�&Q�7Ƞ6�����7U'%s��Y���B�-I�T�A���B*	<��s(h*N��Eě�篫���\�	W`Kf��Ӷ�̆�i����9����yb!�w4�����'�[�{V,��*.T��HR"�ڽE3�ޤ�	�ͱx���y!�Px[[	�}�H�߻o��j���dH�Y�%�d�	w���k���^�]M��C@�CG�=3>�`� �6��m�x�������#]�;\��l�2e�`�,��6�bc�!�*J����kCD�g��Սd�|�9ᐧ�5W#s�R�}��G*����-з���&h���g�����D%lF0�Pg{�����1���N���~��}�qﵹ�Pׁ���F��h�P[���cP�(��0���O�WOEy�>�wL:L*,�[����o~k����oӟ��'�B֕t�Pm��6��R�J�KI��'u�D��sZ�-Џ���+�OQi5�ނ���P9�����z���{���_K�?)�0L4�4Q~@�+,��ņ�3��UfhF�8+�<�� B}��{���
DnT��$a�%�Jٚ1-���"������{5l6B��ɻ�.��8V�������1�ϛޫ/�2ʸ���U�J�MBq�;�����x1�K���Q8�ko4q��ub3�����D	i0A�E)/���Ό,6`�0����c�=A F�b+ ������̾(r������庪���0����6v%"�)���w��7�A��y�Ch�68�й�j���׳��!ɻ7o����~={�V�\��۷F�ί�?��"�>a�yڥSORY�(�
-�Ja�l�1Zs�{P�І��t)�%�f�l
)Qe�,�D(n�9]�лA���}�����бVSg�=9$K?yl�
��#)L���qa���(���b�_5������&��P�����o�И�RVc;~f�&~,���Ȩ5��y<���6��o�?�`����D�(�K�Ԉ%��#m���ͤ=Ǟ�t+�Ɇkp:�U��$��Q�tx8�I�L�Y8�d7F��a��n]H�\S��;������޳���Q�7υ���9B;8r�C�&����d88��qG����;���cP���M�M<U�Nޒ�0�/p�	�?��<-��������e�����n�S�f���e����Ј�V],6k%#ˊ�cb�0�H~]Z����j)������>���ԟ���[;Ef����]|e�][GOD��
;�Uv&I,[Ki��s����	0>����z��}�}*-U%�F`�'��Jm	S��z"�C��5ɬ+��%��wGl��2�����d7ěA�0�
9ȶ��S�x-����{��/���hRo��l
j��H<��xNO����&���KIʞ~��z�(���\�x�o�^�J
��}bn#Q��	e�p0���b���.��B�ɸZw�����+ɫ�0�����d�&��E�.�J�x�DIW֓�*װ�]r��7B����gT��:�?��-�׃Uz��A�> ���s��Wc:�t}Qd�o͞��0}԰�����jŅ�W������0��33p8�KXD#�i�X{� �*)��ێ
GH.@��ڭS	��=9�w ;��������[x����;�g�
͞	�*��j��JDu�?=�֫Z.�=��6ݵ#�	͸]Ysܨ�Ԫ'o��B>ٻ�=�Бq�j��#�k-)$����G�)�S����6�Q�7p������5I�	_Bo�c�65@�|D$+���Ӭ�{ؘ���{��m�v�;�w��+�l��� ��T�3]������Z��c{o��aH�x�ȼT�tQAj�p�;r�c J{�͘˖j�K���X��8����^�R����y�G+'�8�1�������}0Hv�rb���{������r$�/�ͪ�i�5UB)�P�_F�"%e�z����H�٘�C�
�9A��ݛt�ޝ�?����o��o�o�q\m6�6)� ��OG�|�훅���5�yo��;�6Æ�Of���	l4Q���T�Q�jҡU	� 4�3U��3��x�s.�DY6pS�:��� ��jVwe��.���(��n�����	�4"���s*CcڧS�����Ќ_���Ͱ�v����"�+n��?]MV�siy�$]S~k����� ģ��Z��O�����6Z����o����GG�4��"?T�U����0���M�p6�V������ĹےӜk�'���
��7ժ��+��9�D#��g���F��H�B���mJm���=�gt2���X=fщ�s��.s\��O�c�0ui߲i����֨�X��t��\C�����2McM�}��/x�"j����C��򸊞Ex�<R�Y8/Jr�6�1���,(.b�?d�Ł�bgK�������lg�}��'�(R�ԒOx�̀K�3�}��g�^C���g�k�����J��ޗԃ�e���Z���t�s.&c���	�⼛1������R8���gr�H,8���^WG%
����4&]��@1vp���?��fr(O�*�ئ��dq�h�������vO�o��(Q���i�����2ݭܢ��q��-�Et�%o�6�N�Mj���M�!B�_BBf�c��z�ZO����@�=���{�J��{	!n��Q�6� +�IHl(�˙¿B}�;jD�aj�]�O�Kc�Z#��Eڏ���ROe����6埀~���`��G`v��ZC��Ғ�ƅ��5����{���%�U02��?H_�����������_�5����_UF��j�k_�Lp�ը�j��Z� ����<#�W�joi2E�+)�����#tEk�٘
#�`\Sb��l�j�Z��ވQc=�$���>:\�[z%K39��	ߊp�����]q���c�_����kO�br?�Ǚ^�f&ּ�rC�����A P�u�������Eb�d)V���gڷl��U��@����%�i-ڶ�	�e�[8��)���_3���Wڕ$E�7f�<'
�絨�뢴�$Hz!�7����:����"��J]��ds5��ދ�Q��r@R��?u,x��>�X~F����h�hV��a��z�lf�U�X�(j�b1 �����H�߿����[}�^�����Gs8��P���b!Hl�(7[�����0ޓ�)A%(Z��b`I�I	�m�OZ�0RV�;�ί��k�s˳�_͛�Ĭ�DOL0X�'LR�һ4F݀..�]�J"�K��3սC�:r]R�>_��
c�q��T�A�;�O�4��e`�|���֖��K3�B��7��0ze���{�ڷ�y�P�}���~g�:���cM�p���fyiђ5�$S�
P�.k���X#*�f�
;/%>�N�ITCye]�C�Z;���ڹa��bc�n�[Um���M<n�Am=#���تވ��Z��X5O�]��a����*��7���	�>ThEc
#�	c�P����e,�9�R�O��o�$ͮ�9u�!��^ع�ih<�D꾰,>��g�:����$fO�����wFچ�P]�ѻ�ݠz�еi�L�*hj(1�������ܛ0o�~��`�Ô	�����r�TL �!s�B�yS�#x���C�y�����ӷ�|�I+_$��&}�w^��MN�a-�"��v�]0
�7�%���<��JAckr`�u�ƍ�H�x�r��~���5 �r��:�R�f�^P�x<:5�pY�3�b�M�Z�zŘ��������4��y���"y\���,$%e:
;�uǸF���~G���H����/�w�}�����K���7W�G� �5V$Kwo����ڕ���)|�Ih�j���*%�r�㛦�f�$Y�=0R����<��!�������IƣG_X������^S�7kH/���}K`�h �&����/mM���x�M��@Q�^^��x/���Ƅ�O��=�k�P	<|`����¨yҙ}'<�#J?b�R�ͻ�F�ÆLr׳��Qɨ��z��� F�'o�۫x��H!\���^�djǤ0��[�w�G
Cz�$���3U߄N�!��d8�ttγ���Vc��Ka����o���r�,�Z~��+��"��NO�V�Ԟ7��nX!>�CO��9�W�!ҟ���e�/X�hd��k��y�cҾ�ohH'����;U�o�ͅ�Ʉ)B!#KO��!5������޵K�#C�+N�=fh�C�L��1��e\)��]��:��5��r|������/F�n0u��]��G�@Uf�=�M��JN� q��L"��1	H4{|�N�f�?a߀[Vf�����6��R���j#;�"��݂��nj�+�����6�6��>�Wz˽ҁ���h3�f�ڀ��@r]��'��M�1MW�����<S�h����R�˶eK,��I��|%12�0U����9i^ = ���W�B(x�0Z����!P^�:��3�m�Д�\F!u�V	�����������*����dr)�۠a���]И���KW��\���I�v!ͽT�V�|�p�z�5�k� ~mƯ�*h�-�N����ռ�� �@WZ:���%�`Po����Z���x��ٰB������%[�����ʼAC�$-�d�e$�*_���MY���M���q�;�cd��-nQ����J�����ʓP�6a��=�7
%!���ަ�0����%cz�m�1��Y~�%�7/���2����d��0���8�&��
�*BD/,�3*��0��~5� �|�浵PA���.=}�Բ�;���>s���_o^���@�W=�̫�mnP2h79YI�U�t|h���*�wb��;s��PIBƙ�.5r3�j�{���w":�~�)�C)��g_W�mޢ��k&��R�cA�+&Jl�jAmUh[������I?���h~������+�T�	0,P����O����|�Ҍ�AJ�7�T�ӷ*��B�TF,Η�_֭�� ǶW1_�}V��h��œ��ֽ;�X�z�
-�g+m��uTS=%h����{ē��5ƴ�q��xjT���6�7Ƞ�kC�@:B�O�E�>�8(�lm���-���c�SX�h�p�N3���p�������`������i5H�\����
��)~b���;��(K�Փf#���ڥ�(�w����a!y��A���}�20��j.}zI�-˅�D�u���c��:�iP�0��T����!���8�� 3���V�'�8�``�%�O�������Y'譾����_\�~hM3��;����j.��{�g��ϱ�^�l��O�ܟ��.�F����(tk�F݅�ԩ.���	B�0�V#�)���isC�ƴV��V1��������Y�sZ��;�>�ZR��G�����(,�Pҧ~(2�^��,,��B������	���P`k����}9Vx1���y}�sM�FH��sϊ�Yc�8�p����͟S�;��T&Z��pXGL�\"$�,>k���_x�<D8�ƵR���n��es+w���"X9u�U(g��F��*����0�y�n�0t���W���w���'��7`VP�����A��7�ҳ�k}��Mzw�nQŤ(�V߱c���a�G2I8�ɉ37�8:�B��rܦ��r����վp�S�tߔ`j����t�j��c�C]x��]�u/)�W �����o��E����4�n�u�N2;�n�Bd?]�ɱL|��@%<��t|�R>~��� ���/���T[�'][��6��K;�(G7!��e(D�&y��0אmɷ���55,� �����sf��ɞ��̦v�Iy�'V��#<������k��:����BX�td��	?�F�FH��@�6P|������j҈�:1���a��䭍=恵�g�p�2�Α]���z��15l�z��)d$@����>�Wy�"�c�Q�pӈ�TE�"�������Ԏ�{� ��}���|��Ij���~+M|Ѐ�Y�E�`f�Ҋ��37��$"�'{��~r"Յ5�Dp�Vޑ���Ld��l(]�ךH���h4�ب�V;����ŝ;.\m�k;[��T�Ǩ��z!�'�j7J����������{&V�h�i|#{Oc9�/�S"����71�-�^rd._�����&>ޜ�;�5G��[\���]ӊE�%4I����1�|l,��}3F��_��lW�dj��<�ج�k�l�sr��w.�F� 1C���ѳ`@�"�S��QIϒW�-0�H8�3�׃�Z�
��S�s�x�I���[kw䚡�׍{d���uO��KY>Ӹ��ק����^W����d�(u�X|m&�[z���ͪ��r���[{\����rj�?�,��d1s}ng%�u�F���:��<��n$/^��h�Zbi��g/uϱ`2��/ɚs���x��ku���e����b�,-�-芘�~R�w1�"����]��W�����80�k�^�x]ȿ,����~�;��׿ɟ�5^�h����J��F�KMի��`�0�d���ܲآ�9!	�.#��0{�ݡy�uS�zQ��j��'L+���u|��������b�:Z,��fA}�Q+!������RA���WQ˃~H�A}\��??ZU�Y�J֚�*�s]���ObP+J���TOf��3���:��Liʑ�����[��k����M8��.�t�J���/<�qa���)<]��&GNi�K�ԉxJ��c�ghiOբ޼ky&�S����\]bl�,�V�Ҁ6#��}>����3$���:���L����-$��8���+�{�w׌g�E��z�u<<Y	5�����qW�NN��O�ʧx,�Ѿ����{�O�W��1�4K/���ㄟ��R�x~����>�[j<�^�^���9W	7���	����bQE��;͖�9�AW��+���'*�TM[C�+��D��j�R)1�fU��Tᕖx��A���^�A��{���٤�%����a��4J�`F��W��f�K�W��y�{b�횊�Y�'�S[Ds�5�J6��0�%6�=_��������'�Pm`��z �RǾW�>��Psd@��sb��)�$�-���RY}G�Vj�<�K��a���ޛ�7�3Y� )ٹT�=������t��k�tZ"qˉ��,*%�2KQ�Lq��XP�{�4 ��:������U]X>��;���(�K��^	��Qt`��ud�q@�߼��j��zl���ԟ\������)4�
��Qk:����e�-�-�]R����Smwܩ�&~ߞ#�.�Nj�r��uЄJAvJ���	a��_Y��{�8��z�8#�}q<��p,�!�~��,GY_���u���+�d���&����t|�\���:vrU�r*h�h[!EM%����E���O�Kd�͚Q��O/P��t!������}�I�9(�SK��]g�1����}�`u�1J�!vΨ�6�t� ��Ȥ�s��
����H�CV���Mg@3ߤF�>_�-��R��1�J���4(߰%���أ����}���U�P�p�d ��ԙɠ���2c���N��;��l"���J�$����@ 5�A]����{�紏���2@�.F�Gr�f�Uj���A�u�+��'ZB�qأ�;RJ���7;��c����̼֨�9y��X��RM����1q��pҥ����M5�66\���P�M�c��1���P_� ��>̑�|K��i�Ώ�9��65>�y��M\G9U�<~m2�[��g�R�ժ�Z��}����hTz�UU�p��ONW�F�Ix�N��S�c$jBvM0��m�AU�!�������18�lr�D��f���i�^:lL|��N;FtVOY��n�҂X�tK_�/KS�J��Rƅ'�4gt��Ih@=3c��ҹ;��r�0qD�Jn{
��(�&���r%n�oo`�`УOri��lg5k��[���Z�pPOA��%�ɭ���_a���� U&IY�d�Ԁze��*���И!�[#���޾�$٪�)3 ��؈�z���m�ASO���PK�NI"��C��N�A�pܴ4�~�cZ�EV����ڱ��j�A����T�crNH�E�WTA���R���`C���ou`&]J�:$v5Y8�0�d���:����Y�Ԭ�^;������ ��
�f�����xW��NT��}ä�԰��2�c�<���P�.4:���^���iXjJ�d-	xX��Q[��C�Z M^��Y�+1�媶�4�#��]*XG������e�r��!LX0��b�t���y��@�GJ@�@����ݠ��y�2i?$P��YU'��`M e�5����LvfU���z�H��͞4�N3q��X��v�����q���֜�~��Q�`�; kig�$ޣp��Z������O�4��$e�	���C��6^��̯���X��o���8+���LTt�P�s�6f6+����78T�C%���[��2Z��`��ȧ�ٖ^m4�ڈ5�+�6�V{s:���yx6)P1yV*DJ6�io��g5~9I�����Z�]��HF;.��!��c�۽�P6�d��Z�R ��e�Y@&��h(�Z�A� ��r%@mfqt;�T��&��o�#b�r��ג�������R�]f�.v|.I�ɕ�wp&�#JKz�+�
�Y2�n+M2s�'4Ęjc	6V�.3���uI��A2��@'�`Nx��yg���'>��%��Bo�R�2Յ��&H�!f��hS �:���P��t�� -	�ύE��],��T�ЇM��ߜ�*�@S�w�+,=kU{�����}��bs唣}�=�����&�r��<Y��C|n��1%�b�ި�x�Vtƙl P��5\_`Ș�WD[���OlB�ܒ��D����r��E ���������i�P���Y�h�Y��A�0[�l@n��͜&���|�KϨ���N�Rq�6�\_�׶0육Ί&\ܟ��>�Վꀚ��
m�P�IV�ɳ�R��"�	�-`]���5R�������v����p�2{�=��g���eC+���:��n	 �F+��p�	f���ن�F��;tUt��3�cϓ� ~ڈ���~��V��.��Pg�0��Hy���^9�������\���A[�~̡a���REx����9�C�9o k�0 o��F!�;T�G_��~ǿY(�����nܔ�(v���Z����fך�jq����)_�R �&�^H��:x��0a��+)����VC4�R��:�&#K�Q������r5/?~�!&*�&�h��*�+2��v���EJ2o��k�=�4k$�lZH�\1��=��Δ(�7�63� d@7���x�����,Ƚ�@�)���k���������OR��u(0�z����o}�7�b2,C�VՁzO����˰�[y�_I��"�@�]1��@y�2]�X�O�����,��ǓUQ0�g��ʞ�G6�,2�m�S���ơ�A�f�ژN��I�Y<�gO!�^OY�d����-��3�ڀ��5���{S���� ��tft�Ȕ걯�f���f�چ��3��}�R i�P����,)�������Z'4�7��c�Qz}*i�Y�^B�M1��A.�WΏ�7[9ڢD-��bFQ��9YJ�>Մ4����D��,���H\�	o���9�y�	!�k�c�����0����rOr��R-G���@�A%�a�M�)���χ���Ս�Aƅ��)��nk#���-i�I��uP����]�G�^٭J����X���[X����V�����5�����M�N(��"��h'^-s�|�(3�I$��$�zV��a,�loϰ�k4_��̲'�Pwk����@@d0�%;Z���/	�%����u��P��(m�����$��Kn���U�|�#M�����99C���4ci��n�e��
��)N��-8�)�u�a�03O�ɖ�2���-]�;+[��6��(��铣r����K���ͦ�yf��ɲП+�
#�w�8\?�;�n���#�\y笉R�`��!b]�JB�"*g�nC�8����Xs�fQ���뵣��a����4�2����Z��>�y	�U�ո��i<cW\լ8!�<҄Q:���	Z��@���P�o4N1D �% =���FJtvV��T``�gŁ�~�EX��;��:П-k�e�	CHh�p�� \Z���]ʊ��}��udt�l��?�r�_<@��u~��:a�x�g�t�Lk̸��!�`�O��D�0�,���m�Im莧����q�n/lY�嬢?b��,H����f���{#�u�-xe��=�2z��x��'��Gݓ��jaS�v������TN��{  �]�8��X�������gF�u��r�Qٛ��^��.��z�s�U2��*f	�}=�
�d*�>)tt��dlWM8��V�D�_& �XN��h��掅^9)���d�"�?]�@.���9����&gjuhﱌ�3�2׭;�L�_�� ��G�U����Q�㳶�Z5�j�
��c�6'��v��A���;`܃\_�̔�>KFs���c�`��`�?��ǐ"y�+m��h�4��3{1궦�La����w���S�������C�2:��`��3~�bڻ�����L�o��0S�@B�3`#�3Ń�Q)�#�����58Z7�6i��b�W�ٮn½b`���|���D�]Ut�X��7mA�fg��-��^[9騼aLE��`Z�Ԯa�5���� �Ŏ˘��hy4���ؽ�h�,=�j�o"�ӭlPi�ѷ��ƥ��-F�q3�K�U�>e�{��pGv��߳�$�X��-+ZF�w@�� �5�l3��*�ұz0G�_���`�6F�s���@��D�k�?'�iMܾ����0��MI�3j,[]wPSuL��<�v���:�W�}G}�Y�4c	�*���%�?G�l�h��M0)���ޘ~cǊ�.�㏔�0Tg�O���nܧ'u�p::b+�0�֗f�	{���Z5���L�9\�g����2�5�H{P�~�H�G����iF�y�\x�6��d�bL��5��Z������ϓm���PG[����⚓v��0㨞�����~��P�+�^k;}�	l~��a� J<��/���w��O��9�� ��>	L��k,`�?��2���tol6�8�4+;�~tO`Jr�-P��Tݧ�Ɲ2T� T3o�jN�yu�������	�� ���%`��NI�R�=�� ��U{����##@nԖ=���tOڭ�Z�Yc�^�����&��J�m��pd�9X߷~϶��@���ή�6��=����e�z�I � �߷e[�_|?HX ��O�)8֕GQ�:D7[.�8'rE��ZO�V�p��/����)'��/G�S��T-zNg{h�D�f�\PA�Q$"�cC3�U*�i��*��-&�0�����ys��\=��/����%e{(�Ja�{�q�e��Dſ����5��8�)d��Z�������	�����f�Ť8oKm��3�%u�����f�c��k ��e^��P�_����hj�	�q��8�;�2%�xJ5&��$p�q�%���Ձ��  :Y�9j!���όjC�:�a8��o�R���ru@��T,�E��4��d����f�Hi�����0#��1_hq���a֙Jd�K,b���=)�iJCzKZU�1�'6E9����6�>��(6�e����d:%f�� �5�R69�.y��O�!"?t*@�L�Z��� �����]��7����H;�� c�:�p8�F�Xѥ��Qo��i�6TMCU}0�jW��6�].�^����<̬��/@Fx�% Xf(x��b|��r�,q9�Ϋ�,Vk^8g��U�v9�.3����k7�K����9o:�O�y�f2�
��չVx��N  ��IDAT�2V4K� ּ�`|k�LhK�Xd5T_�-*@sc�{̷�&��!�G�k�z��Ƿ��Z�u�� ̆)Yy���x	�.������Ϋ�`�/����7߶Z��\���wMk �]�Tj���y�7#Q����K�.גM�抝:��j���Q��v����&<�A��Pc�tI'��=��Ep6*p�ar����Tk $rNU@�^�P�;�bw!��y�}�Sd��W�;����;�P��RY��9��.�z��*e�Y�}�^8?fǿA�)h�5�U ��,��| ��y�+�ރ�V	��R4��O:��=v���Yp�Mo�r��+V�1p����Jn�8:PF��y�y���(���T%X0�{���N�ۮt �7�!jC���}�.Ù�)�TU*\߰�%0ӱ{Uq�ɳEαG�%Ϫ�D�j�����b�X�M�%��T& ìPkYu�Tr������ʥ�]�X�;��<#Aݗ�!eaɫ�=�y����V�Y@jP?>��!sR�o�Q�K��!$ឍ�~����?M����XZV�ߒ5�?����Y)L������u�*��w�ܬt���@�<�c6�e;��痩,��i�@[V��-2�f���(�29��^w}H�u>H ����]�r���]��r[��Ku۪��=j��ڋ\��<�>���Q��7�>V�s$o%=;!-v:>�Y}.[��>���(����^b��U�x�R�*X��]�����a@�f���ʜs�)@u&��RG�u6.��n*V�å����&`��s��qyK�-��ψg��Kշ���\��.�gJ\��,7`Y��V�c��Bo��d�WnZ�u ϶�.�����	�m�)+�����p<��S���bm)S�qTM�	��
�����R�?O�F�i����X
 [�S�SY���$K�%7�J��<�,��K�?9Tj
��y�z1ub�9��<<��l��5Z�l� /�>�VfǪ�-�w#�e���kE�u�fW_�PK����99��h)�������N0g]��ʶrź��W�g8�yNہS����K�J����p�s�6�����+�{՛�0���]٭h�h\����Kn�t�u�����8�@�n��+l2�J=�kڙvɱ�r���l�A̏����2�w��I�չ��)��A��j:�oa��-��*F�W�R��/�I*1�g���R�>9���
*�S���yb��x����E��lц�٧�t�o�a�W�>��N��tA�X��O�m��&��4Ŝ;/ʶ��ԡ��eV�0{qΕ�=�`ۇ���/{Ƃ�j?M�m	�Y,A$?�G,a��3�_)\�~ ��$WK0mcS�_�㛎EV:�)��2�G�UI5��Tqm)D0� �15v$�������0v�\w�y��Pen;I�ۺ��!oSČ�Dӈ����Ԗ�Nl�u#�v�*�2�s�*;Wʂfp�H��㢰�q[��b�5IAhW��U�rS����n�J��+ ������<C�:7��b�G��=p׫����7�K��0'��8��Թ+�J�q����O{Hk�� �=
��}6�g�1ܧԷ=i����*'��/�8돨'���˛�|]P,��X�L+e���$N�[.� �~��t~ܔ�K��z$�9E^���n�1�n�k��L 8�&�`�	�������nԤ(���̗h����Ps�����`�2�v�UG����p��p�,3-����h�hí���|�ra�_�ܭ�w��|��K����{��x�c.�hK��&���,Lf�M<��-���K�u,�?�%�i�����N&�z�c���G3��7�c9�M��sD�F����k�k�y�C�@�(�1��-��V��r����<�!���P�<�J� �+�&���D���� ��ht�C�ϖ�~�<��!y��P�<�J� �+ȶM�~t`�C�[�P�<�J� ԇ<�!��� P�%i!�	VC #w���,��X�k!$�G�u�����[�I����W�q_����}���N{�{�������%�?��#��e��ҾVL�yO�݀jK����q�mX�ss]�.���K�<W	&���Y��{�S�|�+6?��x�y"��"Lw�Q�*n��{��P��5�w�O.��eк '��=d�k��(����0��*]�&��{�H�Kl�~�m��=�g�;�3�C�ƽ{�@yȝ�P�(K���|�CN�Py���e���h�X=�Z� ԇ����z�C~y �C�\I�z���O�5e<c�_Qݿ4ֵ<�sY��޹�'�$���Ӕ���\U���7�d�y����	1��>�!��5�����1-��L�T�\Ͼ&��� c�s�i]�C�K�6��E���Yڣ������s�}
���s���r5�
<�Y�jVc:���� �Xs����?b�yA��8�x2���,e�3~zKۺ+�{��Aq��d�3r��J��o5�8n$4�����x����x^:��wKeؘ�e�>klt�U��cy~J#�$>[���(������8贿uUΎr�qw�\_�`�Ӑg6�%�i�Wf���g���� �Ҟ߮*y�#�P_H�p�ڡ;�|�3������lM�}�2�7�/���ϸH;�xM�%KIl�������&����"��~��Y���=�� j9��9r
���5�=~�=0��~����_y�e��vƋGr����2��ru�����C���*��1ը���6n�	x�V��Mt�������Y�Te
fUϋ�t�|	4��ʧ��H����2��Z��۾-W��ǌ��oޝu��m��)r3����0s�T~@`���"�V��)�����)�3ݣ��#�G��R���=_���c�������6�$�m[�w�����G���ܞ��l�0���g���o�!w$��^�6�����bq���w=�!���aS偕y�C��re��Q])�x�㥜�(ݖ�bAr���_m��-�*����k�o�Kk�˝���cO�ܮ]}���K֒nw��ع_9���̀XF������{����U���w�,�<����8ӏ;�t5o��P���U��<���D'�1���f'��s;y|��k"��#�� ��aN�5��A���б5&�2����a�g;���h�Y��"̲K]7�T����>���w��Y��+*[f�_hD\�������x�k�����Z��;ƊG��<�!��ٽ�P�_E����H�}�v� ԇ<��G��+@}�ER�C��7y�㏗�>�!yȕ��y�Cr%y �C.�������� ԇ<�!��< �!y�C�$7 �K�����w�D��4�r��S�������s ���?��h����oGN�Q�ں6wLè�8II�F��R�n)��q��X�ۅ
ekZߺ ͪ��oE�?WEH�vh}߭�ڼ�O�Sk�+$�e�m2��I���,_�w&��$�������^�&(/��xj���ۿG��ߌ�LrӞv�ɂ!�TƑ���#GH�e[�p/S��jAV�N�;���5{�9K���\,�Nք	� %�}�(a�t"�=�4(�S}>�S��Mj;���9}�������8�b��k,ݿ�.{��O�M�W���˶�R�I/Ny�[��h��7jy\"���+�{����V��������ϝ�>�$��%��|7yHz8�n#�P���L���� �K�d�#e@���<䗓_Pgj���5V=��[ mX)�m?�!�5�T�[[��s�nlA�]A���C����{
�r�T5���mm
�ǿ{�y��C�(�.�fQ���1ru��_J�B�J��p(��EY����<�*��*�e�כ�&l�W��?�!�����w����
���>�!����W�����04>�!�4�>���;ö�xFJ���4s�ĕTe���/N�,�}��v"Iy�|=t0��צ����>���l�]����E�j��`7>k��8�,�s�=�B~�����j:Uh�5��-�dv
r�f����~&^ru@Żc�mj~��(+��tM?p*���{����w-f��~�:���x�k��jD��Yp���L̼����d (���d`�u<�4�ŒI�����D%mlp3��"o7���۽}M�w 7��|~����r�b˾�OT�/$�)!�E�0��&�A�����4�kݘi1?_�1��K�s��~�j��V�Wz:������?��/�{�Q�M��Zi[l���rZ��X��h �Hs�w	7���W;�.]�o;'ދ̆�Z�ĮQ]�HQk��U����rf�� ?��vL�W}�z�?C$[��k��%R �5��5�~������x�4��m9���(w%?��`�,���S���i�E/�mL��P˶>��r�7/��{���ٲ��3=���ju�2�D�ܻ��S~@Šf)�c��=���`*����q�Ƃⳟ1��r����5����A+;�gۭ�傦�ކ�ikN��y��ֽa�,!t��f�\
w�*�4��4�z�jW��샊����ܛ/���d誜���w]},�Ԏ�w,��K�]5g_o�Ս�T�|o}%L��:��K~7�2��O(?�.���SN���-�pwXP�f�n闯����J��޵L3��#{P�}���� U��b�������N�J���<[��E�J�V�����w(�m�2���`z�m�1�����J׎�_����pSIX���PL�pJ�UM���k���g�I�(z�٭T�{�Q�U?�f!jg�w� W4�7���c�i�F�?廫+L��	�䀪c>��A5��r�`J�j5u���8�pz}�7�J ��ٚ��n�֙8hb!6T�y��rY��@�~�hY钪�^6���zΖ�Pը^���y
~5�~��J��O5O}��PM��,��?� KN��?�\�å��IO�y �
.O�傭Hcl���/�9���N�7����v��y����/�^cqU[{� �w�<��`Yxhۅn�^-o���:������j���}+X��Q���}��ٞ�K	;*5�T6��)�x��mM׉�x�<��r�������T�����;�E�t�ö=�l�~d�95�W���X�=t92H���Sw3W��{�z�{�>�	8�8��������1ʺ~{N�N%��=��jSuȹ3FWOE���)Y��r�3�L=�6������r���n�T�5��h�ű��業�gK~�W�_�N�i���퇌��ߴ�ٿoo��w#����9���Z �a�`6-��%�I��OɆ+����*�m�=���S�^�@�R�L�Wm�ڵ*Y�{�Lr%�l���~�{�~������k��݌�V��%/�EPM5�"�]egs�Ƈl,ϥ�}eR8��Й��*מ2�_n�� �<��J���Z5�^�W���WC�U������&��4�KO�0e������ʄ����K(�..�Se_+���mnӠܫ9p������}��s;ǝՂJw�������=r�J�)7{NT��v_r��7:�����+S�!E�bu,��P�ZyT���Sh�T���x��kl�J4���O�ۜN{��S�
�惂�����２61�پ~q�;��/��n��ފ�T��<ԧ
�Lw9���=@��7�P7/cZ�<g�����o���9ЙyS�塤�Đx��?��Ë/���_O���%F�|s3�1Ը��|| ��{�s�~��x���:�t�sm-ljƀE&�r��Ln��HL*�;��V���g�3	j�rm��L}�
^�rA-�o�Y���܇�7ӹ�V�Tc�.5Խ��g������	o��L�����?�*�,)�A�n3)mg���7��.�C�A�\y�ʪ���#s�i�E�Y��~���ʿ�����0F]U�u���{k�bN�sg��N���\�{c���;�*�I~Ǌ� ��K���ݵ�mw�W�`�������5
����c��c6m�&�|����� ���v]���O�s-��~~���?s���J����X�Ȗ��s[�n��ݺ��+��D�-�K]�*����ru@5[M���s���6]2����5�4�4�o�q�3�/xӖT�sO�i��'�T��k޸G���{��|���7h������eH���k%m��U8n�E�uY��^��;ɠĘ�!3�[Q
1��V��)�9��#�b��p�
��A�͟�t�T�'�+�Z����t,#9T��l��;�U�ڛfq~�~�/|����O��7'�y�_���u]�]�Als��]�U��^�V���qB��w���ƥz�����7g#+��.[�MH�rtyZ���m3��A�Yy��f{^����`�����y�k5s�J��o��]��
�)�1"��_'�y%�z*C�$)�a`��s/�#C�A��
�� �b�̒�h�-��oe3R\�׀L��6�� ѻ/?��0�is��������� �~�z̨��z���+��-�Jkg�$����7Q!uA���	_;Hm����&���� ���V2�Sq�\M��-]1oŊ|�J)�%�0N�{J��:iuK�n��{ x�(�8����;��VY�nbC�3/ %�����N��=��6hf�T7؊�`i�0e��81@Fi�
���ܭ�bg��_b��uY�Oˆ�垅�o�9�i�X�7.����*�B����(a�6���0TE��~J20�l j����^�°����-N��="6DU?N$ݤ��Aj���������%W�%�)%Tf2�J�,W*T��6Nflt�b���K�$�^���E�^G,o�NP҄��cT�=� 3[g��nen���k1�L�@DY��U�ΗZ�y癉 '�M�3��lỶ�VE*.��
��؞�}��rm{��c{�	���v5��^��j_k����)����O�걵��__n��/�L,Յ*��f�ʪvX�k�ca��Wys�^�����V�Y�hQY�=�C|6ǹj��{��^�iqd��:&�0����ڽ�r�H�I6�3��^v�*g��n�%E�.!֔���)N��*���5�h[�������iE�~Z����3��h4*S�+��|	�s�}�ِ����&���bZ�5���F{�h��L�4��.1@����u�Ճ%��U���{�d�*�vkW��V��0��pk�yejm���1P|�[y��-iv%���s����$>f]φ�2�z�fbZ ��%ҫTc�rj;z�]ƾ><st��L����p�X�l��$F�&���>���$�U�@6�
NmJ0-�U�qC��C�zU�]N��JPn%?lO)�Ե��>#��rj�^��ޙS�j[ j1>�cX�sg��Ċ�V&��f��7��|mӛ_u�w1Z��j
_�7 x���Vj���{+��1�/S����x�����p򲭮~���"��d�'���ˢ�r�*�EB�4\:�YT����j?�ڟK�Jhu?�����u����62J,��,��N�U��`���=�(+ξ��i�1���Y)��BS�p�2G#�X!�Y1����e�聵�ߜ���B�����#���g�Y�5H_�C_��±��Kb�S�'��ݓS��Zcv�L��?j�QJ:1e{�ʦ����ab��p��ޥ�l�E�)��{W�M3�c	���8���f �90�h"�SN�������P 68R�Ylp�%�J#����y,�VY���XI.�鉧6f[rj��Ti?,�J����-Q�#��rQ^;z�Mp�n���[��vM$���o_S�{ͣ/`��M���]���/���g{W=��Q��x�	d���w��nEċ��p0�v
�儺��.k����)�� ��_"&�`��Μ��E)9�l�Rņw���G�ٙ���g�yߵx���x����uK�mb�=lr�_�x^�TZ;�-��:&��S��[��'��P;�������S1x�z^�@�u�H���i�ur�>�Mq�6&���Ѣ"��E[���nǓ3Q�����?�<�����9����K�k����U� 6���:O�d��-$��8T���X��f����"�:�"�bEFw���R��u���6A�k뛭��D���.Y�3��� h�k�s�k
��;ܥ�ί�1��;=��ťo�wu�,	H��F��mQ�K�N�%����Z(���Ѷ��������m��{��s���1j�����_6�o�/�8�����Yè*-�:N�O7��]|D�ޑ�^5�Y:zR@��~f�8)Y��ɒ���:�����}��i��P1��[��K�\�Nۋ6杣�a"�B�9g��Ǥ��C�������TZ38��Z��jn��>�t�Lא�kT�m�l��-����gX��N>�%�?W2X��W+��v�y�n��j�HbYY��;6U.�$�#��1T��(/�XR�XL�����̀]}�6�{^�ާ~�O����'���L��d�����zw"h|a��/��R�x�=s����ԝ^x7U�@@9�ӉڤWv��1��������V'@mXf��B���|�e7��Ap��"�S;#3����`��`1Cu���n���P;�(sRc}j�gi��"����Ń��M�>i��;Q���n϶�.7��`�!c���q��*�����͹��IT�K���Pն��#B�SP���tZ����S����LM�����mS��q=~h9|;�KI[t�2Ɍ`�2��T���K����1i�d�|������;)|i�]��"��1m�Xa���<��X����'Vie��i5T�I?`|�ygV��K��,=�Nޛ�7݃LG��H�u�ÿ�������{p{Ѹ"��B#!����2�A��PL�Ts�Y�+���Q��n����:�Q=��~]0M��B��D*p�Fji�l�,��K�L�6�����9�S����� �ǯp���E����2j����_�<t�;k鳙.�A�!'Vf�=���6C/��3Ry@M���Ax,���pH����<���?M*և�~��k-�:��՛����|��gf#2���t�U�N��E@�\��(b@�op�&� !4���N�B;I�If�dv��A;+�ȀO
�]W-��9Z?��T�שnILt"����8��͌1=��]b��I�=�x8�o�]�zu �VS[�v����L��0��e�l��	y�M���m}m��J�:N����G��S9���Qzn'�<�c?����^�uT.[�uR�<G" G���t��:���S����'~gN�B}�j��˞x���Y)�)�� G�1�b0����+)��b`cJUV�` ��͠��uʰ@r�H��Ri���)�ԧ;�����ej*����UL�v��,�P/*{9@�ޣ��uߘA�1.f��'<�b
�=U�9+Ux/���e��S��G�O�I�f ����Ϊ��ۉ<%c:�����>f�F��ji*K���O	<x��	{=l���KW�X_����<P��!&'3-tV��S�5�G��/��'�s��Ͽ�fh'e���S��NI_�~�"fJ��p����k�=�_�u1� �O��Dm�VHE��po��V;!s�"����Ƒ�`_H����x�U��1��J�FuL����K��:���/L$Q�����H�8��i������<�i�' e�����њ����:N)�1uff��bM�H�zrVg��'�y�,3� ����H�WE�d���-�:MFS�"�-ZJ>���t�'�1)��1�'d�,�s:�O�ϣ�˘,!ʪ� �����}�ԌтiT��A!�6T�We���Z6�Z������~N���29�<��ʷR�ɂefe�V�C��`E�l�W+�����ږ�� 2_uu�:CF7���`=BA���MM|�=]��[ީs3Cv`5���� ���jh�L ���@�nd5���4���L�Y���;��Od�e%*.ݏ@��@�ߑ��̠*�4��YY���:Qa��q)�G�{�Y�B_Y`�Ӏߏ�%�Jϳ\T�T�S=9�t�Dՙ�i7�3�ɩ�r�����Ď�IK��YU;�J�_�r@T-Ț����Tv�=��n���D@���lIr�M?�1Tv���gö�"����{�.��!m� �5��1)CS���J:���{1϶=ل;�Q]�*�ݙ�cp<{a�P��FV�T�Wd�v�>h�+q�]��*��~���h�$�D�}�
f
餍Q�Ŗ�f��1O�����\_��gQGɼ���=L,���Kzy�:ϑ���z�	+�M ��I�'@=���j����>R�m��I5��t������LD<�j�S^������kQE�%Q}RY_մBB��k�@�&-�y@���X�bb�>��ebv���'}{�����B������N>||�q�晃Nt��_4*a�)�&��?O��c� ��4Oi&_�|M���O.׷o����ʦ���}�u�O?�?p{�S��z��������v�I��ǍS���B�;5wd��H�r�7���Or��)��3�4w��l����_�Ec݅��Ħ�msb>��j�i�tl�Y՗��S��&�Fx��t��F�_���� >jP`K��QmP,P����V�Z������hvP��g옹�`Š��Zj$���e��zF���#��U�Q���:*�G��C���<=?M�{XT�d{a`�ze�%�Fd��%'���~�2Ӭ�@������۽h�����g�������N@��:u����q�?�s��gg8��8�8�������ӧOʢv��V�u�6���|�NNj�V~}R36���2�:V��f�O?�u����`O�����"�3Y�e�w�Ug�B�Ea���LJ|�h\p�����
���]����4A�
�����}��y�ݙ�Wڷ$����	��yO��J���4�rL*� h�N�Q� �Q3Nň�-�:6�P�E�v�����������1�:��0�����g�I��Κd���6GU�z���%yMpF��Ҁ�Y�U�]=$����Hਃ#�MU�eeO>(O�;L�Qfΐ� ��1.ϩ��C^�S�XToA!�qfk�NK8z�p����qޫ��P �X�_�-vou����;�8¶:�T�^@�8�>�
b䤙�)�;�}w�^�?h�Щi�h�X�T�Ԩ���I
�x�S�$}�[�:��cG�ij?b��v�z�`a��q��#���%}��=awO��5�oFSOe�oB�|�TqbudW5�e/m���$u��{�eA��j�0�؏�l�����R�%Em	�WR��i�=O�[8Tx�5��P�$���4���y0rz��Nl�$=Ox��������noe����x}�����_�k�M�Kjw��`T����L���s�r�2�i�P�ډ���<u��(`��FG�z���胛%�����*�&�kϝ򩲋yG�ꜚS��<�<`z3�[8�(�@�~؆��B��B�"ḻxN��0!���+����PE�g�~J�@5|	6e��̩}'�aI*�� �46�^�1o��D�w�"�n|����7V/���������f90�]B6�����R��zB�A�T��Q���=��v�Ws�*���b(�l|j]!�S�% ���.WOѯ�7��p��`�D.\�?���(�P6��w�Ol���6ޤ�(i_�-�Ɲ{c��7܆\��ã��hl�ɖKQ?�L@0_�3��Ii�:��?�d@�?;zu�a3Mӽ�S�Q�xK���Nm4|U#�Z7���5(��C藩2���5}�T�#��ԉP�]P4(F`���
I<�I]�?O��3ٓ�RJ9d�C���P9;���es����y�f��.�Q8�0��2�3��tQ�^r���GMn���F�]�	/X�@� �j�Ҹ�81�f�KB� �:�~-u��Hz]C���X71e3TfR�	��}.�O*1]���A��5���6&;���߮s�;�y|�������۱�!]p�I;~8#��,��(8�]�Y�HT�[����4�G�w%i�[�r�����o
;���R��������I���B+tv*�כ�A�<Yy�nEՂ�'=��\�کN��ݑME9'�b�~�	��&9����B �g���A��F��ҏ�⓲*�!ZHW�+��ڱ���J�N��_S�~�@��ǺIE@-���D�	T����C�܈�'	����
�}p�� �8K��]�E����F��+�s�pF��L-@¦Fc3�>�D�a����!�8ry;�n'e	��4g{���Z`]8^�
&�$��f����NT&V��"K� =��?��ZtrBQ`?n�����v�Ѽ���d�����$�LU�md> '��K�~����y��o� NF8���q,>�4���Nb��\WM��K8�2t���N ���*&(�'" ���;�U���^dBRG�j�`�R��ۙ�	��ݢl��Z�o��x�a��#$��cRME�����>z����n԰K�9�ǍE@<B�x���m}�Rؔ�J��ԡ� Mqe_H5���T��沍Lla�����$e��$��p�����U�;zJ��d�NW�P��h,�'��Bm&�A�ଢ଼w�ٳz���Ǔ�z>1�$1�B�S�1�'g�)���_��Y�������r����}�Z'�N2�9$L�xՊօ��Q�B�+qr-�āU�F�k߄w+�k�������1����T`��~bL9�}����~(;�Y��J-:�Ϋ�X\������������D�������LB�ѵG5x�)Έ���D1ƨ,W�≏�▟�����+#"�)=��P��|���Sb�-�N��L�d������C����u��ȶ��//LȄX��C`J[�&���XB�LJ;�s>�_C���?��"�� �5�K�#�59�eJg5lT1�\�~�X>]����1}4�I-eUK-{v���A��=5��WЈ��;�46���y�zBh>#x��Q�a�b��̋����S�/G,~]��Le�I�z0�� L`��=d8L��0�0p#�r[�"b���Q�'?�ϻ#F��=�J,�ep���Ӱ�4�M !���������r=����D�Ղ�|�@��W'�5p�Af�X��t��m<���<q�P��e� ���1���LE�<�qx��{��a!z���]�]�y�V��~�@�� +CF����A��L><�4(Y-F�&i��M ͓ �hv����X�c{{a�x����{�m�r��RhD|�ٷd��X8:�u�Yl���t��$od���|�x��	\�b��Y��*5ƿ�5���\�"�_fG�֎Wݨ��\_�.k�����vi����RI������BdERg*?�(L	c*!�y��z�S���:f������ ������ޖ\���&L�m���c,�Dk4xr�<Tj*Xu�:7��x��۱y��18sR��T�g��6�~�N�D[;�g�\���u37���E�V׫��Y
�[���u�.��f7�����󈉲x��1E��;�������������lYl�c�T����9����������[���JH�=��2�~}c����;!i�8�h�}��,A�s.M㒢?^_���`�QS�z�az#P����7�@NC!9C�0�Q�����חW��']VO�th^�1�����q,�+{�ɾ��l��-jtz(��;���*+�tR��S�O��������ET�v:��' zzڥ��ӧ�n)�頁�$��Bx^���M+gN��ꎲ�آYمih%����f���<�����V]#����<u�8���-��� aG�L8^���݃�I�H�|�_)��Յ�U����&��uv�FeF`�sZ����F`�wV�L�,;gaﯔ��K+����V^Z��U��9���/�6��&u���;%VH�[J�8aρ���	y(T�?������E������~�������P�ΰQ�tq�����ǀà�|�c��s�ؠ��s��I��v/BZ�����������6)�t?
��������ҤD�A��HW��%�C���F��>���9mac3{�Q�Ti��C+b���*���7aIA��:�o/~���$�Y��q�'P�z����K� *�E;]~8L�D+Lv�=>���Uc4��9�|'K��C�4��̣jS~�T6@��e`�qq���dC�KZh������1i����f��lp7l�7�� ;vf� a��ⵍ�ƛՀ@�e���:��r}�w�L�񹣩4L}	ͺ�Ԟ�:�����f��ó-����c����%5����?�$}�򒎼
p�+�TC�'���k�l���<ǔRj��ɲ�5Z'N<1%��K1�P� "(+!�2���f#��bap2��-���6�*WM��3T�0C�Xh�����HHu'`$O�d�dE�(��3/)���F)��=�K���yH&���;��n)��auU�Ӭ��+���J���1;�(,ZL�a�L�L��Yųc�� �dUX���u����j�)I��J�]��2:��f�UX�g��N�i;������i��iq�����+:ۙy$禓C��4���@k�US��W��f�:AT�6f��ZXC��"� �rEY�f��,��33/�ռ61�2~e0# ��>=}H�U�{�S��qJ��ŋU�$��b1��Tl�b��i?�Z%9�"�]2��$Y�^���%e;/�����%���ԧ[�U�@�����и���ҥ��-b�]�f�2��I���.Y�����M������E��(��l����A��hI*����	�MlH����=�j,�d�#;��ç�y�,��}�'�����N�]�<ˉQf��`���
h¹歯e[:�=t�O[n@�A �8XF�� �O�y�,'|�&�e�\aW�S(o��L�DĲvh����Ѱ~��xU`'v�As���BTlR��<�����?�O�P���d�c׽��X쒎Y�?}d߃���;O�(��0�{��l�D���zه�Ê/�e�H�Lk��o�
t]�.CM�� �/f�!�Xz�ه�	��N��_!;LR��g���"�=edE�4��̈yſ�=i�y-nOgHT$���{QN�����Q�>J��ab�̲�Z� TJ�֌���?Jy*v���nBY8��Ճ?�@� ��3�ce�u�c|�+��m�P�U٢-1���m��8�Xj��J�ID@u�c�}_��R����X�� �c޾+�Wz�kH�Z������U�y�~ر�]��k�Umh���sJ�+�
��K�-�Ė��r�� Zp�?娙��M��_����n'�*�^�+�2]�#K#B�˘�6�\�o�U�@���=|���h'�D%��B9Α���2�Ny8N�fT�Ȝ�������f�AV�dK7��9Vn�	�������C�d�;&d�P��cO�x�%��G�3�*�uV/�8���L�+�-��jZB�\/�=�����: W�h*Ŗ��|���s�ņ��i��*�/QM��(C-�K�h�Y/��'LT������5�deͤ�چK�[3�l�� �����V���?�W�C��!¦d�� �Iw��QrHR9���rHKH*:�Q1.����1S$��n��,	̞�����?d�kZI*]������{"G�d������"-rߋI�������Hn�x]�
��?�:H6�2J��0�,�վBd���W	u�@d
@g;�4�d�Jd/�hd >~��wz)�
3(��=!Ϣ��W��z��1/����oNt�{��l�%�2���CY��f���~T�MNr-³��zk������ߕ���}*Y]J��F;ހȀV=n���<�4�}*��GV��RW̜�ڡ�Q�9:�͙�	Ydƭ4�ZT=yv�l�s�'�쑗��E���^L�Qw����] L#QF���?��o�E�J��Z��3PG���||�\��~�𤌷�c����������ͱ 1˄#O�<1�>,mpBʶ���r@�ؿ�[EԌn��N�jlʑ��_�R��Ybx5ϑ��R��xm򷗯��GYCNy���L6��PC̙�������� ���*	���i��r�^��eJ�3�c�r���<��`��1+-���'����ȹbSs��njNX]ֿo��n�kN j�ٽ4���j��-�����>1E�����<{]{�X���3��)���\��m����-�ޚy'] �Ʀ8���>��{\�AU�#���S1ڸ�R|�#vi2��tO��ƚ`�����c�9�u
s����C<ÁA5w�C.�`K�D��������0g��^�����e�53	k���ƑArL/���?�Ⱙ���^�D�|�SE�9���?=�/_'�:(y��A�s���b5el�������t�US�qPzv�y�-�3 Ld� �Q�dE�LĞiq �R�N�Z ����Ύ9,��y�Z<>W�k��[�jO��Ug�$�޵3�s�"��}/)��ݒ=�=�-P���T楺��+�B�W&�Ef�P�ZV��.	�w5an��P&7�{��L�� �=�"�H��~�ʌ��D_��L ����C���z0�j;�"'cb8����O���%$G`;]L��9CG�3̑�+&�����0Fc����u 5g�}	�U{���Nͳ�Af+�A���h�%NP9G�X���ub�d�κ�VNH�BL�bP�؍,�j
�EXY��Z�ʺvJ���=�)︣,�����ꨡ�d��dEPQ5�%�y!��b�CF����amB�Ll<�-s)k ����f���|����P`�h�Ԃ�'a��|*we[��}�Gv� ��4���s��b�Q�+��^���k��~�,��%@p��2n&Nh����7�W�܏����r0&J ��$��$�~���=�a+��Ϣ6�$�U�Q�&��-m�:t/��v)�&[t2�iOU���L�S~��t�Y=.�����z�m�IP6��T����>/���{��Q���0Ԣj�4�M
�Z^��1�m5��U��$"��yV�Fq�X@�+V|Q-F%��:����-܎g�QRڨ���e�ɂ�1��d��d(ҐO���2�{����k�:k�PK)��%�o�ɏ���A�©Jd��	�Cd$�-8.���5\fn�I���l�i��&	 X�����ʯ�h��u�6x���L�J�׾���cx�ɫOI��4���J���D'Yl���*f8�I�X�)9�R[���5�f��H�-	��d�G��������������q��)�v���0��`Wc�8�M�1�H�t<D��G���:��/E5"�]�%c?�%4jH�����S~����0m��1l�F�2�Bɣ�`|?�v!�ؙ���=za�e\T�|js}���(���
LW�+0m���P��G��:Q��*�7ٷ�O��B�3��f�R�AN�
�f�3�
]�p~}���*����c~�ۄ�k�JyG��Jc�������_�E�mDZ���:dl�-�u%;���yl� G_�&y�1���+eՏ"99twhpIQv���?��H�M" N�RƴOHш|��L��u-R�:��K�rо�^iO)���v�ݎ+�¤${=E�8��|�3Z%w��WU#�!:^�tx-�Uf��h6��A>�Ƽ�t�e��FX�G9�*�|���3����#�2`�����>C�~ݥ#X�fґ���L39eБ-M�4Ц0���ٌ=��go������f��{T��%�v��V'宿�91؟3oU(���y/,i�����"�E�{�ؿP>gD5.���@O9� Dx��)��	j���՟���Ǚ%"-��;"Q����{�]��=gc#����Q����0&�k�I"^F�L�m� �F�ħ�T�����xԭҳ%��q��'��V?������y����W
�z���5�����(U2�Z1�X��Q�+r���q��S�#R1�!���z%/?�������a�9NQ����{��}���]l���Ӑ�����G�v�K<Ӟm:� E��Q{I8D�{>|Jm7J�5(5�]��D⅗����NA��AT��gSw�~�����_�}Sv�M��W��u�<�}��YL���ߧ�*G1��Tt�R<�s���4z�Z���sLr��XT%�������KO��~~�Ry���
o��x�)!�Ų"�6���q�kS���jտ�4��mGJ!R?"������6����Ӿߩ�*r7���l�:!�5{�b۸	�	�kHN�2&X�2��o?����ǟ�bO�[��!l ;p�M�4%8_�#�Tt��t�2v�0��]�aR��������b��h?���i��ˁ�9�4�@v� ���(eӐG�A�S�o�GX���2x��j���>��\I�^�l1O���T���Hѽcl��!M���WD��=��;�����ʤ���$l�#cy�К��X�T��jw��R� ������vL-76��� Y�'eC�d7��Ē1�9u|�M��׿����)�U%������#wB�Aܶ�)0���s�u������fV�'׸��^�g���U��,)��A���d��\=�)�����]"�9���`dLpi=�Rd�:Ɠ�KdB �"�=*�3 䜁9 �����$5Ř�qAGv��be�F�.��J���ݣ���ҿ��21T��堲C1�esH�1a90���=6a���7���X��c���c��ɎH�X4�G^8n�#�Q�1���D�4������¡^�!ݵ��� {*�C.�b(�;�e�ǥ��Tr:b[^�Y�u϶Pn̲�F�uf�x9����A�f�B��}P�TU������f��*�X��[�3!ލ:mu,�� ���1zEwH=u�v�";X� |����1-2Ј�Us�t���� �WU6Y*3�=	�Y��N8.- |��Lxp*s�3X����0�'u�qv������%�"3�����.N홓�p��Ž�8���`*�D������ ����{Y=8�����M";$��my�0��9�ٷ�A��+`��6��c���cN�Q�m	��F#j�6(	Υ��@����PS5��E`�Yr������y����B�bQ��8��.1�#�s�~�َt`�t+߂�3:eGR�}ll哂�y�qy7FݤZ~eC��<0b�'P�z�:��9,[N�!^V�Px�0���Ub�<�skj��<�m_9l�K׿��D���l���:d�P��F��	{���aV�PΊ��ok�c�R�4&&/%�2O������$l����U*оʶ��v�sF$��,? J��\좴8�?�H������P��Ǐ�x�a�4�o�M�:�Ԍ	���JY��o��k)1�q��j���w`��飏O۱�F�O,}ͥk�������f�qi�-��9�So��&Yg����@��{1\K��vE4��ԳNl��d���f~d;%peU�*�z�aH�ҍ�%5�K��}�Gt�ʃw�=�G�%@�������>}���}�N����w=eu[��Z��5y�G�L2���7���� ��K�S@��b�i�}L��$
�ın|����8�V2 a[��"Ȱ��lvϢk��?�i-^�H�ubˋ{|��4��Z��9����_릕�pt�{�?�:��A�m�MKF�}���M������_��O�N�me��#�n��0d.x�I���=�V�X����TM<�����ۛ���Q+�MAEw΀]��.��_ƪ��"U\=�vh�+W
��PTW�FY�R�b�ˁ������1Ҋ������; ڣdω��� ����d�|L�@Z�V�`UsZ����8zEPyċ�M=���w������Ug뜥�y��qH����_���� fڬ�u�������2%�<� (_|B�U8a�P�*�RtɡP�	��M�O��R�Ez��2�.�$YT�=a��*���EU9.�u��Z�S��t��՟å����4�-N�+ 4A�T�Q�9�)����?m#����	�ߔE�8Ȼ
s��N�t5hQ$u%"nl+�$`�	l�7��<��D~̄���73@�����l�U�'GW�\G�DŦ�cY����\5*: ���,5&��E��.*� w��W��j<^:ZTm�?����P��P�0M(v~l��v�l��S{݁����c��o��9[��>�K�/�E��R,��o���e����lqvl���1��
%�@����vn3�q����M�s���FP�R�_�}s`��AcO&78��jf,3gۿ�z�]�$��=��	��e\dt<�qOo)�����I'W:�����,��z���X]$Ri#&�"��k����/ {9L�����*�����:iy-Jr��H�"%7G,�Ge��<T�������ڒ�)!g�_�6Uy����������P�[��	c�� �*���I�\�j`Q�}T�ql����QJ���u��K�c�]�N9�󇷴/{ߑ�x�$�������li�(�����Y�!g��J��(���c�v�%�	n#���]H؆Γn˒4	���P��=x$�`g�.4|�	a)α�U�<����Y�4��;�Z������L�l��~���P�1UfsF5abՀп;���m@$s`�	�j_=�J����,����̡�|5O��˸0�hQݟ�ڒ٦T�'?���I��N ��,=��z]�P�����_e3L�,����y���M����y�xl�L�&:6s�=ۨ釖i3c����j1DRm�v�P/�_��e�d7oDR��*�߂�lP��t�|��$ 0+���1���{�&R� �S��>:�S�VR��j.[B���$�����i�b�G������f,5��LptE$<�̜G1�8�d�!�e����?���v4�ȋ:'F[�Uǝj�ڠ�Э���B��q�50�fe���Z}�qo ��R�,�(;��qc�nF��0��{v�ו5T��&�F�#�b��QRF/������9�!C���R����*޴��"P�iU;ٍ�h)4%	��N<�K�-���
p{��&�8/F��x=�"��
S-ԓ�y�ԯ�U�Ϛ{�ۗ���y�>N���[,��b�n�yE�t�	��8��gב,�j�����q�R>T,+��S�T@�>}|N�������((��������%�$����7ǘ�E�L��2�^�.��}�����s,vpT�Em`I�Bglɖ%��4�C��2y�&�컇Fo&¥^yC�Qٮ0�A���3�)ոU�f�+c[#��;�;�j�\4}���,���ֹ�ktC�<��H`<:SA��Rd ��T㱣��=�rr6#'��呂�RN��J��oU�B 	�;lT�/��lҲ�[��7h�O�jB���/)�ʩ�~ߛ66z���?c��!�4��bs���L!)U��8�(%ff��+WҸ���)�NX���[s�a����{��T�����1%���=n���Z�u�1� |Щu�#&ApN(�,^�c�t[�N~���'�?�`��;� �a�W�`�࠲�N���R���`�Ps	�$���( �@Y!�j�@��8�8CV2�uE}��]k��w�z�ꍗ��s��E���I�g;����k�x@�N20I�Х��F� ����j�]3�ǔ�u�2N�-�*%c�E�(��N0������K��Ǥ��\}7���똳~�E3j����VS�DE@�͡_Y�A�����%�hҝA�3����ޝ��u
pq�A&u7�ѳ��Z�5���f�� ��,��64��1G�CA�EYZ?y�f�2.6�<�!�R�W 5��mt;�\��y�I81^�;
���d�������������o/_$�>'ya�AR��X���3�0���_���!�zZ��6{
T�$��q��sA������s������9SU�ζ�.�0l�v��QY ��R���)	��|���f�ޛ�=�qR�2��2d�D*��9IW>�_e a`��b�8%��0U���j�27u$B�N:@��KamA�8��� t����ΣI��Q�33m��q����Ef�&�,�n71Tsfg�ΐ�TS�� 3���}�WLJ�2��ƚT;8j⑤m�K��z?Y6ʝ��&0T��q_�[+�ـW�]���I��8Σ&_э�ƜC;��l�)��Nѣ�s���՜RF
���C�(�� /_�������~�"u����矶�N���=H���t?b������f��=f�����#y'[���x#UB@>���:�}`j)��z��+,ԅ�}g��A3p!*w��;Z|���'�Q�R���b��� 9[�,d,o5���d�0#UK��{#|�w%M�� ����w��A`�Ksp`rR����ź�&� V�	qF8>d�c~r��Y�����)ۤh F�[B�z�4	s�H�����|�&i#�g��5�.b=����a��+�T;+�~g
}���*�,�V�t��rOp{�w	ˣ=
������Wh-2�Kj���/ʀV�y�;ԏ�^ڝsb(��f�Pb�2¯$�`4�����k7ה�{�ͳ������AC7(	m1+k���KJ�N,�ö϶v���d
�͂�}�/T�&�B<�/��Q}P�1�����)���4�ai�S�p��Y�6�B����NR r��,f��A�7VU�V�%�X�.xyXǦ+G���b�z� �;{v��y�yx�Zʉct{��d3�/'��&F�YV8JF�:��j�33Q��<I�mu;�nj�w��5�8`�hQr(�A��=]o1��4]V[�r�ɻX�M&����7���.���m�x'������P6;j+Ʀ����A��J)Y��k�h�!y^o���H���Q��0'ڗh���!ܯ��f?��,��$ ~�����k�����1T��vu�*��U�-���,�-��
��\Z��J�s���j���F����N���t�\�|��l[՜�#�&[dB�K&��t�ۅ�~�% �A6�T���	�k�w�B�l�NV�F � }��z[�"���V*9u�^ى66kK<��vz�2�֑m�;�n����W��1!@��N��h��1GD�h��H���ʾ4���Xof�\�M<
!hsxxȘ0��)�F�/b�|��xZ��i�i��q0�ds:*Sۅ�d�4A{6��y�d`@�]Vf&$d&�&���S*�bdA��ٽ�E�1�H9���x0ٱiL��\��W�)0=`,�*���e˦���&��J㤭L4)%�ޮLEs��L����CM)����N���~$�yg�Z������"k���B���U�QUS�R����N���Y���^�`e��\�]ڕ����7���Ւ:�����bL&t�R�d�xL�(��9��M�������ó՛�<����҄��r��ng�s������?���Q\R�{����*��h�U�l ˙�leö��cl}�����p؛m0��\�$�݇�w�B_�@��2��_`��EPUe]{�������$�b:hRO�3Ϯ��]!���u�
N�X,�i	al��JE�w�I_�F������qp��ɪ!@�X9e5�V�_-X��~c6f��l-� �u�*yP{(���)�}�Cm�ooY�Ý������1�7��Ī%\_�y-�f��-F4TV�h��K\wb��A@��t9��z���A�u|���~�CπÁl���*����o�W������z;��$�(��&�'�� ���������:��(�`!�<��j�x�M�O|���MP�RRU���	�'�,�a�i����.:����̪ሔs��V���Ȓ��v��M��r��qe�	�~ gL�0	`���NV8�E��s����Q���R�o�����#��q����@\��*L�1������y4��h�1��ץ%����&X�6V�G��0�4�\E�6�Paf*O��`3`BJ�Q7��9{�\#*�1��:x�Cfs��B�^N���JܸL�ZJ�܏������������O�>3���tK���?뻒�8:�M����k5mڠ^tN�ۃ��w n8�}'՝��S*�>�頵�i�C5��BFNu�$ӝ�ERf2PN[�=,��L�ň� P��I�(w��*�J�#{�]�L*`�����n ��������͓�R����We����NMtoPǉy����n����+p�j?@tIo���OO��?�i�/`��C�f�xW��puZ���Rߝ�C��O�>�q��J���!��cB����>�c"����R4�u��H��dc�ը��(7�@$�e�q"�ŉ��
��^4 02�+��j ��E�]��"��WU{Դ~�(����u�.� 2cr	��^㬔�s���^VI�B*���GY��C��� `o*����ͬA� c�8U�.}����ExG�����{�,;�(��� �/1<����1�D��$�0����nW�e�w��F�3Q�;�:�d�+x!Ѩ�3*�|����JVJ�ڊx�Mu���\�Q��w�wN����[�yX���V��'c1��OV�$Tw{]���hx�/}yǎD������J╖�9��Avr`mb�z'8j+���yO�j�f�Q�.bvJ��.q����<��.h��v�m�)�=��%Y ?L�����7�6���9i<�F0T؝6x����\�����eae!���[�U������,A�R�A�����<�I�$��=옝`�)�S���!@��!{�NS�A�#֙[��9�i���Фo�X�\���&�0��<�e����SPM�:��!�%�'XL�̳X���eo�;o�B�w�4j�\!���*?�{�!h�yb�"Il���f�p�Mw����'c�X�@B��:Fٳ���b��	K�x�M�z�s�5LLm���d�c�2�@N��������Z&��Xm����4�������c&��4�A���S;ӷWJ���T'�S�~���~�>�L׉������;�.v�	x>bZ&�`z�p�^C���{4��9�3��%l��tJ>	h�G��-���P!2T�5ɋX�p,:����q�˟����ܻU��Tb&��aVʁ���-�غ��}n�܆u-�o&|N�Pe����_�:L�*
�0u5y2ah%���YR3CHꗝ�0iu��k���Z�������NUttDs\(�����Q���Gw>)��tŠ�P�ua�"7�����n<R��pLX����H���!�v{zy2���ާg���v�1/0�\��1,�����>'Th�+X}��rzi'\���%@�G���ᅳ�w�ٙ��M7Y&��F��!L*�Q���E�x��%��1sb�����o�ٳ/��+��1���w
	�2v�'�bS	�L?��_$��Q�O|{��&"[�\0�gj��mD؆6��@u[$�:��*U_��>�C0~�0+���d ��ql�c�] z��(h�[�����p��Zfz.K*ȗ�E�o)���kc�̓*`u�^TF�a=�m)(�0v{�m5�����X^�i��\r�X��Pl��5z�FR�(͚��a�e�4�D
�X�u&�*[OcQEvw���R���*�Wʫmu8*�p5Yx\ՅU4������j7E��,\f�m�����8�`we����*o��	ɇG�+S�e�ϲ�A��;[8���#�<�l��}WTYgB%���ʮ��ۇ���E��S��Xꓪ��d�$����H$.[��LrŲ�1�Cx'yg6�M��<������Eˑ�M�Ꝟsz����LuUe�K�	\��F�Kr)2�&�顗��ˋ�6T:hA��,v�i���l�W�V�!`Es��բ>�>��U��q��~x)I\~�^�����W���$���������(`�!*0��t_z�F���P��*v<ƚt���ύ�Qj�\j�U�V�E���r
&Et`��A�ׯ�w_D�� �����]���V[k&����׶S��W3�����C����b �, |���&hӻ�JE$��D�.n��á���^�Mۢ�{_}߮�,o]$>��\���XFO�$N���;��T�5P���!K%�w,�}����.E�T�Q7�-��0�	0���(�cˬ��ܫ�� �{�۽����-�Y��(ʊ[^��?��u����z[��d��o�?�����xK?
�1�f�͞���3��t��s��:Y�SË�bK�I̅�omѦ�OLC�g��@��G���*�Z��
�$��ׂ��\�ye�n���8cz]z�Q*���oZi�m��b�VX��hv�B���G!���8�*+kP�*mԊm���>�9;k�Cǘ�r<S�2Qy��Dy�����Ō�n��f���[��|���f�ySd.).� �]�Iy�n��V��:�Vs좛n�h�;�:�U��1�2� �2ෳ�4r������W��s��������_�>�/M"��F8�YQ�}��D.�A��yI.B��L�DO�����/��e�ì�
$oj�kƘ��ݷs��7 k��C�Y�5�k���������{<���}L������1���H=Η{�`����^�溄@�I�ԞS���'趿���_��}ۀ�`�Zl�Svc�"�{������'.p�N�������?{0�w�C�]0���TU�WXkD�oi)��Di������l���p ��A5\��Ď*'_�8����-l��� kd�W3_�Ѿ���]M�t/�� х@�#U����;D��-���תbaԠjE4�_-��ڤ�Z(���I��Q7κi�_s{WV�����!ت�4�ݒZMao�сB����dn_o�5�ec@G�X*���W~�!���¤�b0)�E� �c��-�E��-bBT�;�zO��ئxZ|1�I}ׁmᴅG�N}g܁�1��R#�h�֬�}=D�9ۥ�r���Ȧ3��-��r��>�>Nh�|g϶Tc���7�3=�Ǐww����곩�>m��Ǉ�Kw�i}��/��C���-X�������8��|Dt��.bg5D6��0�a������j �C�5*|�U�hư��@ǯC/?A1�NVו�l�۸��@�	��v@o�>���z�#�h؟;�X��<n�R4¦��\�4zE6�X`wONO�C-�T�.����+[Kn�葀���a. �?.+r;�£M��s�6?�7��?���2y�8�h�PN�����~��;���5��o=����$zvK]4<cV����܍	�����ݣ��7��؊?׏;�T�<�+O�H_���P�m�t�����G�4��y�O�hL'��}���ؤj�g���� �j�������o�0��K+E��()��\J�l�z'buv�&��%;9��P�|w�~�
�gX�kO9bc���&$Tؘ �3`G.��Y����{E�]�r����(�nUjA�EN�����l��xV�Ab�ڱ�؜ D�9��.���hgĩ>aq�,��n�h��"$fWU�i,��i�����v�����LSE�25I�IiP�9�Ѿ��cXy�~P�LW[�����U#��Y0�-o����I��M��9u�Rwq���Aqtz�S���^���~�t� �f�����o�âA��/A,��@ X������[�O�#ߋ^h���!JPY|�u��I�p��v��w=D�P�Sam0S��:��� tV���c�a����y*[�]�Wz�x�k7	��,bݺN{`O(��w{�8�CL�0��đ���'	���F���Ί���� f@��8���b�����E��ܙ6��(��I�;��� <�A��`#��ۍk�����E�P�׹����`/���cJ�YHe�,q��[�� �S�H�C/.�믺�y�ަ!]��'1�'���?����V=H��(@͕E������Kwo��XY���������X��PW�׮;$W��m��k�p�rk��L�<�n��V�J��%On[ӻ+
���9�U>��&�����\fڤ��?�r��co���-�����
\�U 8�;X�_Ƒ��a��x�W� �6�Mp�y=(N3}��@��7᪤ u��n����0��@�:>��g��i�����`�6Z���;U��`L>�Y���f��>���;;՘`��!���$dE\�!�F�
5��y��{{`|%�']��є {�v������~��q«�dz�3$Q#&|����h!�>�R3x9	�^��������-�EÇ�B��~��?��H���DTl��*��֏�z}�}�_��v�=`.�Tw�J�������f���TYK��b �Il�Y� ��D������"S!v�Y-qZjx��cA�������+y6	q�@���<��J���� ��L��o� 7��ǪC�E�;�}������Ǉ�?p]V�4Lr� F����>�%^oX�=�O�b.A��%�����*����	�>��>���TVK �	`H+���ߋ�ḿv�b�(���`���1"E�EcC��WI͌�`�k��>�$�%WS�U;7N��m1�n�����|i��UC�#��"�P�T���'�P!��+�}���\�P�ӛ��4B]�a�|
u/���~wG�Գt��n7vɍ��vV�}�j��9;���H���V���`��;\Õ�>k�E"fc�X����s�Pȳ0���S_xZ�ب�q/�m�I҃+Wl/.�Zݡ�'����I�l�����w���C|ףE�B��RL��[�h�X�B%��j|�u���I�Ll[L��5Q�M�a'՜s������~��AAsMU��<S�;�o'	k�TY-���8����G����`�Y���[��y��d�T�*ޞ����}�86�o
��oO�J�%��և���e��S�1�b��|���e@e�Wb��ȹ[_�p�����зF�hfb�G�]�13������Of�<�y��p������x����H����Gq�"��`����!�ɂɪ�d;� ����6��Jk��x��^�J�ar#h���ޞ����:�ሢ�5X q3�3̓V˅N/�W[���! 5T-���3�f��y�������Y?̪�P	d�K��_��C(��
�y�2F�i|��V�]�� ��Q�v���$7 ZhqO��a�G�Xz�h��VWp���U�dK�V	�����/�PID[��\-a�{�P�������ZK�1���>}/���H> ��{'l����8���齎�QE d�\ݍ
b:�;3�m�GE���lZ������!+�Ws�)�x���� ����Z=_��7)� غ>�ʈC�����>��:��ipUgdX�Eub�i� �l2$�%�?"���I��D7�����F}]��U��AG
�dwrU*/�Ok*���O��"0>;����%��C�Z��8_�;�VooR	�L����YK��e`���u�R�#\G�4�$�֧L(��V4T�����o1�r0K?��M��ڇ�����k_�j�\��j���6xK�+���Rxϓ���k�#i���zݎ��8D�/���D �㮂]�hG<#���vu �>���>km�6'n��օ`�3��.��� <���t�.���̂��ֶ(�
_t����n�Y�����G;D����+�����.R\ꓕ��!
C�Nn��X���;C���.C���J 1H�.�T�!�B�%��/D��#���S֎�!�5ư������G����6ͅ�G*�JuE����yV�3�lL���yتGP�7â2 k���p�_�.8���q�E�DMy�F���������I�hر7E��C !H���#������JFB= ���#tǙ�3) 6����)��+1Q�* ��룉���}.�������\0��3�DVWD#�("��g�@��Ǥl~�R����}�޾k����U~{�X�烖�Er�	�b̩?>����걌�ǌe.Ĩj���]�.rb ������`uCS��l����]���,Us����?Ę�
� ��p�	[�ĺ�����=^d�����H�v)�$��g,���bn8KvTgUE���B���T�%"��V��6-�����`�n4��`���������~ś"�V�B 1��ƢZ��~��լ�(��8�����u;�o�h��zt��;�a�B;��	c���^���]۽}��:�7�ɶ����b����������\|�������S�SϔB	]�h"sQ��V������)��U��af��14��V����zF�djup?��Ǎ��}�A�T��F��c�����o��8��ߏ�q�\+��c��8�Tlw�i���-
̠H���Hݒ����P[/��5��ky�y�k��`�`Ǉp.�F�f��Ik�笈�f� -?�:q�Q�4�	�z�������)� �5	�p�d>������Z
����oؘ"��.�s�['�:h�>�;�Hp�5u0�0�-(�tW�+I��k��V#���`@���%�����OR��Xq�H�y��,��k���m	�Gx�4V�����G��ߡ��|l�EW��a��X�3�l^k/4~^���Խ����}�P�j���"g��9U}��±��7�^�)�����z�v�x@]�|����&�9D7%�ے��.~�Ŋ�K".j��վq�Qe�zy�\1��$�J��QMITNP½�(��}����9Vw ������/�E23��r��}�)��' &xx����˖0O�0%�:]Pt�V�0�j��<�6��U7 �N�Y�vfr�v��=��w��/�׌m�Ϲ/{�1A*�%\W7�3�N}�������� 3�������s*{�m�=�~�M���ރ`��2�!����f���{����
6�:��W��Y�K�lE<jw�*��d�˥f��m�/:��s��`<C_��'4�x0��r=Q13b(FlNZu��l�e�G	��%�Yd|ݥ����T!��o�
� R�a�nea;�������}]�ܚqRu`���MNr�0oK
�A$�q�;���q�vҧW�	�k�o�?O��9����}�@��S��?��+�a��iy��2���mLF�h��:�l��d�̭�]�Tzn,V]�o���.&� �1N�?h�J@���R�O腗7�]����'�-���0Ԧ��mˋ3Fkao�PYT$$OH��g�u	�Q��z��t���<��=��<zp���Ax����",��V~,$1Y���䖡4�܍#8���/:�ɬPɀXÌ5�S�{g��;J�k�P~8ɻ�i�}�7���+�tk�#,�o{l������f�µPa@tW�V�=Z��������>O(ގ;nę0@b�*��J��J!0�����U_l�d�Q�ЇE���F�<.T��l�O$
�-�>�0	�,�S�: �x��|ϙ�K,�p�y⏢� �[	�25���3�w����Ў\��:�A$K`���ӭ��ĪC (vP߮۶.U��T��]��ZCʩ�5�(3�Y�Ҷ1�|���o��փ|X�W�zQ��	b�N���m�3��%���Ok��vY\ų�	�hz.���"�* 
�`L��i����ܛ&�#�Y�*$��!�B<+.��{18���@��+��0�l�@�T�Q��V����E<X��ַ�A����T��%�qh���4�Ԡ� �I�|-��"4�+IC�!'R~��1P9A֏}.�F��<�D�ѼP}��ΰX�����Ņ��x*\:�E��.�7퓾ǘPi,38�� d`���� ՚�Gu`gx�\�0{1^�ġ���5Z|�Ƿ�b��;��}łG�!�E)q���Q��m�^#)2F��A��D)汪���D�����i)����6�p�q�٠�t?�B֬�	���5;��5����J�-���h~�,����aA�8�R��X�� �� �{יZ$��rġ��G'j��8d�$��N�-X	Vt{ �'O��4`.
I9�t��`5�'�08�|)C�@�#���Y�5�8>&f�j��M���{dt�v{=���᫕�� �"G�q�ya�sKn�`����й� [��]H�j�U��>V���O�,{�-�?�Z����2'�"���y�}d**3zAE�-�8"��ٺJ�L+�z߷����j����I�����?��s�S��ęB�ZEk�5�����K�����"	�����$ʹ�AG�`b��vN; ې$�� T��>�u���n��GA��cwn~�#6�@�6�����c�fL�$}J�ݧ1H�%��?#��3�h��Ǧ�.ś2��}�4b+��	��L>b	ΰ�w% "�+~�nY=��xc��Bg�5������}A�F?pm�z$�H�*�V; ��7���X<�`�c�:��̀��8h�|Z]Gݞۂ��z?��>M]cio1����7� ޑ�`h����z���������	������Wz;�%�ϵ7M4AD"՝J��gⲅA31�`
�s!���*��h�I]?�s%��n�����	1&`6��������OAU�� '����>l�4���7��F�;�b6C�$�/��XUa5
��nA.؄U�M��M��{u��}i w�p�*�W�Mf�����x,�NF[�j��/H�J��blr���c�W�r�lA^`H,I��;����g�`@�6�=x8��%�����?hއ�ю��[�A~���ނ�g8�+��<6��1�}��ڽR�zWZ@v|�/Hϋ�����h�����@�{w�z�ɫ�"�b��}nZ4R\40�X�[��� ��Ĺal��t�o@�"���|�(��￙��w*���n�(O.���&d��E۾:0g�K-������o ����ʶj�g��	�W` ��{�VP/�)����k�@'��6��͠��ݵ�2�.ݰ�sF���ĤЗi,I�����^��	�]��D���\�����0CB�5�>t������������w�����P[jQ�~t��U����HX9���5��O�U��ܫj!R�m���_���Y�A�}�#$�_{vz��o�铵h���[�s'b�3s�@�+�r H����F�x��a4_�f&R_� �$��eI]�N����gu���Q �;�[t�ys�Q����m��UX� cj �bn7�l�N`�\i�;�	�?k��	AY�a�'Fu6��$���U�,�{t��7Z�3��C�z�Σ����MG�E�W���!uIwG�%�=���3�&��8����,� � Q;������_�%ʚa�D!%�+�����K�#��y��;R%��Jǘ,i�p�P��c3۩����4���:ܚ�t�&�Y*�Y�D�����_U�).^AI�IƤ ,6�t��4p�m���s2�7�!�z����:�%��^צ�׈�łI�B�j�����A��O���Ҋ,9/Tp�P���۠$0�B�� MN�9�=�P�� �x��E��_ �D��~��]����u`o��4- 6QK��
�o*l�;��@oOuPJ~�AH��\δ%@��T0��^.�W�?�[�k�]p*��8�磇d�I�)[�gv�ʅ{�/i69�8(����53X��%�f����G�ʂ�>"|)=ű�w�+�6�ۅ�_�Eu�Q��]^HU��+T�0p"���&U�y���ǡ�q=��-P9h, S�X9ҹN�X��hQb_v�	�'���8�ؿ�����+B$*���7���@}#���>�uq@ų���%�]ז]2oO�e�b�P�]H��@��
���e��l�bS~�h�V�D_��$�������6�zl[�]�#��#�S�1��ƛ��{��Y�П�T�?�},��$	��D���3Jބ���� H��9!Pe)a�S_c����U�� ?�%9�������L��z̃��"qR�7�� ����ų~��[k�;�7�$L�5�_�>�ˡ΃T���ثN�~��܎�]J�˂8��v�� H��?��}�-o���	P��3�ˑe�
H�+���b`�D���UN#�EC��!H�u7�i��CeH�S(Sv�Ie_{��.��DT8ދ����a�V���5���j�ij^���t�K�P*�Yy�Zf#�P�U+_��^�J������Q~1&��G�+"��q�9Viq0MD����"�)1X�(�_�w��R_M�U�p����G1eh)���EP�(߮�X)�� ����k����"X��w{69�қ���� TI�Z�����LBWh�#��[	�W|[a_I��"�r\-�m\6����s�c�⣘�$3D��ϓ��l�e&Џ��bt��:�J�I`�b� �$Rs�� �]:Ԡ���h'n3Jc�c��T>a-� �j���?���X�.��J���QH��*����)��2/e�.z�zҧ;SĽ�v*Y�,�hHW*�)aH���4�a��#e�Un3�K���H<��l\��7�X��RWou<�5�&=�ʯ�8:Xㅶ��蓣�v�¢�c���د��:�/ ���_.�����^[�.���H�����)��E@]T��8���U�/VP����-�H����{nT�E��#����X��87'V]R�@�\5Q��EӋ���.-BVMu�q��t�"Ĝ�xi�>
|�K����/�^� J�|�J�?�K�\��:b������m�V�^�0X��]��O9���Z��������[  C	c�=�Y���Xd�G���D�:���`�m�i�)���/ޏ>N�=[�Ꮛv�;��%-~ǒ�KS~��A�ϗ#� 5Z�t6�ăl�/�06M^��O�C]ݛ�Q$�|8.�ǭ%��p���~��߿}����x ۶翉�o���?4pt�k�8��M��s�h�]f�E�Eu]��/�5�����)O��k��c/?�������j�҂�T>"��>{a�|�:0�!��|oL�>X������a��7��5�耶�i�#��POtvO��� Ф{+�A�=�(�t���ڣn���m���#�k�\�8��ڮ$�NB+�H+��E���mQ���ΔR�J�;��w����}�N��k\�(��f������%vi��Tw�|g�Xf 5*�@��� ŉ�K�qn�Sn���D�m!�9��	p��Ѥ�零�@CU���i}���)��Z�e	&�
}���Smt��}RP��\�f�G��o�Ӣ:����������-��������K������aˢHi�j�D%��o����h;=�crK���¹��w�bʢ��Zg������k��nVk�^��:�`h�/EWu��^Q���gU%]���I�+~���&'�H/��	��@Ww@���V�O
)�b=F�S��=HЗ��l �-�2B׌^��b�ZeuF�$���`l/���3�+x��i�X��&jEY�bۚ�3:�Nxa�}K���A�2�;��b����y�J���ZZ�!<���g�*ķk�'���.��W�<n�V���x4×���F[l��p ��t�GڱU���}��{�]��o?�������-`��q�����v²���_I�s��+�� ��+#�c�6�~o~o��Z�~��3��R;�u���oyk����~���wN���D;�mK-gLg���|���uu�9��²'n�eS��+�)�uJ-b�y����F�A7�k�?�U@&B�zা�O$��#�Rl�.`:�F�?��R�n��W�� A�*�b,9(���l�[rc|�4����,z����Hb�h,�z�E\+�b2�S�s�X��mYT��ߦ~�0��
�<�Yz3bd�_8 ݩ:P_g?-ݕ	Ǚ��;���n_�������۷��Y�{8Ϳtv|�f�&�z_��{W��~zE}�.
'ł�=��寉
}�p���6��e��R=��ǇdP�7�H��	WJ�8�.����3�%"�KLxl�[��-B��u��d���b 
�()��m��E����0��/p��8A��v��).GL������d�E�����n@�NU �!��U:`[�.��X�q��y�O�~/4v��?�o�r�;�R�[?�,�Qɤ�E�Ƀ�|b�q��s4$��V DǢ9l�����i�mE���������?�*����� W���<�) B�-�����m�<���.m��B��]<F��ȃ�3�nI��W��*09�1����ZW����5&��70$��{�'0�:�2_���mP������wka! ��y�R�Ws��?��#@�i�)�>zsLTepY����c���P)����DF�+w� �H��B�������x�Lԧ/�o�L�M�u[��u����%ܕ�~$��b]}k�o�F�.��q��޽>���ɵ��/i7��xU,^_�UcwԼU�I�_�r�3�MY� ��.䤺E��6����R"~�����31�mzV��\Yg� �,����0��7�,Vg��E%0M�0|�Lv Tχ�1On����B�3�c�S�|��~x�3\m�f�����?�1�eX���Y�ci�ɠ�мP�πu�s����f�b�D��1b���Y�Q�F�rP����(?m߄���-X�o.ry���bb�8� ���TØ��� u�x� W�~���/�P�ԃ��Uw�!��t�b�8���`��]�C��H4m�+@l��t%B}�L�'�[[a����Vl�Q�gF"08�9e���6��/&�����;Y�oMi���G�8*S�ig�:��d����`��%K�Mi>{	bjy=q�ŇA} �Gq����d �1��Ԕߔ�G~5VJ߃�IM���	��;�S��>=br�&m��*�D_�۰ÑG���9W;�OF�9�,�_P���:�=���ʋM�Â�VG���-�E��R�Ɇ|�c�{��yW��~!=�[/�;V���x������#���Џʅ?��wt��J��z�э3����'��/���l�u��u%�=$1����������,j��$XӹV���}�Tk�_䏒�t�q�l�.���d��Œ�����g�_�Om�{��F.(�"Hw�2��C��HS�	-��� W�1 ��ʈ�/����C�Db�Ī� cL�#s�؉�%5�I* �?�u��/�d9�v4�L,Ę(�#��Kw�  �3��w��f���S�*{�	uU7&j̹PE�n�j^9��S1�P�i�gg�ߪ��#�P'���r`�Yj��n��۬%]��d\�ga.T�=#j^p�9=��}u�b�iL-�w�)�MU�-������Q3<w�Zb�B����"�]]~�0�FI��{��$��b'y�~�r��C=���@�,2b`X�1�R�6%��P]�6�<�apls��.iE�j���mn�����Ǿ���<Q��ҐUf���rK ��59C�q,N&'�]�%�]<�)�M6��@��3������0#�����(j��TV>3
Z�p�]�`9�!_�X��NO5D�*��I�,��H�Jeem+/!х����h�
܍(�����N�p%��ׯ�䤻���z���!^��&�@�*�AZE�҇II��Vol�m�μ�G�bu��v��MD=�^���ֱ�l�Lrη%��h�c�F���ӱ��An����z��~��8�f>��d�0&�6UI3���"�]�nKeLj��3m媥��M�'dv�����2bu���M������-�jӈ�ZH,���O����V��C���J�����~ʰt�\���wL5�n6���h�2����ܦ�����?x��"{��q�l[��oM����c9�L�K��R�~��q]�*
E<�.C�fe`R�;g^��>HaͿ?-���=R	mVF���tcƨ0��W����z�޸L:AM^�����8l��m[�:f���2��Է�����?.�5�+Z���#`<1�З��~�4Z��j�L���T�N}(y��3�<�+y tݩ�~Js]J�Sy��+�s*ړ�+>Wd@Ex0X�\�SU�o�����C�U�P4��Y��E]5�"��^ީD�Ds6k^���n��*��������I\B��l:�<c���d:A%X�O%ʧ����������y��5ʤ������:i�k	��a9A�ExQ��M���&ou�TmT2,�� u�NE�A��W�F�.n0�q�q���ږ���}���BE;���Ib(�b8�d�*cTf��A����ju VЯw��{���@b��mG�r�3�2-�N�� Zt_�3����l��8������'�
+l�����ʸ����|�#q�0f�j�ʀ`�>�I���������lt���5��|FK�,1�3�#M����GW?�c�u�(!�b�q��\�O��7�. �|��`m�(-��m2uu��&֒��d�ݦ]��x�[�r���!�d� 5���+H(����!G�o�������=z܁掫��=�J��S;�3.���� �k �D�v�@�M�Ѣ���\?Tɦ�n�P��y�(�hNH��EP�\ޭ�Z%��ս��|nN�y�;��]+3�F�������y<��կN>m�lHe���^�[�w��f�5���2�_�^�O�m~�ɽ?���w� =0��e� ��F�"�=���ޒ���?�"��=.5��3����"3LG6�°�\֪��sI��%	���B�}c���Ķ	H�@b�j�'a㙃&���g�@�į�RU�ʋ��c�Zz�c?\�w)�&�9m���,�QJRxO`D����bEj��1��~7�X���59X�WD�������um�˃ߴ^�獍?�/�(A�\��e�����4Q��b�������:�">Wù�o��Z�$K?���R���T@U1J;�96c���%v��8���<!@X�N�*���
��j��X����d�@"�����, u}��6)�)FÛx{ܒ�Z�?ӿj�j�R���ሹ����b0}�&e�B|�<�9l���m�zY*�J�`+U���I��) c�V�`wp% 
��qa+�,!�b��A!.B�:I(W�w;[⤚�x�����J�5�	���O���f}<�,��� ���_;��H��������0�	B��l�̬��PUԍ����" �Lz����*��F'}�<�H����	F�`�Xj.Hܚ�M�U��LavR������DD�F���KQ��J?aT��_h_��ק�y�ݣ�;�<Q�<�$�G�G�����\�]5ɏ�ކ�Bw�d�D�����J^�Jz��/�N]�$�K��i�.)ew2���O��f]���zQ�Ѵ�%��Z������nk\�7�R=�tw��P���$=�F&�'���E��~���!	��d(K�yn%'Iv�d��5>�DV�y�_��������WzSTqDW�*�d���s��8&:V7^���aq<=3P�uE%�LX�q���ș�f�|?�6��nL�n5C��?�\{�s���cy ��0i�C8!x�_/D�H������d�D�����G�0�`�"��8���	���q���:��.�L�)>Y�J�#�B��9��}9�;.�<aL�׏�GP�N���U�J����\$?�}�-����/%�#�r���F�¯!!�My(�a���Na׌��bދ��>3w�	��/���C��R9LJ���}B�G�rx�f���D�i*.�0��k��W"E�Lڞٓ�j]���� �xz����+���l&J%0��A[�{Ĺ�
�^�o<1TV�er��P~�$U��Y���i��YD��F��x{�}z?�<�����*.̾À�s�H�$wmGo�9�PU@u�Ҋ�QA���$��g���֕TN��l���ܓD\JùP��(@��#�g�3��ecI�W���h���Hٵ&D;�]���1v�D�&�T�d�s[hU=�r�����r\]�6N�:9������SPn���3}%݃D�ӡGzɃ�|�/�yT�e�<N!m!%��EL���jX�Š�6���<,�v?3.���S��	���Wz��䭧��ӺY�
~��{��G��5�:�Z��bu�o�Z&�:�H��������H��~���@r /��eEk�0/H���T7�s�6�b�4W�|%="��l6�O��I&z���ޙ��+�ߴ�N3�Oyo���-�����%HN�x8��a!�3�S>A,��zتm�3��u����8-�b%-q�@ ��x؂-�%�eT�>��B"���_Ԓ^�l�Z�骂U
��=&�����΄����󩟘z|��y��P+LAd��n�c%=�����0���g��W�������mK3�T�7���M�=����B;neh�MNCK�e��__�����b�5����6u�qe��t����`��j���@n3>��[�~\�������w��խ�f�iQ��|������`�*%�4b�^f�Y쫓�-9=U�`'�;�8J����I5U���_�Y��7�����Ens�t��K9�� ��6��w�'m����L+;�&���K�ܣ�W?����P��mX�:��է����q<�90�LF�Z�1)��%���smw����Rb���s�;�BP7����T'70��-��i��c���`Љ_��*��� ��_��MJ��1>�X��ۅKW)�p F��@8�@Z�%��V�7�ޗ'7fW��U�U�/ u����NC%�:k�g���J�Y�%uLYG]��ab��/�]qp��� (%2��O�P~WĻ.�B�����*�����Zۏo�R���w��$�\+&Tb,���W&1��>�]-{m�d+ 2<���5��s��N/�۪�p��JƁe�Ku��*L�	e��g��b�U��j��A�6�@���H�'��;�O�&�+�i^=�7�nRF��ܰY��z���mK�g���9�z*#����+�S��]�]uW�<{�W��\٬^�w�n��P�R��T��<qJ�2�yy��B!�ƦP,�� �y�����kl��׆?_�bF+UK,�q\n0����C�u㳩��zF����t��|s� �o�{�R_ ��Tc@x `�}(�_L?��;�(e���2���d�=ꊣ��;(AW�����84��+��_�/c� �.��$�L��*��D�v�t-q����v$���E�U�j���	��&+�@�a� �;�He��A��?s��E���if4�~} ��f[���$4�C��I�z3>-�2ރT�Zbw�$�2wtp�`����W�~Q5�*���:���J�:��ŴםWp�yv�	:T�d��`�
�'�Q8�D�.	<]0�a�� (�C>)�ŵ~[�g��#nK��g�_	\�p(��ԩ�����/`wx~�4�H:���]O{�Ӳ�<�u)��8a���L"3�ug]��r�`����-���o繸D��Bd�G���K܋���u�i���'�fAz�`�\����_�x_h�$���۲�(m���
_���7��U;��d� Z+}Q��A�~a�߄j>�\�s�=�B
)G�l%��I�e*�(-�Ew�r�l����f�:#o���g-�tNP	��j2�����������
������W�Oa���e�5���AwC�yRv�T�[�ѥ�a[����-�H��&Hu(S�{-'��谵���_�U��5���$����t�^���WJ��rw[��e�.���n�a�<�^N ������B.��ns�9c�Fu�6W��JRFT�Ol>�|(�8;�O(kh�}�Ɓ�?+�P��f���#������Wb��M,��]�"ex��������*ݒ�S�>D�a6�(���4{�H�Y����Ϛn���}ˋ�P�+���ϐ������Y�g,ʩ; IJL��{���X�]�s3����a�*�n����WD���p�M���vT����R@�O�L���c�O�ߚ���L�f��o�xe���� P>�	�k��a޻���B��\/�_���K2���4���թ~���pe՘�� JN�0��_T<^��L��8��y�Y�2'.|���UZ�jZ`�� �E��4@�w^Mo"��h +���c��G���u�0���N�qE����Zc ��e;�N�`
���3���t{��-6�|h2��]��� 0�5�=���h���;�1�U�|/�i��5l"wԣ�H-�!΀��W��jӿ���(���&��IN�j� i�7����W$Ҁ�|��Y����V�X�F������[o���\��p:��j�ù�V��ӘK�����	�����!WP�a��Ӆ��+���*��,�>V������������9C�23�$��󀾲͛�L_ڞ�ů��N}^6�����AZ ���ywc�2��n9�|�E�=n�z���,����י����������Y>Z�f\����[���%@�E���4���l������;TP�RO��h��u���i�� )���k%:,O� ξ�cQ�	U�_�~�po=���X�vq��{�ޓ�v�{��k)�i�~Fԭ<�Kͷ<��~�dZA	�Qe���zl����v�̘�_��� 'X���E7���#��)̌4����:�� H+�f��^��bt�J����h�\7c4���e=���IS��U0�Tzma�Z��.�mAX���XP�°i;��t�O��?�m
�pN݉:�2�%^9��;b �����כ�in���?��v�����o���&��T����� �Ou* Q���� ���4\ԢR50g)���y7�\�<����C�6f�� ��$������RU�)������Bp��b����5����L�L��A���6�ی�_"m�K��V�#�?!0=���k�n;����l��[�/e��əbfxPz!��4b��٘��
l$�Q���]�2��%�j������R�=��I�z~2c�p�{�ٕ���c�e������מ�����Z`�i.�n�Pg��H�\�>0��������ｶ�1�Cv7<��T�������rõ��Qu�B��sA���6U��ߌ�f�3���>p>��?i�|&��)����Yf�vP	����t�*-p� P1WD~1P�DTK)�wRYh)�b��="�J�6!��s��S^v���X�|��Яtw��-��X5w)����T��5�J<>-���<�IZH�a�Z���e�Qw�ǁ�V������i;���<���p�@mH��7��p�쯅�=��JH4�/����I�0oJ�C�P�q�&��x}�!\.�9QԾ���Ay��:n���h���Ö����C�_O�	b�H��n���{��;�L�%�WJ���{6������2��mꓭXc��*sc�� �b��=�@�H�o��O�o�j�W������o� n���t� >��T�d�<L�u�o;��J���PMi�W��Aq�V�A�h��V"w�r�_�Ÿ��+v�����*ӠD�<Ǚx��Y��;ѯ��4���S�n?�����_(�~.,��w|u��y	�UIa��8���)����m�n��<��79�.��씁��r#�(��xWu�N����]]A�M�����E�����ݕ���e�تG^�����(���J�O:�|������@`b�"1�Veo&�=%;}�˲�{�0����0Vjz�kr�듞��^̀�c��_���m;H�?�.K1`X5K�1�i�%��W7A�J�IצI���� �����R#��;�XT��4�[�ti��7���;/LE��D�:`�l���Le�{� Ư?3Ų�k���iA2��Wl��jBe�\�.����o�t��a0k̢{�n��6]ڽ�� ���"���o��լ��-��ڮ��_72ݟ��O�-��i'z�"9 �y\�EUP{�c�n7u�:�xS�gt���ߑ��n?)�Z�_K�ߦ�k��cE�l���H~��O?d ����`e�.g�g��~����J~� k�][�B mj�jL�wTQ���_����ޓ�}��}�r�Q�+�L�*%B�Sfz4,�>�F�V,������ߙ����%���r�1ޫvu��CA�꾒�����"�#:���	�oqTb�9ջ��9���|������7v�~~d��zO�^>�C�X�K��X�b�Yh(MN�`���>R%Xg�w3�83�
�:�����q���uw�?���X�v~���a>I?k�'!�s����9ѓ�]tKηo�D>�����4����|�s�� mn���HZ�m}�؉�Pշ��m�TlV�I�L̸�������P�*B��t1������L�O��3��q>V��9���-11І��O�ه,Yl"��5 � <aT��ڵ��i�<x��w0��2SH�t}Mq��8����{3�=w\kA;�W��,ӾX���B�٨/�zW�q]��/7x�8&usq��m�",�Rf&Bx�z� ��h�c�xP~��
{ɢ1�/_}��!��|��������`�n�`.%�у���Kc�ti����-�����@�l��~�g:~���{?���D��%2 +%`)�w��O��k?SAf����Iw�q����5@5e\zn.�VS0�a��,	<�������0��p�>c](��*�r�<E����`g�$�８�҂�!c��s��B��z�2�R�+ ��%�0 ]��ĸ�Y�ǀ95 ��-��뷈*؁�Ѽ�:�������?_�j�>�Y�P�y�r�
��AK���)=P;��Q_N���I{o�RmKY�����C�l= ���$�_��_� &Z�ep/�Ҍ���{Yk�� �-��8D��ec���I�{ߕ͏��G�J�Tę-T� z2, ��n�C�O
\2�yQ�w~���-�+�	k��� �����B]�S�k���a��Z �-�զ�{m����Ѐ��v��� �<E�
�]ʺ`��K'�u�?�(�&�+E+���(��.��A�ݝ�t<���.�B���d(�5���V�\]�(����xt���^����x整qs�.;,��>�BZ�'1��K�_��NF�)�ﵝ��<��y*�2�.ͻ��3B>+UjØ6�k�5�!>KMR���`o���H�0���)���4��w-�x�A���������P��8r�����ϋ�_E�m�ڭt߿�va�<=�h�G�8��%��V|��#oD� �9S���H�@���(l|�%��?c����<� �����U�zz�}���ճ@��J�fYT�%��]�"e���f�=��3���#P������>MZ$�L��͒�U#ܮ��p�ss�IE!������4�j���3��y3ϵ\�2���S����M��׿6�^�.@��������� �)���<.\�wF�y�=���Rr���'������芒����5�T)x���Ź���ٞ۠j�h
�kU�Ϧ	˪�b>To�-�-1��0@�IWRV3��\�{'	��ٳ���7'g�$����ג�ۏS�.-�`�j�j�<�H�
��89���
�G)�5��,�����~�nUX� � l;J$w�K����27TJ�`pxֵ�5&�+~׻N��k���$r1��7��W��E���5\5#�T��iܷy���.i$�������l_�ԋ"��Km�>�4G�qnHh��R��\�1T��i���)��zT���@�l�py��V����)ȋ��x�a������	����P�"K���G�R� ϭ��y��f��|M:\��${L3T�������zz`í%3T��c+�Q��b��=��]�5M曪����� W���?h})�T ��5�70��,���{Zֻ���z���n<�t�hb}��Ԅ#�ȏ���f�i@��WUݳ��z�8�N�Ut�gJ�������������t�S��l�H����
�XIw9�<b�������0��)�����:���[D\t� Tb�aҼV7*�>KW�J�'�o�c`�&?�{��-���y��#��9����y��=~�N�&���Y�\r�EvxV��2��e�5Vۛv`_I�StL�-�,�*�m��� w�ߖ����p�d����ǩ>V۳�5�5�\��J��`�#��r׺�:d)	(zI�l���n䕞��YmY<��s��ސ�]�g>��y�^�zפy��ή簎�t�Z���{LyOEIy������M>;)�,�Y�)�L��N�� ���T����fv
v�V��b~)Tr� ��O3��n{$=����>ر�ͱ�����ゴG׍�C���9zQ������+�@S���"J�wi�b;;j�����Ca��s'�љ0W�=������lT8ÿ5i�o����E���^��˦{��f ��~D�"/sI�E�y���k
�r�'�]-��P���
�Xx�Uc�~�j]��aWw��9钦i�m�|!=P�o�N��y��荰:(���� � V���Yƛ��S�a_�n+"����6�� �]�pp-��?��,~ �Ɋ�:�[Ym�@#���2����]\[�|��� U����~�����0�>жj�B���P�P+T�y�o+�����]���� �i`���}��1��I������j��k+����}{�X�W@�����I�D	�ŷ��-Ƴـ�>v9eqܹ�x��p�\��y�Ϸ�!z8��]M���|-Q��+:�j�C1���u>a��s���-kj�4�����+-T�� �H#��N��T��U찜�+��Ws<�k���-۬��㢝��R�m�f%ͣ.�]�8�n�\�_lϼ�X��k�ˆ��}^|���oL��{��\V�?�zO�jYI]'�V�����woJy�ؐRE�y�N�i�H�?�)�}$՛�
�}��WXvJw�g~pK�N[	�ҪB��ub�� %"J2uv Ԏh�������clq���x<����ӇmY]�.I$C�5��}h���q�$r��zGߔP�'����0�ۨ����M?ס�`��*��ü5A<�/����Hq`�դ�/2 �����Ƕ��60��E�����j��`�A����#��
�W-d��՘.0��Y�TǼ둈RA,���M�&����C������|��<o�'�iKO0��-bn9Ww�x�5�X�"�}ͫ�6�ڀ	/�(U~ݖ��2�;�m�~Z��C��c��;��oE�{.����ݴ,����R?3�NcpoƷ��M�bH�#�(��1�=��8Oη�S6�H���c1r�M�ύ�76���%vS��QH�i55 �l+�4g�gy�+nM��C�IZM��;�V�;k�T��z�ch��:������Ü�����ߏ��N��Of8ٔ�ʼ���*���m��w+��w�j��
T�-��5ס3��i�{��Pi��Q'Lt7�q�xvz�](��f�k��Z6�cf �Q����<��h��[O�Eo��y=]�_,T��(���_UU�Ƙ��vf������~jpӃ� Ug��e�E�jƟ<��e|����u2�����-t�nc�M^�1	�C�&d�� s�(.>����j��'����u[��+���@�5�"-��7?O�1�{nz��JWPiw���z[g��O���0��n���8�B2�ew��gu5��BIMu�F��V�F�j4Wq��f$XQ�W����W�s��5z��HB��j� �J����Y4*�u��f]��� 6��J��P�����ߏ���:��u�:�M�"�3Ԧԯ��������z��Cw"�s�����+,�y�7����R��Q�:����	�$`�Xf:�� ��\��xJ5�T�9�m*���AHE്2�u��!�Hz�d�ߜ�I~N ����v�5V�I=&+:o2�]�:fOF�z$9��d��N��a�z�j,Be���=�>���#�F�fn�
���1�՘g�U��n�y������gX�l?Խ�BDR�vǳ74jK���&7�W6������_I^+�`��BC/ k~�)"
Xl��Ŏ=r�)?
:H�pF�m����O������g��c��Q_�SB��u���:�?{�T�R�k�1�w��(��S0�=�"���6�Ľ��g�A���-HJ����qW�Rڧ�~�=i���T��u3o���T�^ ��KNT�2E�1�+H���{��i��a��M۶�A��@e��>~W�S=�F��k����{�9G����[!=M0T�(��-)'4��`�kl;SW�2BV�4�I�I�}m���N@��~�]���,=&=֘�3^���� �-��{��#ž�!>ˈ5�2^�|b�]p>]�ǎ�T��I�mA��1��t�B�@��{] *����@�Q�LNR���8h�,��M%�ց)]�z����9"��DXiJtr�sS>-���:���Sa����Wl�)vK����~�5s�["�:����j�~C�Y���i��J��*ƪϿ�T��2#_���~�_^���[E^�C�LWE�y��}�oO�+����2D�B�Ű�?L@u|H�`�t��1���8.�%�	ѿĘc��n�>>ǆz��6�K~ƀ}C�V?M����0�_j��+N�@?�[\]���,,�֨1�'��H�JV�_��Qj���D�gQ��V�y��x���-(L��$�+�宺�i�N6���������O50`7�x����TI#�ɒ��P!����_u�Th�t�[��yC�c�6%��zX�����!~���`���OM�s�"F��r���������0v�������A����LW�-�|\�z�=����fb��W�(>=���BI��ef�i��E�"�ܞ��WB�M]�I�=��Qb`p�^��w��)s�*�9DpNn�Jnp�}�C5��Ŷ���Wm�%�� �X�P��� n�R�</8��Ѱ�T���J�b��b��V�w��Ѩ��4��ɶg�a�*�l�0��S(���u���DG���B�ҫ��b��`�4�>�[�����i�(��ٳ���.�x��W�[�~�O�z����G���usC�j�u�m�t��^*`_u�CZ��ϯ�4�Wȝ
��$w��f�t�G|���{����+S�b����yLu��bزj��q�87葦էu%���߫M���e@��vA�O݁��ձ#Ot�hA�����~<��W�w@���~�<e�%&��F"L��w�c(9����K���� oE?���u�*v\�������V��*D�Q�U�9��.i�<���Jm|m9-mC�Yҁ������&�����G?�CL+6�1[�&Zl�*��a�=@�����m��'~��-��������ȑ�Yf�.�~��؄���e��V�15`:W��m�����]̷���PC��,Ă!n��u-6�C��\`�����8"��o�=�[ۛ���t�`˩?��!�éS���-�RY����7����r��ۡ����q��َ�?��!��+ғj�������+��hx�X ؑH���9�*[_tJ��ōW9���k��`HJ�;�f��p�p-i����o-��v�"U
��#��(φ��h-R��{�b�G�p��Q�t�T�z�ZɌ�ו�ꈚ����es��R�k���%�B��G�]w ��UʃV��GL�q�S� ��m��Z�d���Q�D�du�o^	�D��3�,�����k�\D1�:�)F��4�0|E<ʛ�ԇ��KI�)K=��5"ʅ8�D}���+�F���ϰ�GW���tZ16��_y��:�p�ȷ�t��l	��6\>�A���N�7M�}��߇�I��kB<��Sw�6&�a��Yx��N��b��X�(�I}�ni�7����^�e�o3��. 7<Y�sy�`V{B*����ӡ@�$�y����'9��:��,m]M�o����yĞ�
��2�=��*�~���~��� �880:9,��>���@50��P�:�ql^����~~߭����!�d{)�K�u�p�i?9AH�\yj�/�\�AQLr�U*��1xO<�L�e��BcҾw���t�����bQ��<4�S�y5^� 	�@�q�K��������}-9����t]x ��L:O̽����Xa��_B���E\w�X���;-�V�ė�?�'`:���e��_SڸƳ��d1��9q��`���;�6�L��0�.��+vk����;U�.�p������?ޟ3��ՈM*	HG#^ʽ�ͦ�� 5e�Ӷ��F��$m��CFx��1��l��7�'��҄�����b?p,�U���~��$N��wZ#��_o�-v13pO�D7 ��&�Ӈ��^ӱ��T�~�|?�սb�:�Ѻ+�Ua��g�������q���;*�L�7���Ȱx��# 7*��J�s���w4���Wѩ��$���)�l"g�D�@���S`������Z��0H,�����)�����5��DC���/"E�:J�<'�y���ߨ�2ߑ�q��
`'�EF�2P�4�]��>�f��w��{_K�=�E�m(>ѓJ���$�`0ݶ�=e�/�^^�Ʌq��?P���49g�jW�H��$Ų����c��u�p�%�5J� a����m�y��e�K�͔��]"���-�eZ���h��;�K	O���jw�w+�b��Y?2\i�)ѬX�F�~�L
M�IQe;���;�s�1����4i�`	?�`���[�90*����EwB��+9܃6���"p��W�cC�G�q�Gw��Z���ƻIh�Usb�2�>��fH��N���A N`��AJn�2�:�,W���2<'��6kL���m,Z,׭?�S�HJ�ס�^4t�aXҟcU%b�bV �f���D
]��x�t?Vס��a!�ME�h�'�3���(<Y�Oj��dR��q4DmSy�k�����$d�-�V$Ll��#S�};� ���]��M���T=Y4~�5B��C�z� W����m)��?�����ޯ Z\�0g��K[�7�{�:TL����p��\1������F��84L����Kb�Ҕ�i���ş��X(�v��+����&�?�,*�%��D
x�0��B�mwCzd�H"�4�*[ro�)�Wnd�ۦ���\B�yf�yc��8{�����y߯���'��;ݜ�P�Jk���u�uWF�)����r)?�<C���祧���n ��_�QX�s$V�l���������
�yI�ޏ��L˟��̆����瞘3��a ���V��S{,Ϩn`��t��J����g��$��������:���㩋/�a��i���y�[�Dqq�� uH����s�J��s��i>v��-$52��M_��I��yG���(�l��Vʶn±ߝ����2kL��ȟj�N�[����E�UگV�"Z��="�Ĥ���>��D��<g�٣�gk� 0R�������2�|4���7�_ w��Bw�_�&�~�b󸩸�����D�<㥩�������g��gG�[�B�u��I�=.�Ӫ)��g�	 E�S���j��V՟�6T>2!�q��#~�F�WD��Ţ���W�2w�O����b�-���*a�	�~�_Ďvu� V4���%��1���Eq=��Y�D[L��ۈ��O����G�ia��h��s[1�ȑ�O�T�r���D&��y\�� �#K�ERd�w��*��o��i�g[���=�V�X�_c���qTO@Jm�Ĉ�[���j��c\�Ѹ�J]$�ޞ�%dQ�]��JOT�T��Wrq+�v�^�+�-�+��vpN�OE�U�5y;\
�vt�R0l���Y� �=�廞N���U�@�-��
��X(�c��@�/dE &�D=�0�;�pmb��8'��XZ�^N�1C�`]Y��>i�f0��Ey���^�/l�N`�B�3(��)W*����``i��s =�§I7��;��n� W2���Ρ���gd�f��D?X�b��q��FZ:\@����e��7����� ��f�����P3�,�����|S��&����C����ЯYu��|����ov����ʢ%_,0v�d�����z�H	�*�ZyE��X]uV;Y��3h�y�+�����=�w}
6gZ+� 1˿�N=pI�Z��f�)���'_Q[��g�k��Wי�Wi�1`d9ZIw{�������$0Ԁ86@ecQ��>7�k]h���lqo�o�}����	G=.i;�i�.�yNP��G�ո�ڰ!�mA_ęo�P�~0��T�;��N�j �� T�h��b{����������+���`-
�`Kt�J@� ,��iT���C�A�ҷ��X�N;���)B�!���B2��X �e|�X������X�#���9h���U����1�Ĵ�L�%Pt��@.�ޮ���_+�T�*�9`�}���%B��I\#M �4[�+pVU�D��_'(�[H����>�i�=l���M2�p�I/���*�[HI�J���Cg�gc[`��#jH�j�*��$x�E������2�n�"Um�B��z����&�AU��6Pm�1�{��#�L�l/�F'ߐv=�p�X������<��y��=�y���j��I�2�g��;�jp��*K��W�.zC:;�9��L$?O��]�g>���6$���~wݪÀlR
�ZL��8YȘDY�ߛ�/Lύ656�S~,Q�W��,���
�����Ӈ�n [hf�����Dލ�Lky�O!*�X��a�N�`kbι�^�g~�F�C��Z0R?��F�7z��N��o͓i�����'~�4R�W=�G�*��g�h>V. ��?�A��Nw�o�����j�l/�	c�i��C�&�H��%/ eӕ6}m�ٖ��E%�eC��n��O33b��Ql�k��%���T �`��V�3+e*Vd�t�g�Ok�8��@`�����UѠBWs*�Z�s�����} IqFz� ���^�`��q��~�#�nyT5�&�N<�����C*�;n��c���~��+��)?��EFiW��yp�]
l���>�������{��z��|zy�d<k��ߣ'}�\��8]�;#׭�����>;&�ׯN�a��xc�={�ua*�������k�������K�A�Ӭ��Ӷ�C+t9���κ5�P���50������Ũ���ϖ��r��]�)���\����(��?(��K�x��o���Uf��;O߄�{��%�n�%Y�Y'Z��\��@E��"JK©��ϝk����_�2�1�rW��0ΑIp�Q^����5�-2�ᒃ����}T4����1���Q*��}{�w�x�=�c�b@@{��-�cZ�ֱ}�T@�n�:ކ!f<�"����Ç�1%��U��g�*�][��3��+��%��>�����@��Xc���_���6�k9@�Z��.��6�j9��ЍD��@��������QkcFރ�X۽����
ծ;�����v���.O�
s�Rs*A���`��K���H��L���rm\ ���X̪8�2�uu;t����r�/Qe;�*�,pl�n]L�
y�������4��&�� ��9�93B���!6��{�H��Z���{���/�?L�}�c��`�^��uc*>�#�=� ��\�z�E��b;��҉a�͠�\�� ��[7&����\��_~������?z��
]hZԋ5�H����(/�0�Dg�)�u3�ƍ>݁�9/0�vH�jb��;�����OX=�Mim�n{zW��5 ��^�}���������'՛r,�~m?��u.1��n�m�A^�k�2��36�`��`���_�g�)�$3Nl���v�X�'�~v��b.�k#��4@]͎�V|s����/�c	n��A�|�z�f�kʄK�g������"�
 	ۉ+7EG�ќ;�U��'�Lo�W�
7�|��鑵/�z:}�c�i5KaU�e�o@}���;�]��M�r4�o�7�j�N^5�
���X����#�3��H]��L��E�ձn���v3��Q3y��]N���4}̟`��4�ZXL�f�K�ݙ���"S�������{������U, -T�+.	T������cF��ߺ*���w���H�Z�K+
�mT���|.\50�������E���{"��M�r�����t=7��p��[60mgp� D�jz�na�����.����Ed�;���V0����]�%�M�g�F;v��dy���C�!���� n��y���flth�\.��/1�:��q��u�=�n���~�E�Z�T�^�h���4��]�vTs��g��w��E�gX���o�.��-��9�뿘����ݥ��p7V���x�y�t�}[X: .s� �*���o�q�������[V����J��_�M?"���SwJ�h��9�72�=tuj����s�F����	�����}�:�V9�}�����%��;�7i���_��ڇ�,��b�&�3�S�����>� U���z#6`� ��"��uoŎ,�D�na�b�-��s�:���D{�58`�3���d[D`X��e/
���;3Ĺ�w��F�J�c1b-��ь�k\˰ž˂�z��P�,�������l]y�}!����c��c�2�xN�2�nGV_w��T�Z#�٤��"aծC;��#(��F�o������̨��X\����+�<m��̷w�o�c����B��w����J����Iv�l�>������������ϑ�[f=�|�}N�.��������8-Ĉ��vR�σ��EI�{��=ABp]��u��!-J���zp�S�W���[ r_�|�ۭ��w��r�d����ڮ���Я.�W������x��2pu�
�6��51�b��y���-��(��!i[V+�M�����9/P�s�R)��'����)���O��F``�R��1[��<�;�˗A���@ԯ�����j��ˁ���ȣm�*L@ʝ��W��*��r�fEBT���e1��C]տ]u�bbw�����Xc���a��0|�wi�P��]�Z����³�(,��������c����q�ms����}Gە�[�u���v�૟��897C�A	¹Ɯ���[d8��ȧ.?�`}�Zc`��O�E`��yS{9a�U�e+z�U�\LY��`��W��75o$ �j�t+[����͗Q~5�j��|�Pz0-t"��F�j�'�12��8��
&�N���Kl�LX���ٌw����c!�.l�BL*��J���V�=���:�*����-cv��29x�ccB/  �����B��Բ:Әg�9^�_-a+)�헒kunj�NJ����������s*�YP���		�\���>S�F]ME��qU9UJ��P.}nk��Ab������m$�����<zN�2��ل+�ހ������v5 H�(�����< Nb������ kc�E>.����>�t����o������3��\�8�wv�����^e��Tb7IN��i ���?dZܣ$����؄��RQ��ٙ��fw#vl9����zp+���UCM�q�� 6�(4
3��G⪪á����	xE;���3V�u�.v���-��k�ݕP�(��e�8.]��Eˋ�g��`�D�G��2-�]Q�Em�W�|7u��g��A<����2>��Ѥ$5q���p���ʁZ� �sTuq���rU���^9���2�X,j�<cx��d�σM��zCJ�2���+�޵����p�Z�t����j:��-��}&��>�����n*���~c*��$�p\�]K �R�'D���aR�5����v�͊�v}jc��d�1�N�WpTp�XH��m�� �*��[�MQ8�2�J�6_�Rwѡ��7��;{�}3��#�6Ϥ �;`�h��Z�K:GW�v�O��x��{�R��h[����{a��}3T�G�6�PS�1����8~����gU��ms�XR�.���G�i�H��/�dgt�������g�/j������#�\�W���:�&��Ogۆ�U/�΀��&�K��lj��E��\��>��.<?|$���1X\`ɭ���`v|Yڶ���쭉�/o�u�h�S${>%�������������wkq&�c��.^&4o����p�����"������Ex������/H�8�'�eҤ�20�]^���̠��h��ʄpu���q���]�Z`ld��ܶ��a���{%Gr#Kԁ 3�!�V�l������Ϊ��+3� .�q��,M�ĒmH�YI�8܏�U8@ ,@w��}¦5�S��;$��h�<��񝱞M@�rz< �=�E��� 0=�f�v��W����S�\ƶ򐌠���������I�xr�T��"���k�����D�q�}�Մ8
�5I�{c����N�I�����w�P������#f���%�*�zѹ�wʏ-��T�<ָD� ⻲����Y�N��_Re�Xp��"5�<�̭���i��Q��x�Q/�ԅɳi��hA�
}DV`a��߽O�Zr��>�����L���D�X����0h�v�zT��&�s�{���w��`��wǺN�-�s��ui�|jFB�db��"����O�g���i�վ�	X��YkϢ:x��d^j�{J��1�Jjf�e���X��qZ��j�LL����b��9�Za|[����w���ݫ��ze�H��� u�4�m0��/Lc�9���G�j�Э5��q��)Cb��\����V��f��r=�Ȑ�V�g&~6� ̧�c;�ۑ�����p�V"�k�~�}G���5+Zk��p,�u~1�1�Z��*r�G ����|(#�a[�ږ�Oڊq"[	�������-��>wJ��� �L�ZI:/a�Y���W���f��X�|#i)�}�����?��4�]0�>@�BZC�����$C����BM��^�SU7����=��������j�@�-�giS/�9�Q�㎭��Z{1���A��q�{��_%���G����t*��GeK�Ico��h?@j�B�1~>���΄��$����q�����H�`{��2:ZG9�ɲ׊i�v�j�M�Kp�dܹ6N��l"�ÿ�N���չ�U�%��;L�V����b?l?��d����y����#�X
� 6K��j*���K3i9�((<ͨ��)���W*;jl�K���I��nG�m�@B*�I�I�EN��E�o秣�Q.�3UC�vR���l)U������`,͸`��1��{��Hd�M�f\B��A�aQ���Rsq�	�~�0P��G�<H(�TK��wa�u��7�u�U��"�8��N�����=�E�{�/�AL~��v�,�(h�{��,��J/�3%W���@�r��'�s

�U�j�N���Z�%Q��iR�^���G}�lB�r�Ip;��>���6�7���Bm��d���i����h��T��~o��$2��@��g�^s��8��D�LkX
߃Z��jؘ�r�'�?�6�����Vb4\Y�Sj��[��e�X]}��jKH�ԇՈad�I��S�z��x��&�!<����5��N�U�@(��\����/��<��Q\�.*$���6do}	y�㬦j��1�B���$��"L�V�{1)܏c��N�*23�r��,����7�L��(M�iu>.6�Exa|3�]&���`s�"���G���Xk��и��e��{+
��za�����a��gp��3���K���m]��B��~����P<9�k����  ��cE��"�'�k�Q9����O���(�:�Q,ˤ�0U����M^��sR���/fm|���U�����H؀�$�~�h�*T��".i��&#�͛LkF8
�b���b"��L���Q>�V��.����mc��`bC�(�Z_�܌�IM߷����y�$��;�����\��I-/���Jz���w Sf�1�J׸�1a	n��������۵��#��.��{�E��L�A�ެ2W�QI�l` �U�����X�v�u��v��(2��}��6�e������bNɷ"��W�'��7n^����}<ǆ���&������Յ�S͑ʨ�
�ZI�-*Qi[(ۄs�q{�Rx���70�t���yTG�3���^�+)��y|��I*"�9��V4�����Y�� �A��JUs�O	-������l�B�5V6o��`�]�����LİZY��C�"7Z��B��^���C�����z�(+�\�JK58$�4G��F=Gjh��r���k��f�^�_sONQSԻ�J�vL�'l�,��o:3��i��G��en�$��$��Ϊ��A�e6%ڵkCL�k�سW��a�4�﯅�Fd0sRԂ%V:��v�%l>��[>�(�xBՑxg0Z��m:��=���%��v�3�}�ĩ���KcLw�ڍ��Z�O �	_r�n�$��l���~|��[l(�u�V&��j��)�s�U6(ԃt"�BUb�S�bNP�lP�Z��F+�����f���H� ��Yc��,-�ZoG��J<T�����wҵD�B�P�l.�h8�ÀyB���e��_����&��63�df{k52�9[OmhQ��h�}{~ƈ�]��
$ߐ�y�qS��T鞽�z��/��X�����������=k���Gҩ]�	�E4��ۛ�i�t���o{���Ŋ��X����{��_/5&'��f�d�����7����SK�Z�>��L�Y�K�-�t|����9�^^_�ӧOr�g�U���&|��;��:��M^^NV�ں"�3�'KZ9����k��;0��m|��07����T��!�r
�wmG�N��A�A$�!7\���6�T��uz5B���_��w��VE��D���߫��,4	zG7�f�m�y�MR,��/���`c��,4�"��4!ݍw�c'���^�ظ��^��8O@P��ٵw����*��
��4i8�<yoɮ�Ld�-y�zQ4H�#��
6����ؔD�\m}��3F1+� ��l�p�}�yie�H�bƯ%!����U�g�;A�0F�r��[T�z��K_�@!`��G�S��=����ˊ�� ��C�}�4�)Qyͅ�Ҭ>����_`���oz��ps(:���3yAͦ�8�<��ps�_�^ߡ��/��4���/���t��/Z�D�����ϛϹ2Y��oo�o~����}̴�� ��}���<��_�H�<�!0���������&��$���I�f�������_3��6�mC�Y��m�Mb����i�D�3�M��FToe�l��E���I����s#�Y9�P7��{��D�(vGi�ȉ��*�����JG뺵�0v�V�0��v��C�p�s���Z79D��(z����z��gĚ(��z���1�N -�W�O�s$R<:#2 ��������م�^EC`v`�X������y�<i�I2�i�饞��n�l�1����1�i^����,뿝]00�%R�l]�U�F� �m��I����l�0:�{�i�؜���u�UD5=;�b���2��.�f{E�k;}�kdE�����"[pX�I��LM+�y�@Ż�Eȃ&�O�C���0�@%	)��*{��ρN�^�I��4������\�3�7��g�̐��HCM{M�\���*�;3}��Պv[�]�#��[xK���dT��e�M���UyV��	���WL�f4��V*��Ԗ9�kê
�g�����F�����	�G�O"�d����팢�V,�Rm@03�_�"�e����
���^��'4d��58u�U[�4�Q�����ov>��(i�ʊ�C#镡Dy�3��6!�-D�n��|;/l�aO԰ ���{u��B��5���iϢ(ۃ�ִL�����r���CF���ߣH2��ެ��_TX�X�aBL�/vړ����o��L��q��,uq����)xΩ��cOa�4���8��煢�V�Τ�#����U���k��4�'G��d3#S�)�Đ����,��3�j�ى�������!3;���]M��s�n�b#�.s�E2ӈZ	/
H_w�w��	���N�
�҈�<���߃�ڒ�^�K��U�-�p��q��3Ckn�G�C��v5�T��)
V�!��X&lԉ�i�l�I�3�[��R����0A�}��3�3Z��Cڳ���C@}��M�1�Se�jDQ��0b�p�>v�7�-���T	�"W
r-!���4��O�� 
�(E�<,�p`���Nr���������L��a��ٜf�7�c������TU/�^h)��|;λ�x��6ҭ��?#��_Ɲ��-B�L}�V��j�
ڍXA��g�>쬎>x�oK�KCH�B8T;=�����n���hvE����q��JHƊPS5��~�	x���A��tH�i�\S�8�ܼ��嚵M�I2H�I�a�X ���@�(y�{7�W*�),�Sf�ؔHw����r;�0�)^�����,s5g2���c>ug�[T0J�4��q������F�^G���5o;�'�K]���3,s eH΋,�y<Ӝs4��������6[�N���OO���4����y@��P^!Tx䏵9��[�C�N��=�Ǿ��>8sU`�-�n���r��-z���l��|[0�:/��r�V��3�'��#�� o]L�3��T� �&h'R�Z��$Z�(�M�����J6�w*l}z�߫%��Ή��w���[=ې_I�P	�a�+㶷6��YP��LZА�{8=2A!��c��9+KL����͝R9�z��<��;��<�%�L�b_��Gٯ�(�[7�{$�M�060쩯���A��W�LFg���:�2vzn&?թ�#T�O�gl�&�s�D�(,,��ζ>�7���v��2���2��)�W5ѢP>��)�	���1���r|�JAN+��z��_Lêh�`���mP8�F�`�ҋ0�'�{�����w+��&85��5m��i�!��j�|?���+���	��֒���#���X�Y���5��8���=�k�iA��m���5j�YǓj�X�ǿ)�$�k��q��1g����(���m���j�ͷKm��/��Mj� .�P���R���q�(eu�Ӓ�ȀL���Cj�`�p1����]��TX�,�:S�$S���c�j�C�w�+�r�%oB�2�tQ+љ09y��G�B�5��B��5#��%\�~ؼ�L*?>���@�����
��j�F��=l|V.��g������M0ӭ��Sv�d���5�k[6�N�����i��B�%�����mM��Gj@r��{�e��c3��x�xo8S`�GѲ��S�	�\����X��O����,�=��z�מ��	) ���ڈO�]������"Q_v&](B�����2��o��VP�S��x�DT�o��>C�����o�gx��4㪳2�vc������	7Uo��e���P��0�8�M��	Ǟm5Vw���`5X�iZ�B��P��Q�U�pT�獵��1�w	�z�����=���'����i��I���(��߹Q4���7[x񝙽$1��f7A8BOD-R��u�xO�cF�u��$t�
�C
/��U���ڜ5��zcHoo��[��ǯ�����c7���P��6<�/%�5�R�&�L�ړ`,�<�Y7�j	��hc�0D}�}b���/�ݷ�#���QZ���D��L5��a����K�/6��6G��{}���;&�R���輡�Mi�RƐz��m[/�ւ>��i�8\�ſ�x������[�-%�H؍�{a�<gþS2EB7�M�~�r[�ͥ�� l���4Tx*�C�|dTGa7�T[�&��N��mj:���3V�6�{��&Ҝk{�@ja�(��߭��0Uf�D��C�1Kk06{��3e[6�M��iv"��S��EL�2�mX�:��i<��'���*�S�O���m[�P�0���L�Ż�l��Ce�۸h���9g����X;�;1�B��d�����:'Za*v�`'mY];��r�P�T�����5Uu�WiQ_L��i(6�Z��53�Ն<BS��0ܾ}K���+Ғ>�_t쟔aFFR�L �����k�rU ��g��~|.G2b0���p��SM���W��=�T3��p.�~�1Oz��,�.�t
�-�)�sꂖ����F��gI˰i�<�`n�p��za��s��(A�W�Af6Tk�tđ�$�bW�j���ͷ_������G��6�ʗ��"�(R���g0�r.������I�y����_H5v'�(�Z7Fe��D���X�$�#̇�=g���M�<���k��D�;���?"LƑ(TK=`��8��g�W�з�9w�����o[y�q�o=�J��7�jo���FǋJ�g$�󫲠�b#���h.d���&�gf��S�`��hP��%Z�Jt�t\<|��9����N�1g[ B�G�F��e���P\i��rU3T�s�&�;��˟�l�X���]�5����C.>F7AM�Ȩ3t��j�1�������I�銨ܟ�Q���؎f!��6W`�����A�v�i��F��Y��v�K��f��2I���#��RR+#�8�풽�/N�����o��/����o��j�H���C]�0��Sf��1����V��)<�(e�N��{�5�s�%_Z�gƆ�{��m��87ŞiXD,�M�y������k SS��Tbi�a��f���L�
s��}u[��	L5��BBQ�h�l��L9F�3��Q&�Gr�]	�3=lz�6#�_r�Z�?i9;L4@s&@"�l�HM�a��Ĕ�K5�6����尛 �s���eV���f�H�L]	%�����,�Xl�b�;-%�
�$�����n�C�"~���tfꜼ��/7���?�I�����_n?�T�I�e4���4	f���7	�|��zW�iZ�6���{�sjz���S?�4�Vm�5� k`���i6��H�L�,�DbQb��������*2�DnA4Z�K���T��M^N��Vr��ڢ�H/g7���ę�:���
�� @E���9
�����2�Tһ�>�IY���E��|m�y�*N6ôU.�L��Jl�@��?���ȕPR2Iu Fv��ӏ5 �� ��'a�kɀu��H�S���6�=*s��]#eѢm�2�C��� jz�����y�w:%��
[s��qW����ζ5���fF�*�{�)�d^��p��<�J̯3�f ��S7(l	� �[9�n�r���E�ts*9"D|���12�`�k�">t���ט0�=5KS�����p����s@�� 0�}c�z|܄ɷ)�h�|c�_���A�wۗ�M4��sP$PMr�駛'e�[����n?���>��`��s
|�� UU�Y�?�P/�a�t�&�%�^CUDq�l��z������E��?o4�'fD[�Z8�F���|�0@�VL��Qh�����|��k.�)BJ���x`c�6)��Cc�om�`0ր�6pGf�VjV�Q��:l�S��цei�T��oB/bB�NhL�����;)�PKXpV֦%} �����u?�����F	=v�&��b��W)~�S�������m|Pm��2ȼ!�ZJa趒Z��t����R��p>LIn�F�݈����Yk�Ջߩ��j]@�z@ڂ�B��S8i����<"V�Q�٫�j�.�h�fe�+LM9}����f�WE���eH��އ'�d��tA��Dߛ�|�rB#ە�jv�2y���wg�a����E��gON=��(�X�������h_�����y����'���~.��`{�)0�36��2cp�HZS �^֙�~�cR4����禮�}-�����_1�U���1�?.6'���B�p
mɨq_f�u���-Y� �B���3;����,�:ԥF�J"΢} �x�1�J�s����s�
��/�?�g���o+���Q9�p����8Y�����-�3{uKsBn=l�`�ծ�����H�(���c���̠ab᳾[e*��@�Y\C��d���wW����bw�X�*��ZD�����֓�~�kG�F	����k0�1:E�~I���y��::�XQg��ժyЀԇ����a�p��^��~~���l��R~b�tC����
d�f�-��.��u�I]P�0�d�M���
�iբC���5�U���.�����s9�����*�RҌ��YW`Ǆ�Y-�0�8�u�0��w�
��S����9�3�D��;���  ��IDATr��l3�@m��'��N�q��57<�5ig�+���;�DX$KCz�B��x��F�|�?�|G����s{���TO�P
�{0��80.����B�f�M2/y���]9��"h:kg-!n2�`�-R�cwh!�.u퐺Z������z�o��җ�����Z�۞7��A.�ORV}3,�3�k� R�}�_s2U`<��.s���5й�$3%��`w�3U	���w�!�����ΰr���#-�S=<�΃#��1����=�_��6.a�)R6�Pw�;��0�CG�@���5�VB�l�D'Q66��
�$��9��$Ђc�9���b�F~��F�lyF��1�\��2�����%4>�_���`a!�6p1R>*ԩM�I���t�}��A�	< )�:1�ޛ_9�$Q>։��:;��3�i5�LY<zx�������a���2�-jJ`�N/^e��zx_��r���D)xA䌎ÊI�)��%����KE���ό%��P���Z�z����5��������ҙ���s�8��T�ڭ �8��b�j�9��sǑa��r���� B6D9N�3�U/G��vg"���"Ҳ���vH!H�3'#ז���#$!���-��f��������&:"�ڜ̐,�!B��>��{X�2�;{�9-�!�:��f��;4H�� [��M��B�[��q��}��u}R�|�@h��;,L�A��[��Ѻ,�Y�3`��"�;����ٛaH3M0hr��yFM��@�x�?�h��<��zO/t4�]MOm�њ�*���Z��6�J�	���	�:cN��%����~���;V+�@y]�&��b��c�P�O5��P!�8��c��d@�2�K���;<Ȩp���.�p�B*�}\����]R���I�ʄ���6n���b�8�g�[n�����,L�̔e���T��8��`�/[,f�]}D��YG�߁�b�
�T�i�]{h�PY���U�f����r�Cd$Sda�G��&6����.�67�XW����'8�I �%��l���M^`�c�`��e:�)��I��{Tݵe};�-��L�h�`>p�P��6�oJvG�v�"���) �f�:�b��:�lC�2�@'�C�|�!d?���lA����["0έF����j����\9)[W�B�ИDE�=T'sqĢ��8j)7�<��	�$�;򖺮����g��	g��9	fӋ��a'>��[�{��~D#w��6C��-T��qSZh��K��ؘ>7�m��Y��#�����X%�1��(4�3&�<ۣ�HYf+l�Y�aᕠ%����մ���	�Ff��;3�w�hf�Nkez*!̕�<g~H��T����^md!�|7e|ӝ�Kdh|wF
Ĺثc�\�����s8�f+.�.p��wYZJ��򈐰k�%fX�J�:��6҄p򠅃��_�H5�$��U3V��R��
y*R�Ҥ��_vGlK�"])��]	aGp�1gyfc��ha�a!�;`�=3�8�o!�djQQ������)%R謌�������`��^�BM�l0�`�>w�3���m������5v������d�/3�c��FMv��L�u��Y	!�-��e�T����X�v��ח5������Mp!A6���lŗݚS���~E�~����c��s�k�0�=e�Ul
�=��}��b5.4�c'(���F%��^M�V�3n���#[P�m�ݘ*��Q��2ir�����y��y@M�*�"f^F�22,��-��Õ�6��]26QB�>�g읅�T�j��Hp�#���
�f��vP�dl��gs�`si�:̎<%��� �H�.��� �&f�U��xOܢ�Ƹ��� 칹	c ��ܕ��	��cA�0��%�Kk���oe��jn����� K����L4�����@}������J�W�t'�7Ӄn"��J�wD�s�?���
�+9�:�nDӘ��+�"H(J�E�%P̹��@�jK�1���C�v.���.�`ȡ������[q7W+�"��j����1B]�B��ݰc4á����4�m��D������=xh�,��#K��8���od?����������ן�r#3B^�
LT��y�wN)�F�QS`��)U�w�\�G� �s��N:�����e[��Cu;-*+C���sr�]SeQ��5�e����gG-���O��l�1� bZ|o���0	a�^�z/d#���Z>�u�#{,��3����ujRskH��Sؕ@b(r�1�����.=��Gh8�L$i�j��-�V�3ή���f��%�F+��%v�
�Qr�p���@��(�}m7��B��o�U���y^���U��sHK�eBK_N��t	E�0^�·Q���jˁ���\6)�w���ply���]�y�//�m�(�6g�2!�y�yZ`v/�#�������N)���71����̭(��B"[ե��lf�\גQI�Ǿ1����/d���U5m�����cʕ�qsN�:r4b�ք��afվ}��[`3!�YL��]���Ȓ܀��	�?L������&r����;�p(�9� ��Sr�X��=�K����ƒ�GV������Z{��h�cxф{��ZOt���d�]�Qe���,p��ʠ.�)����G4����P4� �� �Ϙ%`���h���ט�>�>��t�
�ޡ�`��)�F�\�I��d:+��E��(��y( /M(TR�qd�r�	��2� �i%s%SQM(��ExX�/���	fR�f�Z���Һ�Jƃ���}�nP���`����=&cQ�$72#-�w�)���Pl�"c��������B+�H�J[he�(�9	��%�}�a�k�<�UVgJX3���zh�����ѽI]w:�90TC�}�Z�����j��َ4�NSn#�*fG�����R[�~Z&I��@{ �f�M�L)I�Vrg \hQ�i$����Ʊt�X�?�a�zT���ɀ-쨺o5K�i������ŵ2h��������g/���$O9<2<?aG�`�x�rg{��3��;K��(�W�$QL�@�m�h�����Ьj�T!�(��jʜF7h��Qu�}��7;�I�*5�(��m��ܛ�sCyB�T�!���c��Ĉ�Pk�&T(����"�(;�2rrf��q�U�9��6���%[*r�{X�K@�k�̠�d�LkW�����[K"� �C;n�/�է�CȎH=�I�K����허��`�L�18^YP[t��=�[��#p���1��
[���mbX�H  @����H��~�o9#a����jo��~��k%>���[�g�����T�:�%|+BH{��ԺS�Hަ��(��g; �G�
��c<0������t�Uk5�*��	����V��8����`�R��̈́qe'Ȭҙ�&���+�M�&�Dj�@UsD���v�=e���5*/%g�-T9p���Y��D�dڐD�3|�QMH�ՃF����m���Dq����pAN$�4�<����F�D�I_#��bg�v��^׊��QH������1�H�����^�l�B��w�����`�B����D��-�0�(��b�H���-ь�k1���,L��Q��T�hu~EU�����b,2+17YE��h�.SJ'�Ҡ5�-��G�xj����r�O���Xb�ff��*d���YդLɃgI�#r��9�V��
�ԯ?'��.�'쯤jQ�cUw*X:i�X���s��м�'ߣIV��?W
�����!Z�J���)�_�g� 3d^#u���%S���408����95KN81�d�ް�{����0^3� �l���;�NŃ<L�1i�ֻ5_ p\;�^������&����4��j,<4��Gj���T�֑ tc��^����X���i�:�-����kV��,�K��6��1���G�(�j�#t���`o�3u��s�L*G� P�f��'�R����d�~ �D� )]��	�R�u��ѧ'G�DA��<����I4P��݈�����X�Љ�bZ}��IK@Ay@#0�=��N�&� &
�DFt��A�K�ʕ�1�et,G)D8��erՂ�#���ω���PQ�6����q�)�7�ݮ�ӊJ����s"��9�-��cF�xv�?R����6䶎%=�1��z�'�P�;q��FEķNz;��sGy�SÊ�W!'e�'�8l��52���lR�zE�e��������J�č�l�N�ړ�����ik]��L��}��B�*��
�W�2 ��S�'ơ΢9����L��;#�E��f2ҖP���LF�y�|�z|��4RR���m�?ҖiDH� U���\��ѱ�eF�JZ.�8�2��瓘i��9�lF�z���qx]�)�(�Z��!	'X2B��]3}lx_��e���@��3^��a�d	�,ox��L��:	%��q�֭߅T�i �f���B�`�+ݝ�G�9l|ي��1�It���b�Z�T"���g�{sr�5�A*aв����F�}+��u����O�s� ��=��(^�xо�0u[z�(��J	]L�ǜ{��k2U"���İ)Y�����o�*��v�=?�j$���8x#OY!�5�*�ã�O�a]0���q����Y�l0�h�z\�¨�:��c����G}1TV�	蕀.��Uy̎YS#���8�̀�)�F���5��)4��Ǽ��9~%�(gD�ȠeǺrP=r�=����L1��sedh��Lԙ��a�<g�Q�z-;
����'B�`�s�\n"�l�4s2�N[֖]�]�^�-�<��+Ѝ��v�&��e�ˬ$i)�Q!��0�E���@�n�W/Z}�Qb�6h�ދ��5;j84mZ��em�3v�ș~����(�A��� *eV�I�O1z�{s77�{��G�bc�P���s$�1I�A����bV����ۦ�;Ɍ���,79�1��s%pOT��S�ww�66h(��Os��|~?�X����-ո-��hMJ��^gć����;�o�^�XR���r�Ek?-�� -6�;>��`F*"�Z���Xx2����&�+&a@>�}T]۵�sI4Θ_U Y���|������+ex�߃h��zB�j�T�eV�Bd��0�)�ܕ4���z�1�!�>���Ԟ@�����������zV�I��!�1���2	���1�ѵ���@����}���L����nӖ�J�o�
��br6�IU�/��F�����Xh@gL��C_����D�(��K&$�>l*l�L����T�gc�H��5-o�*?�Ę-�[J�+�B�gm��awAJ+��J
�Z7�8#,���n�I�*�Ph�}�#*�0G��N�'�h"�r��O-�z�#�;�T�4#�Zi!M��Fg���=� �U�� �ۼ��=�z��8���r���XLQ��u�|ִ�UCʽ���SS�'�+�`K�i��R
O����;V��.eG���0U��,@d�1�c��`koO��H��
"ܼ�s�'v=-Dz�\�l���:��W()��zŋ�ֆ|[H�G���PjyKZ{<i�r�hG�{���t$�� ج����K���.�"m�_� �Ň<K�e8�O�<Nz�[�{	�n əaD�4�e�{j� {�=$�_��� ҄� I�q�9���"��������iQ�'!f:�a�����-��(,Q�L,xQ�:��I�Ë\t�3C������F
ft�B�);3�`x�M��@bf��F��p<�"����aګ�z��\��6Μ���_��]�
S'�o�iZ�r�.�[��<�	�ט?󙠋%�7�뢮2O��fWJ~G}B= ����AՂ�����M����a�aN�oKą��e)u�o�����;ў������V?j�{m�]r������3�t�I�T9��������UU��Ȁ��6V�(�%QCi`a[ۑ%�Hx]��嬜ڔ�f0����a����c�ґ�YB8,6�D��d��H�ſ������˘�2�Vy���9����*AEɎy.f'-��-��`ʸӬx�Ș�,�B�bF��Ϙ���f�^�"�T�x�V)��*���Z�%��*y"���F
�L��䈙�Hb���C� �2Ė\�&�=��aK�佣���?���'B-����x�`I�=�ϑͤ��;�l���G����w=��������L��3k|�TU����y�|���5{
^�vM(�+2M����f�M���@&��-���;bky=F�%ڕVhЇ^齹~�Cg�`K�X)D�B�CHI�V�6-���Kdui��&Q�#���q��f���Ɨ㨮�l�ߗ�+zX
�@(S���,��ֲ�ƒ:S�t�l�A�;Xh5���C���C���W��ڍ6��Ҩ$du����[ݙ�f�B	+h�l�`�#�V�E�		��PB����-�7��l�iHJg@����~��UFbV��7�Q�I(߱p
q�ݴ�f�
5ģ�~�M�N@?���e-}��E^_�2�{����-x�N��2gb�=��B�zeb�~��G�#� U�ɲ�ߩ^<������Vu+�{�T!D	��?l��Vɽ8�����F��0�5��}��e�~�6��a`�y���[z�3w�*xN͢
�1a׍2�H?F�S3�w׬jU�1?���R�]�} ��1�����h�]��F��L`!��+j'�LHܜ57$��}g�0ټRZ���u/H"6g#й���������%�,kج`;���QK'=�A/Z�ǽ��R���F�%��c�6���H�m��. ��qڪ���Յ%�zΖ�{C��-ҼkO$o�9nYt�E��e��N�s᳧����#s����f��ǜ�Z��"�6y�j�-coh�Ã�g;٢M�J��(��rc��������O�׿����"�������&�����R��lW�x�$Ę�64�Z�Pa��PeK*��2\��ϑS�ꦤ�b�`�U7����P�0c��a�c�|b�e?���g2�Iւ �왁u�I*����~��':�33@��q�v�wF�u�γƼ�l�F�T������V�������t�X&��:���s���{�T�h��ɰ��ryex�&�g�ڄy��f#��B�7��Q�&����˩���V9״��p���CC�8YB��n���ݛ��5՚�����1>��r@{�`��jS�~� we�z��i��D���b�/o麻���A]�^Ob��^QŮ�2�`�I�j��g|��}+� �|���?F�QI= �>+ݹ��J-2��T-�3~h\��ss��!�s�s������ÊR[�Sx�o����j��`O��v_�뇿��I���/�r�����������l_sR}I���%�Dɵ��~�xμ�%1�a[T���q�-tH�:��og�WG�R-�bBV��+?�X��ɾI��:;>Α�_]mw&P���)�z7��|�����xF8�H5#,6������6�Ѭ}��|=o�Q��lE���\��.��C�$���̃#���G;
���wG��M@�w�.�q�����`/#���A�2�E�Y�L�eӄ@���6z���wS��{+L�8ɟ���L��Ͼ:B�� "3�?ф��ތ1�J�kv�S�s��7k	�����0L^�A��9킩���3t���|t��+Ԣ��ti���#0F��׾��%J%ު����ߺ�/�iW�>Qj��}�\�&����{����kŭKz���Ǔ2�fN�]s�ؘ @��yф�Ƶ���P��n�d���g����b�6���R��2�.����y�T)Wv�
MB��2�z���=Yb�j�,��;Q�X��� {�_Y'6�ΝW�r�(��̮�P�%:Uޮ��QVlct$��	��CVk�*�f[U��xC�����PO~�}������^�={�o�a�s�mm[y�˦�m�m��Q�OY����`ӂ���d!��Bbm=� ч$Cu��b��|����Mϻ\^�ǳp�jr:8���6Yvjj\�Ր���XO_�-i� �
�t�i�V$�ҜeV�15�;S����Aޣ*��$�{�Jl�; ��;ã`�Ɍ�F{I�l�: G�<��p(� ��cߏ��oN��%���j�9C�z�gOrJôA�u˙���dSS0�/�5R�t�t�������S�D!�����XN����\$ ��\╊Q��RH�F�eʪBP���q�*H�}].��Ԑu���eQ����b��!Uc����k��jHZ�:{�?�n5���_�8��K}C�q��ض�*�]J��ʣ�i�8�4�d�������Po�Cf��q�����\s�o���x_bf��JsY+�q&Qg2#�Z�r�ԧ��Z�hqp#�C�Ȕ��蘰f6ψ��%(��@躮�XKx�\VdG���Xr *M�>�Ⱦbe%��A��o�ccG-#p����u�����&�1�~��}-�ǳ���rEHc����J�x�S�6� <ae�#�@�k�i��D��:	/���,�+��hq��:�<����}���S��)X��F���aCɬjA\�GDh�7C�^��1���-|,��P���	�f�͋�|���!x��VO�y)BUY�~������%Լ/�µ�=�2�;`~ "��mANa��0����3Ҹ�('5tb��y�)��������x�9x��oĳ�Y�U
�s|o��l���A�`�(�c4����)�w�5���G_6�j�Rh�Ҡ�%i�
Ҙ@�X\ˉ�<����A��N$bWǎ��p~�		NW彃9��Xl33X�D�s��n� 8�Tg���=�5��<gYh�_��S ��x^`?-`��ZdBx��>�Sr���fz^]%���Ү�^��� ψ�Azά�BN�B���
���wW�Y�۽�5�E��.��������\��qԧ�p��|:%�(jP�@U3�v��M����[t/��$���mp�z�lF.suK��H:�	qL��
��C�#��#m��&��s��P#C��87VHQ��+TdV��.�v���s��;�v��r�Z�9�t����v
��W�68Ɩ�"��!H��0�T�����Z�SM˜�ӧ�3�շW8��е�̏���TO�����iN�V���;���$�]�xdC	��)�XȚPo�t�I����[h�lr������~]�=@V5�H@�:W��s �B�r�$���&���m�����ǹ*ĭy������7ԧ�)�D��I��v��0b���~c ר֎���B��1�^j��W��v�3Tr?�3�sy�>��9�(J�A��g��l�zkU�(C�"QWR2�-�o��f����������l��Q�_�}�<j��U�@�L��Jǐ�҈y� ���/���U.t*ر㎦�����sn粙 V�גr�FvWk��aP��h�(wH5mx=KNц�B$��vur��S�+����dT���R��� 
t�uRL!��^����_?]Q+���k�ֻ���`�ޡ�B����w3�x͌%	 �T��G�`��S��Eӌ�5��(�d1㛵G���m\Ɯ[�������4a�'O-0=���'���STw[�=�+�"�T�{/�_o���&ѿ�.����:�eš����6x>���vZjeذ���03=��9�B~Z�4��*9�1P������J1cQ��V'�������j7�b�a�s���1���Dt���	@�ʄ�P9�a�iK�Su5�4��W7E8�TO�X�����_=�Ω;a�1�f���{�Tb"�0���ֽ˥.λg�8��,�U{cd���g�| �2�&؍Q�Log�h���a.lNj��Pe�_.�S �TW�v�N����X 4 �OO������/�g!���f�)訜����.�}����C����<4�L���g m=� j��>��-�p9�<�Ϫn��i���ۃ	�g-�NM��rc�/b�H�}�ta���V��aX��vc*���M��T���oa����MU�c��V��Ve�[�Cf���y,޴X5�1��m|@|K7�h5&UvZ���{�����c�����n���r��.��4Y��u���r��-��bv��s?�=�;�\C��%�Ԃ2;���M�}1eؖ�Y�c�pG��Y�X�[�c�����b{_6p;�mh7H)�zFE].3AiKP�m.Ȅ���-��Bbp��E�3��Ȱ��k�Ac^>�<,nӆ�7���d�S�y�߄�u��	�ZڍC��F�8�<�KSg3����YVRUв@9j�:hra%S� S�T���z{�n``�*��&� ����4�Z�MI���!�!T�@�>�ΰs��RÀ>L*{<�nD���b�jۘBL�K��"9[�Kr5��+\���s��g���`;��3�S��p�Սi�W9�_ѦH�B-�����6v�^��d
���G{ثA<p`c-�b�x�&d�z2FU$��2=ӄ��(q�M�t3�.fȎ$}���vm�3)u�v�Kh��q]�t~��I�'�F�@�_��Qf��vИ���e?g��I�#��!�̴r�C�Bp��Q{?�!��$*�{F��{`s�d�+��l*)���ZF�	����A�1���)�о�+7�TaJ��Y~�:�:�Q�*0pV_�{��3�'V�����i���E7m��������[��rMd���H���'��Ӧ��=C����Lc��PU��О=ԯ�����U��1��tAe�YTD(�@jc�{(C���	���db{H^SK�>��/�򓈲E�X�һ^#��4ML]!D<�U�!L�*�%p�mے���6�&3B ����f�YMf�á�͕e���>�bzڱݡV��fatD�P��Ib���t�j�c�!Ԯ��l��=b��KA&�@���;�[��%
չ3 	!7��x��U@�_�NQ�m�+:C��	�˞_2��o1�1������_����{&���J
d<3u�>0�9ɐ����sHa;��<�fC5��#ưU��ܔ�U�FS�ͻ�)n ^uF�=�~�*�>}�K�xX$��
U���3��m����*�5-s�>"�deo��Y�۵j۴X?犀n�yli�
ݳp��^�%;m��c0�1C��x��$@��B�'��Y��SѮ;�Z�%�<c+�%�-N$�.xw�8�KĂ�)9|��k��0f�zrRH�%zw��Q�^sh4` +K����oI��/��f"Z2�M5bl�s/����� �P,$����B�~a�D=���D�P���npzҹ���s0]~P��瞪�)��έ%#��)�*�av����=��]��s�4m�*�� -�6����xK�m��(8�fh(0���A��Y��R�����rc?�[�������_b�ZnvS]�J��9��������zH�(E_#Ii[6,lb���Ü֓*z���%��|�9z/E|�p�z5;���jɣ�86.��*���qd�
�odS	u��3�\��6�(�G֔\�|��m96����3<Ƀ���<���f�A7V��4�L>9����ʩ�	Ɔ����'�@�1�
(uA��I/3�Ia�hPt}��fS�( �5��B�M�"�|u�9���0-��s�b#�`��y�����8���萴&C}��u�v6˼C@h��v1T~c��P�R2����<�l���.ծ pV�W���ݬP�6+�X�l���ﭴ
�α�{&{.�}^��۸^N�:x'h]hm7���~�I�O�d�#�z�}w2i��v������ʧM��^q�|FR��c�����Z�X}� �c�����n�Z �wc�w�7�����B8x�,[�U�>RE[�4>����Qm��K�*�Ɉ�e�פPQ���8]>���Z�L(1J�s	��\��u����;4�6TMd�*ԩ�.�j��lf,r��}�y����^��m��3(�t��6�A�����Q�s�@Fv�1�y8R]>����T�1��'3_ܔ>X0�
7kɉ��ywεU5��&�m�!"&�dsgYq1ޗh7a�1�J���ʞ8���Vf%�&��������~�.�o�{\(yش��e��l�HPX�#�S�h۵Ǒ!l"%�8d�Y��
L�$��1R���>�^�x�|���b��[������������m�E6F�0/����V�u����YE�B�붴����<;��-j�*r�}�p�����ZK4e���n�7��d�L)��.���+U
��*ӹɸ��Vrs�9��{�H2��cǋ u2d��,���k�� �IA�E��TZ�#f�d97�={
�0Ex�����͛,�f�>���p��b���z9�Vz�脣P��(��Xh�v�x\:����?mT�c~Q�ϲ��p�kZD����4kiZ�@����-�ԏ�V5`�����gOsJ�;(O��/�?�6�{fI9W	��]���v*���]oj�6����8�bd&�6-�����������rcb�ʋ�\j�i�I�$�Enq��^�C��0��	{1����M��*�~�.�?��@����D�@l�D����֝䎂Q*�8����������Ϊ��H1�Sڔ���#�s4V�wBsp0�q�	J�akY�ž􋬵먧�L��#�զ�uj���[
�$��/HJ��⾡C5��ݎ�#�� ��BoD� �Ղä`�����#9��Vx.L+��y����W�jfBH�Qг%M���kz[��q��K
��e��&�px��"1�O8���}�wA��-����!)���)M��q�\Z�s���TsuVM��d��&��9�*ZJ����� ��q�[~�z��TץA�7�۹ǉ�ܤo؄�l:y�:g��Xm���3��W�r����k����rC"g|���ɶ���M,5�d'��,ccܹ�I�J���"��?��ΟP�X-vM\�ʄ0�A�pTqv�W����L�oOr(�#�7��y<�.�.��0	!�%��{E�`�DUaUC�n��l�s�T���iqb�
ķu���+.[�ŗF��D�'Z���w٣��T��i��$��w��3*`BЎ��t��\/-�MЉx��nnib �O�x>��װ+c�����ѣI��K����E�(��:��6d�]ӣJNz�jxM���Ԟ�Z1�
\�V�d �/%���>�V1���E�c{�Q�#��0w�/��LO��q
o>�X8�]"����a�8���%J%�՚��Uz�ƥ���<������R�@93�����TBZ(Ũ`�T{ْ�.�07/ �b�L�`�PF(��&M����L8�I*o=�փ�z_�v���sO��>�A��e��A�=6S�ˮB5�|r�d�V�!4!��4�*����%�o��ڒ|Y�Ghf(����f��6�n��I��6ԝ���0�}�q��r���$�����¦��2�����Eo��	�p��HA�/����g�},-�ix�3i�0�\�g���b��b3�:��%K,$�mj]�V��L�,�s��=z�g��D�t�y���>%b�E�!@̄r�l��s�<|���gڔ��C(�\w�ѯ_�S�s�!*K�>0��{�ƅV�fWьq'Cd���njo�)Nzfن��8�ZT8M�J0v��0��=��N�b���ky"�P����ƶڻ��,�Z\+S�7�:%�K�q�f0��7팡��h�6��q[{h�'Z�x�&~�w���{���L���D{@��� <q����ٍ�?ec���@CGԴ=�m8*jC��c|w���ǿ�P�������O!-�:��o�*$3t���&y��o�������D� �{nv S��l�'T��k��|/L�B��7s�z,E=Z�	�;G�Α�	
4wKI;��##Z<�4[�$f��|�����ג��a��)�P�ܭ=ƞaF����9��zCh�`�(�2@/��C�{���c���T�Z��#j4�J�p�M.�~~@ �f��L�:zF[fq��!F���D�n���z�*`�traЭ2ّ~1c��n[��Ϥ/жx,�%����D�V�U�r}�kj��UX�W�M���.mt�}]�L� ������GtW�ydf泏'"�N%g('S�o��&c,W��[�XS'͑Wf������ݠ�	�"T��*?��Tl��\�ʉ��e i��ˊ:=�ef�2+	�BJ�M�4"�g�0&SCR�)�i�Be�w!'�M��D�T#�'�lR�ہ�Vj_�hI����c��.����o_Ƒ�/­�;��!�9�`�q2�3���v�v<W����x[[穑1�0߁@�ڄ۽����ƚk�K� �Ƒ��8����ct�b:���6���&�Y����#XMP���C�MM-h��ϣ���`v�[7�w8%�@��}��5��Q��2��r#���eQ��&�����|&��Z��S�ߠ�svޜwk5b}��$�J�^�Iy��k�>��eor�+�L�SÉ�� �a�sV�@���]^O/7��dt:mKк�$���A�>�ڧ��Dᑮ�o�R{��B%{�����裸�`51�
�^0�6�Z�x�BB,�Pm���ϰ�'�3	�>����^�2'�v]<��h@��0A��.�0�S<��N�J�-!�2c�є����S�C�M�����%���n~N��vJ:ט<#�Ӻ-��*j��.L�~W,k,����\I)Nw�44�ƃ��F�ן��N6�|B�n�
 ,�R������l!R`����r�)-Ju����_I{�um�R�4��Uh�5��Wc�:X��?ds�7Oc�`��w{�/_>�_��Wc��?���}����3�ώ(���dFe�V6U�K ���zDB$���MՏlh�۟&��5���S9v��>���=�3l"H"d�I�b��&I�Mb+ƚG[~�y��ACh�1y���T��V-旑�5����9$/<�=$�ޙ����G��1�a�Y�|��ފ��m�٫�?�4�v<IA�-|�����o�.Lǁ�ؘ���5��6�����eO�|2i�Yo�1՞��N�h�j/�����P�4���l�,݉�*�]3��5W�!ñ5�`^�fE��1"��h�?LZj����`��MH�����9����.�U�	��N�ׯ_������o��K��M��g�x�~S��E�l�筧֙�
&�8�fÆ�{�f%��V���b#	*-A����*<C��=�&���d�$}����s&p@��k��t�FJ�*RڗZԎ�J BVw�s���A�(�����/rp��zK��f|`F̘E����.zd���mf�`��n;���}��]�T�X�,� ���f����dt��xl��]6�N�R�,��g�6�pr���-��K��0���W�2T��SU���S[4�0�{��o��;��Z�
a�qn����YǷ	����*�=�<�qKhH(`�sG��e��,3Vi%-du�׎�?�xC526�(;�Oʟ�|���bR��uJn����^���j�6ۓ�=��ç�9YϤ�ʯNU/�a]�����y�0�^:�Q��$DJR9��\L�ɞD��vs-��v�S �\D��6q2�Y��;jq{�ޭr�s�Sի���c�!�I՝噕 X��3����A"�pږ�R!m	�
�Ea��4Q��_���Nh����A�X����`\�(�c�V!`�{x���������6�hO!�A�`Vq������xA�~~+FL�0��N�̈b;����$�-��5�^N�6W����e���c<��� =j�A���n��jw�#��K�-���=�[C+rMo�g8�,��Ѕ� P���'���C:z�񴮧3�K}s��P�/J#��t��t6O��ɻ9K^n3u���.��ʷ�{�+a��~��ח �Ѫ��(c�t�,H��c3�����6"!��H4�y�^�����*ŘPJ�blD�gb*X^;g�G,6�*�=y+�?݆��Y4�qڌ�D�Y�(�0#Pm&2�#���
��*����'Q�1���A��;�H��/�/֑ޅ�v]�tDɊH�b'�MA�z���a���9�IC��k��s�?͢9��R �
�$W�ې�(&^ڂ�nhk!hB��
 ���ɵ1�� z��LD�W��g8t=j�`��y��4q��(^y�s�i�*�n�y�t��j@�]k��}��=G�`���_��̄���_���X��y*b���̟����E�Ү�����[����P6M7��Xp��o7)�.V$EQ��6��/��;i��3
�4R��I��q�)"e82I�j������n�mA��F�ql�"TI�b_�����Bh����N���FfDa�ޣ�����E(�?C�)
�p�G�;QV�����=2rz�:S�*��m��Lʖ,���^��HF��ϲ���Ÿ�wH����X�9*�!�@o����I��J�-8j�#�@	�*�m�ns0��	�z]�iT�5�,��B�84.V�"<��Τ#���q�PG̱;�|"N�f�\k4�έ4�V�Q�(�,y�-�'�
��)v�E�%2jiD!�	a�ӱj����w/�t;O��_@�W����Oϫ�/���Ž�ׇ�@��v�W�h�*S�p�C�*In���_n��f��ʤ�y��m�n��8�nz`�5 WS;!�ň}`��y�n@��w�A.����a�nj"P+���s`d��-�����`#���	1,���l�T�?�/� ��w@�@�@b��ñ���lF�t�̾R����G�"��*�͌�_0 � �����t��;#�]��������@�{��V�]��*��F�y�"?��V�M�^�W���,aO��N��:�FGW�_�����2������Lj{~%�˙n����#yMԹ�EO�p��u�ۼD�X�uBG4G���6����8TV/����ۛw�Ժ�C껕�R8ne������]=9N�ʤ��P�n*B�`���'����q1#���;0�#3�q�aD�t�;^'���?�����ױ�@�"�os=nA}��~�N�Az�N9������k���
�����t��`?���i��}�d���]V��u�}�]���9�������oɬ��Y��yB,,~�j9�ܑ|�`Ӷ�Hj7�����Q��0W�92��P�=P&�}�uX�ބP�xw��o��!��0%�uJڱƂ�l�}��������f~�]B�}<-��%���B>� �U�iqZc��k�b�I��Y�ۏ3�k��K5�Í�&����/�F��ɔ�߸���M�ο�X$�x�ܰ��f2]�i�`��E�����9���Cf�Ϧ��G0J0�R�ټ!˳�lm@��y���屧�u�-,��4�L�ĄV�YϲwcL�8c�����%[�0����V�
�g8�u�ю��Hr�:���0:�4O�}=¼����lˍ��<+��>��x�E����>4��̬h��֞�-�G��p��S�-+���E����:���*��{�C�o�P?�B�ۍ,C����s�ַ(ͦ�e�t������c��B(�p���B�CHU�� @?˵"�p����x����=�S�%�z$���#���Ah�8� ���#�q�~to�g��.��+d3�]�s(1]'Q��z0+`)~�m��uS�����@�yA4��3��VF�
��0�r�Y��N���!i��d+�?�׼�%��!��)�T	�l�3=�����F��"P,8��?'�0�����:��7>�[�3�<�x��/E��R��-�b��]틭Z����u��q����ƪ�.V;U�E%���2Ģ��A��G(�Pdkɴ�x����#X�1ڊ��w��[؈`�����d
Ta�3#�[4+�(6�:�՞��]�s*�9�����	1�dic��r�C�6�-��$���9����#��K�k	xyL�����ga�a&$�4�D�j��4�g��V�9^ZEs葎�N5_K0SC�X;r�,:hXc�1���v���[�{��[��������xC�#	`Qbb�`�~�gu�-Q����fZ�V7$�����&#�ǂ��J�f���m�E};2;����������ʊ`q<�C�Z��Xyc��~�~�� �Ŗj�l��CF�LzA����]�W�f��bF����o����6x:��Ӌ�8�:3r^�a���y>2�ܼ�1��Q������q'ظ�̱$ Z������Av����B�$�=��Q!��L�"J�%�R��`�M����Wj7P�)Lo�9�s����D\U�+�F��߁fb6����A�5m���l��<�x*C�NJ���e�/��� �k��Ѱ��i@\Y����OH_�m���u@�G�d��2�g�6g���5!�)t_�{a��s�Җ�k�PwvC;�$[�G�{'���ɇ��JU������ILuf|��G�:����(��\����Ym�Z�����7�k�wPM9yd���lS�P�%߇�F���G��Q<�1���q��F���L!\�Y��_�(���[;�kFM�m�����%jO�j��rOt����_Y�W)��*IχM�Z������2T��A�T��E���Ơ�+fT��أ[��sTOW��P�:���o���B�#�=��Oz��<&�H4�����|�7^	~a�"9j��[�^�A����1���� �C"S�;Uf(�`	�pf��;�I��8w����=0] �����\�=%�4ց���Z{�~5+�]2hdL�U��<"y����9���w�1'�Ě/����x3���y�Ƙ�бO0g�EtNIg�q|�yW�z��c���ؾ�|�.-�f�L0q�b�8�
��b�#��;�(O>��Pk���@������'���f1��o��N?�ꔵ���x����xQ-�G�/D,t͑�.���kB�|O|wDw��4�2�.������T����31;9O0/"k&����`��Ӏ��9�J�x�3zVn���e�?��nd#���ֽ��4�Ŧ,�'��GJ�ǌ)�n�q��]�l�
Si^��53��>�%5�4#D3B�߲		��XX
�{Y���7�<I�345�._���u�;��FH9R��� ú6I�5:�{����`�ǵ|��\�J�tL���P�a!W��m����o'}R[�����Q�rC��k�^�����礣���k�X���7y�l�����c�G?z.�X>������Y��8	h�����9D�����z	S*;�z���c>�V?B-��������N���ȸ)�bT����G��Fs��̿�<'&�4�qެ�'�$h!�=jǲ��($�����%	AS���4�Qs8�֘7�Bљ\�(p�댽�eS��xwjQ���0����֏;{7�0��8G쥺�7A�MIC�����*�ќ�i�����ʈ���tЙTy\�O�9u�2c���;��ʱ��������ϙw��(����|:����!ʯÁ}��}�L�Xr��C��db6Iح��w�ϱ�\�>`��꽔sCH�3������>
�0��xE���.s��4+c��Z7�"��D�b`>_U�"��nxF}��FrO?����j2T��,�+��tODo�]aYYR
�F�t� �*g6�9؎�bb˂3�̰��Q�,"�Vh�Sc��X1o� YA��& `���3��W��h}���0�SSO�Ӗ��/�G��f�����*�\Ė����^�O����M���낼}��Ջ��.ݔ�K����[b�H�-��{iQh%7\��&][�Ϳ0���)f�`1!��0�'�H]%�g�ji����GS 490�c���I�[=�-��r��c,���_r1i�y1+qU�P�+z>3����fF�?֙�ޡ-���"���dz:
�@jo�sTV���*-�V�y�O�}���١յ�nk�6���G����Tf��&��ZJa�e!��a�$���Z��=�?E�	=.QuL�=�$ kݲgq��GfT8�Z`�|)j�/_�9ޒ�iD=��~
�TA?�n��x<�����jQ�L��^#�z�w��0u�2^��h{�{<��-l�����p>�5%?��%��F� ����=���Ẽb�D�w2:����q���m Hvp�րg���b��K:��d��� ɽ����Nt
4F�Ȃ%.��B�|��7͛�/�����Ѽ�G�q���x/��#E�L[���ڦ�Xe`*�����B�
�3�D������&�2$�-h���<��a�e��l$��0�i���
�У�iP�֭:V&������O��/�y�1�v<7l*(>5��i �ZF�<[�~6��p[�H{ǰ�FS�?�,�ڠ�	F��p�ad�j�MUs�Ck�w��J�X�
�����9�D��	�S���#��jc��a�V�!����0f~7�L�{p��3M���}��y�L���gX�����h���q`v�j�z��5ң��(���(�OR3{�d��8l="���	ƼtCC��Q�}xI/6u�s�c=��,Hԗ�4��tL=�Ǚ�a����^�����쨪�&��,�[T�������i�H���㩙R��؋L�6��PE�Q�rS�O7��!"��7���L+�XRE�h@�#����z�TE� 3e��bb�!&�,BY�]�e�B��w��o��L���V����R� ��XO�'fu����'�ȉm�@N���� �Z�q��|������\3��4�l�MB�nn��A~w�e#��L-^}�!28�~\��>!Gs.y\�v��I	�`<TM�����@�G�奔��I/��V�j���G��;���s0�J��e�!����u�`boHn�C���E�%�Zo����W����Y5�(ş´�Ê��K����X����lD�r��\�Y����61�:�PI����^��؟}��YH82N#�;0��j!3�f�l�19@f9M����p����&@(1��Ʋv<�sTap�[��;b|Y߀���P��9�4���Q���x_�25��=�o
�����q}�������ݽ��KMW|N��MUo�g!�يwm�[���؟�8�kZ��2������ {n�边1�S�Fq8fM��
 ǒ����3� �n*��z6ț׬�d�N����ސ�ke��z��6m�;�t@$�p�c��v�V�B��S�;�&�/��̔�U&�7W�������S��m\����� �9sSa�e��,�'TH̛�W#���L�Z~����լhGC�q@���=鞌RM]G��i�87��fj��<�u�E�ѻ�3H`�z�7Ơ���&�4��IQ<��Ԣ�9�]���9���֨����=��3Tܛ��.к,5�O���V� ��a���S;�L�	|&R���7̗~��|�*d)	MV"C�n�E����7m�$ǱAUs�Ȭ�s�WfegDvV�����/-�[]��nJ��x�#M=�,�.��0wӋ�� ��'Q9���z�/��~��1+���X��wl�f$�ʥo�>�	��d���2�EY����4����ֻ����-��"��_3�>J���Q.���$�����|�o]�2�E����Fj?��.�Σͅd��m��U���T�zO��K�%#(d��7T}�V�)3E4������E9�^X1P� ��lYϕ�s
Skn�����Z�
2�iv} �4�L�ԗw���_�f��O>����r2p9 >�A�^;)|Q�{<~-s�{'�q����i�@K�S�1����I�Z�gq׎���}G�L��[k5��Z���@` �qm[�13Cߍ 2�2�r �aiפ~�!)!����[������(��7�4��|��E3��c}����:>�
�Yq2���̀v����5������AN�;��'9	Y��������DJ�#4�P;���&��^��FP�1�V�F��Ms�V)�u��6����A��瞌Ż�]!�~O�w�@����F�$�ĪKJ�r[џ�~o|}x������j��\�:Q�l�=��Ou*�ڟ�wtD�dҺ������PG2X��0�0��
I�f2 �@m-լ��4h�����ێ5 $�*���Oq�Nm�1��Ll�'s9K�$T-��n;�lx�	�uxO��H�_(g�vi�s� � �V�V����0f�A���W�+ege��g<��N"6k[K�8kw�{�%�^�%��C��&��ڔ��	I[~�4)[�?�����2н|2���o5.!R��ֱ�c�_��n�����`q嗽�MQ�}�K?0c���%������� ����^WG=?=�����'�N��*ǵO�(�� L�Z��R:�����300h�#�,B���@E����}.��{�8f�u��7�֖�Ƴ�E �=\fފ�6��O��SF@̘�R���}��ڌq7a��'�[��uQ
h�S����oj��9��6�8���/X#�M���іvD4E���ܟ��"9��[lm��"B-��`��%�g��퉊�R۞�Q�\��=�)��RwUP_��ǧm�9F�G���c�Ɔ�QG���d���L~�֮.�����N�,'�n�DW5���0ѡ�)�V �{�;lS֬ G���<��]�dCN����VF8��-�֨�YN���0)Q�	h����vt�]K�]N�=#�˛�-�)0��)�W�� GL��w����D�ԶV�D�v[�e���L2�h���u`E��t��4�Q�^i����$�k����!-�K�3�'���߷��$	َ����n-��P��E6�O��<�L�8��Pp����#��n��5��J�� `��>�V9r�Z�h"6Նw�l�O�`:�k�����PUt��ņ�w����E���g�x����P��\7�e3��y�@m��| "�(�7��:؟&�
�h;��Ŧ~B�u�cnqO �1��`o<��](����6�m��C�o�ɪX�f�C�w4����KO�.̡γ�K���hp�����d� +|����SK��RP&�`��)O2�3�{J�]f��*�ʐd�C�@���"��`C��;���[��o�\+71�Y�s�)�k;z���V��~f��W��Ɲ`l� Þ�4jX
������PEr�O����\V���r�ɻ2�����EtA�F�;X�wX?�r�<���FZz����ouݲ���;J�
�1��ۍ��T�H���[��w��F`Nt�EQ��"���2�<)�����>.�a[��5בZٻ|l�bʭֺ��z1���XƠ77R#�x�*p�]0���
�xDֹrhj=8�b��O�3P�-�(!W�E�x�6�?�X����@��H�V�,`20���r��=Y����H �3���g�[��*�G����{I�)&C$��E�^K+
`�L{���Jd0�T�h�\p�c %�� ��oQ8��z&��!�~ޥA�7�ҭ��e����!O�����7���x1�*;� G�
���E����٦ܤ3�
 U��T&H8������Z��~��b�PL�/��ɦ��Ŧb ��YC�w�[�D����`��C& �%���C$�V�7<�XFp���-rN� �ȸUf*��{:�����-�^`ΰv��hL*�i�rU6�9�y����O��V޴e�`�,�ˁ�F��������q�նX��ʄ��>)<n�2���(B�q�@�%�h�� �>O� >����̲=�����&�)�&�v�C���*�p��u��K�� }��)�h�z�u��KZS�-A2�}+vkq���F�`yx�])��GyE�\�u歲Y�$����9��8^�W�y�H�ǫm�䶔������WTe=���F��t<؇ھ�7A���"��Q돓 B��N�z���ec�,�7�>J��ĳ�|&�D��4؍�n:���<��qO���Tl���w�b5> n��e�pzrh�i���2�m�u�p�o�0��G��"�P��4��=��QέWZ�������[b&Bmπ% �g�<=�zP�|�M*���M�1��0���ց���S�vMfo����KC�5�[��� �}Ꞃ��]0h��m~~d7+�k'��7Y?�d�Q�N�wf[�  ����RkU�5ν��0�:���Z����(�u�;������'��p�X���t�98��3�4�^/��d'd���p~/�/'��?)�ټ�^�%s�u쉠�/5wh�-Ι��;��	+���F	 N������ ��]��{�I+�3�ۿ���:�&��c�Zi�㘵��hp�����\3,��Z��I�Mv�\�	�$�}:Y�|����aWKٓ�M�-ӳ�v�]b@eG�1��\]���.��y|�DDƘ�g����+�N05<����;|�b�Gl�����f4'2�Xt��C]7����9��M��鎌P�*�?;�����ZI��X�M~���%�M;4.��,�o��ᬕAe���}fQ�Ҧ ��� 8�A�
���;��D3��9]��`����&v97�4����2�ao��$�yӷ��Y-MH|�A�e��^D��"��H�¬9AjL���v:��ky�e%��(�Hƴ�Uu��lyUz{N��n��SΊm��̴3[�db��������tM��z����W�~1mYb��d�ɀ�rPnx����g+����i�*qF��?��������]�z����.͇�w�ٲ��L�-�S��2T` Xِ3�w����e�;L"��� V� -;��)D��E���BG2�d�����&v����)4�X���v�9F�K��1��4��2[X������P:������w�3�΂٨��Z�N�" �EAL��2)B��	���8a`Q��ދ5��S���\UE��`���U�6~r�{j���k�*7`���`ڻ���US�кD���Cū�.����Yx����.`'���w����P�VT�DZ��q��p����_0 b�<�u�؊�1��f�]V�A�Rm}-�x1�͉0�$�/��WK���z2���t��ܒ��g0����m����k� P�g��/�a@��l��
z^g?h�����j�1��*A�v��0�򚼾M�����#�!�(� #�a��%���*7����>]"'�IfS�.��1�Ysf���T�q�w})�s*Ѩ�M�"R���'�30���',𴰠��l�+@��?혌��v(��p7/������] �k��FoM�Y�>t��G��ܯmk2LҌ|����>t�$v[BR���:�=eֱ����Ɉ�o�3�w�l��v. ��b��q�M;��6T�4��;���� F�u���lW�I	�`M���^{	 �׎�O3'(m�����"�i�KXY��d���	Р��]N1�}޷4*��Mr��U�3����CF�����Y�	cN\�/�o�jQ�Q)��<c�Jj�ű8o0���'�=?������?1!��<}�%�N�u���m�����y����_�������7;��; Nq��`� �b�.�|C �j��!e&O�X$3-h���>Y�ȇ[K�53�;v���& K������f���ğ&t�l�V��=� ��X���D]�=��\����B��}���QC��2b2��X	�rZ���O`�:�(p����.�⩏����\�Ʒ�bL9X-���.r̊tʭ��O�!8����h�1� ���fb��M.�3�%��ju���O�q�f�.[.$l�.9{�{ #G��÷E���O{�����r����Z��1���ƌ٦ZQal1�flF�@j$��!���`����X\i�ü���ϗ��@�@m�Yv7�갆�轶�]Kϭ���Q�l0��j���J�I�����*��i� [A�9��^�2��2K�@�&�F]|Y)�&e�g��zD���O�9Uq��{1_3=W\)�1Pb�k�۳BΊ���3�����u��I��#�qY3(�ƨ1�ST��q��K���[(�d���UuC�r^��Qɢ��!x���e�O[xq��c ���ɻ�@��oU��j�w�������o�1��^�������@i-3&Z|�zTCJ��r��E;��H`٠�z�C]���l��9U���2�uǢd�O`�� t��x�	kzN8k�s���S��3r���i���z$c�2k�j�~%nEBqg�^~<��6��S�9�Q�6�"��޵���#㉹�0�� )�� cjGza���K��dF)�T�'L����xّ��s�=<�E���wV�-���YX�yi�ڲ��Nr7�-Zz�w2yz�@Yd,[� \�
��4d�B�������>_���
�����2�=�8�����p3����z�O7@�W �FPƪf�L������̥�H%g�`�� ��S��Ҽf���gґ�������d~.bb��`�cl TKge�2�i ��b�CdV��ic~6�J<#��
���0p#s[��?�\�a�H�/����X��%�����t��������Ƌ�և�¨��-�4�)�AZu_���@��J����ב�B0�(k	���h����t��6)��Kfl��Q6}��mTm�"�j��	��=���K��6�/����CC(�P��Q�gf����l�K���u':4Gd�ǀǡ�+{t���2�{���H���i�Rl�­��,��Ԏ��ކ$��O�z����/gv��P�^-���� �Nޑ�&�C˚��Q�x�� OA������--vG�z$��M9m+�������e[A��|�`ZM����M��^r��!�i�a���ؠ��p�Ȗ�^"W�wZ��ϲ���Q��]�=��bnۼ������u��^�J�(q�#�4��-��?ͺ��.`3_*a3�܅`m�T�B����[i,�c�fL8�k��s8ɸ�RtS=�9�64��۾l���a�Pͽ�W�rn<��]`t阱�h(h���_��_��zr?��k�?|�`����%߹�V��vmHc���̰��˝� 4�����g��L�B�>b?e7�,o@1;d�����`�о����?")�iO�������Y�3gw-tu��s����`��k����v����X��9�0b�k�&��waHZ�xͼ>cw+�z�
����R����Q߻��d[:��׼�A����Gkol�zry0Y���Q�BvF$4����ۈ��'e��0��k���k����=¯��6f8Y�ʤʌޯk�5��k�K�j��"ë]�+� <���Ɗ�=�xX�>�A��<�RG.�y@64	���}�{�0_�R�#ˍ`^�"W�O���9�ڗ]??�^~���|����|��1� �M}����~;�%�h���'�Vp1�D�4O���~'�?}�O7�_����Z�8��u���.����A�蕱�M�D3�ׄ�ff���lG������4uA�-ٔ�Z$Wix�5�c���)�Q�
oa���������a�)�@lqu	`�M���6<8��t����6��WD��з�m)�s��7���C���I�U(�'�m���������r��038�Y%F�z�r�F!OVOu�ȞTj��=1F�#/��	
	�m�Bж���K��J�\v�+Rl���Y����`�8^JD����3u�[n�V���
�{��r����Z��70�駟�_�/���Nf�;m�'	D 3Y����W+��S���u��Q�><��T�4���곏��fd��߈=f��B����qy�LL s�̀b�Ȯd�rL@���#������ut�Y��'��0L�'�������F�=�N�i+6���6�`��]�	�[��#32��H�����C��6�
�TQ�TD�k�L>OE��:R����^"��t��^m�u���!����2m�A�bJυi�	KL�Z�5��I�G��>����~�muln9j�JLeėh>�X���� ʓ�D|�@��M
e	��$��$c�zd�!V���dۏ��E�)�y���H+��r�en1yc���K�D��Տ?�(?������SǑZ:ۍ]�5c�0�A?L��{�,��uLɉ��~������Z_~���z��%�U�f�_<��эYKm8ͫ
�a�3o%�Sd�cM��7i�~���`��ɿ����X�T}����R�L�&k�$pp;�v��J�� ���u�9[�|�	ܟ �_�TRIրxКq%�Ef	��W)?�}�"���[3�]��\�YY�D􀸩8�/g�"�۷wA#����y����&�M�����E��y���00ԉ��t1D9�H� �zk��;����l�9h8@�Y �2�y�)�^��%���{�7�C�D�0������8o����T(6.Z���� (�u�-,����U)�*�� ���}��'>�x,CM�)s1�{7m��/y\z�j��?Z��(7`��9(O�p��ˋ�[�s16����X�#)�w�Tb�;�5�94�A[��4 5P$fQ�>U(��L���lD���{�k��
[!���ڰW��Lu�v�(s�A�%�޻|����=�MLJ[�O�D��Fɜ���Sk �������~)6������K�,g����ǹ�.�����L�l=��}`ma��ǧʻ�Գ�Ve*B�Ko5Q���R��vL@\*��.-X�Y<� <��u<�ˇ�:��}}Ѽ����H���s�{����_�"���nf��L�y����=��*���2�͟�U�L=xR�Çg��
�zaR
�NU��ٝ�,  俑�؉�=�� >�W��{|#ޕ3��~�΂Tۙv>�Qp��bFu�k]~�����Ͽ�kL8���8E�h�_C���f �R�a~�1��G]20��� �Fu=b�'�ۼJ�M@�&����I�`�2·z՜�G�0Σ}� ���o�ư�
�G*eg��&td�9B1`��5�!E2]K����G����
P��[�m'ś�d��-�7��!�}FiuW�߶��|@y#c�o�rM_#�M
32���ǋ'��v�P�j����s�b"��@=�-#���-�c���&�p^��[D��j�mQ�n${�	�n�o����?�Q���?��~�Ӎ��NfHf�͞�wy��.>T�$��6�D"�1���/	P#g�L�F��&�	��r�F��&��_���iY�(@dF�kƅ���[�yY1�d��0��	-���3�T��׿&y��G�m�#�p��[��=?�W�;����(W��Җ�,��1`�x�"}}Hл���V�+(1;�c����D�	��C3�Orc.�mL;.�k���>���K*ƙ� 4�e����͔��Tq_(�c��n������	�IBӊaAi�d+&�%,��}��po �n��D�����r��[={ж��`�0劾G�VZ�Yv��R�k����n7�e�"��ҥ�y��
�7V �
�����At�,��2����(}�+���x�Z�!�[鉝l㻣��nbW�5���L=�=N�����>%���,��s��fb�dZ��[�#���!��u�U��-}��Y.7!�=r��{��x���ۋ�X��0H�|��/dM��~:hC������0	1���9?�>^��ۜ4ʦ��P����.�$.���*��)���-���'V��?����>b��7���Bv�:	��A��> �q�~Ы:M�x���4cj�}�iԘH9b$�1��IW��t�^#d~��;�c��OX��{�T��8U8��l&7z~�2�@ 8U#X���[�3�"�%���� ��X0ѭ���}���-A���E)�:�ź����PaΤ9�NZ�D�M"��VB�{7Vb��n�x龥���1�þ�
ѩ	�|�	x��*���x۠�R�u&�gQ�ıZ&�Nˎ ^��;|GLU4��_b�g�%Z������_)��4� 0�@���R9Z@���Mq���ͱ�~O��No��� �T�aJ���p��l:��v%�]@�@EÃw'HB
��|�%���7��bl$�Lvo�����8 ��-��}ߣX��}�2��"��{�w�P����SNX~7�X?~���P�b�[�"MĘ���lQ�R���z��~z�~�}qM�0��^�V�ɂ���l5�<��s�#8~�SAh���X[�ϛ�d�*��t�������3�5�&"%���>`���M�� ��1��i�h��/������m!A��b�\ N��Ñb[0��N��l�J�[,�Y>���g�WZ�ä0�rv�����l6���`�L�r92�6A�C��V *�䃵ޞpH<����td#�9�_0zS\:)�O)���E�j�a �� F7')W;BݐTje'l�x�s�|)�P��dF_6�J&������i��\*�3X�a��)�������)�j��2�g[��-a�� -��o��W�Ev~V�bm�Cc����ꁥ2qw�ڿ>�]"�@�Ј�7�l���wa��&�������?=C}�H�%)" �'{
��l2�� z��塝\��%X�M�f�+�:�߉���u �Bbi������,��h˲�>r��ol9	#1���`گ1S�W&��,��ɟ�gmU�S�OF�0��E�{�G)3�i�����
nֵh+X��Oqk�5l_�L�rZ�@��/�J��R�p�J(�A���	��$�i�Ba6Y�A���3��L(^f5�:Vd�Ǭ@'��N�V�ma�(������� ��	�KȒ��_srJ�2�s�ٔy)�`���,��)Y=&�J�L�#�D�weވ����GY&��~Y�-rY`��0z�oO���G���<m3�ȝ�+����gy_t<P��߭W��Z4n�T8��S�2�hWQfLw?)h��=X0X$/��!��8γ���N>"W�������6�b��~T�7��H���l>T�~C�����o�Q�#�F+0�@�6��Jw-^Mv�A�z,��-�9`>{�k����P�b��bx�Э4�9h4@�XR���&�L&��ď\��Q��^�����q�5�T��>$4G=W�jZ��Ǝ�XI�ڴ �-�ϖ^ޔ�-�?��z��R�}>"w�.��e��T����֯�ڏ#5���9WI��Ji�rD�%�O-���3-?iL.AywX�=Z����j>��{Y#V�"i�+I��.�'��[�	� g-B��#՚&@�g� �=��/ C���vb��V�'�L#�>�2�`_Ua�m��o��l?n[��?������C�$�:�#�]�,E�i�&
�A�S�m���V0�\���8�>b�U^>J���� �ۓ%H22k�`6D�ꮥ��m $7$�˛AD҄�?vd��<� ��K�_u��
 O�3"���&�D��=����.�dܣ����X�>࿌o�߷dN
����m��h���X)
 m�=��1mh��Z�xt�G����-��8�����<��Y������ ��P�'5��}s��=�e�vT��Řn�;��C_�j��vuM���L���\��e�q�K$p�c�����rR�'���x�݀�2Q���򹹠�l�p�x�̱y�||��?J0ܩKZ\C��5SO��´��ڬi�W
kÄR�&|�L�2+�U əq�>L�"|y\��K���XP�n�Pf�__�z�[���~�Y]����?��#�����CM?+c�ml)mF����%���5�]�Of,�0�e�$׼{-�abD<]��wmg��4_F[^��x�0T����0�NN�%�O2N2������Ϥ#M߯�uŀ� �n�k�L�M�lP��b\lUˣ���YT롷?�,��o��[��n�:!��_>锸<}|����g{�^>^rr������[���K
��
��J4_��$!��S��aB���qX��{�xk�  ��6�, ���C.s%˷=�MԵ\�x$y2���� P}��?�:��������,�z@�i����OI�5����r�3���7�)��Pp�qWҬq�u�qhUfU�~���r�3De�b�.�Cs��LQӹ7f}���7�Kۻ2���P��Dx\*G�A�N�6�3���e��2*	x��d�,K;�p8;�tg䤤�O�(Hs0�b�c�l�ltd[�qD���"���duO99��_��l7�K(�`���]��BH�&��CN��q�p�7�y� ����e�w��C���b�C*��C��,�~Ǆ�*U�6�g�q0i�Д6��[���[����1F� ӿp� /c���O6�(*���N�Q�MD�%���v���P[�F�gs�0	h��1�>؜�h�Q��M�M��F����E�p)	ځ.p��i�����x�
�u�eD�0`LW*���ā��Z"v�8�ov��j0�+�)���ƭ��9�2f�	wd��W�����'�cw��xҎ��C��M����el^���P�seߊd
��Ou��%�(�swv�d"��}����e̴E��q����$*zN���
��^�7�W���L�)���� �J���
���	��I��MMFJ���x*=>[�g�;�)b\�pg��r���X���cxR����iqǠQB$�qj�1r��czy\�}��o4��.4m��O�4W���Z8�A�4�4�,1�l"�{�HYA,������N�����$����$5�DVҧd��^�	�fϋ�W)�)��Z�}�l���@ 0���}�
4{���>����F@���/��n��SB;>�ܐ��%��!`�(Y�ٲN�v�N�35�yS�u(]�U��z�/ٴ�~[��j	��
i��U�31z�4֖�i�\9�e�ZZ�T�@��)Ֆc������\�%#sw�N߅%�vAR��G�6Ř�?�
S�P�V�T���(4�)q�歲]z�Y��fo�f	|��ӊ�w���˖gK���h�uR ���U�=�������w���"`c�?�ی,:�5�&ǐ�fb��a�}����s�-1N���f�����H�{Td��(�+52��z�$�$ܬ�Kю���i놶x|��K����ƌ�v�K$}���`���_�`s��U�_4]���~�T��@�ա�2lj�i�`��P �rN>�6;��M�V���GI�O���VXkyO�O)v*�9'M����a>T>��K�T8��g�a�όr�.�Y_���q~T�$i�x�̿�,�O0���c�T���Yٷ�~O��>��� %X�H��	0�w{H��Ђu�b��I��w�!��V��ZxT[`��1n�&׾Is{��ϩL��&n2	ڒ�e�\��7ڣ���heV4
�sJF��{��SA��2�~��޳��we���KvI���V�~dK���LGd��c�2ލ�7
�"�&�j���RC��"c��� �(?L�ON&���MKd���~��n���[���B��:0f�G�f�X`o�Ȭ3�ԁУ�G+�ͯ�$���3P��Hv`�|����16�	,�.�HZ�Ͷ�r1KY�-n@��-At���6�g��!�y �s�l{��ʑ�U��\Yy	��ٶ�Й�-:Q>y�dbuh;����I��
�i?	ψ�(��j�d��PC�݈��n��� ��lB�@^�y0�g��?a��r�o���˃H�)�8q���'�h�<�
 ���ol���d��&��9,&���=e1����\�w5ի��w����^����XFL}4+��8�q�Ԥ[B������j�B��Z�����k��$�	� D^ő-s��<NsN�AY������׳9��I�� D�U�Q1�l�js\�=����]�ek`�������˂u�>Мa��bk��z{n�,0h"���V�%�[X�=�[d g#ʭnfm�i��|X�٭�ks��+/%5���w�J�r�
�΋U&7J%_�s�����s]=�6�@?��y�%�˒�MQ��j�{ �iS}�%����kӸԝl��1��1���lp¥J�D���f�{j�xn�V.�b��zy����K<i�l�XfI��Q�d�U?9�G4*��Yj���윯!fg�nQz�~4�#�@$H�|��M4�S0��v��=Ǒ^�r������P�2cP��͗lJ�ٌE�(`�iy� ��\���Y�$�# �����beQ ꁄݡ�l���zS�k�i��ڗ�f���T�%%Z���,e��P��ᰬ��4����Y��~��a��K�h+� #÷^^�n�s�ܙ���9���!3B��|r�[�yj��^	��8񁞱>6�n.G�+��${��&p�f��ɩ[�C���/6�B}(��<���-r �Z�Dg^��b�s}���]����c��������lU���<O�\�%�W��'{5bIqH�.lGq{�܏I��̧�jj%�C`F�#�����x�s;�P�ρH���y����&��~'3��e��IF�HfK��]X��|�k�:�@��F�����>��T�X�i�j���/o�^�4��O-Y("!��_(��(T�*���nB�UJ� �IRIf5c�A�%KjOj
iS��{�b4)���a��NʀL�*�:N~7�Z�:�t$'@�f���X�7K�[�S����_��W<���}����nu�keл7q���y��ny!c)g��2�A\g�J&3tO2��!@�^��N�<�>���
ж�o:�[
W7��S�CU�� ̪�G��E�\��O-�'�z�(}v��|BaP9+/��;�Q�;���rԝ��c��lS�Ӷ։XrF�<�Wq��i��RK?_9��A`�UL��gZ�%��֦��)	�aTCr�����_�MG��#by"�w��B��P���Թ�,�͘�^��x@msC�A�	_0��3�7~<f�W���HK0��ݲ�<���2�s6����e�Dy�e����E��eF|Z	`�)�v�6���qJ	����|��ܥ���ȺCY���䚯�nI<�2;��	���i۔`:��ɥy��ew�D�s�cpc���n	x�h�q4f�3A�V�� ����#��CHqp_CK��%�KB��,�Q�N��I� [�GMe۰b�l�M/�n�]4ź���+�aX)�R���( ��b�����8�+�D$`� Q�\�������?#��D�@[����ʻ�)l�P���J���vq�i�B7*L��d����R�F���`�&�G��.�?@��"3���G��|C���f������lY�MJ��?�W������hP�%�؄���]�E�QҲ�1�m�X�^��e=
���v�����U�`�'�t���{�<b��p��}��P>���Y � ,������.,~r��` ��m�/��d�p�S�pgF�1j}~k�3���XU�ٟ �H ��/�T�������+g��ե}!I�A�8ʗۨ�����{����`{������G������t�п���	D������[�וS���V��MjAI��+��HhK�����r[ka�gT��2@=}��a�>��Ta�ǱL>>�x(C2&A����U��<M00��ޜ���x4����:����k���C&I6��9�ybߝ�Bt��&pY}�S���-�f�/��:����ac��U�!�]k -r@n��:D$3#A��Ռ0��Xjys���|�w��ff"��I���@J��} �y�L��ni���|�;c)�B��̽��	-��w׼�$&� ?�H�� ��Q=�k����m�ݏi��K�A��4g�&Q�����M��6����~�а��[�ٵ�l�ܠ�q*vT��	�(&���<d7,z�>Ѧ;��-�=b�͓��r�k9����ö@9��VOJΌ~�9�t�񉤟	��I�{m���z`����P��Lxlu�A�Ln5APsO����� '�(� lY��O|�u�:��Hz�IMh �k �MƄd��Y4`m�fɑ�@�|$�负ԆN�S�T���cv���i	+^E�4�����;��1�	Pl� �u+���"_ \��3ʣ��ϱ�9 �mNf1h��^�nAn����摫ہ��z}=,K�ʲ���r���dr�[�h��g5�2W�0)
?q���Ѕ��)\,3H6�Gs�ۡL�(����2�X�
������b֣ѿU�w����>ԅ�np�7c�Ok=�A��k=�v,�LT%Vs��6гG��~��!�5���#�)��ւI�?y�o5�l�*$���
���#c2H�j���`T	s�X,����I��wm��gΦ��������"Q�ͩ�s�c�`�8G�B�e[b���H�Y��X#��?c��f
����ONn�. 	����L,��*#���c0�#w�d��}�X�&��A�-)~�M��bsIn��05�e�ޱM�J�{������LҒ��<����G�T��{�t�b������Qm({�n�r�y�Ǌ�_�9��@n��i0Pkئ_�����dV� *�?&>{m�0_}4X���1{G���۟��Z�~����J�T�gGX�:-��<��ÿ:l"�cKs�aH!�g
�}��k�jŉQp6��:�.&��h$$[݄�s�/��i�I�"�bR� �^;��]�OZ�	�Q������PX��6�H�av���d
��_2X� ����+���[f��b�N���M�[�4�#_8���ٕ�Q߻�,*eQ��j	%?W���UMS����=��P	��wvn�Hb���N�k�����Li	���\~����'��Ɔ`�N�k`�`^nά@���3���*;������pO�%���m`lr՝0M'֩e�4�Gf�J��9��3��C$ �fj���
�z�}��7�`���<��P8�'���9�*SQ5+Dn}�>T+�.l�x
��]���Nƻm��7�F�@E�p�	�K�1�)�~��������{�7O�|5���cm)2g��OO�kw�בE�|��b]��=�.�P,��7��*&� ���n�J�婯eq+c�?C�ۋ	 b��c}��ܯ��y��y��dIR��I���@����d���Ԃ�5�`d�V��b��k�V��E�z�e��ּ]�x<���=����J���3-�����P6=g�����=+��41)7�17}[��C�JM�
��$��R�:
��"c_*��1�y=~'V;m�H}���L��٪PyEJ��U�K={O���a�;%�n��'9�~ �m�~�.$��J�~�|�7P�P~����2�k�
~���n�!1������Ϙe�Y�����Z� ��{�E��`\�7�/c��5�25�;͇
3�˹�+�3�fq��}�%�����I�D*"sg��3ۓ�Aφk�10�}���<��C!@ Y^��Q����M o�'�.>@���Lt�O.�!J�@;�
YN�# �1�H���^�حu���v�k=��M���n�rpу,#\N�t	93Wj[�W萵��b�b��ݗ�ɤOD09�|檼ը%6�ji�O�=����u�dɗx�M\Ҹ�����P�E4���8���Q�@<y7�/�&�OX,�w@��O�zg�S��2�A�A�``��H��¦�����11S��4'��i��X�[�\öԩ��ͥGG;\noU�
0�`�}���#��{�0t/��g��P*n���F ᭘(�!4�=���b	k�k�dzU���a�L�� O뛊bnD$����rX �=�#M�YL�bgcG�Z-�n�`���`����2��_�& o);�h�q�E �{�HN&=�_t�������_���C�˿�k,E}2k��ɨ5|�.�Cf~Ac��NA��6��p��/ ��X4�����aHL��V$�W0Ƨ ��K���U�E�σ�*چ����5��:ޘ�ҿ\��4��	�+�����>-7�A	�f��2��l����V[���I�a;��D����S�kr?]\�	*��Q)S�#�m��P_lL���t�T�RR� �M�L�%3������g@�r��4ݖ�ʾQ X��2��#�v��y=f��>�&.k! G�tD�ղ�Ȅ׋��z�L�_v�����b�c8�{@E鮟������7y��9��&�W(7�' J{���~G���#�=4�2���[������/�;
�N�Q���J��̬��OY�$7��j˘3��0贳}�`I����f��A,����KY(���t M���R,8�*.��u ȅ��/�N�({��jG��m��Ѹ�}x2S�Cb��C.�oc��Mr?%����#�dkB�eKc=�+L�9� i�JDHȣo'm5��o-c��g�
��+�J��M�8O�a.��?l��<���/��W���:�e�����<�P��lsȱ���Z) �e�C��ld����T1+F��z����ϟl7T0�U���|����1���"�1+�)țm!'�?,R�Ɣi�?HB�%E�ဵ�~h���Ϝ�٪��+��O�P��H�в�x�8e
v������c�������M�hb�-����7�x�
ժI���NT�*-��p_ni�T3�����
��s�Ǒ���Iۛ�|�~�}E\7��\��.��w @B�_�ը�����h�d�+r�h����y��߂jmd�� �ag@�G�����ׂI#����o7��P=|�{�l���==���o�ٷ0Yd��^�����ADRf��	m�;3F�Lyt�n��3�(ܐ�=|�:Q��s�*dy �V�8��M�I�-w��� ��n��k)G�����B
>Lwƈ�15�6�x/4�����c$� +���	p+X�T�%c��Tq|�Џ��a�<������G~���ڒ��M5��8�:�����ˣU��x��R���HM��Z��2���GE���cR%��mO� e��*��d6w�W+3v[7��@(�;�m��\���rGo��>{�j�l	�h��<�����[�6��w�K�ơ��X����r���]r�'��R'�3��>��GM$����Ķbc)� 1�<	f�z��b]V�dZ��Q~�����z��26Н�t�^���0ہ�c�v�5eq�u ɉ��a�(w,��*Y�6|���B/tO�n�L��� D�gV�w8�&�������K@GL������p.��ʞJ:!��a�X��#��
��*�ɏ��rla=����D�?+{����M�oh�H��	H1P,w�2ӟW�;]sX��5تO\R�9��|z�0P����������Bb�����O��T5]��0�J�vݓ��"��;���E��nޮ��5Շ�9:/�{Ӷl��p��9e�"KF�����GBO����;LC�ij�?<ˇ�oe|�Y{=.����G(�-�ـW|�����Y�4	)����G]/����ֆK�X��QO�+	e�ˍ����wD"쑦P��w���7Vz1e����A~����í�?o�l�0�E������F�6f����5��?i�F�\�+������ ��f\�')�"U�e����'��uI�"�͔��T<����/=%����'�O���m��葆�XҀ� ��@����1`6�@��l+w��m�z&��X�A�b	|:F�D��V�)Z�׮�$7�V���6����~���>9�{��5�c$�k[CVx�nf�-&Rz�%��n��Fɉ��<�s�������R�I@��*��l���[.X���8M�FX�D�n��KK?n�-h��7�1*d����I�,z"����ω��|��Ű���t vA�����,1g��/���V�9�t<~Qύ^�|9��..�<?��O�!�r2G~�P4���D���˵�O۳|`߹�X�o�}٩��z؆�����_1f�I��WS}���֢m��_]߻�ڦw���/�A�p���,���#/k-�v���g�G��bp{Y���'�tR<ify+���16���k�tJ1�f�H�<��b���}���HN��E�c�D��ܒh�jg�$����4�]�Ok�����V�]m���P{�S8l�h�� ��MCy�@��=�Uw���c�g%5R��n��K��ܽd�1��m9!ŘC�y���LSge`�r�b�)��,���)_���B�`����^#K�g�G�?�	��&�<��m8�����;�S=6ſ�b�1|����o�0z
+�0絭h>_�}�fT=Ty�Oa�?c|T��u��)=7"tg�����j�G 8|x��'}n��3g��̃��t#ԍ���L��
Y��Fyx%(=���g��<	��.���n�5C�Y���j�I�����7u-��^(���H��~m����>.99v��@��p��b���40�Azn!M� ���ߟEˁ�N����;{O��k���������R����Y*?��ٳ��b�ϟ�bG�38j31�e\.�&�su�������>���-/*��|�x����=�D���<�Q�� pАok��a�}'l�������5�.V�VPi�]��&1��	�
6=�Ć�f-���?pIR�L�vA�L�=��+�>�9���w���X	��7q++�LP���#�^�zA�L�ⱥ� IY����1"ݑA��PQ^��Ї�P����&�5'dz����8̌�%`����L�X��~��$���w�d+]�| �����dT�ǹ,m9h�K�3g�㎥<+��s��f��a�,P��ɽ���8`������L�
d䝎w�Sj�Ռ��A$�`��Ⱦ�nbTY5��_�Y���jm:�ae!:��I���(�_�ݘ��V�����`�V&^�������q��X3e��o��lJ�l�[m!�ף���>�\���
���r��M%&��'��X������3�[�:�������ἢ�Hz��T�`�yyy����n����W�\��{��
sb��|���l�P�-��a�Ԕ���"͠�k�5v������?�����/�������l�Ĥ���Q��%K4π�m�@����W�_�Ch�SP��k�6��)�v�x����qo�>�x?j6j�Bq�7X�{�S8�5�� ����4��^��c�P�mw�|�,�� -�{��FK<�B�hi�xh�2 �X����C�Y���#6���k�)���x���/��5j�Yg�:|rN�\�4%���V"J��>�g��z�i�=�`C�&��^{���F\�� h��:y���w�!��;)p�O����	�H5;hs�*(zT����R���5%��.���e��ʺ��<E��ʢ_����������������������h�!^&�*�H���Eo�&�� �WJ霅��u@��H�J	�-�>��<�u<8l�?�m�	X2vf�a˝p*(��t�V�������o�MCɢ��ϴ��g"4P�ӬOHkE�<���ұ�a1�J
-�b����`�H2�s�\��%�J6�J1��V�����b��ƌ�8�=�&7�#���NN���o>Ɂ/�(r�Gн4��G�}�ԺXl#dn ��}ϹB��,z((V�([��ٛ�B��W}|�a�!\�r�� �ǃ^�Ƚ���n��al�������	���͟���KL�����|�&s%�a7җw97�HL�nYP�=�n�s���@���0-ө���i��\
n
?�<b�<h�O�����X�(�Jf�u�rxW� �S��{*u#-=�H��A�C/���ƊP�����>$L���*�X_5�3�naJl��� �t���q� ��H���i@ ��S������[�F�Y����	3��%��=��+������1�F�����Y�d�
����ev��?�g���"
�Br�*����>kl�Zv�E
��Gism)��>���N|��[-j�TW<>#2���|TA�|� �>����(�ۗ�<�xj!jI �� av�kH�
���"�d�b���J����C�}�9\�/D���E&;�L�2a$#nss+÷zΰ���U�,w��Z��Z)Å$�N���U4
J��K\sPK06Q�n�yOuʲ�!�x��Y}#P傶�|�ɉ2�;��o�g�S_���,XB�jqt`]$T�̻H�����XL��,�,�?��N�z�����E��{��au�]�=T?�\��f���/�?�᏶��y���
7r"�?�ʚjh�N�F���Պ\&�ڊ�sb�LØ�WLP��͖�[��b�se�������)a��`�Tg��A����r���"��:�]g������L���Y�����g�ڋ�����e&;5H�x���P��ˠx��#Y��?�����&�c�7��9��ho�C�2�평�N�jԏS9�v�����y�P��Z*���Vc�b�(a�9K���"$
�t$s-�:��Em���XQ�G�i�-�ǝ[��;�a���#.sB%b�i�i=�&@3�Ҝ�e�~Uf���Gc���J=�j��,���_X�Lu:���ҷ��
��ɀ
��~��H�U��*�Y%�����G�4)�Ȅ�����"a��O �i�e����;?1����.�u@�k��ו�рX�#���+Y��h�j-�(��������Q �/�9ُ0l�V�������B��e�ڹI�mMD���Zk��Vb�NC(�F�Ő)a��5Lv]�#S�Q��v���Vr_���������K[�g�2��ҷ��[]|Ǆ!^z\_��%S��G����E���EM���6�+ە�N�0)N/v�'�1Iu<�2��W�E��)�X����f�>=d���~�� �2�����Y�������fj�ځD�KF��H���.q���H�nL
*����Z���K��N����Fو)���60^�3�/0����{������"j[H�&
��:t�β�Xĵ{^S�F�����ܛ��9���z묿�U`��A`ŋ���^I&@׌K�x��p�� ��	M�c��	���JX-<£)�P�(�)��>%�UL?��{s��J:����'J�@?/�U;����a�Bs�2��f��:��^��+�E��T5��ӧO2�7��7t�j��p�ڟ�\`��h�א-~��u|��������RI�O5�Lw�ٛ��-���EV�w�
���=��Kǻ0Tf�8�����l�4�a��gڞ~�$����Y
����';;�0m��g'���*�kW�q�O��KT��Ύ���T���PsSB6���_��Cks��~SS��}A�%�p!�ـ�������Y���G��c�䯗��#.�\ѻYP�v� E�BPY<��7����+a_�Z�������� r�C�Q/��TTƜ��n�Wg�B�&�`s��P�W�J��<_����zTf���6P���vj]�Ӓl���J?�~���|��,&�4(_T��ȱ�(����L�O'��*ok_��K����-��*�i̇0�����>����m };E�?rR웯�������$�4��t7�"�����Cү��$8/fAw&��*��g�==��a\�����qH)|<,�4�&�%5r+Qwp�,�5�Vtbm�I������,�\I��Ԣ �$�n0�e@+͚����.߇z��0Ϭ����ϻa��u��F#H%ްs����w�F�߭T~����B�X^amK�i�@60q�nZ���2�9�- �m��Nm��*���	�ԊѾ��o�����}�HW�l��'���f�`�ʻw��M�0�y2 ɍ6ިYa�H`�{�	�9ج�����;5��濥.%M�¹��M��I�[
*̟�6����M��=�����o�%Y��K����}_��y�,�|�Ym� ��1(�L�'�nsX �	,1�\�"�u�q�O&�{��e.S�K_�V�[�?�w�rr5�c���Ԙ��~˷�E��R��5>�x8�z��r�g=c��3��|�c�drHK����z/L��2�q�rG4O��pG�Iz�m��W��٘63N��N����ⴉ�� �������� �Nڋ�&�{|�,�Dݿ�:����YiDn#
�b>T]Ǐ-_�����-}�>�X�7ط(�ob�wJ����e�\S��(S�i㲒�)�"o�9N��ǻ��F]��h�F��/R�� &���䠬V�L���3���~�3����ڣ�vg�zS�F�d�,y�=�	����b�t�#�����_����L���$���V�PJY�(08�X�_\
D,��:��ϺI�����?#dL`�I�U����������X� yv^f�������l�U���R��x�?)�Ɂ�d&��ZN�4�;��9�i���vD�g��M҅�f�J8�޴���yO�7ah��{,�j|�!�u����kQ1��1����d��mS��j�a!�3��Te�����s�%Q� �f�L2V���L1��s_9��S��xC�S�|���c�����]L~;H�Wy͠�C��|0K\g%gߩ$��$��}�� 	�˯��mN�,��)��r�"�#*��΅0��o�&��GlY����M��w�d�׎oQ���]�o{�L��kW�X$�w��O�n��E�ۈ5-B@\o ���.?gvg`z�P���^W�^E��$� �	D���tz|Q����C��1J�%�{��)��5ƈ��a��	h��nsX�T������zNB�T���tA� ��������[�7��̉����g���`�}/ ��ߛ�#��s��"�l�.��	hM`�� �_��A�,v�E+���PK��% ����.�&Y��N��|6+�/�1��òM�/3(b��8cP�	���}d��P�9p�G�����e~��-�n��",�A��۰���A9%aX�ܘ�� �~'Zv����<��=�K'Zkg��=P����)��215�`��x�j9��n��>?[T�� H
,=�m�.]X��.�[�6�epBV& ms��_]o��6���;(
2�J�:�)�Y|�n��wZά4'��3uޘ��e�{w�`Zg���\�%}_���<�N�|YJK����<zF� 4r��3��ݝ����A]�=ǺG�W��������w��廉'o0@����'Gyz�,S��'��F(X2D�ݶ�C]�-��)[߼�O����� ���O�=�x�-P�}���� �](3MS��Iӷ�$�fj�+���ٖ�-Lt�.��TW���Tm`�< (�7��%m�aY*�(��M��v��٨f�Ζ©�|Q�_�dtP��-�U{�N;o"S�&R,`HP ��ūz��P���b�(9�d/���k��14o*��Y�K��1R���5=�D%'M�49�'Ӊ��rjKN��$R�7�h� 1��t~ �V�Н�Zm8ϰO��c&(�N��o�)�`�gj/�?kz�|'���؂>TG��c�B̎T4�?�R*q��v�>��P�n�Q�=��Q�&�Z>��4�D��i`���r�R�^h�t4�2�,���d��/�D�]��%����o�S�ޏ�����S� ���������ݳJYr�[2��]��1֔�hǻ8胈$�=��L�@���鍲K���Z.�k�|���ȷ�@Ւ0E�{�,䙖l����k� ;�2w}E��-^?����)
0���WK4�5|��,m�r{�9f�2<m�냶��Wxz�4���U��daV���I���s�[������y� ��v�
���C~��g���_n�_3s��njh�[jG�,�J+9&�E;��0m$��]��d�&y�j2�R;��!g0,6m������.�ůͽ�z)@�wh����m���Z;5<�x�6�-��k�����v���d�N�������~�w�m�^���)��,{�1{a���-H
Z6��պ|L�B���>Y�J�0�g�bܽ]���A��9�"9���L-�~/�lsV��N"C���xBj��#<gT���"~bɀ�
�9�U�8��?P�d(6�!�2 ��su+?����o	l�M*3���m��
\�\ƒ��^�.n�	mf_g%BbdR�(�x2�����e��Q+��ӯ��*��~>�|����]߯ϵD�1a$)��;
��e�H^����R��s
��-:�e��Fd"��I~�Z�ҏ�^�z����x�O�~!A?��5�f��|;�0�����i���ѥ6ak� "L����A���M ��&S60������ngL"XH]�-A:['�J�4�E�ҷ��2����z"3-����-G�o�nN�?bc�މ���6dR���9���ۜ�n7�X�r52�m;hݤ�����2����i�r�9{?�(��$�Q_o�P�en"�<i_��,d����A��K��})�-`_�c<&�?��O�lþ��I.�ob��u������9���6������ �i�Q�����T��)�Οl1�$vg�ήS��l{��x����@уX�	���2�{��э�J.;��n�i]�:3�kU�מ�$�	?T�@��!��{�UE#���B��7j0���:�~==�ܦS3�(<�� =��o�GQ	���i�6�Q�Oi���|G٩Y+�>IMOU(=��w7$in�Ʀ���5�&��yޞ"#=v�[�:Aig��e�-�v�G~�0c�����-��=�_��OrV\<u��8��k \/���3�������Tn�]�۞�X�rV�q��͖��5 �T"�+,�K��k4.'�-����@�o��el=�����WVɆ-���ҒӼ�b�ǆM�1�n����ۜ�x�q ��mo���&�[l0�l�-�W��Ү���Á��v�߃��:E���б얉X���ڴ�r���ۄ:�C�V�Zl	r�,�P����P�q:N��O�jq���dy��y"��`.2K# �9�xH_��E�!�G��:o�{"%[2��LK#�rumn�MJ̶��^t�V%����R]<�C}�d�KO��p!��#�b�u$c�F��ʟ-X�����]>	�}�-@�.R�M_#��
�K���)�v���P�)��K�R
 ��ԨM�i'���Y��k����Ï?�>0f6���N'�eN�V��^��ַ�>7��Lz�lR����b��l/�r3q�
�tp�391�P�X���_�7]�Cgj�!<��6�;\����6o�6���)і	��H���wAMfv=r��xiZl���Ep��a��-m��8�y�ة�Mm��]�ιJl2��`A���sX/���l�u��P��I��")3�#��&}���F��c>?��C�"�p�e��Ω+�� }�}����m|��֜��1b��]c�����t�������Lh&yI�/E�촱���$�2�d��jO�1*ы4�%#�c솀�G�����q�x���
|<.ub#7^cߐs3^�}�"��r  ��mވ�����L�덥�fd�?��lG�`8Oi����C�|@���[�g��1N�����"KP����#ho#�Kg�{C�U�wO�6|�zs�V�P>ͬk��". a�{�����}���q�,^c�U'����(��ۺO����b�W��V�F��@�>h���K0qc/��Զw������hZ�I˗�%+ꦼ"��,Y�T]��Ii��z�O�_��0�5�H��H�/=�7�kYO ڶѿ�W*�:�"�>a֧"⢂�r�� �
Y�����yA�v����ˬ_�ge�C����q����W��߾v`��)v�	���3��>�`�n�������Ϋ����g
�Y�b4�p҉�����e������!����=���k2��~o�&:]�hhO΢u��{21����Z��AZ�P��'3�} 7�����ox'��Z���_���ɖ�5׉�ushm�훼��r�2���ɮ������ ���O[S�r�N������HR���s��۶ |8b�����!0d�����=��r��6B�ox*���BP��3���-���$Euqߜ�H&Y�ET|�S_/?�.�sn�����=?��E�h��]����\�R�ۅIR�:��,$�p�ڲ:=�/�_r���t~���Br֨g7�ⅽ�r��Z���2)4g���1�{�K��ߐ[�60T��܈����M�v��S0��?�AxfWcZ���`�f3�b�]ˣ�tD�5�<��V��%ƚ~2�b�I4���Ckx0��&�v��D{i[�!+�^�v��5�
P� ��걟-�qa5D���5�����P�#�LUɘ_(�ُ�c$�t�b�&��6��,&��R�x�{��J~�|PJpo|����ܶ����q���9<&$\Z�6�+���������W���#�]"�6��2LOv$�?}������=&&��gR �vODHM?��7*�%.�g3�u��3�}��!w��=�/1C���F~m���EJD\$�4�w�Y�;A&㙕�3��������`�W2cq�$ޣ6�O �k�xO�"�xR	�o�h�э<8-����̔�hSh���.zJpԨ������zZ�6�}��V³<a�k<,��]� n�}��de����� %�	>�� �+�	]�W��[]�L{�$+�.;,�+kD�f���5TNj���w��o�`P�E��[�8z~~��u2�Q�c u��(�N����!��¨���Ev��0�K9�}�P�j�`�M��R�~�Q y���L���5����_��gf{��|��n�z��q������RJG$�T�W��@���~?������pU����tL]u�	-��Dyz��{��\-�,_�|P�+	$�1�UϜ�[�_��/qyA;9xG�V���4���W;&q ;l�16=o����4��b��Zb�'Fm+�����e�~�v���s�_�j)8���S&{֍M��j~f)Lf�UXIާ�,ZȻ.�e��Ɵbyj�v�Յ!���<���n���Y~���w*��X��|�z0��Ӊ�\s����?ޮ?|@��(z?�'���|G����'�Zjݯ�E��GF;p�j�x�va��k���et���A��p�q����}���f텕O�{�[^vg@�%�Ĺ�������~�*�>~4�v�^�}N`/^X������pSD�>��|f�?�S����	��{�����M�cf�!3/�/7`�l�g?ŒDw��i�8�n�����r~���ϯQ�٥37]����X.9+�j(/���*ps����A�5"�r��Ty�$)���m���)��Y!(6΍��e��ݴ�k2�d��#�>:�P��=F,Z�k3ޗ�FFz|�U���Y��AZŰԫyX
��ZP���~�����Ab�)���w�����7GY����su0������	���o�e:����ӧF�,�# ��dn�|}}- ���MaX��f�0����"$�.eM����"(K���Lz���N���V�+����q���>�"D.av�8��a����f���O�b�33oS�[�x>M��r�����(�_Uu�2۠%wX�H0��xy9ne�怷�_d��\ ������1�j%�w����v�E-W�7o����ٶ4�>���.;�~P��������/�����)���7 K(]$I)e9����l�����J�$��b��)�4f�W�e�[(���/n���Ė-�^`��ճ�[~uW8i���@]_VY�v<P������M�iyhC��Y˦)�j�
�'ty]%�)�a�Aq�����\kv� >���=Y+]H���zl0G�R�6q��*c0G�>/�gω�.3�'H���|?XZ��! ���䰜4ۍL�kG�X
-�7����?�=���+���f���؞I1<�!�	�Hs�w�-�ݞ=��H�($��*�,�ʘ�͎r�[c &��{\�\�	%lq'@�G�'��M� X�R�빏?� �˟����[����2��V<_���i �d�d�Pg0m�l��O��3���e��߷�*9� .��n���ܑ �D�E!e���p�xĽܟ��^oZ"t<4۔�6sxG�MF|=l�@�?��Ҡ��'�����QW[������A�N0,���Y��ߡd����a�ϙZ� �-�}�?�|Ѕ��E��9�U`�.�|�V7թ]#��|�b����L~��G`�kL���.(�(f2�

'� ӋL��L-d��%}�sj�su���{� ['���ʜ�]@�cf��-�|: ���7M�	�fj��:/�A���b2�wm\��m��Y���]�}��2|����\���"0?��,��.j�z�{���N������^�q��Ly�왏����u`��o���ӧO��.������ARP_˨�o}�g���R���>�x�]OG	����;ף��]$��q��k��P�;ԇ�/����!��L��Mɡ8��N���!R&�?�|�2���ό������ߙ��F렀�"�ھ�K�Oa����zY�A)oY.�Қ�kk�Nq�`I&�?��r��՟ح��O�)�<|��j>+�&���,���U��%&&����%u]��[ ]$J�m5dcXa��o����"�@M�D���@*'V.M
aBJ�<Uw��H�!F�\�x�+E]0��C �͑�.r���<� 0^�j)�2���+�>�eda
t���잫��R���Q6m�	P[�T���Rx]�a���nz�Z��� ���zcC�&@=�n/��8�l�e����(@U����>|�魁���?f�bU�ޓ��&b���O�ی1oS�����.-�����	�b�D[�:m
��m��M��7�`O�.mK�<�J�a �����`'�F�>�=�����d��5�"\
}
�>�&�~ʃދ	DǣRu$�4�/��5?��G(����6MX�m�v4[4�Ҭ+��:.2L�=b�`e���Ƣ.����pLn�WP$����m|�؂��������������B��ax�3E��)W��,�,:�x�L��
���_��oa��\�; �іקk�M ,�����_q<v��/�r����
e�G����i2_����`>�£��㊀_͡X��ͽ�N]>�we�4
��h��ta�e��i8��C���	�X@>���	�m$@^CȲ���� �W������ �F2�Ƭ�f��l3C��l�Y�/�E�B̞��q$�Pn��z��i�N3�)Gcfj� �k�=+��~����ܽg��F�-\� 9A��׻���x���zoڵ-+It��p��Ar<���h8$4:�>��e~.s��yPY`�����d�������(돺��ct����n���q�_]��Lm�SZ](�W$�#�K�L���޷=�O>�CZ<�7�|����#�D7Z^�,�3�B�W �����`�� ��gÌ�kh�m	���q<]�)a����X�F>���p8��o0�m� �1���X�y���G٬<���&�0ܚh��$��������H+fg 1Y�p�Q�=�����l����ͪVpm����	���sr�D���DT a� ������
Pm �XЙ���x�{��@�ʰHC7x�ͩ��-��<���y�vJ����x�s�ٍ?r_���<N�]��-�G�Wtc�l#�,W��q�{
��{,/61��m�A�D���/�� id�ϛ����jVi�N��> �@t�oҔg�����8)��(���1�+���zg�
5MÁ@�I�77$������~��ɌR8`��0I��S�͘`��N�b\���&���kw���$םf�D1�7��3ʜۤT ��PQ�8��N0�e��`W!�/ �*�%5�9�c�bRc���֮V`3�4����-`�G���Q�%3-V�稳�үݒ5�~���ɋ�Z�����p0ө�T��%���!p�a��@���9iÕHK_�k7��X;�槊�H-�槚���o�/�`����X��M����J�6��  �E�-l�
�
Ⱥ�H|R��9�-u�����l����ø��P��k7;�K�o�O�f�$ui[|�~"ڎ��h�vH�ҀQI�nqI��k˜	_	Q�c��$�@�'�aă�K<�1W[Pj�*\mT����"l��ȝ�Ӝ�3����6ǚ<�[{G�k4[�*(��B�7�C��4��"q��%��0� k>�<��h��q=�?����c�at��f�N�IeQ(��Ĳu�'V��-�1�=׍�{T,��_�(B·'+��SU��sAp{X�]fC ��J��`���8n$��a �k�����Rv5�6�C���A����>g0�5���;a�07F�$V�Z}ײ�:��CuT
��T�_Ir���9Q�,g���&�$�c]I=XO5� ���J��O�CŢw�O��OU�zA��,����9�m�gg��.��ґ7�K�|��'qƿɞ�[�.�����t��@O���Zw��o1��,�a_j�2_qs����L� $aj���{r����0���.m��x�k�z)�q\�4 Xy���n�:D���Е���;��Wu1��
z2uR
F�qǳ��#��"��]��c����� �F�I)xF�֜�KiPYg]��/XI:�I`@]2g� ��Z���ޖ����+��z��zLm�o��5qP��+�滑=C^[!!���`骔�w���PXH����:V��;��qV ՟d��X��늡��J �_�"��+�f�8AA�f`�j�%�Wv��d$�Rl�B�v�٣Ǣ��;��"?�@WZ������*�@Kh���������S��y;�.���&����0%*��:��>�~�)�zѵ� �z?�'���z�؃����)�IZV�C��i��ֹ��<G�C�⤌���7>?٠�8zQ�i����)�k�xt�A�Y?�ǌ��?V��"�/zs�������T7MH�ϴ>PӼPE'�@��9Wp�<�b�C��理�y�<��$��}��5�$�ZǓ�P��Hҡ�+*�NV�g=1�DEˮ��)���a�ѩܻ�j6w�FC�ʍ�H�=�����Ħ��i���Y��I�4}���C�G�дv_KX��t���M�H�\)�	؉�)�#ё�,����zI�Y�V阘�F��EC׆тfb�(X�l��/sc��zCaz]֣�>�`t�H/g9W�;!:�%�Z5�Y��X������ꂲ�`i2��_�R<24fU$zoV��p8Ж�����'���֭o6�\�+MT� w����8��ã���XEu�F�E��R;ߠC�w��3Q *P�t�u>�e�x�s11T;0�[�Թ�㑠~X�Ծi:�C�v�=���O9).L�3��������A�K��]�o���&��>&P #����>�t���ضu)+Q/S���1��Q�Xr+�]�2�j̍��Z�b�?n^z�"��h��D���-D���3%R�aqw��FH�]� U>���z���0�K�)�	H�>�?�{�.8?9#���=�����R��5[څ���$�6�܋��!�y��o���!x�j��9��|H�-�,RB��v~d��~�[X�#136w"p|J(�ٸ@$PK
��~c�E�Z�M���x>�2�~>ᚥ��5㋶�E������u��rDK#� �mǙA����X��=��u-^a��bQ����VNa(�/Ʃ���"�݌S-� �b��L�?5'�>�uuC����/����%�lt��9;���?�z�d�	U0=X�+&Ʃ�����?��d���]�] I���/�k�3a�fK��l!!:�;�i�?�ĸ{�>��Bd֏"�/���u�J0Sb����"=Ug�
��z �Js5R�YUOj�9ct*Bvc
����Ƴ�i�۵{�х4@���Pq��h������ZҬ`E����W��U.y+�U�1� &�?�Iن�Ap6V�5Gvv|G$��X�h���U#ł�#�$K(�����U(N<����Y�Y�:����A�$�SjQ`���qo��0b�*�Mޯ�Әd��D��R�O{�?r<����O��}�C�R�	�� `W��u!���s{�w�����ҹ>�D�33��h�f�jb��=��'�+�C�s���%���	b	?"��c�ú}N)��"�E^���G�ᶂ�ԓ���IQ @�� �_D}�n���y�J+��d'{¢��k���hѕ��{��b\٘�d 
k?Q0�<�zPΞ������d�Z��%g0��@�i�Du�B���e�%"V�p`�=����6R1nR6�$&��B~���iu8�����N�cC��s��h��9M��g��{�ܦ�����H���4�£?���}�� �I�x��Q�� ����'%5ା��	�hq��be�����"�~���X���Y֍J�b����rm+��EL�P����Ը��C1)a��Ϻ�'R5A! �&/XI���EX���E�p#2�X`,Ib\bɞ�luOe-����i!:��t�K>#B�s�Ƈ�˳%�R])��b��k����0¯�Ũ��+��p���T��4����U��{�����u1����w���W�䱾���V�SW-�����y!K+�����g�	"0��L��'>�C� �T�@�%�{2	�5��1/�r�Dp��K���� �t�>���h��!\����ښJ=�>B�J&� �U=�de�Ln������,�NZ��%6WA}\s��	��C��U�R�7i�����i����ˇ�Ws)h�^�|��秤�}��s*�fV@���ռfp�����B$q�~2�1gρi>7��i����`�>�	��f/� !�5���d��i�+j��x�BlK,!���~�Im��ζf.�|o�
;"��_%-7}�8;��U.L!([ �T'�����&�����8dMW�b�U����8�R���<mp	h�Y�����!��,i��v����kx9�$��OnM��1(>2�{�����J�u��2��S��p���9WE�:�`��|<c~m�Ε�L�=���uS{��[�����W��睼��yG��΀���������'�F��N�4�eLpוs�§���v����䀊��u]Q����C�u:��.�X��,.>�H�K�Ɏ���k�|d�}�.�(���xY'��?s��s/X���=�&n=vF�Yl���`���!~?w\����@/��F6(0�������%bi�8��}�����p�EgK_`d��w6M�����T6���Ikn�G�')����ף�n	�����i;��&�zr����F���U�-p�S��'��� K�GY�Q�R�^�8y>�^}?w�@\>���� A��o��@�<�����Tj@��ɮ��ȯ~_��1�S�<+��KF�0̈�`���
���ݡ�������i��=.V��#�Ùa�uTCĊ�e`l�Y�X��a��9�Ԧ�2�˓�A5OȒ��	�-_3��n�؊��^QT9��z!e��Y_�[�X%�=bsЗ�(\�F�P�����_^g	�}x>��Xm�]��@)�=I4��y�5�Z ���:��f�j�hh�{g ʕ<��Ͽa	�����-���P�S�2t҅~:sLu����÷�&o|�m�ŹV���6��j*]�B�>c1@��v#��%��!�̇A��~��$��q�P�g�Z�I/7�$�oov.���g�Y�Wi�|������n�W+Q��#L�`���"4Ry�D}�#%��=��t�x�>��2Eǆ*
DBP�8����6r�,QE��g93�&kvĞ}��:�,�����QA�ޑ͘�Ԛ���B��ԧi/H��S�i���ς�mXH�c�/E!)�!���b�:�����B�Z����i)�4я�6�DL��i�\)uJ������
T�{� � ���2I#�XM�����x��� �Uu�2&�aT�5��Nl�4`eQ�'�*�N����"���NI ���ꬉ��ᥞ���ک!~���-gT��
�KY��. �ޑ��G�9~P��p�j&.���k�S@(9䷴ W�����
B�'9F����d����J�*��?l �`��'9��x�͐�,���V�����u}��[��!5߭䈾g�x��g�+6���)�ˆ�)�G�{X�EG��k@��O�j8�>[��z��n�E2em[�<0耑�'�څ��X�'�������4e;�	��XtJ�v���}S���u\W�'�V&b�:��L�=[�,)� �gq��/KU����H�%� ��>�%���B��+e�������tk��}����|D�A߆8s~S�2�;@(+�]�/J���DQW5wm��rw'w5M�[��:�=���U���
�hub|�%X(��`���X���8\X�v��R�t��Z%��N�g-�3��i�A�}?A�<�$�Q �)9"ɧn���h�h�^�0ɸ�F��ū�$��g ���7OO|bٙ���D���Lі�B�Z�ɛ���,��W���ՊřGٔg��R�$n9E��#�.(��˺I,��yn
�z�m�g(eN�k�4|~�c��gu�2�&�;�[�oXP9�R,�}� nB$��Y�oO�Uҕ�Euf�W�nJ��üYte���B�M�:oO�A6'�K��k��=0$<�<�*�0�ƛ������J
�-�9�����ՐB��A
�I��)l��.DPlH5��\��6D;<�R�v�?t����5�<��h���.
�|���������Ȕ?}@��XCh��E2iO
�9SO>�t��8��6E�̡&����Z�]c�9�T��0 8��Q�Ĵ$�9Y��7��vf 
 y>DdG�t�#��3��"kӲ�?��0���R,֤x�k �7��0���3۬�P��h��JHzQV�I ��p�g�2S���1�O�i5�OI-��Pd�j#���.�T;e�RW�x�lM1���:s�bB��6�xjY��sd�b}Lih��� 
�hPa5�b���-u��:	 j m��?'�&���	�pԬ��y��rT�|D�="�)���Xڠq���8��kU��~�������]���\*����N�\╕��$�
�C��c]c�E�j�w��3�߶ ��關u�Ǧ��.����b�d����m��`C���|��Z!I6�/��ވ�lՄ�`T�V�d�*�����O��2��&�4apq�����{h���H�W(>1nS� _Y��	�?H?�\�V��܄������Ϥ����X���tgo[d�y	h�S@��nc���9��R��n˕,SXuP��Ml�'O��3�O����,�V�E+ �x��^�xIϞ=�g�'1��n�}�Jz鰹��:ҧ:Ч��{6�6!�X6������:��s&�zUu.������Z��p��ݤZ0���.�sD
#�7�/媞��eT^�=�3�����ҝ������ș٩����'��}�;݊��p���kB!3�-H�*f�\x��E���H�b�Zwj�{XY֣�t�iQ#uZ�.H5@3\�lx��d���g�{�_���a���b���(0'j��M�����-^[�'���AI-��j�(�j�H���bN�q8�%kް1OLY��bg�ϑ�i����"%�9\DR��p��"'�P�7@�|Vm����W��A)I���V�|������*60U5����W��j0�2y�d���u��2VشJ���cŃ����/#��6���nQ͢�@��\ֺ����C]c|�MŲ�|$�,V6 (�}8�'�8b�)�2�{d_�:��܄8y+q̓�~�@�u��q�<iv�L:�y]�C��.}TLWfI!����=�ٳ!��%[{�ۖ�7�� �.l���E���A�G�&`����.p��Dy,L�#���k�׻�N�j�n�4ۅ��\��Xf�mtk�z��d�>���5�t��B�6�m�%]vK:I��#_O1'�b���
Qܲ<��\�0���B݂��dL����V����I�;���߃�))��1��G2.�^�&�й�p^
�&���
��n�Y�R���]�!�M���_c����5�'֡��"KSY\E;ec���]ۆ��-��F%�XT�ŇE7�J��'� z���3�L�Ѓ����4I�pd0]��ho����%[�$	��3�EȮ��#�M�"c�3S��$c(�i;6{��,�����`Z�I�.=���نl�L�g�*
����TUY�����$R����K���TQ��LQ�"�&n�ʘ9��h���������<�)��������Tf��C<���G��DY�#m���@��\�ҭ�qZ�U���F1�E{Lݬ֨��2�M�<�:k����� �w��3��$�fn�]]�b��V�p�<5Xm�l�5�'�6�	Q�0��:@aP�OYLlb��
ȁ�&@��BXJ��:�2���w
���K}õ�O"������~��=��R׸O�](����V�Qt�ƨ����=`	�N�p1O>���l5� �˝[��I}����	���d�H���`0F}t7:��댈ն�9k2u����j�����4u0��Q��G��ȯ@�F28ro���ˬ�*������]HL,ʓ͢n5�PҚ]�p2�1� ���Y��@3�J� ���#:P�	��/{ɻ���Ztp&$G\;�\T��j���s��,��f�5���/�����
��4)|Mx������O�C5�oB�b��wZ��_&׀��[&[-�ң��X�^� &����,���$b���zFta���u ��Pu@�=e�����|�xAo��:?f0��3t�E�����K�:g���Xl� ��YDg����)L���^�Hs��-�ˌa.:�H��z8��Vl20��j�j�,�qvp%?ޔb�j5�sϭL�Gu�i���6[$S>J)���KaH�}~uT0bf~�����bLB͔tq�� )��6S�z9��(�U�n��ʂF()�@r��ڮ���З $n	�)�vA�����l?2k���;�:��liʳY�����A�綳�c�TH|��1CTv�J��HHt��	E��>�>��ɻ��gN�,�rˎ��(և����iG�2����y���Dq��ҧ���b��?2��\Z�\�OU��:�R�i��j�n�Ӽ�L&�ju3����X��$u�>�`e��!���[S��;6,�c�B�:N���nS-0�t�L��3� ��d�~ϋ�5K\B%0zP�نd�# @�I��E�9S�4곗-�ʙ\�4�Ҩ��Q�( ���`)����A�
���,Ku�&r.��Ȃ��  �vS�X�|����z�5�=��A�E����:��\΋�_#�]໗�@֝����)n��%j�;�(�X�|��`�sM:�kq�'s��p��ź�e�eFԷ�j�1oTg�O���V5�>���	!TT
�2�'C/��˻֥�~|z�0??��1��5��A�������Jiz���[� ��wZ�n��1Ƃ6��"�Z�u<nnvt�ۺ���y{�}��="O��������J��h&$����h�ju"W��J�0����ʶ�OK�16D,��#�R�c[zh�L;ϕ-ϕ���@�����!�+�/���O6*�N�Dh0a��c�Xך)F@@�$c����R���'�rMXUmЛz�" �\��<� �m�b�4	`���{;�j�}��͟g����+D���_����E�������a���AL�E��z�ֺT~v��5Z2�T�#ܹ!;.`N#��L���|��k�|��a�ј�sc傭�P����:3���� R<�,�,��uH���Z9�a� u��Z��o�F^3q4���GE�I@��>����H�E�&D%!�td|¹���3-#b����c����7 <��p`oD����Xd����g����>Gˀ��I>��K����nS^���!?c�;�ͬ嶇hu�̶ �_�������7�y~OϞ?���s��̆:�73�G�Ry�Q�C~����	����v!�7�zӕ��a�Sr��`
��5�'w���P<�-
.���}�-��M�	S���% `K%����Ui�&���@�LU���`�5�{5��~�^�C�P`d�"}��	�Q��F/�=\����,��X-�US������Q�;䡸����e��.��`l~����V{�bඁ�FS�F5�)�7�7��u�R$ON������\��Hn�Ɵ.�;��I���؞�*͋��u��U@�{��Y��r��PE�g@��O�?��g�R7+IrT#,�����[�[��E� ��:���N�*�`�q<~�`��?�E�/���2�p��Ct�Yep"����PY&���k�X�g��@Tc�����3a��ذ�o���4~��0Z]l��_�t�� ͪ�h�$��Y���dB�KX�����	�ʋ�q�OϓE���Y0]o��snl'�_v���;")��d*��o���+:�!ΛP���U���mߨ^ja��������	]�����~Ɂ}5Yݰ+l���~�B/���u�a��J��~p�KL�0�@���� �X�ӹ��@����`�E�65���IJjj_m4�]�ޛi+��ס�`����nׇTy�H��Tc��˳r�_fG<n�'��ғә6A�i2^���s{�G�@�)�������?�����_�Ub9<��x���^g�	�3�G��Z��y���;�9�0��2�oL���t�s`몏�Z�qp�ٹ��7����ryy�	F�Y*D`��W��nF�y�M$�jނ�lu����k0��9\{L�?{F?<!N�3H� ��(2�YD�	�oŀbu+:V��y��D��7����y��F~�G54��'� �7�n.�d�e�g�YU��c��471t��u��`qxw������}�糓���2ag^�6�2��\���f{�Ev2]�9���~�z�)��[��
3ݙsx���Le�Gug�m�wwN
��Vwi#3c�:?�n"��9K<No߾�òq������b-��ۚ�¯�ڝ����7:���f�-� TW��|�׉lVI�~���J���S��0\���8�F)�\�)3����t��gB����rQR�T���?M�E�d����9d\�A���͎��z�90B !�=y�e1�u_7l����
�b{NR�; �@MQP(���N�Ɩ��7�5W���S,|R�� �E���ea2���je ��$��f4$cj,�N�ɢ�\�nv<�XT��{r{�V˞�!`J<)��C��yب�"����~E���&h���Ƭ� B-e� {�ۘW�����W@�W���'�M!:��;��[ `ll��!5���ʖE�17W%�Q�K?I�R��L� ��Qu��@vA\���~?�}Om��醙$y1��� ��N��	Rq�u�eǣ��S�-e]1�;ټV"`�)�r8*L@]�b�<����\��w�x@�<t�6@�pg��h�cs�6��<tQ@�|�߆J�]C��''�SL$��j��9��u���a�X%�̓18�2�ԇO�#^���y�}4��Uˬ$�(
�Ӭ��ܕ���ީ�<��4���ivI�q���,/4u�Zؕ��V~w;_�Q�
�,�o��a�wd�64DH�D�\�Z9��r��ˢ����]��2��6\W��g.���Dt��[%��I��m�♹�������.�D�M]�dc���i`
b�7eK7�D=T��
�Z�V��f�D ��g�J~���Ƭ	���"�*g��np�|8�k�K����e�dâJ��v���1��Qڏԁ��A�nry������zX��F+ٸ��l@&���m�d�E�l�Yja��Jgq��h8�d	괱���?�x*|�(p�G��FbRc�$�-��G���Y)���uS�n�w@9�2�o���+�����+gX��wLt$cJ>����.��6�{a`�vL]rDVw�8#��0�2�e@BVl11�r�R,�h�E�N�˅^T'�2D�"_�T�W�SQ�U��E51{4
����Z_�f���c�X.Ѯm��{�χX<e���� ��9/;�֘���.l�ls.������A(�򨮏���iލ�*�Wѹ�.�5O�VUtc"��0�am�u|nӘP�nr��^LJv<�K/�6jȔkU2�{U�ٌ!�,�F��QZ���T}�ǧ�u������K�٠24R&U����'䀥HR3��7�ڝ߰gJvm;�zA.V�gO��M�~Կpv)�8Ku��X�9�GϏ"6ts���J-L�"qG,P��]��t����78��b�E��l㉊�\fTuv�w����&$�@(^M��ٜؗ\y�n��q��z��?�T��g�"���j�gb7�ɼ��	�bfU4ۖ�O����!n�n���V�c� ��!/�"�
IgfH;I�dpٰBs��ތUBs|8X�z-����)*u�O�~0jw�*����4��3�2���tR�A��ƨ1�Q7�$�;�aсۤŬ[�RY0҆��}͈gƺK����x����،|����i̔uF9��,<C~�
Nlc�/H��r	;z<��vJ1	;~��ǿ���ْ-�9sR��g�|��+P�r�� ���z�4ՠL���4^[�SUْ����h&����aʟ��`Y�
��kYj:=I-�v0,1 YD��8;;���N�=�2��֨�:U��k	�2��9J)%��y� �gS�9�!����g_Y�gHL��&-���}YM�@��R23���}Q������[�y�<��-�:�c�{�>�ޚ=s����[s�Ƴ��?�ט!#�U�^����m��s ��k�@^�����N6r1����v�Ͷ�Ͷ�cSiU#�	�'�z��2:`��6�h�|���x��N�\��2�|���1�A��D���۝֡�92aQ�����lq��Lo�����¦�%\��!i��m����6��#M\gUX�p)��f5}\�|Ý<�Ϳ�M���x���%���sS���ԧ(��P&��Ȳ�$v5�P�@���9�7���-�qf�k�kULܰT'FL�q�hE$z����-	ΤI�(�Y�;�F��s�nsD7�"��A(mRkd��Ki��
������sHR���IJ��c&B���3������k�5l���@�i�R=D�������� EВ������E~a���
�r@��t����4�؜D�f�����؍���/�&.Tᇉ� T��?Q�,vu�C���Z,|�~�i�������hѩ��л�_u�����P���~�4�6Mgø�ȼ�������!%���|!����sb��|T��f*� 0�^|^����9�!��<ϰZ��!�b�_{$�Λ�˹��*�҈jl��=ȮCXs��e�`�)@}ނ��'t�,06������W�M���
���5g)�S��9+r��Ćŀ�<j��yI'�ҩ��cǓ�Ps��)c���?P������ �+�� QˎPgF�6N��N3C�������3m���Ѽz�#�B�n_J�yә5S>�<k�.)�+� s��V=��������� ��߮)�����"��f�$�|��Z:�����u���������6�ʁ;��I0�M�� ]�	�`�>�x1��(E��~������\�*�����LyH`+��f�}�7خ"����ə6�38"N>��������|��Pnonh�F���O�4>6:����5��i
w.��Q#��=O�qS<�ϛ�*�c`��{:��OV�����QYUCA̬�/f�m��odk�B�G1�I����8�v��|�$��L��V%�j������]8�.����hWl�!������G&��˺�����M������dD>L<rV#�W:��I���X���-V$��Q R-C��\/�T�W�4*�����BEgl��C��Ǯ�∇��:Z�Q'��^מ4,�6��̮'�rS������S�=Þ_Jd�"��+,�^�]L��c��vwt��^\�$\��z-Th�܂�{����.]4_w���~����O�qf1|M|pb�,���}�sַ����5�t��mr$�zv����F��
��ki��v�p��M�yއ�9�`��6��dP�����\�����J eG��i7�=DLdg����r;2dv��?���/D����{z��wz��A �'���UdɟS;Ң]���z-��;  ��IDAT�1�7��]m��(R���&���b��c��G�(���7�h�1�`A���͚?� B�U���tr�@H	��,������h�&�P���F8d57 u|�X�/� }��:Q�w
�Яථ���h5�b��)f�P��=��C�s������Y�*j6��k-�ؔN�O���wǍ'f�({�X{0od,��ou�>�]:0�p�� ?�Hד�p�-�.���a�t'�F���9��	,�l���A�H������L<�3��g��U� �^�37[|6	
��� �駟�?��?������_�)��>~�h�4��Q3Hi{�=e0��ή
Y��`���71+�d���.��NV��jl�ŏ?��ϥ���eC`�q��t>0�r"��>Їe�������A��� �
�	�i>����I����ؼ!o�n�!�*�D�i��`#�KKjܣ$Ll6yc�Pa�Y��0,�3U�}Y:�R-Tzj�eo	�����9���=����1��6�2�nen�"��W��K~/��D'N�	�����pU��h�����5��e��cQ��OL��DS��@G$��&�"�]�O�6���4:�QߓD!��ᢨ1qy��*܈�'���4���	���r��mޥX�)'�`@���/�3YM�Yj܃�Ag��9~CL�c+�� ]�׻��Ɯ]���D}P֥�X�g�������������^-m�_�6뻎ǘIv������	�������[a��Z��A]�}	0@߷x|S���M.m>z!���$Pͬ-��Pb H�L�z�{_[�')iy�iS��5��73�>(��e.�a�
xgF�.t��6|$R���l��^���	J�z��ӧW�I:�X�Q��N�X��ײ�>C)�)\�������(��S��U=M{P��<c3������`a�Y�L[���nS�;��͖���lmA�ގR��BYG���KZ$v�LR�'2#�8Ri֔u�[7�wv�0�����naq�jR���0�h���'�T�8�>&�`4Q��_C����|��o�/_���Dw���/�+��?�.�=v��m��ۅ}�c�-tr=ٝdq����w�R��oۅ�oTE�1���˛��7$a	}a$YF�%�gt����A	wr��9
��,�d	��SھR^-�l��d�}��}��%G�*�������;�÷l�_4fN%�1m���u���cp����Ա]G�6���p�#d��5h J\�kIa�H�y�?�ГW�p��:pˢ��,���A�S��ά��A��x|p�{�o�A:����8���4�?�M��F�h%�|��qX�I�3�p>lB]�BJk櫉�����|�.>��G�â�ra��bAG��6Y�s�I�S�I��J%�KG_��� @��F��ǵ���j�~��.�����/��?ӋW?J���ہ7��L��Us���lWm9��ݝ��N�����X���;�>-������CwC!D3N�eL=�-lr��"��1zB`1� �y�CB#�=:��U����w��T����Y��a�Ho�ͦNQ7��l�9��%=$��^��'��+��H�Z��/������_H�-`U�v�^��GJĴ�$"N���ħ��q5�v3��3��?x���!��V}Sf 2��	�=�N�(�s���^���x��2玲��_�d��U�u�{X7i�1f+(� �F܁̐�L����$�^W�)v�a0��n����⪢��H�]l$�ߣ���yk��8����n���{�*T5�f�1(-�a� ��/�����B?��[�L�n�:Q5����ו}T$��S�
��xX�^/����$�������Ŋ��5�#�D�2 �R'���9,m`0)S+ئ��h�2��c<�����"J5�>�6w���Hq��e�}X�����$��P��%���-.g�qq��_�du��_8�/�S%B5<`�2@�e���ܯտ�-j2$PO�:�o�#y�}�>�u5��E�&�ȏ&�آ����,��߬O�w>�j�]��>���=��Àŷ\�l�3�ήY�L�E�׆T��B֣&�7֘
:�f��I>�����t�q,��9�ߜ���˗�Ï?.L�N��n_�ϖ����w��n��#MM��2��\����NRrb��FY;�����),"g�o�`L�:[o\e�4���K��;6��hd7�d���}�	0,��{�w1��>�R���F���)����ԉ��L)�o��b�>~�����g�M ��B_�{��x��Rr����X��`�6VE�{�ۈ	Bq��!���;֍~���/ΤS5Tq�����w�1��ݓl��[����s3V��G�wVE��ӱ����^�u)Ooױ�c�1�� ꋗ?��W��3�?c��Ç��?�Z���;z��ɏ�O)�Y�z+������]*� ��x)̃= �%�f�w���|E)�"ꤍ~�)R�q{��ޒX��-%�	FUa�U{�0��X1"���h#uB+�W�5��6��^���[���'��q���F����ơS.��oi��5>5��9p�6'�=,��,Wҡ�b�(�)0/����t1����_����ckf���B!���ߺ/�Dm��I4�z��D���(L�8�j��Y�*���M��x����0� ��s����,�����P9���� I=�.��ͻ�"��{�û���ﴵ�/�����;1lqC�v���N������~j5~��^X�$"�^��Qny^��ifwS���'������e_$YK�"4�������~����'��r�}aHhu1h�Ƴ,�kC�M��u	k|=>����ȂT�~�Bš�6gr���N��ϟ�
�v�y�;+��VwT��E�j��hUh\�}��9E>�UJ;��� Z7o���LꮔG�h��K���uO%DɬwS����L�\uo�C'9��A�����{:uH��n32&UW9*��z���ؕ�`�>.�ݛ���۷�G�Y�v�;�������lt��`�U �K%R��i�&��0�ْ`��T+����>����Hr���.i�,�D��|Ĺg˹�%�K^q}6X��7�c���:e�
 i*z?�4��Ȝ7\�����IH/�3���b�8�1=��zb��pi��#���|�5���U"3�6�pD��B]��="�X��+�3�P��[��̊���s�P���.���3!&Q���Qk��θ���$
�a��2��J�G{�;���."I�:y z��i5�V�����ҁ�����fgڿ�ce�XYDg4��,�?,�9�b�A���}����k�Hu�qN�
�m�X���p���֮���Ǐz��g ��)�M��/���3�>G���?ο���/��~x�R�wʃ��.u���?Ї�=6�! e7��?Ej��C#�X�q��kw&
�$�tYl�p]�y���H�(�*Dm���|�:Y��6s��%%�g�ZTq=o�-]:��ʙ��@4O�z2\Y[��m8���c�1R K������)�P�_���1�(>�v-%2�h]�^罨�~�(� }���U�it؁^��Z���UN�]�����%��V �YT�X{", z����퍈�B��TR]��e9�[�=�U�5�J����U-��/��Y�|rӺR�;U�y`�1|�W?��~z���a��g�-�[z��+��_�B?/?\�Hr���Qˑ�;ֿ��Oɚ��eX�׫�(�'��zQ���nN(�p`]�K����A���t?R��6���/�	G���Sǚ��~���U����=��&�u�L��u�v;߅�0����U���I��/��`�N/���h��{t���n�������E|�&�ƹ�y��{��7�����
�ƺ�Xh�s/�E�_����O�M�z��=m9Z��ZB7��\���!�e�A�Esf�H�'��G�2ڵ�)��<T���@��\���u�|�:㴀�Ze�O6�I������N��@���y��ai���.u��r(��i7Z�!��g�-����7td_W��m�����u7s@�������&� �rõ��b�A/���!�a]��T���g���=3��Lh�	�4��q�Zv��}%9��0�v�R��Z��'��7��jx@�6�H]��F��1�kӛO"�P��o�H�:��u�ܧ:霸?4�ʈz�`�M�s�l|8ung��8��4ي����Eey��F�⯃U�F#��HW���j9eu�귱�[*�h#i����3?�S��u�D�QU��}GI$n��Uo*�_vYj��Y�iv��JF�=w��٘�(�L*��o/'^a���.�xU�����إ����
��`50{m��z%l�:U6)�N��j�D>�*6�`��T�[��Zt�@�o	��L�y�g�/iiڛ���Ԕ/>L�_Ʒ�a�i e	PͲp7���%n��Sc����<�q]@-&�z�� �o�
��+t�-1�W��@����@��XX̲$z�-�R�I�3�l��<!�I=)��m4�X�K.�����%�)f��%���ɶ����lm�Z����ŪX�}��!>�rC31/�]�� �g/ ��*Vt����V]��E���`_v�Z�^���}���C
;QhRI��4!K_�zo�������o^����&�/��-�����}����ꕰQ6��'��U�^���,��%�����$�AZ�=��!�K��ʄ@�c����e���ӉQ78��y���#"����A�w��g8g,�|ӹ��h]3#s��a�7�kWT��#��0��yH��IZf^�6��n4�Q��ҵ���dH�5�%K�T+-�PgMO'�+�qJʻ�T�mqT����1%+�b4��|��.�-aխ�m�$��?���o�cf�_~�E�0�����3���K=d�Jyd�w1�a�N���]9Xa���o	�.�n����g�x��J�m.9��\T�)	.�p<����^k�����"�Y������������ͭ�g�A�̏�h	T&�aK��K�,i��/�$�"r=��%�+�yJ$���2���!����1w��ԡ��^���S��8a���I�M��X�%�紞t���
p�Sm�+ �n���OQC�13s�������|V�f�'\�>-?�0�i�k~������O?���L'�dP�2s;j�T1@�������M�,��0sk�a:�����~_�ux����$ᓤy4y�;�D�ɢn`�_�Z\I�9����̐���׀R0��l��f�a�h�݆u�U�`��%����͎�E�X�+����N����<�N����n���"�k�o
�l�������K�������"��⸿���/��˦�x�Qc{x
��4ӽT@�͌�%�*�p��ټ��	\�YB��϶l����A*kACN����
lkv�c�LMf�g.��>z�ӥ�V�R=��ڤ1j�1�g�ʹ�{�R_�����uy�N�?� Y�G���_�C�:̯�e��'n#؝[�������
�k����ʜ����Ή6�m}\������H$Bf��Y��r'GՑ�c�xf�9K;�/׭|�#�!�[�^t��Ã��3����v��;w�ADg��E�?d�� Ơ>�Z���4��ncm�R*�f�|F*���	�g�LH�\a��W��N�$�f�E�,�|�*����|��#? ���@����~�о�����3�m�;�&����h���A����l����5s�	���^,��$3K_�����X��ŋ�!�a�G����� ���k��/�htZ =*���d����x%{3nV}�{(�rf����,�'�����Pf��}M���z��G���Z�G�D��Z�7Y�[;�S��݁?-���� ���Tr������ >g_��uܓ��U+O.W3��6�c�5FJH�p֮[�;D��?\�PK��N�U���a߀�Bq� |i҃b�{��ݹ��W0�>��R��u��[t��G�~�eb�Qc��	�g�"O���OT]"��u������(�L��לQ���<O�1����F3Rx���	�E�.�l��p61���l��,Ϊ���Htas��յgn��y[0���~|�ra�7bH�<�&*`q�Bl�)+~Z�]9�M�����x4-`��r,?�K;-����a����A,9�y= T$+��^6�ya�}BI���s�����d�X�ᨎ���EQֻI�թk��Ŝ�E����R��:�������r�J/*�	�,nw����uM$��s$#��b��{��(#���әK��O��~�̕>�W���t���*ْ?��1a�4�qC�}~�Bexb��9Wԡ�Owܙ�<�X�EK�^Q�"��(6W���Hì��󶋲RK��'
J�^7�ךg8��kdng B�9>�����T��EX����%��+}`�[�$;�W�ɺ٪.��C�F�A7@���Tːp;�Z��������0�0����D)�(��R��2l!{;�Ja�8�s}����̢�Yg����E��\r7��X�$B��a�Kx\��8��r?��A�'�>M����{��n ������Tn�\a{v�ɒA����H)8����q�.z{+Ǽ
���J�sF�D|ͱ�ޟ�]���c�3������=q�����2���Ó��q�j|<��4DTm��qmͩl�vY�ۦ[0/pI?g���j�?����P���ލ̊�`�`q5�N�ͭ���C�P����Z���t�I�?OC���g{c�0���w�_���۷�����>g�bc��t�d�5y����S��{jv�W�u���7���\��o��￳�� ��L��4j�>�;�/���4'K�̌Y�Q�$�nj�3�dvX�{��ӼF.e���a��y�d�=a�v/��(�f�r��]��1�:�N��_��� 5�'�4W��T�r�6}F��(����`�U��yR=���${�l�C72�O�??����.��e�'�
�-��M5��(k�K��U[���ナ�K���Tn��1ES�9wf��r�ׯ_�o�={���$`���+r��{	�/�6)��M���N�����?K�(����L߾}Co߼�2)�3J=�(�nn&"[�@3��T)�E���Y�1z���m��=W�[�^Kd ��@s�=t���Hɧ�X�}�`sQƖ3u����Uu��й]b���n ;{�r�+����W�~uP�S Uu�%��I��'˖��?}�׀��س�n�%r���%y10k<�iY�d�-щ���r�[�͵����{��[�p����3��I-��*c>���|�������X����c�z��-������/��ka˓뢊e/i�J���o.Ë߾yK���?���N2N��?W�����`�ZQ�e`��S��bs�u9�)����wz��K9_\θ��l�|9��:�[�>�b�$ђ�(`�[xC�T#�jUDo$�JuF�8��k���G��p�S��L����F)q�1Cc6Ja^�iJ1���\#=����Çq�z�����^���r��j)��!EOs���g�q�����K���h3Y�Љ�_f�r�P;BG��)�2�
S�O��;>E�2��5Q�9�8���_n�s���3sb��W|)�k��b�}�å��`]��IJ4QI��L�p�����޾}G�?��$��,�`�����x��Փ1V�C��ϹPQ����������"���0�����=�%�t�����GN�'b��������n�Z[��϶�h[*�5�2�@�sO+}b�0�f+9PA�~�z?�:�rξ�N�`��<hU+�Y-��2y��O��IU���XDV.Q90�먏Ɯ=F�&��w��Կg�����|{�ABa�#:���B����O֡Q�����B�M��������sV�i 3���a���\i%JX����g����Pa�қE�eQ�l:c���Yٷ��@��,�KUؙ <��G�����TU7#Ts}/Xi�zl��x�)��$L��y�LA�c�=�75�����m�ע�e�0ڽC�hφ*n����񱱠Tv7���X��oLdb|�R<bh[>�]��>a�$�I����l�ɇlBEY��)
�����/�Qr��,f�3ʦ��JV�6~�o碠�Yl��RhC�����QNfN߄�Q曟s��>Ѿr�w1AO����O]Ӟ���t�&�k9��ܥ��
���8�/���-i���k0���j�rf
�vR�7iȺ��=ji�ٮ��T�c6�믿��k6gIz��6��ɽ� ��4x���쁪`40�I����-l�/�?����K�Ø���~��>�ua�N�,��j�%_�#���7��]���h�Qo�YQ>�f��}N����2T��k)+�^X�d�@�Ռ�Q��j1B��L\�,�ڴ	�%&�����Uy�j��~�L�":�In�6-�cH)ARV�lPxY, ��s���Fj@�w��f'��򳡳�w��wd)���}�����L�ͩ:�|��x��O�2��d��ku�_�=�_I?�b�:�SP����s���>���P�x�Jl����q�Ȑ�&�9Z�Hܧ��0A�hm�M��)Q-��.V����ۖ�.5:����q���'Θ%���Z4�h>�
�R�u�G'q�7�ԃ���8�:��S.o"%��/r��^Q�����hY��۱�b��i.�acU�,W|����]� k��ހ#���0vnR����b�o�H�ctPu�V��6�K��'<2N�I��4g`�~�zq�]���9#�qH$@횈�{;ʥ���gx���]f�eP��u�r��N9́8|�1�Z+�~������zȴY ��j��&sC���32H%}.Gѐ�w;S�ӽ\�`~���=�u���Qf�a �f�������f�����FJ�����A�\~�H4ł&&���8��fY�A��E��I�|����8_��]�
�^PH3���ndH�Dv�&Uu�j`����7+V����_�=�V��+~���\�["�����#��:O�U-�q5A��u�llj�pi�r����z�ێ�R�v�pr+P��Ƥ�a�t���8��� ���>��h��x�l�*�{�|��u�Ϯg��.�P?u�n1:r`���ȹ���D��o���;���
@��#?"_��8�]�ɝ�'�	��C��AFM`\��� �=�wM����
*���O��f\3��,�}4�1����r��H/��7��x�#n�'�(�Ժ�y�PK�(`��A]�` c�Ȁ5Ih�$?��@�N������obo1F�?���r�j���[���-V�Hf�"Sw+Y�Vtn˯��|�&��fŒ2p����\�e#�}LC�ס���Q =��� 2�VuG�{ݯ	���/��,*�{Pݱ��u�d�4�v�@�����}��ga��-�`���Q�ZA8m*ד���P����;ϰ���x2���ԯKyt���LCN��3��+�3�c��� qy&��
c��KX�ԅ�9�c1V�(�^���t��#�]4E?�Ə�f��_eD,i\9�٠_;J6�f@��i�)oV�ْ�0��uH�
�J>��w_MSW}u�lX w�g�SRNS�V�
T��a��`ѕ|��V7�Y2��e���Z\����G73�f�O���	�gҙR�T:ݔ,ξ�{.�ۃ�yJ<�5%J^2��̱�#���.�#�fdӭ�i����O?����<�-��=0��)���5���wǺT�5��_�����lLZ���L2�yR����4��󎧏�wq��S�IT�@�IYR��9�2�_`�1���c�P�.J �N�v�Gݤ{�v@'�N��^?��=#����ǺV�e'�ɬi3����1=��Є�8��c@|%�
�W
�qi���ZMdA���`�q� ���&�*����X����Ⲇ��ߩ��=��DYч02��F�l��2�-Z��P��H�y7�Y��� �32�g��bQ��u�7�к��>zUU��ꀍ}��S� � �9����W�/��H�GRBہ,*�J�E�9kRdۘ�*���.�<��~c�Y�\��x_�|A�����^RQ�i%�<o!g�O�K	�����G����>1*��}��(k]r���>ڹnkGM.9�Y���6>��&"��T���uTRjg�S�;�������>>�k�T{�_���P!@�(��.��	����T1qb ��H�`��`�&]�<����}�>U�?�7���~LBWg�G����h4���~f��U�w�R�s�GQ��~����,P:�6c�_A�\���>G{z�'%7�eB���r�J:���7RD�U��VM'��
���u@��u��N�d�P��3�U�~v�7��J�/��l���3f��Iz�㉜]^��N�?�29
�?��ӟ�f�3�����=��SW��b"��}�I�ɔ,Z�~r��	s�u��`Qg���5�uDu��#��K�ʧ��KٖK
��q��,5�zc�1V�bg��@i��1rhC��	E�YcsDJ:QUxi&&V���䉶E��ZqcS�a�~�MR�'a逃�"�:���q��{H�7��؞�@U����P'��M#"���)Ƴ��@�C4�Y�]�$�?��ru�[M=�H�in�}������[�di|�j�⨂������y�߯�Ǐ��PO^؟��_u�X��=X�EsN�����"N�V�����Qt1.̏��f=���G�ߧ<��2/�Y�It���>1d�	9ky~�P�"`(���rR��st=��� ���	�ì�>��iP%Wqh&��9�e��1���� ��@��W�
Ʒ�����"�A���V+��J���0ZIy#K}B�|���jE֫�U`�`��r͂�����Ү��()�@\��6m���Z�+�]����ck������b����.N�Ǉ�o�/l�WO��������εU��=9�|�~�ޕD�p#á�5)��gK� Y���6�e���Ա�H�<���}��>�S=��jē�9���J������:�&���ۄN��a
�����Uݨ��Z�?|�����J��p��F�9nY�� *3�唽��-B����������b�c܂E����Zϻ�`�FF+���|r��ì����c�4?�,8aw5*oJ6�Deqa�mf!)�{2}���l0fjnT����O\��A)޿�:��CM@
p���y*��MJ}P\nW3%�g�������(�P`u�D'�W\��틸���>D��}q���fBz��,��U4�����L&��Wύ-=�bd\4�ڨ�z���ٓ��)��鬟�l;�5��fFn�C%�dȚ�}h��Ǵ����^�Y%J��ל�폢ED�G�ݭp_���ђΐ�+!���e����v�����*k� �kx�H	�5�v&�Ƙ�����7�fٖ߳I��c�Y��-Ue���"ϭE}yt�%i�"�+ï/b�_A�x�8���~��.�Pb�W����(�n��t}��>u��K��|�B�c}����x�/�����k�|wV@�o.�Y�	p��Յ,�B�2���,�0�M�ϲ����A��w��ʠpX��^͢�*ڧ�;��!�T�E���'���Kx��Ef�&nw�( Gv��d~��(��+v�}*[����b�J�=)�P�5��iL����������)�@Zn}`���^d~����Y��D��v���j
�t�S�<�^,?�3�����p5CʛO �݁���P�4D&=���5g��3��}��ƀ`���w���/��ң�vح�-$� ՏQ���~�*�av$1]�Zq ��E t�ł��r������m#Gͭ���,T�OV��b`Y,� �Z`j���~���;�p�I7�'zţ��2k�U ���-�D��-���I�zo�*�I�>�ǫ�כ|㾼�������:ՓOqL~x%�c��U���c
��_�Ṯ��'p8n�A�>��r��%�}��M%�;aϫ��{a��7f��r�e��j�z�p�n�e ]�G�t[O|Ĥt!D`�x����hCAu:�;�`���5���L)g��E�ʐPC��7*��^/c��5@��9E^u^��SO
��0��ȹ~��V��&>f
p͇I�=�Y3E15��A* �½�Ĺ]X�����ˋLu�?x��V�w�`�G�戅^qARg�5pe���Nic�)�ЌY|
�Ւ�=��z�|�a�@�Il-ᓯ�USӃ^��>�*u���@z��������*�"����~x��;��s�aB~�~��PĞ�ͦ�zT묊��NM ) ̟U�%`5nXkZ��b1.�Y ��tw��'� 	�:�r4 v�YB�57���-RI�6������h��[�� ��O�r���N�� �`��R�����>O@����s�bUC�%�u���3 ���D���#��x��?R�@YM�yN%�*���<I�׻w��Cl��Gv�-0�=�[Hx#��~��4��������J`�'$ ���u�o����!Ɇ��?��a�<���|?���eӗ�N��~��s��X���?n���}�0��߫��I�Y�a�
�!X��ܱ_�������	o"JO�@]�LV�Bd� �q��u�7YL��P�ذ��?�����|�H�Y9GE�":b�^nû�k�D~A�c�tw}���=��*L��K��u�T��栏sX'���\�K<,�Cƨ@j�C��Kw-'��u��ߎY�&+���v^���񍒣�G��񱮇?�/۾�X��L0q��MpzI_�F������ǧ�� �:�c,��,4c��1*��g�]f�7<�X��Lf�𧫓e���ȯ�DZ㪻�
��,2�����ߟA�"ƭEyLm1�3#t�t���%g�'b�;T�4;QS���U����m9���bO*1M�|�}ڪ���_�|z��+��G��yXj���*�-'�L)MXa��Fɓ� ���eSDj�;"�-�����]�D��f���-��2��2���ܩґ�蒬�h�.}�X�1��;~ן�>��P׺'w��NnL	��z��ĳ>B�+[�VF�փU95������������ɏw����%2���㰹�;�?,�$(��%�>��zS�(��"��ja�E�+�v4�����P�6+�B͢�����bg�h7c��;d���c�
:�4�<ߦ�9�YP��3�Vu%��9�S��&�ɲX�վ��α%C����#AT�=k���۲��NR��X��,�ME��nj�R�h/ύ��60��/b���Ħ�����̲�H�,�l��n�~;rV�㞞��ԅ�a��.XE��J	�)���@�}x�3�����y���SqY�]��I��: �q�ń�[s�o�q�z�@����m}<�� �ݖ0�N=|3��Rz/]<�$Q�fYTY�k�%2�%���_����wfӗ ��t����C�U<�=��t�A��ňK���#�.@����PEN)���A���2����	�݀(w��=* ���0�y�h�R��Y�T�:U�)�S�V;���Р9ϯ�G4�1�i���|R�����o7-��T�!�����qb�c�����
_H�C~U��x83MBd79�����2��v�5e��)���_��K�)��)��.ǧ?2I�G�p2%q�0�Q�����KWL��)R>Te���],L7�2����h�}B�}�s�R�Y��/�5�����;a#�F�r��W�~�ϑ|��y��+��n�?U؆�]|�?��A�&�\�S֕�~������TA�vY�p�W��)e[+9� �s&j� @D��{L$�/i�����κ��	*��k���'��w6�8W�|�K&��3#�AW�k!q �^���9a
@�L�ik�r�`� B���|��\�w�߸��k�R.�Tӳ����7+��d�Ғߞ����A���Zr;9�h���#K?��y�L�W9�����t�H[隭��'����Ӑt�,`������tE�&��r	g>�ml,ᆜ�����������ʖԽV��r�n���DO���K��e?���i����}RmF�Ҟ�K'�F���CP?�Ey�h-n��1!�?D��?9�������f񎯉�P$��{r���@�[� �#z�e3q�#$^.�H%��qO=mPWy��O�ِq��7�,z#�s���L�� }7��6.�O��);����'V��g��ʫ�� �Q_�M� ��퀚k�b���E.���)�?P!�gQ%H٫$Ο ���=��Ņ� |����3�+��`2�`@����nv7����?泻{�-ٗ� �9�ɘ'e�*�O�!5��ds1#R�T܆�`X�X�\0-eP�!�z�v㌩��'�����T��i�(�i��4]i�H�LdN`{DTs�I`�Q#��<�H1@�O.�X�o�6�:$�i��4} b$&�~����K�G��e+:��̐G˴U'O,���"ѓ�-�%�bc���������BfQ?�@�-]��f�1��zljP��Y��!�^���:��'2T:�x=���|J��� <�n0�̷͵���c���b:���ݭ���ͭ2�4D��P��O)��"e�Q�2����8]>��m����fúZ�[6�-����=Gˈh�9��O=r�"��(��K̟g�	���( �^'m|%]�D���q�H&�~�̾�l�r���Xn���z�R|�������4��>6�}��*i�J�!���ƚ��D-3i�1]�Ly��d�X����:�<.=��ke�`Hk	�\�������z��+߮L��4j0�/���D�Kb��"�0�>��������a:����F��|�v���$�8�s�Q5���
r[K?ǌ����#(���Iۻ���s����gi��Ǌd%��Qe��
�ie:Q����L���D���e��dA�i״�����f�� ��f�k�N�_�~�>�5K�޺m`O�D����w��6�� N6W9P �&�sT�Q	�-�_���9�M�1�(��\�NTF0<{�c ��&RN���Zǟ�P�� ��.��b~O]����O�:fz��s´�t��Nf�� u�g�5(�� ���%�6�* 'T��1�.���{z��%�x�B���۬�*߱(�.դ�Ia��[�QwWf�q�}�O^�C#�u<���	w���+N9�Y��>���'jy��$�4��\��x��}.IOˇF��m@5%�FI2�[��(��"�5F����=U�z�0t�14,�á!}x�Fi������y�?Pa�]������l�����E�(I�z4/�񗎳���I�侜v�f��]Zl�OЫ%#)����r>�P�HXd�
823�������_~@��!XX��#Bҧ�s�:B �t�u�٠�li:6i|C�j �BD^��G�y�\��w���&�ɯo�i�V�j`��$+th�;���5Oi^]����GiCT���}�}�T�(���[�|^<'k\��7��7"OQ�G=��p����Kj��Բ����d��P������b\�x��D�q9�%���<������/}>(�NJ��8ß?�>���]�R���d-�.=h�V�dCP��L��X�>J<�֕Oo߾���rʌ���	��/���T��fʠ	�������s�����+b�a5�j%���SN�~vm8���yx�+j� 0�<?
%��&���\	_ݒ��/ �Y��Ӹ[���.~��������W��@PdD��"�Tζ�4o:��S���oQ����-x~��y�+��XU?�or�6��G:<I
��'�Kˀ�s�J�� jZ@�[��2����y'�vY����6�˄�1�cя��iN�j�l��[;av X�-�F��zo�p�8�c���$'��o߼�)�΋+��hb����={�̷zL6�I�j�h�:K�;�뽥#���� 9��p���}/� �;N�fϤ��0̶�'�f��:�,q�Ci��+�5��l,~2p�� �D!��}-5uX��[�ꮝ,�b��,���K0>�M��&Y�w�A|�%��vc:�4璔��nH@c��^������؋��F�{�=�̇�)��J͛��
��D��tu8+o=e��������ǏO�����r�S-,�`'�]7��y�V�m{�PY��G-Aͯ�����8o�1&0�$N�?���D���S�zޏQ���T�ZB�����z�����>pdmy3�s�[��"|	 ����	,�`[�D����Q�p�XSZ�k�I�=U]�ⷼo��1^���I� 0�<,磦d,�e%�՟5����43t����q�?@������ۖ/�S_��9�o��#�/��`�l���"�3��z,F�.g��Ey�}^<>L��޳͑Y2I�i�[-3ұ�ew���ؽs�<�̌F-��wUE2�x�!���"�� ��L�D^��J���l�L:�q�_�✮:�b�ȓ���$��"8gbg  ��=�'�E� ���<��>w������������ᄵ��#'~QΕ�}3�ɻ��5��
(�2w�=)��A$Gv]�̚.j�@��*I�U��w,!��Z�w��s�-�Uﾞ�L�o����q�u�?��Y#Q½�ſ�&u�m� �t��̂%?�ڀt�6l��QL�Kb�닚V,�w6®i����f�-��\��ȋ^v]�����W�U�������[�k��>�]�����?���]�K�G�\���8�D��s�e ��ǥ��f/���HX%�O�
����-$���&G�A)���e�R��ԇ���D��h$*]\8��+N3$�L��'�7�N��H6�E�]%v�.u��x�;��n�[P�~��B �/�N�e�ҿ��V�ڕuV�O�d/;�[��֠��X����=pܾ�:u�⅍��j��q��q�>��`��Vt�׳�[��zz�Jm?�,V�K;:��%8�;�� �������]����S@-��ۘFX�3ڸ�_��X���q1Jm֯ў����!�\�ջD�z��G�T�<����:�Z�iT�&1��-4���%��ZJ	g�+,.K�yU�?��E���G�E�:���&�7/����5CN"FQ��܉vq�if|o���>/
�p�~dR�q��Vz��DK�?�zgl�� /:Y_�[���������/�t�z\������ҋα�?��	�L��Qv�>�۔���i�������Ƌ$�7��m�i�K��Ns!h)J�c�Q�p�������q
���_ �PL$y����&-��G#i���W��-�F�j{?��J%��%jKh�[OW��g��*�E��1�W=��Y^Ċ�I�/Z_W�S?����z_�zY|��MTc�-��.ʨca�vD��4բ�}������}�~r�a��;�Kj����(h>E�"��l�zS'��<����P�rM8���]�b��M�d�*U�\�D�*qS�ʥ`��a*r�e,z��_�
���� `���j�(y��S�C,�~V���!V�-�B�\�1��'si������z_w΀U��X[O��\my6���>йsF�a�U��w��@exA)�3m�R��g�/��rS���.e���0���V۽��ۦ"o%��ߪSu�J9,��s�������i�ZOt��;ʭ��u�'�R8Eٳ�>��5�T"��}���ߜ(�D�$ǝP���� }8����p�ݟ��[�Oo%�fx�-��9 ��흹M�a� ��yi���7�C���h�1����u���Rur����z&�X�Y"򤠴���"V8���)w���z%�����G�k�)Z����H|�V�}�0D�\{�Y�r��6�Bm4&~ѿ9՚:3&8e��l�`�3x�4S�ip�XK#��������p�~���K�W���_r���&� �:kgƭz]���xB��A4�Ȫ����U�N��p3���	E�rS�$=��~�C��ȸ�q�t�
�����_�o� ʡ�s�h��R4O�ў{�:p��T/�:�LP��V�<�z�Z��uJ��_G��K�c�0ձ�Eu���1Pm�G���M����ZZ�͋����=�?��~~3jE�:W�z_O��8��(3zy�+W���6
���	��h �sp�s	�d���DeM\&J����<$�|g�d(�>�FX��<�Ӊ%�N]o�w�m��f s��:�Ps�)H)�Tq�|���nLT'2f�w��Ond"q!����n��͸��ӳ��V`n
\zlR&��Ts��gi��+���VM@���uۖ�Z�Mp�Z��Ӊ�5|=�{k���jYNwv������"��r�_�+��U�➰Sn���wܙc�9��<ƙ�59� ��Lq8���KE�ѿf���b�4��^D����'����
.O�b�\V,�>�t����@R0h�����i����6ս<�"+���[������J�eMhb�":U�T��"doL��hA����@+<z@u҆�[lwIeT��S��[o���J0���/OM��?�#�"u��(\�tT��t�oM�7���_�E�^++��;mQ�� �s=�;��>'�mb$3cA�m����D�+q�Π4d3�/�0�h��0�>4T�nT��.�I�'�:(@��iP)	H�q����b@F���N�����њPK<���ɽ('�,W(�z�=O��u��nME�E�?v���*P�s��U�����DI��!�h�Aoam(���؊�1����Ƥ{�ܻ/G�@
��Sq�aw��M���)b�r&�	���K�'0����|�5�D��r�JP'v�&�'ɍʾ�|����oI�V&8�Q�S������Mp�Y��8��{0���b�n��(D'���,���C_*˾�J�(`�8�)�q)I��=}\��$�	:QB~�W�a�����u��c}�@��?����-:'��z/�T���N�o��~5<��Ӎ+Cڗ֔��K�޽2� k���LԸq;m�V��6ʗ����i�!}A�-�+���$�L�_"j*�ᷖ�hE�F5�����0iZ��x�z.�����e7�h�smk�G%"%���DMB��X�P�zhxQ=()%P��-.:�yQ.��S�#�	�:��*o�g��U�n�X�t����a|QA$HZ�f3� �"h���X4��Z����9��U���T$Ne�_T�K!�������Չ�&�s�ٽCu�V uпX�D{�U��X�ݤ ��D^JvD�MS	(�8D��w���;7����m0��+��I�o�&��Q;��Q!��DܥZ�䯓���$���"���4$Q�%a�#y�s�8M�K�!�Mg��	dLyB���O��HyF�+���u�<Ȟ1�1�k�~�g��4��g�"��m�]A>��:��^��q�~�7��n7�� �w}eѾ3���vY��;\ >2,��'U�� �_hfuA�k;å=��zC>���S_�Z�V6ǉ�c���
=��&��F*0Ÿ��;h[T��������_�!�"o�P�_���JD�]��BpǺN@'�}��
�ׯ���n��DW��/�X���B#q"�B3�}��?G�ڵ��9��T�e�R�T"�d����u�yQ(����N��Lf�D��M�[P�Go9�Ǯ�,��y��z�t^�ό)=F�Q��x_u��w�sc��E���r̀C�k7�L�~=G��Eْ�m�y ���|��]%e4�w_UHm*ѫ/5O����_�2�9���s\1H���4��|>%Z<e���ʸ�wk'�иN5���<�4"Q���[ؘ�ݺ�o�W�ǝm�rV�}z-�n�U���+[�s>�>����:Z��x���n1B�<��'�8�9�\"���
��&��V1@�����H����U��fl�EU���GV�c�(k�?$ջ���|=X
���B�p��q]$�kt\��r����\��9�
!6�X���<���N�r�|Ba4�++�Ή�'%
J&�iBK��%�
��\/��\
�k�Sq�#��ƁXgpE�n��h��c�]*����z�7�y��#�h�7P;��[�So�Ͼ�_�ѻen?����a�x*��~�ƺ'#t�oԘ���[�{}"�aQޥx����ʠ-׈�6S�X����}�f��>圱���>n��0녥�o�xT�����Bsծ�������|yR������~z}�X���X=h%�����VI,�>�y�t��uy�xޛn�m߱_���5w9¬z��y�q�	56����'h0���)���Aa�C�bs�j�e�l���Z�]H"�&�b\�ߏE����?
#+|ӏV�~9�;�D�(�4u�y �(���>8(���cܮ\IQ_��.�'F��N�U-
�׫A_�jI_�UY:y2�49P�g�ݴ�t����q��(�Z��B�[l���=�3`��dȡ�}��@0�l��C�?���*���g@)�`;�a���y�FN���C1)��I���Kt��H�Ro�0�S�U��+���)=p���{,�g�\]�~�
h��9����2���{�_���c��\h�d�L�\��v��<YsA�����M�Q��:_��x�P��ʝ����{�ש�C�����(x�?=��bR��	��}����z���>�~0E��P�Ϳt�fzbԕ����Qm�$��[]�ĭr_}ł{ZG�<󹨻̉j�$�����H�7�3��� 5�R#,�{V#�i����J�^�6�����W�icE�z�� 1�!q�o�B�^$֖<��I){��V�PD�N��"\�-ѾxP�3��To�i�%zXyVG������x˻�r��w^�wᐼ���'�6�>
���獄���b��T�aS1	qp�O�>[����a�U�:���X^ZF���ڇPQ_�[���j�&挋<g?�&'8�
0nR]���ל��x,�CUˮ��װ��� 1����µ�oiI�7��j��⣣*�q�3�ܵu����`�?��;���2���W�S���|��,�o�8����&��=X���sDs��#���{��\�?�QsǺ�"V(2��PD���q�ol��c�r6��=��:��Y_:�G<P�\�n���cl�*��)v�q�2Tв�)���nK���Ձ�X��~�w�U�vܔs��v�=i�����&&�^�1�_jϳ���:��E~�w1:y]���/nb6�(\M�5�f!9ໜ��e0P��5v\�;_#���\�x�ۦ,>�->ɭ�Q��ɺ��No����8�z��_�x��ED]�F�R:�=\5q��SZ�ܫ'�@4w�W}_%!Uꌾ�?�g�@�cǈ�5@â�]��}��a"vD.���K>R�wYO��~��\����2��=6�M�fJĝs�F+�ôfQg�7��֡�R�$moM�s���{�RFn:��l����ܘڭ�����{�����q;n���I�]�ʥ�d��]W���=�����~Vå-�3ʵ!��yu�>[5��0�	v�[}_�mu��s�x�:�/�C׺V�(J�ߏ1�[��7<@e1���k��F�;j���m��LK"�Ƞ�-Ke�{��f����S��'\�����z���ޙ^X�L5NA\E�z�5�}lJ�6Od��r(��@������+8!�{ml�8c�(H��8����_ O;vd[��,)Lk�;�rO��]�7U�v�g�y��S�=��*ef���5��
�j��,�I�RF�F����.����>���`��uG�|@ã�s7��[j
��=�O(�H9�d�(���LF�lb�Q-\n��ZVޗ�("`�~i�Ȋ~��9qi�N��r��HPcq�n�K	dK�"�����i�lJn�Vg�^�R%�W�N=qL��\����J$-�}��T���+�@�^��6�
��g��~�A�Qш�����n�x�^ߓ#��� ��62N~��CV�K��$\�hW��1��O]��O���Cd���G���?W۝��)��c£�+G�^�����!ۃ3nU��>�pD�k�oĤ�ͬ�:a5щ��:�a�i���'�f�׺O��[T�v+�Sݩ����g�K����g�!/�WV+<�ܟ{V�w�I�^��1��\��>8���q���]�k��9W@\_�䡭�N�n$5��B���.^����Nr �A	e�g*}���F�J��]����$ب�0b�҇�Q�^�;��0u(y}^E���gLWm�E�*�V�7#�#�d���wд$0ׅj�� ����kq�M�POp�	ݜV���1^����-���fQ�$�8��z:;#"����9BӃ��=,��(c�ǡj�޹d�tPW���s��JU��$�6N5j�¥֎���E�MR�M�����WO�����W)-����6w]c��T+�[����|M?'B�Y���ÍYo��`C�5�Y�Tʋ��]L�0P�����wb%0�J�[��s��E��L�}���>����W���@�h[K�i
b+���x����	�g�	��K�;
f��8���t����m�(مl�4����"WO�Qܘ8��a�d�v�B�1��+�!CD�L��} <������τ�x-�>�d���R�����{Ml�W��ӡ�g1=�{w�mS�t?�e�Ux|���V$'87Y.4�m�6�a�����z���"Z`�>��S �R��R�ґ�LTeP'?Arm�^��,�v(!t����*s���=K�0���Đ�MJ�%
`�Z%a�u3V�k�S�{s%\���]=�Ym;���R�59DF��/�B0��T���&�M:�t�^'���^J]����&��R�_�O�
 .�iee��K%�q(�G�=?��)�y8��'�Ƨ��ކ��^�w�X3(���C�Gm$M_�XAUK{p�o\�ܫ�O���!�M�n ^��F떄��2��-[6�Q߱���<����2Imژv����y���7�}�Ǹ�Ҕ\l EY�C�P�"�Ƴ����쯡��ٲ)��Dّ�R�vږ 5Y�G4�"��_l�q��p�DG{'�_d1��}���}�b�P���8m�|4ݿ�~�:�]�0[z8�6��݄�y��Mx��yx�����ٔt�L�黯moc�j)��JvPu%���J����)��)�6Nʪ���9�}hT8�{�Wذm��q�x�҉�v���0dc�\S=f*�8q�c�X���a??��4l�l*��ծ�PO�|\kۗض���W�X�vPrd$N�k�)u�)��� ��P�b�D3p�	��+��c)Is��T�^���$z˻���E��4V�^��/���tvp��{������ɓp������c�Pg�=�J����.RK���r���j{���Kq�%,t�Q�u�k�6&��-`귝P��j���z7�aj#�[�S/�6E��/<Ź]�C����a�o~ʴ��mz[Á���i�ѡ�D�.A]� �Zܹr��$�-�]K��DK��Gp~r\���N�X�@&1,��B���4�r,r�"g��&���L�	N�DS��'>A�����w�����>Ϟ=#МH)5<�=+@5(PV�����	�U#N�.ba�L���u�d�{�3���f*���|J�|��uZ_?Z�xA�EPF��1@�wN��ΥT���')��n"�[?F~��VO�s���Y��LT���
� �tR��O~5L��&%�y�((-�.�l����r17��Jd�L݇*rr�{�y])1lr/�{1��||�rI��0 � �s�&�2�x�X�g[p��H�K���,��tt�^�f0($3��S��WN���-7�r1�� ��~���K���c��`"�f7ٌ�-�����n
��O��w��HZ���{DK�S�0�/��ө"N�.��Ż�Ho���m�.է��:0��P>g۲��P�@��7o�Pyߣ����[�{�9�Y�~d� �/ `��O,�(�a��T1�?�s��	D���\v��ŀ����P�@ݢ��s�|MO��e ^Ȣ�����/��W����}�ƥ˗��T�?�T��fL��|Oť:��8[��<��Mu�i�N�F<�d,���6}>~}�6F���>��:)P(��Ѹ40ũ�Ե�~�c�gj�?}�Xۮc
�%�!�-��f@=��������ի�>o��{�><��|���'�C�N��?����9��* V{��uˮ�P�oh�,�ͪ�;�cݵH�V��Vr�p��KZ��6���H�D�|�F�_�N}�޽s'\�v��O�U9oT�i$�2P�(I��J����6k�quzJ����,mد��s肴ɳ]�f�p#�Y%)���w����w�~���-�z!���<"�h����q�4�T�����})\��c���L� l1�0��\��,�{�.���?���>��dN�$s� �y�����h<g��A���|S�#�d۬���tF}�cُT�9��9L<��o4��0��c��$���0�!�Sz��S�����xx���1V_�u�v���[��J �V���"��N�2��e�z�Ę6���Ʒ�,M��!���q��҆����Z������sz5m�V[�.U���D~mc��9D�3[L-k�_�n�ʯ��J��? 'X��"uppnݾC�I-����(�������l5��@k�Ne%b`N��Z����q���RUjıP6)�@g����q�網��@�ntJ`�J+��^�.]�k��V�$-�>밚.XU�t��O�d<Ne��m��]����:��m5n3�e���Q���T��71sݦ�H��@��t���1;�b����ߟ|��o�mPe��U��p�3�v��Eڅ�0�t}&�%��/&��s���Ws�W���v��k(w��}�Κ;�{����T�!�S� LM���{G�c������%�B�~���\�?'Q���DU��Y���S�sV��V7�69�\{6�O�����6c��S��O�vw�=b`�T�F�o_��]�F5���b�&7�I�g�����m/j��Z����.\�@���ǧ'=)�V�:[�= ���NA�sM!)��+��@f�|�#�t�$)�8��Փ׫�hsÃqˢ�ŧ�`�w���\�����Xv�RW,��� �����sp��e*�gN/�L�fT]��(?]뜳���[�Ul�8'����2I�D<�f>�6�v,(tɬ���er��Yѥ�<�ꜵX~W�wr{7V���c�S��|�������8Ԩ�9�X2�g����U5�)����u��Q�_�8���2X8����-�$pSK�.���U�>U+ n�&���K�x}��4��.���-:S]��$-�1H��} ���$'ꮅ+�ϰ&��� &��z�֣,U[��
�����M������*P� �I����Q�6�G�x�QF����5�g�E��������t�u�G�qSN|��0m�AtX*LR(>�^"-N2�`�����\7����(o�(%��θd����������]	'��Lw������Rr<��{�]~�N|�i� 4�����c�(P�P8pS7d�_\��X����425��F�0
��V�K�Vw�g=S�W��e���~��o:4�	�C<�n ���H�u��5�W�_DGƤo�?�%�!�]�W(������s�>@A�mt夵�$96��f��Rn�cy��E@MC�WiMW�S+�#���a-/���������J�ш]W�MIl��k�=X���җ}��
��c���ݘ��تs�1��r^r��'l�=S���v���e���>�{f��1�4��L�1��%�2i_C�%�n�mJ�� ��^5�|D3�g����,�B_�t�Nű˾���mYAП�U�^
uI�?�Λ�zQ�������ǥ���4z���/��Y�}1�V��G�e�/"w��Oa`)���ʦ�j4�Y�~	�)��a.�/��De+�;�W�mZs� 4�����7y�}P�M`�&}��U�+
w��f�D׻�Y{
AT��cPk��48��mk�J"�H�ʡ�I��"�cZ	�&'ڦ1�U�������l�=���m�����ݣ�S=R��
F㌶���B���1Nu�~��c��O�=on`���2�=�Y�k��f�Z��	�j4�ax�3g��}�l]�O}�߶�(:0�3I}�����"3xP��8
��D5�z�zc��~.@'�
�t����B��ڧ����ԸV��(�Z�_��͋�!xZ����FO��l�
&����n��έ��2����ǵ���`j�iϿ�EU=s�<�T7_D?Y[���j���V�����|��m����(l`*�j�h�7�Z���*ZL=w7v�9�q�A��m�������yUK�㪃6jt�f�/�i����1 5"O,;m�����W/G:�jSoУ�!�*��۴�kL�3OX5�[M��B�6�J"�����뺱�?r���Ʈ�y�7��z��h�s?c5���_�M1o �$�_�_VO���ډQ��K�a��B�t�n*�9n?9�s���h�Z�\i���9�Յ���K��0z�x�o&Jo1�w�#�ڞ�Zmc��U\�*Q�wz��D�I��]��Zf�G�5����v�M߇q��ES%�(�b5�}j"��e���	���5^��U�]��	쁭�M8��OY���ȯ��cpˉ^!��F�����0��-��W�-��e5���>��U7�!�-:V�-�=��?��h��]�R�5*X�Ł�Yȹ�;h[T߬��Gx�l��$�U]_�n��=��G1����U���0`c�� Z�r����\������~Ζ��j�����]�9Z�GsT������]۾�_��y��������&W �G�w7�O��+B<>\��JN
�(ɺl���������vnE�J�̭vvm}N�r��+�0�X�Y��� ���eA��\%-���q��r�����x�Z=���%ɰ��-M�O��#-�X��izڱ]��V@�)��v�b3����N��x�j_O�.�������|ڍ�}e�rA������Lʕ�3��p�a���S��g��z~�r$Ϊ����0K��
#/���JT����yH�xF*��?�ǔJ�����˔�٣�$dኪR�-%y��ݿE������Y��˷L�g���:V������lY����#ъ����ci�T�H��u������s��c;�V�I�	�я%���m�t��pr�����/�����N:�a��Q�sxy�0*�ڢR35���g7��^��Y��U��j.�m�����(�b�{S�O�[���d&�&��'��&^g��\]Y|���S��L�=����s��|��y1bɶֹ�\S�����''�ou�$h��]�.˸����t�k��}=����
���M����뢽����Ϩ��1p^����U�ۖBx�G`�D�\��Q��ɫyAHV�Z'/ˢ�e�פ۩J��V��\g�	���~�H�@���v�Dw!�d�"��G�i�&���Ⱐ}
�>/,g�~j�C4M�=[H�W��E(���?�:g�{���^�>�z#����zlx�ݹd>��t��R��q�7^H�����k��~G�NQ��T�HѤ��9X$!�8���N��� g`��Upu�ȑ��i
W�!�q�a�uێBO�mi�����Db�*�8 їǃ&^���(�����S��P	���ϱ��`%�K�6��Z�f��<�^tbN!Vb�Of��X%�}�I������U�p$L���L�)k]ƴ[��'��g�H�1��&�V�_R]V9aMTC���i�|m������^���;G��ݗ�QV�"	�-v�1��At�9ްt@���PB�	ԙ/1u�r�E� �ܴ�~����D�Ui��4��Z�3�|��_�>3�*6��PH�+""����Bx��
j���x:�<֔�Z�V �;}���h͗s�����c�I􍭉�ZVş�D�Mǃ	�c�Z���K�l�����â��=3�Ef�^bL�g*p�A_���
��O4��F[�ȶ`�EG���Z�?T����ߌ3M�oC+:�@���]��/j�;{g�y�;[%&NK��U-��.\����+&��B�`	�K�O�O�Z��+.G\�|څ�'
\�����(y��U6�g���˩��4�K����y ձ��ɿt��k4�/��o��rp�S�Qi�ϵ�WRT��"��9@b�	�)Q��z. ��Jb[���DD&��YT�05��,�*^uxғ��#�0_��Z��!G�M7 э1q�2�t��I++?��/
��O� ��3�D㡞���^[L��Ts�]�E��=�}�6��O�`&�k�	���PR��{zW��|���NU@�H��UZo�E+uږ�*�	�
e�`�E��nى����a��A��Y�X�ߎh�q�cJx+"`Dl���5�P�խ��_�6Q�5�9�*i�+�e wܢ>
ㄈ��+)/ &RA.C�K�qJ��8i;�S�l�W-��i[�P��n$�]*G�6v/oDS���M"	ՠA���>��r�:>8��`??��kj���h�>pTin��ڊ񸨓����óg�������Ix��u��̍����Ҏ���Y�x�R���'ݥ�ẁ��fl �d���Z�ՃA'�$/Jҟ��h�f$�`�/D�H]:�U��[Qm��};�t8k�:TncR���	6���h��X0�ɨ���k��^���
��������3Q�Ė%����$ �ϵ�_��Z8U�T����8��G�е��OĄ��^�)��:]M�.���&��{]�~����ӣc.��r� }\%�����CA-�P&@j�g��|��J��|���z?�&d��|>s��|�I>�M~�c)�rd�*�b���жS�:w;�~�m�a�m���;�65;�6��^�
��^�w{��C�V�e�[���� Q�:�@�y�ƍp���pxpH�ڋ�T,��<�`��~�,�����X-���E_^�z>dp�	�~TS���/^�Hۦ2��V�{b�N��;���^�\�C�@P\2�te��Bx�C�L*v |3�J:��0����R�O��<��G�.T �)�P:�i~������T.�s���>d����Ho�8�^��gb!����Ȓ��y�o߅��A�d�~!�a�����{z��TA|�._
7oޤ��\��+U\cd�A~�w�އ����丘��f�tg�%���I ��ǏIt<��߽G�{�}�v~�k����t?<����j�����"����KVټ�4�(��g�.>��@`�ğ8�㓻F��jb�� /����y�Ύ��T�@oO2�\̴��A:�ٌʭ�C~��Mx��q� օTV�~f.����$\�r�\�̠��͌]����g��H��(��֣���Gl�Qu��0u��ZtcW�8w3j�'d@y~��?������H���PEx��(d ;<��"8̼
_�p%�# z&l'�P�{� a���������߻w�t�� f��DtTV]�NJEs���ׯ�O��>ND�z��"F)��ɓ'4y �Ws�p=��2h��&W0����E����������<_�u����N�\�0���<N�3����Z��p}�V�T%c2�k��?���Tei|ߘ�u����
}%
G>}�� ���q�׼ 7��֠�"Ť��� n�KUmb&�MK �?�Jt����[�*�z����_���<���ǔ\���|��޿���^�v��c΄���0�C	Z�r�"D~4{������gy�j�D��Y&#	�ݍ�Kw���U�Ko���%m[�n�T��&�P�t�Tu�Wc�=�bO'��f�p^d���?o!����Z\A�Ġg�|/"�q���]ȠN��H�Mqo	Q��os_�xAAXX�nD�0"�}ޓj���K����%�>�\������_~����_a�y�9��1��ϟ�>�/]�d�8\�d�\��zԏk1���DǩɆ�w4�����!���7���Vu�#h��Z���a�j�/�-^�~�>�U�:>|Dt���!1]�v��	��a
��T���+�a xE:$�lhL5��P����;"���m��畊,�XR^C�7˓T���Ҿ�}b�zM���I|� �w4 K�5���؄+.D���\2Zk�`n �_�5�: V�@,�eD�s�=B���F4p��tP��/(�{J�"���5�t�Y��q��V8<<�F�}�;���_~!.���؎k���h�^����S��ܽn߾MtsX����~M�\�����Z��6o�8�{
����,t�cH�Y,L�Cq�B�j�][֧+���
�n@�y�L�X��k��,�p�U��mЕ>{�T�vn޺�}u���G	hsj��Y�z��%-��2�N���*�yAӢ�ҭ��D�rS�/
H�=�%�NCU�ٛ<�<��:����`��@ \����%pwy�O2�%���oџX�MR?5���~h���J���+�y&"��W._! Ұ�N,� 7��!X
������N��
���}�V3�B$S�< ,�^'��_�sA� )��m%r���^��d �J��@1�ײ�?�Zb�'�|��5�MI$�T_��*��i_�;��-Ĥ�sab���G���o�y~����?�b��I�;s���f>�=iM��KX`5d\ã��t�m��Y6śFRK� ��nJ�c}��L#Б6���;�L�1�͘IY�ÛL�/�"_�v%���K����L�٦���W�3W����l0(�g 
��,�迿�!���j�i�2	�xD~�K�����IbjTev���/�[��y�z�?�3���l��;�3�<_$�$����e��r�z��'���!��|������&�������#epM��h�CW�U`�s��e�O������;$�R�C?�-f1`�&�,o߾	<����a"�p�Ѓ�#iE�S�����Qg�<)�dB1>]�+���^t/���T���Gp�X��5���ac#�Y>��sߡ����$.���3�~}�^�z�*����L����>�ܹK y�/���@�����?���+����l/�*g�j�y�7�bq�F������G�@[m8��� C1?�ă��B:�{��S�1�Hs�LCqMd#p>R���~�4�a3-�̏Y���^!K	 X�}JX�H�3't�9�� A�翳)/�)�L'���>�P��IK�ӝz���������fJ]d�~<�&I�-r�#��.��_)n���;cHCWJ������U�J���ɍm�L)3� >>��M�b߽�|ٽi/�.b���� �:�a�?�{Z?�j�z?T��O�H��jN��o�������$#��8�|� "yAXЊ�&<����}7�� �}��ع>�b�G� @ �k�3������I	o>�'$�-����-����	~�ӿu��(�NX`�ڿ���t���)��Wl0x��I#>7�����߶8T_͋�
���	M<"G��U<�A��(h*�m#G���$����c�C�=����sV��Aq0���C23��V��!�d�@�ǔ� [�FB�Z%���$@�Q8ݥ���:8�Բ[p�[T���rN� ��}��r�X��HtCEFѶ���ԉf��{��ۉlG��!��I��. ƍ�y�h;�: (��F�$�G�8!�b ɂm��N�@�}��ӷ�\FX&��,���)o!�������y�n�W�.*�M����AU��)�-�)���A3��O��фO��\�[����A����'��A~���T�����2��B��ɋp��
�V�Ebiv[I���c�͒��� :���3���Yl� Q`�}����B% ��ɓ��ehoܸN\(�8jLU.ĩ�*�x��ex���j�?���U}3��h�M�$�АX����^�I�m����J��G�|Q�ߦ#�E@U�:Ъ�eC��h����@۰������3��G�,����M��fW?1��3�Ry�T�X̡�j�`� �tט��[��Q�>k��0a�@V���������ﬕ$����x�����U���j-�P�I^�4l%��b�EW	�����D���@�D^r�tX.l�P�Jr��u�C2�l5`��$Kgo(���	]*|�<6���I�]"��x0w̺�VR�a��Gs�3����}>И���֘R/^�?�t��q�[�n��_}���2C�}EՁW�E���	1����W�R@�� Tp礯������⨙V�6��icnO>��N�X!�IM2o�0�Ӣ�Ԁ`F��?K47��$�h� ��_d:&���`��A��˗.S�'G���YR���_IZ#ϑ,eMg��X��g�&� ��n��|>?T����ѿ�� SpZS	�$����>�9p�'DnU�J�����?�s-2��I�7�4�b<�Ħ%w�X�Y����_&\@�����`t��I�K	$��������W��#��kWIQO��D��*���]2Q���`IG �S�o������ŋ��x�W	"�c�_��͛�X����f�cDN�֘��q�G��u�ac����W�P�����VI�=��;��J�:iu����*�x"���	T��oM����r�1S]�.^�Hn�� �~E�	�=�CsMt�<�yo���	Cm��|���|).�C���| ��--h�(8eo7�#_��Ԙ2=�"�k틚���#��"�Z=��+�jS8�*�_XLO��V�׫�-�2�t�T�X쑸 �C�pP��0�@QEY8���J8_n�%�bפ4&�h�����?�"��X�[
gј[���gU#b .+=\T�s>&b��?�B�?L�|���!\vZ��(�A��I
���ϘxSϟ=���5�ql�cd����8�J��s�y5�I'\g���?Q,��&�y6�
�,e�<�h:7�^�s��s||��Q��<�S$"�
�ɠ94���� !��ܥ��(-��H-yu�J ��TՕ�[�q��6�lvj}�S�7ש!J�����ޖ�5�˪�D�o�.+z
�f�$+y`NS���ZNE�ٶ��L�%�&���=|D k��C��_���޾��*0weLl�p����x���q. N���q����G�����}���'h�;8�j"�3Y|�O�����&������ha/S��d�p�]_�7WC�/
CRl(�0�/���%Y5�p,��T�>+>K�|[M79ɏ�A4���k�|N��.:TNn��b�B��&�~�+���u	��s�Y��]iѮ+�L����P,�
ܩ���|\G;�b�U�_[���ѷ�Yl���y'����F� ���� 0M<@��=������ �R���[���c	��ʄҡ�����y���(�lP�����ݯ���|K�xGǒ�Dߩ�����Z^XR��U��p��?+E�<e?�K����9{�/���L穡�唢å%;�26�v�� ��;�a�9ՑB]��E,���	d3Mr`��I��e7�߸>����D)�,A�fc�)Z�l�}V@5}�nW���o*bG�7"�,���T�yr�(ⷲ��=�C������8<0�6��f*��c���Մ`�0�#4�:C�/�L OP���<���x
�Q��>��D���W���'O��u6�g&j.������8�VBi%e ��p��z��a�HA����~��3���`�~����	O�F�� R?���n'.�ێ���D�?�J�wl2b.ڐKR��*q�/~�D�����C����m��p�����'"uQb�'O(�|�����WwI�C )`��r,O��E�B�5ʎ
'�6����M2����mʚr��"��L�K̰z�d̡�m�'�wɉ�;�(�+�Ke���F(���e�㨅(E��k0G�}d :��i5h��uP �8j2Pe���h&XB�G �' Ap���u�V�m#\�eZ,i2�mc�r֖�-:O���~��O9kD��Ȅ�{�=�,�#S�f�{%1���?��� D2 ���O��AD􊜋t/,���Ç<5|�~(���_2���u�����k3=f��� ��e����C�7�����a6�,�U��}K�`M�\��������^S�����{ugrǨ�в���{����I�|���[�q0���� *���eՇAW;�,hp�T��J���lU�$s]L��fUG�At��mJ�P��(@:%D-!�� _T%��J
�MY�����\o��HE9[�����\z�t��6&e�!�=}����+|
�y%w.	�����?A3`u.M���2����c^<�.�ER��/u���9U.������pO���/X����B���p�WH7z)\�z���@�a�(�)�}-])�	d��~*���f�8Tm�=w*�6�2�6�-I���E�����B�ĭ]��?b1��j�E���ͺ-ٮ� �z�  W�n�4����2��Jy �z}���;���8�1�SE��O_������f��Di�:��)bKt��O]`ba�G�R�y���P����^��O)�_b���U��Yp#P`���ỷ^� *�&~��S�G�J����U�V=�&?7ݽ��V�~�ꍽU �h�'b$@��ר?�\ɋ+\���`�k���n	u�4h_\��Mk��Zi�<&zR�Nr��٢�����GM9�J�P.-�5��{�pw�(J��$��8	H`�J*J[�B��T��{������8SuM�Q����󂸞��zO����	/]S���ϣ%�U'�\,e����[�|?~B�>��_}F�����Im�d%��$�ل�ƨ'�Z�.�s�HZ4�+�A� FJӖ9U��Y��q?�wd�� w��*
�}Q5@� ��y�P��eo�ri���^����2�A?Z��
�,P	8�����m�Qۀ�Gu�RN�}��3Ƃ���f�\�H9���M	υN�H��b�e�IA����#�k]@Ճm�.�6$)�G��e@u��Dyo�ID�g_Α��D �bi.7VA�ďNqI+��A�R�,궤uċ.�s>
 K�iߩϧD%�����K,=��9X�5'��}Ho,���G�4E����."�!�g$����Tj����V����=Қ�yA�0`��k�χ�)"Z��l�H%(5�U�>�W���~��|�·n�����RA�ЉB�  ���N�-PB��r�Gj�7���?�L��:
��0�a��4�~%�a���g�����-�O��H���q��m�٫o:Ozc��8��@eB$)��J�=h�������9�:�VTF�"��%N�T�d�~�S3����m¸��w� =��V$�hQ���΋���D�)������Z%�'~%OpҤLI��{[��k�r��$��5����t�<N�V��P9ߏ��+F���u��_��$�`�g4F-ł�L�^�R�7mf���:I���@I�ˠ���)�������� ��W.!���T��T�R ��
����o�o���R�a�=z�J���G)�+�����0����T�<^剢b&r �W_��	���\�����%D��%�0���8v�c��~��a����.�Vq�P)S�M^��cB���ف��˜��a?jɣ*ю�AW�"�4AϚ��И#�?��GK��R^ P�:)�s��kpj�R�y��t�����t��[EE{��r���&����6g�������UZt�Q!Jl����K)9��gX������Hp#b֟s�Z�@���� h�38�7���)% y$�J�b$��}����"��<����wT3����?�~��{��T�p��W�M	��>$�0M��u��ăWqx�˭dQτ(�����-A��Y�w��i&�u���$�-8����I$��>�F+A#��M�O�Z�����k1�k�^�~�C�odp�z
����Ph����ܧ�t�4��ᓭ	R��U.)�~��5����<7m�>�K4W$cWKp��La[����q��\�[D���(�a�/lL4Yƅ�c� ���W�������NY�N��4�H�R�uDB谊~�ݷ�Mp��GE��8���Wh\R(I
�mT[�������E�����O�]�ʩ
3�� �9b*c�+&�Y��B�I�s9x \&	&,�$�e��>�-�x�2{����+E�m���b��QM��׵��Z�q�1�ۀ�8�rC+��ds��J�Sw�d�@�5���+2]�>5E+��r���@�VC�Պ.ׂo����$�4�tþ��}^$�?�i(���r��N�^q��ߪ7u��ؗ�V
ߏl�nR��(�뛨�۝�@iNu{�D0�w�㤜��ߵ�m+��=��S���$�(��1�(����a�9��!�<�``G�p� �?}�}���o��e�x�.Y`����0A)�+W_��"d؅L�!G���D�5�aq���m%�~>0U�"�8�U�/��M���Gދ���*��Ze1���zo�9���y���H�ʘEaZڙHV����<�,�2�%�0�� �]l�v�ND~�<[�k�����ʁ��Dܨ�o'5>�c��NW0�w�׵A�}�)��C��ѥ��S����}EYv@d�� �d����>��	D��@��Du���k����D\�"��D�D�ą���W�]���}���0��\����?SF)��p��k\��	)P/��Zo���_��F%1q!g����+;<�q� up� ~$�=��΍�f�+���Vj�INt��&��Y���]�u�$���)��[�b)!ԇ$�PJJ���Y���m�;�X�t�j�0�y��K�� �cb����-��E��C=��[D;s�PMU����
��'d�'�(�ۦR�s��c�x*5"r[���9�/)���D���yX8!j�>�����mJ����	˵��ˇC�t� �� ���L��`�W�5ĈX}2BeМJ�Q��(�B�Ir�gR�D"��op��,��h��)�D������O4/�7��,aKb��&#��4���/葔�P�`l�po>�"�Ph���ϥ�u&���U"��0�a��?��@{�O"��D{�v��c��qց��7Z��~7�^K��8P.ָ��mg����ۢ[��X���>�/�uΒ��j�	1a���=�(��)��Ը�$vqJt^����=% "��;�I_y F�jW0ItB�H�϶%��)������K��Ԉ���(�/T/}
УDذ�Cω}|m6&�p�B@�{I�lW�T��1��ip�s� .^�㔨f���
+�\Z2����/���<�>kSfäJ��?�^�T;�k8�J�2m?{p����t�h?R�}��ʦO�mq�fI�*e�	�HtZ�H�z�(/T��
!�i�d�T��(�˾|������h��%J�+"�Y�V��#�Y�W�q���xX ��787#m��R�=�rʜS��F�������4r�H�j��<�S���H�ʼ�r*���ω�8�,��ZvB�@P��_�J��p,D}��������Jɇ���u�&jb���"�:U��p�Wҥ6��T�8���Je7{��F�S���nc��V��D�X�����ӏ�2��D=���	�������jw�T*<����r�kN��@CK���̽K���uN�!��(��.����:r0Ew���1��~��;�B-����(\�r�is��Q�D�� 4 �v/^���/SkL�o�9j�C��d�w$�E�\G~`	���Z����S��DP�#6nH_���\� ��͋���jRe�z\��'��w{� �Cb5�_�^� �Уb1�7�}��.�(�8������*���BC)�br�_ ���7�~NPX�h�� �1U�X3�R��KT�H2O�gJ
�RДh�A΢�����^9hQo�)}�B�"����]9V�ay�纋!ߩUCG�  ��x.��W�.�+-nTu֛��e�K�(VO�9�E�ZXXq�%��I�Of�o߾�?�Hw�"���3�ׂ8�g�=��z��l%�n��Nh՞͘�}�6��"�	��huH1�7�|R6�ٌ�^������I��suע�������1е@a��}Y�%��%�C�@-�A
6�b��(�d���ϝZT��>w)�����"T���ӵ<_
�C��H�8��Ą�����xu���k��Ƭu�S8*�}�&��rC��ݮ^�Ծ����e�sw�����*�=�_Ǻw���Ƣ�Q]e1h�j�B:�ӹ�8�l��c
յ��\�4;�����RJ��O�"-��'�(�E"���rQ	+������	*� ��8#YPs��$#E�@|��E9�����uQ�P�.�믿���)%:�����ұo(��$���x(t�l��+�Q! �8W�o��`q��	�#��%1��R�q.g61CY\��ҩ{�#��~��2���ۖzÊ�#g&�K�R�Q8T����!���4q�f�ЀlgR�ɬ~BY�iޖ���.��DA��d����	�}rV 1K&q;�轶=j��͍�1+�dW6����I �Pt���T�����%O�P52C.F~��[R.*�r��er%��Z̜��5�������+��1�7���ʤد����Y_ ��ף��%Nެ�����D��ǵv�b��.P�;�K�����tf*v�?wnߥm��Zb��!Yt$�#'jp�y_'o�,�a�9}a�$�V}�ơ�I�P�K�
�M?zRԍ`�a��j�������⾃�S�8#�m��CN�����pbg��md��6E���"R�8�}�t�z���a�@g�Y���Gq�O"U5�&S(���r�
��Ld{���@L_�I�=Uj!7�}�B脩P�V)8E��I>���t|�@E2y�Њ�6���0t�X:?f���R]*���E�_�@�=i�xӨL��%��bj���~x�0�.;N5G���).R�+��RJ'wjo�2h(\G/��(J�\P��ɩ�x6�T?,:K�ń��n3:�ǃ���r�h��I2��1-�3W �C�ir-�r�
�T	��ƞhE	P;�`�F����<�9�ⶲ'�ۆ#(��� g�-%K����PC�R�/)�0�ri���X�p|�o��� ��w�Wtj�U҄�R*9�^p�CM�5 ��@&��W����m¡����$�Y�LJ7A��h�6�V
:쪪�Ez��E;A����� ;��\�ٯ\��̅h{����%Q�vn�<��|Ga���|�>g�~㕊���A�5F~K�:.����?��[��	5�X��B�/Ǔ3�8���ىN�Nլ��8qv��Vs�$K}q��'iP�(�î����?+�XO�LbIe5�Db�<�apb��RU#&6նp�@���Z�(�TC�-��r	-/��T��ઞ+J��7��>��*z�>�&�V�T�Ē�@��0.�0�}�/��~��9=�e$����1ZXW��T0:h��$�����?op�mf>J�|����1E�>"��G��b���ytrL�!=$�&����{�:ʡ�-)�s�y!Db����<�y�$��uA�Q�Ч7)��b{M��3;�ǵ��Y����GU(�hAߵ��]�cR�l%�u%t��B��-�ގWZ]m��g%(AB1��S�N�Vj8Q*5�9��2a���jYH'�A���IXo֌+�C@t����5]�����2���E�p�8��v��'�z���4�{��i�����M����e�H␜�E�)�.nB�X��4x��,�,�r�t$���O������U1�j��@]fM,��T��Xh�i/p1ᬛX��6�gT��7;��Z������@��`\,sjC�h8���x����r���S��FVЇF-���T]��":��R��%��w�| �� D�7�x�s"���5c��^�ܰd���=s��"bUn�<�:~���<�X�$�+`�	����t��{'z8�z���c���K4�-%>X9��q�;,Q�A���D�`�L�MU���h���­�����C�G��Z�:��Ad5C "_<{N%�o����W�`��iE�2�]{2�#Y���t815���gTav�mX-U�(�U|�D�SR���
�)���]'��{0I֐�R9�"��k��H˹A,�K��p��VR�� M��u/b(�a>���8��Œ�Kx@���A��bT؊`���7+lb��kD�B��Dʘ����8.�ol�#�"f`��8}u��\x�犱)\QƕV�$E�"p��_o_�~)'��"!�`�>�T?� �Zo�Ҫ���:]�%7���BQ}pˋ��%�5Wf�I��b�3�b����<|� \�t�\
�A2�N�j,X��I�J_K���:�0f���q���������PT3]W"���B�����U�`�[q�B
NG��S�zTNH�2���9.��׉�M�f�e��h'&����L�в���t�HO'L��,��Ju3������=���@�l�I ,!�I��;�O�X�V.:5 v�0V#+zm����+��4�M�`�/V�R���\P�r��j��m��Dy�j�;{z9���"��^��Z�)D��Z����W_ݶv�ќM�	Ҙ~�'z��
"A�>�N�O��?'��˗�eP���$ę�1�1�y�8	E].w%q|"Z���
�CJy�0:��L������c�ӪA]n�$V�Ӣy�#g�'�g�>r�� 8���-��.����� 7�E�N�G��n��1ȭ�u��fǱ&����v$�u�z�E��.h���4��ou��1`�f`f#���$�x�+���]%K�
r�f�I�Ul7G󶔳F�-E�:ӥ|X�+U����P��tq��,��v���R!��7�1S]z6?-�*�P5j?E֪��b���oI*{�����"�L�V���������|��K�\���?�{Vs���,A���N��@ߗ�m*��n*J-)R��Dy���4R$�4�fd~6�]z,�*0M���x��3j��@y�F(�ĝ���T�>��̉D
Gݑ�с���Dm$u�4JF'���LM,N!T���������+'����3�/:U�$R-̦�8���Fǅ*pgqg-��X����IX*��w���ʴ�:��FE�t�薡�&�r��0VT����ǚ�	�� VUq90�@1�w5�:���"90��d�T$��ܙ�Yw��d����:��>\
�Q�w.�h�	�)8Vp�0h���yQ]@�x,��~F@-����aV���W�薽������1V/�D�X������&(�1���v��
uĽ#�
�x�2�{󆲏/]-%��#W�<�2����	�Fj �(�3��S�6k{`@%"_�)�4�q���DY�2��0����px���Bb���}�D0�E��iEV���7|��i���(쇬Wȫ������_�,Ɖ��DNH�o��I�)�k���J��S�jL��C��Q/���M������-�hl&�c���7�����KT�pt����D�Z�K����eࠐ���ܢ �W�^���*eg�
 ��
�`H�s���⅋���(�Vm���-��]�/�(%<E�*x{`����!(C�/��m��^}5���g��Z�{OG�R\���!� �����r�+x�8�Ku�3� D��i&��E�y�)�j�dj�n�N'J:6�dc��)?P��^�krgy���~�;�4l�ʧ )���/�
���%��n�D|�a\j2�@9my�ՋTH&C��>�`� ���}�PO��5��΄3�a!�� ��a���Dn6�V����Q�C"F}��JW7��L7dj'Jԣ�NhWY��T�cE��N�*N=������TLm)���J_t�x���<!�鈀��:�J�E\ʤkM+Uɉ���v�N?�QjŮ8�U������9�������YS]D7����`u�V�J�����u��sr��N�g�@�|H?p�\���m2��9N2p���D 1�	tMHf�lU3��T���gQ�܋J#�z*���x�D���1e�G�^��t\k:劓 ���iJ�5��vBݡ�'s~^<#R�������B���
��^T]��3���G�c =�EYk�@O���%�IA�e�����w�q�⨊�6R[A��{�;W'zS�ƒ,��+4���($,�T�4/����}W=ӣ�̌B�8�Lf�����t<� 		��f��%ȶ��J��&�T{d�?F�0�9ǋ��u��b}&�ڱű?��ױ������%����}������d�x������Pf0{G`�(��.C�A��G�*㐹4ҽqJ>*A���n��d���	�V�`�����	�(�����C�v��G�U�h��?�z �;�)b%�;W8�Z��Ľ��6������N޿dP�����jU.�.R)y���i��9��T����AG��6i��޸�M�X]O�>-��XQ���``�S<�qn*��7o��\ �,%ݧw�a�¡6���!� "�n\�A�!�p���.��·�����3T� ��:���^3���D�4����jl?��P��f��r�>k�R[O�TSs�}Db�#e�Ղ�~����Q��P�9���B���xL%�) Ȝ�;q�	� +џ������~�'qs ��t.��3+Q�ϰ4gf�y��ɦ%�Ŷ���N�h}�^��ƇI��ꝉ�Y-ۻ�o�+����U}�cZ�
`���H��B_.^�j�G����3��~H�}+�ddbF�N�	�Zp����?¯~%5��?q�F��K���M����!���u�Ë�	j��|ɺ��s�`4q��3�(=��S���l�Q.j2U��R\���K�����$�4�q�;b�cc4_��D��Y#"�T����۲$����΀۾��3x�[ݔl-�X璠�5����"��HD���3�NJ6�̫�s.{J���_�I8TY�N!�8$��ҡ���w�۷H��=�C��Z�a�ވj�}�T/��Պ�}������ ?�uo6���?�B�����3I{F���)�������ЗH��2w7τr�^_)ɬ\�Z���de]���o#���0��ء/l-�L�N[q{��:���1q��8���d@��'���Ts&f���A�
��5 ���g�u󖉄���A������O��
c��/G�N\��+-�a��Vl+$�F@u��s�3�]�U�����U7��۸�U��W?��L��A�]�p �s�������p4�����S#ゼ�d��
,AZcΖ+b@�\h�X��fK��޲>�}nSk4�v����a�ߨ�%�FV]?Z)}̺��O���)ZI��"|��4�u�~��>��Y�锤P�>鄮4W�Äo�V�;Ҍ9V� �_~&�< �{���������q&�I&���o�E��G<nZO
��ݿ?�����N�	YT?�> c���wI'��U�NP�VW*��ͭ	τ� aH�*K���TǊ~�\"a�֒.�`�Y�������O�������_�9?���|.'��{��ܔ�0�8�R�͹�vJ�F%o�>7��h���W�I�­�b�IUCEE�)9M/ߥJ�W���&���
�$A�Hb���^�|It��û��6��%��	�!�@]#$��(/ ��]�O�������g M��l��A	�����ȟJ�F.7��Qϥ
���O�������&
��e�=?��)<��bȠ���gfd�a	��MXu��4�|N�Q}בh�� !p��|���H&qY���^<�9���`�d�J��"�i1���@�ʍ�R~+��{�(c?�� � �h]�Ɔ�G�н�en�`Q~Ic���K�.�kD�	D@��o�q/�{Ρ���0���L����-���T�������0�EK�;ƂT'R���ӫ��pxȺ3)_m��(>O��t� �F�4m]k'�PMV<#�Q��d�k���2Q@���k*^+A�o�"�jp�>��0ׯ^���&q�P1A��~x�`WO,���8|qH ���_�9�RMctB6H�MM�Vsj���F��X����<��K�"�]�����D�%�D �x � �J����DR�!94� y��p3�%�,��{b�gC�}���3�u+���4�?��%D����[C�=�<2Xv��Ŀ,��e<Gt�b8��������T�Oݴ@�t�Ŝ~�m$�N�J���/�d K`t}+H}+}/X���@|�� փzVp&�}�]���L\&8x/��X��Zd���*�����ne R�4=Y�1+l��Ɍ�����ǨN8So[��:w[��`0�X�c�Jx�I"��0*H/D"�$�lP�]c���$�<~�<:`�W���Y�Z
4)
�'h��;J��8�p߿#�b=�ܼ��#����"�v�� �X3E?+B�Z�v�L�9���}ōf���X�E�E��1�?~BD�;�3A,s_�A��D�K�1_�8�`���b��{eq�����  d���A%NP���ݯXG�Ŝ��  �1a�#�z�d�ӟ��~u�V2op$]��b��� n/�� 0��������	�}������P���5�Xd~����:QZ�Q$#^�3������������Z!�k�`���P�,�-W�]�7�9�_��1��Gp�cb��6�"ƕ�a�ſ4��I��]�=�X�(y4K-32��c
l9��� ��0������;w)��8�,����cq�ӟ�#��|�[2��[���'�����V/�z��T��[�]���jrNhјxM��Ǉw�6FUٌ�bT�9<�[px�TS��T�LA\�^���#���Q9�Fyb���2����_�
`y,�s�;��2� O�2�{�����[�'�<P! �>�cp���|����@-���=��5�4��D|sBqSB���3B��q'd 8�q稥�\[��TJ_���)~�1b^M�H�ء.@ZW.���[�I��%�`M�RAdW�Z2�a���E 
]�0�c�!Xq�8�ܴ�T�eM�Eq!�8m�r}1���7Q�)[�S%��~5$���i(Z��N�;�շN���,p��NA�; '	���3�����W����X����b�5��Ot�D�?�J��/JT=����S���(OF�yyw�~3��+hIxbnSd���P\��$Nz��M�'�+B����Շ����'R����J�VR�ㅼ���)|�.KI�9����V�_�!�f�)�a�{a�s�6)tO��#h��譄�B�@M\c�-`�3�QT��O���q���I_q)��Cu�:(�o������\L����ܦT�"_o��*s��NR4P|W=%�n%�����S �;��� %��й�<�mx+@���T�HD?u:or��_��NݕF���I�
�)E�-?bq�bn���V�V(ã>��Dq���h�%�����J��\+�K�td�w�y��L ��v�����/�鳧��Y���!�tG��䜒�Y�7���)/�����2��\��Y�/�MZ-`�l�Z
:DX"1�A��nߺ���Lhz�p` 'r��ۏ)V�D�qa�8������:��^$q[6 :D�����{rB�D��� I\`����lA�^+�ҋ'���'����WA�G�c��I�!Vc�8q?�`��vp�j`ڧlAd�SR��>���J�pe��"�>���'.��m$ �����{����%����
|��i��
ԍ"����L�����}�s����Rӈ��K"�P�w�K*�WjO��mHpI¡6��|Fa�"]g^��aR�<id��{�zh�.�Z-	
��W�FU�F����Ę/��Xh�L�a��~C�j�l�����K�cK퇻��:V�x���c0B!&�T}e�ۧ��*��\Vz��SB��/I�F*�!��M-�:X�R\�����U�i�@��\R�U �
�%�I˓d)�����?�՛Z,9 �S�Mh�87Rl�8U	p�_JZ���	���9rI�%l
xoF|00���F�,q ��Cc����صʪ.TM�H2����97��J�XX:IC��Qj�}�#x�1jo{ٖ����0�S<�Hs��&EQ��X���To�fҹ���dqo�;b��B�����_�xBRc��B��o�rN�w0��n��� �42����o8{���+��E�S���0��6Ki&�A<X-?yL�������r]�8��=�D7GJ�N&8�tM��Du��9a��/�C�D�/�gb�R� �|�	e���"���S�|�B�:��Z����R�&��*Rb&�j�3��j�1 sJh"!�b����alR�b���\�z��"��\ ��g�Rғ��Z;�~�~Sq��{c2�0&!��+>�N�A:kxQL�`�3���?uL�y):�3N��0�|ڒʈ�ԺQI��ʤ�K� �D+� ����C-�)����_��
���oo�0�KjK� I䊇œ��_� �;�O0	`0�ozFz�%��L
�oaWm{���YjH�׬��>Q�R�P�&����H$Vkl�-|��[��`0�$4'%;>/_<'Q�&��X�|�-qa ���٭�L�~T����U�ZJE�?\�2v"� t�~Š2�1�*�����Mp��u�Y}�~���\����"BG3��oݾE�DAOW����.�g��R%����{G�%�UER��ڼ��~��������~߸۶lI���Y��� 8DV�VѤdϝt�EV�8 ,���.%��>!g��uSx�V��~zc)�s�oq6:F��׬���q�g�x60�BV4W];4�b5Wg0[<g��^�a��&��|'���1�����ߣaɴQ#���j$��f�|��C����xt�R6�A7b��{ɹ?r�ݻ���+$���+�����Y0q��#��3=\��e|�n
�1�r��=��+�Cv�X6�U+�tV���j���Cl*3�I� �մ���z�'�����ʘ�3���ZV�T�Ȯ5�IB5�Yu ,z���X���'�;����_9[`�p)F�������%)���}dt�A�f��3_v��RB�h�����w0��U|,��*� ���F(�sI�u�����[wn'%_Qs�aW)�Yd [Ӿr�P5���H��*��h �}�7.hU���M��
gYi^eh>�j�M?����:Pڿ���2�PQ�����8����%�����J(�32^&w���;|�u"7i���ϛ>ϵP���
�?-{I?�6r�*6R>��=��_w>���0K	c;����*�)z�=�QG$���/�ڂV
͒I's�mFE}���E�.Dp�������ü�
�=��n�am������M��{�����GN;[5�2���B����-���S����0X�vS�I�V�\�f:
�β�+H�cQ��i̍�a1W,p�deϡ[%���+g�S/�x�L�J�����O�j�Z������0��Y��M����Lo�G�� ���t�R�^whs�88<��4�1��_�k��@���tx4��i�Õoz��)��O' 0\8��ДwD���ǳ �i �E�QG��!�A��5�?0��k��+&67*����k��;��$qh��x�Y=g�9x+���n����9>4ݔ���>F��M�n����6�e�9�3*�߁�k�8�fF�Cj�*ʘ#�;Λ er,L�?B�#x����\���/]Lׯ\MW����/_KYih��P�t<,w´SD��/�a�
9���v�1�p�,�Β�cm���㐣����P�y������N��%z�nɅa8Ii��쿇�wZ�N:�i�Z�U˙�~�RL�s�*�N����h�E���>���߯UPU�nY��������/丠-Փ�T�LM���$���g2�5�5{A<�?�Q��BWxL��7�l8Y�Z�N���P�E�u�%DM���ʊ�i���8(��G�}f�%��sR�x+��X{F�b�*(F�j��1O�
ܨ�u�模w��{�x������l����̴e�@w���eg�#皒��R���?}��\�>N���:.[��(g��Y ����Xh��R��g���5�2! �1�z���=[*�8ą��"jB�zX4�����@��"��ϟ�&(�	n��F�h�2%�����-à�-u�/Y��R�׬x�H-�a��i�e�x����Oq����yY-m��^\pRY�"{Y-=�7���Z��<�#4r ܚ�=�"����c�Pɯ�(Q�2��g�8��#R������V>�6%��R,�i�����2�I�M�R��RcJ�r^mbi�dO~o�R�ǰI�&���uu��$H�q��������-:�����fpQX��y�Vb?AM���sq��Y��Fl�=%�^J�:2J���'H`a��IJ�'���5�aӮ��čB��<K�ǉT��	��x��	�P��ug|0�� ��F����wn��-�Q�%������������Z(�؀����J�}�␠���>�� TA��#�0}�����-�M����Qw����/�m3�X�;7<��|cwe�t����Z�F٢�2e"ĶiצsS��N��i[��ʎ?vx)��f
���G�l
��x�#�	�3
�{d�c���g+[��-dl/7�~������^�MG�7�U�;����z�X������gJ�Io@'d��ci�^9��n:��6s����cx�NA-K�k����Ɔj`f���h�G�+)�H�U�U���˗U�J/��r��& �]�"�YbU*,�����8�7}5�?쀣�%�5g�c0��B�������f���)oǘ�g�Q��Ń�W�$i*�9	-dF4��0M��+�A%�	�wz�����*U�sJ�S���搚9�f��{��1�`:� L�ǔw�@5�ʸj��fsvJ�r�®���!T�3��۴	!th�:R�ws�-���N.n���b�@�.Wi<�
J��fc�i���C�P�q�ڍt��5	��ֹk�T�4!C�{�z��+E0�a�7o��y�Ze_�3�������<ix�Dll�Iǘ�ĈN@���MY��l�BH$?�IIR1m�@��G�M�^<%�F�Q��2�r�zX �	|���M�eҼ�]����j8�T0lM�m:m��>dW�e>/lA�#��M�Ks(��i:������؁�!) ����Q�9���F8g��C#^f���Z)➇ٞfޥ��Bl$��������5�?��?�ݻ�$��t6�������.�K��D
�?���<~,d8Hxx虊�H�X�����F��`��v�$~5���>p���n�-�����"P��D�D����q�t����)��������2O�q�i�� sRja>�u"������S+��	n�o��N���w��D� ��5g&Ou���q��z�'-�WMK�2H�G�����m��
I���/��/��N���y�2h΢觠#��,�,sy,��ת��˔�n����?+#�.�ijh�T@�zE9pE3U�#��)�\	�q��RA��B��@�B[ݱJ��O9�����MB��(�����Y��vQR�KV�t*�}�$� I�R��3[���<��-�y�A/�C׼�(
_�#���K�(�TC3����)��c���rjp�"�U�
G+�$Yk��B�����~+�������sp�B��!Z���2I-����#[Li68#��M��Z6	��[����Ѧ<p�����[K�H굇��M�7')��h�� �<4�)]b�j1��=+ H�������ο�����g}�m�;��V�c�B�	S�u\�ٵ��j�� ��B��*(4=�Q�)��]k��l�0�7	�s�T�<A���7K6#�	���'O�� ,@��޸Nq>���VS_�.Ꝗ�~�>l#�Eg�$��+3K��!<y�&������F�ϖ\h]�������a8⚈	 ��T������2��0	rp+!�I�����i�m���5�k�����G�
9��+���0YU���+Z�zy(�R���%P��Z�6jETٰg�͝R]���G����ݟTVd�[%Mɲ�"�S�$�3�&�Q=�	��UԢi�FC6D|p�N�2������Ҁ���?�xc/x$!-G�I"q|�(�w��myo�M�}�i.�kK4)�G��dcY@�%��A�-+ьg9cb�zK�{Jۄ��;2G���M���X.��_[�w��S!�r���_���j�9y�
��P%�H�gn1���.em�q��W_K���'τn��۱��]%g��7d<���:,'���}�k�0*@�������(P���ݫQk�k��KP�~N|F�Ӛ�8i�㌛[�ڱ��
�$�`�.�QR��G��ɽ�t����4�\��(_�&Ę�.d+��L�_`�Õ�QC;}Z�(�ZPl�L^����U���o�I���R΅D)������_�@$�f��H^Ѵ��	)|���̞U�f�CŴ�iO����}����[�'�������{�;�fI̪+��xz)�Gpȸ��L�.:�4Fl�����j�R~_I�0�ף���L~�u�
ԯD�.��r���g�8h�X�FQ��/�G�M`r�u���]�v]1�2���z��
�3��p��ɓ�I�'�7��&4�4TmD�g�z ���Q�@Ǭ%�gVMс�`�g/�[�փ�𚉖�o3~��~�2nr	�����lae���1�II!;�c��8��,���&l����]MPʻle�w-�d�"R��*Ʃ��\,���Ke��&|q��Χ����R�	��Q4��pU�=�>���H�i��}��Lˑ�s7�̬� ��P �F�6����p':P۽�Vx�tF�����)J�!�[�Cn$'!++�5����-���m���):��)��O�0+�>� ��`i���~#5���@jp�v?\����%�/��*X��ѝ:�ׯ]���}�>��@�Ii#4H@9q%�?%�I���~������y�UC}o�$nײ)�����s���P)l��9O7%����&�z�<=ML�j����<���M��M��K��!�WE?�X��It�m�;/�{�MRzKSXP
Ǚ�9�~!�{������g�vH�j?f�3�e��;��4�z ЊY!���=���Xn�� ԌGL����i���Nb�`�G�^�_W�����d�c��8�XZ�pc,3��]lr� d4�H�Ki=�s#Qa�8	�����G0Q��r�Cˀ��B�'n��ɿ��m�FKheT�S���K��a�t�n�U�p��M0㑉�zh��@�	�+ -��@�Ar�B%.0�Y ����]�|�wp,����KWd��$C�Fc�b	*:3��k��T��!��:��OJ�g�Y�`���g�O����9����O�}�	�p	#A��m�M!{��^�Y꭫�Y��Ġ�״Cm�z�?\T���bĕZd���$�j�9���@N3SD[�U�0�p��L<2�w��:�ciB;>_J2[(�(8	=x(%~���	\Lrh�0�P$�)0+)�b�>��!%�M�Xh9���p2��;ڦP�0���*P�K��A�炀Ƌ�k��c0bk�pB�g�>�z���1�_>���W:\�&�G�$��fO�:��pn����F�|��WŁ�7"،��� \Q��ʪX�X���7��J�H׮^������:,m^�.\�|XS0���s~�XY,2���"Gf��R�iD��s�����L&X����`Z�n��g��&Z
[�-v���q��h"Ɗkn�K���W�?�1� E9FY�Hj8���N�Ѵ'j�q�nm_�<b�8�V	�!%�W�'U� �2�'�=��P�yӆq����B�)5S��E\߮�Ok���o�J���?E�"#
�
5�K.Zg)Zd�,��f������Ŗ�)����i�\�r4G�hCGK��j��~f��c�k����ګ.�?������ڦ���,8b�tnъ��VJ?�tW�Ik�鹘��s�źcm+Nr�U� ��~	����K���`QLh��{������6�M@׉>kfZ�����SO'3g����q�m>o2��㹆*��7�g�p�mX�{~��0?���F�X.���^/�p�V-�,�ì=�5٨-Z"�Ԍ�0��@E�Lt8 X._ޗ�;��(p��;E(��<��W�D;�B�h���IB� L�;kC£����ߊ'f��@��BJ�=m����0�#b׫a��2hy���(�L��ʰ�x�h����!PǕs��v��H�y�n�5�a���bS!�?*�r��N�oq��lo�x�ŦNO'$]�{�A�Gxu1~�?͚�P�*��eK�s0�A��]��a���7c,0�p,��8884%jaT}:wD0�
��>E�ߔ�����"�/^�:R�Y��>��M��ٔ��Qu��B��?�5z�Q h�KR���V�O��gr��`�A��]'l^A20$	�Gk�3�����Q�*�I�>i�X�x-�#��{�@RB�%�_Y�o����tD'�i1���H)}�~��*�)�X�0y���;��v������l�3Yd���`״I�C!�u�޹9�Tƕ��]��Ls��ll�;����±f�s��TE�s^�B���e����v�.�+:}'�G)������2�Q
�mx�`ަ�K*砖���ٯ�`:w���G�� @�"u�6u$��whP�6�g����Q�3u�
Q8��܏:UדV��1��΋����Tn����f�3��-��y׍i_�y�-3���üs�Jw�x����26��Tɴ���-ޚ�d����	��N�b�0؎w E]n�:�"nJ�K�哛���D�ZQ��ǿ���yIqO�>�m':�p�������>x��<y"�?��,�?K���B��p�]+�&aO��Mj�d�j�4ŵ$���Ę�D60P�C_OM ��el�T
Osč�pĒ~��S�;��%��A	�!��k���P��O�Ov���`��C[��+��s���,js��/�l|��%`�h��!�Wu�~f�$4+�������h�0/����(P�86�A���Y1H�j��w>��L5�|�]�z3�Ï�&� 8Ҳ�D ���U�:C)�y	:'��"���-.��4��s��)��[��:�(P/J)�]��vqI�{���=#�V!ي�y\j0O�MW5�G����bE�K.�+�l(%]'#��K�S�ٲ��"�ӏ?���	
MA���{@�a�7_�nߺ-Z�6�cc(��,����V�<�cmʘ����%<[�er��9�~�CK7�+��\ʹ�U�6�%5�S�㦉ϳ���X�t����P�㜃PaC���_[걯�:�ÿ�MZ)�BXb�'�P�?�8u3���9ax�`��MR
O�0ƸA@jl7B���.5^B^�e6w�VF�0����G�M��Cg��~�1��cZar�h9%LX��M�,�%��Uc�_u���_M9m��"t�x�
�\R3���>�`w�\�i������v}�[� �ϒ�ࡘ`(��ة��/��9w�3̙[��Ջ�|������$4E����D3ŏP�	�E�Ф����0��KMW�dh.�x��f�<� @��j���4dj��"�,f{}4�)5|h��I�
�Yg���H�@t���18�'l���~�-��@�]cN͜���y��h�k�{{��ˌ������}`e�A�[�N��@�H"h��&��P6\\]�G6��ӯ�~����k,1�G�s����g�d�*ԑ��?�QM�����0Eh�i���t.4�_���tW������{�fr�����+H=R�U��5�df!oM\�O��5�'z�Lg�����oH <���QwTh���$��۵2�1�<��0�f.7�d�$�ڠ�C��j����&&��.^��+��l5w�����4B�`!@��A�~�}��=%��ZC`V�19'�K2(�6Dj3��Ա��S������Ov�W��`l����\�����<��˞V��4p�'�PF�g��fs���~,|�HsrB���,�`?���ƼA�n	���#�fjZY��h�$����}]l���X��r\�@�c`�`sݳJ�d��=4��gq�Bb�޸~��~U�%�b�x8����gqd�
���;w��cOxs�)�q4�q���Y75j�n�R�� �P�p_����)�B#��>��?f�8�k�H�gv,j���Y�s��{��Z�b�?���H�����)�^��.rgT5�_�	�����)��!��ф�C��Z�__��u�
SU�NX4��������W[f��W��3�97'd1�G̈�j�^&�8\VM� �|�.΋�/�%�~r��2Ύ����;&�:,	��b���d��a��Ӑ�К괿�N�t\�Թ� �l���p�j޽e赥���J���:� `��` >cq�#)e�^�Ï8�����+���#e����?�J	�C�/ugw!a{3ې1���bӼz�����6�l���\_����æ�9J��i)�P5���u֧U��=Y��UQb!���Ԗ_�q�E͘�^���{�{��5�N=�X�Y��ʸW,�em����]ٿ���L��4�<�
�#�H�{F�=ާgϟWa�D����3��Ki��7��, z��zk��O�>�f�C�`���ʑ�����!������
d�'�VFlb���ciy߸�0�l+uvH���0�U�&3�G_"����.&?��&�d��y�M�Ñ�%ơ=�M��ʐ�|�&��u�m��d�EPt�i���8��8��M�U��l�"r%�n�����k�G��{���טgBJt��GÝ���&kۈi�{/>�b��S�[��!h��_<7V�ך@b0Zm�UHh8G,��6P%J��~�Yg*P����b�`~�:h)r��Z� ��s0�$&'���311F�
+���\VV"8�"�Lv��;!���&����L�	Zu���1P�^<V�e>����uǼ��g"�`�H��W� L�g�����`U��['���(�1z��dNd�'N�U��V��G�ՋWR�g�8_�h6�P�
��
S�.�r��`�/�?�l���=Gk*f~�&��;w��ݬ��H��h������GKR�Y�s��Lܚ�L<sR�Y����{���>|eq��0�/]�)z�,��^}���s�K?�ZB�9�7j��;�B=i$iIbcK��;7��̏�S���ͺ4�}�C~|BԆ7�]�������m�0�2�:_ذ�Sv��j-\���F̜�X��V١��q��{H�:�,�ml��a-@5�Z����H�.��z&���woe����z�M��`6߂B<&X�2�?�`��z��(����N�ח�6 �.�U�HL�&��� �l1,4h~0&!xP���	)Z���UbEp,�uGf��]��]=O�3\�5���s�Q�N׮_K������￯�Ӂh�R޸NV@���]���b7]�T5�K��e^N�z���dY�%"Ӄ_���ߗ�Q���;�L��C�`�~V�	�c�`G�AdA��5��� ~�*�͠%B�ޫf>��nߺ����z$��Hj���n���E�H�r�Zk�3etF���oG2�TCD�6pց�zy�5��Y � ����Bɶ��X.EP���o�ԫ��o�/x�nf_|�U5��9Ɯsɕ)I��z���hu5�|'��9qf�X���|�����7��3��	��>
4QS�y�gY��t Yt�*ԮݸZ��-I�x+!yi̮!ʼ�:�l�����`�-ϾX�1e�|V�zb����.��]q<=��?�0� x��V��RB��@(}Avє�Aփ��I���[�nF�Ow|�T�pB�S�i���}�d����]1eׄ��X���r�؄6Y�A�OZ{rg������Q0c� <�Y�<�o޽�Ҹ��D`���䙤v޹}'ݹ{G�|�_B8b��N,]�$8���˃RC�D��>�x��^��n߹%B�Β=b������+�;����#�0�!� d���>cB�dӲ�[Y6��C����y3��� 4�s!�Z%	�E���?�����.w�M�\�0tq����0�|�gYhR��PY�`�"�k���+���a�5ee����Kt8�כ��Mן~y��? /�Q(Mk4�{aJ+�8g�3OW���q^J?~��W2�Dq��G�il\�3�j��Ν;:�H��%��T��)�*a�0-]-F�XKu=$%>�p=�H�mIy��5�1�=u���)��z�'"�&^Xl �'D3��v0�[m�B�lp���E���xA��oAb�ih���\A ����b>�v"���I.&0ǥ�������|�B�W�Tv�-���%���e��eK%�� ��UP��Y&pX���,�^C��=�Ak�E���:L{�}�
���U�W�A�)8����XL~��`�V�W�"���[|������Ǝ>$�
���"9bh�FY\�X�r���qh!B'ǟ�x�?3C�����dEZJf!lb�q@ bIrG�����j�����@�{����y�g���]��0.�U$⤮�K9������3q�NTn�����G�9��3�����M�ib���r��j�����$�+K�-�c�Dsڤ�d�ɍ�X��^�~��
�גƉ���A�"c�ƅ��(f�M�U�@��Ź�$���������O��k��c� ����~������Cqj7=�����b�"���]3�c�Z
��Q�GHk�o^�y-׃��{sY ��|��	95��PA����������/h�O��8� p��n�N�}����4X⊍s`��"����x�Դ�d����Қ��"�7ٟ�ҟؤ�uW�{d*�>Zj����GI#.�s!D�8GEt:�!� �N��\��t�����!u��l�W�W9���?�@����n�)$'���V{o� zG��h��Ip����eؐ�K[l�+WA���%=��az\M�w��o8L8��zY�E����y%��+����E��[������7��;����?D# D�WZI/��IrAV*h�0���8�ќc�$Rb�Y��J�F=��Z	�ܱ0p���&�I1���D�����|��1 ��p����qcZJy�#u�9ś`��}�o\Ow놂�ܓ�\dy_�������3��&��ZHU�X��'[�/Oj�ʹ}v
�ln,
3�~�^����L�͎7�D�ږ D=�DA�yr-NC
=	�$}�x;��0
�i��,�2��V�'w�e6�3>>�@uAy�ˎs�I�F�i�v��E��kY�'B�����s6(|ɒ%��2u��/�ᚈ �=4�*T��y�N���Y]�Y-&MQV{`�z����5�;9�Q��?��?��><+�gox�����d����V;}%��UH.Ŭ��й8�>�\iv� B�L?y�Q1k+,zPR�I��`6XM�Ɖ	m,ڍ��Ç*�DM�  @�����kt�w��M_~񥰷C��!����5���o�����k1�S�z*a�9��Lk<m8��=��J���p��]R�T¨Bi�(�M�.X��/-�1�1�����(a���lU9���x�!�ֳ�pd�����F��8-��i4Ԭq��O�)l��05��&��(P��S`��&�����5�m���X�衱�C�I&�k{`Z߸v#��_ߋ)�4Th�B��z; �w��L@l/_�pHB&᪚�R���ś7�7�~#���
�m�vBAB_@�W�!�,1���0�!� �!pᜒ8NI�\y����0��|E[�z�YcM���^� }	��u3�^ūo�7 �[����sq��7*�r3ea�R���-&���u�	�����:����ֶ�t�M�h�V��xl�V���E5�1���in�jՊ�)s?)�|`�l���>_"�;��h>�X�������j6���0��j��i���
��{�_.lj�c3vZ&���߽�
���i��N0&W艹f^�;&N՟���W�RGf	;	7U`}!���Ѕ�A�pX��G�2�`2-y]*i��52�eެ��� �}��i��VE��ƥ�_�!y0��K1�/]�SzoG��W��shaVKK?ݱ4�,���LP-ĉ��]q04Sx��6���9�9 ����17ě�1����ژ�L�2��ʰ@��p��X��1*�&��U-uF4�q������Ι8��=Ne�����F	���aR��J�D�q�Z�|Y��O
/
.
�lغ?WM;f6N��<�ب��l��s�!�5����2+r�-C߳
�S���П9>�S*�������=]�_��[-�����~7�x�i:��c@C��ʌ	j�Bh�/�x���~�(�ǟ&�ޏ�1ߓ<�V��,�"�l3
�ݻ{OIF,f�0� �/��)�V�vBcE,b�s@1Ghtv-����D�gi�AԿ���g3�Z�>� S[��>'��.>���G*"���
H0�Z�@t�l��pH�E���}.x)��X6��^�K-�(�Hh$�bT�T5��ZY�a>����ƹ����s����q&����"��'*p�Iǐ���H��(��2�r�=�\*4@�H�|$1��L`���������+��]���0J�fˮ���:�>(#�*y�e,��Z�=��m&�WJ��NC��=ۛt�/���l��wr��b��̴Q�]�|Qr�>C��+��I�X���͛��)j��C3�W�(����X�'���Ȭ��\ 6{�\Ⴐ"�:�)g�2�q�ʃQ�����z�����X��:蚩>rg�\����S�%_�6����0*@`��;��i���B�Ҝ�Z2�_�� �.U�����$MS]߯}������':�����:�m�N,��g0�KgD�}���f}jk���)���:�~��$׎�
P۬�a�]c�z�w�4�by�hm�;���N�~�:i2�8�(�rZ����:QX3�u�Z,�� ���M^�61ΰS�d(�����k�fx@�b�\`�����,�N@kՌ��A�4��'�J�j���p-J Y��*�3i^q�:>mݕ]d�"�F��X�
'���0����hP1��jƇ��?Z����N�"�m\�D����8�~;:�eMi��f�fFm�lme?u
C���$���V���"��M�M�I�W�27�VR�41OAE��m͊]�Vݹ;���`Bx��a�	PMi������w�8M���Ͳf��Q���Zdw�$TsnZjbg6�+.~�V���'2 ��P��2x��CR��"HYK��Aj1)����Q�,D��b�?�|�J�W�+�)����,������;���#�y�@��$�$�Soּ��0"`
/�<(��(��ʲ_f!dep�#��24[�:�,��"�-���`��Q�hԁ�UPc0Lve�nE����n���� � ޵n]�!��CU�pF��W������IT�6�-�M��i�y�"d��_L�侊��u��&iO���t��5��N�Lp^ͨ����?#F��*iNNFT�'� %��ʨgu�]	�J#SU�)<��-�$-���N��A��Z���*V���.n�����t����8$�a��h(�v;�,څ���k�I��$eP�ՑYnbΈY�4)j�Z�~��9��z�	%vg��7��L$Nŀ�<1Yv�V�,7L���LۭM�#�S?'�DP��a�ʘ�Zx����k>���~@}3�>-�G�z՗�f)�S=�����5<l`��(���}�w���IװƱ��2����i;aɟM�y�N��8��g85*-L�RZ�/[o3ü��H��'��b�U�Q�A�i^L0.,�~4\4^3�K���  S�k+S���{m��v��L!�g�&�3j����t�ٖ@�R��h����D�����ꔝ(�y�m}R#Ӆ�va�NS/�����z�wơ��=#�2?qB{G�K�y�ڔ�(��
6�*�X\�!e�`6׀
!h�M��q��^����_ � �f�����6�-wPLfr0�p�Z
�?%Ιql��F�O����o�P�Q�{h�c�&��&`�s͕�T4a�]��z0�O�3�s����w֮a*&�-�L��1���y�:ޅkf5j0b��e���_�­/���{&�4%��E�&P��J�{t��1O���2��=���^:��`��?��V�'�Pه[M��Bj��nM�� $��pSϝ���q�Hr�kKa�ۯ����$�H�K#w���-y�"j�]�&ro�f���V��I�e����'r�	�_��p�I�Y6ez~�m���g��X��ht��.Ϝ5�q,��{v���X�h�ك�R�c,rL,YZ�����>���fz�ƾTI�N��.����K�`�D��f51d�ֈnP���X�K5X�i�_�:���E*�Z����������s�';�;Wj����N�(����S:�1�`c�;�6�G�{�F�f�&j��1�⚑�N5���F6�ډ��/�����&�*:$U�Δ'��-��0�8�~Ӧѷ���L
�:ng�WN>b��`UsW��)|0�8]�f=��.�fOꈖJܼ��͖sQ�,cM[���6���K�������w(��1�=���16�=��1�I0����!�1�7xP#�>K�\)�Bu0���x|B�:�NrX�&ͣx�F��Vj�&��v��5g�����;J6Am/�����ő����,��|g�G�m�6JQ�3���R�>Sش�������k����2{>��~/�+��Z\6�M>�Q���Q���U��|b!���~]鼢�q׶|�f� ���ZC2�� �ti�C ���M�vs����{���J	�dC��,7���*������55�lʫ��\o~L!0b��ߦ�#�2C���w|2�J荇�R�IᜢN�o6;�/}�C���k�ײL��w��co
�	�S[��^�{���L-l]�C�Ѳj�N���Ԏ����0��̜�3͜}~uh���D�}7�I������i�8���־؞ܵ��H����:.Tد)!��"*�%�	22A�!�&��y����%�۸d�ćB\���9(1M�M�Yo���q`�J��䊙���l�sd�ny�f<̊����{���m�m�v	N�.�>Z���;���7�9YQ^R�[ω'�ߍ�����l�8M�Eۅ��}J���\jl:)�v�V��ǣJ*S/g��g��qǚf9�EY�(HHG��2+��w�[K�0��@�l�,XWE;�c���J����l��߈�*�"	�����C��;剛2U�A޳궹W2���&<c�����`��dLV+KT�2ވqf�b�b~��ϛ�4$����J/KR�S������&Ȥ��)���������&?��������;�:F���)/�}�QC��K}�tS��&��ѡa�E�`ݔ��4%3hg�T�.���b�l�pL���~'[�b^cK俓LՍ�RG��]cg��)�Ԅhg��!L;K~V;��+�����$���3b��Z&�>l�QR�N���LB�+�d�!�q��#��P�9%i�$Fؼ�y�ɴQ�� �Ӿ����kZ�b�Bzs�^cw�~������f;M�7���~j�!������2�	Tj5퓍&wIs�nz��4���&n=�_�m�ꎟܻ��"�lh.�f��*��5�7.�Ιb}�ߏ�4,�=v!X�SN�����ф�.�4��'2��Uq���k^v��@�������w�peXAg����~����5V���l^�8�M˒�YV���ۿ����py_��f�'��埕�L��/��l�N�\.�)���f<!�h!\�3���К�,Hǡ��Y�o�.���m������Ã���U������'bC�A�RgN-C�������f��"e�Q(g�����&�\t���TM�5��ؕ`b�1
��1v�6s�K���ʉ0bN��%vy�G�k<��P�4mś�~��{�_:�`f���%��Ǽ���k'P����o�H5���������*��W����l��,��O�c�p�F����К]`��q���ܨ?��l5��IL�a����<-�����Tq@�X��B�1����8 �}p�*��zdｨ����G��/���P�m�]�� G���
�5)�^�8va�W<�RU�T�IL0�^eh�L�T Bc�e�S���'&�0����9��~�-�;��w�(Z�RV^�q03M��qB<�<�:$(z��qC�[銈m���Z�h3�ᴻ�����Yk+n�ӑ@KG=�v�0BÛ�%{��*b:�Q�W�g����ɿ�$i�d� �f��S�����+R�z�TV��Uo��U�L�����62��&!H����I�=X-�	�h�S�C�{�>`�����ϟ�H?��c���ߥ(��؂6��E�">���P<�M!���&����y�(v^���υ8�j-��t95r�'��X �A8�&��{{{��w6��q�5j�����SmF4��o�9(������w����qV�s��aG�)&(آ ,���lLAӶ�pO�0ul�4��`��CLA{r�����xm�7��Eq+b��F6"�S�u�W0�Y̧��m �[�������1e6����٠R�M�y���w�m�Y���C){�
�/��J� ��_]���bv*-����9��&���I
�`#Y��n��H�δ1@?Hs�\.�m��؟�]��+#���~����ÿ�]W�2R��ϟɜ|�����v�:g�g�q��
��2�����m�N���v�"/�)�_XoR:��?��H<O6��C�L���8�V�JOv�L���$�YH��3�UUU2+Ⱦ0�9C�|��ڑ�þ(�,Fi�O�p>-����~<���u��˚���(+u������Fw$_>� aP��/z��N�Tt ��i��;���uA:����q1��j )�"YI$7��*b��B+�t���ى~�ju��2%
��[���<pv��Eud� h$-�>���.�s���+#��B����a5c�	o,�U�	BKE�&�i�=��%<!������|���ψ3#�_�z�x�G>t��?6Z��fV�Ok���R��ѣ*��X|�XV�Łs�5C�ីӅ��B��U��:WQN\�SU�ʤ�v�D)�a`��-"�qS�6�9�	[�������M ?P>Ƌ���B�Z�b�}���ˮ���3ժ>n ���H��W���m�ݳ�����Q�oi	Q��b�Z���&�H�V�iw�+��3A�3��MH��&�iO�4�&({���b���ga2jg֓'Zh&���1&����[�{!}��w�̺��J�͙kd��[�5_T6�v��������`��sF�#��A�ᅛ�0くA�٫�p��D!<�s����(d$4Ch-tj3��ʨG&tD��+�:����#���L_5�GL�"��Iۄ��~ϺP�Z�.#&����X�+�hj4�"�a��(�\�<���y��*�]`[U5O!  `6���]}�����=��ϒM�΁K ���Ȯ��d�n
��y�K/Hd��^�CÄ6�yۦ�b�?߿_��j�ߦ�>�%�`P� ss���'���G���m���[�"xv�VVkhge�Y����Ê�q�γ��c���H"�UC8::�~��<�\�gl>x�r��0��ԱAM��H�l\��cw
NUխl!!,M���)l�vN��8C��Q˜���	��?k��b��hL8yV����d�"8L��/��nE�i�1�;���b�� ����^�v#ݸ~S�l�!0�I�9��ɭ�U�R�-�PZ��`|�♘�X��H.�]jAؘFub����,�������LG�8�Դ��s��u^\�����ݢ/_<�&$�O��͛7���:ai�ϴ"j6B�2Hi践��xR;�#�� �J@k=��܇ڐ���Lnct
�4S*�q�>t��@����s ��g�L�5�f\-�}�c=^V3  ��IDAT!C�`�d�k���я��qГNn/�R�CC����m�"�/��&}�ͷR%�1�q�S,���~+N���f�3S��F6N�V�h����Aύ}�t�����V�֠W���F)�K���?~R��t�
Z��.2�χ���kL8D8�[�y�	�ꔊ���c�S��bh_��頶���{6'�&[*�S�f;���lԌ���pX�EB"��������٠A�#+1���I"��g;?L=hy��,m�%��;�ơ�B�������h�h��-��}��1��}���Â�V��ѯ��_�Q��i��d��h]�W�^��f�WGJ�Xt��9pN<x��am�sߘ �@N�5n�?߯u�	eйἛ�O�T�9tf(�) h�9��j{���d�駟�K�J�hl)Ê �Y)V�Ǵ�%������R�y�	o	6YR%R����s BUo���˪�~��.�����>{�X*�P�6'\��%�d�Ȼh��n]�����@-6l�Z/MQ��.@��K��m��u������V�9�������P'�r��99���GJ�%�& G��pk�Ү�c���:l�b����
ݖ�T�)�٩	Aw %E_��b�-#K,7�K�Sjg��>��k��4����*�~/���`\,�G<��N����_b"�{�X��Aͧ��oR�ߡ�43�;>������W�㵇�P�a���"���o�ݻ��s��fgWk:�C[p/��k�E����%���[�����pk��ls��8gm�.dmb��Cn*̱�Ѧ����w�z)j|��j���l\׮^K{Y��$�&y��;�i�U���kR�ϊQ�&���B��!��ի��!��1>�[��z���?cr�Fl8aUh�+���R�����k�D
���ul�^��@�X�FAI8
J��s��>��bs¦;�_OW����R^x��Ku˴��9�,���m�w(��SJ����YT��}��*�Ys��;}&U��w` v�p�R�!�v�����4Tmnl��pbL��Cٍ�ѺI
�EH��ʄ*���6͜:51�0iQ[���R��!9�i�f������j�%��w����@5Qh0��B�T?۱�kj�8"y0��'�l|V5Shh_~�����dTa���˪��*�N��:x���x)� ��/�H7� Z˓��Od!�=���\�$�e�5j�dG�z���}͉gK}��T�-�x>�0�ꫯ�!�xh�^pܠ/��J�Yj�6o[ll�w)��R��ʬ�tj��v�A�g��A��7�y���^7�Cl���;�Ox'l��X������ăE���b�B`�mb쟿x�~��C��W~����!�;��846a�_���5O� ��~�}��+4v:�R��VdLnq+?����8��%S�N�������l�m<��5�������i��Bi�U�#�3���"t0����SN�����Ζ+ ��gx6c|��w�>�(o!�R��]��R2a��A�(��}(<�3GM�{@��q�
@:�o���UJ����b(���&������{ᜯ��*]�rUڠN&5C��Θ	�ʨ�3�&4Q����ݷ�	f�k4�Pq���X��wK��Һ�C�(�k�_ntZW��R	1A��8���#�c���P(I|HI�D�*�Fh����|�^hN���w�eĄX`b��U�� m�)�sf�{���s�E��|�����nb��n,��2��IE�ӷu#~R�����_����6�բ�PV��Łv�,:�$@_�[l�h'�SD`��~�p����N�R6�����A��4�?�(����f�S+u��7�uZj%N�L�5�^�R���MQC��i�m;���-Mܛ&���d�J��#1�TL���3bk���^%{h����/D�@˔r�A��ϚiM���h�gp՟K����Έ�{� �K2-Z%2j�-�"A(���z]�/��P�GՐ �	\�����B��`Zu��ćb�e3���,�Bh ����#��� �$w�H�ZJ����Ii�ݘH@�����*��ܾ]��KҮ[�o���e}'3�I��C#H8>�%nҩ�.��-���9�#�y��I�}���0��"��+�l�[M4h��,4�	s���Ï?ԍ�7qV"��*~8���^D;��ע� ��`ΠO�Rmm l�؀����V�e��ք���G:��˿n��Ǆ�����n�7���薾�4��̻�ACQ��~~9��hj#�ϴ�S��I�*��L�����'�b�I<��˄Ƥ�{ﮘ�X4R~�$�tZ��ɉN���>g���X/C�b�(&>4��z��.�h��D//5k�7�y0'a��D�v���8���Bx�T����kMj¬�	�w،I2����u� ���w���" �e�z�m��+�?�͍@ &+�!H�R6;-4��۵Z���U �+��e���.�o��V��P�=��Y�5����ܮ�ĝj�3E��82�~!�G�;̿������`� �M�RsJ�YU��	��_<sE�P�u�M�1 h���֍�V��B5]x��8��V�l��Al�a8������N����&7������2�Nʮ�L=��1�O<e�l�n��4G���<��:k:&&����{	�A<߷�~+&<�`��1��0��&F���3h�4��C��d�BkQl��f#$G��f-[�e�!1a������a�B�� ���OC;^%DBŗ��`VZ��ﱄ%{:m2S64�tfI>���3���7p;���Z������X9T��"*v*|f���������|�����q�`)-�z*\�SB����9�����mVX��,��#�	�Z�)k&�
Tu`a�={*��6���~�{髯�V�{���wfC`�0�/4��JC�a#����[���Y�+'�kG���c\�l���[�G�~:���0G�7�.�6��0*ӝ~
�8�Fa;يE�I�&�Į���n����J�NYv�&��CXv��	�)�(��^���\h	�ijb I2px���LC���Th��Ы�u�P��u�`1|��g�A(9�
Ly'���5������l����0!̰�mp�$�:�����nH��s���U�ͣ%�|	�12%f^C��6�0���2�Dê}�_��_�Շ%��jGpH&�vz�[�{V��w��5�l�)�-&O�B� {��XJ���J���s��쩻w�v9��ٕ�����G|0``�/���>�����w��G���o$&�m���M��גz��魪�b����^�sBW��L4��W�ӶG��hU��|$��|N������g����S��.�o������)O(�m����z�b\�:#�A	��Ǭ'w����B���|?h������qw���J�f7�:Z�����3���U�4�Is��6�X����@�pюy(F�2���粏�5��H�x�:�5�g}����M^��&��3�f��.vH������"�]d��6��8�'K���K�I�-��06h�B������@mN�v���w�/�<f���`Fs\b<�
��0]ٿZ�-��I��y�+h��T�'���/�fe*6�;a|'�!7�����Z�}h�b	��cS��aZ1�d�(�
 "8���؝˽p=���k��s����-[�C��1?�̝}�o~g|��@m����uN�m������9�JUIi*���?ٻξm��Z�h�	^Z|�R0/��0o������G������vp\��h��T���"�V�5b����6��gfAC�f+���^�D�3	m�� Li
�am��@�a���)·�L6P�a�}�l�0���B�����G^�Y��H�i�Ԝ�9t����
iE�m���FK�AA��u,l2�ú�R�7�e�xg��6d酥՜b%jJ=�i��o8�[���Q7���|(��_|�e���?��>F	�x������	bLp_D0@�II��ʆo�#
�=�TX/p�}��w�p��U�<e�f3�{]x0?��@�%�W�HKqo	˫�DS�q��f�3���xS��� X�O���Nq��@�	��Cj�lX=�X�G�f�x�C��L�Ri&>��3ĺ��G}�p!3���yhG+�"�A���]�/��DF���M�)�[T0�����X��!%A@D����N�_L�b�"�	YDX�G�
!��/Ne��[f��.\C��oē�E �?��3#���o���.��
:���H�ڪj�*�,�o�:��x��i������߅�ͥ#mE�y�&���#�sF�؜ -޸��ԲП4�GR����	9�"4R&馶�C�`�AJ'"$!��}�^�p�0������R��/.�(t���Mep�?��,��U��y�x��{A��/�@U���r� ݼ�΅+�Ly`���8gO���w�w#�PC���4�Z�3l4���P.j�p,"��]=�w#_��$m�!h���7u
�La��r橷6�b-���c�}7��h�Q��n�N+v�F��v�)��3��V-s��7��떡5rڑ��d�0��Z̦�6����*�{�E����9*D %�!5Ar��m_�ZOJκ��D�9�BegxF�J�P��B�L;Rh�����+���K3M��"f�O���z�/���>���8���2��@��.2a���}�q�{FG�^� ���Jd�����tW�������ٔ�yД�	��eUF7�hV7J=�V��T�
h^um�q��?��� A<���B��zdRI�R��<�Q1�d�,Fx�9a�,0�7���_@�J�_nߺ�>��s^{ڭ����k׮�@E��C�!�y����hd
��(�&�g�R��2*F����Z$柰H�ł��"�&>6a��������'X#
 �1��ي�  �gB1�Ïyr�;��v��?�>��"��"��L�KM'W��f���~��)��V�COk����p���ܞ��뜭q	�V3G�i	�wL�D�%�~>��"2LF1���T��S[��=���.*,<h�8���DB�V0S�a���V�-&U8v�܂Z��&MuZ{��}Q�nf���9�dYv���*�H��-}T�M~��ר�I���P���+����L/}&/B���2�v,|��R�i��oA�4'��Y_L>%��(ϤO�p:6�lۊ12-��N��k؞�������@ӆ�!LY�YW�cX���N5�٥˦�&~�E)p��5�+�I��V`R�!;X3�:@��������L���[�|�Q�e�c�aRqImN(d��!��T�d�o<�2���A7��$&滑_՟��a��^|HLe��|ؑ��Ǥ�1��3Ϝ'-�(��I�L���g��9jՅL�&�f��?w,@�T�KjZ}d����Ex�^�cq�$"��W�h�a�v!��/3��V��-�kV�H-D�Cw�L�Qkh�E)ˡ�j�a�{Sc���+cjYSaC����6��J#�^��J~�Q.Rj%{�>��o�	�Y6�$�����P���/��3���	��s��lz�g)-��E���>�Ӯ���d0�����3��!����D����v~YL}�7��� ~����+�}'B_b�_�w)��eD)�I�4�@j]-v���}�x�� �p��t��U�"����#*\_짍���.
��L�F!X��i�i��ύ��^k�gߑ.ܬ�6#��~{�SIC�79ޚ�NɤE�D�)��_д��XwGL%�������鄠{[8��a���.w� |o�bH������4X#���
�eP���*LI\��ba�Z��)G*AѢo�O����C9�W�U�Ь���e�mf�]�<c:�����t�39����^N#Vy)����D��^A��o5�t�x/�A҇��K�ϒ���I�<�^�Z��B�lLsj�"(�F��f,��3% ��h;zn�1�����M:]%؜L���?��E ��~����<�{l��x5�X��L����/���pĵ�O�ޠ��}�N�/����ŝ���_X�=��y��O���A��.4�F7��N,c�J����`�-*a۵]W�#���o�Ҷ�q4�P9>��aMJ�A�xV�GA`B;`J�
͔�|eτ7�}`�ǂ�)���;qF�x�B�c8.�,�]'�{%��R@�l,B4��W�"ƹ�%W�C�D k�8�A�T*@教���I�+IMT�kɮ������!��u�~�/�q�1�E"�Ԣp,��~#��FR.%��Z�����SM����cO�	���B0|��vZA6#��Cv�m����m�Z8�>c�>�Wh�Z�s��`���P�0�U���S�\x6��_�5�y�Z6Qh���1����RH1�����%��Ν;�/pU���0��V�u5"�^j��z���i��/���3�s���Og�c�N��D��1��&e�*a�������h����¼�⠘����L����ґ�c�
Ќ#|�q>�y >ɔ���^�o�"��W��»:����K/�(T�Ґ��k�Xp~�|�R�\��R%��
�V�6��(>x���~4Ȩ�=�|��Q�j�,Q��%�g�p�j3��)he�G��X\����
:���e�ءO%u:>{_�M5��iR̴b�0'	6�����m��~z^;TTæ��~��\�h4�gCt�$&Yl����S��4�e%�=7�V��x.0�+���\X8�^���Ҩ�X��%uWRl�r_�����@�H��ۺ��m�-�/)A
�MA3��K
i��_~�p5@@3\ߡ/R�w@��G{=�Y�g�N�����<�*t�2>�)�CBF+�q�?�\"͚����(�y�����F���L�UT�������� af��ӄ�a6�gf�)0��1iR���h�/�-$������������ ?ĳ5���W��bq�AB��������Vq �x�=@@�M�`�e�0�+�
-�Wq��F	�m��x�����o:��	� t�6E�$hs+�(K�g1�-�"��ˆ�MЦ 5�M(��M���Ԇ]bL `���ƥ����R���:�^̌b��ԣ�/�@�	T����7�ފ�g��U� /�>L�	����Il�!W{l寵P�:��`�@��x�L+6�=�{:u�p�E5Ә�k����Q��fa/�1�bI�Ɏ�Gc.�z�*]}wU�%��-�Mq�щ���`��wpJ����1ԖO��/Wͧ���Q�X�=��w)�؁��d3�����zM$�+�9Gg��[�M�#g$��\�Q8.M�V/6&>Bb�!񄻻���ZQ@����M��܈(�y�l �%����˖,@���xBI �S��c�k�"��(8����(+I4�i��3��@#$�� -��o���ǒ_oV�J�0�L2�`��KR�!���	IS��ߋ��m�[]�ёnn"`j; nߺ-LK��4{I5^a�s��ȱi�fj`���+"�IƲ�G�(�$����3Z��z�j!6��	샿5�t�bUJ����Ԍ0����]K�_�L=T���,��B�r��p2

�K6��J7Ø�y�1\�vU|�I}�60�=&4%�֨��9�2Y�':��OS�$������
F��s�."���Qn2U��D�	6������i���/9�Z$P?T�7�"��ݛ8�Y�L�������\�}_0֥NV/ng&"�g��W����ԯ%����Q +оV̤'�L9;3�
�U3�M�#��>_����x�j�W��]���U[��x��eYL0�h��z#!ipP�R����jv�K&,4|�4���|���A4pFC�w�h���,�_���RJm�� S��YLjw��|�&MW&L+�27v,��E��P��&(-��A��ٷ��W�^�[7nҍ�p��]e�ߕq=x��8�`M ������*�d0�|67��xB��k6� �A��N�_-�"�%��0�̪c9ouB��r�bs�s~�M�'�P�9�wq�ell�A����k���Y��M�mtٜ�d��R��K�㦅3�=%��T3���,7�v�v.��D��)�NuQ@�B�3.5�i`�^��K��p����G%�5l��炠��/�t�����L���k���$%�n	�a��-^Z�dh5���xЪ��V�;`h:��Z����㫑%h�]�|���� �f�"��|!i���o!�^u��ņs$0�a7��k�8��*a����'7JGl`o�HM,8�0���K*��J�!D��;6Dh�S<,�*�:Y:+ݾ���9�FP���߅}
07Zh�p&�v�/s���|6�HV+f�$��BK�HYȧ
���gZ�!:{mM�&a��)B��#�)�iGn�ױ�5�})���f��������\X6�����\T���P����GpvqQض,��͋�Q
�[�d�̈5^��B�7{�s�E{*�+PRt�$���l4aK� ��څ���)�ͬX�Y�Ҵ���/ O�f�Ɗ z�´�&���'���zd�ȁ�_R�;�B���٣f��#����6jL� <�1�/s��fie��?H�Ms6tYP�1����h��2߼Ѫ��+:��ǦY�Moq.�8�T��A0��~�@=88�L7� '���g��ŘôVrh��	ݰ����G�>�'�Z\���+�� ���%!���/{X�B�*�u�Ю����
!��'����E�_�=A�~���gE����sgW��הAa���aS���ϸ��h��(CcY�l`G�r�u���OzC�s�q�g�4E<D��7u�h&o��Q� @:ݻ��29q�h�+�3�0����@'�΅XE�=~���aV:�������eq�INm��SY���;��<�/p�jUQC�?q�(&��Ѩ�wr��H�������e1Q�	G$�f�X\tR/�����K#5a�?=���U�hR+�[�\;�֊�9�qҨ	}�H��)��,p�LwU���O�1ycsd��+�ߠ�b�D{ȧ`[���2_�OYa"`�G ĩ� �o�j�ڃ }� 7n"��N���aݗ|�CT�,��s���+��|Ŧ�kT%�iO��#q����Q��j�W[������0���bp�(C�枾{����[��Ķ��o~�=�XC��R;�Ƕ�C +��~t��㵋��RD�Z�ѫ�N\���&3���Ke��ef��;�X=V����T�v�q=Z�/,�03���Z�J��	�Tr�x+ON�s �X�� IP`M3rZ��gE٬�K7.�,�>��g���ދ q�3[�Q��9�$�2�"�.�	Bءb�C�~g��<�0g_D�g6S���뉡��/�e�b����?Xj6�Ss� ��=�y����~�$Q��ZT��}���B����[��Q����H�K�\ZRQ���E	���3�qh��:%۬��e�M�W���^h��N������?���~I��ۑ�Nط��I���ݽ#�'�⾸wO��f��l�#nH���&}O%_��>��Y}���f6ؚ!I5Iv�)�p����?v���~_eFݱh�ĩy�q&U:i�����Sn��]�� ��ގأ9��o�	HU�"�Ò��`�_%�j?l^jm�C��m�mj��), �@��{�v%ڥih�4
=;���HNΥ�'���q5I�Ӊ�λ�s��������]%Q(lQL�x�	0�B��p4><�7f�pz�vZ)�|��4uϟb�à!cوy�o�ێ��p�i����{:Ϥ���jM���l�b�x	e��zn}m<��4A��ߦ
K�V������mr#F'��������ŵw��Y>�pA=�L"��h���%qd�w�j�RP6ɢ��bG�'�|n�����9%��6���n�O����{YC�Ȝ$�9��%��fLa�i�ݩ��9�����t�S !����p� FH��&���rK�l
BX��x	��*L�^8Z7M"� �g�<s��	���&5;}���u��P X~�9���6X����)'&��ɹ8���mLܭfo�ȁ�vP 3��� sW�1~t�h̩�c���վ*���e��ډ��8ęA�J�A&8�e���B��-$b:4�`�c�)9���Jؿ��-��fCs��}DhY��j�U\qD�lBs�	b�L{�J��|�`qs����w�HF3��-��W,x������t5j%����m�XHr�W���^?���f1�j=�i��䁲��7S���F���f�PjJ��t�����Եk]��v���L�ܞ�YJa�e�j�����T���3�u�{�M��'߳)�*�����'y2��b�p��쇕�^qG,��lV�e �=�װ,ӛ������<�&�)PY?$��}�V�XK���,�����Hy��dS(�f
�����K�n��i�А[z/����SbR�ʲ��h�E���H�ɛ��� �6ȨO�Ώ}!)o�[�w|����D�(F�T�L�G���&Ƹ�|ԓT��n%H�y�y&A��V|�	n����}��ŸZ*���
������Cԛ��E��ޙBe݄�X�_3�L�i�)�G�N��{���:v��%�������u���f��F�L��m�9�a��������x/�k�3������X��8b�N�[��ĭ���'�wd���|
fIl�unk7��A��6�:����iz�d������e�HKioE����v?�u[�t�:��Z��C���@��M�e� .S��߮i��G��:Y|��͆\�f����x�a��ͥh�;����ǳ�	�%��$ǐ���Q�1γm Mȑj-j�Qh�g��4)j��6;��a�'����Ip��������ۻ~��bM�YkYx���\YRs��yύSK��zD�<�9~�{Nӥ�Ԣv7�3��0ju�-�t��v A����M�����VY`i�U��侦�T0,4b�y4��6o
KZ1z�
�&���ݜMВ�"Z���mN�U�m�+��S:q���/}�3M&��|�r����^g@J�ݞ�2<���	K:S�`{G
�ɋ��;�������ɍ�]�G��ǹ������i�y��i�p����"�]�E�i�A�F���/JX��� ��*�K#R/��{�&cW4f��E|xs��V�[	�Af~��Za@
��36���y��So�SG��o/Lo9�����Ni:"�bN�a�c�6����Yl�>��Ij>��& M����-9k$�
v������km���|S|�9<9��`��b�Dੱ���P U�@�����4u ��s� ���VN\�y㯛�ik��(���K�N/%��?�M9�.�~��ߡ�>�ot�����ޫR��Q��{���hK��� m~f��-��J��YBp6�f@+u>�StP���fq\X2�F�yܛQf`�V��)��
B�Ǿ�A#�&��q8��8�R�=� ��`��x}����H }wM��z����SH�����Vp����G����2Tb���gO�5Î5�tTGˤ����c���8Ͱi��ҧ�t\,CCv���a��柷�i���M�(������O���kMs��D��M*���Qyg�fk�o�e��
�4i�n)!{���GIA����lRI��*-���k�z�:���Dܿ��h��Ў��֤i�blEh�Vdq,5Zz����%�Gl1�-�:��u�ǧ�)忘~D-��A4=\30�r��5�?�ny0������-'p$�m�˔�4��oN�a�L��Z�e�-b�x}{.ئA�]M��p�?m�s��n�����:w���]�<��%#v�n�f�/\����ڢ�\{�<}-$I^�!����i������ڙ����78ַ��Á�Y�,�Kٸ�t�U^H&Dyt�0td�"fE���	7���17Sj��1�z��߾�y�ֵ�c���F��;co����
����ݺ]�ػ�U�g�L�}�5[���C�E�%.Dy_�Q�	+�1�g	��ĸ�>�3�7����$���]�	���Ɖ��t�W]�Wo.��Y3�8�7	��,�=h=�ݓ�Mp�Er�'�#^gZ���(e��̭�<��׀�������m�@m���VG|�b�m�dn=�i��8�Iؤsn���;'Js@5K"���s�����ùM�H��~�3m�LEjp�DY��:ǧ���0q0�/�bB�q��Ʀ�1Gؑ�;�+p�0��"���@#
T���e��uc����&�\3B����u~��^4�z�z��l
k�����ЛY���֎Nk����5޽Yw����R/4ܒ	בe�sL�-���[ zj��!�������Y�W��C��$�f&j�����w�K���8�4L�����z�i�zQ������*'�L��a��hJ�`��n������>,�2X��_�8�V��g�qߧ�V01ݹcE�T�+\`0+c4�0Y�U(ʦ�SA 5U4�0("R���N��)R���wg���r�B�8?֏��?T7s�m1�Ȧ�B���%S�ܹbfX��ڂ{ʽ������r�Cq��4{�8Y�����9�	_ �o��B�O((��*�r���!�=��V�>��Ӷwq��a��S�O�a��{ns��-�c�{�'ZBܬK�*eΛ��M��v4�ʻ��qL���������>�x5[��L�ԝ֜�\�Qk�Mܩ�$z�����2����q.u}:��]c�/�&֏Ql�P2�w:�\3���	�'�L��eZ��f�M�Q��VNoui� I?�^N�:�Y��ƣ���M��?������z��֤�l��c���	̊���?{���ȍmA2��Lɴ�6�u��y�o���'s��9ݭ�7%�MCk;l @&�����e%3���E�8�9n��[:��5�����w����y�I��ԁ��n}G�_�2@�uٌ"N�����b'�^t���cqV� ��_�-d^:
�w=��d��G�b`Oo�T����P��$w���=*r�B�ĩ�)��B��\Xft����w���=cO��,/�*��?��}���)��j*I��8F�)�.ʶ.WޘRZ0��:g�~C�r�T�:J�.c���e���%	��/P�t(bț�yNc�������Nl�&:������Q~Չx�k�mT��z�""�p]S~g�6"�m!��Z�C��Y�c0w;Nl�0@UI�'�E]���޷b�W\.P�^_���zƶ���'��H��D���c��zc��[@�	В��ri
yv�2u��}��$>��3f�qڲH�Nl��W�`�hoi�q^����r��Uw�aٲ('��i�P��B!�H�e���k ��c����S�F��ω[�2�E�jz,�� �٪���*����f�՚��&U�Cq��͔��m8O� 2�Y3b�'�ύ�����r[���|^_�欚�y�:[�s@�\�p5����z�d#���,c,�n���h��;r +/ɑ��/����N�2���&�hJ�b����P��>�Nf�K�x��������Ь:�	�k�3$�>sOj����o�]rnL���X��YO�g#[�@��埵%��j�#�{���E�}Q�^�?��<���%�K�sM
�F�ѾX'����������駟Y6��|�}�5[�Ю�`��A�)��o_���)�$N���_Qc]��V��E��B1J�X�ӝ�o7Gu"}sA񕕿�T�c]B俤F��B{.����g lF,<��`V�0��:? \�Vi�ЉrU�R��.���ӧ��~�!���/�/	P�������<c�-lӭ��E%���Ъ:�E���-������������A����n�lr���^���=Ǩ�!�m/6�k7�CZ�'O>歉��f��M�i!��\��3s�ظf^�:q+�,GS4�ܽ��}�����a��g(�θR���yx�����Y�ٷ�����8��/ip 굔�+C��}��^��}`�V�T(�iذ��5�+֡��q��}L��V@�i�e%�7��a}�	`�Su؆�t� L�=�#|��7�Q���і(�g���3�Ruk�A�����i��� 1٫�fy�0�/���YW=V�f]���4z:�=�ݧT*�@̋�yx��%�'0U��;"�)n���so�ͺ�Q��2WG]K�{��¶ �Z��|�1�WQ�-^�	f'j��x���>4q�����4�`��3hb���ǳ���?���E>a���b{�'O>	O>���Š��H6�H���=��ڻ�׵�e�^�vs�a��JUD���4& �c;�3�1R�B�Á���slۗw�4�y����#&��߬WR.��7g��q*���׫H����_cekq��|X\�uC}�YC�H�Q��m�yK�{[��qB{ů��.,s��Zė���[.C��y��M������a	�C�! �M깴���z�;rL�`��W���:Z�xpbH<@m������̊pe��m�K�o=g���oq�RN�c�I�"�LY�V�����he�-�� o�T��y����-(�o{sК����� ��4ȑ u���������n�����a��Q��H�6�m��\�����u�%S��닂[�po���ǫ|e�ͤ��8��S��Q��.�Ey�h�!������B�^�s��&|A\���֣���zM�CFU׭qڪ[��v�㮄6���lDd�8�#q��P��~﮷��ߤ ���*M4¾�QS8�U��\�p �=~/�AŘ�ԌHN��2�-�m}'H�U��UDW�Y�aT��^�����U��n�GB�U�h(�0����FITB�' ���_�-�
���J�� �m!;%b���f7c,�V��K��>��5ZcXR�pԴN2�b�u8=;��QX��!�;� ����0<|��H̑K�>�q0�0���~nQ*��F�Q���
G�iW��ːN7���Q��I1̕�
�>H��4MwԤ��$�	$�6��O �&��ld[�D��,BCf�粋��ZS���)T6O���huLz�A�N3�C�c�G�Ċ4�6�f���&���xI�:y}��6���|���ܛ�m�X�O~[�s7vO@�8x����D���\K�zD���^v|O��^1w"�e�@m�������>_�ϰ�0��CY�TʡEdaϨ�tky��ryL�8��o�?���NQv�]нy�1�Q2���.V�54���/h.�䶾wt���UN����az��n����-sQPjjŕT*i�KdΛ���'�QJ_	*���+���wEXA�B�4�	�(&k�懗Kf�u�*�*G�+�� �� 5��,V��� ��L �<�h@�Z)I߂l�k�'��<	V� <�	��3�i��X��o�BI6Nj$�Cbf��D]�s�<G�´0ᏗGR(g��<؋��zx7,��� B�9����(�7�%��8��cX P�	ȱ��h���k�]:u;_0���ek��M�y�@j�Űb�9��<>e���gd�BcnL?��V�9,%�P�:� U6gS���q��+����+���!��դL6�!��脋�7�+ԡ��n����%]�9Kg�+�t���u�h/e�)��mla�D5�Hm����u�:d��`A����s�a�R�ֽ�)G{A�B*����d:m�J���m=�:�gOq���BT�U�R*��3�H���^��Jq%`�ŉ�gHw*.���6�ӿy�ִ�N�`Yb+h�eJv��6K'P�H����s��P���i����1�И<�e�9O����4�Me��uCAa`�����S��|�	�e��!�^f��dp8=���qJ�fU�ނ�Σ�H�Č&�h�I�π�����-E"�ԁy� 񘪍q��)n(y,��Ld��e�Q���&�&w :�LC:��2���(�G������KuDi
�I�?ZbxI�d�-O3�~}���C��z��&�&Κ�PKh�3[����s�\I����Ҽm���X��~�~�34���7d_zZ����˱rmW�)��L���̓�S:�)��Iv8�{�=h+sgeLz���4EY�R�NK�{���
-m�a�{��`�7Ib��]�Fe+��2���X���X�v4
���#�����a��E3�Ϻ@���XV֒�Q{'�:�uuy0!G�ZS�-�I�n4@iYg����rq
4��
i�%��P�TV-��,�v5�jN)�Ny�g�:����,,2Є�PݯN��NVe;kL&�����2�s���P����[&s�&`p�P��u��@ܧ�����3������A�Z]��yzr�N������x�����cѧ��e�y���������g�4!�$ q��=���L�m�_�z^�|��U��'��G������=�������� �\�l ����\\s?�be�yK�ٳ�ؾ����ً�<��z�*�I~�M��>]��G�=p�˗/�N��6�}wt|D����yx.�'�&��7E�	���f��P��K`J��U:�9���}���!'K_�b�2z��u9��ǹ��Y-#S���.����d���qU˚m�cd�gꉠz`���w�Ők�e/�{�@�4�A4�х�����3��7���o���dKvf�݃�j�� ��NJ�؛?w������O&��uL$]E��ցl?�/�N!=dR�I"���2k�=H��P2u�3�(���R��z��c� ���a�Y�@�,��
��5a"���\��PY��fz�.3�^�IG1��&��< ��% ��D��e�H?J��E�Fshl����P��,&:��9OP��	��Й�gy�Cܼ���'@-��\���/��?�~���*�{ƅ�����f�{�� �a�{`�G��h�y @?��s���o������D�F�?��#
����Y`d �P�������_��Wx��%-"h �|���!oǝ�_z��ze�nLO3���0|�6���;TV�������_)���X��P���ۯ|_��T6��x��b��\I/2�L&p�":W��t�:/��lx,�z6'���ws�S�����>��ʔ|U�T&�}�k	<�$b�z"�O�MݿX��*��v����k9 �U��T�R� ��	���A�Gz7Z��/�O3��#9�y�� �¹u�r%��4���t��H~���(CjU��k��m�RE� �?��GT+����ϟ=Oό�_hR��K�5�����O?�4|��gP ��d�_�o,&(O�d�S�/D����	��ӏ�Yf�p�"�xW�- �����_�X�J%�ڣ\�����"� �,�ϟ���>����d�����΢u�w�.L4�s���d���느^���?�`l ���q%��>f0����O>���Ԙ%�
��������#���s��ˌ�_#����(ba�h�*��+�����ȁ��WT�'�Ë\�?r�������ᗟ&VN�23,����o�E�7�ɚ�m���������Lv�(LR�2Ii�`{���X��� �֞i�y�̫d$<��}��h3̙(���A��P~/T�ǪaR��X9�O�* 
��窚��[R�V�OoP�B�$	A�B;�ty�?zp/������$f/�X��n�%Wlg�휼zV�ð̬".�h�}	��d*��Q�բ����3�^
zP���{�߫�o5�	
�!��8
=�	�7�������w�}�Y���b0A�nWK�_AO|F�	��}�E�?���n�(i�bq�"=m��`h�e������(�?~'�ƹ�E/�攐c��w����s;��x�����/%�d|���6�G�UddR��m��� �W��e:�5'�QP&������>����<�5�{W�%���[`���;��a����@�s��Ԟ/:X0y<� {�y���9����o�E$���ӧ� K��E��D?<��)1֔�M��6��0����9Rc���^L���KO�����	r9��S���ms�Kv������-=�UpC�P�^D����D�N-90�m�r�xu��oPKs��"�#��r �yB�5����pz�!}*��2$��1��>���1B�	�y��%ۊtO+�`1J����4�N��Z�-E�$����e�������B>�}-��A��#�x�>��?��A�{b1���1MնR}a�p��H�����}���ٟ>'VQw%��^W�vҷ���=���g�>�7��wXO�����69y/]֤r`}�fŢ�!���ܸԊ�����u�>3��E�*n4y2��t���YE��K�68��mS�����("6����n�|���PųB@��b��ږ5�2�g��?����u;�~�w_���`����:T�Gfu�N�i\�[�5�V~5@����x*�I���So� ��\
峛��I=Txw�p��b�����M��~��H܎��CM�!�]Y���o���CF}O58�;^�p�eRr�ץ�gN@��<���*�CĂXy��UXg6���l�V�db�3=1�<hO3;Zf� vx��A	`�N��QI�Ʌ���)�C�`u�	���w�*����U+�Z�5�%>� ������w�~Gb8�k�|ad%_��%��,�`� E��102 *�@��-* �^���G~���,��8��t]�=C�g� I4]��$0S���w'�QX���O���s�;��32�A��g�ŒM��-وcTXh Bx�(�#Ó��#aC̙h֋A�f*�����b��Kx��_��\� ԏ�r=�=<�,�ۇ���~�#�w�� i�;�~�{�)xweܐ0NN�߿w_�\�]ISuRHl�:�����*��NĮP#�H���Ѡ~��LU
��U�l|�L�5Tתz�GO�\>�'��ĭ��yZ虑I+{�d@8��QV�%���jM��4�s��͑��E�wu-
�o�q�ߗmЊ2��z�E����<���v�T�|�y!�|�� >y��C8�$CƢt�l8'd+z0��&d���PGT_vb���`#p�I�Q�)�-�����4��e��&��MDLcf2���F�?���M�L����q�e�����R[�� LD~\W���	������(��1�,�S��rE�Nݤh��]
C���
m��MF���1酿����y���t`q`��^�2�|��j ?  ��	��f����xb��1P��»��w�``��t�A��,	K �/WˠN�`�P@����C_r�,!m���_`w4�k�,$'��8y[����w��s��@Is�(A�+���d��ҁl谁�	c	Z��8��n�8h�T��Q�}�NEwځ&5~)0[���4�y$�]��0KN�f p�EB�͂e/�l�V��JMt������T�%+�s�<ȃ���GF�!�C�����Eƽ< 2��fѕ({ �ҩ1��8@�%�8�ݢt!�ډFF���F��g�"
��������瑷��X
ۯ���>e�/3��(ޣ4m�Ly�'�-z*���o���xQVhnb~	LpL�� �O��za� �6I��}'��;b��lIb���	-�+J�XdT��$��``�A[X��q U��+|����/�_~�e���O��}HV|��y���t��	��$����z�nq�:X�Y\�A�ܚ��$"��O@4���@Gz[�*����ft*,{-lXT�� ?�� �ot;��W�ﾥ��E���5��>~��H�Ņ�ƻb�Ӕ��e�B*#��Y��#�"�"R$�hH���R$*2bnJ�_������H�&���YI����*��t�;@e�l��I�J�e�ѐ�wX�H*���{|�E��=rM]����ZÂB,����PQ�QCŴ���Hs?b��E��0�h��FdP�`YFV��i�9YE� �y`�����H�b���D�ď�As�;2��"��*8�1Fdف6%3>cR�`q��B��D��b��_�����_@�8�z����T�NEQA�IaB�'YDV�ƀ�d�B�W s���3�h���믿�1�ַ�:�`��XT P d(����&-.X<�`ȁ*�qf�����_��ȿ>|@�$��~��G2����O�f�z&����(��e^��3��#̏ ���y�����f��^����q? �~�X@��UYQFq�WR�o12����t8��ի�t�G������S2�)�ճ�oP�@�/��m�"^ ib-FD�x @�����Sx��3$�u �&6�I�}Jcߒ�Ś�;�:Ό���BP�U��G��dzޖ	Z���?�~qa�>A'k��X��~���`(�Ev��~x���Q^�@��}>y��^��.9��r��j"C,�!�P(�8�x"�8��XjDF�2Ơ����iH���w���I��$]C�g�����X��yp塚W���K2r��>��R��6e4P��Z�,9+�dD�1{��R��1[��
v�V⨿��Ւ]�4���,���S�T��>��qDbj���x�c-u�&]�Z��������W�3=��T�����j�PQ'��}>�@�ş�D���}���߅!��؛��1��=�=K�IEE0I�3����%�V_Vb���x޿���q��*T���2�A<�H����;�
@�&��F}9�}���`:���G�O�����9`� v�45-�G��d��ܢӰ����ޕ� �@��:��>�`7�����D}�'�6��y��=O�5U�# ���Ə,jþ�<?������uGK-#�pS�*TQ��Q�O�;�y;p � &dW�рiZ,"�9�U/�{���&t���(it^8�Q�S�w?��a��,/^����B�^7��-w��b�����\9C�ΐ���Q�dV�?�u�D�(�Q����.8����GyUBƩ����~�b�m��:�N�,T��AtN�ٚ�9Ƀ�E��z=|�(��,>������ zV�q�z�!�Wpp�Pj"�#tlQT��7`t� �D�R��a����5D]���O' RH���'�Yd |FL����ڳ�uK��q/ 41�?O�[�3ƍ=��	�������z`P�;�1%速�9�xWf�P��9:d�/�:�(A��C&������$ �AW��CL<��?��?����2� M�H�-�[}��"1��?7���:F�Z�9�{�9#w-���\�`���iႤsĉh���[ڄ��kQ5��T&Kƴ|?��g�}�%��P�+ s�U��ǟ��K��(����^ 5QۓKj`���ʿ��c8��- ����"�i�A1���g�Zl� -X�i��"��|���Acn3Ʋ���ċ�B��>�PQ�	T�w�� �X&��E�x=��ȓ!3�\׳L~���瀨�G��'u,�yp�FD~29Ex�Y�BL(-��`/=Ϋxe��p2f�V���=(��V]�0��Fu��M��YXg�|��3���9
0����5�%�c`� �$X�3j(�����J����力]�T��%�F0����������s��|A�X�� �+�_�,yE,8SX@Y��t�`�؈��\r��a�%$� �<Z?$Ƌ���ً��u�����e������0�ί�rcZ--�V]_ V��7l@�D�
����0� �^�+ꖍ�c�I+�(Ɏ �Ѩ��V�f��+X���<��}�ДUm�&�j}�`�^�J �v���ɓ'�P�3���dĂ4 �q���b�J<1x؍����4�GN.��3�b7�Y�[
�_��ڮFWU�RZ�["ŨٙDX6����6_KQI`�B��֡2��T'*7�azO}NCs��1��������d���(�QV��H��	�Y�p���t��s���-���(Lh���^��h:f &�f�yp̆
1��41>�_g0���D���G����V�3����<�n@d%y�x���,�VL�����H���(jf0;���8���
5��Hb�1i9��1���ù�F�7�3
��a�J���0h���L:gU_H+MZ�<�9����Sz��(��*H$�ȣ�������-1bMF�F��:$B?�0��h��2֦"��GH����mX9���!�F��g��Ң��H)�,�F����Z^����I��?m�'��f��R��fѲD+�U.An������ʈt�>��"?T$5�Q5��_��������ŝ�U���1��0U�Łk`f��5�EKy��c�$����RY����xǅ 0�Ml,WQn���>c��ʋN�-y�t5;Γ�񇜾���,<?G��(]��X�`G}9�y�,�'�B�E2(-��Γ_��%"gp-�h��N�슒��TwU��_���i�F��M4M�K.�,��Ơ�Q9�tN)�ǚ&�J���(�2�X�R �E�	a�d�5� cU'���G�̆��[���	R��$Yuq41*��fX0�o%���e	�\2�I�R�W�O�R@��&��L����������D�X�L��ɔ/��R��m�@��ho�����>�XNn;�,����#D�8T��3و��|Syw5��v�����hL���uBe3�?�̾���פO����b���Om��ς$�1���X>������wNT���A3}Q@���1H��h�J~,����Bq�R��Ƞ�C�4:���r���H�u����(I<ƴ&��WV��+��Cz���,���S�7� �4�7"�Ujm�	��L1��
��r>Er'�˂|U�S�a^��CQ6�T�Re}:�����sb�Hp�J �D�������4�i��u�n<xPG�Rg�VlX�1�e�1�ġNYp�+��d`�!�?��y|ϡ�`�e��<dRJ}!����^�Fp!�(�,(k��u��p��'��E�����J@f
0F�=I��ekoU��b(��i�aZ@5�Fb)J���={�P?
j�䲖 Օ���;)���Ȯ\P������'�_�{�{�����^PV7?�mf�ߗ�/x<���x%ޟ�Vs�O3�ܠ������w�Q,��LN��ƍ�g����n��a:D������M��D� �h�9�4��sƲ��эǅ��Q��U�T/"�飼}f� �I�@�,��{,A�E���`�j}FII�SA۶�����R��>|�E��$7�\�C��fm�.�B�ۢ�1yCWR�&P������}_&��Tjm�0Q1��peO��]���
��xr?�����|99�ǆ7{��T�_���rLR�~���0��,� ,x@��M� ��Mـ�DE�u��E~�x���J�|Y�MEeʒ%�](�^/�m2hB,Д�=ܕ5�Jj?S]�����<�H�1n�n�HZR�^����$?��\��0$�J�(., p�A�ls�]
� w� 5@��@l�U �u�Aq�U���.k�X��j�	c�*n���e��t�`b
�݋�� ,�Q�s���*�"g��d�C�#"�`�Ԩ>���4�~G�]ӡ�T�pRxu�
|h,4J%Η'�*�ԇ���������WY�Mj�r+�.NI%�E4b?�5=�:r`���q�h�>�Ě(�G�qh�V�Z)�r���5���b���B��G����c��x����x�W)<ً^��Ǚ�|��禗��`��D&������A��C7&7�)cC�T�-_�K6�b��$�ą�v���A �թ�(G	�u�D
�_)��I�6��0�T(zRMy7:�����R��,(+X0ݤzN(i#=��ǓS�yo�w�l�$����W�YL���+���V���ʍ�Tp��XP�Ht����xhF�(��,?g%?d���8���Ye��R^���(X0�,Be�;pL�=tbTsđ�:^E�[[~��^$Iu��0��'�|�>��BiWz����@Vd�����W��q��ӅU�"��G��+7��hT$�]
hp�XS꼳<H��@]�8���4���+ʛ��D��u_뉳�����nD�"�z�FT��-���:�p$�TqEg����${QLam>w�3	G%��#bG��34�.dP@��r0O���Nп>�����X�Ŀ�2�AIca�Fq���L�Q����)��UaN�(��i�8ⴟ���QR��{��E���W<��NSu���['n�}���[�-���t��.4s��}R�����/���$��R��Ou#۟�	���RG)f]� �Oϖ|��&4�aL�����*jS�睧$���L�M2�36
������;U����ֽ�m��y�Kц M�(�z@���K*r�1�y��,��X���#�&I��4�_n4۔�F�ʉa�$�Q0�Qc� �ny�ْ��#����E>~���e�I���"G7ɺ�*��a ���gu��5��4Vz%3������Y����\�w�"$F	�����'��	C���	 �+C�(�
�S0¼��E �3�t��o�����G�e5�/�l����SJ=2�p�8L��S��)m#3V�0�՜�3١�㨝(Y�hRl6��HZGuvq,q��܏��E��Q70R�꟒�<�R�>�/�Qi���:�$�je�:T ����~��(}I�s��S�,��-��_~���&�����/�z"�h
��h%G�(�{Z���$Y�x;��l�#Xd�
Mz�>����X4p��.2�"@�y�SF_��P�g������:��hG��vzm�F�w�8�N�d�Ň�5/z�٦��|�~��4�8�|��e�Kɨ��e���S*�J7Pe]K�tZ�b�^'5�Wd��������>���0"?'�,�ؐ�^��X��>;)��"�F�v�ӃA#Wr�P�!c��A]�6
��Ⱥ.�U+o>�D�Jh)tjH��Te��D�v͝J�P��JnL��! �(��)2 	��*�	�ԐW�!ļK A�R�d��������Sm���4����Ň}<GۢE�m��X�*�0��,/$�L:P��EHQ;=�q�}�7X$(���I�B�%j	�"�lL��D�1�F�:�%a}b$d�H�X����pO�%B������N}Y�\�E�¼+�.8}�
�h���K@�:�E{s�|�G�(�`'����s;�"f~�fd��X�E�Q�G�K	���Q����'{?�.���u�H���Cs]�unk�R�Hz盁����bu̞+ N,����k��7�V�ݖ�S�)j���,��RfƧ��F�[g��$�ʋ�`y�8<>zB~��Xv�������73�;σ��ޗ"��7�D�VЋ���ف���Eu]b�`+�m����O9��(�P1�G��B���a��/�D��R�K�K�3�iF��P5IE�P}��"7!t$>�+�jL�Ȏ��T�3Bz9Up�MfwdHf�a��$g.J3�8���-���B�3�2�B�p���(j<��������� d!b9�7E�eвJ����ͬxc"��t|�xB`Խ�ث`(�[�@Y5V��/ʢ���C��.X��8�R.�~F�b�+�.eAձk~���l�҅��i�����>~HI���,�:��X��dҮT6�H��0
Cg>@���w���
��� +����j?Y����Ư,���!_����#�I������V>�������$Q	\�
�j u�`l!�����;(ڐQ�*O���v)ڏ��#���4$΀�|r���Ӏ���`b���q�����-K�3dB
�~����xvt̫$Y2�V�'u�^Ȩ�	C���i���%��~L���>e����ҧ�`B8-9z��o��	It�Q6Oc1鈶$yD�
H�pġ����~���9iL��bQ>C���'��E��oQŅ�,L�P_?sm_��~��%+����Wf����_�=��ӏ���&���i_�Ȫ��Y�F�̚���܄.yiM�(�Ӷ�⣸��Q��i�3�\�V��";S<���A���-�E�����x.�W��ҬO�%� "�l>ಏm?�MIm��8������a��셅�M#��2G� ��DJ�����`���*{��:�������C�K�=�yPT�7�:��j�/%�9}|đB�����щ�8��n5G�=���.*W �Řd��52'��l�nUo,�ڈ����4�
|=�R� ��ºA�X8<
���������S8]�)�	T�>��l&?:@��ê}��q8z�0����p���o�H�'0evA�āqi����jE1�eP�DĨ��5�������o�ὤ�>%u����0 ���)^�w}>�����W_RRҡ恴L�����>����!�o�����ݷ�&}�H���N��#2�I��l�ےR)JT��,���p&G�֍l���D&8>b0��aM	W�
 ���������Gg�_���������\�u,9B��Cc����&#�
���(�������A���&zM��Y 9���Y.���2_�zj���d����>���~����ܿ��>���ꑤM$ϋsk��qm�<A2�s�FzM�A�z ���T�?�����
���R<��$��"�o7���ϛ�iS���0Mm��U��z�@:�)m��Lj7�9/���SA�H6m���J'Z����R�T}���ʥ��O��3��]4��Ģ��MY�v"[�+w0 ��r_�B<����p��i>��SނDҟ��|�lQQD|�|5���ۃGI|��]#�p0K�VK _�T
c[:�R~(�; $~�ظ�a�Y#�c��ybS�)��$��,�5��\L,JG�(�\�O2�~�����O Qh��Ĳ�~��aaQ�� wv���d��/[c2����Y:ʒ$��u��f��c8���>���y �.�]��N��ɀ�\��O�D rUGp���8��%��2$@}�	�b�6�Ÿ ��%���Ph+j��"t�������]�<���>����{�d��?Gs�?�Q	���p]{���&�L� �s�4f��
-���=��p����69e�4<A(0l*���ȳ;�\$��B��;��<I����ѕ*$t�5?V{�`�b�|����
D�"3�J�^���>��..�+��}�
�uF���(D]��9�\���Z�?���AD=Z��q;Ĳ�B���V�̪��AD�Ɖ�1�$&���K����X���DY�(��&�) "b�a�03�jz-����"]q�!m���T�|�)��[�(�R��ǒ�6�Hj�$����XD��dF��g�_�=�`��W/i�#�tx�*�y4�R���B�)��f�gk{1�Q{�* 8�0���e���ʜ��X��e��,է��B��e)�>]�{�5�Z|������{7�)�����4���C���<�,�ȃ
w��(��I|��myV��)8#�;�oІ����``:$�������g������:�B��j���\���T�L�AvU�Qp������j�-���b���T���P��*p�����ù97�߅���]�J�L�0C$���r
��>,0k��W�)|�w][8��&���Q�2a���&�N��5+q����EĤX�P0�('bݧ�=F��/H|G|;t�p�Q�
K�<�����9�J���T ��8��(1�%b��}�p��d�G2�ӳ&8��[�������	����_���H!^�|pݲ���jit��u�E�W�c�����:ޙ||s�f���\T��	F�$����l�
V$���G���]���J sV�)��օ�r���n%�X�������ص�}�(��X���T�C�R����J�|�|��^�B��`��R��������*�q@����&�905]�����F��u{��[�=Ь���R�=ǯ�^�}��|L �E#]5��p�F���
+�$��/��p�6�px�O>&�vOE��81��9>��q����1&/�����>'1@����/oЍ�$������o�{�X�,c!�'����0b��uf�����CD��h�l�K�$돲̠��!���?��Yp��PC,��i�ح���d6��\����g��"|(����4G9��	j�hw��&��PPR�[����ԿV�y��,Us�
�������4����@�
pl36#u�����s�����!���9�9�b	�g:Á�N�h���Z����[��f=� �y�h�g*.T�ۣ����]��ۍT�6��)g��Ki=��b�M�F��3Q 5HP���  �u�x���L���爔�`���!�T�Ȟ��i8��ڌ
��(���i\�$R�(E?E��k
=��)[��QR�X�3�ń$�}���w������_�?��?����E���$ʮ��m;�\w��H�c�'/{ ��������(�0,:w��$-U�d`OD��fxD!�N=������h�3�;t�
�z� `�lQ�F�Eie�F�O"3	�e��^f�7M����E�Fc�9L�HRu�t(�8
2^e[�q��]� ��Ds�ڨ��w3�B痛8��ͩ+�'7u�p�i�:�{�(IV�L��4��D�@M����0���%?@����z�y@yk ���0!��������^rnx����"�}�*��y���!2C)�pvec��?G+��a?�$�Zδ�:Z���A[q��#=�qY�L���]4���
S"&E�,I�A�MI=tPN}wB�I�y�"���yXhw ٱ��Q��8��	q
��ZP�G��f])'_Ѿb�����Jˊ���IK���&]!&����>rޅ�L�(]C�T��$[HN3�������"����"t,҆�ܨ;����
��������'�e�����a��a���t��x�`yv
%�@-����,QEzU��w[A2&�.fR�喷
P����q�4�΍�����b��.�N.������jwh�Zk$�5��j,Q=�r��?���g�g�X�녊��/W T���]�M�8�rFF����� ���R����ğ����dː��_�O�#.�N:L��6[Pw��F�z�f�T%�o�6�-(���N��Y�&yO/
�3
S��3iT�M���E �Gf�2N���y!��d�O1������a
=WA�j4�ݔ�&�OW;yWהe�s����Ws�������
���j���lXltc�nh��frt_\Ry{ U�{'�l/��zKS:�R��(zid��� g7��I ����j$��%����D�$B�@Q+���'z� �v�'e\�(�7t2�	���@�nVPA��~�p�����g��NeK��=5o-R�N�sU�wAl�b6h0�}���b�:�M�p��fM�K[�(�S�*pv�w=��V=N��6ʅ�&b�Co�A祠*�X���6X�#N�wߗ�̀>�
�[�+=��alIK�2*'���<��)�3%:21�<�䕬2_5����'o� �a١+��\�g�9��:D��C!Q��8���� j�1	�ǽv*�ys>;n�0Π+�S%�ߡuT�N3(�I�Dw5�(�"w ����B�a$����)�冩/]
�)[y/�'�̀�X�4:����C�I�ȅ-�)w����b����lw��-��($O½!�#xV�G����9�A��D$�Pq9�������X���`�[��k����(8�+�#����c���Ƚ�&��(� R3�Ҿu[7��!k�.�%L7u�q"�] �~Kba_
��'����ˡ��̸_�~7��e����4y6�"� �毎7}����LY4w������ �/���z�|SYC�@U6���IBB4�Irh�L0�O�~��ȥ$_@Q��:0��C���J��P����qK�-=؄7�� 78�q�w"7(2�q�z�� P�M!�_�^��Sث�<(��gl�����7r��VӜ���O:d�e��ʾ�uH"/�eK��Ce]�>W��T*$u{�Uo,Lu#nt�W3�9�Q�5)l���)���׫Y��~U�X�'t �C�c����z�%�Yno���ԑ~��O��5����o�5NR�����c^uW}[P7D��c��;Vj�S0-5/m�n���}�j��R��m�QDΦ�bTv��*��d>26\�1���Ì-�	��"�D�aЭ/`5?'B.M��ſPҜ)�x�EXϠZCEI�z�����"��>c6�M�� [�˿��or�W��)E��3��4����u6���'���K��������S�V<>�a�sI&��V��JU�,/E蜳RM%7�W֦C��W/��B@������S�j=ϒ�S��s��T`���"�=��4M�@�+�G{5�H�U��@�Mw(��TE����z+������%�$wu[�
(�Em;�mj:�n�q����"��Յ�3�mצb�{����hN���z����*P���ԈQ<�T�cO��[�V5�*�+[��2�WX��6���ӳ���8�jl�d����:{{�B�~REAU�6 Z���8R��*������A�� ~`wQ����"�+����2�b�A��W_�����cTI�� %^>q䘶ud����dɧ���+��N{�(�:eA��d�ɬ�6h{9uPP�+�Jr��� nR�]J�bM�.["�:���ܩ�m����4d�s�.3��ɵ�EW����<#�����>��-��I�l�R������/=����\5�?ۉx�Yd�0�n��I�I�WzD�`+������b�2�ur�OKǗj�ʽu����( ���qJ���B������,�1�S�T�s�V�G��F�@���E%.�(
�?H�]F��������g�hP"��{�d����-�iK���Zr;Au�w���I6}f�Z�\���.��($v
��6	�����K
P��}C[�I=��m'��ල���������u9�v�8eX]��rk�yn�Z,ˮ#^���AљN���˷�&�v��v����u�_-R���(�«��]뙢��&����4�_��p񺟺���*>����^��$E�����`�R`_JX�&D�mP�"��� x-�wG�VT&���7b�oa���zYqU�m��8U)I%O/��˾�Vj�}2�5M����Kq�z�$M�y�+H�K�2Q�:H$5��h��[�Z�����Uo��+�k�)���Fm�@��G���CK���^X�%H0��T��1��� �f�����x-(�f�1��� �͟뵩�{���}Tg5U�*wMl�T��O�n���Q��� ꔃ)0y�>�[��]�N�K�����-������N٪z�b��1���y��P����^�g��H��_U��̯WǶ1�r��1
����o��'��s�ҵ2��#N�������y�	�_��~���^����1���L���ggＭ�_�d���p)�Jt��\�8`Q 0PI!Գ^�qt�	�q��>��gr7;���_j&�7��:���wQP�q�ȏw�.ft������H�ff/��3`����M板lz��&W_b�I���a��Ŷ�Ü���?�f���y���y�y����09�㝥+�2��N�/��N@��^&f��4�R#'J���T�|�R�[Q�������N뮫:��׻� ���V�ru�'�F;?5��?=�B*�dLTۥ�&m���~������g�TU=�b8��Ec(��j�ھ�Xxqu��r����������XO!%��4U����9^���c�A�iH��d�P���$�d7'ש)ی�5�APV7��T�+Ы 0��hD�N�Aag�]d��<�hT������$N�0����	��&rMEC���tǛ���@ʟ!��F����5��ޥ����zm�U���W��ߡ�a��WnP� j`5|I3N�7�2�Q�[��� ��r!U�LX�"�^���º�%!�c��jߢ��[4�R��U,��&o���z�#c�U����u���?}�'���CWY�����W�c���3��Y5�}�$��uI��g�oo�k#�������K��g�MS�t)�`���tu3�?;�[M�T}�R? t�ڤ,��j�C��.��}�GեvX 1�����jyZ=�g�Y�ŉ�*�kJ:JhKa�>�@^�A�Hu]l���m���U��F)�絈�3�k����p��s��Bx.�C���?�L1��xb!��.��8�ZQ��؃�<��U7�}cF����b/��T?�nR�k��ϩ1�^XCp����*� ږZ���z�34�Ԅ�5���إ�2B�{Q������}(�W1CY=nN��+�U*�ep����!�p�����Gh�IUF��Q�I���?[l
:���ň%!���4��Vn�
�*-����2g*>*V�Y�j��d%�{vӀ�dm5��{�vP� �X>2㖔}�p*c�]|�݂Η�N��h$�X�V-c�jðoK�W�j&zťK�nW;OK�ͫ��e"��bsY*B�z���\���ġ�|v����z���_��i`ks]��N�w7_�:>_� M�0�ϱ̦U]�u��m��u��(��U��\Ԓ�)�ɹ�<�ع�D����D&�Fa�a,Y�ld�e�e���[�i�^����N:����������*��?Y��0������A�:?g����R�Q�K;�P�"�܈�Yu�1t�f�ѐ.T������꒩p7)�����=�u�&��Yҫ����k8�^"2��UG����{������q��ƶ�����i�kGC�l���Ӫ������1T<c��ܞ&��e��x�YC�������$���n�4��>�By�&�ְk��i�f�qb��c��l�lY��3�R�&�g^����")��fR\�s�J��:����.���gR0��d� �@i��y��R#g�J�	b��7�m*U�(WB��<OZ�TU5�%�Si,�g���r�5徾.z��53���ô����V �H	5S�7A��բ�@��J&�R���+�jU������l�^����Ǣ����-s75��;�g�I�2�m�u��J`�E��F���Rg�a:Dh�k�VQ�� }4��z,N_@w�����dI��%�HP����rjS���D�'[�ͻ^���M|��������!U �?O%o�:[�J�R��u�طx��m�Zܚ���2�N��wi�ʉ^�������9��MYh�n�G�6��J`��zB%��0��sj���I��g��H�JHR������?�l�sկҎ�d�]JNc˄��ɽ�+ﻡ_�,@U��M=�T�{M;�{b�~J�Mc(ɢC5���6g�{w�F
o>��+������Oг��c��q�M��܌��`�e(6s �{�����0����B۶ȶ1ڗSUQ�V�!^�N�Z
#�)ex�`�����2�Ԁ�'yT��ʾr��<$�1Qv��5ZE6!07�Ռr%V��
R1������
�{m`��T@՟�I}륭�[��������K�~]Q��iJ�q���s/��~�ֻ�*����t��.��������?���0��,�y����� ���f�n� ��;��l�k���׺����F��
�m��U�u��j�d���-t����.�U��Q�{@$I�Ѯ��BhZ�(4\�k}1�_��]%0e���a�2{b]�&���<���@5^<@��wh��t���x �\��nז�-}7	X��%)�YCQ��T����һ7�H���Uf|���JNe������X��r��!V.P�Ê� q���@[� L��fկ�S����Ӷ﷨R�����x@��\ݤ,�3�c~z&�G��/Xۯm2�^�S�NΊ���<��.��{G�q�S������S1�N�~�m�:t�Jj�-�gG}���/s��;���W�h��)*��mL�0��%e�s�j�8��-��������,�S�C�("��ɕ���N͠6Pl��C�3������f8�TS�c���7Ӆ�sϦ���攋����k��|,�mt�,Ց��Ew�\�b�mc�,�H������4��m��w���(�����CR*�kRI���\��;.}K_�U��	"�r+W���Kd��*��t41/�����UXmx[��sU�eR�E�F\�)kU�5@�_��4�UQ7��.��n�������X��WQ��y����]O�7v�Y�"E�93��ۇAk�:�����zJ\� T���6h�]���[]�y]�F��R�F���������m7Q�`96V W�F�MgZ=���,���1v�c�rd�b�}�4�1��K�����K���X	U*>bv��)�_�|ޘWl�F�6�B�n�m���C�W�V�vk�N����=�U�?.�t�g��:��v���7h9�[�����jV_߰e�}p���2���?|�Hҙ���ae���ۦ�N�E���'�'�__[8���}
�J�u
�|���L�M�ɛC�Z�	P�GT�B�WG�����{�ݢެ_/P���'�s2�5Ҟ�=�ju/�i�����\G�f���d���h?k��,���8s��^O�,�kU�R$�H0����|au���͕2@�����^���ٵ:^|s�t�|�Ǹ�dWTUȸg�P5�ް8�z̗]�B�1�Y�5��4��n8��T��.���FSF��d�$ �s����{�Gw�֬����Ϟ �G+��w���ύN�X�|n��V$��8Z�"E,����<�K���R:��cRݫ�*��tNyKV�5��"��{,Jo7��5u0�؞o��ȼAf�f�TM����X�S6���B��8��E���&[�Z�߽����+	3�2�鸞T�{|�cB�U{�-�mc��8;L70ٟs���͏���
�+�l���)�����2W|>�ν�?��y� �3� L7���7`���<K� i\�[tk]������� jG!�V%n��+�1��z�	g�g���<@Aš׈��Cnit�G���T���)j �MY�[��.�;�Eɉ5�w�"�i�궝�t ���ݶ�����ˬ�	�'�e���q\���mEo��ں�(犱��s/�_ד|W{�q�e�Ʈj����]ؿL]zZvX�M�Ϙ��ֶ�w����&�x���*����2��]��rv���Ç��G�	[��,�o�q�lƌ'љBp��\/�M�5��.��*��]�]�.�X���A�t?ϫƫׯëW�MT�K��<�M1�Ta���1�%s*�̌�mb�-�e�i�k(+��Fub�<�O,���V��:vX����I.(Q��0�z:QO����:oCYI�Ju,t؟�6��vxQ��m_ұ9��� !���a�@l�V���ܹϸZL��D�(��|fkzO�Nq�HwX�qQcr�&7���R>��p����L?|�0FU+0�\�q��W���1�+�1��k���u[��[��qa�Gg�����Śi����8�2�}*�}[�_�� �Et��;��-u�*"�4�T<�-*��)�𮃵N�0X���u2�[��=]PT��_S6����\�� 8�7A!�eBy�ej�M��.�}(=�k�+����ӴF5�U\=����Gt'ϥ�x���+��5��|㪢�{kq�`�[���;�s�4�W���^w'�U�䤫�1@��`�V��,O�8�	�Ș��֟PO�<ۡ7��N}���+p����nxZ��R���/�!Ȁ*�����P�3��GrM��1X�_�YZ�b���i�Z-��`oY��ܾ{<`»�-�|x6�:{мھ�N�?�d�V]\W������Ť�Z�VL�߱�W�V=�'�j�����Lq��oϹ�r=���Cڕ����}� 0笌n ՘$�SMT+b[�X�M��j���v�ݘ�g}n)Pw�R,)��\n�T��!�rM
�U��͞��f����������|�6W��nFւp�֨���D��P�z'�ϡx+�ya���k?5�^�Њ�- �D��:�:��ĵ�Gkox�([�Uu�������_([ ׄҡ�K+W�ؐ�Ы�a�F^FJj^R�9�$b[;w���gd��U�a�n�7�8�� p���ϊ�P����ir�]�"���+��Q�:�y�H�m��)�E_�Y�� �9������j���{hK��x��V�"�x��By��o)n�{�����P��s�D�W�-�'�{f�+�	��x����k�Sʿ� 9	u}��06�c��&���^ R��d`rƞP�.n�ru�Lk�Ɩ���'�C[�JVB{��H� ������0Pݢs1#��L*�*��}&��N�Q&e�MK�����[*6��b��[�_Ltj��fC9����uW_��s�$�g�3���\����Jv��)���QyX5���ݣ4�U�P��n��r�r����@o���I�܁j���"N��ګ�_�v����E��mפ Ã����|>D�6?�Ut��̒Z����P��&��r���p7qJ74+������*`��S��R2ޒ�-:T�r���ɑCQ��M���������Wr@Z�ğ�>�v
�����y��֗\.P/�cjȇ^�j��֨��DA�Jd�Z�T������$����ؤ�A����щ�vw��5hb��To���Q-T�L����&�-�=w.��Y�h$
��:�- ����2�(����C8���{�f8��[�v(k�r,iN��������$� �;��WT����&�a��Ƽ�7q8��4l�ϸ~t����~���a2	ZQ���m�7�}ω�w~_|cs�>�vP�1�CY�z��ae�S��I�@����Ŷ�.�s������� �}k���T����b������>xW�2��lR��$i?i�++����`���#�z�GdE��!v�X����J˒q�X��j�,P�
o=���;늘J���[!C��e�~,/�Q�����\���oN�n�GLv��QbT1�����e�W��ڭ:���V�+%�^�QNq�[�hĵ3�-� ��k�{T�S@�-�
������qwU�}�5X���ƅ���P�v��+��[KahU<�^<ӥ��bT��0iͪ.�0YU5��!H��Վ��b�'���-��[��_�U���e��{�J���qQ��XH�c���+�մ�:|1' ���r��TQ��y3i�	�"՜���7���2������e=)Np�]��tѩ���z�%�K�C�WD�ڥ��y,���\O�&'�n�N1`t��X�3T*����Pg�D�9�u+l-bLU���-w�a@4�Gb��[O��"ǵi�M��(UTھU�-�7���������g�.���ݦ�1уF����5��N1k!���Zx��_B�~D6�}h�=ѹ��HS(���	��qw�9�ڞk�%^%Cu�r��0э�DJVʋ���;�"���
nn�4Z`���
�Mʪ�Q|�^����bl�oE���CS��M��|Ҭ�᥀��Z�Tk[��Z��E��� 9�]�]��Y*��}O��P7D��?�~�zВ�f�v(��|ة�a������8W@�t�2ed'Lu����j=��K�ޠ\����R���25(��T�2��&��C-�FÔ*�էBzb�o����mk��I�2�I��#d_����ϊ�V���}�53H��/<pq�{������^���+�`/��nQ�h����(`��j�Bɡj�|~�r��v����k{q��e���]��8t�h�׷+<��g�W_'��=鯣vs��m��5�m�~]M����-(H�|�����]�+w�)7
�*�V��� ],�L���8���x+�+(�{�m���U�������}w�_n��v��f����@񚦡Z��]��ޕP��n[�������P\mM��x7�w��ͬ<�^�z�1��ݘ��������ٖ�7x�m]M�ʥ��b��>ʼ��E��[�w�10�����6���Q����(W��x�͋��c�7QD�p7�.���"f�&8������נ#Hs���,ݕ^�"��r�"�������2����z'ʵ�@� ��j�[WnN俍�$�I�_A�p�D�;��]�+w�)7Tl�KC��]�+w宼�� ��J�K�Q�p��/1JXj��R��{ڳ�jxj�,�t�~f~��dr��'^��y
J���ͧ��1k�*O��$pns����#,�09c�zd�����w[�����+�Ҿ�wir:�6�2�&�4[nWyS�߬��&�I�:�����7��/1��Ų�+D���4e�lT�7�68��+�q0
 ؖ�5*ڦ�!@�s�O�u�.|^�Ua�CR�83�������ҹ�;�+�������~�ٙ��n�T�N�:M�A3��)����k��I�'I�^��(R���k� �%e;$~�&R�}�m�ٌ���L��M�+B�[)��&�����:7�Q��)ny��5|�\��k��N7L�1��J$U�sћ�Ɩ%���gܖyr�:�9E�Q.íb_�;]��[T�?Wt#ȫ.=:I�޿R�w1�U����=�nv�@mD��.� 0�ģ����=-��swD��0�d�Nt]�pc}v�]_��������h�E�e(ٞl�͐�Yg��)��u}�m�j���c��>sǝ�.����X�`��޿���@��ǀWTV�� Ce��&��oy��e�4��)�*��I���ӡ]���+�zJC�+��ݏo3Y}� ���	魘o� S˧fv��|w�v�x#��	�`8W`�M������:�!I��[�e�2Ӊ����Y3����ci�Y��3��Ԥ��:H���R;� �쀶�;���x<l��E���-`�R��z��F�
��W@	��U��C�v�i������pn�׾�۾��ޅ����~�Y�*��]��]�ߕw��B?���{r~�Q6�t�Xu���o ��]_o��0��{����+�Z��̻�Eu���� L�w��o����`�r+ u"v�A���1��R�������{��u�9����Tu����<������jEKk��1� f�;����'�=�u���8�?�����Qj��T�TU�G�u2��� �=;+n#f�u�׳�1��:�7)�A7�~pMni�܅�%61�%}�1$��:�@$O�~�}Ռ��[?u�R�T��Ck�D&���H-�-1Z�YΟ�{��'N�~]���%V߫��7)ǠA>%A
����pq��F��Ň��H�B�Z�dǉ��43L&�՘Uu~�èC䙤�a�g���x5U��lذ�� ��乽�t۳��y��2��7߭��_�i���Y��n9�in��$���L��\x�do�<y���75'x�摛o�)��涕@��ܢ"c(�������]9�D�);�%���8�(�X�P�>�N��"�s+]����O{�ls��ˀ�uu�m��g���s��2� _��v;��)9�.��ͩ�?w�ui�ׅ�%��
)h��k-7�5��l�`�����%*�Tn�2�]�� ��Md��vn+pW��;^T��TM�قjU��S�W��[v�L�`�r�ϋ�ܱ~�]<մ�Pv��������������c���(�S�O���,'�$R�>B*ʋ(��ZG�_q��i����(�NW��+-�k>Zi��]�ۇ�7�6���D�\�~�j}/�S�wc�@�/'9=lt��ѣh�j���ݜ��[��I���M5kg�L׳�Pn�j�T?-j�JUդ8(.���˟�Q�g[�������{�=e�2�S��>UZ��?�T&vI�7QnP�n's���3�����'S���K-H��tA��_�3{G�xѽ�t��{[�/�j�X��^��z��� �0�9��Jt־-nȍ(б���b�����jە���MG?���Bxʜך�
���.��V���ηuYx�c	N��P|#�j���8����9�ҭݽ��TW�z�ө��3�X ���V�8��� x�+��]ٯ��D���PQ�hcaf��T��ސV�Oow�{�^.Ƿs�C��P�����A��u�R�k:+�+�X�4���u�M-�u���k�����*Ó��g�.&4���*�Ҟ �v�u����~�X��]T��$25�_��n�y"�Ξn[o�&�+�w(������MJ��,�h� �3>i���E�s�gkr�+ԏܘc�/CB�,�����S�z���B3U�T>���4J������Ӽ>U��.;��RA�;�%���\�-�nۼ�Vf�8�Ք�XnϠ��'�;;jT�7褪Mc�X���F�}��#鰙�nc���tK�Tm5��b�mϝ2ʭ�;�$7�2��3G)ʜ�#gk+t��ԯg�*��-��og�Ҏ����{��ԅ��P������z�����T�)�߮R��= Z��Ǌ��K;*z�Ns����m��E����b���>ZR{ǽ��%Ӽ��jS��F�]�+��h8xl�li�]�ݛ�7f�ߗ��^&���ܕw�ش�8O�!$X�٣�y�ʍ2T�-�z�:����]��2SОR��~n6n�Ӳ����=���F_p];�\E��H)V�֢B��v-+oѹ�:SY���y~y[��]��e�H�g�ںe�ؘ �jڗ?����鷱�\�T��R�#�k�� J+�h9�^2��z���}��b cx�x�-���&��������kc��wP�r	���:z���>��+�p���z��L_��r�<2��F�"��*�񵽊���w��-������1����s���N���49��,7�i�ȯ�c�mn�rWޡ��fu�>f�9�[�wuF�z?�x�%�ܕ�r酁0�l���E�m ���P˞Q��\(e���v5�]}��7�Q��A;�%��[����?rg��'�)Hmt�>Kȴ���S�(���|�þc��w]��W�X�!@-�GK�-��=P,�h�T�/��֯�3�5' �c9��6%?����{�������ɌRɫ��M�;��C1ٟ���;�iݺ�!�^A5���x�0w���=�?;nѳ{�s�� �;�t,�˯+�]��f���'�䯩Q�J6��&m���t��,��Ǵ�9����]hh�\��I���<�C�����8���d��~c~���
��c�1p�n�i����W�E��m�U���TjD$I�Sѵ�j1�M��p9�����߬��9��S�	]���3z}[&ʎ�U�֒ɴ	6Y,)L���<��#,�m�`��&Cl��&&&�X	�L�,2�W�v�&�$��ԩ���E0��ﴽ��iU���ru�Q�?;4���~��4qB���<�K���v�v.uύ��Y�5A���DG�����Q}b-%#U(=u��L`����{��V���U�M�~��Vv������b.�3 �c\�q�`�)m��jB�PrL�N�5���YX��	K���TB'Nr�bS�󧓱:/�pQ�j���X����A���?��͢[j�|���1R������b�֙��b9o��&����X-*ժF~s�?�=�_���=ԭW�	��wC��ۿh
�R��p�W{&�
�&�������AT ���>��+����vb�����=������}7�~Uiب��HG�゛�ᛞ�V�Fcl����IiD����N5�J�lb�sw-����(�>�
Xv��`��2����ɓB����^��D�}��tM���wy���XU�+*�T~��/�1�|�hUw�lB����}^S������p,��xWq\؍���W�8��CV�\'��ݜ_�(e��Q���+��{\�����{��u�wPM���	5��!U���ͨ�����f)���M�;�����δ����WWby�"ѩX�vi3�kI��5(�t����:ѳ[�ՖB�k���ם-k�lpAQ]o[�j!��/��yw�~�}'O�,����j
?�&Ų�dѓ;pRj��V�S�cAN����x�@}��4��54�Tvg�7��>7ޓm:�U�	��f�VZ5P%f��u��3���;��MF'�� �J�k���c|Y�gXR��_��2��N�n)��8�w.��WW�9CKꔼ��y��$d@:�o��m�a�u��Ȗ�i��S�o�T��|��2p��J!K��W����;�j��R��{Ů	�)��b�Ϟ;�4F̡�q:�+W/e|]�#MQ4T�b�0t�f�
4�Ӵ���0<��̴�2K���g��Rέ�	��

Oi^[G,N�[�Q"�Y/�=�nִu��;�{��|���"�du���Un1�B������J]m��Y�	[@��;�V<9�RGo��A�����G434���b]�(���S��2��"�'Rs�K=9[z�O9��F�M��$UgGj��M�s�O�>wǠ���TD~y�y�i�Fb4bj��ɫ���j'��c��5�*�ރcs�ͩ8Ħ?[����H̶�[eH�E��+�4������X�ߜm��/ħR-n���Ks�
4�g�|t�<�Zo8��Dă}˖PR9�����_
f�jݦ�]���u��"��o��M���~�|N����I��9�W�1�
�z!�d�T~Ӿ�w���'7vk�]�s>2Fӕ��d���������e�i@E�SvZ��#?m��9��%�z�5�I����^.��v�D�nA��2��)�Z�4�2|��O�U��xl���==�������|�)K��s�wܷ\4N:}�݁�{˹�[�ں&�][�"P3a[T��+C�qK�8:Q_�Z�U��T%C�T�{>��܆������i���޷�����ԎT82S���ܤM�,�v�)�c}ʶ�J63�b����DA2� o��kw�{�Wi�W��;��Q_��.�����p��u���&��o:��$c�`˶�߅�:��H��R�_�g{M�P5�7X�WCy�h����++���������ڗ�B�>�Ԛҫ�9)Ճ4��
;)a�[K�9-�����s�X����X���P������y���>"�~J�b���Y�S����D�>c��?�'�cX��-�ڂ�k:��qP�J;�o����;�I�_ԩ���dMNMAYaꂣ����m�+�H&zNy�S)����,�#(l��g�w��Sׁ����jkj0�6N'-R^�8�ά���鵠Xn\f��X;t�kI��`�w�	�{�*�Z|���J��#��?��^���S�0P�UX�g8E�6�]�@W[��umݻh;��R�5��4w>e��*�LMS_Ljc"���$0����}�b��)��P�s����I�X�aZ���@U�L�g��A����9F=>H��''H�?qp�9��,]s�.�k��Ğ���cE�0��k 6�xu��4@�չeڇ��,5U��O[�V�,��S>��ɽ},MF�Q�a�o\�zO��~�g��AW�+�f������[����������7/[�c�ڞC�����eM�)6�b�b��k�N�µ��W��+1
P$�h*�^O��
tS��:V8�~�+9]�������x�>�2C�yÍժ�w�r��n�g�i
ݦ�caپ�^a���+Gpz�V���u�xw���P���j�z�ĸE,��Ȏ��gZ��VSd)Z[XWm�N�
�E'�c��?{o��ȍ,�U$���}�3������9�x���RK"Y����H�(���{��e�%q-�Dfdd�-YaK�.C����?Y	������7��A��=rG�ۭO���dgT�ٻ�]���>�6�ǂ�����^P��',�����"uX����"���mϿ��B>��n.����G���(o~F����G�w��Em���8m�q�A�'ݚ���'>��6��uD��(��.�ޣ�����Qny�Π6�D��x����v7B��Φ��3�o{��Wo6�N������nyݟy�0ѡWz�}7�U�筧(�ǧ{�mP���.���Q���������蟂�E����o�L��/z	~h �?�f�����8�4-��L��YC~�j̉�)�o���O��#��#������j"�{[4|��������'Nؽ�LSj�tYB�>k`�ˏj�WF�fV�{U.¸����p����Y��6cz�|���g�HޞҡF��_|�������O��۠�rf�o�HR�u�{zx�b�R����R�����|���ڧ��I���U�����xysC�|�aTrG��=��֤T�J_zz�{�)i��ԃ#8��;oN���ۼ�����3��&ͷ>��W�}����:/s�A�n1��X�RnY��w,�]�)���/º�x���nE6T����#��Sm!��g��cڛ����~�mP��7����l��+=�o���ɞ6��sn?���5�Վ8۟Z9xM����ݎ۽ѻC��n4��w<��mQS������E�����z/�b䛶#�>;d�F"�|m�_v��-��mJO�Y��C]�Ӽ�o���4����R�x��V0������������];�<�c�4�K;賨�������
;�?��,���7���<��-�A<-T'n=�ÓhI�|����]砋�?��9�4��fq�F�'�9i��*��d�tP�}X��E)�������O��V����v7lr�%��w��Z֣��zCؽ�T\�~�i��~�O��������j���y�X�z\�����irU��z������OA�ǳ�zj��V�u��u� ����{꼉�����}s�� �r��'���w���h��\.��uI�w=|zi�g>�*=�缜��al�����}����~_�V�{��:ͦs��q���uH��V<����⒩N><c�·��;�<榁!è������{aTm�����R�浪X�#/[��gr�/��C<G'���"ǿʤ�5S�ˡ��ǁA�+fM��E��vœz�GL�C|�nA跘2��6�+����XpO}�4Ǯ��n�b2���s�U5�X$0���Jj>6O;;�uN�O��-b�Ms�?EdlgJ�Jᾡ�9M��r���L��0�Y�ڗ�Н�ͽ&�&u��G7$>,IC�8���`b�ٳ\�ˆw���U�[*)���m�oit�fa」��C��Q�s �����F�a�|�<�uH�sf�� >>�����\��3I	�3��3�C�"��5�w�F��6ϧ�͵B'�<��A�F��NL'Σy��N����I�?">7�i�y[/T��1�ں�������d�y�����u��)\�������E;�>�z�Ooͼ��`�IZ�MS��Q\�z�գ�T�s�x?.�����vK���2���f���uZ���8?O���|ͦ�wtt��M,��5O�z��r��f7�����9�Z�@��^A��۝�_8���ɭ�{Sg%�|��%�t�f���cs5$|�����~�Y�P�}�Ӟc���Ҷ�vuw5b����������T�F�_�b�7�}S�{�����v۴��Y�+4sx�v[��n���j4��������5Q��㺬ߓ󯾆�uM���&����e�ut�(�O3�)��� 5cO,oΒ�����P�pF퐷>���zsaLo�b��^��M;��X��'3,�"�0��q�]_]�@�ie����>���������'O�e}��{������1C?�
?�3��jpͨ��2*��txΝq�Kݮ�����IN����VG[X�]�c���wzp��F�B=��̺��n�z�yF^;�6«:n��R���k������#n�8��\�QޯE 3_�������KIO�H����|8������~Z�\�e%8(�g�^��Z�k�ƣ�T��~ S�~��g�����L��Π��g�徻ͬ��=��,꭯�(�~��pi�0�{�-�{�&��F��u�8q���3�����e���]]^՟��ɬ�06GIڐ�'�����]ox�g�}��Q}������圦�jl��6GVx�a��/F,nX�k��/�Rx��*�:4w]��~�r׽����Ӝ�G�i�C��#:�M���S������Uz��E���7�u������_|�1���X7TFm��3}_��gϞ���/�#l�0��f����߻?=�����7�C��)��}S�g3p�g�������J��8�{�1��^�����"�����	���.�f�a�]^í�-�m����y��Y��m��c������=����lI�.�T8s^����^�{���c��)�%z�o�׼��?<o�����"�����NO����sA��Ϟv�ԓ�z��I�yT�o�������F�ޫwV���fޛ{��`[�#��Q�q��;�C���?�rS�}�us&�����?��ܢH�y��MNn�`�x�����@a�^�9���+/s���6u�=>>��uʿ9��|�ͰN�{�8��^�_0�!�4z2��W�?��G�=�h�����tT7�f\��q�w#�;��T��G�z���J��P�j��U��dR�h�k�bP07�����9U��rݮ�M���������;c�L�bW��7o�1'_P���g��A��87<�NLjS��FϡNp�3qк��߻O�X��ׯiD��.L�c���rr:�B�����>��C@Ux*�R��A�W?�{�7
��Lt��2��a	�~�Ds3n������rq��\���A͋��m�(c��^?a<Y�5<���_��������F�~dn������<¦Vmf��DC�yq}}E,u���ؼ�����3����3z���jd>|H��>�s	�.���yT�+�6!���z�!�%)
tp*�λ���9�&{���_8?p�_��r��,����G�}2)V�]W�t ��g	��!τ���.�e�L4��G�E�E��ull['=qRܷ��㘼��gi8�3ī��v5��-T<�W��O?������D-���I���<#,f�	���=�^�g��^���y�4�Qz�4�y���xc
�A��pl�E-nn� �B�����;��vުr�-@�-r��]�?a�h@�����3Du���%\c�Z=S��H�K��c�+cl��}��"��:'\�g0��Z9fH��)�����A���ߧ������J'5�'��hk6�}����AR���֡"^⻢y�|��y�B�{ϧg�,?��������F�,;��f0F�m0	��4����G��b�_M���)�oFf℆G�&���ʰV�� "���z���3z	�W|�{]�|z�Ր���ӳ��,� �1>cf���Гe�8{��!�zhH쯾�����[�=����k[������z���,w]��iH���7�pۤ{# x�KUY/�L}���[?8�ǵ�GDR��v��1Q/0b�G�\DfH\SA+�S�x-j�����)Dcs��|���å{�{�;�����0C�٣��� �U�΍b�(+�X�w��Kҕ�`���m�夛�x>��|��$����N,.�^W��}���ȋ�E�`A!r�&,i/[[D�=a���!6:�WQ��KOLM�W�����G�^�����s�=�~�����o���w�v�x�~~^1��k�f���X<x?f�����z�8_���a�Ӟ�(�J�ȡ�rn^[����k�m�܎��xSb�,���r�U�ł�)�ю�a����y�������7�\}���Wn��%n;�'k��Ɂ�V�;��*
�&����������`�T�@ct����~�HXT��'�I՛���#��?������~cb�˯�L�~�m���/ҪV�\���,M��G���Ѣ�C+yäf=�y#�Uk�
�zo,}��#0����ҟ�������n8��;zV�d�a��,97T�, ,�}5~�Q1���p��ta�P��Ͽ��~��Gz20d��'f��D��;�;=�z^����� qXsQcq�p���9ɘ� �W�S|_��z8���y���(���]�tc����c�7!E���nQ�����v�M��n~������igd|�,�����hQJX�&5�1����߽P�竗�hH��㦓��ZW��7ǆ�qE"���,����wڒ�jF��.0����>���������?�����_�[�MծA�e��[�sw�9_r��0I��df�&u�1�m@�L�����??>�z�����!����em����?�dx('��Ƈ�?d�O,��߸�\Px�+3���A��J�Sx�{�f_�|�dhT�� �蠞�8���P�{����(�İ�i;��\s����ǘ^o�ـH�IV�����L�KX�ϧ�"Gn�)�H\�m�V�I��nL4�u�ɤ�jɥ��
���Ƙ��zݼ~D8ú������F#؈�b��8�� ���#�DA��a��
��>>�n�?b���_���P�;�ϗA�< �����Ϟ���;]�X�s�u�Bp�|E:v�{JT�MXc(�Vf7}ds�0�B�R�H��t�>�oY70���'��B�����D��^7��Ճ'r=��y�Ϟ>K��?�K�4$$�)Żc�Ǫ�	�"�))�$&��D���&3&0eNiQ�-/��씆��?������ﰽ2s�'\�oa�e�`�������I<Ԟ�]I8�Y��cc`�ױ8�m�Cn�s�EU�;���X���-�Y>�G~bP����
�k��$z\#�[R	�玕j6�`h 6�79��\�{]ǙI�q��-�\�$�msDX���iئ�9���?��������Y�~���
�'Qx�����������` ��c�0��x�ѯƀ1�_��(�����1��h�E��&c�W܄4x�aϛ�gPs�ᔬauY��j��`��啛F���?��s୩�^:��`�v�eZm�L������l���~����eڑ��%=�� ] L��2}^w�髯�C�]Y�9[�!����O��'O�pa� V �'N��"S"��bc���jؚ��xOL~,��u�]�p��c�k?��sR���>xh�=[�/��@Ba���]6\�8�n�-���l��h	K�����NQǛ���_Rm���w���\��!�C#K��ե,\S�<C|O<����9��y�����=����#�{g��9ܸ��u�T<Gl�q;ZYi}J����|	$�K�� !`�U� ����	�5x��&�=ǀ{�� ���=�
����1����_չ��v�y���`�F��\"�!
95�Y�A�j�$�W���Cg+o���7mش`N����j�w��?K�[vN\����zɭ�/t���8����gj-i��L\����_XU�&�,&]��W"���_~�%���)(p+P�~���:i��=�yUB!<��A�I���9���X��0��������������T���q��4�;������=�0�eK����$^���yY"m���@�-��/>oz��O���_��P;"a}�6V�/���H�����5ƍ	 �О�?�����'�j%\z����_D 0�0XJ4a��q�0Ѩ����׫����� #���"��c���rS�c�q�\�y�&��>7YQ��]x�8��:��,�M�0����?�0�-9\�)I�׿��B)��VX�&Bd���v�Yo�^��B��;Z��ciB��c���Vӆ*/�e�A9��ӖIf�I3:�D�a��_������äC������8}��W���G\�=8��K|��9aKL5�Cu���X*k��X`�d���jᅧ*B8�Ғi0���0����\��J2R��u\V^'�c�R����|%���Y9��c���m��Řk����f�Ɓ�a�L_�2j=S�$�aԨ��d%��lcv~nb8�`<���S`��/�x�^j���0Ѹ�DUK�̼��3@(���%B�hK���x�	���0�L2�7�d��ܼs�����,����py���˚+�ȖPG)clJM����ךQ�o�mx7KO������[֜B�e���h���o87��O-��Z��T�bb)��+��!��&\u����p/�5'9I���+�׳i���p�y���^�BQ�>�±pyv�6[`􌧦���98�rx-�yM�j��aW#n&�|�ᳰ�.�W#t��L!��둊�k�[c �]���?{������1X��R��P�z��D$\"X������Բ�^�Q�4�0T�����\���@&���܀(θC*6ʕ-O3�9
+�n�(Xh?]
E�����s��0ϺF���s�3�TMᵛՆ��7�'<�z�(�������z�<|`	��c'�츪_��wk1��Y���W����w���� ��2h��>=�q�lj��[^�%S�Q�����0��a�WB�I|^�߱�T>��sz3�X�Gs�&LD�j;z>%���-ѫ�^�����2���L�4��-|�����{z���
�
��}	>�}~�%'y������C%�����y�ej�m����?<ߣ_�
Y3�=��v�؁������48V����I!�M��mYŰiK����5+�.�9�4V�_~���6�'����?���*A��oA�Qhs����"��9fJ,*�+&X�cl�*�&�*#�Ǽ� St��5o�@A����^��Zu��	,'�udF�폃����ti�?���y�o��E�!�;Sy`h�9��K0�L{�l��%�܏�h�<0 ���f�'��h�@��6*����Ù�Jj����]�+BÅ-����B�P5lQ��4�[�F�I�k�[K���`��.� -�^)����ҋ�=A�A=Y7�����c��K�����K�xg�u���,���LB��~���}P����k ����㹣I)��I�KVnz�ST�6��M#U���_�A&���f2/T���6H1�v���iqf�9_&���ʩ	��Gi�{�z_��;��-����X2�W��L�������uz�t�~"�GU��^2UX^�j��k�߻���M�I5�ww��?e��s�^��&�7=[F�m3�t��Bj���� �#��0{ݺ�sX0�h�u��sd=��g"��c�h���ł�|^*����:�8��h���YE��p/�Ax���
甇jB���)xh
/-��^49�9�-���QX��q[/]�XR����?5��!c!�/b�<��QL�1��qn1��+��1�l.'�d��
ùu�*�Hlʗ�v�`��Jx���+�&�6pN�:b
�ձp� �#��!��>�u��.J��e�=J��:y� ��|||7`�j�A�w`1C5�F��&T��jt�t��/Q�!0���N���滢VY��l���S�a�-�2B�[�Zۤ��GY����%�������ѯ�a��)Iٛ��<B��ָ��]�a���w��S\ST���c6O�;1c?��<��2�T��=l���F(�K���e���k�_>'���E��G(#��c�L�ƽ)W�@n2��`���rS��U��	�uy�+�׼�Ss����^�~�P�hL똁�ilې�u&���@X��a���c�q}G)�c��'w�B��uI�`B9]��m�X�ţ�7�+6E�cD�	��P����i��c|�k
�\s\1�8V{ƣ%��:���&C��?�`,<{���L����o�1����m˓��"w�w��X��/)u��S"�yv�@�r��ۭn{ngLU�4YF[}� �D}`QXL4X{˪��S�)G؂y�?��?���;&��e�7Gkð�xpt�"���e�3�0|,QD�~��k�jE4z���ᅡeߡ����������U�:�B֏UQ��'�/G����A�_���X��JzM�+�
�`��i�'���c�����aQn$m�o|?d��A�k�Z��<|h�5��q�HO��q\��3W/Y|�p�<~�.�5�ѹS��F1��z����QB��/�(~��VfjFW�_l�ڰ����+T���Z�`LqfH<�����ƽn���Fԅ��rl|'l�=~���G��\*�.�������<�"�Շ�'��pؼh�i���4���\�9�:�ՏH���'��!��*C|ϊ__^��9�e��b'���aF�J<��x�"���?��~��Ɨ\H�Q�w��p�2�L�L=qa^�5'�UI�+����)mcL�_PU��S�w��NW��ΐ6y�Y>�d���D̗A}�8��M�ӈ��!�]ֹ��������Gt1Kss�7m��H�2DrN������(���k�4��`5X��X����dq a�����ՠ^9���̘��8X�����%S�8�}O��Ә��������㨀y��@9`�2�>��fr$��F�.�#�Ӧ��'/!�#B�65l#���2����7m�ھ���{8>�Am!K�<��)����i��f��0��'�D� ���X0J�^� 4�����Q��']p+e�-;������뀙�=۩����3�w����B��D�hU�Sv��Z	�d*Si��hl��Mň�|�4/mZ�^Snp������+�W����01�r|<�pT�	!$� KL��T��־�/?nZԤ�6]j����.��b��~V�M���X�6�����)�y�J�`,������_T�z���Ye�G�p
Ci��a�,,������ɼ�✬�t�$�%�ګ)��K���=���wf�SQ]2COm��]^V�?��F��b������3$�6���R�@�.~/aX9M�n��>�� �_r�S[��=�8B�;h��cz�;]�K)3����n�/%Z�rB֝���=x�_~�=d2���?�^���u7R��D\��Q~h��S���5�Ƴ:юhx��r
�!&�y�V������k����j1S�=��Ő`���e�װa��l�6UW/#�����<��C�u[��)ϋ����dښ����	OL�:()-��H������qN����E�gu<���D|���?2�"ã�F��o�!�FU8�q2�����%��V��/��9 ���6O.�`Cx{xp�a��r���;��h� �O�<��o���@K,��"uo���xs䚺��v��:/�y�y��VJNf��^�Zb^j�)Yٕ��{�vB�������w�I��^lCU?�i�`-P�����|ݵ�)S���TR���u����V4���Kvޘ�x���~K?��_�i��������2�����/>�q=��L��&w�����e� �X%����)�d��}2Y�������;�b�b�q;v+,�s��z����i��8ۜ1�0���x��Yҳ�=޿G��<)|=�y}�BQ,�/���%}�h;X�����(W�jK�tl��x^2�ta}x��S�j�xt��s����؇�A8�ͩ3v��P���ā�M��Dc:�1=��0�;�W̚�p{y��U���'4����6��g���%ꀝ&��_���3�sK]܁�ð�Gׇ�ދ�]� �W�e_'��[z����i�O���[:Z�9��7�x�F�b�R�//������Xˊk����a�:v�PU�{T�4U���hY�L�,�~�P.�� &: ���}CmW����S	m��e ���>�ٷ�#�+�Ŭ�L�c!~�ヅ�����3�Y`t�u�^��F��mY~?���u�rI.�`��8��9@�◟~J��h�D���s���a<��	
%H�}��W�ޙMH|6 zx��d�N�i��|$���4�s�Y*̎J�j�k�aҟ�;cu����7�'O���T,��aXׯ��уtV���l cs�vOc�IM�`ax��_�����{>_Ђ`x��l�\�7x]�U�AA�F��_�W_~���z��at�VݸhLK����RY��J���//�Q�cl�,��b�hy��y5�?�s���Ͼ�A%��R0��_�����u���dҋ���/�-*�͛���`� ��ōцJH��iQҴ�`��"yz��G� �P0���*�j/�D��5��LD���1��q.1���=�ˋ�.u~-XW���cu..�����g��չ�)���K�"p�^��̩qg�(��U���_�ǳ���:�j�w��%XЎP�����dPs`Xm)��%���Nc���<��◹a�u��ӏ�_��?� ��l��% �d���&?G�S �S��5���=�k���w���),����1h2C���������Q��S���?t1����㓓��&ݘ���2N�N��B�//_Z�Mz\�u�d����/�\���zy�0ԒS�v�yy�ka�XH/��#�|�勨Ȳ�/6�YI�n��v@m�w��M��hwu���ю��M�ߝگ�(�Q��{S�S,��W�=gB���º,������������[���ٌ�YD3��;x�e�),T8�哒j�(��yV2Өw��F�{\=kT��`��8zV�[�#V�Q9*�(`�g�����'��c�q����`a��t�<ej`ۀ�����i�	%0��ުK����,��|`,�}���3���Tm��o��|�O��*��A]Ȩ��p墏?������aЩ	L
8W�XW�����=��{ϑx��C��k��;¸����b|�՗��;*M"I�/���l�WsN�d���z~� @H�٥��k�E�� ��e�[M�,�!y���v�R���V�C\gL{��w�x*ᘺ��`E�{�����Ԝ..�K=G��f������aCٹ�H�"�C��ί���:cU3(*���e�����e�2�ڄ�}T�L��V�J6x�S���X��a�T��/�;�k)g�|,R��N{��\��Kd���vk�mЙ"ƙ��vg�Ux���#�I{@��9�����; ������ow��1=����-������T%��(D�
2�����?�Vp_�u�Q�h8�)�crҳqI4k�'!��Vn1q��hR�ĔZEC��;0+@LF�J��FWܧ�p] W� y��)�mqRE�R֘p�, ��T䵾�r����H�q,d|΃0�܄dp�`��Hz0�W=ug�$)i��M�>2�=���Vtǁ��}�{�������j���:Y>K����5ϓA='��m���Ȏo�C*S�d�3l�����j�a��1e�owaр�kO�����/`�Әl��{�����5y�H&}��~�d�����Rl������l�V�[n�k(��1$7�[BлO�k�!yEW�VX�`��9W��b*XVܠ��{��YMɩU>�-���<T�o���n�v�bn6d;�JS�߻ʸ�U{��9��{n�pō�3ϒ���V'�v���IYn�{�΄�����ghl;�����ڗe�%��ٽj��Ym<x�x^�E�1:��"�#��U/0���x�ꝷ8�"&���Ȉ�]�$����◄�KT��j�HAO<�'������Zi�=1�G��W�Q��uS���!c�1����ppt�vV��=�z����lhC=wP�gV����˦ %���Қ��d�y��C(YὍ����cc��q=|� ���צ��T^����:X��0Γ'�'*�369`�,A�a\�\�f��m����Z\��1��^Ub��vHȋުs��&<M
U:M7���
树��!(%����f,f��"���!�bP�0�����û�-� U5��p��T/31Jv�א�����ֆ�������>�ۙ�@�	�B��pD5�S)�,%�WL>�����bY���D)�1�-N&�<y�p�4fR�����B�'/��:A	�]!�ra�$Ε��J`������o\��(~��\��{��coܧ*mZ}R��Z�=V����̠a�ej��+�� ���RGM�X+�Vj�,���&��bb�WM8ƥ��"�P��8JT�y�4�̬�ܛ��2�-�:��|l�.�훈6-$�pM�|	���^�6]��1�;:���@nr��Oη.n��^�a+��&��i?9�P���+�?⣞�_f�]?��5�C�@ʆI��{���ѦҊP$�n���hשKP��:ƻ�hcƷ�zO�M��},)Ռj
#I����]���ɝ�s��{�\��^b�|�����ce��:���b��6x�����KR���?l�Z�Jo�&��ݴ��������������*���p��$����C��P��n�Ņ0��Fa= ����y蝭�b�K�`PqQ;�Z�6��F�_����yBp��Ņ�Azfz�mq$[2J����G	������FBJl
�@9�v��4N!ai�k���no��1oe�o��rx�}_����J�I�J��Ӭݢ�5��"�`�ޣcoN��fm�WW��r���7�{5��v�q�ҍ䞺�%f��� �a�
�^����ƅyڪ��xN�.�K]mN�5q��}9��!|v���;W�o/-GLחo�d[��`\?lO�[���i2�&��f��\�[<�B��*��`]=5!N�g6�h$���fٱذ�c�-I%X���CcǷp����RO$�>Z]+�0»��:Kpx���ɒ���Ơ��=�R��+l �H�� %���Fѱ4|xhX�ye���if&�S�y�̕�q�9r�s&�����ٮ�P�Ia��bs��эtP94��	�K��
0��6�60I������L��<���<-��d�K(껪~�u:�6�<G�)�З�ð�<�n�[��KS�R��<���Tb������`�D�
�L �'Cʹ�rYB��Ґ�[F-�Kһ�ǘ�QXi*ڷZ���lv��ٶ'y��{ߴl��vڼ�y��E�:>l���94���;~W�p򄌅@%���idm+��]m6iK)hE�)EX�5��iL����N��-t��ӄ8����Ƞ��n���sṺ���^��^�)çE���3���$ķM���:� �i2���B�kq���UC���Sd��1uI/n��\��o�ss]Q��R���C�sygN�U�$y�K#�Pʌǿ�	�E�!�G�3u����߱�險��%q�+Fl��N�ӡ�GԠ�!B{ݜ
�0D҇U��0^8�>��+
�lCi�X�l���)Z���؛��ϭG��i�SҧpX�Ds`X7�0������o����E��ϛ=d�Xtє�t^7��5�ud`��,�SY��Vݿ��i�G9��9,�������fY���S�-�c�zC�:�։�u�!�����P�0�T�N������}I^jx*q����d6â�A=�JL�Ͱn�qk�^�ȫ�	?�!����@#��}��.�)ş��L-uK6��^Y�%��Z7VA��ܱW��؁����'�}, P���<A�����3X�:�L�77���Ux�0N
��Z��n4����dI�ŵ���{��(���>���M��Cv�z��w�� ��J��9�Z@�:Cg ���)7�:�j�>>>�e��x�~Y��!�i}�\35����Q�[�u/X�ڼSa��ԕ&Y��qhÏ�K���G�c�D�su�~���21�r�j�Z4�P�639vmZŚ��<(
(�m.ESn��$`'�ɓ�%���{|X�T>����P�[t
?f���)�xȼw����i`�#1����E�B����|++\y�悲��u�X5j!OT۷+v���g8�І��.@�6(a�wH�EIJN��ʍ)�db�O���wjj�/�ha�7kk&�w�D&m��������~��Q��o�}���oz��q:���cz�2��c��0hC���[�"?���'�E����ƴ̗�I�GۨI��O�׫���VF:��`bq�"�r�+�=P�(54�FI֌l����Ҁ�M��Fl�J5�R&����IW�hOf(�!\M������ުA[��0��h-�I}%����_��'{���ug0�.Z�� �E�'D���1썦]�NT��]Ģ0�=[ԏ��z�C��M㺸'���y�J�H�L���>ΚcbT�T/�xfJ�!헇�!E�;:�D���1���I5�Sݵ�J�I�{�Q{
�3G߽	��.��k�.EZ�j%�T�rd3��8��?3�!��o<!��H<w��P�b0,qE��x�XX����I5�/�����M������]o�DU��=����jY)t���_���a�}C@#_ޓ�؆a��|S��$���˵���1S"�3��H���ySfD�����6Pݯ�Bn͋�"�e	3ۨ%2�"����{	b�Q��N�	��"��Mn�S��`�f�LB�/��X�Se������פG!��g��"m���N��g�,[�4u֕8�����f��*�����e}�n0�8�x��i���( ����1Jȅجl������_핹x��EY	�H�ǐ�����Ƕ�������ݞ��tDx������	�%�O��μ�$�R^PK�9=��հ\��=���(2�Me�)ݺu������X��r/W�W>�e�������'���I��"s���7a��p���n��%�0�li�5��5��_}�T�
���5��]<��'~��ֱ?�Ɏ��{_wc2db��#�=�Z���j�i�."_P��l\[�0[�O�� ���~nZ�֒m�Q�sa/U�P�4zE��'e�@v�}T�)[/�-���Pr�Z���7Y5B���'2MVr����XR�I�V]�҈���ɳ>>��k��'�;�o���� L��lp������&�Y]��K�㫵]���u,��VR�(��]�㡍l����SDtL��(�t�RyO�{�m��mc׿���ν���B��z�~9�͕e�"?���-�KC55|����rpA���B�0 |���yzZB4�������$nUc�)$qx�E_��4-�1y 8�*S#1je�#	�Z��	��<��� f���`1C�P]\ס�9�����Rj1�EKj�/�c����d�ϯX�{���$�#���(�X�U��˙[�Q%���lf�s:��YĀm�H�x(�0���^��c�W�w]��2u�ۺ1ϱ!2$wc��17�c���3ePq��DQc����Ӕ�$��n,�g����j�������0�d�f�3`Z�u��^SLi�M"1?W�b��rOW���2h`pn�%`'��sN-��Rf�I5�!,VY-_��s3�	(�F�P%Z?'�i1a���#�e`��=���ƍ*���rɼT�%cQ��[C[Ϧ��*gz��g�Aw�q��<S$2Vο�N��y�1pF��?{�%<�����EV��M7v�9p^t)�ƨ��o�ؕ�o��o�ۦ�4N�lN�L�&,<kL�c����F,Ta`���V�L,{]�K���� ����� F�c�><"I������~�S
4���$�t��x��6o���6��I�J�G;V��~S=mz�G�������{��'0�8�GT�$;)Ck��M��sPsr\�L����1��i^'͓��o>��S2Jl16�gK JD:x Cm����	\I�a~��9��0��@a�qhדE^��j�,�<g+�\0K`��w��O��(*�7�Ӿ��At ti�4*/R3X�l���H*^f��:��\ Ye����0�ĉ��H|/���jMC���HCtv�����zv֊ow�����n�WfLGL*�l��IN#� ��@m�Ou#<M�?��P����$v�s�n��+��2� F�!-O�Ce-�`F�X�'�s?���Kb�P�BH�Ey��VgR��t��xˏ�>�Is�q-J��3՜�c�Y�Gc7�9�o�6M���K<q���*��F�����J��:����.�=7��a`vL92��宛�h|���I+*�*���!]��m��7���r��N2��Aul���T�JN�a>���0�E����q���(³2X�N�)`�G���ث�(���w�Ԏ�S*�-w=��޼�KtȰj��KqzL���/�/er�� �j��h��s��8�Q5k�L�䔡��jp~�����]X`�ɯZvz.N��1-�)2�2� ӹ�뇮S�\Z�ů����LA͒7��P�4�%F8���z�_�����D�cQ»���n��9igX`�!erK���+4$�k{�LC�sx�2�9�������^�������d�g���|H6nw���CiqZf��\ul��=��T��#`�kOD*4��^��m��H�*~O��c^�fLo���Z�R8?�|Wv�G�eH]?�6!�z�IH�H^�p]nHN%�1��U���׍��I����z|8����� T&ү��U�D/Nᏼ&*C������u�.�ɳ��ؐ�wĉ����b�j����C\,�(W��ʘ����Ư �Li)�1oKB��
�S��-�-^��� 5�_��6��S���#E2
	8��ٳzo��M�����Ɣ��� c
o�����i�徘��9�0�3��skF'�;�fKˁQ�qtx����h�%C�Ҷ�q�0
����7���X�&S3y=�U4��!�h�Z�&y�s�եl��Mx �x�Ba�[�j�l���� ͞aO%6�my��'D9+��jq��Ql���~�[���/�u
�x�nu�VY7�x�NY��%����9n$�8��X��)��$�o��ۨ48d`J�[7S�%�:qP�@8<?���]m-T��Y\~���b4�b�&������C��$�[2�l�*R����5t�I")^�\�\��{�����]�veZM���.±2�w�����K���y|􂯣�
��eM��3�������C�q�V��xn�k�)��s��ޙ����LP�]�!Ef�t����4��,� �1���Z�X��||a�J/!���"���e�Mg���������"�[��h�h��������0O��0{^ +3�r�J�a�J��������ئ�k-\l�E;��c�V��m�1����T1C��-!�>��:C{X���vDN���J���E }ܽ���JZI-��J9v�ɭ�-�dFŲ�r��z�quf		'�_�t�d��/��w}'��r@�k�g���&~���3��=%�Cx^�
0�y�P������F9u���"����<� L���	����[%%�3�����<QЦ����J܏�L �J*%ON�Gn�E�e���w�X��[R�,0�P]�j�k^vNf�����x_���������fu�l����}q��X��.����qC�����
S'�n����)��IA�'қ���1zYID%�0ඳ%k�-�bٵ�ν�����8SG/&�2Ĉp}���������y����Q�G���*�K�{w%��[Mwn�4EF89:�-��Di�c&`��#��g7dj1�����u��D�UYM@2V��k��i��I���M�2�ϲO�ʳ˿��R~�!�X1��S��z庬�������k~`�}�
x���c�=O!��:��o���/��~��jV0@�nL�,�/Kh��+zV�w�FQK�F�vU�<O]r�]ѩTZ
�r�j ���Y)(6
$����!�����`<��Jt<U��Ū�>%6;���R[�!�KP��&B>+��p[��]Ɔ�_�q����،/����
QFO�aSA��cks����vЍf�͆�כ�g��&�SW̑Գ5��Y�hB���6)�i�/B�r�[ݑ��}�1�����X�Ȃ��!Ns��i�A]���D%�gϢ.������Ⱥ}��^o]�ޒ[0����R�׀C���rHyV��	����y�����5,Q��ϳJ�*�/��m�.�Q_���M�{#qǢײ�w��5�}�s��a��ӧ̔��\r�oB���F�h�^A|+)�SU���~�)Q�M���м�(E���)�<q�Y��ݚ1���N�!�n�k�K�X؎q�������yB9V:�G*vH\��	r �f�!���9H�*�X�*��b��ۀ�w�f˦��>����q�1O���� ��0�l��<٦�����i*�L��o^ɖ��V�i��e�WYuaG��vҾkcќ�T�j���p٧�|uƘL�Ą���#<���.��%�T/�R��՘��su���d�*<����ExjJ��S�����	
��e����<C�J�Q�����k�*��:��D,Յ4`X=z�.��G���yV=�Ǐ3�3�&���mh�:ˁ���˶��+�������y�nLSK�L2���Kd� ���;�G���mF��_&zp��Q��9���2|.ǥ�g5�33V��9�*�@�nOt.� -�fΐ��������sn�}'i���G�3#(V���d� ?�d^�e�EA���W$&�<�C�׎�S�/�F��H��$�o)�7<G�7K�ۢ�eLEYi����2�����Yݦ9�x��l�d(�G����>��F\�䋃��j��%�ϋZӳU�>!�h9���짦u���)���F#���R��?ϙ�3��i��`�R��R�_!Lw��)S�BtM�@#ڬ�J
ڱ�� ����z��Y���M��u�"yny�m���?�΢{@Zn�s_�SJ�~���Q�+J���I��9��O��7�;�\���.�;�tc+���0�x�57m]��L�HZJ�������ͣW�Z2E)���*%
X�z���7��+G�v)C%$��O����ĺ]=+��Q�k�@s�=�;a�|���ߛ��H��*�S���ƹ|�ﲞ�H�݋��pW�ǘ�*" X��w���d!��Ah�"c����O��g�����w/�p�����}�b�����?#ކ�ޡ�0���Ķ*Û��A�}��:�6y��L�j�3X��2�k�dF��I�Q����	r ���YuCɻ��jH�alè�__�L/�� /C��jt��:�%��(Uw����;k��"O2�-'��e.*9ԤYF!Q�8䀏z6�
���d�G��J�E�bI���Ȼ�q���Hv�?+|�j ����N'~��摧�L����)r���F\]��D�ֽ�9~Y�9��W����I��!|�N�
%�!�V�f�yl ʁ�4��V��9�JDC���+���0?����ߡ�6$À��6���'��dǎђcy+`�7�K��@ļ`�\ph@�RY���A}sv.�°���Y ����c�6�W�L��R;�]�4w�i�1yPCN���{�����嵵%��2�$Lcҽ�d %��Yy�o=����O�s�"l���pȗ/���'O��\Hr��	�/�0�ae&}��S�w�~R��C(����)�7�(m���(��N�CbF"j�ih,d���6-HB��r�s�C)ј�N��Ӏ�ؒ��n�Fq8�-�6$C��1���%_�%y]m��n.�k�x����엋�>�ב��1�^8�����JTq�8��B�x}^_W�?i.&�S����k��>}�Į{5�(aUC�k���{�X�6iܮ��$v�ZEI�w�8�T��vrM�c�������z�����AQ�a���H#�8� ���z����������}@�zAg s�G����D<広�""Z�PM�֤Ri�J"sۅ��%����X��n�%�~������~!���X��*p���t����b�2+�a	�`��UA|�ѪX֙s,Rx/��8��\]-u�(!������>wa�_��XBcb��>]�X!�&�H�}����M�`Pa��8��h�;�G��
��8�{O�`a�mYj9�wl�c#z3��g
����&������~���r4�Sh���b���őc#5U���G��v޸�ղ�}j0�0F7^)7��`N�59�Ʋ+&��:�h{O�U�mo�7������N���zf��VԘfp.c�Ę {ǆ�β�R�8>�$^�i�nPw:+�q@�3	%�p G�u��Y	;�#��54�c���c�0�;���+��J����g�fw�0'��)��hD�=��f�Qda��|!��R��U<[Y���jod?���Ը�X��ü��e�8��
1"\�7�Z��� cLP���ϡ�����ie�!���o�R�S�x�ko��	zU��N}J<n�./7��J\CjF�[iL��:�$Et���ʵ7>[;E��<9��m����{���{xX�ۼ5�#[a�a�����#F����ae-S�'�L_�U�y� �0�1��u]x%�6�P�V����']ڷ��  u�IDAT�mY�o���K^�u��k��'kkJGLy���9gr�T��}�5T�i	���J�qt�p��6��D���9%�u��}���^�5�sk�b%E^�7��6P���6a�Ѫ�����n���%07¹�gƆ����R��M0�ޱ�[4�fN�W��S�"Ӆه�\���QM�/�uh����1���(K쇭�.1�%�]9��n���1z&IAi��j'�%m�5��Ϟ-�:��[O)�a�� �	'(�����K-!a��UEȞ����m�ZOsQ�����!��E}���}��
g��h��8��QQ[ �6.����,q�-�b��rN�e5.��fD7޽u���T�䏦�N���~/�E/�=�D�����Xvp�s���3�en�����#����$W��w��6�K�!�pɧ�s3<;��MT�tU�!�;�J�u��rcqX��3��K�=��0y�ɡ�����_|�%���dl��m�mj�|��.�E+�"�tq��W�q����b〱D�j��FwS����7�>L�]!�./0D$�X9���e����y����E�1�2���T�%.z�v�����.t[�T�#�N�3ǋ��UkEl�L&I��n`�V�'N&�D!3����7�K���l�c��?f���w}��M��=�[]�S�Ғ��|�����$/f�6g.Nqf�^转��U�LadI�)������זD����=�}��w\K#��"�L����xڡ�Kd |�/b��I�S�e��|Z����CR"�������[�:���evHu�1%�=E䂤���|�����?<���_,ǵVݫ�� r�ģn�Nɓ�1��m�Cr����,lH�B�s�>x�0�d���9��}��l]�1̓������g\^���ǕS�t����H�wڊRH!rsq�X��al%���U�R54=}��&��+�a���q|2�J�qc�ia�A-|T�Ju�b�S��@�:>9J�n"0������lB��3�k�aW%?^&4R
/�	/�Q�_����
��z�-�޻������(�')q
}G&�<,�R�����'��ʦ���DWTӼ�J0,6���]�NJQ�r���v2;]�a��y|p�X�6a_vu�R����.ø�Tm�}�ҿ���T3`��W��i�u��_*P�����v����g�>K���?�����E	.B���<NW+�L$��7l��a��=8�T�o�n�g�~y��^�y96;�����pup����ztie�`%T���ܒ�����;�x.�Ga��9����kKJa~�S�>SS�����A-���q�����bg�`ebnT�w=b�������1��n���-��m�C��� �E����;f^g��'����ⲳ�ȍ <N,H�Ѡ"�c��\�C�yժ�f�l1�SiF�j��J��6&h!����"�f�W�:,�|޹-�}��7�SRk ����%�L�`�.�a�,���7o��^
�F&xx�9X=��c�릑�����og׭M�sW�&�u�9ځ���[K	.r��c�x�:�m���!q�u�8�ǖV�A*���B�~IC�D����N����~���K����O��)�c��:�U17�a�)���M��YWn���1d���ȵY�񁎥�w(`S�V/�/��y�������ŭx4�s��;wa�t�u]��sD&pV(R��M\�a���?��$j�>C���dE���+�"�]"���a���_�_,B�n���qgJC�C��ݚT�:1O�����w��ێ��� �+T���P�uU��a��*NX?�
�|Z'�#�u��ȣ#�!^\Z���ΰ]d���pY���{�
��v�j�*F���?YV꺝;�lyRcsD�`�X�ֆ��1�w�wZx����x��zh<5�w������ߨ�[7�S�J�
��P�J0���R`-?ʐǱmt�O����1U
c���z/[Eqý3�ĩ�3���+7x����EQ��0B�����y��O�)�qP��)p,
��/.:���qx�J(i|a��Qn�0<�:>�i��*���O�䚒T��@Kc�-� ���"�C��R�2�����8�t�$W����5���IT\WZ~�,�n{�zWp�3�Ɇ�=�1}��j���o�!B�ao���3ǲ���/�=�1��Ļdz��!�{w�s$�����yP\Ҥ#Mil�E�ڣB($�e��?qF&1��e�,X�y��K��X0���#�V�]�~1"�b������e���v�3WAwṡ�^݉����?���{�A�E1}㝶k�F^3^�[ꆑ�0v�?G�jI��`��^�m���gw]7�����Y�Icؔ������Z��cC�a6H��3�Ք��I"��s������7��\���O��Yy1�nm�ܼvË��#���_1����c6�$4�a���a���*9Ĕoi",�ڢ���M����GMކ'�$s�)�PV���8�@IԹ�ǃ��b�D��^��]��#uc����_||2u�����; mhQ9���$���i=���CR	�ї�_��]-���J
��<s!��.Mm��	�X�]��H�",��93Ϯ:���4��U�X�j�Ke�P���?�Y��\�^��W���W�<��D���<~��]d�'d�'f���	s�5������{�m�Į��h9GG'4R(��u=C�Y=4.px����bj���7~�iP���h*�kh{*7�QEf�}�ZD،^"�Fc��q�26���]7���S�m�S_WJ��_Uo>��9�x[�^I�������ù��ECG-$��8Ys�~�����ϿDe柕���([�36�5Bq
Qb��Z����qQn��wx���Ob�x� �@~�^�d;���W^��]M��'/����S�v���a�)T
\z7��T�.ޫtF�/>>�Z��Het�e���-+�E�W^.&/k�!��6}���ߏ�2L�Y{+k[eS�G����d�V�V�-y=�	J�P�)�V=���5���M�ަ��j��ڽ�S{�ㆷ�P	�*��;��<cѱ�o&`U1�/y�Ź�������۪�ۺt�M�jvpr���x�ɹ1�OaD�-�3��(6�.�؏S?��[��.��c�cb��e(��8��sqW^�i����3��^["Ί1�C5�q��:~9���-���B���&�w�9�Wt�!0�]�&�/����WUn5�?��on�8o\���:�	�Q����pڋ��_u-
�Z��5��Ki�R/,񈹂s|V=d�?5>6�r�.�y���+W�W4]M�C�;k������Q��g�������Ŝ���c��P�Bo�=T���Eb?����M�����-���u�H�xHF@����ڥ�^�� �y;��T�]`_X Z����K921,�����S��b�n����;7FlO1x�� ���k�}�Z3�� ���f۠�`:m��ګ$�XK=��3�ȣ&L�P@T�̅a�zc��V�Wz�&�gL��8
|�U?+_X2��T;�,�U!��bF�ߟHj�b�LM�^X(z��ۃQC�¤�y�(�m:�X���۰h�ph�}���#�CF�T���D�+��6�j��񔉬�f��䑅�
�cEDc�U��Z1N����y����\��ʐa81�p��g����M�{==�e@A�/������r8����$ab�5,Ugޠ���Ko4ǺV�%��ֳ�TO�f�����������a��s(��t_s'��_�T�¤��d��>���A�����堓m<�b!���ρ�!��n��N2�~�H��
��*\�k�k�^J�u�]qIYai&0��عOOΌ�rte���{8)�R����>�yW|=8�_�5=x&�}�  �+��^F��	ҮD�8��$�ܳ�"���[�����,���`ԇ�<N���+�q� JB�n�F� �>*����d�uLe�六ʫ�<��n0H[t6>%z-��q�Q�9&n�+������*��&�2N���sv��Zv��k��>�o0��4h�^�R�+ֶ]��T�f����ai���)X�Gy�������ֹ���]p=f��c+�H�;xg�q�_�J�dW�\���'�ކ��k�X�c-6��D�Y��9���(Rɭ]��%��>rRKD)(Y����8a�o�c9������M��8�/j��p����a<����2��/2��&㫲%��B	'7��������JI/��;�0�\�$���\��t�x�� ��z��٦���ԛ�|��hܤ�
�g�O���ɓ �t\ptL�3��P�hԖW�!���+���k��o2`��0pX'#{dm�lT����`в�H��|�`S���V<� xM�LI�G���L���!x��Gy�1������b㾌�J@@:�k�r����8F�A\�������� ���K��BO�C�ժq0a�؛�n@8L��� �J���96m�de����E�Tr�s�(�M��S��8�|F�Q?���Gi��57���\ .
�U��$[Hml�.��Z���cl�>U�)���(�_�.F^�^ҒP�^'>��oʍm��SG���Go:��;}�(��1iX9��_�~Z*]�����,%�}�w�����0�R'<���fP�DC��2�Ԍw��W�3ݸ�=�o��B����\3����zut�Mҍ���㯣y <!�d����xu��`���Ħ�Cfć���f0�X�3���3k�I�r��ex�{6�9��8�Q��Bg�)3�G�[GM��K��j�lR�Jf,�KܴM!;2ÁaӼX`��!��o�	�@7vg���筪�*},1�s&�U��ݻ�a���~@*�ސ�8�+�A�<\�%먔򨤾�,���:Ȳ���FL��%��}���:���sS��7�^|�5�����&�C�ȫ���țd�2�{���Źy'ؕ�jWQ��c�)�5��!>/�1:�z�����A�!��7��v��_"�b�&���%u{zM�a5�6�Ff�>x=V��B�y�.l�'U�jx.�t-JH�=$9!*M�����S��sO��� Bhx��:#mI�C��^{��X�	7�����y�h �l��"��&��8����
#
���{m<�����l#�s�k�V��s�5���nY�Iy9�L���z�~8ۇ{����4��ԣG�.�C�`�#��U?o�-#'O1T�`��Mk�����we�<DT��b��1|Fd��*)<O&�<$gAȋ�$�kF/U^qc6=�GaC�;�����]D#�K�]��Lt�U'#����ykj�Rx|���b=��r��Xl@yr�T�Ul:� �xhc�G(I�fi����q ����q�d��A��y�0 �,N-|�y�^�.΋2�jTO/N�㶽���e�U���(�0A�+��*����J��O!t���}�p@�v��b���q�_1� �r��".4�����l���ɱ`,�k�;�J�cu/��τ�ޅD���ܠ5�3~�)3�N���*���W݂1��u5�D���	O6��6Zh@��]H�̱�#U�-�S`{^�̏������K�E_Z6;k��������++����Ɣ���V��񑉱�|�6��}"!Ai��2e��Fc��®���{E/�(����2���m�̴T��� �}�^�*?�Wɡ��
�^LcL�H;���� �r��U^m���(�@�`9^Q�z4��DT��L���A�I>�0ٔ���)<��u��/�e*��CB"�N�X��N��S��[MY�<A��F�����x�z��y(���IJQC}�-��O�~�K
ϋʙ��DL�_�/KI6L��c��fU�0f�l!����-�xΓ���"|��q�N�0��������z�=�FFD'���w�~=_z����\�[IO^bp�J���+���^�we?��ǒ{��>����).�\ޮp�P��X�)ެq�Cv�:\Su�=���x������w2¾���K��νX���|��"�禓�J�B�{�^�'����$$����.�ub���S�
=У������svͰۍb��n\�چ��j~Ҥ�֞�� �l�/�5���M��F�ע`�����4�e`?��0���k���9�Q[�Z�j��mt\�j��H¡^=+��`ܻ��o��J׾��]�iZ��<;�r���IZ�F%��`�G �!�U�}��}�͔/8�f'X���3Hz�\[����	����902Q��F}�����ƪ$v7YR��5	�a���6�{��?>�h�}��G�C�E��8�9��ql����ϝgS骃ɠ��re�6c���<Ӣ�sN��t���������v*x �2�l��Q��Ǽݰ��[2�*���[]�B?Bj\K�<N�����U��8�9�`<���~�š�ϢoOz�`n�]�#������s����l���!&R�� Pay`�*�EF�Ԫ%|��D$��sE��;/6ەws`����ӂ�C4w�~��'aPq(䋐Pi|-��@�g"�<5"�{������Z?��0�TD�]Kq�IS{�]�O����[���p�6T������ ����I��5�n������#�}�a	6�l�j���l��v��U4_������C"��.�kx�p�{���d�����Ttk�S������1�y4aDs7�%�t`$�p��l�;Mͅ��$�=Q��Y�<iP�u�m���g�Z%O����i|D��<k���GB6�NK��&��>~yl�=5y��D���(E��a�սO��к�bs]�ˢ��e˓k/��|�#!|�kcfI&���Z�x���6�Q�H�m9��7f�� ���M�����e��>|Տκ~2����L�})p�¹R��Y��r���ν&9��%v��(�&�s`�l�|�5�G��?��e=��62��Վ��K+Jǁ���θ��'���QCS�WKe�X�����-k��Bf����EDE*���ʓ'�1�x>a$=���t���j�B{�LJFD�C筈#�d\[	��wY�ҩҭ���QnbC��D_�'��-��ʆs��sV�g��s�;t.+�@�
?Gy�����;��l��u��GP����̔܊��j���T:�������߃A݅.���~g��4�{���{�I8086d|�w�hn�;'
Ĭ���ڄ�����#���;�#'�V��G}��C^l���5}�nj�#9>-�څ#]T�|�qݤ�D�Z'�~�oe�|��S�Z��%�Gi�rg��5����8��j*�ٽUw\yr4��l�.�0���zx�!5u���UՉ��/�G��C��p㸁�#�%*�
��Ӳ^#k�q�
�By���R�5��ıɃ�nH#�`x�B�l7��Gح��e'Y�ep~�X����V:��TAR�˞O�l$��O��}�ز�~.�AF)`zԍ��7�����6A�QT4O�'���=r�,�@ˉ%x�eA�|j����]�G�(��/�md<9�ʅSt�A��ì��R�Mt�i.qpE�/��t�Ԋ26\6_�	��p!��̍$¾�c�h�}%@D�Gj�K�܈.M@�}l�iJ�����;��	t5U�w�>�l�w���%��2���Ȓg!	���&x�&D�)4L��@��1���4f�ܚ�U��Ty�p�h1T��ٻ|Nֻ����w��hdj�,�T�:X.��á��6`���$šl6Z@�oI������/5Y6��K���K�}����Q���H*Kc�����G�N�6��rj�hc�����<<_ն��)��\��D^�B9��lz��5Γ��lFr�����MyW��\F��"���"����l��ޙ�cG{��rS���>P;�
��^� �D��
��׬m�ױ�F�B)��g�+ˣK��a�ᴷ��Ey�����0���ʟ�|my�ؚwjJT4���V�?4'�ϋܺ����OƠ.��rn��v�a��[���	2+�Q�H$)�w���IT�=�4E����
�j
G�kGAv� ������@�+#������%��H�P΍��!L��:u�<��tE�W�I�HpqH��=�g�~�2�6��y� �T�Q�N�xe{m,��=������駲X?}8�~L�"4��}�!���6!n5�Ҁ����Af����"�<� ��x��a�ƩnN`U��4qC/�Lb	8]M�=�s�1>�@o)�g�z��#&q�+/ع�8����� ��zU�~��}�.��ՐD�"�PLMl�mɩ%�J@5���9i>��EMs�K�U��Y�X����E��[���Z�0=�����k�jP������B
}������I��xo��`���m�=,��2�O(;�wQ��,��I���הI�� a_���{7y7H&�'|��Ԡ���SRK�������S��<<W��8s��B�٩\�<'*�Sk��Α���z��2�c�f/%�n){����6�ka��Qac��ƚ�U�dS��ug3��5!t��5{ge�,�{�~i 5�G�K�`�-�g����q���!6�w��;�4]�mn�P����y}i�
J"RHĄB8ր���݈ԥ٠��P�0���-d�M��R��F[n
�A���^���%�K�Y`�Yy��!b��W�]�&75�F���z�V��
(
�9�0xuĒb⬃m�6��[e?j1'%���U����"�0vo�8��F��G5%_8�j�d��DZŝ��Δ�[�Aj���7׿4�S���t8��Fև�Ss<����-1���KÉ]u7р�85x�G�|���j�cKT��Z�!�������4l�2QS5��I�R��

�d.�����ў�R�l)��񺐜��Ǝw�}rу�Ҧ%�ӖL�O�XD�\'�tou��W�bE}ކƖm�W��
�pEo�Ǎ�;Xe7�u4kk�\ťڼ�ja��M��Q��Ҧ��+�&ו�̠���3�������(È���1��o~��*�6G���Ş����m�[��y,A�v�{f�ٙ���og���׸ �d�NǱ�*�N%�u�x9<���\?<8H5����#u'����|M[����l5�����\��M���_���f��iΰ[��K%�*�����$����-Vh�R�[d5��b1>�E[D}���t�j `lQ��U��ށ�KNX����S�7A��$����	:nt�--2�ޫ<����!%0�O��s�ͺ����vj�=Y���m�"�KE�D�*�P�t��L����"�O�JO;l:�^�x�3���2Y���S�e�=��̰���3C�l5� �d������^�1O����04�8ozB�����_�	���4�
�	�)S��^�X�g��"��r	���.�������8��L�(E��&	��~���k�.� �t��i�i�#����Q��I�#��M_-�O���b�$�x���r��;����
��͐Fl3�1C�VL<�.��G��{�Su�u�^"�䟶ۉK��d.S�틿4�<m���[�a��c&��t>@���x� ��	7�*���}%��>�L������w���T$WPqmJ����A��N4q�W��B0��VkQ�s(���&4��uGl���zx��Y|�2�#<O�l� d�#�BgK,&�;�w���_�C,��q��'��$��5��Z�w�I��6$�z0�iF-8Z�:u�V�v����R�*�<�&��)$�W-�⢴����⟡/����6ʋ��wyW�f�Tc�b Ǜ3vU�hnn��1E\�,�	���60����Y���cf�`w�xpB�@���g@�,0����6���B�i$�9�9�F�X�����U��ŀX����0:ɯ%*�?�E�ڸ��Q�Vd���ǈǛ-)� '�'ASv{�`ߐ$a<6��RL���$V�$�?\~�� �n�0T����}��B_;$yB�f�2%����s�����G����Z���S�j�8P4Ip^f�si��E�Kq��PƩ	�d��I�tB�kA���uŲ4öՕ��^�+�.�lau��Z�WT�u?�b�e��4Y&e՘p��~�ѧ��dV
�Z)��f�_�06���\价(a�ű��(/ �w��w�|j�f$�ۙ�z>���O�`wz�m��{p�!�'��؟������ח��r꫐�4��5EU���($�N�m�ئ����xN�ĪVg�t��_�f�z�sp�j-v�M�4��m"*�9�'���*��D��I&�Qo����aoyd},�^�$�	�u��U(�[��ȁ^V���,r>17l'�탅<�)���dWg���!�lHWX��" ����z���+홹pNw�i�&� .k��.�Ƀ�D�710hX>�f��,�bA?]�lS ˏmS-&��r�,5Nx	Ls���X��E8��)�g�4mgLJ�eV^h5{��.0��>:$LU����Pw�1�����g��m����-v�HhF��f�O��ʂ�p[.g���qr��U_I����w����ձX� �(7�:���+��鴖-üh4b�,���(�^����V3J��dŗk��&b��!��kFYiuw:/���!�狏�k0H�ML�<(���<N�J�A}�����!.c�4��Q������Y�̖_q9*>�ePUr�f�A*����[x�x���G:�/����4`��<�%6��[�+�j�_�9��ߏ-���_��	 �-����~
0C�A���f�A�d���WSrϛ�K+���T1����)�H�{`�m�qCvn\��Vo�yŞp�D��y��b���I�=� � Y��]l��{a=�HH$���S�1��b k���mk)X9��E=���e�l�t�2���H��Tӿ2C��R�䯲 &bd�v�ߜ�U���`��dÃ�}#�;�*���2�������T͢�P�ֹ.ѕLx�Jn�|f���3C��j����P:��M֬�l�j%�ݎmEe��ƕKٷ=�ῩF�Ӽ�dos�[8����])�v;�����
������d���aAd��R�x���j�?Ҟc_����v�S��k�ò����Q�7�Ef��4|;�0��n{sW��_""��@L�ӛ����tp��f���n����B?\��k�.,�Am5�`!Z�h7�N� �M�cv�Ϝ�_N߳7\�t3Gxopq�j"���?���|J 
�9�da>1�݂�L����I�+�(�������e!�ǌu�u����},�N<A^44c+цYO���̓�wF�ب·�TG�o�����]SI=�uⓖ�2T�7�ek	r�i!O_hb>�� �N3P�}�O�V�ک��^���֎+� z��;X+��XgƁ�g��ǝ��2Ў{�f�zZ������bQWs}���<������<�����]ξm�ǘ"jLV���#Dz�F����#��:Yw�+�J�3�(��{
0�M�wh���[Ш��K%�)�FM���x`��	�k�d���|��1ѳ�f�yuc'/*��斂Q��ٓ� �*�Θ�ϛ:T"9zg�LB0'�c�`=�
0U/��X��S u�q�Ԩz0c������LY�T�~ɥ-梧��)���B�u1$K9������Yvp����c%�p���?k�\�@�^�=W0�4�a�uߛN;���q�F���*��` ���A���� � �b��P5`:��� u�8�<^�Ytu�wd��"�ۻ'6��[SQ`{�$m2�N������?����H�uc����3��Z�8?�^U��ș��Cz1��J�9Rq�Z��@�KE���OF���X�m&���F��&$�O�Ќ���I)��q��Y!#�4����?������Xʿ�X=F�e�ǰY�_/َ�7V�"�[��Tc��j��B��/O/� `˔\�N��'@��\�ĝ,,&Yp;����� �ܗ�!�dĢ:Sݧo�{M�.�%�Cd0��+�-���z�<f�>���s[�!��������v�E)��\�
d^��MR�2?v[$ql��9��-�U G>'Յ��8�H� ,�;�+�۽��ǀ��X`ޝ�4R]��Ì���Wb�U�W��ˍ�{D%�]�ٮ�^U�̀}#ޡ)	.d{3�E��ߕD\}��ʰ���XT��CC�� ��6$L>^Lwf'B�j;�f	/��Sr+�􀾡d�5�Y�}��o/ [r���b �Ҧ���٬��n�NY����� m��r���O���NxY>Gb1$�!&���֗:�l��>�YƇ�j'ڛx/?�d���Jemx� J��jL�8�U���SjRzU���qvk�` �'���\�)j0���}ɍ-�Gs&�C7Y�;�Q�jD��&3�pY�Z̚����z�Rk�};CĤAO̐7�@����\f�}y�]2/�1 ;dД���;E�*��!�o6�w^����[��ۙJ 9j0�Ơv0��U�AU�"3�y ؘAI����OLNҒ����r�� ��U6km�j#�d�8�p� n�д��gQ�GT��;��x�Ru	0�9��{���ns�]��[�� \5c��߹�~�O�((b�`�������[�f�m�yF��l���q��&Te 0�Pe���:�ج�{�7� �+�E�Ɖ�$�E�3>��O��-����E�2������W#�S���Źjz�7�$�A�<yP
�c���G�L�*M՚�f�����(��l��{G�"F4g�co���{���@դ�.��Yx��G��!�#".�ȑ�ESj!�U�5�9�-��{g��nj��`�$��?��z�0܏��֊�W**sb��|���at9X��(� ��4||1���'GE_�&��o�}�x
 |�����v�c/����]݉Z��n3V�0�	Y/
0�l\9�b�˗3O"���Y�������,��1���A�j����;��۱�\tʗK�LX
q�nfl,�Rku�kf���!�����,b��H�4E�K�Np�E6@���kr\��4.�՘�.ތE��"n5�����Q�P�JͣI�^X벘���b�u�`�����dg9�_^^�\�9��lC%O���A����r��l���� �(޶��$�C�Ӎ�a�>rY�o��n��b�������G���_�A����Y��,��6�������<}�I���/s���uz�W�[�C{�6G�u�(�ኄ�} u����}��X\�b۞�o��>�/�Z޻�U���!����֣�>3S�/H
��d��!UY�T��0 <e���\U1Jw:�b������1TŻ� ��F�s�U.n�!?U�d�)k�P@UPL��|{��n*��\%p�2�_� "�.rA����{����y���xX��E�X�-Vhe�oY'��� e����5?�!�������K��YE6kwnD�½�Ō����n9u�ɡm�30��0;��ڒA/����޴�8�G�-dU�]�|o&~.P�^H��96K� �c� �X\c�z���v	��׿|+��#�+2Q��D�W�Оm��m�����%��Aj��ҕKikqN�[\�]�P�خm`����Ь�{��%[������s��\$���"6��:!|��:��Ӏ�1u��S��-��S�D��~��T�ln1�?�͍ ��X��z�zU!�=�?�Y+�L�8�t��ۊ̮RpO��A�M��~�a@w��e��l��T�)�E����L�mh�W"�����E�c�ڤX;���,�����=�=
��L˶[Rk��G�j�A@`	�<�np@�d;Ih]���Z�%nnֱZꔬ_Ƴ��.b�]"rT#�oF�2~� �h9�+��{�?�3�ܠ��x�Hc�FB�ga����O�c����P-5��;�Fױ�������+����|eU�X�vB���uj)�E�r,f��I�8�\$LB�\�<�A�M19�Ų��)��O0L�HE�7�K�����%����p��dx������,��"�[n
�=X5Z���S����08�0��ѩ��y;z?��ҚwFk��Z�=L�]$�+cq����V�2��Mnu�ķT�=E�W�q�l���	����,d�ns�B:���,/�b�7K}x{q���&˶ ��ٸ�{t.YLw�ܰ��VS~����Le�����4�q)���c��j��'t�#�/�\�X��"��5D��WT|:a�$ˆI��,��M����H��u��xb1��*��ѦΡ�k��!�*���~���(�Z��s��RLu�wBJ	�1]��bC���ښ�0���������Y�;Á՚��iP�|���z�$m�c�{>R'��!��<{;��8]T�+������9�����{>�fXDE����u6�'��kI-���0(��i�S	�㩽�U}� �"\�bA_#��T%D����l�n6��  5�Ֆ\�?g)}X�u�Cm%D2���?�9"-5�=����
�����~���:Se� �)ta��x �gS���u�\�XFVæ���B<���{ ʒo4F�l���}D[��9����4�Ё�:�>`(:=jjk5�7E~>��a��^w?��n��Ȇ7��G�E��'�KIQ���b2�B��K���j��������E-�UE͂�(k5���	S���,�|C#���k�[y�(�i�L��]�$'������ܠ�~�$�������L����J��FU����Ã������5U��E,C>"u�i�%�SҠYJ�*0 S�u'2�֖N�Vl���(L4��Fjb�<N���Μ޹�}%r���Z���
FԠ]�1ս�0��,L�J⃤�������Y�>�n|H���U4����QWx��D��0P�� 2��?_�S���dY�K�%�g��-ʐ�MV�����5��`6� �s_���>@97 �~�h`�D���F���|*��]��' bZ�k�\�UR�o�����T�!:�y�6�AaclQ0�{O�oY��k6q�uFi��l��҉f���f��}�d�P[X��.X�eҁݒ���sd���х�K"Y0Q�g�]R�o�>m'���9ϓ3�QW�~�{ �s����Ѭ= �8��� �v|��%�1�<��aq�p����7�L�t�19��ۛ.��[���^;���h{��'l�Hf�Ѝ��:oU+G<ߒ���[���iM"�Xͬ�Z`�
i->bh���s����Jk u��nY�O�~1&I��K�@ߝkϷ)�_$�$t?%��'U�X��7�hFGܓ8�WK�+���j�"I������ox��v�z/-�d�V��H�̥~v�p[��+��,3�	:�������*��n��Mk	R�����O+���*K��F������A�Eފ�!h��'�T�ݴ�JL��.?�H��}T[�mR��OX��O�h ?�k��6
���H"g3v9�zZ�ɷ� � ��H�m�O0b׹NC�F���G:ïQ~m@-ɲ�_�{J1�Q���E�K��)Y(=���	T�[��DΨ�8Y�J�%�ݫ[;]'�wH	�����D��H;w �����jz-(1(X�MyVIe:�	ѩ ����ڔ�۹����X.��M����z<Y*�[�TO�Vr�_�����%��t��7H'�9Ö T����ƣuu�͢��	*��g	� AAn�&�P�v�K��q:��p�d�LAO�C��5?�7�,8|EїJ.�(Ā(]]���jv��v� L��J�n��J6���!�l��r�%��ݕ�H����'>����T�LJ�Cg,v�u�U]�jS].�������Ez臷����r��/*G{���R �!���A~��4NN�0��Jf��u��&��ug=��>u��;�j�=/������x��~T�Z�F��*˞ ˿nȡuQvUM��N� ���E����y]��z�͇g�g��9�Cc_���v��B���9WG�b�u�o���6���V��q�V��̫��3CGF�CG�Dׅɐ@�E#��
����6Ɏ��Mѿ�΂b���"a��D���F���S7z�`��}[<$�Tl�Q��ѿ����db��rdv�M]�{(�T����32#�7)0�$0�,��%��fJ�Ek��U%�N�ۦ�[s2�$!��#�����ܧ|m�V���ΟΏ��-�UUOhc08,�`��X(�C?� Ms�=�/���^��.��p%�	م,�;r��H�@0,��wb��t�C˗1�\e�J7��Y��̙���8x�]�m~Q6�� �ј؊VF'�NW�i��e:�8t�`S� �Ha�K��l���fu�h�'=�#g�(T�z�Ƒ`��Y(	�~,��Z��~\|G�X�l1ӻ����ġPo��s���p1�)��h�]J_�ģ�y[�wO�[�]��~�v���q����4//n�K�,�M��DxE�`�غ>���!	��J�w!ڣ�"������>�ʑ#*Y��S�q��BH�6�;��
0�\m�^�1x� GJ�3��T��;o��=t9���Y��0��~�gK���k��lT��w�铦�������x�Yc�$���sعC�l�z}{����QZ�L�r ���ە��|J������{tK(صAFn��h�'s���I(MVʉ�,��n>�tSn�>E�@ީ��|�q@������l�l����4@�j���*���uꟗc�V3r�͖׷���[�-�H�"��@GNb4�\0X u����nLxPk��ml).�����;�g1�bǔ/�:�d:غ���#�g"�RH��ޮDp��r��^�_�%IcA$J~����3�5��0mgNn�&b"�TF5@V::���Z���k��Klf���܀d" E�d�3ؔ0I�Z�@`wΏ�����,�� �(1��!���F�spI�:!J���<y�XOA�D��^��ܗ�oW\2�������_:���3�,�5����:T�'<�l�!@�h����DrV�D�?c��o��ژiX��u�b�����J���/���ڴ�#qp��K>to`q�y,z��ګ�J�F�T�
߁)��By��/.��)�`����Z��Y��E���F� )��[��|�&;3M�&��� 0�\��Vb���ٳ8-�gjq ]lv�>�,i f�@i�A��"��a?�`�8���Q-�vbsVzt �[�"b=yY-������2� ��1K�\��s��fR�&�[d���ϮtOxH���V����ڻ�X�~w�Q��Tk<Ìk�ހ��}k��x��
ʞ	�Tn�o���z�ӁiX�F+7��'���g��G]��d��Kr�
�h���6�eB@������( ��ʾ���In�;�j��,2[&�Llt\�T�2 I�b���τ������U���q]���q�$�T)�⦩~��ӶqS/�t����N-���.Õm=�&���c�J츗�Zԫk�[�=��U�U�J��L��P# \���v��w<6���wS��<Z�[���㯶ɯ���2��.x�y辫��0��&��`*]4���ZF�3��'w��X�ͥ�ں?Eq�?HE75X;Ia��r�]��RR��T��5?1I�fzp�S��?2ԩs֏@�.m���Ń���;��֝����7����K�2�p� .
tD���>�01�Z&��+a������y�,�ӧT�9M�l�ce��uP�C�:�1�-�M���x��C�O#�z���O/�/�X�'���
OR��!�{�n��dC������>�����͸7�e��D��^�t�c�D@�^X�C7�b���-��3t�C6�Mf�#�c 5�-���'�n��ɐl��v�*����; � ���!k`���?���*X��N���d@�	�@ߏC���').g�0�.��H�wU��W�m��i��0V�l��[p-[WF��z�G��;��'=h�������:�r_�2�/F?��z`��⭬��*>����6��^ :�� *V� �m��?���{��� ��~�V���r �N������f�j��֯�����T	Sq��i��ǧ�fF�Ty`h�;`�H�|'���=��l�f�+�$��I�ߚ�?�^*�`�@7����2<If����+k`���p/�,�ۼJ,m����,��B2$��0\������߸�>1��ET��x���u�Ym����>���||�~:Q`��SJ��:��*�f��8�Б�|7z8RH�S{&l`����ը��JA>-ub[��4�#�R����6W����e/�hX�F�3�ݱ�}�@3	4��ڦ����E�+�D!��IC���Ӝ-�Y�g(�+t���a(�n䆺3��y�I��n局�(�=mМ���Y��I`R2:2��qHqqn�t��p�U�^�k5_�Swi���8�����םc�c� ��B�p0�s���l�����������P&��`������}�ܪ���-@2�+KiQsv���}���"����liy�6��Ę�>.��~��<u��5s��T��*yE��н�������s<����(����>���Z�A*��`9u���LQ�wX8� ����8ܻ���6�su�χ�C;�/�y?���i���T7D��!���gl� �\/� ��%���'���ž�e���w
6Pm]}\�����R�P�V��ޙ���f�����big 57 V�j�w�W*��v\fVşG#q׭n�I,�`k��]���w��������>�n���K���OP���,�r,�w���$��:�)�'|Q}�6��kcx4(F%l�v���<&ƭ�x��E<�`ց�9P��t�o��,�1���5�؂�⧎]*�`q��45Dr�o)j�|�HO��±=��Ż�۬U�������/������� ���&Ȳ�@̆��$��^�dS�a������1�M��F���&���Ѓ�%�g����g��_�a$i�Yy[�Yw�����kiz��J��/��/����!�h[���P�~�n�4�ca]=���kT,��A����S�JS=i��^����a�6���y1<P��գk6�=�n嘾�O�c��Y��1mz*|vy��X�����S��w��q��s��hWg��}�&�N��I�l�b�,�m�`ѭ� ���kL�8�B�E5�83u@-q��R;�CWJj;`�Fl���F�e4ZI[�m�6|Q7�d�wݖ�+`e�l W�Z.1*cy`d~��35<�\]Xa�����t�t�W>*�H�W���
� ��嶌J�����S�<Գ���h�WH��Y}�yR��w��.(X?߻<����� b�Ev]R|<1�y6�TUI�W������:M#^-�GH������ٽ3�1��n��.���h��,�2����;�uɥl����R�>��v����X��+����ccP��eZc��F�����$3Fy���S�~���^�i ��A%N�Yi�lX�����/�J��LR�AI
��S�-�Q����y~ j�bBtr{G����f_)�����w'S>ֱL�����2�g��=6(�Y��t�+��E�Ygq[=�69�� ���<��Μ�=���q�r���xPտ�y��@�C����ѦVx�!�}��eKi��(A ���A�bT�4�q�U1��d�r���-�K����}d�\fz=�'�K��`F\"Q��Y�{��i<F�S���`0�x�� �V��\��	3�8�����G�_L�og��R�A��fU��/:��|C�X��;����+��g�|~����|D���ҩ���>�<�(uv� S\9p��Z��T�[q�Vx럄M[�m�� }�_���q�.e�䄣7�"��擘�:4cʬ�Ⱦ�=[M*��	��\��� <�[�8�d�+����yh��F�d�PԘv�=��]s~��@?�߹ �5�%z����ùd	 �믕�p������:�]l�.R�p}�(
�j��.Զ��W��鬻��K���j�0�8�eY<�3�!>�ﲲ�b�i��7 ��F�\;�/28�}�ى.�}8&�m8��C�����'V�]ǆ� ��[�+�����{܆���y������5 ���ݝ��z�.��w��R[�!�r�otc����p���@��:���J���S�_g�L@���=�?�/O��p0�e�"9r��Ψ�/�>B��8�%i��/_�@�ئ�Lq�Zҽ	��,�Jr�zO�� ��F�<�{��Lee��ރ�k�tӱ���O��>+�ɒP���6t�m�^6?�����A��ꁁ�����]rS�,7����$�,aD~�;�΃�M�Ck��Ű��k� ՘�h.'����VM�ʠ�zN	�V ��c(�QI�dK���I -Ѳ�� �ky���Do���^֟慨��v�&h~�yn|��� E�J�[z=h.k_��"?�c��kz�´�}M'W )�ں��U �����q��� cSto�_�]��� )������6����a2�(�{�\CF�e�Ӽ���GI��T��<Qf��[� �@e���G�D��o])�e�N�� &��8'7��[�3ܣ��Q��1�E'���n��&ؖ���o���ư��#���Р���6������8��n}����{���x&������V�W��P�������5�>=	ew%��9 3�9�X�O�8�-8p�(�T~3�	Z�v��wI�L� ���Ћz��=}�s�����休�n]��\c����]������Dt.*���(��yq?T_X�l�o���X{���	�s�P��ڒ���XVX�����;��r+��S�
�-��?�u���*�0n�qӎ�6�8���h͒7��`���W�6�}��X��N�6q�w�W��x~��իǎĤ��ş�Y'�@Po$�Tn�hT�\��e9�ֿ��Z9������W�=�T �ʺ`�7c��gV�:��ZW@q>����ά��ߙi�e���T��~�[%�m`|W+l�%��h�=o�t?��7 ��2��_���݁>�T�p7Β2�R�!^{�ۨ����^x �.��蛼Q��cq�����׃�{g�܍W=,��4d�����>�㻡_�����cp�yky��b�#N#
�nj:h4�3����"�ͬ�d���)}p1Z��?��4�����t���#D-߭E؄��1�Y'k��9�z��ze�x���Mn�w���΁�c`>c��e�,�˘�4�ߑ��2
�������n�\�%fhC�o\LK��96n��X��ne/\�YKW^��S�(�y���o����kW�I:6n���ȼ�4Ie�"B�i��o�ݯ�$[Pǘǣ���ÌR�)��Z�'����,±�[m�}�������Io��ߥ� ��*{���a ��Sߡ�[%�r�[�4(�5_;p�c�禜�G'6��K�Fπ�6���=r8@�3����z�ܧ������R(�p��o]o-YgO�d֧\�}��^�)v���X����2���Ѧ(�&��8Q������ƂC����~�d'���)��B_���Ѻ=�%T�J��;��]��_K_=�4З��Q��g�=�����e�!U]8w����.:$�1j�L5�#��ιN�V}g�`T� 5��`T���o�*ق�Z8?��2E�W�VcM6��PM<֋��i	l y�P�[�
�wN)�!�C�����|~q#!����!S��|��n��ǡ�����[��R�D�N'A�-�K�Y��t��M��%`-�ɟW�r�����'����j2�V����ʦ[~���rI\�����6��W���}p�2��}��/*6wZ�����%[�o��nZ\H���"���R��m*�p�l��ˍ�޺����,9��'�R�Dr�԰�g]�F����؁��5Fq�!i6���i`}�t,�z��ì�m��\�%��jL(��1�:�cI���z@}V]8�3L���#���هzܨ����
x,�B	����Qs�-,+���`e{�鿩K�%��[Oe>�$+�{���Jᜡ�Y�]G\����׈fƆ��- �u�lQJ�w�`*�.w(��r���n���D���l�����j8�'g�΂���v�*�2��~7r`d7&������h�o7��V�m���@'��X,���Z��mj[�k J%�9	X��D
w����ʕW&�y���o�";�gÚ����w��X/&�߻�
��º�@u��8-���ه�����p9�]n����	�vŷ�7z��Jo�7��a�(P$�RV�6~�}}�oIE0ia��Vb�������v9������c�ނ��(�̠�ߢhq�e�z��o��ZaL��o��9����<h��*0�r	��p?췣6�>_��T��|N��Ƨ�*�ߠ<,�~w�H(�t��Y]��
�ӿ���~���^�^U����,�3[�E��A�$�/' �x�o��(�����\�PS$O��@���鋅���^����^�<3�:�k�(B�ڱ�!
���������Q4�RZ3��������o��v�Ks�NZ%pB����z������7����@�9�+T��6/y3Z�Ae� UϺ8x��p�r?T ��{m�
@�
��=�Et%�%��u�s4�i�D��k��	dw������w[�ÿ�Fy�c�pG~#���H�^�A ���u��R�dw���m�DV��Ce�|}�!�ѩ�S�fP%	Cݑ7������F��̡�xf�6�3�R,�q��d��K�'����D�wQ�Bs��`����N~g��\����.F���~��f4dA��{f����d��b�U��8�����E�(
Ĝ����{��L���	�q}b�8�g� *�'fKS7@9d�g_����>�6'� xw����o��@�I0lX�-�'��=o���쩌g\8�%/�ݱK��k��:/�/u������s�7�,�v���1�_�"��z��#"{����M��t���H毚3�-�������)�D�<-}בE�Z�T�F@��<#�L>e��N��b>_Æ*>���rt�b ��P���jTc��վ%���: i�
�	���V���}�Oe`W�5�V���ڏl�:;�[���p�\�c�I��8�s��ˁ�ߨ�5�M/\h�O,�r��9���7�WY	>[��?�}o3���4�jn�t�;�)'DnQW���Q�s�5a�CF`|�z�$�"��~�z~&mS������c��������^@�J��΂j�|MxZb ,�&�oGө5^꬀�r<��~.�ӳ��z,-�M
o���6���>P�Ľ��D�^)4��{��X�Xg���c���{�N �m@(��b����/�ז� Բ���n
0�[sh\^I�'@=A���b�N!�$�����?55\1{=�O z��%��e�)��f�*"1����z���G�~�Y~LZ�<�ew�e���߬t	&I�:�=k+��h�����=WF�)�Qe��t��O/��so"p��j��6�L"�yw+�8Hh��߯pJݟX$��j���f	,~Ǆ���ܨ���Зφ���[%��14ꪁ�fe�ʀ�l�ŎMS�s�@5��F*)R�;:��I�l���j�U����l���ն�<Ի�Ȣ)V���-ِ�4�u�P�O)��tK��n�!m�S	*v�3����3���y���GJ)׿G-���2����P#ɇ��*�nN�آL	7,��R����Z'�ָ^=�Bqխ1 ��ԇj�SZ�?Y�16�IBL�@�&���lTU|ہ��N��CvR1��Ӈ�,z�{3������a/u�Ջy#��Ξ�L����{�
��ܕΩ��)اӵ�3uF�.���2�v�����������`*��ߨ�u��l��-��l �`;��o�l�绥���T��{��f�ԙ�BM4I��2��b��%66�����%Q�
Ñ+܋��׽�b@�/�lUe�G���{ey��^�C�A�/��yت���]_�x�+�[>�_�F���xf2�ϴ#�1�]�5eE��d�RJ�5�P��o�q�N}�	pW�$�B����L7���c�'��-�>�r��>�<��_�q����\!������t�ب�),�Gjn��tG[�5Q_q�*��F�~Q~^O��u< �+��֊����O�n���jj��U C�Ѐ�n8�-��Fq|@T�':F�������Qt��K��f��>7���%A`�n�=��<���:��x�Zj�����d	���{��˰�j]�<�R���<P��	F��}.ZW��Юu]01�eJt~�aճ]���Wv(�p.� TI}M�^/
p/�~���v�A���5�Y�u�W���u�)@9�Up��>d0e�U���X���/sC}��P��<���WZ5K^��s7�0O�r�XLL��x��Ub|^�+�?�����\u
&1��w�_%ӊ�//a�wW[�kUO�סH�����F�1a`����|�X4�=iAO�^�Q����Yr-�|Ր�fN��3בv`3�`�`}&�1��r<�9 ��P��[��m��g?�p|Б#J�|�:���N�Ux{Q(�(��u��u�ۋ�~͝Љ��=�&e�#�#��{PM�V�	�8�7��HTd`�4���sp�
�nl[��`������2t3;͏��:����8)�)Y7�Z��O��t��w���B}Dh�ߑ��u��ӕ��'/2��6��`��1��w���fO��;���������������L��:�ћ��V�5�ۃ����:t��$��(���H�Z���F����UEP"¿�j�m[�-�pϲM��X��X%�4hh�����v8��{pT�GO��\�`67����z��y�u7��C�̰�ϫ����9����ifxd�@~�?��G������g��h�s;�bn���W��	�`�<��9�z��
��i/�+�Ղ$$�Q'�q��V����
���`5���G��3��@��
^Z�f��b���N1�LS3T	��"J��-J��(�����qzf�7� ��ʹ��?����g��3��j�9٠
�ᚆ�/���U�X;aU�3��b��ts�|��g�>������V�%����ӂ�#��^ۭeu�y���j�qq*1���祡�.�N��W�b����v{fKs����z��P���o�>��|����"���s��~�Q�����h�f"ӱrǏ&�5"B�������ig��N��[���'џw���i�T쒢z�"��dw֣߳<c�t)E;����U, 5Kr��`�-^�[��?��i�
��_Ӥ��D�+[]��Ka6�i�=�wc���7�n�9���]%���=L{ ����Ҫ.�o���}q����
i@�e&��Fã��}��D�S��o����"����Ӣ�e<b�J�L=�����~~���r�N�16R���XT�Gb?�H����zx��m�났o%�;ϭ�*<���Y���c�S��3vц�A���n�� u����Yw�N"Z�sa{����P� �8�� ���6HKl��,��3�Q$����y�)������I� �MS �n�d��w[���*��Սt��u�0l����s�>���WL?�`Դ�ft9�|2�Z]d�d�ͻ��`�h��oZ�!h�JoÑ�]!JK�=�F�:��ꟾ�7��o3�
M��-å��{��2�4:�S��Uۋ|��@{x�]bI^/�W-KZp�@�؅��P�;��� m��|�-��#s@JF���L�dAW��w[����1ԁ_wl5��udB�K��B��C�v3٨��O��%L�(!��T�����m'���$+�B.��-�u*~]]��C�D�Xd˾� y=�F-�?����tC3*;��&Mx�dfg� ��pʳ��M�� v� �%��*�Jk]��u �f`ZOma���ӫ�K��ľ��kd��u��ޡ���0�u�.~ﮯ�z+�	�s�¤k�����3L��i��7�ˠ��&x/���q��l]���Ii���v��Kg���P{�=��!�]-���r�tC��h�5'j�j���7����K7Dd%&Ͷ���y��ƚ<����f/e�ǧ��<0����Id(���������t����Y�<j���_ ��<�PwU���n
U�U^Uז G�[�BΉ}1"t[�������QҔK���μY������ ���?Ix�x�=?��v�>���~m�_Q��*����Mn���%V��o��A���Od0����;���%ݥG�UkV;g3fD�ڡN�7�xZ��q�p,�)�����$)�s������J.3,O�1�څ��i�����o�\B��$��u��$ak�<��J��j'�`��� ���ȸ3"y��+��02��B��T׉�W�J�	L�!܎�2�@e�Y�ud��%=�I=Q[��75�Y�&؎�ǲ� ���K��2�b�� t�p��ʒ��j-� Ҥ�����^π�����|�+���*3{�1���m36��q�����P��������xX�~���*����gHo�z�m��B��	��G���D��6���C�������%�.۵��������x_�5�|���� ���9����*?GN5�vV!����Kj^t�g����D1I�z39<��'��/����v�ݣ������o��E�_L'J�Xl;*��Rf�^��/V��*�)n�c��	$1Q0i�>��'��cM���G�p��2���sh��:���Y�\�GK󎟹Xϝ�
�P;����Mq�� ���Ys\�ȯ#Oʈwsv�t��F&����"=Q�P����6j?QǴ�^ǭ�x��hA%���lil�z*֮��F�m�XZ��3���[��ז�2T��V�9�g�d/iF4�[�Tk[R��Y� 5?"���vA����ύ���Ϙp�� ��:Vt4f%�`Ө�� 6T�`N���.,A�՟3`�OSu0���	|m6� �Q���[\�R�:⃱�J��N,�E<k���j���q��
 ��O�U���`O�PѦl��������u�Y�k`�9b~|�$��G$����=�j�i߹n��^GT;�~,լ���3|�4���:,�Н۽O_�>������^X8���5�0ϱ)ht"УN��$0��<�<L��a�vG�<��i� �<i&��q���3��6�9�R�O.uZD��ϣ�H��]�HE5BKz��0�U���M�5�j@o������ju��^��d�����s�䅀lҵtj�̢7��$*�^k[p�Q�;	@�hZU�3�OF��Xg�O.ԏ��9~u��Sl��>�e�t�V�������.�b�������YP���w�j��� ܮ�m���4�p�
e�+���+[�Û��-���FW�<4k�X5�F���b�Xn)ПV?nج�a��{U��7�AHA����~�n��K_s0C�Dx,>OK:�(��a
J�Y �u�):������:J߲
���欄�y���a;��]��8��NV�U�g�^��bɦA\s"��}�b�Q����,-/C(��y!Ȋ?g��I5 ��O3�OE�n�BWȳ����@;Xb n�#���ق�rYR6�P��X����#;���n�
�p�H�uR_��1�6|�����ڕ�|�bl��K��K�3�>:�MR�v�@��`\ʙ��h�IZ��c~���X��&n�K��g,4���?vbTt�J�˽��3����x����hi�"��1����":�d�&�M
f�M���^q)�-�����^�<��F��:3!}���x=�30�,���B1���5��H����H��������*p ,E#Ȕ�S������(N�[�Θ[	�e>y��:Z�Y}l��S�`q��C�Y[,�k7�h%<���J*CR:;���6 �Jǚ�O�Xs_m�B���}���T[0�0LƝ�3}�E���]r�E�;��,�`�w)�Np���[�f���*f�j�;1���p$^��.�7�ҥ���~F����"�X�ॻYNPC�dlJ�B������-���߻�����]��ի�ATfs��u$����G&0�h�0�	���hI�j�v�������5h+������\���s�ݖP��kP���8��J�
z���T��f�K6\����}�1H8(o�K~�G��0t�����e,s]��w�[�k�̺��a��u���u��?M�]ө%�ȴ8�}���Oq�\���A��2F��1���K���c���>�N�>:�wX*�����_t84������¿D@��F�/N�F�4́���㖺�tQ��<�~7�Ȯ�`�HKJsbz(O]k��Ƅkq�d��J⽶T@����t:�B�5$@)�n5����[�sw�~�VH	�Ԏ{�Z��y¢�"���-�ܿ/0pŽԓC����Y�M|�S�����0i�7�#�}}�9���C�u�=e�bYdG�}��X��c�Z��c�fĚ��ñ�vY���}F�x���^�G��ӵ�9�-[\E-H ���J_�\�g�J,e�<#�;iC�Nfi�:�lR֭^�u��nr� "V/��T|�.�����:��Y��zݥc�W7���(�� �t~g�$,�}��z6Gμ��^i�wLɥ���I-�X�O�=M�=�� ��$Jͳը�nr�eۍ��6'�6���o�&��}�gW[%
V����A�����]~�U%7��q@�5��[��s?����1��u�n��|O��󌠊*�q&��B���==�Q��xoh�����㧗�]ESl��i�����kʕ���/�������R��o�n~� �����J�o�G�k�M���w�3p���U_�6匕BBe`*g��߿ ��g��"������tӧ�����(�"n����ޱ��$����������~����Ӊ|V2�:co��d��%��~��f߹���2TH��~���ݖ׳g�A�g�__�?��V�_��-�ώ���|�$�c�'��R�]'��������+������VuOK'���<��סn��.��޳!�*b�Ź���%�{�GI?�,_2��G��������{�v�^��%�2s�E�au��K/V>��K�񳗒���������xQ�	��O��9�}P{2�B�L{�b�.��><I�U��Sӹ����O\Z�X�|����Uz���| n��}M;���ձ\x����蟗Oԭ5�ry�|ß~��z�K�����Y��(�oy��L�-�w+����R~q+����. ��Ģ��qe?|�Y�������ӷ��|bmw}Ї�㱓��"������B�B��dں�+b���ָS�o����{t�<P�J��WO_�v�~�|���#�Vל�/�ț�+�%�'y�O��ϖ�ǅ�=I����+��}QG����K�'._��lbC��E9s��y�/3��,���~�|Y3}����+��V����?*���廜)�X��O���=߀�]��w�.�T���|���]>�|�w�.��|R����]��w����~�]�#Mi    IEND�B`�PK
     mdZ��S�  S�  /   images/e5551f5a-2fb7-4493-9527-57db21faeaae.png�PNG

   IHDR   d  �   ��'  0�iCCPICC Profile  x��||eE���Vx�*�g\�$�{�R�f�IvC�]�%�lv7��l��U����E�4��)"ME��   �4AiR��=sg��E?����d�y�3��)�s$���_�`Ψj�̝�h�{���{�U�J2:�T�͒/�,\���Ց�'�~��ǒz}���J��~֝1�p I�W,��K���- �~��g?G?K�0��g9z�J�'�7q<�ݭ�S�d`���>Iƭ�?�ha��������sA/=a`ͻ����;c�I�*$�̚�x��ch̹���A��$c�\�?<+I���g�\�FЭ�m�Ϥ�%�����2���L�Ve)cͩlf���:�����y��C�4MR2M��4�1�5�kʴ\����Ӕغxx�ඝ�{Y��"��t%,I��ݒ*��,iƫĿ,1h�HZ�Ix�:��&��;�%�6I�8S�ׄQ�u ���M��{���K�<@u�ǵ�1c�%m[��&���_��^[�/X:<4k��j4m��>o��Dғ�,�6�~{��ǆ/<�����,��qA��m�b��(I�x0I־<�m��d���䶶H<os
?>Y/�*����������\�\�ܖ<�<���|аJ���a׆}�5��pm�C��Z}T6jڨCF]6�ѕ�;���ţ�����1��yb�cg��b�?��qG�{`�F����J��x��V�b���X�UN���ʌU��j�w�ֲ�-��կZc�5�Zs�5���'k��k/[g�:����7�׽�+����p�m�y�6Zg��7�k�1�\���6���͏��~1��m��~�u�J~��[l��V�m}�6�}y�/���EM��w��W{�+I�ͮc����r��[O7]v�v]_����w�񀝎���-�M����I��y��[���>���w���η�n�պ���K{��6a��ݯ�c�^S�q�7���侳�~c��N���L6����۸�����l��O����[,9���.?x�e�|w�CN>l��O=r���>z�1W�k�=z�~'�;�SZO}��#N��ߞ5����\r^������{~��ŏ_z��G^���Z��p�'�=u�/n��/�~�˭�ܾ�����;���{ο��yp���,�����ɦ�����y~ʋ�_������ޘ��No�w�����?���-�D�X���3�0
�]�ɇ�׍�`�a��='���W�4n�q7���Ru��W��r�*Ǯz�j��~��׼`��׾}����z����kn��F;l��&�7=u��o~����K_�дE˖Ӷ����m����^�ts�ǿ�B�f�o+�5�zzc��m�n�f�o���;v����>���']�v�ΏM~i�w�>v�M:d�nS�N=������~�w�i[M�e��{�����7��+�Zѷ��[�o�ϔ��s�<`�wf3��}/���9��}h޳��\���*7^Դx�%��ׁCK�t��g,��;7}��C�=���W9�z�8j���8z�1��=��?8�ǟw��?���kO���מrթ�/������'��s�g�z�~t��G�sȹ�w�����'����-��܋g^���/���h��+߿꣟���r�:�nv�6��׷��q��7��r�慿Zv�Q��x�Y�_t�տ��o����w>����z��w���������?���{���{��?�������?v��?|��?��§�yzڟ۟��/��m�����?���^�����m�+����߫�h~m�ק�1��ҷN��eo���s�~���><��?��֏�[1Ɲ��ɿvo�a�&������/��5�ͱ���t�����J�\���%��������k���kݼ�=�<���������������	�]���'��֗�M�p��-w�j��{o��ˇn{rӏ�^��+���gϱW���ߪA�7��5�[���o��rǖ��|��-�'�z��]��o'?������Z��b�W��N]�u�n�u���Ҵ1ӷ�}�{�y�^˿q�7��?}�����o�O6�6c�`�̡Y�g9tھ�w����>5����ko��-j[����t�qK�9誃o[��w���|�f��#ڎ�����;�裎9��s��q��	w����>鹓�?�S_]��io�����=�3�?�}x��|p��}t��?^q�xQr�'?}��]�Ko����O���+�ꨟ��S�>����~q�����ȍO���/_���z��nk��r�:���7[�6�s�ߵ��{���u���ܿ�s~?�����8��=鏧>���S�8�O��?=����L�ˮ���\�����~a������}������m�^������.~��7.y󊷮���8�����{o�k�k}8���Ώg|BH�#�Q�Zä�s>����G�ї�i�_{Ӹ�ƽ=�ܕ����ʯV~�ʕ���ڙ�����k^�ֵk߶���>����_��FS6^���Mo����/nո˗fN8|�s��q���~y���]�i�扵ݿ�o�,;���/W�[�=�Q���v�n?f�uv�b'�������:鲶_����o����&����;�N���[���ݳE�iӏ���=~��s{����ߒߞ�7k�C�O�犁�g<8��̧g�0�͡O�[mΦs���8�kA����p����r������J^{ل���~���C�v��q������Ǭ{���Z��<a��8���'|ʲS����ӎ��Q�}�1gsֱ?:���9����;��������p���s�~�����K{��.?��<��~v�Ϗ���kN����~�ˮ����n����~y�����<s��r�w������ѿwW��U�Y��U�w������s����`����������cW?~�����'�}j������g��������=��#^�ދǿt������W��ο?������k���[;����}�9����]��߿�?~��_�譏��ɇ+���,/n�$����]�b�No'�Ӯ<��wW�x���a��R���k�L�R�H`�k��$[�̱j�Ks����#u�l�)y`��������%�Z�Љs���־w�N}'���ڤ��������8-I�w/3������u]�N�������x�ۿ?���x�̞l�����񊜡�!�*n�Ff�����+x�O@����D���W���������M��Fo�����/�����o��*_��'���c��㎡�m�W��#g �N��޷S��a�! �~ ���C�B��9x�-��|K�_��	�v7����x��k>�b�|�x٘.;�LaaB���}�A�U�����߭+Aֱ4�m�'�lP���T�jK�$�����o��ȍ�7"����T>ukjA>����AYƀ[ǀ�	��ݴ��P7�N7W/z� ���!�)U���a��&��u~����X�~��,w�����\Ɠ˰i�
�>w%Mu2hQ�IԞ�m2�N�Q���c���\��ȌdD��q���C�&���Az���>$d����fh�Z�'���t|
�RY�,��b��O�!�/��Mg�5��d�!e�l4�W�1���,��6n������>��m>�b��;��bNV䝽�Z�V*��zZ�ۻz�vW[�g-�3���?gh���EC��U{��g.���^T�7s������2��}r����]g-\0<�?��������6���ӿ��ٿ��L5��I��d�:Ј�������v���T'��tu���X�i�2���oR{g_Oo[�$1��ή���m{m�sZGo{c���jc��}�Í�ޖ��m�}�Szz��u�M�6���=�h�:�U'a�s��v�o��Ο3�s���B3V����wϮ6��sw[�.��)S?�-=m}��o�X����jk��n�ȻuL�Ԧ`�X\_�NVm����̘�jmMp�XZ�R[˔��4V�L��l�h߫mR_�Ծ=��4�6����X��>�mj_Ǵ޾V0L�n�m�:��kjOO�Ď6�T�؆�����胈����Lo{*�K���Ϯ6��T�[���ՁP��U[q��gTZ4;H�Ty��l�W��ͨ�'���Se����͝8�����6eR�ܕ�{ں��A2˳>�4HqbGK��B;�G��6����o����l��Z�X٥��7��x��}_�Wml���tN�ڻ������]�z�v�ֆc�6N��m�{_8a��5u
��}��V�L���݇�����1�����'�����L��[�i���pJA�������u5ɾ=ܿ{��rB�{�=m�=�L�sT2�v����Z&4�#�dk�Sa%�Z�״jT-���U5�Së�ո0�����|��OV���g�"X�E�1+MZQUvSߏՌPR`M5��Q�)SVWtU���/c5�,SUY��pK�	&S!*&J��%3�GGX8��S��ظ��~R�D&9��(-m�*��J��t,�,u�gBXj��GF+�⺒�И�?v4�yVe�k�a�c��d#T��Q�Qe5w��"�i�0��2��T^�b���Yn���2)-��M���(;��1���"���L1[5�$�}d��������יѴ���(Q�T�1�����*V(3E��A�d��8F�4V�Ɍ�c��:�d��wj܎>K@����u^� �h���F,˔��g	�	�&B2�II)�
���DZF����f������D�љ�)��ĖZwdҰ����X��L�-�z6)T�Å[�)�Q��pH���� �ɌT�&d��Y-���:S#�z��!�&�f��c��3���VO` �rͱZ�o�Z�yjmN!�0jR�z�՘4�\b��6�*�ak�����$U�,�*+p��aF�jR��	N��\#�q� �V*���he���5�2)�r#`��=PY����	I�]O��X�m	��b�ؗ�}a	Ο�贄PX2�P9U#�ġk�R�
[�X6�hN;�#�feʉ�ڹcq�O>�s��#��I����N>'��N*h��,�B=��$�!�Ԓ|)�Nji��n�c&ͬ'���(�p�b�Y��*�5o�uDF��Wd��֑��d4#����� mWp�ďȝ
Rc��0h������ؘ�QW3�0PZ���P�
���{������V0v�c���P�GW�4��)X6l�,��.�9X��
�!�
�9�[G����9~��;l�(HѺ�f�S-S�e�)!x p�
6.!j�T����(��?����g�(�����"��U���6U�TBR�
�#�g�k�C�GX�)q�>@9�(^{^G�PEi���p��A3�6��[=� �i�������a��hH��K"�:�+���疤
5�)Ed@%@�f�0�Ԃ��@�pĄ�2�+8#�j�FZF`|!Nj{���6�8Z���7VuA��BpO%N�W�)��J���F��* M(��JI��p\���mf��RZ�@�H�X�V+1�_G��Y/!��R2L�,ڈ
,E���u�$G��¬�z8;�pxX�2�����$M#,�(nY�$����q1����% �T��qdX���i�F(%�:��f@V
SK:@& {��ZJG�CiZB?&9��ٚD�68����#��B���Bt *��U-
K�YOh�m�f�U'U�ۑ�`�F�wrHaL�>��@dX*2-�aF
VO�&a���dH�Ҍt�֎��0Π��a�a�{p+`W�ϑX=��4�גpp��wX�EE���!&: u�"$\�%,��(]�5D�����ı S�c� ��)����W2�>��E$geK2��[��4�I��L�ɠD�ӒL��H~�4�L
���<p0L�_�+Dֈdڥ~��5���e{���*e����8t�đ�U4���u�b2M^�B9%��W-�=:��Q��:H�'���j*��b�����H�#+ ��'C2���U}GA����#�t�^
�uI���(B�(��(��g��z�-�'�X*2�|]8aC���
$\챾#�#<�Qsʩ0�Ó|3b��%eq UC�AHڎ�,EŔ�q�9��!�������{8VSVȉ'�����J���LX*/Q�(.8C�����<�BF�E�!GqQ���cF�f$�.Z芑%E��! ]�<���QM��|ᨒ�#� �t��
�����[�*d�xc=�g >H�E���H�tMZ,Ք�1�����Fy�&B�V1��Y��%�֨\J���nIu'�i=��u D�����Uj5:f%�@�`�P=red.��paι���� eU�:p���:��d��/�� `d��i�@x6+�XZA��?F$Y\80��2b��T���9e��UB�����P=^���c\*��8xPޒY!]� �V��Ǒ
��"�{��b��2:S��& �!�:�hH�(�� V�-q�EGAZ�H�sN
7I�V�Ҳ�S4��"'g�z
"�U�Ҭ�g\,"��J���L��|�
I�GV�Z?�MK�F�\�5�r���K|kT�T��|�����@��%�5�pF�.��\��\GU����\�l8;CU$��'\zH�=���EO���\Ru&���qFs�U���%�=����� ST=�j�EONY���*ydEU ��1Z�-�:~��6p�)%��r�YL�d���b��e������9a�Գ��{6v������M���'+�& 08���34�=y��D	Q��a�������K(=E��B\Flir���irƥ�lG֔�{"IǏ�'�Hwa��o�T%�&@oq��q��ʼ8_M��%3�ۃ�b��V�9��&S�l*+�AظO��lJ�3��L=��9mI��R�|"	@LU"CY)���be
0@CN�ƔH��
��²��b�p����"�p�1V�5�e*` -�s��6N�SF5錕=��� ߗRM2/��:`=\`��g$�p<B9-U�Ud�J��%^3�SQ��rߔjT��D�r�J�f�d�v-�Ne�ڒ1]�5�JPq�lؐl54����֔@ˢ'U2*i#OE?
��dX����k�U02.:OH�Q�N%�IoyiS�l��xIFu[x�n�>H\�����)*�k*�"�PO%��J�Iт�)�r5Fኍ�)�`ٜ�)z!*N�*�@aX)=yL鑘(�&QBS�Pw���fS������ğ��fya3��ss"��<y�����%'8Nk�uC@���� Jz�����?���\����l6��T�'�/����^II��i��lѓ�}�]	XC@N���e./����?9˔�G:Lm1���\A�	T>���y�U�'�,�����9HZB`,�r)I��5	5԰�
���5��ꎰ.W��*�ɍ��e)|�I��)0r I=%�������V�5�
�R9^I��=� uTCr��X0C���2Ms��}Cڢ��R�l�}�O�Ӕ���27�M����C��
[�oG����U�YQ�Ӑ��e�5�Q��<5ݏ �q�!���[f%�6��R�EO�$=p��D��IVҳ �
�vT� �ߑP)�[�K�m�	T�b�S�`gy����S�[��(�
hKF�`��=�Td��~����]ʧI����Jz��39��T_�G����2Y��>i�,/=��J�?�GOS�ocO*`[Jv32q����0�Q��I�  F�ψ9=n��JCB�4u,.Уz"C��j��V�a�L�F����B�\3�S�+�g�%��
�8��È��`�);��)^��O{��y�f��H�4^�%D�J;��pY��H�M�,�a ��E*3����jUYRU�kK�\:w��9���.U�����n``�0���m��}���7R 0x�D����C�C_�!e�BX�	˥{% R���(��2Oغ� �]�/��'�YHH�С��p?Tc��VL*���0����H?�!��j#�I�:�r?�8!������TN�tY�4ܕ�'�7-J�1�r{� �	��T==�AX��7�DQAf�f�,.�U�&��݁�4�dh`�SWa{�/�_����{����IlXn��ɪ��ϭ6/r�a��q{�6ς��6�̈��-��Y�y �K�U���dPt1D4�;`����DO�讑�HXmރ��5{�������?wh��>&��x|�������}F^���*K.I��K�t��������4�:dP����H���H�#T ��{�JIǫ�S~%y������ h�/��\+]��ܓ\�Z�R��x)���"���D��c�����U�hϵ*:u�I���"x#^�������i(�ʽ���v{c:��C�-F��Z�I�����YF����7C�ܓP>'(�6�KK��V���rNbk������(�V	hH�ؙ�� xG���'vҩ'3����>�@J�xuJ��]�ͰObe~9�N<W�M�|6hDrR�r#����f�5�(=i��$N �t�HQ�o���M^�j�#�*_��õc/�A��)����O.(���� H3?��t�x���4�<	8�G���+�$\���f�̌_�R���r�p�9�?BA�7�F�T9^�2g�)��'�Hs��HL���8A�� ��ۚ零,גe䋤��61��taF伂�3g�������ʜ��o�z��V�F�7+�n��.3s���K��]�|�J��Ѝ�8�;��q�/RYDG�QE/�u*�Z5L�g��t�Ϗ ���,7͜���'��Z�x����r�.+`�ĩ�n��Q� !�UH&o<��7'�4�U�+��kԊ���@�T��eF�����^+h5�!�;^���{�X�C��C��� 9�ίݑ���@�4��u��Y�9��+H/�&�nq�2�	�ȯu�d1��+9�M�l=7�)xh�T8��M���>a
E*���b����
�IhWn�E��j$S���o�.�K�+��X�R��
 ��"e4���ר���?�"��I8O��+DՉ�Aa��'�:�zI%d����ݞ�ys��[--���^ؓ�Y�\�D/H�DR������b?~0I�ϓ����C�k%���Q��y)�z^���!E�Γ�%�$t�xYD+oR�@f�P{�y�!?�%��t{*'c��%g�[�t ��n e�������O�I�dA�G�xe~A�Z�~0Lt�H�����ێpL���T��*��y��`B~9V�`�y|b���<�E�k/��כ�je.�y�Yo���qs��j��
I3�I���y������g��z}`)=%�y�������R��/a�[-��� )� S���]�k�>�_/�f�	@f��Y�0T�5�T��@�ԯA���,�K�t�5�<���;o��̸�6��Ht��r��Z�]�Ԇn�3^s(�Z�(Ȭhu�s^�_���w� Y���cO��10	�)�[�)�7r~0�% D ������A-��)��L=��0��n\x���@�5�)>µ$bk �6d��Y0�	r�y8R�\�<bFK�ޜ�U�[`F�@:�8�!����pR{�����GÌ���	�H�<o�a�h8X�d�4>��aA��y���*����!�����F6�*�y�0ٗ�cH���Z���a�n�$O�g1�����P�D�j����Ѓ��7���"��{$a����6b��-0���2�;fȨr����cz��@fao@�1M+��9�[�V+�z#��6��b����O���0ئ��	2�L�4�g���0�KY��GHNI��[�0o/�p��yxeP6La�#$���pł#��@	£�z1��}��ȴ��ĆxН�a8%�~�Ȕñ 'h?n�0nһ�i�:Sx�2��@r;�!R#�a8��c */I�a=o�a����Mʤ�k�ƹ����0�),�f���խ�Kg޽�.����<��X�v�#� o&<o�a�~�
��o=)�q#���r  ����E�"<�'2����rވa�kK�Dz?)�=��@Hʻ
J�6-��T�⁴<�J�x,"�p�Ap
>fa�J�q#�4Ͳ�aCʺ=�ټ|#�����D��*#�F{���2�w
 U87Z�_o�0�|����7S�,�mHD5U<�Z�CNJ���a���y^)����SE�04���
�~�>:�y��a�=�,�l�y��H�b�<����d�tg�������^��0��>���a��� ��ԍ+-�����މ	XH�T ��ވa�+B7��@B�r9Ȉa�o� �ӤB�����g�ܬ�,t���(1t@z�����Ւ
��>Ȉa��ZRp�*S���1�D����o��/��LF��5`p�������`��JŞ�м"��T;��rO���@d�0�����
#�u�[`	�*�*�I+�<VFC�-�@��W�,�Sd{��^s�C9o�a0�I�$G�y��?��a(���i�f� ��a$!.H�2�|<>��H�_A�*0�1�:���'Dw��"�A���R��{�,#���)yH+�a>���H�.���9I�L��"b��0.`uX}�Ï1ZC�����=�����:tCLR��T~àU��
�WF��v1�A5`�q%|R�HJ��,��4-�v�y3r
8���W�o�a��PI�,ر�F��e�I�:S)���Ak���2:�"��-0Z�<�D�g��sSà�����������yC�}_cR��>���|MAE��>H(`�i�k*b���_Ae�O�gY�&�"��O��@���1���BE��)x�R��ރS�������x��OY�:ӾN�"�Q���p�W�l<o�aEw/>D@�;�U��8*bEy��K�t1�x#�Q��^ri�~�=o�a,(���8��vz=�F�~�!�T��G��y��Tg����0
��?'��Ǩ�6#��v��/����/߈aa]0�B���X1�,0hHj�*b���^��@�P�R�`��0h܊���a�~�O��\�n��>1��9��t9�y��(k���7S*6{���е��`�' ���#��pm~o`��`0�sH1�Ί���{Aj�uRGC��Ҥޤ1��8UGC����T�����a4}7U`p1'��up1r���K�ky����g:b�|*��^$�uC~� /1Lx�����g:b�qo�#�q)�;�h�>^5�i�b�3���a�^�Oa)�
$�g�7bL!y �GP�i��-bL�|��y� H���1�PޭhE�<I�sވah
xU��Q��c1C�FS�ɏ��w�1�~R�TC�1KG�)����ݐ�r���a�<��C87#��/t�0T����i±y��#��!�j��?��M�wL�0�>���[�U�L�0hUAa(��Wf�^J��0huO�2Q��U��(B𴆊$���+ӷ�x]7�P�wx����t'�-0�zC7��0��y1�f��>��I+<^7�P��;�$�{�D��"��V$���SP�e1�c�Fp�H��&b�
�4�
�M�P���-b�J_7d��|�Dcx�쀀����j=~�à5�����p ��^'M�0��K����㐉*lP�d��&b�߇�TW�����>U�ݕ�a��W.�u���;��F�1 ���&b0J�@NH��xC���� �I��}��Dc�{����k�����DCu�`8�Ӡ}�a�
*�=�F�c|��D���zhv:�q�0����w����R�ve#�!��^+��QXl�-0dX:�V�[�AFxc�1e�!y T�9[��)|�l҄q��ue1��/��l�O����xa#�J�>�b���EK�Ҭ�-0�ʐgY��#?�Kp���06sϸs�4�4��h#���4l��C�|l������\�#97�y��A$�BH�y��t���җ���s�P?e>^f���}/,�y?��S��>Y��
Q����-0��Jc�P��;��[l�0�A�0�^�2��8��X�ҍ��B��7�I1��YAH#U�Fj#���c���.Hӕ�-0�h��?�q���ECu��7v�����ك�MgA|���6b��p���0N*�-bk�2=�N8Һ�Q�[`K���y+?�Y6��.Z���k��պ�3^�N��� WuQ���   	pHYs  %  %IR$�   �eXIfII*     (           >       F   i�    N       %     %      �    T  �    p  ��    x       ASCII   Screenshot(/��  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:exif="http://ns.adobe.com/exif/1.0/">
         <exif:PixelYDimension>1392</exif:PixelYDimension>
         <exif:PixelXDimension>340</exif:PixelXDimension>
         <exif:UserComment>Screenshot</exif:UserComment>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
����  ǸIDATx���$Iv�<"2�ή���ٹvg�b��hF�J&��Lf�*�>���>���H`���ٝ{�ﮮ3��p��;�=�2��fz�SSY������{�7]�E���s4�O�7���A�h?8B�>^�HkY<
�w��G�_��}�� H8�:��ȓW�x�g8�9�>��ÓB��El҄ z��Y��;�[bϧ0gP�^A�hLQ�5Uv�\��nru�@_;����9��O~���]���w]O�ŜNNNh>�Q�u���3�Ni>�1��J�
B����x¿Gc��Q�?L��ф&���J��z�o0A����oi:;����� ��ތ'|Ѷ2����9::���}�p�&�ի�hē^U���d̄�CM�L���m��ݣ]�=ij��f�|#	�&Т[��Ǐ�	O��l΄��ʟ)!�u۵���*T�߅O�>�G�1�z�|�c�'�an��],��e�4��ss����6����b¼|����7M�,������ղ:`�xzx�Y�)s�t6e"t�!3!��/���%������d���q��mnn�(�Hk�3@|O��?�}ʢp��N�:{��{�0|(�E��F��bd����E��1����&ƂuH+Z��T��pV38�.�(�A?3~o�?��)_�����f�Ҍ��ڢ��ѽ���ÜRQ���oq
�Y�a�ȑꂕ���)�9�6v��1���ų�zs�0,��YO���	��n sY�u]	���P��������<T�ގ�p�Q�� +��9�<��?4V�)d�H��T|��mml��/��J�a��
��K�;;ۢ����D�=d�r��]�L\�6s����X_�|�����TP�u��o6A���Eʓ��+���=���+��W��KL������{�f<�@N8�By��'"�	rt|$bp�����Ç��`������}c�i�#�5�O5�*sk���+���.ݼz�a�X8F�ȩ��$�1yc2��fE}��u�tbӴ<�?�?��?�����;����p��o���GTc\Pӫ/�B/ݺM5�+v�����L�Rxܧ���!����A�<������(\���Zs`B��U��oP�E��P�v���VxN���9�_e΃�`� ��"�����7� �'*���Zt$�c1�g;9V���U�#���ǢpcB�|���l�l3��Q��~K���$�rU7`�*�1=!��`L�t�#�_�儰5���-r2;��!�z[����E�Jꩅ�� � ��*ӓ���X�#�m���>���d�t����9���3�y���ٔ-�y����.�>��	D����Gc�(�&����.�{�ŵH�1�<Χ�1}!���2q����	����>��cz�����^�I�s�y*�Ť�?FT_ܿG|��k�6K#�*7���A�G{e°��7�������?��7nJ�̑"�@��(�/�_����4���ǂP�P�q� U�������+$.�2.���M*c��K�m������������[w��?w�n��5�W.�X$E�;��&�q>_��ֶ�#�⏂���	�0�����0tq�ZM�X�O����
#>���|e�Ŷ}z�`�����L���v&����b��{ e�2aqs�ݽK���ّx��,6:�d||Mx�Ă����c���b�����,	PݼyK�w8gE�w��B�i��ϙ,&>�/�t~w\�f���x�3-d�Fu��K��N=�_��h�z/�(���#}~.l	(�$ܺ}����Т��9u<�LD q����G��FB�-$^a���FL�_~�^~�U68���rΌ��a_x�ga*�\9AVX�xO��U���e���?+	s|zBs�j�`һh��&�3:�XT�!�}��T���	��F���ߘ'n����Bxiu���l�!V�Xt�1(��R4O.�jT' 4cV�x�k/�4L����(�$ $4l�P��Q�͈.s�����tFǰV�9����R������Hl���3/:ԏd�I���I4&F����[k�	��>�>1k>JЩN\))��#N����ʘ(�<[�a�reHb�r��ǡ3`sd\j��"�ܢ����(u&����:% ¡��b٘ �r�-��Gq�yP)7�o�: ���KB��r���0
��Y�&bq-�K ��Sх�M�:��z�4����ct���ϫ��\	��U�y4sI[B�/K�ѐ��a�C�R W`�c%���5�AH#yv�9���f?������U2įdfm��wo"� �O��y��#-h{kK��V�DW��$^b�-���r[�9�7�}�'�)x�[x=
<��{t�c5AxP��N�Nh�ga�6xh�(P��d*C�Zro�� �lY�KsX%�T]��X��\���d�0e�������'�W�������M����K����������� �P&MƄ���𺣖&�?�;}q��N�@~��rP�жQ�%'�C�\�4:ɑ�� �d�yR�Lt�]b��-��bF"�@�d0�c�����|��xT�J����O�Ν�d�5��J<���)L����f�h�b�Kg�>�V�!z�����&B��#�:�	�_i�!XS�k��R+r�i���>��666��W_�����CU���H��JuKWB�>����$����H�Iq��-h�sg�
==xJ�!M�J���1_��	�D����E)p�尞HC𢩪�c�恣Ưf�x��ұ�Oy�AD\��K��4���.s?�%uE��J����9����"��{��	�Z��,u��R6 �cU�h���,�3�&�[�1�pQQ��Z����x7X�x���Ǵ����z ��8!��s��+Yf�x
��&�1`��HT�W*f]��nȗ)��"��.�F�WI�{n�b��I�n��٢s='�8Ӊ.�ϕ+WD�!J_�qCN��R�$O��C���1�nHDȋE�Y�p��,�7!2���I�'�2�7X41�r�*qA�p����.��p�FY醫	���zC8�$/��SLi >1���rY^`��ݢ'�.�h@M_'B2�B��@Q�Ϩ5�F�Vɹ�EsIYe�j�e8�9d���ɣ��@!����W�Ĳ�JX��U��r�ؗי*C8��A5 UAg�$nY��&MP2TWf�+�9�y%b��Գ\���,#�L5��	������Od��� �k��'(d�g]~�4y&��7 �{�zU�A}Sn����>m�h�ِ����>�������}��(���M���qO�&HWD�(�=>9�����ޡ�W�"�ϲr��֓1cr�����"��t����`+Ox������ӢKˉ�AFP�FIN���|�k�Q���C]�ɟ�JBE��P�3���B�]6<���}65� Āa��c[O�g�*9���*����pD^��y]%���j��?���|�,)�����4�����mߓ$��d7�5r���q��Q��8�)Q�'��ұV�Sz�J�y�����zkkC�+=L�ɜ-d��a�lln�R=|�T��Z�z}��� �����"������ə�B���������r6޵|.�#�m��+vʥ�9�q-�
��'cqa��y�"�F�M��G�.I�5�������+���(�&����܋�wC*��C��CD�1���Vc����> -���2�߰�aԁ����~��)��H��K=����� "������+1whq���l*��|�pz|D'����,��+爡.�b��\T��Y�2��0�uX-9�t�mmo)f��W &��p(������J0r ��&��X
�`ۻ;T�c�+�+�n"C[�][�#O�<���C���T~f(Cూ��PЃX�[��(��c|��U�.�[��ń1��
G�1��L����3�1y,���Z4��V;j-���ȃbՁ(X�""�Dd�9(9��ꫢ3�P(<�X�{{Wikg[&�\��K�0:;������}�tX�O��������c���`Ԟ0!��, |�T"f���ի���_�^ ;�7
M!�I��GV%�*�@�@{"�(s��s�ITȨַF�0yw���ϱ���#���Ipk.���)���xX�;L &f�t��^�f+�SWM�א���*���Z 5�����C���������O���;�����]��A��[	<b�=~�^�s�^z�e�q�,&����]�F�PW	��	|q1TƵ�(��~CƢn|�ɾpr�0��<��I��#�|�(���G̖;q��@<��۷�&?p�"��	�x���g���E�� �yҎ�<�O>��~�_�o~����L(���ߣ�B�)s;)p�����\��c;x��N��B����z����W�\a�>���+V��~�L���ļr������V7����7V6V#^?z��޽G�<���B��~�7�HP�E��M�����������d�H(����I��=�Zv�7p.������k��O����޽�Ro�_�����L�I<����t��=A�o�񦈹��{_��.���>f�vI?5�͢�⋲�J.'W'_ٹ�bʅ'���WT;&`@<����C���E<@q޸~�����M�{e��rU��i�_�<���ҟ|�1����-=dN��;�0���c����I'�B|E���8�U)	� "���O��#�޷^���wK��,��?~��P�h��Eses�~��~@?���D��g���'#)��ؘȂ����$���ʒ�s���	C�xˬH2���\��>sB���O>��>��S!��^�W^yE"f��)]i�D����ݱ8
�88B���@��/>O�Xo�����?U�2�OFX�%�&z@�/>����/���C	���#��1� �{�!f16��ڵkr= ���(O���/g�S0~\�	D��jĨ�},;V�X�����B��Պ�fu(A�	��?ؿ������w�cA�[:s��@.S�߃8�W`����ŗ^y���'�|"Hv�
��bbϘ����_����i~ʜ���=z��!�`p�A��b�����8���7�8�}�&^���p=��
��d��t��f�;��2o}ᠤ�C���:���ON�ʂ+0��ypX�x�	�	i{��6�`�#�T�� �b=p�u̽�w5w��	t�)O�w��]Y���|�+qc�ĸ�G[&���n)q~F�/�����E'�o\��vö��77oܐ �'�X����a���Ct!�;`���r���|��y,���( (������G].[�"Ab�� �@�۱�Yy�ޯ~ŨE{��^9a�|��_����tN��) Lu��WĜ�k(k������$�u�5z�����?W�΍k9o�_�<yN�t)���>��^�U�!+���pL����5o i��a^h�x��[�fx*��_bpp����<~��������S����x.�}׺���I]��Ѡ���H)�ho��!�0�;lW	F��z��u��}��Ǻ�q���Ao޾�,r�o���^~���������WR�4�x�2��\c������b,<�n����g,j`�� <@t����PY��}4���`��8�~[3�>�ЗDY��C�ʋ���≸��L�'���3�dU�uֹI�}E�>�:��� �e�z? +qƱ<Ɗ�����ؚl���҂Wrz�e.&J�l��W����X�w�z�-����N��Sq��L��(}A����Z&
���@�<�ڬF�8��a[l���LL�L4,} z�w�b�O����ͯ-�q�<~�evF����I���}�a�O�ܲ1l��BN�{�{��������"��_���y" �o3���/~�D��av������f)�P���S0Y�*T��f�,AC�Ufb�n�ꄛ���N��k4�Y��u��)�)ԗpjP�Po���,,x~A,ɨ��]���>#)�^��\n�/_�#a�L�j����y��'���'S�Lq[�`QN�a�hl�`؈�-�M��^���$�.&m�>��3�Bh�d��=�}�����l��9jS�:Ei�(�>16xR�����LI3j�P1U-4A��O����Zý@D�ۛB$)�K�g��DJ��ڌvKی�m���_���o�N��(�����ՊT��4�^���8fq�ڌ>g�E����ӎ��=�ʈ����x���s�5��X��3J����Tf�XYA��ύE��6��g��m�G�V0�+<�G@5��Ome�S��H�L�t�ސ��ٞA�*�ߖ8~-�>V�c����
�ؒSVr�jI4@��M6���;�)�'�����n ����ߡ�_�5Wz��n�}j��>��b����X��O\���hEac|��;2�O�}�Iu|n��r���}��GP?7�(��,� {�}�Tϋ +�t��Cf6&�eR�=`t� �F�t1�x�gG�(2Zy�7İ���g_�O��oX�?�*��}�{�j�� !<$�yf��oj����3|o���~�0􅱩1��x�5[?Z��T��D' �q��%\����N���m� �X�����[�!{.	��Cؒ�A��9�)"	��3���W� �
ԅoAΦP*?�_��>����k,.����w��TU���$MX��1�rT)n(a�^�1 ���8$9�n�G���[Ҟ�n��6x���K�Ӆ�23�?�VX�Y��b��J% �B��Zy�R�~%�~e�H�I�,�^B���$�X8"	��0UjG�D���T�&1�-���&O�|!py����{t��)�?�������o�K������Y+U8��خx@�H�e��'�`g����؎�h��7b����CD�0W`��|,�ƒ2���0�nr�b����M^`*b�a�ci�)��n4g@����#X��W6����LV��#�����M?��OduI�a�ڪ���G�lmo�_a�y^υpG��� 2����}[�_���d�a�v[Z]�&
q}�����q�!�^�c�'�g!� 7���<�c�� C�J̠���'J��⅀ژ���b=~�̮^��P��A�=gS�.s������?���`����������>�7�z[2Fn�D�5�����槴�l�@�A8:�;��?�w�N�X��MQ�����˯�B/0�x~V)	4� r�a���w��\�3::=��-�ܞm��_I�B�@�XD��7�^�-�p.$�B}�Y ����W_�#6��M���M������r�:�'`���K�gFW����J�ӄՄ��3���������o�@���>���[f<����D�Jp�[̅/����v8"յ�[��L[��]���/��~������?	A���񓁊��Ap�/#D�7��D���L�;����`|���bh���H��6���Ap��Q�� y�s����=�^KJJK@��m'�����}���������C&�(XV�s�X3�j�E X�+	���߫� ��KUB��I�������������D��i���P����ċ�˟�\�B?<��6��D�A�b!�$�ϻ6�)����G��;[t���P.�����LH�GN�[�[v�P��J��	?R-
~��?��M�����|��D������s`}��w���Ġ!�g����7^g#�����<���{�Ͼ��d  ^ʅ��v��֑�� 0�/�տ�{���1��m�#*��oݠ�c�C�}����5�� ���g���2�T����w��o���gn���-�RX�M�$A�
���u��{V0�&UC��H���^`�o�)+��u��WX>���_�k7��ہ'�֋��ã{��­�����/
Zdz�n�y<-)�"�*a��������/�����^�Qz`���7/<���0T�����>}��\{����?��pߋ��l%���\�9�����q.A��ue�	b�z�k����A��w��bE��?�Gz�_��@��@�7�}9�2nؒ�[��������$���������B�eL���[U^���`��hr���,2��B���G����O�#{̡���gn��(]�- �>�HԸ�G�o�F?��w�����/��:R{��$�TȨzE���%ɼ�J	�ߐG7��mO�>�������?f��%��?���� D�泩X��$ �N���N���������N�r��$e5#):��e6.��Z����ٍ۷��-��_��x����?�1Қj�-�? @$�!!��<���">�dD	��sb�H��R�x�/x$��.�F.�:�+_���͉��|T��Rƃ���?�_����|�Մ6����6�Q���.b��5��M���=ԞG/G��c�y_H��b�be��ٛo�E���=����JB��|�$��g�\�1|��7��̥�� g�+��E�r/Җ9Mʏ��~?�CB
�g��J'eY@Q�s�޽k���86�����*�����s��ce"!0�߾���&@T�7��k������[�Z��\w�މ8+���tX��~�;�o�����a����Aa��G^~�eI��v�m��M�؍&�F�}�(���P� � �~I�8����T8�r_W�����N��ѽ��Lv
�[o����@F�SP�#��������#$��w�O��-��Eٵǲ��Q����2��(�f1�}�;���;.��#+D�k�m��]��">�RW wU³a��<������������ڝ�paY�	0�6��H�6t˶�N#�5�D���:�4�
�Ţ��i%k�o��B鲇����ؼ��>� ��r_CH��\���:��^Wh� �$Ҳ����[8��e�ेT�n�+n�Y�.�U�  Ψ���e��k�D��A%�	+��ioew�F7�2��+ԥts��X��H,���[�)��Wg`oL�E��U�,�֬�����;֢,���D��v�o�X����U���e�2��[ۢ�և.d�L�Ք{�`V��Y��u��Q��c&�-�'�锽sV�eo���)������w���YC~�}������E(䖀_� �j�k~�>������U�<��D�^�T4t�+�w�&�+����r&y�t+2����uq����<�%)�A�1!���?T%HO�ABZ�Q[�4-��(��EN��$}ˋY�`�_� �(Q{��]�#��z+[B�Zc���#{������±��*:��6]GA��C�I-��e��t��ظ���H%��V�lib�SŔZ{�g�S�~'��_]d�{���C���)W�i�25��I����J�%��D���1�3ܓC�V]��r����=Nj�䟅�8!�X+����o�X���R�DU,����9��{>b�&RF�h��^����dj����+��	鰕M5�I�����yw��
�	������W6�uA��;��r\�mց4\��G�*I[jP��ˢi�y+�H%����`[ �<������
4��řn�����C�Mn�`};i,+��o^ޣ<�a��s�w^(��W�Q�(��=)��瘣���P:QS^=�*u2�i�S�t��:�~Mz#��??��ׄh�b8A��N��1�χ��6���j���/3	��!t`�ڊR�2�o��Yk��ET$嚑S*Qv��)����<��M��,�x�����>2��t�`��E��G���2��ϋ�K��^+~)���W	���Y���YUt���A�[Ɋ��1ĳ��pE'�ťP��%����#o��� �OZ}��� g��}���_#�[�DRR8e�$���v���t��Q��Z}�u���@�\����*�9(�_�l7!��-���t��!�M�IG������ϼ�2��h�|?駸�����j3���y���[��s����� ���a&�*d�ǹ�.�!�?s�$�}<���]b�=.2ₔ��ʥ|��t��gM�B_�{���7�xn�2�[�MT������eb+_ױ>�J��D���ɸHg��]ĥW�ԗ���и~�N�e��n�++wώ����c9�0J~v�!�^���%���x��n����#[X�AC��]5���p��]�W)�"p����YA�@�f��{H$�G����|f���g*�����:<���Y��o�B�������}�sˢ/�)#������]8gb�۫�SH Cq�x�e�9��a�������q�\�M:���%�?+
�V��|B��
�LI��Y������tDg���g����6ID��s�c}к.Ëg.�^�����7�lQ?�Y�y��.ow,����N������.s�{��岾ş'���E��aq@���8����9Xɫ�]���_u��i)��Ķ���znyK���9%m�OKڢ��C���Zo�0s�?�m�R����#b�/VF��]t�r��O����.��c���Y\�x��z�@۸|~��>5��Ĳ:��]'�BJ�;#V��9s#�o�8'�zh�����2�xdL&�}��AO����l�h�K�Ń��зH��������Iٚ�qY}��<c��0Px�2˯д�d����i<�C�O�il��_�������-�pF^Vq�!E
�Ͼ}I�<Cd�U�:߁�ş���ϲH;.!�pH�OHu�ϊI����r6ܸ�м�8tT.�,R(>S2��3[���Y�c&���I����yw,\$�~$$�k����-]9hh���J�%��@fյJ�}P ��]�r2\N��l�f�i1�"-W+�jh{�;�3Uw��V~���2i�>K!Lq�'��d/��6͉�-��Uֵ9�6��2x�ٽNV�y0��zXz�4_�����6��5��(<�̶Jƥ���O7J�i��K6��b��Q#��R-�ͭ���	��sj����{ai6��q�w�@�[EV	9:r��4{����r����䇳r��IRr��3b1!����r9[��9}f�<���w�v�B�/��S����I�&�A~g�b�s|�����+����$^���~��a��̔�Pv/+�s��dm�ѐ��I#8���B�9Y�t�Ϝ��}ͳ���&p��y�i���RiA�0��w9��vw-y�zo��OX�5�gՀ �:'�n�Թ�*�B���s��,7F��)WG	��l�T��UH;�{���i;��_�+D���	O/�ՋY�}�2�k�,�ӂnE+��]$<r��ד�{k�-z�����(�����{^�T�38��� ��.���0P��Q�_ł�tD-�������l�߾����[��ER�wu�D�uι_������m4��x�AdX��TPm�R3[�,Ψ�.)��[+։^�;L0F%�t0���pM��}K� b����ґ��W*����h�^��votc���UQ�鏎�ڪ����LD�g�����&�;q�n�޶��y����j���t��m�f�1��]���'�r?D�C~������E��w��mp�ŷ��M�����K�RJ�BK4��?P҅n�*"�vC�G�� �W碆���{��"ֹk�t����Si�!��G�%�t����(S�h��ߨ�G�H��*�jk��;��@����I��믿&פX	�5�Π����F���r��zJ���r�1�����1m^�J�3����dF���-OS;x�L՛�o��u?©m�����.�x�)�����^[P��ڡ=��/D�m�(wB�!��:��*�zhT�"�\?>y"��\�����JŽ�����Ûo�\I��q���wy]=��{�Ԋp�Ź��۷^���Ѥ��TfK�}#+���CQ�~��v��؞2q>��s���|��u��sE���A���}�x|@-+��1��������՛W�f��������������ͥR�6C����X�&Z��d���Fړߌ7ebd�;^/�������t��N,Pa��.��2+6����v�e��iׅ��ފ�BE8�1���������4���%��&�\&}ww�9q��=x�s�\TO}z��$�n�o�AT�v<�tr�m�H�-Ni�=�'��������H8�ڵ��V+�yU]��l�C���K/�@���ZQqh.;�$^:Cs�mG������>�������.�C��r�c�(1m|�V�A�tM��j�w4�������}Aw�=b�tf�/���]�3���k,�1�<�Fs��	�lT�-�t�s)�D6C���vI̝�+Bu�(���tK�H�GҎ�weo�&hj߷��Cad9!�U�*��^�"��K����H'��,��'{�O����G���B76�j���>��c�W���+���b*�. \�s�QE�vJ��Sِ�ʮ6���-_�X��ye��G'�窝3G��L�?x�7�,b4t���m�W�	�r�b���ū'��+ t��u�2nA�ob,��Ë�V{�o0����iGF�o�cL"��e���h�t�Џ�X<��O����H�.��[&�tz��
�nD���=�-�����]e����O�0r9��т��m�(A��cFs&��
�;�mn�HK��m���;�U33���e^�^DS���pG��r妉676d�����#�gW?Q(��N��\c������G�0�?��um ��4��\�/4
��-��C8Yy�!�g2���f�|�Mǰ�W�T�l��AQ(�@	5Ccl�-�sZ���O�y�u�X;�������AQ\�$�lpZ���ъqJ��J�-E����������r<�h <�v6����~���߻+���YFj7�#p?m�6����T�a�9�HB���\}�U����}�!�0vw��b������#�˖�dd#i�i�ؿ��{z���o�(_�ER�i�*�A)���H��ޖ*�Ѿ��Н�f�9�>l𷷞\U=O4�����W����
q�b��-;)��b�޽����]���x�m3&��l؈��bH{�/F��������EH�����)� ��uM�ܿ+��mb A�,Ʋ��DV�CA�6�]kH��DU�E��I�֖��c�=�;�|����G�����d�Ȉ�&�旓]������p}$wP��j�6�Ld%������j��ڶ��R���G��g���6���0�$�%��h�{����+$��P��F3�q:(7 ��|g2ސ��z�_(! E�.���o�9p���g:����x��dSǊ=�f�m�<�}��v�Z�
�k��V{s��H���Zl����!�H`g&�G���<����{���V=2�/m�:�B�Mnc5a�8����PWI�b"*k��M��j��%��@�e���d�����CF4/'U�c��6Y�C7���=*���K%������H_��;!o#6Gٍ�V$�[��6��*�˶N�/�)�����)���ĕ�m������d��Jj�4�v��d���,O�
�dW�Z�!�C��d8�����["u�>Pp��b�g`��Đ��W�ҫ�T�t�W
�^�p������Ψnd��@Owx�]�q�J�ʔ�"M�d��6�#O< ZQ�cSv�Q�)Ȁ�1 ���@p�p��eߘ�H��,Fl{���k%z� �>.��/���z�-le6��1��C;�IY0���T���8V:��5���a ������'�%�Om����-���5?����)b�U�X&i�WOu5�g�[�`��T�?�p8��L�@g%
�jl�:pވ�ȸ�N��Q�.E]�a���<�P\�T< .�����6�nc�'EF��3yyp����H	��0�vc��yb���U��9*�]���f[�J��^�L�m�����	��o�W��c{�Tf��uѫ��O��`a�o:��e ���mX?��K�V�P�>��	Z���̀y7O�Q�х,u5�h�8��?�˓�ӭ^=7��w�@_�c��7�m�v=::�A�t�5�5V#<��v�t)�"!��ģ�Z<�����8;��TBi����;����Qg�I�I���ݷQW��4���gp�x��y¥2��ql��L�y�܉�(˛�$���9���*�X�ط	�zg{��-�aU9�p�9�͍�1j�'GW�K�lK:�O�_�Ŧ#���2$�X3do5��b� �l.����o�����[�l��ZDܢ��c�U��֎n�Luwk��u�8�H��	b>��2��P�cV��҃�+���ϱlT�6o�`%��/�N��4���.V��3�011c햻ay	E�i�5ڇ�'2_��h��_��A'%����=�e�2<m�20)ň �X�Q��b���=b]�1駧3�y����������'],��.�C4�+�>7�Px��Q�¼��K�HvS���b�kyR�*�>�1-eEF���܃\%@p����R��;��͐w-P�Ge�C�:&��̐�;�W���-��!:������l�K�k���Z�ksc[�ۗ����GʢjT�b���E2;w�@G^��&�Y��ãC�zz�l-���>#jG���8��
x�����nI_��1�0�X��Q;�m�>�Ő�$�egJ߼�řl�'�F���]���wc�7u����ͮ�%���%._�LJ��e�!8�����A���:���vK��)��r�6Gb#rK�(63��bt�^Uw�d�l^;gzl���e�¥bPAenV��_f�hK�WKO�pg��ed�Y^0X��Ƃ�2��8n	�a*��AʀØpз��(�i���+�
��'#�7/�lt]٣��m�pVA�7����5PR=�+lG�d)[�5�J��5w�M�(��vz�������������DJv/��%�=7��ut%�m&����mf��3���ʍn��[��g$��GPt>e�*��Q������6$6��V��������U$; `��� .�m]7'OZSn���t�?�CI�59�M��f��G�7Ţrq�{B��G,�W��z�����(�m�1nl�h���I�%��y�ߛ[�	ek�Ⱥ�"�Cv+�]��沽����wY��H
��$1�?�r���U1	�d���w��l��gœ��0����!���R��H��7&�����EZ7f��h "UHa74aTV]k�!�C�g	��*)1�l�Ӳ��Ԇ˝ �ņ<�û<��ֽ���LYF��!�
�'^���?�`"�b_���?���h���,��H�()o��6�����P���S�b�g���{��+>�)�{	�e�*�mѠ��97`0dpW'\k�m��d�V��?i�� sҵ������
)C�?@�-L�~P�!#D.	���a�bro����`��7��i.{~�O㐑������]�8��y��5)�-|�H�q���½��鋭���˹�y���s�Z��y�Z�Fq�3�&�[E��^~��u��G@uZ0~�O�[������_�k@���:�8��Y��±�_��ڶM�����{��0��X�u�R��'l�^�h�;���х����ҵ�=�o���__����X�PY1o�g�E+��q���.�ʀ�3-B;֦�����S���9�==��|nѴ�"1�EN�7	���cik�|Aq�dQUܐ�@D���y�&å�S���=+#�Z��HQG�B$�#��u:Vf.�L�Kqu�+����,�RD�	.�z�J]�+��l@s�=�&�$fP����]�2ǭ$B�99���;[O.W�1��bR�]�C����S�X�)�Qz/���w0nA�p>_������m�Ήc��IVu}�0o}-�PO��٥�e}��e�L�x�l��ގ�#.����I���2�#Q�M����9K�\`�5vX+�o��(ɘ#�#�f�o��g��]�i;��q�\�(���^!}V�����4y�]$��*��s7+W���#f�!�!;2W�wu�NP��rJ�!�!���".��Qo��M���L��D�����
�V��tK�.�%BN�+z�%����� �W�]��f��ԙ����x��Zaz��:=@�Q�dx
N)����4��dD�pV&��Fhf��>��c�Eb��m/���y����2�H�*�g:xTM�̱s�'�ȍIu�6*�ڋ+	sֹh�v�*Z�MU)�b/���PCZ!]G9ju�JW�_�8��b���]��Pם�z��lW�m݀���Fѫ��#+�&.���9�����dz\�8@�N���%�G��"���e�EGT+�]��ι��`�8���p�u/w���XK�leD�� �C�-�lAH&�/�Ե�U�ΪnB	g���*̂�������=Y-{G�=31�� �-����`��9v؝D�E9K�Q�=@R�
8�h�m�%����)xY�x�������5��ؤA)�h�<X�l��\c�?=�&%)Y&�{���TI�L�9�+�Wk��r�ui�H��n|V�<�d2_8db��3��3�0aF�����
�+Q� ��H	���=��8=��b��G)���s������*|^Z����p@'3�3�NA��{-Y���L�/���9W�q8̴�ʘx&PFK�	�n{d����H�I?�9s�(�C��x��		�\Pda��c�w�\٤�{��4�(f���\�3S:}u��{���NTw������g_Թ�,]#v�Ɇ���=.O��
��K�P���m%Gy�Hyc�$R���!~nk��Z5�.n!���"�1��jP>�3g�au��&»7�ct#Y.qhݯZ]C�d�`3M�C�SU���V�]Ht��57����l��a�0�}"�K�^��g�Rﵴ �tA�Y���.)���!v�m�E�?`�/_K{ )%�Ī][��ZN���!A�7.�X��lp.�=�/Ti��}���6���k��آ�^a�_���m� ����jT�dH�|�D�W���}(�a�Bu
Q�����4��8����G�MV���>��=|���+�������Q*.x
�����]wf���c���EQ �K�՝MR���>HO]��I���c��Ƙ����nOQ���r#�5�[r���y��;�l2��m��=�4����
�S�A_Z�ꮷ&8��!Q��B@��I����\I^�Bj��8��J�AA��>Xs�HR��Q!��tf��F�C^�Z�Lw��IG9�By�h�Y̢���&���g��z	��1f'bL"�av����"7&�������ɹ̜U����
WAH~�!��[R��#���J�X5<S���|b�=F� Q�%��|�	qH+ñ�=_��eٖ)}Yrm�=O,�G��j>����|��R��N>�c+��Mr�d���ڹ>e��}����\����C삳�p���3�L��+O溭���ͥ�hϮ�<*�R�vȉ�n����Uf�{i��Y�.�{�J#P����.7�$��zI�S��a�+ev)��T �B߈�`��M�P	/
��2dNpc�Aa�����MϦ��aP�+Mg\_��:��U.�g�~.�BY8���'D[��(
.�ͺ5�JcyK��<]nq�b%���J��n��bN���@\��Rb]\��1'*�T�Ø��5�<�4���+4E!+�G���-��G�g�OxX������#�T�Z�țx��fa�z�����R�R"F)ˋ��Г�V�P��^&B��^�ԥ���jQ�����J���@��F�q����9O�K3^�H��>_�	㫎�M0M�yU*�����w6h��fS�*�$����%hw!eϋ6+DU�R�%���8�'e�t��	^���+{�H��K%w�˟!t���VL4��S�0x%���r7q�0�|��)?�"q�C��_� F
��XD��N����k>��fDG��$�2"b(� �N���6F3ea��fªc�_"L�g$C^�^�*{�]HVr40�(l,�TcS
�����9�C�~U!�x0:�U\�m�IHWkj6���oT��H�؍y��苲�]l?� Q�s�}h��A*�b1���#:A�%�Ç��=X)rm��9�g#�|HU��o%��^ߐ���SZ����s�e���mob�<�֍!�8Qʭ]/	1,s>XR��?W�����*h�F�$����?��৒��Tc����%V�.�.���K���0�^T�0q�Jk���c� "�6��'7�$�3Ag����'0����۬XAj�[��XJ(b4nk���l2�r���sO^P
8�X��]�R��X��[��l����0;�������"k�&�2��ʚ��OQ�L��:�ʩ�*<�������U\��8+w.�)I��>rC��gV�����	�I|iYC�DK�"B˂EY$T�q]�`�s$$����Nf��x�>�
(G��y#߱�(d����h��,��Y�Y�E� ��"B<D۵.���b?|��>8~BO�<�I�_WQ��G3�&c�Q��BJ���j����ȚsEY_�=O�sJ�ER��ԉ>!�����B�Q3�#���Ѧ0X �H�W#.n�,��״���J�U;�j��.z��m���3�b��1�&��Hx&ABFE�j5���%���'�bz�e]<0X�Pb����jP�+�(�g�͘����srY(::<aҥY�Babk�@&��F������I�s�ͨC9��;p����h���:�m��-JP���[(Q���r>�����"�ƩsD+�Dtr|��0�z�YdB��(�:�������\~B�X�>������&�vĞ��0=(<�I?9QH�"I�]kU����� 7�V�
��Co��xq��/�)��m /�Fa���V����h^Fa���{i���Z��8�L�gjm��R�kb
c��ٖ�׮]����'X*��_5nt1�ҵݭ��.{��T�_C1ml�⁏Y)�Є���J��E��^����}z��q�.�#��Q�;V�I��#+�� Z
wk;�ɱ���Q�A���WA{��E���7���/zs6�������Fe*�P��\LB<aqI#F�����p������^x�Ez��ԏW�Z�)�5���s��y�£��Q�,!�O�lR͊mc�M�͂��ڹ�r|�H���߿/r����&�&�9++��M�w�"9�أCQ�.]�V>͜1�TiU�o�Ҍ�_�$���f֛r���5��	�"D�d=���[��N�f\)�֜�xH���O���H�	�����9���xE�۝�e��v��넖�ѿ|҈B�^V�罗l��ׯ�8�I�����QZ����m6��-��Br���s�t�F�C�1�G�Dי�1�U(-��\3G7��ǜ��AK��7&��z,u���Z��S�Y��},�����v)�q�ĝu����hi�tڜ2Aަ�L�rj��Y�n��t$*�Ty���ϭ]��i�[��J��2[�^]dm�ð�R$/FJE�����
yÖ��v�b��=DQ���:qnH�D>�`��bw����5l�/dNz:=i}����m��ND�Zb	���<*�t��$K[�i5(��	�> |C���F��h��,~1�yee֪`�L�1���d��u*��F���M��27�+Q;��f�f�9E��I#��_oea�Zapt&㫄�iL�"�_�(|�X��%����J�R,�w�!T�6���*	�ɟL&)���{ ���}318:Q:)A�y2�6�Wr��l�w�:K��Zܷh�ZU�����Q��T�Vy'QY���X]1�p��si�R=�UR����_x_��C�8No4
ҚusuІp&M�\�P:W]
�[EK֔�ή����r4M�(%���t�ȈTq��r����;�m�ށԓ�jM`�Ȫ4+Z��mۑfI��6�ӊ����t:1����.��s�>�`Ī6�<Y�A��j_�(���h��$�n:F�ag(�u�:5����)Q�^%�A[[lm;���8t�mS$-��~��`jmm�܇�	ж�B�L�BЙY�
mq��t��Wf��Ĉ���|b\g�!���љ�q}��5H�W��?쳨�zؚ��'$8ed��ec��ڪ��_p��t�c��8Q�J�͍-U��ne> H��\�������D�ܼ~��<z��	��	oMay�,������i�TWS���-�Ҡ��@�?O �?�o���K��u��$�G�l�{`��A\A,�p��#�$J~2N�Ĺ	�[��"WI���!�/F�-��o�/�9�`�ш\�sg������0\�=|AY�Sy8�-��B�bÉ'�Lo�	8商�3��f'kB�V�v��qp���.�1��>�̀�	�U/�Ƀ�nr4�n���B��T���$F#����Wj�Q�ig i(]W�6S ��"�����mۻ;�c��9q1��Q�@Lm2����5���1=�*ry!����9�E���WKW!\C�8>��N� �7�&�:GN�:�\�2�d�"s6�<�m��o#F�����,�@EzC���X��
_Vj�	PQ7B$w\V�ֶ�u��Q�Md�bBQh0*Z�K����U�xYI3��o�;���U)� h����Jx�I��g§EA�� �ܕ��Au��h�j�ʜ�zN-m�tK�&���ģA���E�T��c9�&�2G*�L_����v��[p@?�X�����3�u��sm�$i�	��fn"B5)d}4d��.P����� �,=�G���Ї���T!��c��J��?I�fe����^3[̣$'��I}ukK+�Z�7_�kG������q-Ҏp��r��3,����i��lK�i��V���!D�`���܃9K��Ԭ�]��.bk��D�4���ͱ�teB ýc����������
v��t�&M�s��W�L�1�Gs�!�;Hdh���&��o^:MW�����j[=�� ��ʓŋ�1���)+�6�b��"Q1�}���d/�{$��!5�����������C��_�C��z��ڠ�޸C�?<�vvJ���%�<��	:1�Q�v�ӭ����"�AW�2b-3(���?�{�hT�I+XSh��=^Y��C�2yu��=f�"��!��I�	�[b2�F	���$���'E-���gm
k�%����J{�j��Kq�(M�ѓQE/^C{?�~%��%����^,j������(�[�)/�7�����5�#�ɤ�����+��	ʝ�r.���b�R�6	!�s������VV� �>��U�R6�ު^�d�'U���0�15g��������0��"��֜>��7���{4�b+�iL_�N�I��m�</V��b#�k��{OM�s�OU�dq�R/91�)f�q���b	
��Io���z��]T��"͛r?j˝�C򕩧Am��V>�8hJP-Vle�ϓ����v7�.�!��
-�$�?��_���ϦY1����݆�2�����O�N��e�e��N5!i]x�J�Kp��:z�ʝ�� ���N�b�Q�W��PLܵ��t������8Q'Nu.p$�yRO?iT�N�w���-��$���	1�M�%�գ�܈�v��n �d؀rN���}b�JY'2I��������5]d՞�c��o�B~�rR��bYt���^7�q��$�шW�S�坸]�( 0����Ur�{�LN�4ڳ�}u�Oͩ�8ް1/���MP<&���]�c(	�r���y�V|�Lɔ�O�'���ԣ.!�}.J�Ğs��E�F�)���fZ��1�"��-q'h���g4z�D
���͘�ؐq�jr�S�[���TD���Q�n"�L�Ę�(���&�+d�����7�\A}"`��|zh5x4^a.�d�Q����$�T̐�.@�B$�(e��ܴ-9M��}O��ő�mv�X�=�AM �ij2�z�p�Q*���>"�f�O {0y�']q12��_�)	A``�G(#*M@hs��K�sC_��uhr�תX��o��#M� S�9�N�;�r$�c�=h�ۆ�b��s�������y<3�ԕ"��p\M���WW�%���䩯���K����yVk^��&O��M�)s޼�-v�1�K&�5V�'�9�탑m@���vE,�1Uj�"��Q��_�h��mO���=l�o�,4Z҅D�n�'�5q�U#�?�f��� jz@WW�5�^%��CA/�\�Q噸1��!���iux1MJ�{*�F��������5�q谜���r�y�	� !��֊L3��m�][���zG[d�⸂"��3���AY�ت�L�޳����֐��9=ᠷ����/]�l��"UnMQY-�\��Ý��h�۶�@�x���ڜr*�є��#�0A��e�D)(m�Qiv<�5(�ܴ�����!��X��ܳı���l������ż�P.S�ԞNې&����#��e�#(���3'dE�r+zwSt�Fq���<�G����4�#e�Jƥ������1�l!�;dT�a�A�JPM+�֛~�E"@%�~51����4�s�,G�JNf��9%�2.�e"ߓ?s_{���eg�[���Z�q�諶���9!��^+h�;�s����܉ ��J�J6i�n�R���Ĵ��RC4J�(RW
&.)�Aco��[[\��Ot���R��Kq�F�&������.���RcO�7m���{|,�iMk�4�@��3;>�/>�BW���>$vWVG\�V��V{e�ݛ[%�����;�'���M,�z�)����,nߋ��蹲\ �1�-R�/&������A���>V9ggg���ZZė"�7]��|�j�е���ޞ�)t��]�T�t7]��J����{�z�?y"F�6��[����d-��&�|b\?$��s��6.Mʦ�6�uRV G�%�9
S�%-a�<}*�ԯ����V����?����x�]ǈY��m�\��G���1��H�"�/C�_��d�궗M�%9��V�f+���.BB]X�ya�(h����Oऴ�-�<�Ao��
{d��Pjk�&搉O�"��힔��C��"R��E$�z�	���P6���A��Ƙظ%ֺ�;j_�;��Q�õĽ�D)�dAĐ0+�4�G�A'�I& ���kS�����l�AF2WD	J{�PK��R�X�~���n$�5�H���ȶ
&P!��M��N�l �@&���.�@�c}J�KyQ�ve/���T��>oic���/�P[��ZZ'J$�*�n�d�����7�sE�>Fȴ�/�!m��S�Ѡ�6&nާd蔇eJ�t�y��`�n�����K�4���l����ȣ���P�
�Jt?�p�<!��+��f�;|N�/�n#���dz�-l�}WR��,�S+� cF�!癉�"J�A���i.�_<�;����yGd2r�~,�N?J�.����}R*�˸�ox�U�%��?�kf
�3d������ח����\��b��dY(�('�Q�h1y���b�`{�����H�_����qC[>����p:�LGx�Mko_� ��`�����0 Ro'�ۣ�W{��:K��IѸsm�{�mI9q��\�`+�7�D؅��N��8�c9W����X�jj:�'K�8��\�8ս��%������28���EJ!m/spD���N�]9�#�h��B �XR�B�6z ���Tө��]i/\� ���H���Ju�yKQ��Z�>[LU�z��ww��B����܍c���<p�]�~OY�PZ��t^%5դ>Awp����ھ��_#��DQ�(�*%�m���K�i0d��NR���:�6����E�޷=��A��5��$b�d�:�i���Qb�e»�a��Fck���v;���G�,�C���������ߍU��q(K^�zj��ݧlE�l��V�!�X��D���Ŕ�r�%�q��[�>���Aԁu��F���iL�:�J_Kϯ+��e��c�p��o�Y�&kVz~Xٔ~6�{b��9�e�*� ��$F�*��c�ɾL�B��j�Ud�B Mf�P��,�������T s^���gz�";�PW]��ݭF��:wa�&���L+��byz�:��-A�8��4�����fH�3���8E�.���Vּ���.���P���G�Z�-�T�UFun�&�)X��ib\Z����&M0��V��+Qc��zCS��^�Fix�vI���Z�����_� ��cR��p6s�պ�X&P��n;b 6&�0�j�`��ֽ����Y��4LŲuw��G诠���D}O�Y���3=P�<�>�D9�o=;���]�w
�Bɭ�g�a��Ů��|m�^ mT$���M��`���B+$�y�Z��N����8�Ӣ�D���
��+ە���ʲ�cZ-P�Bt�?!�c��~��_�Ri�g�x,C3;}x�|q�v1E4C�D�))]I��]m�w�龜���ճ9x�[r%Dj��+�<%�������g�Q�� �!�\EW bh�)���'�3�0���s�%5�&u��8�X$�3��&��a����ڹ�5B"���!��bL��n��JH��µI�UѼ�
:�@i���IkI�W�]���-�vۇ(/���̺EkT���7EH��E	"�kϭ�%�.�1ݩ&统�.�"��<w�6��dq�J�P�t0R���B��&G&]�PjE�i��uE�U�.q���Ȣ�-U���d�:i���"�)v��"�N���r��R�ۗP�u�~�B%��!^&J�m�D�kϑ*5��AHE4���EۢA+���壮rZS��;ӵ�6�!���X'"*zpY���N�Y]��E
�4RsNZ�@s�%/��V�e��D�금���2XDSa���V,K��4�F�:,�pb�*g�Q�:s�;�����)Rwq���A����hH���X�,�BH��sZ�!�9+͆��Y�:1��EY�#�IP.	f��|u�{��Y��sW�:�F0�h��\�D��"m�l�kkZ����޷���ˊ0�������o�E k+�h�<�o-�Ҥ%�Ɯ�J��DR՚TMEYE����	�r���%E	4����	V(j�F᦬�@)�CR�C�^j�~���r*ְo�͌�+�t��\'�;�V]Y���
 �o���e�?��u��u}��ƞC��SC�ucr�9G�^3�J]S��9ZB�hI�k���+Y��R����	)�b��&���8�*�{�6�)���Z�"�%�d/PZ�z/(UI����}Q�Y��F����%�Rnׄx��0���>�&F�%���#�Zعףxx�o�����4[�������b�k��˜ๅ�Ooݾ<At+�6�yK��Ѓ�ǒt�
£�pND!��pl���#�{�!e�ܒ\�75�c�o�,D�$	���	��	TF�#��T'n���ҾYA]�]�+�<��`�L,$�#�)�S�vXBGy/�d�TlL�̭�1���[�_� ��/��%�
A�*���a��9��SFC.�o� �fxT����)V����M1=�Q{<zR[�5qd"�]�{ac��	�ݶ)�$;�a�|`�fO)�Do���&z���+�E�H#��2��DG���4�3��{ޱ��1O���1��N�5
g�S)�|��Wu5Y/��t����"��Ӟu�aMU�#3�<����J�Y�Ŗ(�m���Z$�KX��u��� ⱞ/���dƩ{"����S-�46�l�����F�X������:K͊��?��Y<h���;;;҇�L�[���x{������L���S&���y��k�R�Z!��ʔ��T��V�'�sKtS����2���  \&3��pauċe����R�5R�<%	=V��a޻5�4���ab\!%�d�
/C,�o)���Y�&���{���tG�B�oy�/���iT���}
.9a��Nis{�|>���j ��ZY�S?�}^��hm[DRz��A;݉�B��iV�,�!�mq��Zx�2�M���
��)�*��M5�55�Wj���b=QE�&x��0������4�p>�f @lQ�Y]� `F�!����i�³:#d�{lܳn��h�$m+��b���˓�i���zKn��=�+ :�v��Xb�GD�"����ln,��(����~X�D�*
D<@%�	Ć���z̍JO�跘�"�V��-a��֬����97�wl����J���O�I�=�x֎ħ}/vs�td5(U�|T�:���7<�x�+Dɟm���#m����<!�C�50�Ѧ���c���\�9 I���r�f�;%q�i���md��p8G��O ($�{������Q{1�)3u�yy��+�Bj|��n*Vs� ��#%�{��8E�+�R��3Z�=�&UC�Q2b����XB�M��wE�2�����C���B�]V꒽���.��,r�ֹңt#U�p�횑%L�ַ�Rb��?g#R�tsW�.%IW��S� ٛ��U#N���ĸ�5�>V�z�,�����5S�¿�an�{=&Q��y�׀����L�E
�6f���0xl
P���IoK;8
B,��a�;�;��F�Κg:Ry�������Y0s���[X��Q��=5��$���Bx�nAY��h����6"������|�O�TS�R)g i�歕$�;���g�g��A�:	!�-RMz�-L�'k�d�P�;��n�[ y������eg��碞��a��(�#[��3���z�[���(�	����\�*�S�����M�[`V1�*����*X		 �G%)���ZiU�BV"j^�%3����� ���'dc~�+v��s*�1�PT��S�򹕻^z�%Y@ ,�ޕ+��q�[u�M���^����MiZ����Қ;d���5��7&I�/�~�9dSڧ�X�t��Y�hQ�իW����Ф��}$s��ڂKW��u�����MV0��4�	⎑|0�!E��Z8�a��w�ޕ4"��]�C���D�lܹsG~o1DwX_�ښ�\���W��&_#ZL��]�4 �9::1A	�(1ܓ����F�ͭmz�[w�.�{M-=M�=�ٱ4��saB��s��*�@~���aR��N#}⚩��8/{ݚ(�i+W��1 L�������roND׉e�Q���r@k�s[�@�i"b��6U&B]W?� @6]T�Y|Q "��WJʹ�XY报�K�*�^��>
����ll1A*1'��Ʒ� �Q�G�>�=��%�LФu,�����Q���fUkO�ʈ��81{E� L��T\�F,���F�>_��{c�j�U���I�j��i7��s-u�P#hJ��,�b��"ؒ�V!�䁻l�W�#,Y�!ؖ|��(]IZ��w/�5Opt��M�6��1s��:H��^R�
#�%�l���摹��X.�[TH*�\ �����1��R�s'nח9��Mqz��
�>c��fE��FY�<���p,.�i�X�"g�;�3�I�\���!'��1G&����V���/�W�V�x�NV����N���w��ڜl��==~�>�ͯy�3M��:F�K�O��t�S��(絖�����,x���ɜ���d��_�|X F��@����da�?k=Ax�hj���c:>�j|��ĸ�(ocD�-ɝګn�y�JTs�`%�8��j4������Л��Z��1�������1x��!ȍ[�Y�n�/~��4�oK62���]J��cB�nW]������{�����a��J�`����E'h�ՙ�C�Ûm�^��sV�s�� ~��[.̭lM]�~����gƧ@�L�rH+���R���2M�r�)s�w^�~�?��?�#^4=/�/ܠ�����+���GW@,Z+����M:9:�V��MD�>����;�ߝ���P[�6���ɢK����7����Dod�� Ip'�}II�v��v[���7o�O�f��{��ݞv˶lY�d�I��I�b%P��]""U@r���� ��2##���~Ϣ�h�9ي59��e�g�&��wb�u�Qh�� �Zq�J
xN+"� �1��8��*��H!�%�D��r�R���>z�d��NS/\8��|2�+���������hp�0��E���/ƹO>�r�z�(��������	���ŋ�����a�eL�*�r#��Y��hPٖaG��0�G��֓���~�7kqq�&L����y�]g��.-�M���{ڤ�rUY.�߯�����z��h�ĆjF�S�4?����0��!���>�jr�x�9��8Lw�_�^�PB /��������҆Ԭ�����s	WS(W  ���9Ym1���5,��~&��FP��C�XpJ"��nq�uZ��Y��i6��o��>��'���'z��NVi���L�|�p������&?qs�`N3�;���E�����γ��ѣI��=�	�s�h~i�f�<���E#� \`��B��OQ/��@��^�B��B���dA"��%���Erњ�},��)-�j�0Ƹ�����2�=CI�J��.�@���.��G�%X�R�2��3'���>+]��6�������瞣�c��ڻv�'�S^~\����g�j)k榘��x�Q�C��a�#884��93;�N��J,��%�xtW�F�4a4�Nk�����N�k#�V�i�Տ6뎚�+�5����O��?��{A�����4�x��d�����w��{��?��v��M=�=�e�ڵ����^�}Ė��{��1�Ŷ�*=�ߙ���܀i��C}�Ƨ�-f�d5�U�������N�+�����#_��e�a���(y�k��\yWD_�+�����-��cw���AÚ�f�"Z���������n�"%l�B3$Y����1{XR�#Ti�}�jt��Y�M����g��ChFj�� ��8��$���I�F����`�B������]|�dyd
��Œr�uf�o햆a��y���(�3̼�\������O?��'�rI�GDu������B85&V�U�/+�3�W�
U�5I��/i��( �T+�����] �\A��ikg���K�M.)�pD��˨���U��8�\=�q��K�B���Zʢ��*�t|��8!�n�S�ɐ�rj������5�G�����ac��څ���R�$�U�$ɫe�		S�).*P#�4��VT��KF��N�����-kM�eq�)����%ԡʑ�|�D9����QHM�A�€�2m�)�~���8��$<X<��U6��͝��9�F���z���Ӷa�i�'��45H,�|�i0��E-q=���D�D�"0���ՂOl�B�u(	l�|�8�@�
���nG��&�y��;_XwlԦ\��]X��9&�o`��7od��]V��^��'B�C�P�2R-�����Y�L��˚��q���B�j�[d!݈]9�KW�*,���Oa;`E�ޱ_L��
�^5>,�֞߀sp�H�g�=�,Jk�W��Р��D-�lzw��!E!WPB5�ؾ�*/��!\�5Y���w�?��U��������X;���&�ѡ�A
�gee�������]�d�X8]��֦�����9���6=-���,���B���ڂ�i:��2��u�1�Z^$�P�,V �"|���G��:�y"�Q�����������Ӭ�"��	nȗE]��خ3G�mt��q�	
#U[V���ұGkBj��vy��#�~�$N�x��q�����Yj���/��E%oW�!ֽ��H���H+�iLt�N̳h���
!����3�E��G6ӆ�P,���i�I�j9�8��~p|E&  m����]!CG��[���m���8�p�L�4�����Or� G�����Z�
i�j4�!�hx�Ɉ���$l]'��/���0�԰k�ڻ��j1�a4��`��|_P2���`Hh6&�9�ɒ���R�7�˒��A~�:ߞ+LW�t.���1s������� fI�c���YB1�_v��{���Ώn$9 �%Ӣ�ܮi� �i{ؽ핶��HY���
et�I��dD�N�q�A�qن��'-���@S�"�K�yM�͛EU��������0���+-N|/sI����53i]���]�"����j��b
��*�lLV~��2	�ARu%��b)�Ȭ�è���d�Zk�l���5/GB��!9d���� Qo��BhC:��}k���EӞ�P��EDa�A8=hQ�_��)g0f�� E=!�ܹ ��=C\A��<�N	��"]�+���T$%��(�`o������(����_�e��9m\Vj�5��z$N�,F|�>��<,�E�����6��K�,ءiY j/��ժ9���KJ��;uXgg����B`���ϑ����'&fH���3���փd��tw{��K/yN��]@۲$k>�R݊�"Cl���%����?�Y�q��.�#`Ω��+������!�w�f��Y�wU5�,�/qQ��������^��,���B��̕�/Š�=t@�3�n +���\5?�S�r+�^B.S��ly�ZU��D�U���D�
�v���$���p��k��$Ysj��SE��;:�������	���H���&
&����m�S?a.���$�W��}��zS��� ���c.��Z�ȝ�,���l�l��/�\7l��dA���)��#�����9�\���o��cϖn��])��:p��������(H�	:�e��?s���\K�k����Τdu������K1{Q_v�ݿ�rB�����*#�t��%:x� ����)�UKi~`�n2�|Q��{N�i���`�+yv���h�)ԙU�'�&���\��W�<?>������Ú�/_��cw����49��f��x�qP�Z�+�*���db��.]po3z���t��޸Q!a��C[u;�<���S�������JKʮl!�$��Ƭ,Z����wY�v�b̦����J5�in/Nu��տ�_H�ur��T;�%�h���XN�*4���dOE1`$k|����^zd��*�֘7�Ѹ��P��|��ͱ�n�ɯ�W���,g�QL9�4Ѣ����WWo7o�+�H�Ǭ�D'�p�`l4-���*�kK:h�G׆��]Ix6rǥ��f�ן\$�?�u~�x���]d�[t��(
=���J��	2d-j/1�X�����^�(?Xb�7:�+��j`�l`SaK'�ͺ<�QLY��v��+�OE�߅��z�����n2/hz���2������$ѕ�L�k�(q>�]�vK�%y�V.V�u���kl,��&W���PC�!*_W�Dj���LU���0�|4�1���>�)*	Ts��$Kp��1Y֜�H@�&+��� �W��9��06;�,��#��C��mvx�"�'��Uo)T5Δ��˘�r���H�ʣin�~�ˬmKKO��=t)�-���]��2���B��=iЬ�]�s�$8�R�^J��a�a�(k<�v��]o�.����-_ n.{&�Jz3 Y���A
�&�����6�mYS��꽆I���<�d1�E%�BR[4�I����j2�Obc�Ʈ��IJ�?���Ү]�X�=,��϶{�µw��c��u�6�;>�������lָ�#y��)��	�L?����6=�xě6�7�x�����Iڰq�3.a6`)v��M[�l!k8��X�eE2� &ߛ�%�#�q�u�Q[�	6� gϞ�������jt;#�>u���۷o��~�;��������� ձ����>�cǎѩӧ衷�~�o��_z�/�z���xG��/~Ovz���T �‒��>��#��p�GE���g����g��K/�Gę������'�ҙ^�-#[�f�<�M{P��Y]ج�z��V��+t��Y�=-hh�v���IZn�pj0��,Mqq�N348D?��9���͛��G�������#���i�t=�8額6Ѿ�=t��k��χ|@�=ݴo�(gȿ�⋌�s���i��Z���U�|��YY?�b�JI�P.6SEYs����֘��-�z����?�W_{�����wߥ����F6aFK ��Ѣ�g���@���ԃ�T������s��;H��G'���_
r�2��v����C~�o�E�ԁXv�����=t�0�4n{�u�[��w��o��QƟ���̿%��ѧ�|�.��J�ڱ�)Nm�f7gERUQJ�4��ϕv�b�az������5�I��/~֡!ř����/��N,�چ��t$�S����S�Am�����͡�Ǐ'=O�J�7o�}��ѹs�h˶m�9�
vp��	�_�����s���m��U"{���
2
�
�s��K7T�r�l�yA[�B���2e������C� �����v��S�"m����NP�8�ȭ����०UIEp�����)�}��y���L;��e~NOO���,uuwyj�OW�\�l'-h�z{�����H��z��,F.n0�j	m����{о�@짻��2x 6]w�TQU(�I�yA�Ø���^REU�I�sne��`���Oa�
U.Ɯ���m^{2�N$�=s�$���w���@� ��{���'�-��4�*P�����m.|E{=uإ� �E���K]��/�uw����ίpם�y�ꏟ7n�'O�<ݻ{�nݺɔ���ghӦ��y��1ݢd�$��cF�p�Y�E=G,8���� dǃ���K���{��q�}�՗4t�_�#/�!c�絓K�.z��)匌lf�ו��8��٪����6JFS3~_+�9�3�3�5���C۽B�8�Ů=�,KX�+�"yEa�<k�����_�~�~��_��A�bR������;hl�6k-7o����!���OyF���-����s��~̀16Iy�\-#]#�rQfE���Ā�)ܭ� M�5�s!>���A{��e�%�!��KS���q�T'Gs�,{4��Яi)�P�
!Z$����6od����:~��xj �m�Zǩӧ���mT���~ސ&_��?����S 	��OU]�8��!Y��w�f)�lĵS�"�q�JTE�D�V��e��e�P��j �%���H��\���0�km� 
}�����-QĬ�JS"(v�\k2�n��d�r�_�4���(B9uF7�ȃ��@�+�!|�"/����2�'�h�p/�2@#[T�ꈦ�;{�e4Z�~!.�S��Z-</�����O��;f���7m����f�lg�j5�6I�_|����C��� �d��h)�y�;yW�M�����s�L�ݝZ2�$'�&��@�����U�K�s��J��8�T/q�0�)ҋ*���Z�\�H䚈�~��>4ˆ!�h��x��}.\���7䰷��r��?��&;D&@�|9��T�&�!�>$�E�a]�+�����/�c��v��;�Ax�F����qn��jav������0���[YX�����*�nݾ}����;\o���G���c~��U�(r���o:e5���$
M!����C^N";���lsMM]c2�5�RƵX�XWGIVEEC�)bgψu�k����I����N����4���<ݹ3Fw����~@;�����"�7�o�|���Af;_�݆ɇ���E����	��_���ݹK;��.�/�{^u��^�4z̅b{�A,�t$�w�����F�O�*�qȽ.oc8x����7K�$o���H	/fњ���"kjŬ�,pӌ���P�E�������5�|���S";�ɠ��?�ȿ>d���>���:w��x����k^Ki�w��)������ϝ=�Nǟ��=���df�~��3o�@��<2���������`LQ��c�'�ې���͛7Fcr�c���u1�B���"���ƍ�&��V��@��BhW��qFY�[���gS�7~�3j����;���K��ֵt�����~��nڲ��4��s��z���)���7o��m������B�0��/�B7�^��[�r��4$g[��u_�n�$�М m�BH뾧�`�����h��^�L������7�]����Jp��I���)L�d2J�����%l��o���xgw=E��Ӧ��ğ9y���Qֆ]�k�N�qld\D˿��2����ǏӡÇ�>��~�6n���wn�	
|(/?Qd���QCq�DƂ�ͧ������6C;	�`���cw�!�X3O�9Wmd�f&2k�!�/[zMC��%��su�@8�u�W[^�.����e�\�]/�g�|8A���
�\Ԃ}`]�7o�Bol{C<�^�?��~H6�t����ܽ^�E���I6L��{8��i(�F�jO�ր�ooϨ>L�p��f�\��QTl�|���B���ڮ klJ�?a��4�~fz�o
`�U踷��n����[�Վ��IZ����z�5�9W+��/9v���&�"�&*��V�Lu��Zxc� �y5qK|嵭+^�9z��ܿwOZ�utg��"J��*$����>���P+�4k�k84�T�SX���}�)�.��X	���������m0��X�1WC65i�����'�����"�,MXH�<$YC���-�W_�~�h�6S�����T�nV�2T�{Z�X�o�x���2&*���2�g8=�?�\��������޽k��%M#�K&[9���0�̇��5��q@	�t>˂�[OK���v����o��4=�����o��6!�Vh�Z�l�k#4���~�nr"	���G�a��\c"��R�+�6��I/�^�Nz� ��#P���*�u����1�'tP˭Qvg��i�JA�<�%8q>p�Uo�/�F�&q�"q�5��������O~��Ң��z]}�&B�N� ��<<4��ŉ{B�?�e��W_sh�TjWݠ�%uG����ʵ���o�����O����],V�v�`�uh�mރ5-�.Dp��Q%G�/Ӥ����o�O
jA&�
8��ޞ��D�~���f��_�e�������}�����u��2�A|��ȞG�yr�̗vHi{�d��)��ڗ��:��4k`�C{Z!�ր����K��gg=�Eܦ��ݻK�w��_@�Z������Qa�[�N�Zq☳�q�� H��Y��+WYӲ�+�
�:�8ǎ����}v��������χ��*c�ט�&�[�eg_�ܢ�/0�D�zZM"����)΃%�����w�~1ޜ;��\�B05����;�,�1L�ƍ�L�'���M�݊��J�%�{�Ȥ�	����9�-�L���|_$��ݣ�鋳�Ӆ�.��M#t��!Am����[��{2�����=}��m���9�?:J�����D�B���	�Sݾ��裿|@����y��W5�����m�m^��0�3�\�����\�o�h���JR]D;{�m�@37�Г�'M��^e{�W>�}�$c@^�����NÛ�Y;4ӣ�rע,:���xt�Y|�K5u�J��!�g�}ڳ�?��O��u�[�p�M{=��o�a��^�}��1:��__�|�;)��?�OI!�|��/��2�9s��{���w�66>μ�it���%S���k���V�~C�O.��R�X�X��}�嗂ܱ�ܡA]���9��j�� �iO�&�ݪjoPI�Xi�q�ׂk��@����cGyr���8�Y��{{z����{�( �0�� 0�H�54���2�P�� ���2{C(��_�/�en�%����]l�Fc�QЗj�����a��Q)Q�ӊ���#_��gZY�Z߂��mᨸ�%-&�D����sž8��3�h���t��ֹ�9�%C�<o�ĚϲjC�>����Ň����O�c{yY���f� v�����kfZ(J�Q�dq���i�J� '�bea�fc�Z	�Z�Â$�kշ�����m�
��(A@G���B=�)�:Ǣ	@+N�y���� ��]�K������bæZ���7�J����!�;&vg!Ӿ���e�0���������D�,(XW΅g��=R�c��*�̓�N|V��~Nm���%Y�/��.�99ět�7\�32yw�k:�8����dJ�cc�MH��N
�@��P��g����T��Ɓ_i�[����jKag��J��H7��hra���3�k�>��m'Mb(/��,���^Z���eE�gŞ�U��G&�M7�J�X�K9W�Z,�-�ھT㴧9\lBw¢j�~Vxr]�|��J.)������);)��3��+ �K��)�8��'�^c����#���;c��M�D �ˎgAG�-}2-��Y'F�a��ԭ��֦��Ԗz�6&v������m�����HpU�A�,�u�����=^�d���y��"��=ӡ�}��@+M�Ak����H��a�p�>�%�Op ����[t���R棰�*�o��oi~n�)�c�s������eUAyxN�x�y�������Bej���.f]0�bᚻNTe���`����ʍVt��Q*�в����~�������B����^�j*$(C@~��g��1v/�cX�09r�8����|��e��Oz�	/��\�,���C����F:w�K?�3�Oڹ����u!s^@���Ů\��.�_�����ի��}���?�|9�ة'Sls�ٯ^��ss��-ڻ{/U�# ZЪ�b�8KkYgn�`���QXNo�l��e���jb�E:0�@��XE& ��������1��[�h�Ν422�I�G���v4���/x[����L�X���N1�!�*�%:XfU����\��E�hHSy��6��-[����,C^z�ea��`Ŀ��ijz���'G����dq��)Oy78�6�1@��%�'��5���jY�@QW6�IL>c��9��������l�tQEz��w����Z�|��n�'����E��.��o���2x�_ë��4�{��5Us]p���$�0��ǎq�-v�qOa����IW���#���~�o�����~���M����7������l�\�|��8@��s	�����~�c<e�L��"/+�F���'��`O�Zx��YKi���{Y�<�Z�~r�߱�qx��򀅸�')���&W0vɵ�$��W�6u=u�BA�H����Պ
�LUk��*�=�R^=��/�SX)�9r�nx*x����a�ݼy��ul4���:��i���rd]����P[��XU����,�J䩋ř�C�%�u2�P5.�����-[�2+飮B��EvgC�ƮDY\���[��١R		��{��7LMX��?��'�Y�XU���b[`,H��OP�YƑ_ⱌ���q�U�s!�po$�W�������\�%a�R��fk 3��j��� M sa���(��t�P��70�g�y��>�<����ܫ�+//�x���y�+��������� ��];w��/β|8v�hJN:�U�J�5�����Ԧ-Q���"3�Z/_���d����:�j������6m����g?�g�z��������,�0�S4����p��֭�ͫeB����K��u�Y1z�����Jc-����CL��<߇�?7;�ٍ��|oݶ5� "lZ�d�?�݌�2�;��< 7Ck��y<<.H��I��7�������_�С�L-X����Zӧ�}��xP2����� \�$��Rn�c{~�b�=£܃��SQT�� ��;����0?oV�.p+h#��u��	��燠 I���B-b��j�Z�+8%��\�f��VW%�\xhnu���g�xr&yd���߈���Ѕ+"+.Ĳ��H�~��Ƶ�t��>.��>w�4��w�`���=}��� �x3撤�wߨW��cd4K[�GGf#Bi�Jj6L@�A_Y v*�X�]r؋I�������3�p�pO�0q��?Y��Y�p���=qf���"����i��!���k�\j�Sɪ�?���e)��#[6o0���X�ͣ��&��G��"I�J���o� 	itV��T���X����Tė���֖kI���,[w�s��o���i.q���ơTP��-����iE'3h�cnS��?��U�}��^ظꇫ(�^OjOk
!s���W掗�@%K������.����!��#
�sp�(C5o���ũ)~��͒m#-ԅ�]iޗ!q�S3L~��#3x)����s��.��cv�4�������Vm%ѩi��5�u��G�]w�LY\0��-![R�q!�~Nn����hKH�a&;;��6xȐND��\��/=_2����`K-�Poi\���"�o�lJ��;�
�����!��T����6N�F~i�v�J��e^m�\o�]a�"�O���񺍎"쨕.}�'\�3D���ua��B[���7k��B~��R��^���n�V2����7X�
{a!>����ߥ�Ϟf�B�·��sg�l2�3$���[L�K-

���N7�����!�/��3�;C?�Ꮘ��d�MC&
V`ݢ49�V��4@`f7�b�_��hc��Sc����.�&¬��Os�|�����{���\QhEo���(���%�r�@�-�oE�m�Y.=zC�K'���s��L��8���\�;t�Bb{	`�Nٞ���T�$eR&K
��As�d�����cm���N˟��U�z�Cf<]~�5���%r�%Ub��5	�����������G�A����j�4�\Zf���pI�u���v��o�ݻ}�ݟ`�ڱ�S�����?�E�8::Jސ��W�3|�W3H�޼�a��uղ'&�֭[��I������1���t#��ꭄ92�fV�+�.\�C�}�;�BV.�:}R����X�Uo-�Z��[�S���
e*�#��JN~ږq�L?5=C~�O��5��d��f߁����&����nߺ�^���;|�#w�:�|�k�͚^���_~��=̮��µrg|�~����k�����PN�'��Dj*�Nׯ^����M��ũwZ0Id"�j�֩����q*<e;�Я!���xTR��B�.yæ���	����,HB)Ɵ�����@���i���/�,����}�u��r�gtI���Ob�!�g��B�A�5�駟���A
�"T@m��<�T4L|]m�v���Л}�Ν���|L���d��@�1j�&-Ɯ�����nݸI;�m�>��j�3�X&��g���'��S��_ˡg�$w#���A��~�,�*���V0��Wj�7m����B[�|o� R����h��[��՛�X������{@��>�A�L�T�o��o�;<̊e�uT�>$$���; ,]<XT�^�z�:���S���
=r���6蛒QO/|F?��/���ѿ��_���@L�
ˇB��/~�Kz���-}�c����B�(C���ߢ��^��S������t��U�$��i�s� �Ξ[�j�������*�r�S��3�Qg�j���zA̢�E��{xdM�W��PW'u��^�����U[�h�����EޑHzˊ"hQp�c��9�8�E�
o��`��.����&���K������H�<�<7�Tշ��p o�Hp�#�`�ܙ�w�ʹ\���&'����`�9UL����K���S�rÿ/��r��3�G�l��%JG�M����5-Q�`Y�=���v�8F�"=�°�����	7p4o/�␥�H�4�f߾��E}-����cw蓏?�O<{X
b��m�z�}�9)�l	^^8-9�N�kז�WS�1\�Y��I���6�,\��XOEdb�S�����*���Y��@gY�F����Y��2JJG��7r�w��Ӳk>�.#߰����/�ݝ���Ǟ�_�"~�
fP����?O��ߡU�������/=��^S��إ�g�(OҩS'�_�.,�sq��=p�*	��z�]�tQUu�c
@k�E���HN�g�7~�����G�ywpXMQ�%!3G��~����"�������H*�$�%�/�R�Iq^��� ��A��S}-3�
2g�q��	MH�������5U:zh��CԷuͣ�tq��<�k��%\���.�����z�嗘� U��4?���h����-���z������=���rΟ����2������6 ��ǎr��G���<(��S��� ?���Ƚʾ��~���� k������K��8%ɿ9���Ȗ��������]{uM�t��I�_QC4�׈�$.vB/�P.`vպ����4t��q����A}��	Id �������
=w�Y��<��~z��W��z��	pW�v` I�Ѽ�o�៨��L��Y��i�&����W���#�T\��;�C�G�'v�������=�M�F����RZl&��>*�7�6
j06ѕ���O��Sߙ�0��в��4�Ή1�7�PJ��P�R�r�7��4"~rQ�Ɯ���,���jh���~�#���Ѯ�հ�2�LLK�����fc��4l���$�B�J XK���F�"Sj��M���
rF��Y�xR׍�s�Aj���L�U�^�rx��Aj�d=(��8﷢����:5�k��X��U���J��x7IN��LPwc1kd��������,ߦEv�\�|p"����ŉIFB��	^i7C.E+��(��ؕ��m��}���Y�3ۊ�i�~��M�Fq%����C͚��S�IŸ�>����s�Ʉ��?��st�����vhoCk {&�1q��Z����LYD�P�g�Peն��av�
f/&~��Xk'Rg��ou��m,KW��d�\b�:x�T�H�*��/�%k-�Ү�B�I��hWJ�y͢�y؍�-/�UL	�nᕭ�T[\��$��J����J���������-�^�s���nb���p���)�-H�eDC�2~KJp
t�>fl�+Xۼp��mK��4�����$�w���d�b�\"K����8N�{6���|��K�����,�SG��d��t���"L���X��x��g0y���@:�� �d-
H�J���c\� �VFꊕ�ڬ��X��wJ��5��&�T��hbG� �L����vgdg����8Ν�\&)'jJ���!�y)m�?�n��
�ڜE[!��
�p�N]�1���~���K>c���T�N��K	k2�UT�-8�J��3�c�Cy"�&!}ؒ�6�B(��D0/n0�E��6�c����łv��.m<q���j� 4��i�X�9�R~/�U?��]��(��0D�-ZB�󳼀�S�8L��XM^�
��@[1�#��ΉI�J�(�"&�5�dQ"��S�UJs�Z���pD�V����N�<����T�&#�6�?�� U6v�j�͡5Hj��U=���_w��eq;��69��n�!Ι�!�9�/-d-/5:q�&b�����i	�ik$�f)߇i&����-���Q���4%�s�5^[;��n���p�G
G���f u�wv�S>��o���D�j"�]��
yHI�bE'4��&�M��6�AbM%,Q>����"�h`�i�Ѫ�P^B��e�Qɂ�A~~�JI��lٜب�xp��W9#�3���>���a��m���|�h���!��QC2�U�f�:Z�T:Q�#����N�+6Pr]�9
��c�\uf,'l�ɭZ�E'7��79�r�!�^*��"��Z�E�L�#e�_��s�]��i��u R�9-%g�\v�]�&��cEk�(��-K#+̹TV`�$N�5Y&6
:�ӝ�j��A�6^���Pm�B�,��,AR]��4[YJM+X�y(h�+�A�CN��(˛D/��I<�haSu����*�� ��N�1;�?�$����S:����?_��=Vequ?�r�-�������7s�u��49��z��u�s�V��b�����3늇���e�Y�:xJ�b�ֆX��Ɣ��!R}�X� �ǵr�B�f��ԛ�jz��9�V��|���Lf�f������i�j�ֶ �
ʋ�� B���n2��XŦ�ӭ`%��~�#RwQ�d���]����N�J���QH+m$0(U�[/ɷ�ڮI�i�vO�-�n�Q�N����N��o4�i�M�"��(�ޕ�����|�W!�u/Hr{�Iȴ̝�p���5R?��Q�JVA�%����&P���<��E8/�;�N.�k�!h�в΍�rsԭ8c� ����.R˛̈ҿ�m��Vy(�L�HR�0��N���Uۺ���Ӣ�3���m0L쯡`����.��U��Hɔgf�����gŘ�$L�_�h�cZ���)9���\�c�-�L���x�־�p��n�Őƕ��RP(iH��?Z��E�z"ף~��)	�u�S��E^�a(���ҪΝ�Q���SIv�Y���ť&�i4��5����}���b�4n�Fw*ݧɇk�A�j)�$!s.��E�����{�v΋b�S�����6��'�S�j|����
'l:q�( ّ��:������X��^Du��~�zv�ד#��G��[��RN*�wd��X�b�	�[� E�w\݂�m���G�R�JY��,K�	V��cmϾv�b:c �.Q&Δ���jr��-�-Fa;���,���6�����LTέ�06nC\�VC<2�<*7�΃�a����"� �$�[ӚG<��[4�5 [ˊ���3kç�W���a3k��*�̓<z�8��
��07{L��!�lĆE)�Ar;G!摖mފ)&�}'�"��&�Uȧ�;��o�om��k�Fa�?�R'���wc�D؊B=%I`��=3K@�$6���^��yHI��ՙ��@͵�tK���z�jV��b�N��m�ූ��a��zHD���ʣ�3Q������	��dP�yv�T�M?���%�G�0������6����QL�0�Z8��1�{���o�T?[�+w]��:��*�*\P]K*��WX�A���>#}HvZ����H�K�\�JklsI�Q��.�o]���k��x��,�~n�d���@:�M&��D	s��V�)8U�<PQ�e��Y�(�R�M�$jY���꾓F�5��ߦ�d���Z��R=Q��5�A�$��.\0�
�d��Z������eH²���Vy�i��X���u�0f+zMM�I�Ǻ����`�T��A�֔x��Y��(k��x�6��vG(���F�F-���E���:� ��Ag�0����uj
]��p����{�ɑ��ٙ!�S�2'�E0�jR��yh��'��P��� m>�oc�A���G�;�2��	�F���BYLN��B穠�T=8��{r�1ת�C�3v�6n`�ށ~�R�iWV~P�s��ȵ��ay�gp�����
����ѣ���������--,���0�!���{2��rZ!�%��Ѽ1�z;��cw��2���RP���;O�f�3'?Q�	ۇ�id�F���o��/�BP�=8����8F[�m\���@���%y�-8XQآ���T4q	3Iw`-�P��>� ,�L��g�qy6�pQ��c�.F#b6��Ď%�s.�se��y��ˊqf�E����ׅ�S�����皾��>?Fg�����Ο;��0�pP@��Lp
4�G�(�O���`��K\�qp0�oE��M<x�`�������8��8�h����wfj��͇7n�[�oч�ŏ�,�y����!GA!A%Z���ku�����B�e?���k�-�'O�`W@�h��^:u�U�n����4����`��]�˾�ט|��Y�>�?qo�F�졮�^���v(��%Y1~�7`�1 ՠ{��}t�������mz�]���E�փ*�ȿ�������
�����^y�Uz��3|���F1�z�"��)-����L�
�j��`�ܴ��+���;��Z����j�D��̝j��W����s����� 
��e��0�(������Dn��� @�uPpO Fp��%����Mbj�'�ט�l2`v�D{p�����������&���������0t�%F�
w�i�t�g�[Q���!��-J$��N�\�wa~���߸q��Z�q�� ]�t��:�u��Kw�*m![��S��%A�����ڕ��������366�]FF6�=���넙�.�ĵ�1�r
��_`�@":�Y�_�{������@�&�����vڳ/�z9��Ǟ������&@یL7X�&a���k]�NT��e^�)�.?=�`�߾9Ʋ%\�`��6�lt<,XX��rg|�*�H���橢�Q<���#�<Tp���G�R]o�׏<�I��勗����ڶbq�?{����w u���ԓiOM���+�(�Yi���VN�~y��<���G�n-�"��f��;�;.���р�azy���)@] Z����kO���b���w�.����l�����=����ԦM���_�����^}�5������k��n���&�˵"ԁ�R7�r�f�ܼz�j5�������t��uuv0�D�l��NVB�3�aPo�U).���5�-�4��H;���E����M~A:�����3?�w��aO��X����Ȓ�L��e����釬�c��
���]�L{FGQ�����y��b�H�z�c���k���o�}M>~�؈��?�b����Nf3����?��^=�����P�^D�1k�~" "P��M[���$w��|��l���v���Dz�t��]��1^��J��G,����_P��L0����q��Ӕ�O�0��m����1��&�6��c�:���7 =5�� 	(�%O���'H�	��	#��4<<����~�@��[��-?�c��0�	�Z''����]��;ζ�*{�rS�f�8��PVg�Mi��<P&�T�]�
H��6(��@�h��T[��kv�W�o���|�kzݬ���@ol<�Yjж����\�ԹjUe�kV{)a|d�Z�7��A�zp�>?Z=<��3�|��6"��a�`��?:F	�����pL����
|�-g(�^x�;�|��Ǭ	�����]%�s��d7�W�=�A��=�F)�+T�./�&�-Pk�@�X�-R��@-�� π�����=sP-�aSU�sA+쁁K�s�S$y��4��"�Ф8u����@q'�e����	�=L��ݧ��ׇ|�Ͳ�ْ��Y�2�;v f�8h�h�=�Gِ<r���h�� m�8���M������~����;6�Xo5}�f�P(Paq&���DP�{=�V4:<(�{ Rl
 ��.��+X����lP�q>�V�A]��|zb"�U�d�xYE���ĝ6���C>�V���\h3
����؁`Uv-C VD�c��Y��O�����v@���2�d��I1������"yM��c�>�S�������A����^�*i���r��>4f1D����î�:���񋰸$(v�G�~���:�Y�t彁��Ѝn%_�T���(��Tݵ��"��XV��;���� ����>�1�r`M�(( �����۹Q�]�K�^!�x�O�4�ۿ�SI?��_��R5���P|�]�3�D�e�P!���V�O_��Nx�㚗a�<�lP�����gՊ`+�5==���]��ĳ�<�I7Ri��EhNi=Z�ֺ fQ��a��7���� ����nO�PC��i«���Җ��x�w{{j��~.�$	�� ��N�����'���7fh��m��~��_ѠW�a|�c��-5��Z����\����-���<��Ը��S�T`�� ���Xx�:�?�����<c���,�7&�]� �Y�.��'����yԒXV�*[&��YGN��9 �xk�r�˒[^f ��ĉ��fp���2U�6q���|+~������2o�^,��̔�����=��۳a�qv%^��߽O�K;��|�G[��G�i�N�n��d�	���`M�~�OO1�&y��~U]=]�-����C�5�� c�A	/pM�pekW�_���]���Y���-8���,��G6Ӹ��!@/_�L�~��ݿ�w6�U�mصೋ�{��	���E�����gOpU<Y���c�,,+���$��ħ�4�
8�v�
�5y�������mݶ��}�9��[o�W���$��q���`
�Z� �w���=˪7Tn�%�>/�7P<(���;�Y�	\��4��/Hr�Y��]'�c��]�ʞ�s���o���;�-����������� Gh�[��<���I�Ȃu`��)pG�nc �$��\@W!�ѣ���]N��׹G=���W����^mF����?p�
��/��u�=���_ee�7F!�aM��A)��J:�`�q/��*#I�k.EMjY5�+Q�"�P4�Kj��L�����t��s~'-x���wӹϿ�ݽ}��t���bڳ`��z!��'�p?C�1�l���l������.ܺc'��K^մM�Ij�
�
Kl��_�p�S�j��]��9ׯ]g,�-ޮ������}�?4�<��M0�	o'!�������HP,Ӫp���������o­��x��:����s���{dh�0�>��)|Z���:��Y�?F�lea���N��72����(��a)wV=O�Aj��-�p��Q�4��:=B�\7�<dA�&YfHW
�y~��ȃ\:x�}��gt���^��o�ځ��T]�,���K�8/�����l�"�^˗��~Q�zJC_Gg;�[�����
n�6�(N��Q��W-����=���P&�i�8�'r`�l����vE��y�0_~�p�#�_e�����$�g�-�*�8�����7� �{�b�l��w쐟�N/s��\�c�!R�l\�vY���1A����%/&i�ˈ{���}=������t�S�j����s�<���	�q���E_���h ��!��c��%A|w;$9bh���;�n���$��^/KF��g �ە6�� mdiq�n>��w��# �؞�<xP��A������mF�_�C?�w��t�b�
0�XVX'�p)��0I�5`�m�~����r�+p������/�8�x�G��ܾq�Qc�ܴ����m���]@�|8,w����]A5䚸�\��,��Jg7�T���ϣ��=48LK;���=4�_����lᇎ'A?��^�#�)^V�^?q���EU����lgW~V���FX��q���2�������wqם� ��Q�M]Q�k�S^�aQ�a���J��{������D�������v��v��F�����(�)@b����F�	i:U�mY�/���'���1;	��@לo�!e�=v��GxbA5�=<9�Q!ɡTj��莃�����������Dlĸ8"C:x�繟�<���f�,в��sO�3lz*,�G�Zˢ�� ��]��Ӂb���U^���9x��u�W
��ɚ
vRV��Ѕ�n�̶$UfI])Y�,
"s�^G���v��_��2n���5������O�"��� b�Da\6V�h���eԓ�*,-��"򤽍툁���� `Q����q����lȘV� ���n��<ec�శ�a�J�[�XP�&u��hL�36p|���<,���p,DGO�'�o�O�"�5�z�����|��-SW�6��YE՞�p������~��� Vѝ��װ��ׁ��
kX^`s#��Bv`*P�=�m���H$��pl�ވ�rd8�K��2l
�)lBll�Я�iQ�J~��,˚��*�H�I�CfY|���#�U��݈��8ǲd�YV�^P�1���B�eg��?Ь��< ۰���O���=b�Mh`pC��������kI����d>�����,\����͔֡��l��e�мi�~�XR��dʚ.N�����0œ5�_E�z�/k-��������݊ICpd��Y�v5������q�*ٔ�9I�����nP���|�-�� o83��Axs�OP&��-/זⰡ��	P���PSbzy�:�K���뚼�c]��M��i}q��� �=l\���~��rA��q��Y����Ⱡ�P�Q���D����2�1���&+�L�
c�DP��m{L8�rq��j�!��(�+����v9/ת+Z�̨?V�:!�ׅp�m�"�]�Z�f��m�vpÀ~�L)�5M279_5�J�[	!����������#Ƌm�-W>��%k�W�,�Q��0b=��Dw��0LA�KXJ��ĸ�����7W��W��2mՑi�bE�^�T��-��Z�|\
�N7h.��p�O.:>'2kƣ��%d��������E�C�j��/T���̩��T(���1�X�Κf�;�<��ܢ�U����ֺ�mw��$)�+�����$'*0n�&@ƕ�_^R| �j�j*E���\�����x��4�F/�-'�&I�9�Xw��O��)�.�
QQ�_&�/�����5���Թ�Lz�c�a�&k�\�+�[Q� |ε�E}�:*ժm<!	��4}�T6��F)u������&�����ygU���b��z����� oI�]��۠�O���X�B��.nv�h_�]��8�����}:OZ��le#b����Ws_�''k�b��8~p���LvgK˜��b�`���$m-����NŅ�pB'9ˬ�(����9DVp(�@�I�m��k_}x��P�$�\S���E0�¨��Bh1�]�U�����QќZI-J������h���L6�ǯ㢁��E�Mg��f(,���r-%K7�z�<S^G'���ː�e]��%g�"<�xeY��b��]m��f��.t����Ƈ�Q.G���(�^��Rt+nDE!��48cG������!έ�i�u\s�h��nWp�xM�EP�;'��$�=��'$$���g��.hN�y��E�4�"�4�����J�i`�� &F@iva��+��b�3����u�����#�2X�jG�3�Tcrs�Hh/�0t�UQ����H�Zc�\�QG=��Aǜz}��$J��	�t|�2i�lx��H5Q�4m���Wctk���`�|U._�
���l��YW���(\�w�Q��;�(o�X�hlL������A�(y0xX�߫o���X��5ːT�;�/g�{v�d7���6�0�n
�奧�y[Qe����$�i�P���O>x|cJ�-J�Qk��cu;D5���-���m��\,�@��|e�Ч�,��G����0j�V�\I>[�����6�� �˵ؙ�H�3�g6f�<�R�Q�/KǓ�A���b��μ,�Er��)�5��T��֠jy�̡�r�� �N+i-��< 6��l�D#K�Z�%���9+�W�J%K�S�bzݕ*oLf�y�R_]V�.��WP��2>�^�,��xHq;Pj&�y����`Y%:��+4/�+NH�����2�D�����'m瞋~*#-+3��e�6�E��RO�:$��x���Z����Cxk��I�vv��B[g[nm^�zU�֬�R��"�� q��:K�4-R���$&��r��%-��2/~�����$��^���J�BNo�C���fN��v�	����8y�����kxR: #|+����@�'AN�VT�K*����a�;Q�MvvQ��@����a�R&系FUl���K�k��P�0tQ�P���.HGG�D�_Qг�E�v�s�@���i�i�uƘY-�]h�]H������~�-�jg��&���,����0.S͸�{�\2���3��Bn���p�M/.�Ȍ[�����5a��6�y�tf+�8C-9����-*`O�����Q��\�L��"���^[��[]!���W�O���-$��Oh����M2�@�"h]�L�.����V�2d�[)y�X�c��m���Y`�\�)�e���K2�/�Eܻ0���ιv�4څ��?�_Yc/Y�œ�K(�YR0�
˒���	N�U-D�qc��b��Xb��md�V�KfoFh�л0����-L�W���)� �Pkaj�3���������g{�w$�@Sv*t3�yY)��Ei<Īz�-�i�pQP(V4-���p����K�FZ�U���k�	�IpM�(��ge����FG��
����m>���l%�[}w������s�8�"r8�n�B�4S���&�7G��[�e���6�����p��he��0FMWYE�k\Ҷ�t�|�%��Q|�����*crk�4+/,��r�Dҫ~�ʻ����q�N�7��l�G�Q�.np��t_���K��vvI�6��wF�����Z��v�5���1�^��2    IEND�B`�PK
     mdZ���I �I /   images/ae036c7f-e258-4627-a75d-99715ec815e7.png�PNG

   IHDR  �      MI�  0�iCCPICC Profile  x��||eE���6�G��y�]�$�{�R�f�IvC�]�%�l�l#[`�H�"Mw�J�"�T�"H�&E@`��3w�N�]������@��79�Μ�=��{I���挪&��y����L��ǞՕ^IF�u����X�����#�Ox���{�%��H3������;sp�@�4,¯X0��Q����- �~��{?G?K�0��g9z�xǓӛ8���V�)�V]20}�n�$���^�0IV�O���Ṡ=a`ͻʅ��;s�̙I�*$�̚�x��ci̹���A��$c�Z�?<+I����{�\�FЭ�m����%�����<���L�Ze)cͩlf���:��լ�y��C[7MV2M��4�9�5�kʴ\����Ӕغxx��6���Y��"��t%,I��]�*��,iƫĿ,1h�HZ��x�*��&��;�%��I�8S�ׄQ�u ���M��{���K�<@u�ǵ�1c�%m��&���_��^[�/X:<4k��j4m��>o��Dғ�,�6�~{��ǆ/<�����{Hl;�$i����6�Q�\�`��}yl���d���䶶H<os
�R�^�e���vLrjr^�<�6�-y y2y5��a���D�.{7�pfõ5�6j�Q٨�u٨'FWF�0z���F?3f�1�c����M��{�������J�4o�ߎ�x����<q���X�UN�����U��j�w�ֲ�-��կZc�5�Ys�5���'k��k�θu�Xw�uo^�{�W�?�~��6��l��F�o��&c6�vә�m�ك�[m�b����R��~?�-��f�׶�f����ŗ_�撦��;�֫������fױ���`9G�g�.;mۮ�������p���|�̖�&������4~�;��~��]�w���ִ�Zw]�}i���'̘��5���s�7.��ߞ�w�^o����3�ۇ�:b���6�7<�w�6�Ȃ��wZx��K�?p�����!�~w�CO9|�#N;j���=f±W�k�?z�~'�;��S[O{��#Ϝx�o���ܕ�[~A������{~���/�����g-WO��랺�7���C���֭o_�w~���w�u�=�w��>���G����d��G<��s�<?��/��ʌ�����oLzkǷŻ_������p�G>�+V�~����>��kWrQ�aCo�u�6u��7F����5敱�[w܍+�3�:��o����q�������k^���k߾΃��y����x�57�������MO����_}�1��&4Ml�b����Z��q_>{�˚nn����W^H��>�b�\S��76���m��j�ݶ��C��{}mA��Nk�x�umw��ؔ�v~��cw٤Cv�:u��.����Wz�O�r�λ����=~��/���7_�֊�u�ڪ����͜3�p�f}g��C?������s�܇�=;�����p�EM��[��{8�t�A�|�!˿s�w�;����;b�#�G���|o�cf���#����x�'.��U']{�/N��ԫN���K���r�yg�u�i���Gǝ{�y���\���2|���ɂ��]����.�t�V��uE�\��U�|�Օkֹv������冎w����C7/��!�}�I��s�%w\��_���>|�ӿ{��7�~�����}����O���~辇��í�\��������'���'>����������n���]��U_���F�<�o+��ګ������׶}�o.}�^����<��'����m?��Ã����n���c��_���a��Fm2��Q���Yc�{ĸM�ݱ҂�ی���wU��rƪ'�v�ꧭq��W�u�������/���Fo�ކ[m��ƻm���'n�|�;�O~�/����Ħ-v�r�V{m��ˇmsJӏ�^��+���gϱW���ߪA�dV�kl��W7�n���-;N�ڷ[�O:����?n�f��Nyt����٥���ίN흶���]/뾻��cfL�m��{�q���o��[��{���x�l�m���}�f-�}���^���s��Լ�$��1��B��m�nKfpЁ�/=�퐇���w�=l��7;��v�nG����}�ǝ��K����[N�������ϝ���/���鯟���>�ݳ�;��s>�ч�~p��x�G~��A��$�|�����m�.���/?񊣮<���v��O���k.����n����w�#7>yӳ�|�����[>�������z��l������~W��߾gֽs�s�������>t��G��GN|��?���鏟�������>���9�f�_vyv�粿6>��c_x�����ˏ���Wn{����������eo,󊷮���8�����{o�k�k}8���Ώg~BH�#�Q�Z���>�ר�G�ї�i�_{Ӹ]ǽ����g���ʯV~�ʕ�^��٫��ƅk^�ֵk߶���>����_��FS7^���޴�3��_ܲq�/�3ሉ�mq�m���o�n�6͓j�}e����v6�D\-oU��G�3�o۾�ݘ���a��k-3'�z����~�ӟ���>���b:v�\:�G�n�z�{t�����f��Ż�f���\�͍�%�=�o�^�������|p��}�����7�>�o�9��m��������?|���-[��%���_?(9x�C&|G������X~��G=~�k�4��q�/�o9����0p�ܓ�r𩇜���;��}�1g{�������=�S�?��.�鏯���~�=���O,���G.��e?���+N��ȫ��Q??���9��s���/.���n��������7��WO��̭�����o���?�͊;G�n�]��W�g�{W�o�}�����������w<rˣ7���]���O\����<��ӟ>���<s�_�x���������^<�3^��o��r��w������X��-�����o���a��޲���]���g���Go}��O>\�p�����$��W�x�+v|;i��v�A���b��$+���O��ϕM�i_J	{�?�d�3�9V�qi��=8�?b��}oJ�2<88�?pm�|�A+6i����4�����c߲$�UW����Q��5���3�%����e��@����o����	���u}��_�{������ہٓ��z�7^�34<�W��M��(��y�Q4~���	�Q�x��׳�
�Q�uo�w4�)_������������=�� ����3�	���1��ch[��������1�����;%}�y��H{)��P�8|�/G�C�9����c~B*���~-~9������8�$^6f��(SX���t�{opPk=�#?�w�J�u,M[��I2�,�;�ڒ�I;�lż��[�{.r#���F�m0!�OݚZ�O��c!zP�1��1�g�i`7m��A����Ջ3��įyJ-#w��	�x���a�i1ֱ�>˝8�A �!���2l�¦�]IS���Gq��k��m�')ᘉ144�d�2#ѹj�g\������I�$�d������I�3�)������V��Io18�ªF�.����S}H�K�y��o�9 �fH�#���a�_�-=z���;u�e��O?f��>��/�����ygo;�V���䶞�����i��Ɩ�YK�̩����{����y����Y������U���3xn��X���>�}j�Ȯ3�.��Xi�nk�m�\m��_T��_Ze���m��V2Wh��3�[��Z;Zzz����{�:Z�h���O����7��������nZgWߔ�=�6�9������cZw_w[W��{ʤ>���JoK���޾��=���;ۦ�Vwo�Z4Xʪ���9�K���7U[�ϙ?ܹx�~C�����׻GW�ݩ��g�j��i��ˤ����v�7k�ĉ��t���v�t��:�wBjS�s,��ur'�6ZQSYfLZ��&�f,�f��eJYf+S�uw�t���6��wZ�}Y�V�h�i��h��6��czo_+&u���O���5���}RG�g�Lj�I�A{tt�AD]��v��=��%���gW��{�ͭX���@(IԪ�8�E�3�-�$�i��fj�ƫ��fV�o�쩲ZVc���N���Xi�:�t�ʴI=m�3ڠ?��Y�t:�8���ul��so���v�7��?wwC��i-m��܎���Z<s�ҫ66�xz:�M��ySWKo��}=m�NoñT�u��w��/�0��6KþHE+S�wNj���Fvjo��S�^ē[z[�v�����tvu8� M�v�Nq���d����=ܿ{:!��=b���ޞj��9*�;�O	ae-�ˑ�5m���v-�kZ5��A�xժ���U�j\�TU��p>�?�'�y�ʈ�3�,�"���&��*����jF()����(�?�)�+�*��헱�`����if������Wߏ��폣#,R���Tl�s}?�j"���^���6j�BK%KK:[���3!,�X�#��Tq]�FhL�;t�<�2ص�0�B�1�T�*SȨ訲��;�U��4g�E� WX*/Q��Q�,�R�V���W�&��Q��]���L���t�����Q��>2Yr�E�@ڌ����h�N�c��d����SS�IH+��"}͠yZU2]r#w��dF�1C�R�V2�C�;5nG�%��P��:�D�l4��b#�e���؄�n!ӌ����Y��~�a"-#���N��L��RCH���L��t�	bK�;2iXfhaIYa�jk&�L�� �*s���-Պ˨�e8$zTPB��dF�\2Nrˬ��W�p��=Q�ϐ\a3Hڱ�
Ù�֌c�'0�`��X-�7X-�<����i5�S=�jLm.�GB	�rH˰5�u��J�*\�N�8b�0�e5�H��'OE���8t�tC+�b�P`�2�_G�@��K��h�(��@�Lׄ��'�a,ܶ��H�Y�K����O|tZB(,�Y����Y��5t)K��p,�|4��`�2�DX�ܱ�����9����`�$�J��s'��fp'4rYc�l��@P����AjI�X'��TX��1�f�`Ka�i�q�Daͬ�U�ۚ��:"#���+2xr���`2�G���VO��+�|�G�N���q�
�Bp�N��zlL���R(-�Xr�U����=Z��z�R+;��C��x(�+lj��� 6KDHN���RؐU�����#�o��?B\�� 6��`�h]i	3ѩ��ㇲ< 8T��p*]G�L��
����3tU�FZY	A��*�����*@*!)����3�5�!�#�8y���P���#���4��G�Q��a��m���@��4�O�b�Va��La4�j	�%�����sKR��"2���I3�	�	djA@a�z8bBZ����R5l#-#0��� ��=[M�� �O�������:� �}!��'U����H��	�K#SY��&AJ��BG8.V�r�����3@�)�E��n�H�g���#H������r)&N
mD��M��:B�#f�VaVP=�� 8�
,� X��zB���S�,I�Le�uոF�u��E�J�82,Ug�Ȋ4U#�~c3 +��%� ���R-�#С4-!�aN��W��lM"��w�u�~�	!g	�}!: ؊ʪ	�%ͬ'4�6|��3򪁓����΁�HR�z#�;9�0&D�j 2,��0#�'��0n�V
@2�ei�:
Gk�_Gg�wZ�0�0�=��
�����H����`�kI88x�;����TI��:x_B.�����U�.�"T^Aza�X�)�1r��ʔdqFV�+Ek袁����%�Ṋ`�@��$�P��dP"�iI�St$?�p�Q��a��`�8���"kD2��?	���SV���=�w�_��Ffjd:d���*�����:B1�&�H��]«�E�ˎ�H��ړ�E�p5h~1Q}G�S$q������!���ܪ�����B�p
���	/	к$�ǁ@	��q@�̳Ba���e,�qF>�.��!�Np.�X����9�T���I��������8���!� $mG@��b��8���j`�@�
pP�=��)+�ē��QPG%a	J@&,��(L��F�C`^[�R!#Ќ��Đ����`�1��3��-t�Ȓ�����.P��I��&CA>�pTI�u `:Npy���RE�-f�n����3$��"��rW$A�&-�jJ�gGNF��� P�N!Q�[�b�{kT.%E�y�������|�: "r�EsJua�*�����\�h�C��22Eq���\|E�d��*r8GFi�zd�by����T 02��4P <��a,� {՟?#�,.��Ud1CE*XŎМ���*!j�����LUt��XU�1.��~� �
(oɬ��K ]�K��H�R��=�T1J�B�)q�Q �F�{4�k�Qj +ǖ�Ǣ� -l��9������diY�)�F���3�`=�*ziV�3.�TQ%OQ~&U^�L���#+q��ڦ%o�H.�z�H��%�5*\*rzF�Ukx�	 �z��U8�`�Zr�H�r[���^ZVE.V6�����P�.=$���eu�'BO@.�:�		]GO�8�9�*�q犒?�����r�)*��e��'��APM�<��*|���֖G�ZJ8d���K9׬	�W��rr�
�X��^�x
NZ✰s�YVO�=	;�dp�]�ӦH_ѓ��B c
�M���x����D����ʰ��PM�Rg�%���Lu
	!.#�4��l�49�R@�#k��=���Gғk���G�7z��Q��8O�8eje^����}������i1�xA+�Pe�)X6��� lܧ�Q6�ٙBl��Cќ��g�L)U>� �*���@���2	�!�ecJ$YZ���SaY�T1B�
�rA��Q�R�F��+�Ѳ0���9�L��)��t�ʞJ�U��K�&���\�0�.0Q�3T����*~�*2T�}�����zO�oJ5*�P�`9�T%^3j2K	�T�2N�mI��.�Q%�8H6lH��@v�D�dkJ�eѓ������Ch��AO[�5�*�'$�(y�礷�4�)�6�Y�$��-�	E7h$�?Nn����5�|W�'���d%ޤhAb��@��p�F���	�l���'M�w�0����<��HL�x�(!���t(��t
cq	���SD��s�OHN������9hp��FGM�T����ܺ!�AHka %=�j���z�Y.[�|�{6�~f��ڗj�
�H/a̤�$\��en��IپѮ�! ��
As�2�OX�QퟜeJ�#���Sde���*����<�*דe��dd{�$-!0|�����ؚ�j�Y��d��WKuGX��tr���F�y��>��EX�9���K�U�r�h+d�q�j������x��e�:�!�zF\,���V�P��9u	֌��!mQAO)X6�>�'�iJz�}R�����@�	���@o�-�#�	�j�m��(�i���2㊚��@J���G �8�Jz�-�Ee)��'U�8�s"�K�$+�Y�jP;�R���H����%�6�*l���)k��<|YA�)E��-zRI�%�B0Տ�t*�S�X?bvʌ{�.�ӤU�C�T%=��a`��ӣ�|NI��,�Cq�4g���m������)�'�-%������yM�Z����$W ��gĜ�QO�!!U�:�	��=��s�|�XV��0uT&U��_R\�G���)�г�F�	�A���aD�L0唝C�/�秽	��<x��E$���D����j�� PL�,�E$�&J�D��0 My֌�"��E�h��,�*d����X.�;Iݜ��J��k�i�a70��\�T�6��>MY��	 <�D���!�/���e!�Є����=���{f�t���'l�c�.
��I��,$�G�P}O���hr+&�~Nn��n`����i��פP�f�b����jt}O*	�L�,^���ԓЛ%��I�� N ��P������ ����e�� �p�L�*t�����N\240����=�����z�����^�$6,7\�d����V���0�{�=V�g�YW��Ɉ��-���Y�y �K�U���dPt1D4�;`����DO�讑�HXmޝ��5{�������?wh��>&��x|��������G^���*K.I��K�t��������4�:dP����H���H�#T ��{�JIǫ�S~%y������ h�/��\+]��ܓ\�Z�R��x)���"���D��c�����U�hϵ*:u�I���"x#^�������i(�ʽ���v{c:��C�-F��Z�I�����YF����7C�ܓP>'(�6�KK��V���rNbk������(�V	hH�ؙ�� xG���'vҩ'3����>�@J�xuJ��]�ͰObe~9�N<W�M�|6hDrR�r#����f�5�(=i��$N �t�HQ�o���M^�j�#�*_��õc/�A��)����O.(���� H3?��t�x���4�<	8�G���+�$\���f�̌_�R���r�p�9�?BA�7�F�T9^�2g�)��'�Hs��HL���8A�� ��ۚ零,גe䋤��61��taF伂�3g�������ʜ��o�z��V�F�7+�n��.3s���K��]�|�J��Ѝ�8�;��q�/RYDG�QE/�u*�Z5L�g��t�Ϗ ���,7͜���'��Z�x����r�.+`�ĩ�n��Q� !�UH&o<��7'�4�U�+��kԊ���@�T��eF�����^+h5�!�;^���{�X�C��C��� 9�ίݑ���@�4��u��Y�9��+H/�&�nq�2�	�ȯu�d1��+9�M�l=7�)xh�T8��M���>a
E*���b����
�IhWn�E��j$S���o�.�K�+��X�R��
 ��"e4���ר���?�"��I8O��+DՉ�Aa��'�:�zI%d����ݞ�ys��[--���^ؓ�Y�\�D/H�DR������b?~0I�ϓ����C�k%���Q��y)�z^���!E�Γ�%�$t�xYD+oR�@f�P{�y�!?�%��t{*'c��%g�[�t ��n e�������O�I�dA�G�xe~A�Z�~0Lt�H�����ێpL���T��*��y��`B~9V�`�y|b���<�E�k/��כ�je.�y�Yo���qs��j��
I3�I���y������g��z}`)=%�y�������R��/a�[-��� )� S���]�k�>�_/�f�	@f��Y�0T�5�T��@�ԯA���,�K�t�5�<���;o��̸�6��Ht��r��Z�]�Ԇn�3^s(�Z�(Ȭhu�s^�_���w� Y���cO��10	�)�[�)�7r~0�% D ������A-��)��L=��0��n\x���@�5�)>µ$bk �6d��Y0�	r�y8R�\�<bFK�ޜ�U�[`F�@:�8�!����pR{�����GÌ���	�H�<o�a�h8X�d�4>��aA��y���*����!�����F6�*�y�0ٗ�cH���Z���a�n�$O�g1�����P�D�j����Ѓ��7���"��{$a����6b��-0���2�;fȨr����cz��@fao@�1M+��9�[�V+�z#��6��b����O���0ئ��	2�L�4�g���0�KY��GHNI��[�0o/�p��yxeP6La�#$���pł#��@	£�z1��}��ȴ��ĆxН�a8%�~�Ȕñ 'h?n�0nһ�i�:Sx�2��@r;�!R#�a8��c */I�a=o�a����Mʤ�k�ƹ����0�),�f���խ�Kg޽�.����<��X�v�#� o&<o�a�~�
��o=)�q#���r  ����E�"<�'2����rވa�kK�Dz?)�=��@Hʻ
J�6-��T�⁴<�J�x,"�p�Ap
>fa�J�q#�4Ͳ�aCʺ=�ټ|#�����D��*#�F{���2�w
 U87Z�_o�0�|����7S�,�mHD5U<�Z�CNJ���a���y^)����SE�04���
�~�>:�y��a�=�,�l�y��H�b�<����d�tg�������^��0��>���a��� ��ԍ+-�����މ	XH�T ��ވa�+B7��@B�r9Ȉa�o� �ӤB�����g�ܬ�,t���(1t@z�����Ւ
��>Ȉa��ZRp�*S���1�D����o��/��LF��5`p�������`��JŞ�м"��T;��rO���@d�0�����
#�u�[`	�*�*�I+�<VFC�-�@��W�,�Sd{��^s�C9o�a0�I�$G�y��?��a(���i�f� ��a$!.H�2�|<>��H�_A�*0�1�:���'Dw��"�A���R��{�,#���)yH+�a>���H�.���9I�L��"b��0.`uX}�Ï1ZC�����=�����:tCLR��T~àU��
�WF��v1�A5`�q%|R�HJ��,��4-�v�y3r
8���W�o�a��PI�,ر�F��e�I�:S)���Ak���2:�"��-0Z�<�D�g��sSà�����������yC�}_cR��>���|MAE��>H(`�i�k*b���_Ae�O�gY�&�"��O��@���1���BE��)x�R��ރS�������x��OY�:ӾN�"�Q���p�W�l<o�aEw/>D@�;�U��8*bEy��K�t1�x#�Q��^ri�~�=o�a,(���8��vz=�F�~�!�T��G��y��Tg����0
��?'��Ǩ�6#��v��/����/߈aa]0�B���X1�,0hHj�*b���^��@�P�R�`��0h܊���a�~�O��\�n��>1��9��t9�y��(k���7S*6{���е��`�' ���#��pm~o`��`0�sH1�Ί���{Aj�uRGC��Ҥޤ1��8UGC����T�����a4}7U`p1'��up1r���K�ky����g:b�|*��^$�uC~� /1Lx�����g:b�qo�#�q)�;�h�>^5�i�b�3���a�^�Oa)�
$�g�7bL!y �GP�i��-bL�|��y� H���1�PޭhE�<I�sވah
xU��Q��c1C�FS�ɏ��w�1�~R�TC�1KG�)����ݐ�r���a�<��C87#��/t�0T����i±y��#��!�j��?��M�wL�0�>���[�U�L�0hUAa(��Wf�^J��0huO�2Q��U��(B𴆊$���+ӷ�x]7�P�wx����t'�-0�zC7��0��y1�f��>��I+<^7�P��;�$�{�D��"��V$���SP�e1�c�Fp�H��&b�
�4�
�M�P���-b�J_7d��|�Dcx�쀀����j=~�à5�����p ��^'M�0��K����㐉*lP�d��&b�߇�TW�����>U�ݕ�a��W.�u���;��F�1 ���&b0J�@NH��xC���� �I��}��Dc�{����k�����DCu�`8�Ӡ}�a�
*�=�F�c|��D���zhv:�q�0����w����R�ve#�!��^+��QXl�-0dX:�V�[�AFxc�1e�!y T�9[��)|�l҄q��ue1��/��l�O����xa#�J�>�b���EK�Ҭ�-0�ʐgY��#?�Kp���06sϸs�4�4��h#���4l��C�|l������\�#97�y��A$�BH�y��t���җ���s�P?e>^f���}/,�y?��S��>Y��
Q����-0��Jc�P��;��[l�0�A�0�^�2��8��X�ҍ��B��7�I1��YAH#U�Fj#���c���.Hӕ�-0�h��?�q���ECu��7v�����ك�MgA|���6b��p���0N*�-bk�2=�N8Һ�Q�[`K���y+?�Y6��.Z���k��պ�3^�N��� V�Q(&�[   	pHYs  %  %IR$�   �eXIfII*     (           >       F   i�    N       %     %      �    �  �       ��    x       ASCII   Screenshot�M_  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:exif="http://ns.adobe.com/exif/1.0/">
         <exif:PixelYDimension>512</exif:PixelYDimension>
         <exif:PixelXDimension>960</exif:PixelXDimension>
         <exif:UserComment>Screenshot</exif:UserComment>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
ǃۥ  ��IDATx���#�q����]n`�(�K��%�
�,9��c����؟���e�z,[�
�dٖ�s�|"0o�����'l�������\wUu�d6��P��'��⻊����Z�ON���1�R���8T�Q�s�(���ͥ:_8��U���b���~HgC�<��L�^�0z�N��?+��������m1�N�6��|f��ǧO{6�鏢�Yʷ�|��W��{������Yw��W��[ǥ��8��-N2��>�#�ļE���h4Jф|�<x��� ~��,"�<�d��a3��#���*4]N���ĵP���$�H�˗,>�N'���W�U��p�>3Z�<=hmQ��흠��>1=���g�Zz�\? �_U�~kݭ�"�
�
:n��-A���D?T�z�
�րc�U�]���6]����U�e�.Ҙ�?0��~�f�����s���VX[[K�Js�������[�ӫ�F�_�$\��8�L��c�TNt0�VOv�a���|�b[�����|������/�ЅwٽӠ��|��>:Ҧ�\�1T�~P�bY9.'���ӡ%U������Z�����;�y�pKZ���\���<�w��;5�;/���+_/�.�g�_+�W���<Fu?�`k�N�x:�+A~W!�1T.X`���=\�2݉�_�X:�q�`L�c���r}�1u*yz,���i�f�gss3<��c�ܹs�Y�-M�g/\�z5��λ����p�捰��_�t|��4�P�� Հ�N2���Su��G1��c����Z�frK��EU@��=�)N�����3��νC^��F��$t7�! >;*M���iUO�������30�V����I�[��� /�ʻ��)/�Uˇܰ��ד0;�LZ�$��w��ቡ���h���1z�����>ht��e�[�=�9?�7a��݃_� 0�
l�o��b^��q��X2����˗�K/��~��p���4gx�P�۷wo�~��_���_����67Z |��	.���i�nai�@s3 N5'��8�)-���'+�h4N�߃}*����֝i�Y	�	���5qu�f��_�zH��L�&x�L���x�� )N�����A�� ��ڟV�>�<�P_[�����K��-�����oЋ5��_�>��  |�v�r������YQ�]��{H�[� ;�<�� ޽���駟�7�|3I�ڶz�|��m=B��a3�r���g�Mװ�766��1!߃Fq}~뭷��~����[oD ����f�a-���ͭ�1YK�Qc�;o9>g-�nܞC��d� ��v}x�5���{�����5��VR�ș��/���S����YY�:���e���4����>��о�������D�)��=��]��t=.˯��׍�]}��]��A �����Z{��g�ƍ� ���,�C��>����x7���KН��#u�Xwem���b�ʿx/,�s��q��G�w�}7���;��;E}�����Hrun~�wvv��ޝ�����ك�o��W?�$�5�P�s[�a{}3L���H���:
0���w�m��z�d2�@�`�wn�����"|� q�\��6�Q���yb����_fNi��$&�t%�5泚�\��W��JJ̓c-��{�t����?���%�>���ԧ��,��!.^���Oj�+	7�t�F]v�6�΂�R����Eui����	j��<�Hx���+����[�� ^u�q��s[�GN$�UZ������A���>�����M�x`X��ӤU�>���R�a�%��_!y�<o� #���{'� l�Uam�����h���!ovo� x��#�򗎀������724����������X����3J���Z�[h"���g�Y'� X���_j�U6��{G�s ���q�P	�� ��T��U4Q���åHvՁ{h�ܥ!��vq*�w���{�V�W䯣|]��޻�ƙ^;���4^J֓R}��Y��g�B�4�zh'�K<X�~������4tO�}~��q�i_?誳��]u��(���^z��
�,����R9�gi������gK y�K��{�Yg"wg�����d.�E����D	�U]��;��r����9��q�=+Vb���`�&���+���d�.g&�T_���g����I|)���De����d���\�_	��j����d�Ű {��Zl� ��m~	���l�F`;��*�O΅͍I�6捛a��t��ٔ=ވ��~��<������L��k����;��@����!��P��?z�F;�ׇt���u�~P�8��Kx��Pu��c�	���V�w��!
������R?�y�&P��_F^3k��#�>Z�Q�"�׎v���K�Ք�n�c%_�r#B�˽e.�~�����f~�A�8-)�ğ�������eTj���rH{��McW��K��$�x=(��]�t��a�{������x-�?�}�/��<�?���JϞ%�r�燮!6P����K���R:�n��������������m�X�U?}k�W�u=o��`ݻ~�zq߯�Vk糖��A��E]�� ���W�l�ݫ��Y��*�ҵH�� �!J���)�:"H��Gv~S�+;���5T6Z�,>ݮ<;��rC��|�f�� 'Gc&�����L���@�L�ur_�Ų7�VXh?��N&<�o}��g'Mo�O2�l����n�[��aZ�c�'	E���a��Ԝ��X�����=s��z�Ĵ� �Ӗz�����:	��XvѴ�>C���Zb,J`�-��ɧ�*8\�|���C%��KNX/�siL�	�}�]�-�> �E����կ�e�٧���Ծ������2��oɼ�
 ��ǧ�2�Z ����_]�Q}<�{��>����'�qi���6]�<�w���y~l�����N�|l:�����궾�*&|�]��T'�G�Nu��ǰ�4[�,��n�J롵�x��y)�Y��w��E�_�[���=�*�Y ��7!,�dJ��X}�g����J|�B��m[~�J�����K��h�vm>�@#�6���ߺ��и��0��`v���V�Y�Z����0�J��o�[7s@�Q�����)�*<hћK�m���B��ζl1;��t�А�ى�.�C�9�2b��>��:
�Z.�{�I�p��Z�&���a��8{�-/	A� �;Q���l_�g�X���*?J� `�;Cv~����U��*p)�H9�v()X�,����<���UL���-����u�T�[շ�&�mo�Yo_gMj�E� &�+�z��d�g��.�-��Q߸��i��B�Zy�ȅ]����??|�_��O�����=�u�(��} ~UZ�E�3�A���|�i�~�N�-�%re�M ����
��Vm���u�$ =��x����$�'0�lT����,��a�Ϊ<7\�bk1�r�-�V�_FVkۥ��sǥe���,�g�ZWa��U*�ݒޝ�U�7}�:q�4�$�'�>p=Ԕ��C$���<>��!��V�� ����oJ�Ew���|o�'^�0��þ��,��K�(uKn��t��}�:�?����s?��oyź-�O�N�=_��U�;R�.�W�W�U�|�Ix���������$��F�b/�+ ^E	����RV/�t�U�c�c^ã�}����2���|���c}�ħ}�?3��.Z����\6'=�'��&Ϻ�M��}�c ���t&���ws=E�^�����D����N8����x��zV���	n�| �^8����_H��:����&�}�i���kq몯�Z��
�ǥ�L<}4DYR�= R_V�U_���4�����G!�!=��P_��C��%Z�>Y0_�C�[P}p��E��,�\K�^�K�����Uz���t��=G�oY��_���O�q'�! �ӽZ֕��ܒy\E�C�
"�3wr�6ߌ-��3gm\J}<X�1���u�« 7v�m\��u[���	�\-<Q�V�6<�c��z�kas�N�dU�Aճp�p7��������:L�JD��[v�=��P�m�u�Hi���U�N&|�|Zց$2�wi����q�i�]���t��� d�9m���˙�j!��d��	��G��T� L�R�,��<�Œy~U���IP�E�� �:M��U��l@��'��9Z�����2��q4���]��p�׹�|<�Q�xj��.����z�*�<����g�C}����U��s%�/�����!��~�z�U�U�Q�#�(r��ݸq#\�z5��
��u�����~�����gM��w��Dw��IF��c��͛i��>א+e)��0,���?_.��$r��y����GR-�Mb-�ۃ�cU��fweY�g�g�d�iM"��Xas����gaRM㇀[!�>�,=����<�r$��Fs���`~��RZ$�4�&s&o�3|pU�_HZ}�>+��� �O(,�q�ɲ6YF��k,�R����k׮�� Ki���[�#[��X �Wά�" ^�@�k	6���_����W��zDp�ڊ{y��-��N�o�{uQ��rde^�mK�WRT˒�jh�kW��"[6��R��<��.���w�eW~��t_m�Ǐ�5;����"��`N�d�tEж��Wd就| ��J<Z>}~�~d�~�+YF���Z���+V���æ�<���i)�JT���EB?��C+[.��%ߏN�\��4D���ѽT��r���q����U�:�|d`a�9a(/%9� x��u�O�8
���O�$6k
>��Io2�� �l�1'sR�	GIV���NA��>ߪ�uh��Vurw^_��q�܈1����z�X��'!E������F؏�wo/�iS�e>k�6���</��=C��w�z�tL� ��_z���3�$w��k���w�x�ôJ�9��ㅩ.A����=�G���n���2�o_�k�Y�Ӡ�]UZR*ض�ڰһ}��
_6��˗�ŋ�{�^��t_��U5p[����F�5�&D!cgg��T}�Z��y��CY��k�-�I\�H��I�7eT�}�
���'���X���� O��-'��t�R�����^��ޑ�FW���B�4�했Rp �_�;]|�OzޤQ�S��tIA���C@�T��>�S�=s!�O{�zRTX}�G?��:JL��Wikڎ��oܧ��|y��^�O,x����r��D��c�q��4�~^
NRk�A��W����y��D�3%����)O�i�,c��M[�c�22ƴ�L<��:���HSc����=�7��.IG�6�g���q�]��n���ն�S7v	jC�-���7VK����م������?�0��4/���D:��?G�,���h�]ȧ k�6=�G�N�y��dh�ɿ��Ɏ��ր��1$�e�Uc�O^�>�:�$O�� ��i�������m�i:)?�N�YA��m��E͞\�=���s*�$$��9 �k}�ތ���$.\qT��(oEP��HX���(�~r�f8��:�1�a8�� k�g�2ε��1�=�s�q��H�G�c��������7�x#|��	Pud	ڥ�$����t�m�E�@{g2o�?m*�!����Ĭ��!T;y���u�/H�:��6Z�j���],=(�˶�/_��|B{�t�հ[�Ke�%��G���|�+_I�@���)ݣ @p5�������>^|��������GM}�=X���������I�F�ꩧ����/~��ʕ+��'�̀׶(�"�~����^���o�@�U�|_�P��������I4�x<*�Iڀ"���׿N�HR9h�r���_Nc�믾�j��������.	�Hٳ�,H� Ud�َ3����'m�����S�׭`j<͡\��I�����sK��f����]�T��_�� Z���^��ַR{��'������-i7���ٟ�Yz^G��'m���v��6�m	x꾵<��ݶ������,�'���/$ ?�s��/�}X������{m�⃾�H����}�k��7���L�����J X��6Wi� ��d�S&�Q�����i���K��8|!��/������������CyH[i���?o��vۏ��:w�:.��[�ft�>�Я}�4'VV8����>�Uʺ�����X��+RV![&� �N���(|���_��ϒ��� p	,�|m}��G�cUZ��~A��,�^JsY>�i���ݯ��#�
4D�-��%����t�C��5�-|�;�Pr��q����~�^��E$
��J6��ֹЙ����#p�{�����|��z=Y'���w}��a
~�QH�sD���F��&�\E �7�4>7ۍ	OHo��%ñ/��҄o�*��[�Y��o�[d; �o� ��\쁅��I*	�>Z��:���Y!.y�G=��z��[�TF�]W��o���W&,ȵy�c�ҡ�R@�Hp��oq�����λ4w��G�?ib�� ��+�\�B��
�r/o@���_~�s�KB�����3�{&�x |(w+���F�Q�з_y���o~3}�.���K9b(@�,^ +]�I�A^ƌ����I�V�� E�f��x�	 &? 
B7�l�e(E�PQ�e�O��U�L�]�PB:�J��������n�qiN�}����������T�3['uZk��Mwk��²���!'�'���vPtX���+WR?��� r�ԧ����5�+���`���m�)[V	��\�?�H��7���|3����)�,X}��m �W`�y�&}�5`i]�UVՓ���,��t�Cx�1 �WD�%Ɨ�[z���yW<X��˪L���dƯP���E�ط���Y�*t߳�u����3���X�����~�Xx�'�������S��4.���P^��+/�߲���K)�Ө�ߟ5�S �_��c��%?� X��P�6$�㌇���Y��J)/�j�o�����A�k�<gd2���L��(����O���wTf!�����
�.����q����r���n�O��d-��( ��F��m��au5T�3��]�!�I;�gLp�+rV���j���oΉ
ᨦ�n�]Xd~����?��!>����� �RK��|'�{� ���@�q�%�z�o���x�tX�´��u!$|��?%��R&ͦ/K��`�}���Z@d��5�zhy*��ǥ���>
��!aW���E�DX���O�#���� �L.]�Jl�& k*��"�x&扒��<X�l��
� �����HV9,�X�x ���pN^�����SN��0�w���/@C�k҆�w�}7\�v=$����9����$�"|�ՇPB�k����T�C}U��;����q�Hm�t ~�_�>(�� ����T� `x��4kW?��S{�tOʉ`�c+��j�Ro��SYJvQ}��P��>V�3�}������c�O>�n��8�/�<,��#EƄ�W�x��J+x�?ұs�z�M��C�P� ͭ�O�ؼ=pU?�s'颸�?��{A�Q��ۄ>��	H���'�=ڍ��7�"|Ka�~C�<o�w�L�q�/��^��S�ȸ�l�޽[���q�y�@���%��2/��������-�iX>�<b� oɒo��R
��B��[}yڶ�s�_�|�C���Qw�W�!K}�t��j��i��k�;ݖ'x�\�l|w��7�j���v�=rR�T�{�Y�^o, ��c�0
��aInv0�� ���m,���8Q��zC�Ո���X�pn{��r�U�J>��m�T	z5Y�X��G�����ݙF!��nޞ��}
�s�&C4���]�6 ��oYr%�'��E�sj�%��Dأ��@�� Wľ�f� 4��g�=�>=-($`x�tq��i�U��L[&+T���Ez9 !�7���,| |r]�>0��V��;`H��P�`J=S�0�ǖ�
Q�u[iv	%˯� ���xF��h/�-e�9@��R�����(�uM�|��kڟv~����:>��t�>����*+��#��E>��r�������^K.���� ��m�5�4 �ԉ�zEM��r���~���P ��C]� ���E���/�DVC���/^­���3n�t�~c��o9��.���C�~�L��\�̌�J�G��{!=�#}��G���l�[��v��<�4��+Bc�׍���e����ӆv/��7�����æ��}���M��◲����|����e=����n��>m6j�@��Ϩ���ui>�B�ʱ��պV{e��ԯ����r�*�ER4���"omm�J˻��T/�3x�:!A��Oj�,�������K�ui~� vxmY,0�T���w�Ǧc�W�'��B|�ս~{O�*���M=�[�Cv��Z�����C���j��mz�V�sd>�-w�F;���;KF��5Q���ſ�yPPg&�[aa(򹹎!.� �:�N�� mr��A�I4��f���1�D}f����i�=� "90V���m4�#,Nq����Fu\|#8�~x3�eO����U
2�+�I�|V��Rm]���G��W��KUڝ&M��[��x��p_��W��p�p Ṵ�N�'��G?�Q�?�ߤg]����u�I��_��_�� PN�X�x^�5�
�"+���� ����/�2�;lJ����W�j�	�UP�KV�8/��=|����r�g?�Yڏ�}kV�n'���r�F��+շB!��n�K�}����G��
��ީ��~k��q��F Ex}��˩�P@�7�Pq�%[�<�#��' ��E����k꟔�2#��mK�Ҟ Tܘ�䵸O��=T PA^{���O��O��ڀ:��Z>��bY�e~ȏ�Rn�%`�	�]J&��\Ե7W��� P 1��@"]��8��S�♼Hߎk~ÿ�+�(�
c�|H����ɇ��7��G T�RQUIW�H��〴�G�ȩ��󋢳�*��/+��SҁOx�G��y!-rq!ݹ�>����]�}�w �|ķ��\����Ǆ 3��
�Fy�[|�5��@@N{��ԝڃ{�'ρ�|nn��{~��UX�+��������ǁ�7�)c��	���W�_ xU��$3�,)����Z@����vYյG>�)���[�B�+�炽fA�W�����j��ѯ%�i�R?��v�k���ȳ.��{�!_��Lp�<K������]1IF�Qg��P�C�|]ƃ.*)TV-�C�7��0�����jK�oi����x�c��~�o�8�b=u,~�S � ���QFə9.R�D�wx�V�ɫ9.���<�<^&��	'�	;p�=�����{��Z�{��n��Řg��f L���&k�I�<_��>����%
��8i=�=�3,Ur�fo�F�g����],����5yOhf�⎀���#� <� �V'�1Yb%d�R� �~+	�,ܗ@�V-�vA���ٗ�0�� �*�k߲]lĿ�R:�X�VP�B��A$� ¾S\fD@�.�yR6��> 	� ̳n�ǩ�� zꇿ)��o�Ic%B��IT��3y��F����f+�h Z���gd!�A�dŤ]I_��ߺ+z����(;�\�z8x���[>�!�|�~�e�����C:vo;��(2~��~J{Q��� ��X>ڗ:���On]��XՖ׮_K=�?mtc���/����������ܗ�ʺ�Rf�Y`�� ^I�G  җ5[��e�:m��Cc�2�?�×x���'�e�����C[��RvZ��
�iJA#�t�@s�~@�GI� hv�?Pn��j�>C9)���
�[�� �KI�D��]����@�x�7��=����~<�B�#��xOn�(c(#m�A]�kD��m��i3WP_|�k��%ڣiwʯ(�/o��أ�IO�C9��_<C?�2�&���C��[�8���\�r%�	������}R�0��@��hI��Z�EA � �o���||
�O�x�y���0+h��]�`�J��y.'�ȟ/)?��Y�=�)�A���,�ڿM�%�%�{%}I����c:�C��ҽI^!��V}��2i0�E��e4�k�o�� �-��J���$/�E��a��������6���&.L$+�8f�w��c�`���g�n�B6
��q��r1K����қ�Gr::�V�,��ɕz��ѭ��K�"?��ۺ���J�8L���y��2I�kq���s;��}{'-�|�م4	Y����Z �j1�����B�Q ���I(ױ�~�{�kݕ�l�䶊 ����M�ɥ��� `!��A����H!�K_�R��P�4������ UG�(_	�r	��^GdHx��B�=�\`~�<��T>� ����IhU�,��zN�Ԩ#�<���}X)�7 �K���O�@�/��5FV:�&��,��+.�\iK~�?yX����([V4�ٛm-�^�P�:?�;�8�� �� �
�����B�O���3ԝ���}�w�?>�a�O�,��3~˲I��]��?�I�N?��_��n���έ�hEXx�� ��ژ��7����7�=� �I��|蓌1�Dܣ�H�q@�xO�G��EٹGic[�n��-���?���/�՚�i���M�YVTꞺ����{�A�@?�]ȇ1%�_�?����$~�O[ǤIy�4���h¼'w}�Ń����\����칂b�rqO�ҧ��1J|�������'̐� e;h�t��^�e��d,2��Q[��}�S�-�[�Q���pT 6EZ�̴�r�k�KeMd�hS��L�ﭦ�(y��'쪙��\ؕ[7��|�� ��P�'<�����<�-���𨠯���f�%�A۠8�_<M������+�nXg�'��qڏ�~�v�Yk��gN)h����<��@S�KQ��	m���<<(W�~-n�E#P�9D�i������A%@o����n�i��6.��Q��!`�	���[��Q��ݥ���e�����UE�C�?ȷ�2�H�hq���\���m��ǥ���������=����D{��Oi��z� ���q6�$&��a���0�x-��ǻ*���d��4�Zܥ9Y)�y�.#��oHu�)�ܵ�/�&z~=<z����b:��YU8�@8T�q�Bc|���sa/�*�>���}�:OTnb��FC�i�p|���'z-�c4�y�s����YUR�<e��6] e� B�,B���%�ĸn!T �q���kr����\YI|��Ւ�*��m�����Q.z��l!��>n\������7'wR{��.K3�#44x���q ֥Ng�R��|#@�)@^n�r�%}�"]}�� ��y�)/d9&?�B�DP�_"�+������#�PG ��Zˊ�d�y�Rw�Ӱ_t環)��Gm��O���hb�O?�tx�qod�J���a��~S~���J�պ9R~��Q�\�x�b@
�.�~+����i#rMg¢�tR^�D��_�{�2�����v�b�h��y��	mŻ�-�0���Љ:��:^�H�@��'�I���Yꐱ
�L����]�%_�5uy�=ל��=Yw/_���2��l�d�>㖣� �
�F��/�W�4vc=P�:�6)o67R� XQ/�%7g�#�VSnU"��M���\�A>�cY�C`�y�jS���8Iq��z�Soʏg�h;)�&���(u�|@�Q��q��{�1�B���XTv);�+�C[RǤ������R�6 ]�&���Ns�u��V?{���bP��\�9����苾}�M4<����~k.�{8��/(
��V^}��`cԡ��l���@c��a�tZE�*­�=V�CxZƇ���5�*c��
�d)k�-GU�gv^�Z8��ӻ������C������ՃD+��]��J]�.CH㮝Sΰ_��v g��b�������F�r3����6��f\�'X������z�:�H����~���݃ð��u���dE��(��@4!~����"v��A:p)Ez��wF"Qo��n^�� _o��q��*@6�oD~�b�>�������DJ���,�T|�mV�.�����E�Te�M�y���_W�Ka��i� ��do�N�rSF��M�#e`�;� tL�pRL�X:p�xaPV(�f���<K�S�� � b����'_��r)��uҥ^�� XBy O�}�5V�C�X�x�g�o���;��A�x��)�%�G퇳�~��a�"_�2�K	)u�@L?�9:�^��|��z��%�p-e�����?j��,��|�.�?��j�^B�����3�K=V(����C��}Yۨ�#�WxF�ʨ ��g���!e��ְn�C��Uaq���rѷ��is�.e�ǂFIؖ����4�#훎e�Nȋt &���/S���+���_�������w��_�{�0ɇ4�O��G+�W���Us�N����@��Z�s���w�����_x���y;���w _� c�6�����S��g����c�~����FP�:�/бE�D�R����*.,��՞�L��@X�֒'�cȃ��M��|H�v�������3ڄ~M^̳� ZgM�>�ɋ^��K���2�S���w y�ԛ"?{0%eϨ�(�=ZJ*m��y)�J Qml=�P�_��|�]�����i��P는���)����F����u�B�4ֵ�"��?r���qO������S���g��@l���T�}�xϟWy����u��Je�Ͽ_z�$$��)��Gt�RlZ��>���Z~�<�ķ���Rz^	�W�C���`(�餖�������Y�Ϛ��WR�u)�:����j��̇�PoheQ7<��R �:~�@{H$惰��b����in����;����a��]�;�+�r����ڎ��$R�BFAq}�7���9_� �8s�oU�h����x���k O���i�qa�u�F��c�Cs��Z�����Go�H�I���J�K���9 ����j��-_�b��8��ל���ͻ\"`�]x6?FD�U�N�&�*V��~<�������}&R T��
��󼋰�`� ��G�<��<��ԅ�7��V`�K�΁�W�
��&��d_��LٴwӞ#�TW��ZVC(�m���ٴ��z^o,��!�C�H��{q�G*C�N�Q�����J���(8_Ku�UP�_I�2�>�#�y�=���HC���e}��;�J�����������6�D=�O�
 �U��T���3i��׵A�,IIa���G;F��-A�zuX `�Ժ�+-�`Y9�e����r�
h��d$�-.��� 0�>r�^}�2�(�H8 H��z�y�����JHZ
�E> ���9���#�2P�����qO�ѯ�3�^J����B��0#}���c��9 "�F�bJ�x�y�b�i��@A�l�y���� 5է<]�/+"|iϮ�xQ��?ˏ{; ���0P�P?�)�р`ޅw�˅_x�9�m@r���������@��
���E����<��e%k���8�M�Ѷ��'�	�EY��N ��-�=�H�S�8y�g�ğUjɻ���G^s��֒�N[�- ������J�D�E�4u]�pI��GmZF����׷q����q�ϣ/=�;�\"5wM�vjo�G��kB U��	ZOK�47�5��-�i�`��P�%�@�n��,�$����|�5Ov��R�)g�g����߫�� \5��pV!���X�p�N�M�� Ճ�q����#�8��Vr�$R�x2�GY��,8���Wk�5��%λ}*|��Ǣp})�?�~�}�f�WW�(t��W'��$��q��e4��6{�nD�歃d%��
�zr{��y;	߸�r��IpA�D�A C�І�d�3'�w���}M�}\ų�3���Ӑ�������"L �a�@`�� `</ (�� �\/���B>r��7麗����Ә��Q8���g?���*Kl-�7�VY�a��?�q�aa�!��k߶�a���-i><ϻ�b<*/��侀�y�.Fh
ͤ�����7u�3Tu^��,�/�qM.�Xv$�!���
�����>�/���p���R�k��(�o+<[+Q���C������G�
|F�����+����(�\��u;�|
�£���{�e��ZA�*3����G|ـ;}{$m]Z�"�Z��Ϳq�g|����{�c����J>��_���s %YN�(]_[o]�e�J��S��v�����4���k.��3���o����2��mF��f5�����j��3�eŤ���
L��y��h�><���	B(���gP)ڹ��X�t�~/ԩ�����8��^���z:���W��R���R"R�K�m��w�C��+�=妎���?�'<ۇyU�)�Jԟ�zS^Ə�Ǔ�׾��4gG�{ޟ�>{6�=ݎ��������b�OT>)EQ,P�ӥK���۳w)�R^YZ� ��ߒ�fO�p �A��l����W��w���m^��=����]�xO�%k�}f�u���ur!���{�N�On��z~�����@PW��_��'����+��uX�XyHw������Ί�r�t����O}���8�,�#�)��}|����u{=�U-\M?�g;� gov�����^�͞޴�wD��:�m����8�Momm���kam�R�<����������Q���"Cc!��5lmgK0^b��߃)֘�p��p��4|z-
P�82�f�ً@��"W	�mmr��d�˂R��ǒ�'�
 ��䳥��+i#L���6j�UU�����^�$u������$wO�Y�~,�s�<"���ŉSGs�D[7���5�V�-~,X�Ĥq3���w�FP��6�BE�C���<T�^r�~t��CJ(� z����Y��N�.r�J�Rm�U�>�	����6-S�^�[�oK� SWRL(xuhR0!��=	��O��6�ՖRX��
���[�Ɛ,����Ҥ�b�����v���0���r�]TdEI��B���u�ߍ�C
@&yP�<��Rf����G⣉@����V⾬t�X���ó���c� �Pc����s�zAy�u�	����<�j������<���(��Þ�l�E��>�ɥ��(8K������	^��}|Y[�u�;r�W�2� �����u#K1i�eYQ�i��>���oVB%����l����������y�:���'�LGL�e�m4�� ��W@�R��# ��S��������-0�i����O���O]e�A��k��]s4�k����lU���W+t-��:[�3J\���0,���I�iGx`���t�_�^R�x�n�]�f�՚Qʫ���:sZ����w�S_۟Y�/�������_�o?v���9����q��R��{��@��5�9�6VK`D�q��	��NXq���,�xo}#<u����O>�R�M«���}���λ����Z�w}}-�?�Ν�lą!k'���xk�RO��S�<ӻ����>�z#L�G�q�0�Ӑ4뀰����tD�N@�>��#d>��g��F3���A>�㝢��wܸOn6�m��u:���O>��������G�V�J����X�pa����u\���|�f���#y�!�b��o;	���?n*�L����>�!l��NH�| 6ʧ4��$6i+��)7A����l�W�ldʢg�u͂b��~5�l,K��_�]�*J9 ��s��Ӷ�}.��8����Qʥ}�JW��I}Z NmA�*Ye�Yp��#��ݣg�>@4�xQ@/> =�\��^A�#.��ĸ ����d�~�#���QO=�T��Z�)eA+hcA��Z��o6lD[���r<�g�\�=���)���o�����|Ξ],���̑���O�]B9m�����}�z%$/����a������?�Wc@��(жnlY��T&��C���u������@�:�1��� }RnI� ��g��5�xcQUtn;�ԓG���S;؈�60`�����s���k���.^���f=��������Z�=Ƭ�:nJ��4g��j�쓟���6���(~��$���l�y�̹�z�\^)e�I}���Y�6�{��/%0f�;���O�i�+]��oǴ��*���b�������n�w����e㼯����4���,�?D�q���PIizDq����S(��V������BY��c��?� �b���:z�v�KS5�D���%#=������O�g>w%\��D�qk�}�jx����{�A�Gao�z��q����v��}n3��n�ߏ<�A�#Q�:vvq}�`+
X��:.��A�A�8��
i����pc:��.��ᒵ}n�=�Bh�e����O�k7&�h�z� %׾ �f:[a�}j1 J����+�#��壣 tP�G��t�g{�j��@��L ��I�{%�'m�������F^x>GXŪ��#�R���CG��Q	UJ -	۪#x�Y�lQ>�'�Y)�\�K�X���Y��"ܒ�1e�0i�F���)����(*>�(�������B@� /�7��q�
R2О���-����F��Կ�ᴷ>�h�b#=������dy��I���^ڋ�{)�0����*>t���|ُ��Ϊ&}��z���Ƌ� ܾuۜ!�)M���~�����Ⱥn][���6Z�w'׻zަ+@./=kӰ�*��>���r3$]�s��R𮭤�r�~�5�jǀƳ��Y�M��U�����a�+�� ��\�8?r��d���mZz�ǥL x�n:h�.S����z��̕�2y�����@�X`�VyFiN�{���k�C0���Y�|�EױU��ҋ�D��3��ev,���m	*��?�btYw;�wU��>2�+ɹRk�JK}ƻb/�W�x�Iïa]�ܕ�2��x�J��gK�K���ٿu��7��=��>��zXs�����0�z�Ҫ�׮�'�cd�Q�z��xu[��P���<�R��jaڬ�^�i`�DH�`�_
�>�B�/��_�ֻ�����7�
�n^���`�v�Q �Ջ��f\�o'`;�[���5�
g�;JG3͒��(s���,�N����'��׮�{�E����Ih'
&�IxC��֙S�k�]�8�A��W_K&���w�}'	���0X &��P�b��0P�N�cVd�@�EC���P�ˢ�!�(% ۂ��н�h�?�y(�3ϓ&� &eH���f������,��*O�V���`��B:�W�L�J�Q!�׹��%�T�������R .qґrK�e����H��H��ԇ��_E����] 6rS�����v��BT��-�T$�4)�-u L�� u��*���~c��>^@2��R_�GM]S^�Β>ߊ�HQ�ʲ��k#�r��q$��W�Z�a �ʥ��Y�L#;qN���,���ZսuU?�]5��n��qמok����~�ׁ�JغXЄ�E@۾�����Z~ӟ_����/i���"��L����������*4�|��ߊ���k��W�Q��r�] ��o�x��	�u>�G��NR���r�KѸm�{t��7Tf�����c����\XT����%z/kȺ����MRF�c�wt6�������Қm��� Vv~󊝒h����6�x�.PJIbݾ����G�׎Y+����+fJB]�P����$T�}�iI ]<��C�)�Q��i �������P��}���Z�J�� w�[�%:~�D�=�����Y��P ��J���3C��zsT���9o�<�LA՗F�?T��z҂�#�.���ڵ�ŐL�u��fn8�詧�	/|���d�������W_+��Ȏ��X�QX�f@}X����:h�q�kq�g�s���Dp]�����4]� yՖ�+�t �\�`��R���TdU��e5�|��d_���݀��ͬ��� ����۩$�����O�&aS���0k�G��&p&WT���+�Lʹ���X�� ��"�Ճ�yJ(��<�<'K+?+�(_���"��o�#�B�Й��!��:�o�r���k����<V���X�Y>_Wm.wQ)H�G>��oC�f�tIK�R	�C{)��n��n��uiL]��Z+� �����I߂3�Oڈq  �S�:>L��|�*��r�J����\@��Ѧ�������+���C����:��|�u%��Z+XwYt�����c��u>/
��#�\�Y�ڿ������g�]�m�*���i].N���a׻�˭8��3��dS`7��Z'��<7lh��B��aqQ�e�J�4�Y�uF���9�:�(��Iˎޥ���qE@g-`]�1j(@tl})��n��S~>��b�PP,�HgA�--��`]�H����S#��{���j?�JAu�Y/���F�c�|t|��Y�qWV>6
����ٲqd���T'rL�@�/��v���[��)�<8^I����ީ
s��r�S?�-[�	���և��*�\�^W-]���*�/���<���P{�����:)�-���o�صt��Dg�>+�z�B���ԟ�&������������Z��P���R�B=�ىΞmV)A��.��Lu[ѣ[�Y�#�[������ҋ_{q���_�"��O" ���V�I�I�)�0}��Sk���\\�g����D<�U����qߪ�K�I��P�#��#���'?In��s�:�}xeᇬP9*re%��1�z��\���2Y�q�P�!��R�!�ɽ��b^�B����@��G�ڙ�;*l�UO.��C= �e��̓`zp�>�>V��zW�"l#�B�p��:�|$pC<C�Vk-������coHa^�]�L�ؙ��5���3�q��BN���&m�{R8��ԓ?��։���%ɂ�Ћ��o�/1�QY�s) ������ �|����.u��z�R|��'�� ��V��T�9�R,�8g�~l�ض��R��X�)���20��z�/������~3�m[!۶��Զ<5iYk�u������1�s[�kvA�.Җ7�7c����9Z��Ӿ���+��)7�R����^Q�ħz�
�& #E����ƍ�gun�<T����v3�`e�q���П�B��N9��5���γ�׹���D�-(���ˌ�0�"m���ҥ�)@�\�����t|P����&uOz��5���i����9��%c@��p�o(���<L�������R����G��@#	�FicǓMxD���/.�{�{@շt����Ӻ��%��Pa��u\*)���v{�ѣ�"p�|%����Wx^���8v�!�[\����SI�f�WH�j/Ջ��d=v����Kr�B}��д��$v��{����ï��]5����E���M�q��#Z6�{}J���QU廋&R6��Ѳh��_�6�/�_�E���.�d�^z����>��4Y/_{����믦��5�ㅹ)���z{fm��c�eR��3�}���c�8r����dɜqm�Y�@�rۆ��otX�;,�,��;��,�Ǉ���I���ÅIxkk;}䞬�S��!��
 a�<h��@�"M	��3���6��HǠH�Up	8�#�l���<���
a�^�ܥٗ�Ż|j�)�τ���y���:�D{���!�k��:G�P�������_��I?�Eוּ�jG���>Ҿnw�����f���
@� ʻX�li��6 㗿�Ujܤ	6E>(�LI3���i p���12'Ck[Bi�S]� G��%��x�>fޣ_f�G���bO��k�¦�K��kg�E����L�xk���ϭ˨U����|i\�g��(-h#�Y��h�G� ���q(�j��Rޖ�Ң�]5�5.U&��>&e��'e���g�e�y�*�le��1(�7���4?0�$�3�~ļ���藊p~�9��`O�,�ʗ�����NO�c��Gjӑ����Cs�Z1o�cO<yP�(luV���>�<����^(3�x��M���~��_�?�\�	�xi��
�W��{%˰����ߎm�g�y��ԅ�(�������
 {���sK��uO]e�@��sa����Y̧+�%Y���ɻ>�-Gvl��]`���5?Z����-��E��.pZzήh��|��J ��ﲶ�{�D}k��<Ϛ��l��pϔ�V��ۯ�v���ǽF���g����@������Q�6��*����=Q�Aŀ�a�c�@���-uQ����~.�_P��/~����(,|�ɧ�p�TXU7�Y�L`�8[G����(x=z��$��c�&U�^�o��'y��⽽��ٹ;��&�$ni��@��]�ٝ�wђ%��?�i�r�J�YT���0,�+�F�+�B�V���½����V:�xcs#��f�$��9��f��  ����c����dj��!�gy���0��/})	�X¨'�G8��c��ז�ԕ��j�'@�@:�!x*0��T�jʷ,_�O9$h�7�K��@�вi�Cҥ��Y�A�~�+�Q'�+��Zܷ�b�	Sw�,�оG�tH.�H���T7��O��j�N�eTQ�� �<G]�������8ξ��o'�y(�'u����i����[�:{������PY)X�������|�U�@�,���� !�G?�Q*;�,��{:ig�����&TI�� =g�&�k�����/Ph�K�_���+ �ⁿe��3��XǱ~6H+���q��cQVX 
i�����2/#ێ�c�
�k�1Y��N_U@=Ƶu�Թ��yc�
����W�W	�������JY~�ȯ�bH��z@a��qBߎ}�ʋWR_�ٹ;����F駹���2�/�@��@��[y�صI�r{/���/��+Q�����g���xDP.�:�A�:�H}�*E,��/�vN�����,���o}+)'�x�����i됏-�,|�h��J������.�t\*�v�Q�^^0.;�Un���N����kI��)�+~��j]�R����}�G�|ڭRv}R��\ik�d(�-a�Է�?]m�L!S�}�Ļ-��˔Q�.��v�<~4��I~Ϳ�d��zYRJ�ER
[��i�=C����� d X	�M4˅K�O'�oS)�B�;3B���=�@0�X��^{=��ƛagw/.����6߷�'�Ix��#m�#cΟ爆�IH`�k�k,�yO�9_6ʈr��A����3"�� �ܾ��X�_��[�IR�(do�}����3@@�dr�-6J��SwTZ�<p.�;�����SO��8nʵ�M���ZM8����.|�aLn��	 3�
�0�y�=#����h���C�IZ{�d�H��������J�?5y�7���G}k���R �𫽴rIV4g�xu�WC��H���ڹm|,�PDS��]�0����i�0�ߴ��g�y ���J��)�����c*փ�*�P/eG>��	WS����.�����,Y!�f*7rD�HB���h:�� �Oڒ<q��[�$��}�� 
 Z���"O~k��Lx�7��u�>M~���w���8e�����3�xO�?�����Ku/�q�.��&�S.k%�&@@���Q=M����;��s�gM�+ҐeM�@�)�(��M-sEcݞ�L�]T��^��;��B�o�e��<#�����붎W|j/;e���o��e�T?b�4|�@d^P%����K��<"��b��ʥH�RʳB�\�����:���.��Cj�x/��8�9��/~1�CY���׮k����<�	�.�Q��WJE�"O�]�߭0�s��v�����F���N0Pz%����\�8N�y�KiY��K ���%-���[��ci��Ζ߻�z*�U+d��Si]���|l>���_X٢o��i�բ���a��X��C �k������2@Y��n�7]
	�L�yD2��V�`�'���D�ښt����=�>[-�!:�U:'����d�u�a�0������D������阡�^���~��ߦ����~�q�V���*�<�8c��أ�������sX7աy����>�0�Y�����t��N-�����#?
��~�l
�K�4YYp��G��'a�g?�i��6��\��dU����i����uja0m�������/s���Lc�F�@�<�5 �ʢ.�"#�3�
��Ҋ�,!�o	�Xd�7�e3)��#E����rP��T�h��"\�X =Ey�b�=���e���$�Œ�ɗ�B8��3t��(��-�Lj[�a�Ad�R��_��������H�$@D�TP�����Xkń�9��<#WP�hb-o�y�ł����CZ�HY�}Y�W �<e������4�ƾ�*q&v���y/�/E�T�,��������GxF�Wg���ϴ'�9��]�@��.u�=@���� �����	dQ�<O;I�3�m	�� |�,i��?�C�U�@��Q����H��0��# 5���Hq�����4Q>@�jO��H��	ս�"�2�e�M�og7Yn)��((�ܟ�LU^�ZǤ���2g1?��<(+iI�!e_�{�oXΥPa.�x��K9�M��3_'��A�������=�e��N��M��XǸ����?ܮ��_�5��;o��}?܎kJ(�x��x������/��f��,ڿ������n�r�����A��Xk��f}Q=��D��_�UN���?H!�~d=��:�5�����D����;C�̕k����+ӽ�������n�a^�
��0�p2�4
W��б��o��%k�0٥ظ[���!��+PJ X'0?��:FU�C��=�;G�pC=�#Ϥ�?��͍laLB��GҢ�֛o��_{=\�v#��'��{w3t���~ Xr��C�'ι=<84�7�a�]�����4�#-�,��8�"R��rs#l^��������:9���f�#  �&7h��v��S��W���	�
$-�΋8��f@�E}�����W�'m=���Oe�E�HG�D���oYO���o�]�[{���i#��]Y�$TK��p��:#VQK����Ϛ�|�畯u��Ed�G2�Z���	��bB���ӥԄ*�z���s����FN�z4Ey��UϺ څ��Կ��R �׺��,�!L��@�ƭ���2i�]���X�Ir��u}�Fڳo�ӻ		���&t�QF�K�B��#�J�:�Y���c�H[�Q��Q�R(�F�G� �#�W���,�����ڌvXҘT�6�%J7�e�d�g�al**0�(%��$��Ã��ʡ�j��S�������n�蓅[��
����87����pO���e��� �*�b �m�oI)F_b~�\���6&�~�<{�� �����i\Q�|�Ma���gU�}�V���IZӪ�<Ea�����E���Ǳ�>
��>��{�H�:F�1���y�B��_KԯjQ����JC¢�</E�]�T��cP��U�Y��m��bShζs��Zi$E٦-�ϒ��2Py�ԺqvTu��?����9�K6L�ӳ��E�֑�>�gG�]�`}*���]���r�On(��ū�[����H��f�q�9B=R�A��f˳l�죔F�t��q��, `��`�`��<yx�{ ���i�7���w��ҳ�I��m��>XW�L���[���O?�L�u�V���çGװB�#P�H�xom}�R��=L�G�gD����f+�l4pyf��(�;^��;-�⚿'�K�����,\��bZ8�p���s�������&I��1C\��n�
-�AH�-�5B��{�׍+���S��F��9�����]�3:�R�gN,�p���	��Ig��,��79��A����Z��³�z�B�Br����	�%`"dq��,
,\�ϑ�Gh�\rOԞbݚo�W�X��ܕ�kY����}v����Ĩ��n��XeB�������r.k�ʫ�� H��3���v�@� �����F�\�~Aձ.�O@Y�H1"�ؐ�al���Β� O߇,��7�����嶞,x�^<W������7��4�q;mޱ�Ӵ���W�>�~L��>[�N}�j�!�k�m0��H�v|J�P�<)ФdS��I[/��i��ʫ������֊����͂���s��J�T?̫�Y;k����ʍY�]m,���q�+�n 2�u@l��oD ��al��8Ni�F�:I����^�+(��~�-�?|��8�0O۽�⣋���mc"HAj�9B�ׯ>��P�*�K)R4��^��8,)G�����nw7�]��Nu^�Rݥ����׽M���m�p�(��=���}�N�GC��d(��"�؂P�]������3�^hG)+lz%��y�Jמ�`���?�inb 7!_��_�Z���I��v>���R>^��E]<�
��z��t佪9b��R��^ ���/S�t)�������v[m�R��"ڶA��y��	C��I�p�i�,3���5D�y��{߮!Ch  v��Ց��T�JYE ��J.r�$A魷�l`�H�UD�nn��}�x4?��Si��4}�i\Z�UZ�'y�/��$F#Ŏ��Ѫ�6�'��ētcgg7�;{�m����&[Z��}y��-O�����b-uTu���"ZM�(̅C�9g��������Cʾ���쇅_����k�h?� rp��������R/(�F����G�H�eu���ON��!	u�J���þ癉�,Wi�����w�����5+ wiB����[����d�	��1�`�n�:Qy,`e�  a���-�ј�YZ�l�z+q��,p��>�4��U��|��pڼ��?�Ѿ;W����\j'pJ� ���?e�'��4���OR�X!�֓��g�MG}��i�s�-��dܑ��ֳʯ�k������+
�8�} .T�xV�
D��0������ڲ��@�I	��3RlxŊWnA�8�؟�W�����9Y�G^1���my���V� o��� �֭��5@���Z�RT'�1K@$���G�}��Ó�n֍b������ �g+X��yt~�.�Y�lP+Ճ�Ԯ6�oK�j]=���k�����QS���~���i�
=����1k=���m?^6��9L���Ǝ��v���}����<�t�{���;U���z9nk 5}n� e�[���s>�`�k� ׏{_g�k~��u�>���}_�}�X��E�T>�Cϕ+WR���|��I��9��3=��*Ճ_=}<.�����A�2�{���x()5 ;~���_R �d:^���}܎�.c�2��$T�����_����o��ߪ�t�}4 ��P;8g�DWu�9�����v�/^ �Ux�ͷ�o����5��5(k���w�k���>���������	0�`GYF�_<r��dn|��ﬞ�G�!�d�$!i#��{�֍4	��yp0���G�%[$�|�����P��W�l7KƴPDU&�1����FY|pپ~�F��nG �~i�lk_ `Qt��
.�� �E�Ac%�c�E�I����\i�/�Sp�=i)2��S�v�� �z����Ϭ�#vd����sr�E�&X���}Ȳ�@ʓ��9	J�ɯ�k�x+�Yˑ�8K��h�����`�*Y���g�]�GIP�J
	d���7��?���$���-�޳{�O�
�%�U"/P��xk�U�@RJ�=\���jW���,bJ�.Xj
~��F͑R�Y�m�[���.�-pU�؀B�����mA��G�)�b��s�O��A L���x�}˂8��a]��3^AR"�,ň޷m���q0O������_o�<yA5�dN\h�3#-~y]N�)ϨqM�F)�d�V���6�wj?x�d(ŵ�vn��t
��:ט^P��z�}��v>��1�[`�F��"z�v�Rv��`r��kǫx����%�x��N�G�M����G����{t�Mu`��3�c�uc!h��@�����t%I�u�c%�Jh�VNQ�`Q�ʗ9��L���p��Ұ놭W{ͻ�۾k�ڦ�缲E.�2 _~���o��x�?�4J�o_9W�]u��t)|�O��i�i�*��km��1
���Hq����n�,[CN����l^�T��3-��
W����N`�rM,�k���G�@npk�� �d\w�x�ɴ���nni�IQ�q�^�G#!\��w��c�Z嶓��L����I��s�+��p�g�R����7 ���?L`�(��1�/%-KP�45ɯ:�B^��O��Y���|��V��,h�/�_J�1����վ5����=E̴��]�+6���QAzx��\S�XY2�F]{�$8��/w�`Xԩ�G���V8���w���j��V�e��,��`Yf]@�{~o��{�|$��rB���O�)`���?dr��{����w=q�te��h����y ����s�|�^��� �lr��)�To�U��%��v�ԸY+����w7�}��0g0v��2{����[�|yJB��X��W�*�W�+��W^HH�ɳ�;�2�y���n���ۋ�J�QǦ�u^�ж��c֔W�7����d��y�l-J[rҘ���hc=y)ፔ��k�e��w���Ҡ�P?�J�S�i<٭&�j���� �����s�+�~�Ks��;�4�|�X�&Ő�x͕����k�s�\�e=��ӕ�*!��r��]��6��0k�Y[�oG�]u�����w�s����swi)�s�U�(ϗm�la@����b�`�qM�7Z����iZ6�k\�Lq8�N'CD�}gw'నd���Y՗����SRv��#��߲���Y�C+����%��tV��
�����Vsu���XryF�Gs�3�`��Ydƍ�Ur}6�ܚ�;�we p���]�	���2�ٝ
�\�?x��d�z���Oeʮ_�!���k)�&�A� � 0
��OBv (r*����O,��%��b�a
��G�+�4�XDh����Au6&yʲ,@-wEE<��$���С�_����B��)�"͒6i���@�K.��f!+���)?���Q��4��>\/���.�|�tOu�`�w��#���0�<�qD�e��庬wd�8��D!�X"t,O�
�xk%�B����e ����+]�J�[ʔ�����/O�$E��DZ�̺\�o��^1Ҋ�u�� �R�4S�Uz��>��	K�}��X{�5K_���U��Q��j��5S�:o��?�q��s��G�'�';�;.�� poiV���K%�_�Z\d՗w��)Z���%��{?] ػ؞ w�_Rh�����9�慦{�}Z�h�U~C��]�2N{{/�*�qY��r�N��3n�E��22�]�d�qߘ�ϗ��V�恫W`��_���m#�ζ�O��1Hp�:m!��B��Ҽf�����J�A�{��$��nǭ��X��
�Y�H2���Ev\�)=N������! �өକ��WXr/]��\e?� �ʛ����S5��K1`
�9��WP�1�=G�{M_Y}@̾���Fj�tH�Wӈ�D8K�"���p>��X����dq������X�H@+E�e�~\!�&�O�&Lܔ;l��ג�lf�a�҂m{��v�3�H�7<�g��_LiP'�X��Fj�ZS�Z��}���H[N-օT�O��p��J�k�"����� �U~KK( �69��K��Уcx�I�kۢ��2�P|��/�U�@ˀJ �=k�,�O+��*������������m]E���޳�lz�J�j-斬u�$�yp[��1�U&��c+,�v����6�ś
�O	ۺ-�;]�蓺S55 �Y���T��5�c�[ "�K���ReK!�̵O=�Lx���Ӈ��G,�KJ"0��) `�m��]Kl��G XQ��X��-��, �^-� '7��t,���
}���+���6c�^�F��ȺQ�H.2@��"���k�zNS��ߗ�4��GR��Z}M�ޘ�<�O{�R�KOy��UO�����{v��s�'/��k6��R�W���\���2Ӗ�R��G�?�7s�2���i��2��e�,���j}�W��'���J9�S��n%��]{>���(�g�T��3{v�ߓsm��xd���&=��M
�1�b����L�ơ&M�)�>��_������p�E��� ��F#�B����I�h\���b
�@�4�jo)[��"�e�Hr
�Ϥ��o|�$ԥ5U:v�u?+8ZAU���UmF}]���%��[��J��=˟�خ`C�W@�K[��lI��AP� ա(l���Ug��U_6>� D$(���P�����s�F7\uR�#?���<-JBQxoNi��>`n\ ,���w)�����*�U�Y�<s����Ƭ:U_���EϻPK�����%MA�s������wOo�Yx��JV<�6�Q���4@��������n�s~���acs+���׾����/��� ���q�U`�O��s��N�Lr�� ����ȱ��
�e�ֳE <���DSjh-��'}��P��ٖ{�ƃ_����+��Y�xݥs��K�Y�1� ~�F�b�o�7j��,�W)k�u䩍R_k�I_�b:ߛ�ʶ����gh����z����m�%��=)[ �R����.&�6���8�Κ��3 �!����z��-�,����6p���5V1]����� �����1T�
���w=Ӆ!����)[���9�0�]�o6��j���Β�G�T���ܡY��Ux��p�1m�fv�.�N�9��l����Gõn9���r�M��b����B���3�k�����pW%��c%e�ha'm\)|DӒf#dB%�_;�w�T
fc�:g����='I���v ���bSҺ{ AHiX����
�v�=r��T�6
���R^���@O���|��M�<�^?¯��A�%R�Xw���*d����ӳ9�x��u=�}��u���gA��+=-� ۾a�� �N��{6r�?v���~�Q	`���oE?�����.m��xX������t�+�z�#g�T��tn�M�_VަO� ��&��+�Vr������SO>���Ū�|�����< [ �`V���#`���m�+`���p��v~��� ;��x��]c��J��ď����Wx�Q��(�l��&PU�*�8��:�>:0�̼ ���G�ٚ�u2,�>�|fi���s/��H�/c�J��������Y���~�4����ռ+o>�%�{�O�������E���� �%ZqZJr�I���R�/�J}ϟE_>�4O ��k�:gyRm�]-L
�����8��d���$�s#L%�m<2`E:\�`x4�X �a���I���Iz�h�#�i��t�r�x�j��؊ϬG~r�I���5$�[vgȁ�H��jHV������ꫯ�O>�$����o��Fx��/�Z�e�%l�	ks��hT�ȕ�ҷ镨t܄xU^�jm�o��R	 X���h���w���4Q�4m������|˗��B � �fQ��R�z�H�S�-�2Y�ǝ�}�8^��;~m~����7��r�ki,y����q`��=:l$r?�}��r����+��x2^ X����?�X ��޼�]�/��!��&�)T���J'1�F�3z�/j
N8�>L ��|��(��j�͂�T����I�?�O��7�|#���?L��r=���Ȼ/{��}�z���.�V!c�+��@��K���u ��v��X� ����/��*�!{RF��*Z�:��ԯR P����1>���3)Yrp�Toc�gV`�r�Z��*X�}Zu�Z6�y�*�m���m�k��j�.�}��˶9f�f��;A��l�/�wҢb��AX���R�����Ӿ��'˛]���Ji�>v���ԥ�Yy���� �܍� ���O^����K9FB^bgM#jЄ�)Z׺4!�{�67g���9��	z5w}n�G�+7����ڿ.e���|.���v;������N�I�5m��%o&`j;��G8i'��b��~���(��}g( .M�v�X�������k�Li.X�fu�y�I��%PO��Be|t����6�����=���g�5�-�n����U�NR^H�㙁q���ϟ�� ��Vs|B��k=n�E/,�(��R����R=�ŗ�% �r/��V��g;�u� ���RYm�vL[E
J�>��^�`ǰ��iA�[�,?�*σ�FIK<
�i���(s�G�qM���u�Xk��$ ��F��L8F�B^Gs�
+�j3�Ku��Ђe�M�`\j�l���1& ��F��^,�?;�]
?�m�X�S����8�%ZgAC>�Ki�XPTr���X ,^�X��͏�>�����BK�C6�C���8�O�S��5��nd"Ev��2eȍ���a�р~�{�t��њ��'�0�b$٭q�N�^J~���8Ʉ37�t��е{Y�*�j��������������Y����Vyc]���~ԧ<"��ݾ��KF*��Wv_��ï�����܅,;
��i�����|]���K�L�)1_T��#W��t p3ɭ�m��s��1HLt鸞��p�歬��F�O���	�{3#�4�Z9�s^�ۏ@� WVةB�~l&wrn:fv���*~�j��u:jHܝ�yK*٧��-	W:���{��H� L�]ь��mb+@�Mj^P,�/�r����AS�2*/�[@��|~6�. ��g�_{m%�F5W]��'Yv�����ǚ�(�J X��U��&O)m��+D���Q,<\�C��(��B����F�ْ���.�6� ��,�~,��+ϐ�Y������(�����R�f:��O��	���pa~���,f�Q���4m�Aٕ��D����
��l/
Pa׷��(��>]����E���L�p�ƭX��~��\\��knՀ`��[��ڂ�l��$�����Z���޳�q$I���R��J����̚�g�s���s����?p��1=۾��7�n��0�J���JU��F��Df"M�a�܀2���r� `��K��F�����:��0I��5� �₠�P@��B �eH}�,�@]ޘ*2W|�H�0��eȎk���� �oV�bAd����Á�ϖ9�X��+�:�4��h6xL�Iohp�?���!��z��i���"�w���\�4:t�Z�cjLO�5/�qy&�?n��/��`Z�Ǵ[�vO����0Z�ᮻ����]�������oϙeϸ*���ua��M��z�R�"}�`�բϞT�Ĳ��i�^<m]���@E.Z V	��s�$�@@(�^_f�T�3�ěj8��(U����7|!��d{lR�q������$����� ��wee������%���q"a��ڰ���m@]�>�a=�Z�}K�S�"���}�����q��I��	�E|�*
߱&��)��i_�I���Ѐ!Ś�!i.���[2}�����Mڈ�7p>��Js6�&1��T��P�V1{U���괺V3 ���e��d�b}�txpJ��80��E�8(��dM���j������ݚ[��Iz��l�s�뢢MF5�L�~%��`��_��k?����Y������V#m�A�cnS⺛���a�l���B��o�c��[�T3<ЖY7봵��cc}Ռ�
�@,�1�R��7c�Oh����m��:T6϶����ij-����j��(`�Du� ��K��q���\U4HЂ����	��� �I��Kc>��_'��I���H�w讏b�����w�{]��,�O�賋��x�4&��ǅ� �Ų�n���fj�<��+T�����9&�dC��=�꾔�� ��ҠY�$������v1���Si�� l /<�Z���ԧL��@"��#/���9G�>=;���i�%-	t�7�%-��)Yg�@����
� ����8F$�1�e��2b��xا��eH66����:ݻ�Mw�m�c�67W�^�P ��QFp���}z�Dϟ��~|N/_� |L�V��u6������5iW
�Efs��#��$i�G���s���>M����y)
�G��Z���ˠe�@�\b�>�f�.ɰ��7N�P�͸�Vw�1�5V*t��}��zp�|_���5��  .3�Cl]�nH�Gg���������g����h��Q�}�<c��w,_�<�0�Ƭ����������.�hm�0�. ���&�Rk��q�,=��JK��]Pt|��y#�p��\����[������ �
���M"�;��*��Uvȹ�1tI���:�C���;q��1�fϪ�s�i��Ӏ��`��Kn3�W�_�F��D*b%���E �^2�-�����ڴ���H�6���0�h�حT�n�P�@#	2�����eP����z��)��1�>e ����,�&P�	��ITD���O�d�6�,Mo!�{�������8 d������10�Ӑ]t���՗���g��w���ݤ��k��V7{�BD	�(�U�v��{�n�K�V�m��n���)��w؊�`9�,�9�AT� 	�U��Ve�K�%g�����ֺ@�t݅�����h���.�V�ն�)�|a�<�������a9�Z�B;�����C�=�k��}ڻw��6��Zc3h�1v+ ר��5�e���Z���?����C:9=�N�k�L%ߥ�6�.Nc���2��,KK�ߡ���ιefթȵ7���Ŭpǫ��ehA�+|��t�:H�v�G����#w�'4������?������(_���\m���d� ���(w���o҄
 �?W���$(Mu���oi��u{
��=��^td͒b|�̶N��0% �16���2
�Z���a���c��E�&�i�� ]��oIKZ�dψ��[-�W�" F� ��U�+H7��vis-0 c�~��m��������f�5{U�B����4�G����2���5eVWig�z��6=}�O�����קt��ª��2��lmp*XH̴�P�o��i'fYK�}˵x$� ٠c�A�W�J�~L�v�*�
��٠�~��������gwiu~�1���˧�k�iЍ�8-f��u��e���z�^�v������=|x�������'���[v�~�f�|����#_9�o�S�@�4[���Js�j��y����-Y��-󦑫�Sz!�$.������")�YZF��>NĒ$�y��\~�ޱ����eUMӇ���� �`>s$����A4�`+͎�3 ���Y��-B�(�A0*���"�/�%Q�JS M��"�U�l'��D����-)�>�I�%�\Ғ�ts��$����B�ԟ
�#h~#Z])�έu�����w߀�]z�p��5D�X��aǺ�$���t���kՀ�T�������j��)�ӠQ�c�Lb_�P�jM�5����B+�%.��a�t��|�{]̀�,�KxW{�6�.�{�R��I��x��7{�}ã����!g1� �c��o�~D�������]�����sa����MA��{lZ`�̹�±W��&՚k��Z�j�������s�r|�2�(N���]�b��@��h�q�>Ԕ�K:`���M�}����y}�k�y�_p��{g�Ez�h!�&ɧ�ts���������&%��]E�o�� �F	H�X̡A�� ��w�[����g)�ǿX�f]盓E5�Y�fѤ��d]P���<�،���t}RX��Y����@���Y���]d-�� 8��lTg��#0�XE�&��$y����a���ms��Ҫ%-iIKZ��%�8�c0���:���>R��X�:��"j4���ޠ�?�C�����~��]�Xp=6�.|1{tKHY����"�RRN���(H�MQ��<��`svb ���^��I�jL2�Ш~�>�~v�´����3��"���1��Y�ɧ���eM*[���2��N��y��m���P%���HgU
#�\[�/>@�������#�ڨ��sn��#3/��7x��JA��O�C�)��S��������N/e������Uҁ��o*�jд(�E��{�����ߡ�����ty.���h�GGG�	KH���!�+}�,kN��5(,H��^X��]M�K?U�v,L���;w�������'~+9��}�����y{���9�
��Ol�����r�|^J-�Rë�:u���2L ����i���?iY+m��D�ŝ�=p@���8N��O�������!rl�'﹙(Jv�8�`��榏[����L�¥{�bs��_k�&\�0�K��idՓ}$�n��-�s4v.�D *����Ƒ�CՄ���kD��f�I�ݢ�~�G�|}�=X�hpl l�������
�Y�ao��ÁA�Up��ڻ�I�����Cz����N[l� :�бP8��2Ղ95��Q�\���_>-���R��i��ߊ<kr��n������g���</@�$��g5?e��zZ]����m���=���=����uOi883eu��At![Յ`�lNj�#�e�*15�5���N����b3��R�oSV�t��6jͣn�,LvV����X�E�κ���3s��|nӀ�E�;vu}�D����� � �ȱ���n��`��P�9��_�VT>Q�<�^�r�L1 �x�d���,)���I�ϧ���F�;�����Y�����yB�ܿp ��1?
�"��/����� �D3<��$�@W6:4��;�G�D��	��~�X��m&a�� �vK���ȍ�,֕J��R��vA8�n�K�L��C�@s&�H��i�M_|�j">I
\-Vq0Y���?9`�%c����=i�,��/��)��?��t��L�?�a�� o��H@Z��J=Ֆ��k�&U�����y���c���L|��}~ҭ�&ժ�D}��j�Dǰ0�+K��<�q����kg0ܥ�f����>]�cz��]ƶ�	8o�e�7�Ѐ^��)u�\�r�B���H��`є������=i�Җ�ed�^�&O諫�=.��˩<���K��o�-�`�ڥa�g@�:=z|�>�����e��1�'f,v+6`k73,(�X��@�(/c���+�Z
��/�X9���S�7o����C���t{���G����f�n�i��v�uǪ���ɗ#�-�=\�-Q�u@X���H���vJk�� W��4��޽���:<<d���.�_�u��r��
��/ 5 n���uL��`�0���M�s�J�w�g��.��>v�	��Ȭ�����L��N^�⣅`>1�@#E;�����.Dp����03n�;<^0�����CQ���$��z���R�&@�����˷�� 5@����#Q̃Q���RgH�..��џ �J�j
�D�-6�.�E47�&����� {>��Zȗt��2�I��D	����د1��=�$.��'�d;�E�+���?�OrKbj�s����eZ_���{;�wg�u\�5���y����F�t4m�g8C�5]CJ�Z�ĩk*��l��!�0�[�+t��ݻ�E�g����;}6���|����5�<'c�]{�PÔW�{�[�,m�.;H�iB�m�4ZA7��%�e��9$�����2�� < �[]i������6cמ��3�*��v�?����//��xQ�U���UA4�$#�g��6�t�vv��ހ��nӋ��tx�6c��>m^pӾH*"\q���mR�\3��0V�Ã���3 _ ah|�;���b���q��} ا ,��R7��7`��<�pB����X���e|h��z��-�N\a����Y�d=�7^}_��,Z�B�FN4�
���tA��e6�1��4�����F$4�׊$0T�\�א|�ؔ+d�-��%�;���8���4���O�^L���39}�����x�|y�R/Lx� �h{���MfIKZҒ�t�I��4������mр;N����-8A
�����!�=��-�{ך4�-0����[���1���\ZՀ��f�nm�r��F�0��=��o�3�Us>d����)�?����S
�+��c�v��z����P��d��2���|�����t�V��\��"m��w}��4��z��U|}���X	Q2�����0 [������da�W��a�� �����tmz���~z���E}k+u�X����*��ޤ��:��y\�B��f�B�[�|�6c�m���И����<��W�.5X���^���W]G}N_'�������E��9�������7o�x��5�͚�j����R���T�y�g!�R64ˢ���� V��O�>���wvw��ݻt��}ú^y�7���kk��w��JLٳ̣���E�Q��i-$��4���TFL�11�q��DKh�0ghb1���6g�i�_J��:XA� �٘���������������9á�x�������0-�{��IĹQk�f���� �x�-@�<4���Y��P����H��tI�^�ּ8����x�r�g0˂���gY�/'�3������f���j��R�����b��ط����('��g]���m�V̾�(ҫ�Q�Q�"��1�>�j!mm#����S{9^�!����h7��|OY�
���E[{�.�/�j� ��[ֳ�Y��,v���,AB����ި���A�z�y� Zߨ���[t��mn5)t9XZ��Ȇa>������cz���N�zf̴ o����ȌM��רT+q$�th#�7�e�7��5�4H)9@_�ô�)����|��M�-�w�jh-�p>����pj���D�cC@Ήo/x_�:�}��?��B�1~Vq@����J�$�^k�4E>!��!��0�HL�%�.����c��A�� �����YWM�B&�|F=������q{I'��h�}�^���<�����]( �@��dM����,������2̣E�@�9��r2�P>$�I���H���b����O#�c���k{O�Ox⟞���k~�U�,ڐ�#�����v,�+* q�L��^#MkZ��c�{���"��\�[I��:w�:�aN�[.����0�HN�u���_�}N�W5റR��&�º�k���6��< ���O���S:kG�A�� �>�[�Tk�� �r���@��J��i����\7��M=��ʊ�E�$�3@f�0�+���s$��=(֏����EhS��sU�x��i�����ݾ}�>|�uО�a�
 <����i�W_?�{{;f��P��̌���[eDͼˋ��zuB�^���iD��:2��O�6"��is�M�z��fp�ÀM��� 2`�D; om�Q�Z�t�_q_�_%s~�Iƅ�y����i[��W�^ѳg�������@�(��<�՚E�i��]��|��D3-��^�����|�_|A{{{��:P���y����7�4?Mۏ�x8��%"���m~7I�M
����a�otRİ�J87IT�1���a� 
"� ���3� 1�Agk6�#I'i�k?Q�ãC:<�O"۵�'�NI�+� � ôe�$��O��r �Ou���$Ӕk@_şJC������ȻΦ�>q*F��%��	2o/H��<`�<1K��� D����1�9J6h#��0_ܐ��؀�.���tX�~��R�)u��MGg��Q��WRb#Hc���٢G�*��u:=��a�S�LBc���ݻ�X^M5CZS��1�2�y�W��wmQ�j��zFZ���.K3�`�&�Y��o�<x���P ��z�� ��Չ������m�7�`�	h8�V�0896 ���vݒ��B���c�:�w͘���*�i�|��a SVX14�O8NMRG��m��Ǻ�Mgƚ���#n�+m֫�������<�kvrMK��<�n��P��|��M�lJxw� Mh}�ʻp{I����W�־�t����R/h��!� ��	��!i�v��$�2?�z�;�t�7�(3���z=��]��"��i:�,������I����ω�s�ɂg���ٺh�����mm��[e?#��/7J�ۿ���7�����c>av���vL�H;�����_,��?+6�{��)
f �,IN4|�z�_o�%-iZ���!��;ڹL,�M'�d����'��o& �� ����C��/�� ؽ�Z�a�o~hs��T h�¸���0&HmS��Z6x��B�P""�ٯ��>���\��}��Q �{Y��?آ��*=��D�~�`�X ��+���=z��}�q�M�%@i8�5o�MS��e�Y��\&P�к�f1`>k8�|��@M��q�V0�_~�%ݻ{�c��­�f��zf,E�\hs�l����y��>��	.^���f@S�ZPe�(�{��=f,�����X	0�$̶��������Va��6�cR�W�`k�%�<�����~�&
�������[����$����A���	���f�/ 0�3xvX7�J�!���۫M��R�����Bn�%h��ݻ�@���`M0���[�X�0��7YAU�i�Td���^zn�rn�=�:���\5M�Y�p�� I> 0&¨�*�6�W�զÃC�u�˕Q����,ʰ��s����VlC��#NZ�(Y�)�r0���$E^h�8y�s�,��D# �`��Nq����/'L&l0�X q�G � \��K�Y4iQ�=��p��u3��b}!�Th�c�@ĥ�[�J~h�v�,R�ϯ�&�l����'KL��iI��}��Z4X��E�Ba� `����)J�-��q�i��k~��a�ׄooٜ�%��y#��Ṟ�Je�W,�l���˦�[@�Z0��QX2�}\��!`h�a�%��.��'eϥ��ӧl�NQ �5� ��u��Y�f���e�Ou�zJZJd��o'��B#��.���
5{U�{e`S?�	_�!M‭������Ps%�2c���V�a�0�s�hdǀ�<���\��LN;�E�A=�t畫�����Hc���r\͙��Xe]�����PR3�����Д�B��[Rqw�����f��w~��s���upG;%چk����"��y�H�E�W�|�22״����=��^��!��Y�����7�6K�@��?�_~����X�L�T%jw�f���+��[��!G��TZƉܱ�����xD[�L9�.���8��m=J5�p���l6�$� �o�Dy���x���rqqN6(��/@2���br[S�&=��'�<�ZҒn�69?]A|w�A ��_�(�7�j�@U�K��P �یt�F9�>&OK���f�]��W��MvF�?�pG���&�;���h��#����K�Ǳ|�W��0o�H�gX�:� WaP����׋�E �>k�{lT����V�5�sg��Û��&�lJ��==�F�5���;���tp� \uJM����������_�J�ww�J"��L�4�m�����'o�մ��D��J��PG��Y3�YeN���> r���?��O/^��v��+�������g;���>�?�ӗ��SMy�R���l'����{�٥�v�y�
��ȩ����(Q�Y&�%J�!��=:>;����"�η��{��ɟp�C�,p�7�H�>`�/��3bgs�6ס�u��K<W���ĸ��_�Jϟ?gh���
(w0�d���r���Y��i�֮k�=>����@��s�6��7����&���ԥ�`BG �~K�K�\�����ӂae����t� X* I̈��ۻ�t|rF�Ng�q�d>$����sh\_���r�dN$i�pG6eG��xY����H{w�n0���q$Rhp�����S::<2�4a�7:�Z��l�F�����M�w����Z�%-�CQ��_�5�XO8�+$��$O�m�K��&����_��E��!��$�MH�,�bb@���"76c6o9��x�%LL�06ք�F��Ѿ8�^D<z��H���
\��=�/��K'�v��7���������eޗ�h����f���yg���E�΀�F���+柝[+���j��pJ?�%� gf�zm�~�������?���S���1���f��˯��&���=hzS��ߋh��c�e���8y�n��Q��Ε"mv�%���|?��3����t~zf@l�M��sj�V(�6�vh��:�Զ�dx"�ā��\�iU9Bx�QoxJ��V���Ӫ�����z�sVC��k	�3 S_�;�6���@_�(�vFd]ۦZ���5&�Wx�^����rN�%�NL���Tt���5P0 ~���@�+�9�[�[�<�=wN�Z�;��r �D�-m����h�&X�ln�M��"�S��B��,�J��x�� �g���I���`>0 t�X����`f����9$�㷄hʽ./�`X1H6����lǇ��, ��ɵ�D�Cv���t��Y�0����b	�@���{z���M��G���C

@i>�_ }�\��[�=[8�%-�i���H�f!^�`���V:�|�1prʀ�?��0��Q9D�Mx�ph�c}�p�V�t���\`aаf�fN�V6�qr54�R�V{Lt�®�$d+��f'��(���u�\��&�ǔ7vbϧ��  �1��0�`�����|�Ak��Ck���p���y�h�ꆹk�=�4H�G�Z��f�no��=��� W�~�4{V�/�i���k��R����LX�#��м��O�7��`�r���ç%s��Yp���9!X��1b	�n�a�k	����z��-m��h�qT�m�aU��j��o�f֜z�NO;<]4ks�F;��}k��=��1���K�6V��a��]��B���}`e=��7�΢q���ܟ4��`@����1.����/�O����d�S�����y$ʳ�w^u��j������m����~������=�EW�E��B��3�n�;F�x����n�2���p��?+Wq]�	4�����O"*����Y�����>�nwY��v��Mh^W$�`)�X���^V��r�Ȍ:�}�C�4X?) �C���/��� �p�Dkl#?��-��������I��F0,���KZ �T�8�����j.`�M���7�Fl����k�Y�9���ئ���zww�H�!t�m���uL����f����>'�$P0�Nl�M%���B:�K����G��%�3!�ɸd@��a\[�� �{�Ը�|�u,�1'H���Nm��*U�%:ouy
�Lz�Q�u`Ve��������L�֐��Z��݉y�	u;-������}��`X��,���M�^�d֝�Yg��T�&=-a�	�V�?¢w����;��U���T�#�U�����;I��j�L�=�ժ0o�i}���ϥ2b�؊��*�:��2��w���Szp�� ߧ��n{��jq#�^%iM�O��
7�����z��@����GL[!,�>�4A���;4��?�'�
�7��)B�݈�/�G�b���v�~����@���"�t���W��z^���.���r>���"�(��Zx$ќ�;�##��+$.�������ٰd#,�b7����3�p~ݞaf��D��o6t{hZ��Ŗ�h��� �$*}-����ߣs�ا��^�����3~��6���t�	���> ��T?���5�Y��fw�9�5��1�~���J�.K��8`S����߿����gi���PQ��d�b�Ft�G����:2f�v	��;PB1����� �E�u��߲�L`�hU���̺����umD�0��A����,k�|�c?�OlX!�M��![2�|v[}:>�Ћ�tg�I�;���^�{ u���0�r5dFnu�B����@�[7 f��_L���\m�۠~/�ÓSz��=�y}�&����#Ic�y��`8H��Ƕ�����=?ـ�G�D��\l�A��ioiw�I��ޫF��A�U+dg�[]���H��C�
k��+�vl���Nq�FǧCz��}˟<3kKیY*y%Gb���*��u N�v$�hv�[I���/�Ab���5�R��Ǿ���z^B
� ����*�/�\����L�����2\��G�ӵ&�� ��}������߳@Y4��V�|"]�D�G2Vf������ϻ �ṋ"�K��mZ4��O̳���k���0)0T�h��յUW��ty �.έ��:5Y�f,ʆ!;:>�ޠO�n��a^1y����v�Z1 ��Iׇ�TZ[��^������g^���ko���86L �$p�S?8[Hɠq���1�P�G̾��lI�*}�R��^�|�<Y ���C3���iig~)}��t��&a��N+�MK�ʪ��y���Z�u�*�U���r|�X��؈� �rN]��z)PbT�ҩd�0ں��+Pwo�����i�QO��l�Z�V.B�*5��Uh`91ώ66F���Ƿ}1�g��ѓ_^�wF�=�s��0.�Bݨ�7o�[Ĝ��A��0j%	�W����^���}�h��W�B��c�#6#�s�\ �|VJ��nA��0�o�<�e3�ʫ�܀��<��|e��>��?6|�o�|��&���h��j�����iީ��z5��(�)�M����[A�Ƹ~n�H�4�3�]|�"��hFa�#�tE���k�S!�w,E8��簿�/�W�G�}��wӗ5��9}^�?*2��7�Z~��� k����?Y0V�"�w�����I���AO[��Ħ>�� iFdf�q~ʠ����dc9x̀n4��#�a�8gW�����4�m�3�=??���:><��ȚC�]�X���%Bk�+�/&&�����E����M���Ƀ�f���D���&�碚�If\#� M��n�7�^��1�s�+���	`����ڧ���l��kܼ�2�I�$Y��xNVu����#�Xm%
������?Δ�'[p�&`��W�nӛ����3��h�h{�J�:�v�]\#Θ�S��'�u����5��B�+�K+��/���^�w�=7��9�;gE��2�!�|���%}��Aab� ����o��O�T��LBK�w��v���~��!���^;���,\�6�T*7��E@�3��_�П��3�}{lx���+,�q�^�u@)��+��j��l+�|�� ���?��w��h���4D�.�\�?��#�x��U���=���<���H�ry�z�k!���_�F�̽m[xmP�΃%,���U9W;;6F�_8=�1&����y�|�E����_5����Ȫ��_�" ,"�rL21�~��3z��1 ��<2@�܀P� J���L jkD�^̾|�A��14�ŅT��` \K�d�Ke�l>�� >a ��v������Y#�%f#֌:N�$��P@�SÇ��v h$H��r�	x�r���<�upH>	�����0�b�5:oAD���7֔��|�A�UK�E������������,L�����̌]�2PVZ78פ�tP��v�6�?��K}�������)5p>�l0�|��X9��&HL��Ol�� _p� rrvJ/^7���^3@��[tgw�V��W� �d� �k�"�yMr
G�Y�ך��f �5pO2��Oo��^ӋW��nu�v��VI�T���LaáM�Q�&��R�2�|��$�"�	ͤMz�r�ڡ�v��2��uǼ�{1'���}��c�����+��>!|�g�����H���_����Q��n�^5�4(0 ���$�:g�mЭ��0)�T���B�V�3���^ѷ�>5��:?k����R�t��y﶑��3�yti�e|w�����ss�/}�{�n�/
���iww}t�cy�0I[��W � P�D?�_�?|`��P ������_!�O�^W�*>����_�e�z�T�@0��(��h� �s���Ǣ�׬I ��[}�&=KGD��'���K�:��WK,�+$-���F��P���������9�J�2�}M�ͺ�\e �V�M'�'l�\13v�V�(��)?h���)P������D� /(�R&�8X��T#9L����Ǐ�� �g� �	E'I�4��x��4d>�˔���w
�ބE�S���K4d6:%rE�i_��0�����������)w��Ӵ��H��!�@a
��F�x�1�z+�
i����� �ln(9ťk�<K�����3N5��ڷI6Q���9'�����G�o	�x+0&�,R!���-a�qٚ� �A7��WJ�J#R�y�(��%�kA���C��gD��^��� �O�ߡ���.� �X��Y˥:u;!�S|D?��Ҁߗ�Ï��|F0��5���k���� 8䪕�V(nG �Ն��4��Y���Oi�ė�U�c< �k����͑��n�u]�U��:����.3���{���E\��n�3���,`X؃�0(���9��??㔔=T��c��VV�4�_�9o+��eb����e�8<ڧ���_�O�����%��?1�Ԩ���B��6���~�pE��ӂyy}��Իc4�� a�{��[�SAXv�ݱ!�h~��EO�/ !\����dM��v�p/ #,%�;��uݝ?����HƁ�O�^������i�so�Y��Ý`���g�����yXyV+U��]�H�~6o��x_��3�[E,|��:��Ф>�R����dz~�i�|�0(ᇀTG�[�j�LH ���#~	��Dp� &(1�b��u�ӎ�5�t��	p5�s^`N�0��x��T�&���s<ч6�0�E �}��#��`ʍ�B>���A��I�x	TP��9A�>�F�2ţ>��@��[�ޛ|��07�߯q�� 1)�>_�}L��{�~�f���k��:;dF@�e4��F�4uٚau���=n��< "�7k����ؗJ��샹A��׍E�.��c���R���DC �8�w�u�����g���nL�n����H�TfW1g�`9��qHg'z���~��}��z�r߀�S�}���Z��&&��� �l=V�X�w�=�4K�?s��Թ�iZ3�&D�c�zMys?KÒ���������4���X?�$�Y�^u�^�����~��Z����N[�/�CB��f��BEvU�l�k�� 4�Y��p]�'��?��	���+:�?6�G��
�b�Cѥq�����[F֡����c�E��^�%�џ��+=�F��Y�[#��+m�>Ư��J�_��/,%���C+
���fO?����Mz�����u�;���� HF�������6*@2�CK~`���/M�/i�����,�1Kf}և�&��Y�~���0������f̘�;�v������?������1AK5�@$�^2�B�"B~������kw��o8�D�D�Kj������"\��|0r�f���#`LH����?���ϹKZR��i�8O�j�
�R��)�����߬�����{?erA�KW�Љ�Dk�E3�2T�)��e��C0C:4��_�%z�����t�����4ǖٻ�.�4����0x]���������y}BGG�n���B�W�P:���UY��}E�~��]5�k
E.Ya*���
gb��< ��I��2���. �[��0�z��g
����h����/n9���j���79"N%4d�J��
v����tl ����/���!�}������u��mz��.���ZȦ�2���C�����o�:���'tz���j3�+]��"���߁���-�}
�u�t��w���eNȱ����K��A�	���Ϟ�f�N�{u]A |���7I[��c�Ќ~��RҾ�w�`Mn����]L��I�]�~�l�b���hM��E�y��`e|^?�"Bp!=.���Y�u�(I��J@�4�|�T�i���S�Z0&̘Q�յunC�z||DU3�N�$<?���ͬŁ�7HL�P��5]��@����gX�٬9��r���]�!u��Y3�Z�J�+��`<|���/&лwo���ŋ����_�%}x�)�w6R�^�%	>�v��w�W��`WC[����)J��[O�ᘤ5\�$�e��k�=���1`��ٷzfR�}@'�'t`�Wo��`�v�3�_  ����~p�v��{�޾1��s=_Q�Zc�}z	2#T1��!�2�bG��>�ai0�Q����%�| �X]-�f�D� ��w�i�!*������I�R��S�����Y��u�1rY}皇�~m��4%�Pb�L�d1u�=�π����^�4�����;�ԍf����{r|� �uѥ� ��ce8 �0�6��:pux`'m�dq䳉(F�Ѓ�ӘYq��C�+����O������`|n�Y�:�\���D8�6����V��E (�z�`��5���'�^̤%���3|k �?P��7~C��.�_��m���H*((��^�'����O�>e�����"����o���S�u�;����UѼ�-� ��`��߬	>����_���~���[�W��D^�۱���LD�a��S��XvI�!�L%�Q���Ao`�r QՀ߭�m�������X�U5����������{Hᇝ�K��g~��)P�z��ӵd���k�"�ᛵ�_!��x�H���)�'N���n���'����",4缏��g�9��z�n����3चhlȘ����=6u.���
��"3���BS�"�G *��Ӹ
��W����*��\��]����J�c�u�6��$ �E�v���N��� �/�� ����������4B�����)�K�uL�p�%ܾcle� �}1n��NY����)=���e�g.����E�����s�<�T�s����A}����Մ�U �-�c�~���"̟ټw�� V���Xk�dހ��!GA#*~��kW�EZ�(k����/�h~d kWYA�JR$Ah��Gk�<;����;�t�� �����[6�3��X���~�f��h�F��������46[�V��7���RU9��DƉ���9���͕j6p4Si�|%��}���"=��� ^ҧE)���Y��%]�3�Ӄ��:<�v8(x.���r�YإT.N ��۝��تР6��0��.u{:�hsЯ �s8�4�p	"6m�s+e C��"��FJǵV*A�����@�/�jkk�vvn�=��$���<Cf�@�2�Z�,Z���\��O�֤߯hz���(�Ԩ�n��"(�i������s��Čs��$��x	j���`ƊC��j�{=��l0|B�*��$1�f��1�0����O���^H��u �?�߃N~��\�k�>�cږ�%8Ȳ���E�7d�Ck$}e�Q��A�����9t@�z��	��5�A
���]:b9���GM0���`ݦ�t�Q/h~qH�>��U�- ����vh��h7�	<�����Zw9ܽB֫�јg%wr#���,ٓ�ٝ��M���,Ͼ^ �0=v���������f���4�_�5}��W����kz���dRS��EַW&o�n�qR~��;�0+-�X�ך�t{g��ܽÀ��ݻ����/����g��#m��L�������CwI7���#3�[�9�OSv��h'��	i-�d>�R{]�|[�XD�����fNc��.��/���R6n��Y��3J&�d0��S	�%1����e����j�*����� X.��-�?|@�Y�S~�T&�@L:��0�|]mN���i�����Y�)�FNS�2�:z;�%��X1[[!H@e'�F�ͦ�X�j����Q�J�FWO@�)l�{��,��ڎ%_��DS��˵ӂ_Wङv��\ ,����h�.`��*/����xE����ǂ�Cs��P�`<�q�����rb.xO�(>�++)���:A0+��{	ڋ����X���Wk���Bj8K~`dxA�0� Ɓ~�ubn^��y���Ab'H������9$9���{2���>��U�I��i��e�F3Z�s�8?�H�l�e6o���|ek����*�>;;5���9�9����ρ8����DIx~���*fc�q~`IQ�A��f ��m>vͱ���/�؀�ϟӳ��x"���v*%;�A,�&��� �3	o!�k�)o%�k��k����p\0뾋,���ZM>���u���<�)��%)g�[��A�u�,p�Di�[Y#8�M�k�	��l5w�v8J��V�&^J�GRE[�p ��BK{{g�������?cF[c ��nd
��� ���� �4pE�u��q�-_�w5�>��k�O�~���
������J�K)pI�*�#�9J��鯬�-���&��1����l`��9s��e���
��7ig�@�:�D�"��<�%s�r�?}��>K�����"�B`'c
�,�4� m ��`���
Xd�tA�(��(�vU����󬻺]Y��ڋ: �KRh~�DS-eh��?�v@��4�@�h���A�]*JE8i�1���Q�h�\[�� ��^ ,`Ro�����)=y����駟؄g��.Ke���k��7��������<)!�I��u��K8���H�[�[�@rks�՛���&OdL~��'6s�#�L����Dj��H���7�XҒ�(��ML$���U��_1�����K��^'�&�F�Կ�w���M����Ä��w�1"�e�I��M��-�=8�6�>��Y)L���CC;<�U�{��,�T8\5 ��Ƣ�3�%�um��Dk'+��s����_�fk�j���Cأ�֬fH4��Ay�,M�Fy�s��A���X���y��+�W.x ��" �����$}f��ۑ����]��,,��l�� �䳟.�������Z�نH��5�����	����)g��at9ұ4@Z�% ���pF���C�^��������FO�O�R�M|�Q��#�7_,`M^n�w������ߤ_ŲB��˳$��*��+�_�M���uB���º [|�E#�����婧�<c���1-u�����NTs=n܈ы�k��I}��o�s������ ˆ��zz��C�<�x���o������r9�5y�?o� Vh�ۭ6��=>W*�x�,Hqj�:ߋ|��9Ƣ����9o���� pD|�"��&�X�b����󗴤�ȵRH������_ŗ��%]��6�r7�<�$�0IS�GE v�y�=o�L1GN�N�2�|-�R����/m���G'��P�>�(��$kHh��<[_k.���{z����Zah�p���3��j�g-#��E�?��$O#T�Y�5z~ ����V|hd����$���t�dyB�č�y�t,&@W�j�N*ڕnI:}`L��7�'�G�X�@�'�#'�$m�{����40�A�����φo���2}y�} Xʒ�	`�E��#�-e��"��Ȉ�cJ/��5�������Hl/༘��LkR�"Wh�N�{p�\���۫#����ٰ���� W����WA�����胙@�R���I��=��g6��OK�	I�7vHf`���
�4&)^$�:�fB�h��<�v����tr|����߇I%�(��#I.�*�gK�Thl /G󒮟��f�j	|�$�2K�3+�����@ɭ_�f���^M�S�X�P�W�ӓ�FO������Yb��x}Z���I|4
c~`��$�M4B����c-}��&���o����y xR݋h<�2���e�_�_��`�����\u���1q9��#�l���=hM�e�W~1���0i[�4VYm����<*����YQu��|��� �"��Du.��
�1� ����Y.�mb>ڀ?�4���f���h�u2Ɗ�A�����Z��gC �>����m.*�}��k���
��}1��[���*�m^�n��d���A�n:���r\ޣo F-#3i[��;88����&������R��@��I�0�h�|Y}�$}�� ��`���X� ��9Y�{���I��ʮ�<N��VmN�"�%-�R�������]�i �0�?�O�5����f����|Ou�S�w�4���ʔ_ksq�0)�U0}F�,<��A'A�(ӇF���q�p�	�{n��&�؋aY��u����`��"��� ���i���ʘ�vX�����5��%� [A��}���4Z��2F��ϋ�F�#�\�'o��`����_��rލ`��^w4�Q�]h9��@��|r�'���
�����mwQ��½ ~?�D��4�t��f��;���1��Q�߳1�/b�����yegQ��$,T@��a�~���gm�C���6�FW��
�|�]A��#Y��UQ^��L�S,�Z@���� Ӂ��"�t��A�#K�eA)�l�;l���M�c�Ȁ��k��XX�#�밇�u��=S���@V�/8)C%	�)(���ZҒ� ����.�����6�y6rͼM� /��¬�2c*���x��R�$ݽ=����3	xU✯%��2��KDI�!NMC��9>L�X�;T�P�8 |���7������3>;;�Ë ��w|I#>'����0�`���������2@F���(��	pM��J������V%����f$��Gq�e���H��!4�������d��	�|���0)�c1������-g��΃�Gy�\�!H�S%�7>�ǎ ��9x�5M�H���i��v�#.��r?�����ё������s��
��@K=���V\�
�楉k3M_���	��\���0S�d#J8x-y-�b:����,��)���0��������G�}�\/�����������U���k"!���,��&_����8Cj�l��zt�~�=�ȵ�/f��_|�YM�q$�a"�ƳB��ā.q$��Fa�b~R�9[ZU����t��=�����f������Y}�!���I��E�M<�Xx?(�+1�􇜧7���#�ݚ��X���hl��c��|�v5��g�b%�g��7Eƕ6������e�����5������O((����8h=~HE[+y�u�-��{�q�c��Ԛ`�K`��c�7��;�g���y�����L͒�wu�s���(�`�m ���"5�z�ԟWiᤅ����=�4��
�p�}��)�3���8� <�<����jne}(��w��� r�����_	/>�lya0z��_$j�d��e�咖���)a���ˉ��#��I�W�|ݛ�<�����E�j��6�0,��;I.@/�t`��'},eZh[-��/cD�>%��phuʌ��D`�XD�IpH�`�<yBo߾������޼y�P���h� K�{��6o�y���j��kD{���_ӿ�ۿ���,�" +���yC�i�,I��uV3, X�ta*��(��	�G%i%r�~K���c��h�Y$����a0T��Q��6;����o��傇��r�h�-E�_���� ` D�z�5�Ӭ��k�u�SiI���g���.k��>�Xc8��x��=��	΃տXk�aF�˨ �̣yH@�p��y�0i��`���9��M|������.@�W�hӅ���P�:�?�
��5�8�$bpN�N�P-%�d���5N�O&U�y��D����A�X�������7A�3?���ddw�4���㥀h�X�>?��X��E�ބ�J���ޠ,?�i%�g��\��-�����yp�E�X�&�`�)��=Q�W�)�d&�81a�0U�ap�ꈭ�8�I���I�V�8x\���U�=4��uB/^������={�2�n_΢5�Ңfi���I)X�X�̸�|^�|c~fнf��zK�"���G
�Ե+�]���-Q �Z`�"$����p��0�
�A-<N�y�#sƖU2@� BX@ ���x�c�-��z��OE�Sk��8{��TQA���{Ek�}��>��]�wY�t�ݱ�����I�/��"y���5��Uc鮟:�4ʇ&�`< 4�&� a�h�]s�,�{����xJ
��$u�h~v/7�x�ལ/�6N�zn���J�g)O��+iWBZ"}�\7%�p}�u
$)sVZYm����Ϣl\�~y�]�8��C��H��p�J�3G4�!
]�aO�e%�?Krql��F�	i���#I���4b@�o�E�|���<���sK���E��1�q��~�c��H3F>s�yhQ��f��1/]'��sE���{���~$��c��`$p��5�hX�0��~��eU*U��V��\�7�&�#�i��3p�~���D�']�{�&�^����C�2�WQ�\�r����k�LK[����aV�"ZS���Ӵh��(E'cѐ� Sk�Oޏ��� �cy��"���Z��?~���ڰ8Ă`� �2�_�	 ��a�Jf<��e��*���	r`���C�h����Xª�*���Y.O8��>8�y)vנY�p���ɷ��sa0�@�q�
�̷�_�
�ߊZH�V�#Љ����Zd���_���m�ɚ�zdnhshWÙ�.�O��ͯ�=���3���vZk�g%^��X���Ǻ�Ԭ�v��8W��|���:O���5�nt��u�0,�t��]�4���~'E�v]���Z�1�Α�_�έ�0M$��K�ǣ�ċ�������w���EL����%��UG9�r�|�4I�[�\�o�F5���g>��(��{Y���{�_���8H��k�p�����>__���m�J�F�+8�Ԩ��Z�B]�S �J�I�nd�3::i�����C� 3�_�h(R�dO�)c�m�葦�0���i�`eiJ'=a]��0�Y��1暺j��I�X3��0�y��R��IGw-���[Y�a�V�3����mV�^٤f�L��_�
���Q��r,��ڽ>���զ�Vǀ�J2���%B��r�
}hl�j�fz���Yk�X�5Ӛ^}^�&p�:��N�~�z�k�F��iޯ�s�_�`�͙Q�1� Q?+�m����E�h�,��4i��~�2�\�m�����F���<�BE"?%�Z��gA؈�W�-�:7�ϸ���u�=�2"��_�����2�Ղ���g��+@��)�`�a�A!c�FL���' �1>�KZҒ���O�\�����y%��E�]�묙?P
�R�
a�(3�d�R1=�vY˻��J������;�po���n��Z��l���i pX��E�Ooߝ�����'���{Dp�R�0t(��Qz)����J����=L�vW�f&1+ �g_��< *��W��p�<_��p��P��fH�Ff�Z�R��Q����'�2���f�=s]��W�t{k��ݡ���6im�N�b�˕��д�զ��S3��ū}z���O��M�fdꨑ5��z��.H�':]��j�| k��\�!Yy��Ɨ����<Y�.cR�  :�ɤ�`MX�u�-B�����ɳ��/�nAs��,��%�~�kОׯ_��3ڃ��w���g�[�iɮ	6�> }P���[YT�%��`=��9�5N��>�k27!�����O<`A�ٟ��gz��)�i� e�ut�~��KZҒ���1�F*����h�e�nM�����L-.�3N~�0Td�h����0k���5z��.}��}��=ػE�w�h�i�̙E� _�R��݈��l��f�m��	H9:�H�;}U�$�@�6�Mco�b�f W��j�&�9�FO��<��g	@f1M,Ri�vd'�Y�p���j��6���z��}���ܥ;�6 F����e��J ��0Y5���l��l����x���<{G������p�c�B֜^��h��(��Ƭq�ߛ;�|�����qV 0�C�Ҋ��B�E,���n: `h���j�]�`{�#6� ���y��/�/� TW�7h��� ���k�<��,m��.�k�on��"k���H[.i�ckY���1���#������ �!$����s@���u�GK ��%-iIK�,��T�I-�A,������I
������u�a��J�����.��]��6��ߦ�翣o~�Ѐ�ZkF-P����!�qD��l�5Z5��v�B�����z{D?��������/'֯1���m�����~Z�|��G:0���~�y�p$�H��V�����5�>���Т��h��������}���Xr|g�"�]��Yis�������o�����f�V��/ca�5��Z�1�6C���ޥ��ܥ������^�_������_���}�qXf��K4���Qy��ѵ"q��5�V��K��C=G��hK��_�[������[���E�"$�B]�	 ���&ۋ&W@�-&�'X�P"�D�_W���X� �<4��o߶y~����0�*�":�2u@� �gZ�5M� ���I�6���o�N���Y�U�,s�w�{��$sZ����ygg������o��/�L���Ǐ�O����|��n�A��r6gt� /iIKZҒƨ����$��$��cd]M�os/
�]��<4�F�)�(	�ȩg��6�PĦ��4h��T�mm�3������y@_|�C��a@�K�~��A�`�A��i�X!PVV�\� ��I[5�7a����)u�m`��X����/3jI~�T[x�6�tYz��>��A�=��Ƭ�'�<�,�2� �h�v��q�S#�6�j�W���[�ۯ��x�`�j�>���F2c��$����B�������Xߨ��M;99�quz֢n��>���<�o�l�ꑼ�'��j��}����=o��em�B�
�~�W)T�>���("p̖����>F���� ���H�	 �}~�M֚_ d�_�*I�����B���#l��I�t����+o��[���������a�[�n�5+�G���s^��q���KZҒ���1�p.�yy �H]}����0P��KL6H�5Y�j���n n�Q2�������;��oҽ;M*�-j]�R<l1��<����e��a��A۔e I�Nam��Vj������#��暗���w�f���#k-~��=c���asxr]5}}�x��$! �M�S�GխKV=gOR/}��-�g��xX�߹�s!�G��Ѥ���3���N�o5�R�ҠNèm��r�-�J6Z42O���X���W��K�R�>�����;�w߿�v�ĔQ'
��ӚE����ӿ.��@k�Ƃ�D�w��<�I�E��I>������|��ө���oQ��"���B4� %��.@0�8f���� ���ŋh��ý�J��n�u�O�3����U`\�]�P�c���_<�X�]��ub���������w�X�U���C�dC@pH��X�q2�/9o�| 8ȕ�\�vIKZҒ��"ڈ�b��YY�����Иx�u/���]���4��4:f�!�Q<`Qo��ݻ��/���~�>|�*%Ì.h883�6�.���ym�*��2������VWh}m���os� �G�hY_M���A����6�����h>'���@�&�q.h�گ�Q�� �:�e���2eX�O�mȚK�g�~�i�]u�g�3���@`�о=�	�T�����I�v������mZmB+l�C�2���FeQO�9`&f��>���T�4i� �������q5�w���ٵ��)�=+
�&w��gi5�ӀFޥϤ8Ok�S=N3�#�F�P��s� �m/H4� �8���{��=<<L}{%�����lmm1�Κ���H�o��DX� �&�Z9�w@i�iȷ����]�D��F� �+D�ϝf�M��<�-�+�ov��(���y�X���O /�풖��%-�&1��)�� �g�G��4]&tC�o����g`�l�#h���F�m4V������w����:���`He�Z�t<0 � `|�
��a�h�1R��nQ-P�V3eާn7��/߳)"�GQ����pds3�QF��<F�h�$W#�l�~�w,>\.��r�4u�r}��j]�O3�.hv�v�׌�c��428*�H�����T>� ��.�WW�������szx�6��Oͻ�`�_
�d��c�?l�Ǡo#���	����a^Ku���!��/����iπ���i��MY�L�s�>�%tp��f�:���Gc��X+Q�@�)^����zK^bhru�`h�;�� 1�ja�M�[��F�BY��>p糞�V����w���i�'�("�F��S>���ݧ�V�Sl�E�p v̶���y�Eߚ���%�]Ғ���E�$fS�[cW�fՎ�l_%�8P̅�)u�yxYk��c-WJ��ޤ�w���mZ[)S%�Q7�RԀ:��lw��c  s���k���5���{�1H�ʬ�{{��ܦ�����1���,�(�� �H ]��W�ܦ�I~m�������E�I*"��AVD���n58ҟ�ݭ��{�c�9�a�Oa�݉�y���k+u���}�x��6j,T�`c����8v�}��< ����
ՠ�a-M���81c0�sU��ڠ{wn�cی�S���9�o^|}���H�&��4X+\��!����>}����>����J-�O���h��Nk�� �O����Y��=ןS?��1/a���rо�����P�r.�Q������	�&}W�����r����~�+�>r ��%-iIK�J��>w�(O�����(�F�{�P:�B�#�Bܠ���6 >�ad l�K����+U���P8���wg���)]\�ث�V+��j�v�V�޽-j�T�^������&�P�A��^�;����:��P�sN�*m��{p���0<ojf,����f1dn�\���a֠La�W���]�f�\��,� �)e��f�m69=��y������j�6W봳�F��ҽ�M*��}���|�>���1�%}ppJ/���y���6k5�\[���u�C]7�Ѱæ��IGJ.�6k�{{�n��:t���?�݉�����Euu����#�jM��5���⺔�cA��+���:�aP�b��j���|v�]�����f���X�܋�`��p �J��g^W�|�üu��o�zդ��U���_V��I�x�y	:������΃��h	����%-iI���(|hЛ�	p���}��'��̍�`Dׅo�`p�?���a�h}�n@�)�[���"*Q��3�e�^�2 ��	����0 x}�B=SVcu�J�2�e�ۍ�6�M��\c��Q�:]��R752`jh�B� �����;b�c�?��AѴ��sZ{������>��I� �w�,� �x_вh�jU�Ҳ)�y��ww���û���-��^5��u~�V�R�Ӂ/ߞѳ�'tz�e�g ����D�z�<���J!�?��ҕRLk�*���2 x���8�1+O�o4c�j����L�.O�-kͲ��O��t�S�[�;v\���r�/
����֐f=���a_M��I��#��ĵ�&�+�K�D 2+�kˬi���k��]�\�I=�����A>�-�<?�U� /iIKZҒ�t�R�O�S�K�mJ�џ��	�?�+`Vhsc�VWj��O�!�� �vwH�������0����5m ��JD�� ��~� xc�0��3!��5��J�L�=ޣ(�R��n�pה�0W�P����������ݻ���h�|~r3�N�	�$�S�usjO|��9s��\A�����9��F�A>d�q��-j�[lp
!�J�L{�7��/����m�X���B��������x}F�_���Áy�Fj���N16N�_�����G�.��_h�ڤ� ת%ضH�v�>��̠}��>�sai����9[@h���F�:�� � �Z�pi���>V��7���{]rʦB+�ܫ�% ^Ғ~e��ҳ~IK�P
���~sI*pZ5`�f�z��ڻ
rRrHg�q�����a$/�ttԦ��u��A�5�%SV� �J�k@m� �*5M*Wlp����:��ۥj}�V��2�	æ�O��A� x{g�?~�+�ſORhp��3��&�Flv�w��$�:��C]���5\�<�[҄�� ��H�Y�U5 b:�h���9G�=5 i\��;Ԭ����
����Κ�}����)*�DMy%��wh��C�N@�~��Mό�A�C�ʅ���66j��ڠZ� i�eʉaeP���&��������퓼��e,�}�1���bv�y�a��&?�ۭ����3/�T�($c�y~߱N`,�/0>�:	�a̓���Mo�&~�3�Rw-s�k�X~�4�Y��]7e�fRsy:(Y�s��Q�jhs&��% ^Ғ~U�}	|>U���O���W�:<�qj�����o�o̚��#��d��b�9I���Cq~S���Ц��/=���h�w���M[�SnL�^�2��T��?{��%�q�P�}��G3�(je�^��w�;g��w?�'�]�ER�f�c�{�����_$d%P�v�3� k�&��H��u�w���[�Ͼh�0�X LM.w84`�?d��Ç���^�x�L���T���$��</�a�Z����T��� ֦�ڇ͍\�e�����RY�jp�/"�~�����_��z�3�|,E}6O�Cj���)����}#@�(�,�=�2���y��h0��y�Ogg��E����Q4��F����:�M}�����uc.s�
;�2dja�]�������߬�Z���<T%�j��R�0� n766XӋ�#�����9�!�<�$�}��i�����}e�yv/ZV�I����,�r���j�ݵ�*��\]����+�ͷ�	�f xF�.|f��6Ӥ�Iև�YC�jm\���L�B1]U�O5��?A�~�1�e�r%�ei`|գh�u7>�W>.�:-iƶȟϞ�䓘<�����Ξ8H��'L|R�2�F9 ��F�b��~p]�~�>)��C�>�q��G�z:���3��9��l���g�LN�h>3 )K��A
(�hз�ťE����'.M��U�/�W�8�V�Ǫ�|u���������Z��v�!�n�ߣӓ35<���g~��iЎh����U���<0,�k̘ds<��7�n����q=�C�c&��Р<�Z����9��!��Hr�aG<����i�{�������8-2u����%��&������d�M�\%�s��o����������E�+hz��ZM0F�&	�ý�`y�>�؛��}���.[��wvI��
��u����4�_�7�&	�:�����|�`R}f ���e�������{{5�zՁSp\�e���2�E1���&4j3!���	��ĥ��"�!��`�i{4S[��t;���l��y�gɷ�[K�}רRR Lx�#���0�q"y�`�6������sZ#h�a�B;� $��(4�7i����)b\����)jڴ��1���Il��To�Q�٦���z���b����;���Q�>g�kr� �����ۿ��VVWC[#��_�!�ĸ$��>i�F��nJ׬�np^�;�9������u���I��׸�.�[߃������觟~���M3��YkjǑ�;�=\[��_ܧ�~����a�J��72��4Zh�i�ұ�q�&���:h���;���b�;4���ha��{�������6G+�`&f?రETEH���$����O���[��yw�Ӊ οw/E�롵۲�]�����N��H�X z������~�����Y�@W� e\0����40��SZ�_V�I�����<�v�,��X�Y q�#�£KP��M���h<ʺ�S��ْ$�;\�S�\&�K�7̷K����s\��"�4�[��� ��<t;Ό����q�n�����o�fL'E1���LS�MG�tjp�>GH6Gwc�k���c��꣟-�|�o����i�F�3��xU���6��>���/�	(���X�=\Ft~�3�d� b�x��AN0d?�8��`XZ�;G�gC��=]+Ԁ�i�ѡ���$m �B��p��� �Z9_�l��nc�~��9���<����7 �a���0J��9�_�gͮ���n���L�o�T9滿�L�^WE���{�8��Q�r��|�����׏����9���˗/������k:;?cr�@�{���_������JÌ�e����ENjNg42 8��{�l�����9�"���o7���EZ6�kn�IA�B� �{��c�؀! r $ �$���Z��Y4Nr)](?Wq�~��L>�\a�$��GW����}����Ʀ�YWH^PB�� -���c����e���S�	yO�*�&cD�p\#�ʞ]�.Bz�@_����
��q0ݻ(�UIҢ��o�zUFz�����������}�'��h��>����ďSi!'`�&њ�q�2M�� ��f����P���Y��z(��k$�x����(�u3�Mz��Ues�� h?A!���ѹ*%'�0e`��U��n�6k��M^3�Z����}xH���\%;�l���l)U)����v��������Z�����җ_� �@o^��a�}���,.�����.���i|�y�Qir������=���s::8��r6�j��:�й�HIS|�HU�34��@1���
�G�����>��c�|̖f�]��|���N�#u�T���21�D��OX�vxt`�J��P���q��\�[ۏ��}䌎�Qm}FC�ؗ8�_|�����>��Qߔ�<�wW;�f ���<5�x��@3Q� �Nӌ�Ь�Èz���G#�-v��"�k���=�s��!�E�l���/߷~?ET_a���0����hA/JE��_�Xǃ&���޽{���%0��� ��o�g��@�&�o�� �5�\�.}pϸ�<�����u ����[����l�}]��w��������<��|�3��@p������� �ь~F$`�{.�J��J��Ҧb�Y��N-&�E�����y�Ϭ	$nl��l�I�f��2� ��\�o��BE�F�5<Z�+�+H�
��R|%@X���;�l�wyrrL�{����.�=�����7[4�� L�MP��/P�GТ���Q���D69:��2f�75�R�4`��y72������ F�ց(���(�m������`=& �( �t��%������qY��"0*%����
��������X67w��Z���ܧv��b���F#���s`���R� ��;+[�%��X����Qh@��g}�?4 ��0��ħ��mBEI���ķ��~�i��ְ���
{/�"���i��u�� q� x����= ��دp����h�*����]� �� *Y��|�WMz_�`�� ಹ9&��PM�~y!�;n�<Oܘ ?��rE� A���������w[ <��e�����Qk�Unn��>�0Vf xF3�э�^&/-�+M(ʀ��#�i0U�����/"G{���r7>9�r����	6�����ﺫ ������I0|k���L�|tC�["��CNa������iu�.ͷ�p=4 ��Zu�n���i6�o@-
�@2�P�V;d�_as@��[��{Bo�lѫ�[����Z�9��M��1�u�~�F]�|�2&�v��E�	�|��|@����Ǟ�M�1������^����|�f\��ϙuc�¢$MQԧ��>�}�Mk�;���<�{��Ż��*���4c�� ^5�Yu��<`����&��-�u:<����>�y�M�wX�So`l5�>�Ӷ�}7��͜Ϧ�q�[k�ǂ-A��k�}����k�+�Hjmg���d ��	m��y��M����o߾ek E���w�Z;	�W��Hz$"D���1��y1����:5��.�gF�D0�����oi�~�G�w�e�ߤ{��e\��c۩��O�N *��L��o�1�_M�a�ux>��eBz��i���m֙^�z�^��r�8k����/3 <���R��"�����Rh��c� 00-r�-�H��I_����I��`$ܠAr�*��4����{�ް5�
�ǵ6�f߽�sD�Rsg���d��x��df��Č5f�W�7@iуuH�.�E�!S\�Rk�A�"�o�!����2"D�����xH�_�����'��ڣӓ#S�j��u�8�G$3,.�c|��޽�"鿋ꡯ/씑�F@���� NR�p:i�5� �� Ի+M��36:�lI �@��AF�	��6�G���Ј��W`�C���;tvӛ�mz�|�^�ۥ����ز�ӷ�
���O˛]D��]��	F_=j*(���ИZ-?��a�^g:$�4� �8��	Z|CQ�w�2��M���v�|�ם'Xƍ��]k����4<�O�Z�\��(�@���k��4P-�#�q��B'�p�ZD;<<���z��� ح��^� �hF3� 䓘_��wD$�"ل�W��=z��4�v7 ��)�D�O�e,|�H�hm.�r�߿ςHse��Rz����â�{ �]ST�/> ,�c���+�<��Kj�$u��d���'�mZ(0��0��u���Z\�{�3���=��{��9E�>�c�Y�m���i`�F���A5n�`�thw�=��/���|����3���Z�<��+����A!K4Ѥ�C�k���f�&ic��2�P?_��
S��T�����[��zal��@�9�z��
��_f���;��! �Ç�����}h�5�Q��A?1[���P�È�W~d9�l��~Ԥ��}�����wo���:<>1c�e�R�����]v�1 w�*#������_�@ze�d�)+[�.Q��c {��KV��
�׹� �������ڊz`��?�����E��B@2�ٴ����	a뤋Կ�y�2����0�����:�j �"���v�#�__��y ~C�2l���~�4�>.Є_���|��������s:�I��\D3 <���H̅��GC�lwX'���+f�u�ٰ�yAc��L$o+i�L�xٌ|f�E�̈�@���y}�$p��
�u��+����.R����Q��E�% �s��Զ�ռh�k!2�?ءW������>��ݻӡ��p`.�c�s��<"yf`�#�fۀ���lf�����z��-���&�C���3�Ux7V��� {w.�+��n��g�G^�)�7��+)�L���;5�[T�.>���ُ� `�F�Qb	�s�eßw�?���}��Nmd�0=X_0��Q�0G*�,����7T�Z���4��C3�6�����/������ǈ��e4�@���i����{������������6_T�2*�\���6@¼'��9T5jrQ��c�:Ͼ��`��N]ͯ�K�|���M0�4�A�v� ��'�W�U��� ��?��x&��"k�i�[d�PEV��"�e�K�g׺�L_�{!\��ܤo���Ǆ `��}��n��ޣ��R�߸ `[^�zE���9������$����gE�`�u��8�7H�զ���	f�UH��,κLa
ˤǷ���"����D���u��"fep�V���e��i�i���7w�3�z~ȏ�}nk���P������џ�<4L�1����~��c���a:�4��h8 A��^V֙�5�C�͜h�%������/��^һM�/"͑a�;��W1k�P����k�'7����w����
�'�V����e!�׶�:�{�U�E�D+�O��� H��ͻ�'�2����C:<:����u�m #
�㇫ ��3����w�4H���W�:�����hc��������Џ�|O;{'�	0�o�g��� X�\��<J�  ��IDAT&-<�����h��*��}GE�:��U��n��yn@@0޽쁾y�[��9��}�f��G|tEx
�Zt����3��o��\� S ڒB�����+h*��*��o�h�"Zm�O�" (�\�+�NJc����3ɂ�2��T��,���?���򗿤n�}����~� ����<Ӣ!���RVY�� ��f�����e��UY�|�n;S>-]DJ�Ɨ�3�t�� �*MS>o�����W�f�=��2�T�ν�L������Q�%�a�h��"�M�#�o���|y'�w02��is�^�آo���^�zO�HiS3 ��<�\ΚBS�@��'
`F|�NMb檌1��L�}�������h|���k�[����˼�������q�? Tk,��#Q��9`AG�0�}�����kq���Ӟ �kD'g�k�	���5�����逶���?m�w?��/�x����������
��$�6�a˪��I�^X߻􍏢�E���v*oQ��jZ�]�� 
?\	�'tѵ�J�@�6��1kHq\r����O������BȦ� 1�F;q� R����
�B�B�-Ϫ
Fy��}�2�iU�N|J�8�vZ��j�3��v������Dũ8=k�^3ݴh�����	2�h�g4�}Rt���S!͐�n0��P�Y�|�VNF0�`��0�̜���ӷ��nЫ������ߥ�w#�isd�^��3Ø ��hprD?|��^��e-��i�lL�6�(�����W����\��ߋe��*ڑi4�^RL�/�#u(An9 ��.c��0�a��r| ����"y������z��I�٦Z��d�a,>�V��Mf���{pxH��F{�l��,l>�+��
0@�<���ߥ~o�ywvN���-z�n���1 �7;4o����\�H�䇻Y�������1�e�i�gW��
<\f[������Y�z��;b1_���� `h�E�/sR���"��q��SLOQ6�����vp&ψ!y~]��~|��:H9 ����Abv���y�����v���溠��]E�A����>�x��ڸ�TS���~��2
�X���A��iJ�8��\���(ϙˁ�ٓ��Xuߥ��{伮��}4�3�ьn�&0�Be�6��4�4Ŭ)
��qPK� �	����	I������>�ãSz�}D��ӽ{+�0߱ ��3�b�NO���c�5����w���C�'���4׆��F�&�����q��W�6b�V���
�,�N3V��U�(�`�zj�����\�_r5���WI�TKa�$їف�+��_~�5�Q<����n�����-��w�t���_��z甙e���#��� �����^��6 �����Ma݌�ZÚ�Ǚ�T3P�^%�c)	�V�����u��ӌ|ƿ
�2D�$�� ^�> �r#AO2�u�!��7�/̐�$ў��SP��iǻ���`haA �=���ã4�������dA[P_D�_Z\bm3hR���|]<~����ϵV�e� �>~]T&P���$A�K��`��ԭ
� ��f4�%f��i�v�i$�3���R��\��h,&Z�8ј�͡C��uH�aD�'=�wi�����ޣv�i�_�A����3�G@��������6(|3~��Ǭ��K�ؚU�fhE41eZ�I@`�v@|�u�Ia�]�K�0K���Eǋ�^�a͉�Ւ�C:X�u�C��ͻ*���ؗ�$c��o�8�q�7?ztv�`@G��ۥ�7�Ԟۡ�cHyd���Fl�?�M��ܚ�5)@���z��i��Yn�8��\i�!���/��o-l��J� W
�� �	�f��8�%ƃ+��"���)�-h~%������5о,�	��i��stth�Y?]tो����Oݬ/ �K�K����wNhBŀ�G:��$r�pU�m��q���E�̊����>�>(�Ѧi�۟�j��k���hF�\�^�d�
��ߋn3��(}�%����������$ܔ���Kd�����OG���RX0�&bC07�� `����8�f�I�9��-���?�{A�Z˂�j '�����T�n�l0È�^5�zU-��2��_k^�-*�_��@.0��'಺�y]����b
zQ�g��!z3����m�rV���E-qb���Dfl��HWԥ�vY�,�$#������~�3b���Q�øn��C�|�"���6�녈�=��P��U�in.� �\	4Uٛ���H���,�0 � R⓫˞\ �L���j~��p�W�iH洞�b,��8M0��4�!��̜�����:����g\D�h���Q��H�O=�u��I�W���n>��eEk�o}�4g xF3�э�I״�W��	�4�ӑ˨��>8�E�M��$�|3����d3g\��6q���7��r�޴A�BD���+̝a[�w���Z��d��	#D��(�����n�[�Q<��|.y��P�vM�  v-,� ��<O+��
3���VCyq�:a�ܼ�. ���(��'O��VЂ��G�Y��u�Y��F���-�������j��Aa�֔]G�t���0e��id�h`�#�k߷q	��I��0�k��4tU��L�4�����z� �9Q�#@B)i���>��	�ϯ���h������.~}���0��Zh�s��	i�`9wB�A�B��<|P���u�!E�p�YUH'B7hh���j��ˮ�c�2�rt�&Yi�4�WN�p+�S�-0�	.xnF3�<��[�>M��=�͏xz&)�2�\��2�vF��6��ocv7Ut�{�̾(7&}�)��L䮏%s��(P��5�,�A`��I�?�9H�m��� ���x%П�Au�o}�ڝ���ӯ�kf�'�i�<�Hk�ЮP1l�$Zl1 �v�\��v�H9_�`I��d��P~2> 8h�eȭ����Ǐ� �o&4t�zhM}���q��6�zZ������5�<Ht��=$��έ3 ����@��ˠLk�DǕk�4��X	�t2������H�=�}`�p�����֍�kiz�.�l:��;w�}��+4��ܜ�\�]��(Ȣ���C���D�v^t|��J�� s �#�2a�C���t�.X�6��� ��B�C]/_ۮJ�>M9y�;>}QPH���ҧ�|��5��0?�>3�WN�<G֞�����hF7E�����%�$����_Q2�&?�� 5GL	F�D�Ϗ��6��>��W�6���Zo��������[6_��c�En�;WQʏ�X��f�a#�'��3��S0Ϧ@�L�d�7"�z��(�4�ڱ���p:aN�&Z��FA=8<�ã#Z1��޽���?���Pi��n�����h�W�^��=>F_4���D+����}�9�yM���,&%�i֠i�	�W���������Xj7�ٜpƚF�1Dh�Z��c�c��l��D
�A��7���s$�ĸ@A�80XD9A�?�o�Y֦�����������2&�H �s�_�`&9zmTJ�BIj�A��^@]�&�bh�Ӧ�RO��XGƘy��}��WR�[4�e��W���ehM0� .ѵ1�%@����j-�om��K>[���{�6����e�+>ʍ�UƁ\
U�>]��I��o�u��7}��Imq� �N�㞛�+�I/,����$�ьn�d���
]X�����D�+B&�eZ�� �1W�\�i6ʘ�2S���j '��j��O��c��{5�u���|�D���5�Ή�$�8���`'�%�J�@}ү$�4@H������#�� `�жtisc��/-2�f�V37�n��Y\��I�ƊF�S�ɕoyoU p�&�ƺn���|�lyFU�����������۷�����B�D���r_�W,9��z'V5�YA2.���q�D���}�-�� XƝX������}al�洽DyM����(Z�5Й���U=��1��jg�� �����-C��I (�K�gI�}l}�Xu[��|sX|�v TQ?�`��F�%}�\�+O�������chaՂ6Kt�i���)�|�~�2~��7_������?p�GWxTv�$r�E�ve�3 <���FI!av�RB>���q��ۤo]���$�U6�i6(���Iur���3�|��B�%�0�̴��(�ˬ�Ƨ�Z��.�+2�@��q�>aJX�8���yD�_<���Cz��477o��e���$�ET6��$��*���Dy͆�5i�]@[�� ��&^�ͺܓ�c�'��l����G��ꛒ!�0��X����,���Z�Xͯ��%9��K�t�o�&�y-�D�����i?yۤ�[�:�D�N�!��y��2��.����Ǟ={ƚ` 9 E��B��H�'\������u�_�u��"�n��sK���<��G,R�}�f�<w��:�b���v��i���2�X���"`��>��a���|U��w]��D�����{����3 <�����*%�Y���
��<�GG7'��2�:��U�*�����<SG�����K`��j-�����
�U��yͱ�ҹZ�4�����W����p�� �>�j5I4�b����M��Zg��g��h3r�x4.���9�f��:��I����&<2�>-�� ��^�mR&A��z�f^l�����_{g�pӖ�o1��$y�ƒ{��	��A�-p�;g�Cn)$���-�lw�	,�ˑ+ �j�����wƌ�[Z����_����_>��w�XP+�t}��p��L��Q&��x%)��[�[V�o��n �2�a�@{�D�F;$O��?�"
�c�}�>��3�}�pS>��gR۫����o/��Y�X�L]�>��u����]_t� �hF3�dȂ^�|y͓M%Yha�YŜ�c"����|`qZ�nYyӞ�DU7l7(����$�6�ˀ� ��� ���&L�5Ui9;/-�$Tӥ c� ��{ai����)�������o�T~s�niS����F����IoG��"AG��T3pZ���e׌�\�j��Pi�.2��:�91����������~@g�g���8�7G'O@N����q.);|D��~��rL|��c�e|�9�)��R�`N>|��6779]!�=b (>� �ŵ���~�6��s[�_�/7�V���g�C���vw��M�$��1?��������x]-��[Y/���:Wl���k���W��lٴ�HA˴Ⱦ�u��� �ьft�$<�5��(�@��ƌ�j�6#��_�Q*�_���nR$0J�J9~u4%�^䔋�p�P����R`N8���5�/���^¬��� ߵ�5���'��gO���л�w�q�3hg����P�8)�>�{^���mN+߮���j����D���6ż.B���)lӼ����[�Z������Pm���FL��^�m��,���%f�9Z`��/�I��)�ఀ"/�]M<�n�����M*��[����(\~O�:�u>� ��� �A�Ч���}�y�_�����U�_	<�
~t;o���I@.@,�.��� ��[k��7 �@>���~�o������4�����-��T~\���,o0m�����9������<� ��f4��8s��ϕP�qn�sVs�<��4�-���Iz�`�e�\FqR���) ,�0��̄�IDI]�*���Lx.�$q�}�軖� �o����I�t�6�p�^���6ϱ����ۧ?���lv�
��.krM�w���E	c�� ���h��Z�ZW�����Lc-���/�?��?h`�x~�� (�ԓ@U����C&�Ʊho���ǎ�(e��� ����@4�
kK�<o!�t�����t>!��b�!����|q.z\h����I.N���L�/B"��� ���ұ� � ��)���4  @"�)1R�H )��Ԃ�~}sG��X�C[�.����6Z|@?R'����?��?��>��R��h�MZ��Y�]����b,'X��cZ�	��89��hF��%��,��j��|�M�~�V��n���UlD�<�Dk�\p��=>�1�
&o�ya���?��2�Qd�Ϲ�m�\�jt�O(���4��T% .�l��٣4�/R�� �폈,� ��N��8�|�<_jV���%�L$.����+���8�(�2��������n�YO^#�V�X����5[�6��l����>r�w��9⻮@�o<������=5���g�0��E���Lۛ	Rl�����Ќ��0Q-4 ���S�B�)��Uq��9���!ũ@E�����vw
<�����i��"��P�Pŭ����+ө�e��zlB��&���f@Ë9�y*��B8�Wh%�3H��^DXpT�>�.RW�M&h����X����������=�=i<\��W�a�TI(= տ/#ę����ơ�7�"U����hF����z�J����X0��-�2�B{����ڴ��M�
Db�ېݾ�H����Z�2�!���'~� ��3k՚u��X�fR��;������0��V��*����w0��$�����F�Z݀l�Q�ވj�&��zC��Q�q�搅A��6�~o� �4XKH�9k�/f��eH'I���a<���L@"��G��v�l�U�Z��
(\�V�:k�X
�q��kc_�|��53���r���u �H��ۚ�42c`0�(�b~�`7J����]S7�Ȏ�^� Hi��ب�w��c �g��F��ɩ��u�1ޠzh5qSq��U���-�OP��yg۫�|�ٖ�O��������9�\W3ꂧ��'?�����M^+�:S�_���<7��G�~�m��FK�K<Np^�*�����}�#G�:�$���O�^?���c5¡��i`8�X��گ�����0�o�UU��{ݴy���x�]ׄ� �$afU�s��~���H�\���hF�a��6����x�n� ��۝1�"@t7"lڐ�#XL�į�j]}�a��A�a������=oZ��iiu�����5	D��}z��h<٦��#T�O�g<d�Ҩ��iP��b�u~�c���j�-(Y�=f�����)��٠6��j��!
纑1�MI°Cb}�آ,I�"�U'`�:y' ɫ�W^��scPWr4c��(�ܣ5��[ ��Oo�}z�
3�/u�ur?���v�{���k�Y{���}���߬��aϬ�Cj��4�5��cj~�I�m�:l6܃�d���Р�n�g�tpxD�^���w��8
�ڀ����8�'�s�5."�q�����@�IOи\/��f��lm��dp9����n	��X��8�.����`����CG�G,�� U��H� ��}��H�^��`>�6K�c�
#�|�������mE@\��6�M���#�ϟ�5�ƫ�oV,T�>ޭ� �ь>*���a$�A��j�C�n�vv�5�-fl��1���6m�R�w�ү~�+�Y��kz*J^]0���)��T.�e\TSQ�n�����y�iC�$ȉg����:��� ֑i���\�����_�������}��"����s݌�v{� ���ئ�o6���״m����A��?3'�cI����$��S@���LCz� X��*cb]�da��P� x}��$i�f<u{��:� ��z�R,ϏR�� ez�h`ւF�V�:t�ުYo��ޝE�c�Whh4�lU1������6����g�i�����k�4�x0�����:�, �r9�E��ӥ��X�@ =���i!��-��f�u���O\�- ���{�_@P���K�QW @ ?��7����{��  ���^ ���ׯ�8�����E��&i-�����t��ǵp�T?7����4�% �H XV��g���c��3�?3��3<����ŕ,����~�#�N�/�p?Vs3d����Qza�ׅ�3��œn5��A�4��43���0
�Z<h�����<LkʹI��$�~�d�Uf
V���E���EӘݗ�C�Zr�/&҆��f�-��ܡǏ��Çw#w�V���gڎ@G�t�jt���_0@�M�5z�v���Oh���N��h��k[���ũ���MZ@|� �5��^ �7��m~A�$��\%�b�ڨ� ׬?� \K8	#n֟Ĕ7�<C�%�f�WJ�� F��О�ۛ���B�`k݇�2>����`xk�R���B������
}��.��-��W��Z\Zdc�ߥ!k�k��g���u�1�Zn��N2�Nm�� �%��5����A����~�oߵ�9}�]_�g�@@�s|�Xյ��>=�t�7�@#*4�Am郿�	 t��1�O�+ў�n��)h~�<y�p��Xx�k�\����"`wϑ�9�O�w�HٵB.vA�o)ߞ�y�<w���A����_�ɥ}�14	S��B
<�O�돘��a�g,�l�9dm ��x��V��1I� 18:u��Q�7��
H�^<��� �f	�՚.}��5�J��hS-z�4��I��e�ꙕ8���5��qu���Fs�Y}��������~D�.��rӼC)"6��X�?p�@F�Ꝑ�����%=�|��n�ӳ�����?��^�ꍆ�>p�� ��� ���Z�$ �b����<���j��+NMl�{����)&&����u �}�C�gFa�S � �3��Rc�v���ʆ���A
v�F�� +AN�Y��ږ�:V ��U�ܺ�9g�W=��\HOޣ��ǯ�_=�k����2��ʁ@	@y�ϭ7�Q��tg�A����={k�mz�*0@��)2kr��1���E��B�p@��y=���O���v�WZ #뭬�hA�o�ʺ*u�����"'j|�=L@0�����O��� ��b�a��	}!� �v���l��O���>� q�b=�?H�}���z�|���|&`�|TfQ3X���_�	��=��	� ߭�� �(;��[��KW4�s����xaUMg䣘Ҩ8�po�`y	)}�o �=�A@�aHy�G��Q�TG� )Gݚ��"��:�5=
���޹��X�czr͝�ѫ*)�rn�w&�(ҾĢ�
���L�=�^�N�3�˟r�;�y��A��!u�����������봲3�!�g���2P���� �h��&ͷ��/��:G+���mq�I'G�4�і��k�i �����rT�>�E�2&����7�8ѐ�jH�^�W�!B3(�PPs�q䔟�# ��P�&¹�'�U^p�EEC�m��K����%�O@��c�f̘�yWޡo~i�׿|F_}i��JӀ_b��(���U���C^Z�{0
��nН�9Z]�������NC.����3���&�K�^u�3�q��^����ߕ�sg�4H�FI�+���a���H�M�A�8 �8��H�Ʒ�G	dw��x���`Z_�|�6���mH�/�����_'�k�q�IUڗ[-��׍��^�Q��+ۗ'	�'���_=���3 �3�t3���dݷ��W��@}W����NxwS��J����0��� #.|E�	�	W�J�Ö1�[�(53�b�ܨ{g|Qt4÷��ķ��LB\�f�sS"i�2I�.��&3qʳW��ʷ��^�Ʒ��� ���_� *"pq�e����,/-����)���_������`�S��Ā�3Hn��1m���2�(j�2��Ŵ(��2n��b������6�1���<�ӳsP:�;�Tc-���
���A��Fq�|QW˘,!�+^*�RG��<������.��H]�d��I�ȾGG�'Y0$�F��Hq& ۶=N���J�s�,�E�X���4���/�,�j �1�,���K��o>�/��17���9�6 �}S|D��}p��h��Ԭ���Ֆ�O��j��ɹ"Hv�����W8p,�(�9�(YMm>ʸ�����2�������x4���q��'ÑS�*O��	`�S�0
��u�?h ?�@��"}��g����"��T@�$�c"�|wvv�������_�>��Kޑ��t�hM˭7���cB��t��\���'�����WF*f����³�s�]2�f �S��1��!�c�N���	W�yX�{Z*�Nw��r#t]�3ɘ�>>��2mP,���h!�ߏ捲w���<��@��7.�Bbr��R���ۥ)��fM��"�T�/�0v)�t��K��Qs/R��4܈�>f࢚ߪ������>��2��~}�����
��M�Ʋ�%s���tگQq�$�/��\�I+�K��[�o~���z�Nw�jT��09��Q��m^�0�[@đ�REr �kˀ���<}�p�~����;���9��k�\F�cj�*5-�3f?5�T��(ן#����ݕ��t&%=%��;H��̰1�~�k�g�̏U����봶-e�b�a����Ӳd�I����H�������~Z���L;���
8FC�Ū�����~��Ǭ�]�3��p�60�q��`��"$A�#X�����s4�ߡ��@22�i��KŤ�`Z�}ΝI���c֌����r����o����@��@��ȫPnQ�R2Gs��%�0�>;;��[[,�A�C	()����e��QA�`k\ ���}?ҿb�0�_�-y~�
~��r��:J�^�n����+e �I[	H?�c��{����\�{��|��q����w��]R�c[�wN��ƹ� ��ilى�0�h� N���;�4����Z�Ϧ�E�*Y�".]�.C>)�;����]�V��{�@��@E�Ẁ�?�m�:'n��!-��E$@V�?�j3QJ�� �P,��O�%��-����orL8�K����ːo|���H�������}��U��
��9����2O��.���{�(�cv�������'�8�aܣ_�hZ_��`Hw�,��_N�����twf��N���X��%vu^C.kl�?������a��g#��h�֤?���/!m�ۦ�]�(�Kvq���Bq�4f봤�W��뮱E��I�d?�/Ps;��ŶpxceP��R�ܗi�6-H�[�܋���q�ޣ+�}��/bik<V/.��d�H/��Q�ǛݟkG�����S�B�C{]X@�5�t���u~�	��R���1�{]�̠��!�Љ���ߘp�e��=��vz�z�F�Ю�o���\ۢ�3��x��K�(W��[��B���O$}��{��7���	�������s�\L�|�ˈ_	�4X�1h����:s�776���7��,�/�,//3�� �ZH�-�t�Ջ��s5|nn��]��Y���F�h����f�����AE}y��s�.�sF,ܱ����A�ۿ����A4���G_4�(W[�I��f�Ϟ=�W�_�����O�
�@5�k��ng ��D)��	��pԅ�O	�����4��Q��`gʚY�ۈ`��EJ;�E��(�+e��R&�� $��0#��NF�ޕ8_�
q�%���P������1wu�U��N^�bs5�0�P��)�M<.�߄��	��
���h���f�q{�9Z� L�t9em��~��}@���ck�hJ]�L �$#�s�c���	k��4o�u��u��ڡv+�A�g�Ч�fu��(�AoH�����Y�Q��ap�-���X6k�����Ԭ/ѣ�{tt�N��Wi{g���tޅYg�	���(`ag �M�&���"Jw�D0+~�: ����
K���a�;��d����i=<�haY��� �7=i��#����Y���=��8}�߅�i�zo�VH �>V c����;�!�\�2kaތ�����/���/��J̜Ck�<2@��7���!�4��u�k�fٱ�[�o��1G�V�x���-�=8��������F
����UgQ�5x�Ѵ�5�h�������Ʈ��"0q]46��gs��a
 >� 4n��p~K�`��Z����'$�4E��~_@DWC+_|��u��}���G+�`��sT��h��q"sC�=_\К^CA�;�9C��>}������ܸ�X�u(S�`��t�T�9�yx������"�^;�?;���@G�]r~[��I@�$��'��m��l�;t�,RKˈh��_��X��K��䢩�D���aD�� �:�~�< !��>&��S��|��;1W�K�&����|igg�	�(�
ۻbUF�gfR	��9��A��fm,����>���C�M8�O5�}c#��[ɚ�
#��8�Y ~�i�E��0k�"=0 ��
R��P-�т�8�^?2�)mn��I��V�IK���,����ԨQ����3���-.4������}d֔m:�S�i~��	�2d_��G�6k?�� )>��Zm61 ��������+��i=���ƈ�M^��̛ �8��%�&�����$ѡ��nvή��ۏm���H[��7���:���7��~����?�C3lL?�1����Z�?O_~��c�	Kw�N+���֨Q� g��o���7�t|2` �0צ��y���f��f�Ce'>�CN������$��ks���1V��Y?���If�h���!�Jec��:*���4�e�xь�k�E��"4v�+_@t��mF*�0XD*<I��~�V��Q�ݘ.��l>�b`�`[�E4��'�cq@��X__g��]@�4��MR���:H�S�X_y�r�^S�׮I�B��s����-{H��ੑ����^,�:J{$���4�?K��&�kDڙnP~�Y�%���Dy���G��>n�$��~��)/^ �:/��/��2�X� ���0����dQ��d�R\����f�]O�5��Á5���Ʉ��ʌ��{0}3�0���ə����HC���5���ɍ�K5���1l|�`S'���㿜ie*�񉐫���H�s��s����]>(H�.J�Z�U#>�~aa�VWc�B�K�	N >�a=�8m��ـv��hs�^�9��.��j5��ڣ� ����P��®IAhs�v�5���b@�=�?��(2(��f ,ѡ��63(����v�Ƙޫg.�����LH�����B�$�2V�؎M����R��^�X���Q1��[&��4K�'+���CG+��[7-��p
E}�-�cW����n�����H�0��t�y��ԤG�l.��;�@UCN��76?�����sd��� �j���#����)��-�6"u�sP�a��IA �����j ��ʼ�`Z#��MO.HPk5����[���?- ֚�Tc�HWF�
������O0����-��8mNݞ9�7� ���B�r���b1o�1 �9=;e�E��:xG�+�v�w�Ѥn�{����(�� �;.}V
nZ:wN��#�|ɑfcG �ܧ�`��� |�ܹ�� 0�;��֤i���B�.&r����h�N�M2�_�ۘ�Rpc��ew��(�� ��l
�+��������s����ڱ��`|��2��d�E,�0�`<f 8i���O�|��5�f���38�)I�L>�?��b�#��)�W�r ��������j@d�/\�D��#��c�';���\�<Gr;��]ݔD�*��1�!�j�@pqi�0�4o G08�h�c�����!m����.ml��L\���?$j����Օ� BP�pd�y��t��s ߥ�S��-v ����	��?��r{�wr�*���OP�Z�y"�˫�v��Yʨc|���n�by+��h@��x�줘�G����k��>y����y����;���i��|��kt�4|�C�������~��~|�I/_�����λ����3���3�Βk5������	�f� \��ԞC
�y3n�<i�#P�^F�;�j�j���z=>��H� ��i�����Tx2�h��X�<f2��l� L�h�EYI���!zxπ)�f A⢆�"�̝a��oh}ES]�meFWC���~^�|�Q�!(����}���4��Ѝ�	<8rq���ѻ�w�������~��.��»����bg������/$���-��:�k�l��<xH��v�â�O�Db� �}V�o��},�� xs�`�$ڥ���w�>k�=|Dg�6�����sk�d�A����˴$f�̳�����<��ŉ0"H�"i�Q��|Y���a�׾p��q~L�o�,�c{ft�H֗��Y�s13���2��Ɋ�5�Ȱ��f�|�]����7��'��N���7`d��N����cz��#�vYY96�a��� ���9��Ç��Wh��gf&���A�����_��06���NS�\��^06կ�[�_�|I�@1N�.'���T�J�r�J�Ea"+��)��5P�S��[���W�j����3bL2瓖k����(�6�[�6l�/�>��G��9�{�@���>4��F�,���.�͛q�?���bM�;���K[;Gl}ګ�`��V׀�s��m�?�������5�sb����=�m>sf,�Y?Iۂ�ׅ�5���	a�cʴ�zo���em>]�.Z۪�-Ӿ.�Vf> ��. ��b�qM��0@��q|��2�������Y����y�]Sh}�D�O���ٔ�㜌�y�'�. �� ����&��˥�.�y_T��_��Ec�ҝ/�c��3ow�P�w�]L��DY>"@�ih}ͻ���[�,h�����F��_��~܋����
Pf�A�{�{d�?q�l���R&@|M���b슔H$}������}��K|�ki!_��MCb��F=���7��OÀ L+?7�Q?���/���~aA������k��㞐r���l_��)�]]]1}sJ˦޼��I�DQ�O�/�0lj��J��iD<Ϧ��D3�ѧG.���bAlJ�I�&�%�@�gyu����#��YJ8���&L"q���x(���~�PQr�<�Z� �����s|�O���0&���Q�o Lc����1}��*�Esb�, fm4�k�J��y�0(���y��OK�/�����nV�k�0rv3a�9yw�7D�JAG��!�[JA���"S����P�5��m.0�<��r��-#��ܞ=�-�/Ҳ1^V�W���Z��B�M~����W���i�]���0g�T|D磐�&Q4�TZ�!�k�=Po`�ЀSF0
9���ӝ�ݿ�43��  ���3c�N�V�ZmN�=<@��^.e���[��uz΂\�ȏU�q������*�R���A>M�n�>'|���1���Ȕ(�0E�&���X�i���`��G���ן2������������*�߽k��e�7���@�I��s��L�]aDU��^��n�}:���w�[EcvS%��/�LHS�?�%�����w��?��O�sC�������w�}G�~�-�>c��%�74 ϵ�k� �LH��<9"ر��_^�4�ǜh*�g'�k�;0#�/���E�L�c��Bz�������%1;�Z ��lH&a�_dh��d<2�v��=0籑���ԊM�>{ �.,���|N~`ƺ��=�1`s@��ٽ�b� �n0xl��m����i-8���,����)s�M��L2b5��2��p�$�b�ӌ>q�.�e��|��|���eZ"����Lab/æ���!@�ՌE�gH?c�'�.M8[�U�@�a�M��
�L�+b+v4��G9_�$"036adׇК�őM�I^�:pz�(EÁ�c��z�zKgZ3�Gp�7���$ۍ�}'J5�j��wgZB>�AD�`׻�qݸ���Z�ȥ/J�x�䎖��E�l?��_������`��� 0�On����\��z��Je���@-���;��g4J�%�3�c.P�K���r�>C�Z���j�]K�B͐W[�4��3|�uYE ��h�竿6��O=�7-����0�7����O���oC�&���@��E�������������p�>d�H�����<es�&\b�!=/2N|c�"�J�T�}��-����^�_�d����M���+�����?�I����͚_(�~7����Z!� �'O*� ���D�J�g�8c�M�nq�p�Y6 H#	��놆�4W���%ɠM�y˄v�QgM+��j"5�|����"$M �b�Ii�C6'r`���ߣ����_����yvv����'�����������uf��lh��o
0�
`Z�駬��ҿ�1�Q�EA�K��|��[�ϋF�5�6uR(�`��i4t�3|',\��1;7"QU��0��8��O�n�g�}���藮�G��9�H�I�u�P>
t2�� �g� "䅙7��1��$P����&�ㆭ��5�d<aX�/�����-h����D>uHtӢF�α6�_����ӋW{�  �"�}E�\�S�?���f��Q����DkT��,"��n�ѫ��<�<�ٍ��v�K�I`r��j�W�
x�+Q����~v 䯍�;m H�
���/@ʛ7o�ݻΟ�=���L���w�̘��E�=Y�_��>�Y	y��H�!�/8 a� ��р���wY\FE�Ӫ`�}u��Q�7c�1wךf�'::>���S����Q X�'�̥8	x&@����h�yS\� ����i�5`�|�"��.�y�>�:��s���6����*���k7�R�[4����� E�����1 ]	�$�W~��͘�7,lͳ�����Y�Э ��E ��8�}k�hfA�+�eǨ���/���ӧO�_��_�o��� �'�����߳���d�/�/�#L��>���O�3 �3�|���D۞_�$Zf}�0,�S�!/�A�I��j� �����A'#��Q�D�j�!����B�RI\tY�����m��t�'��R�9� �8�$�/,�-vT`��a�����f���f4�AC���x�ʦ��1w�g��Q&��a\\�W �6mp���"9�jF���;�S�w��{�{F�6���������l�D���`W '5D*"�*r~��|�#��6�����lHp��`0�t|:��#���F`�!�ɼY��3��g��$^[!D�wG$�����A�~����\3�:�)�z���0����C�[�v��������W��ڔ\0���K��K��� 5��+J8���~���L��='�Oʑ�"��n(5� :��I1��xo���.E��@�~zI�'�4��0��O�Վi�~��@/�EԬ/S�f�k`E��?sf�ܿ�b�L�OL��l��4�:mNqtou�SnAP
Mo�4�֘3�An�g�U���Y��p5������'�P"zg�:^�]k�����i�� Y�-���@�E �쑁Bܾ�I�h���릟r� ^h��O�/� �Qo�V"lI����6!I���_�0�����?�H�nY���A{�w	���W_�����#���X�9=@����w�ހ�w�ޱ����������-�i�g4F�'p�����"eFh��">�[d��3Ȋl�J(9����G������INEѪ5x�.�dWLY�� �`���ٳ紷��Nh|�,���[��l�{�{��#G&+�p�%�!3�0�Ib��7u��w��uM?Fؼ����:�%�?�Tb�R�]M�����Q,Გ�s]��L�;����7Y#QI&c9�
�{�9x;�Eq��h{{�]2z�9j�1@~�~��0㭍8z��?��Y�޼�5@��Z�v�F�u�w������\���R$0 �^k@ܧ��}z�f�� �~��ԧn��,%�[M:>:����t�1�sg��&�.-��-A��#1����P�[�$�R�%XU�&��9	x��YTy�)e �ސ��KI������ �̅:�_m�۠��8:����[�ƈNN`m5�/?�CwV�>���G���ڥ�}�d͌)�-5�m�kP�Q�53��<X5 yɌ�����"6˯�[o-���F�0@)̙��v}�D�FZ��e��6�uǮ�a�:�y�>�Y�����C�;��O��-x�u�M��&�@��!�x)��o�Z����5u�D $���$��6��s淎��c!m�c&�>���*L�5�t�z�&�(k!�����������?�{!L�����gcc�-&�o[R���ϊ�2�3 �)��<�N(1+d�šA����$e�M�B%��T���:[�DjD��6���"*��)"����ǾRY�?Rǲ&T�ܓ]O�͙Lrfͦ��bs-h�9��&>H�t||����(H�����A����ˬ��0��FH��yom�=�0�`��Ijz繛R��T�� ����A�M��;r�
2*P��x�k2���|�{�'C�я�P�~I4�ZU�X�03��c9��������㐎,��Yk�u��e;�����/����0�� ��v���ԡՕ�?u���a��s�5:;���{�]إ���OL��V�zԭ�}������̈d_��o�f<&���t������jy'<Ki{���z��}|o��:ż�H�l�zzb3+�s��TD!��u�=?�ha�e �.=�צ��<u�5��z��f@�V�A����" x��"�7�SF�X�!�~݌e\�3n�tx��=`����vڤ}�O�U�7����li�[�3���-��{] ,�5��{䢏lզ�B>���(j�R�Dѵ�Z�?>��#��/2���_]���TPݿc�<�Rv ��=b�|��|���` ݝ�mx��.4��&p]�d�����e��/�}��_�f ��'g�����B�p9̀�ͨh��sw�~��Kw[fS�s�*�Պg�*J�Y1���4֚�إ������:>�/���!$��r����aZ3�Z�2�T��.3���$���u�D��S�l��Ȯ�&i;+���лH��Vh}m�=�d�K��%�N��'/+ 	�u/G��C��}�}��Nφ������xCg��Z��j1��0�.F���*3���>����GsZ�y��@}���K����0�/�U}4�isk�v ~�r�#�=6�FC^{���.�b'��~<���Y ր[	�?�����6}ppF[���;0�[�<;d�Mh��dO�oh���S�U�}Jo���2`-w�c�`Xb�{��w��z�֡w�!n��(�3���kB�ۢ����y�n�k��nR�Qc�j�/�wGT��ѣ�yFoD;;������:�Ok9�g��όn��Hk���.�}����}�Y�ύ�]$��\'T�-��
]�9e_���T�����~���ӯ~�+6y��Z~D��7�1[8Q������b�3@�5�g<��hק� ��)�j�^�x���(���p���gq�M_~q��~�Ns��a�l4PD�)���X�\�,x�Z㐁e�j�y��>aM��i�����=�T;V}�*�t����<�f�%� ���O/1)�K�q̻�1}9d���Ľ�-,>f�}����<}��=���ӝՆad���L?!�7Ƃ��7�7L��w��2�d@�=f��m���%�l�U.h[��s|Ӄ��`4�~��6��c��3��^�b�͛-zp�C��-Ҽ�A���H�tF�ύ�Mo�l�٘���+슆���|o��D=s��z�j�������Sq�.HA�@e��:�+�.�Ik?�ع�ן����D�wm�OAE��M��p����g���g�{�G��}��DKM�@p@`��� �v+�V��{?L���&]�bN���_f������C�����ն����1����ȺybSSr�(lі-7(�O#Y��,+�=�c���'��r��4��W-d�i�%��GL�9��ڬ�:�X���+�,��+tJ�"�>#�3R�B��
M.��A�����r��K �PDAc�C_�L�gt	�iǉ�o�U��W�_�Q�M�Glep�,�eq���d���:��m���֡��F��4��&���j�)�ғ�^LV�Y��\4֚�^gf���`��4�T��C�7����a���:���2=�b���7i�op|�Rz~$y�D����K�|m��`�>G�~@;�]:<�r4�k'W�;�}r��uq���t���4eC��v�����@�]�N�IK����h�kn�sÚ'�56�0k㢄�B� �,s�A�:<9�������_�����X+ȆA��e�"�{VK`��l�p}��5U-I�$�W�H����/E����� �Z(��~-I�G�ֆm��n��|�Nא�a��jw]<�=æM�(L��̙�]�w6{dB�5[+�?�ѳ���~���i�vw��=�� ��
�H� �\��Dhͽ���=^ D��T\ׄ�狩S�M2�t�IyeW�Lן��g�㚁�4r�:]N�)�&__V���$Z�l�4���	4���Ox�G�/N�� �[�}=i u���qI���<��߾Msk�4���\�j�eD�F� Ҿ�Z3菂�b�5=.G9��bd�X�`��׮��B�l� �1K{!�e�0�	�����{�~\o�4��"$�-������q���>b�@Y�)-t�Qf~c#+�8�����D(f� �;b�� `8��bտ���E^�ns���	.���4#2?���]n�Xu����K	�� �>�p�h�����"�E�M�}Cj�a�����̷����D\v��	�*u����c/������u�����em��/*�{%�7i�|b���X+�KF��y�]��ݦ�f����+^s�~�F�f^�EsM�Lz���o���6�eD�� �_~�`�N�Zp~h�ɫ]��o���M��?��sô6C^?�t���8�d�4i3[�XUf�5#V4�q�5Y�l���/3�cЮ؅�s�bْt��
 [���3T{L��-ڻ҇��k˘T;�4 L|�ɺo�z[4���w���^�k��� ޿�U7��f#cr&��/�_��V���ev�y�=�ӫ7�_Ӌo��:3�+4�a��E��h���N3���5�o='iz������qC���>�.��T�������{X+n=����w|u��g�4Q܎0H�[F��=�=�^+}�K�Fh ��U2�.hi_�|��^���*��r��T4�Rg�=ヹ��䎫i�/h�o�nX�'�1p�&�9�vB�f�A�{��??���!E3�#�"& 8I+a��F	�5��}Ȑ��\[k���%�`���L�d�͙k6xS�3w7U��8��O�MG����.���`J3	��d!�ˤ�&��36�o��͏���~a�D�L?������m�c���e�a�H1期u�h��D�`�V7h��V�=FhMYU���4~��2s'W�kT)���i�:��z\�q�ĤLzv&�'a/����ʘݾ���:�Ra���2��'�GU�ۍhk{���_?���9�X~��Ǵ��B��V�5y#�wS�9X��L�����hJ��o��t������/�������]:5�%2u��)l���ȃ�1�#�&#ZE6�I��-#�'e��^'�W������&�'ҥkڱ�g$�Z���(st���;d}��(�)���ܜ,O�#����ֲ��(��3(��R����ptk�����,�a���;���_}MGg������A0Ř�>�7�7bW�8q���G&� B�6���~����/ikk�M�[�ql�X��ٻ��c5i�tl��L�>/�5��ej R���帠L�v�+��� �{)�\���Kr�"T�ˀ�"p��eW�GS�ه&�ZK*� �5���#�Y[θ�Ѡ�� 4�;�cS���Gf|Z�2� ���seh�u�*����q笀Z�`Z̨���
� ��҇��	����\�&��X�ٱi&����M�	"��F}b�'��Alˏ א����T��E#L����h|"�k����vc*q�DAƌ�o�f"��'	�̄f�H���ƨ��X�0̞'2�(.�@��#DY�����J�!���yW���a�����0D�� �=����ţ"���i��)���g��q�1�e$�i�FMb�o�Fy[h�ٔ{�Uh���r�2���"�X���"@��3+�����̑���u� �@��{�֬�pO���~D�ݥջ6�;�M���b=�!B�]���1�&bw�^��3��5={���p���e{�歃v�aR��m��D������S�Uƌ;d�xAZ.@�GoTZ>�s��S[�t������se�����쇭~��.����j�XOYw�Z�j���A��^'����W^L IȦ��� ��?�4`!H����f������I����9��A$x/��#$G��ß�_���v�kG(,K�LI)$qc��9���eUVe�T�{�$3�Guu]��̬�k��hb���oq�A��ڠGC�ʲ��w-��t:���ᔶw�Ӄ�_�O_!��s��ET�5NӇ�S�"A��l � �r,����e�\�崝ϯ��%WѶ��z�������A}:�Ч.�3.�sOB����^VN��7�6W�h~���xQ��: V��4G40.ʀ�vg{�ǵ ���e�����޲O�a�=<u�$dD�G���q뭮�!X�'�(am�B ��9�� �1�g�S�\���g�<�OEA`8k�a��f�O��*���4G��g�{'��Q��<X�!�T�eV�*��{�6�W�g�C�K���F�����|*,�\����
֖+��+���~�E�?_��t0�Ӳ��ԁ��t4��7�~O��Cw�M�ߺN�=�֌J<��ztp8��O���_�_�q �����z�|�^�ءQ�-�p��<�\79ShVkxeRnK�uS�"�|KM.ܵ���Ԛ�^!E_���d%�.kI��3@���M��NJj��	���CIp�ց���F�FR����L���s<r���s����������ߤw�IoݺF7��8��d�U9�v���'�?�}��cz�xρ�CWޘ��X)�+oJJ�ܒ�I�i�֩��R��'�%�Z�Ϩq,��GBI��f�,Y�  ��={� H[�`=+���� qQz�Mƞl�_(?=z���� u2���	��/?�J�@`1Q����u��fP��6u��vY{�c������ �Q����\�����4�@֪�I5#a������)0�����Ma`�0���Vկ(�,A��	�e�� X,��Qב(�W��ɞ��ɘ�%V!]V�PDu������3;�{��GS�-Jh!Wm�B%Lp]����xe�=:���U�y�gm�u�H	���6�k�͎����R��5����ҋ�mz�s@?<ݡ��[oߠ�k\� �t����pL?8�����g��r0������qx���������[-B�L�`�da���_��ױ\�b9�xIYぽd*������UU�l����5yi����J o����Ϩ�!X�����3
j�Ⱥ��.��V�C�Hm&����|���1M�@�����O��zo��z�&ݼ�I}�N�G#ޣ>�s0�v>|B��k��Gn|��q(V6�s���G���V
, ���$������&�Gn����.� @?��ݹs�#�jW�^6y�+�<�Ǒ�w�EV���Ǐy����z��ț�>-Y����Ҙl� �*#_���z_��GI��)�2�-���&]�!5\�/X�tJ�huiΏ)kCҊ[�qq��7�A"8ΙVIio�_�>MD��*� ��CM
���^�������ח�\H@<5J}���.��*b!��f�7�+��ӧ�]��;z�PP��~�ɶ��`��tB��;t�t�v�1 ��_����!m�8rtm�J�S���i��-u��#�!�@yl�����-�O��&�R�o{;��Bp���)��z�J��B���У-p���7��m��MU
��!�"�TV]W�m�U�w�5؊�vӚ�[QXv���DKt�{4�Y~�3�	{
H�YK�R~i �H����w� 9�x���/�4:~JϞ��_�yJ�67�:�a�w�s�h:�A��GGcV�����~u���pq���-�_�e��ǲ�?�. ��HyZ$�����������K��^!]���\�f����m���>}J�ӟ��͛�m �及����"�bI�� x���k������B#V掞�]��\��ʞ�2$�3��Q��fQ�gӞ\\'��U9/���堣^� V�UW�#������ƍ|�MC��l��yt���l0R���ƯL����fwuZO�h�s�I�Z�MF�n|����"�oU%w����Ӫ�j�k�-�H�wf��g�%=�j�s���ߙkNX�dU�*��n�N��U鼀�I�� ~A��\r�8���o�n`+Z�j�5r �9�Ǉ�r�������������j�?������1��Z�|�gvE�kg�S�m8Ae�U �g]7��� `m
�"H���,sA ��3U�Tޅ��di��D�&�ӆE�$ŀW��Z}P� f���U@����8�.ʦ��u�~<g�EYeeE �6F}LL"��o����"���v_�pcf�,[����9��|Z�����6��.�7�Q������f؟m���*�]:�UwYg�r�Y�r��3�J��w�@�>}��W���P�g%��}e�4�g���װ�~����?��ݠ�2ϊ|8�[���=O�䊤|^�{������(v>�����ﾧgϟq; K��i�����g������?���O�䞄��� ��3��&;XIÜ����+ݹX*u�t+D2�d�O��jO��TYyI�H��^�j��MVn��=�W���_ Yǔ��b��QYm^SZ֝銖�60|��7��ew$�=�,V��>����p[��1���O�������5'(��"�����#�'UՏ�z,���R�t�/��(mmH[[�N��M���\���|��A� |A"46���^�%^CZ���.��@�S����~��m T��d2UB�j ���ʼ~�:m�~`�`v<�ã�`�I X�ƾ-��U�����G\G��Qύ��?_�s:_�A�����$`�e >���ԏX܉�������<����VƲn�Mкx���_�eD�����}��=��ڈ{2��].ҖU| � ����?�����J����@A�es!^��PPŕ\��ڛ�b<t���~��G�/��/���?�����~�;���kr�uº��'����������7* �s����
 _��1!7�H)�3��6�H�	m>�&b�Iw�%���v��+����Wi���V�(�:k���+�i��<-��P2(k�ٓ��"ձ�Oq�v3~���-���h�Ņ��ai�y~�ӗ��nXm��a}�LH�<���g �J;Ñ�{!o9���எ�5�r��	��=[�k�̸����I3Z:��|���{�.����w�y����z�����L� �A�Fq-[��4a\��ا��rMX�l�O۬����>ڝQ �/@F�������-���o�O>��n:�q��j~&�i� K�,�X�>��5D�p�EKX�;M�LUpg�!��A {!�[J-U����۱�YJ�߫(�Js������w�����c�������-��x��w�K�v�W�+:{*)�J}���7gX~�� �����>/���c�����Ǉ��W�y�i���I��Jjq��g,����~�� .�p��T�^X�1���/�����<�),��/,�/�!o�R軮 ��EW2��,l	�snI1�O�r`�EICbC�&y�h��g�&��e�^y�-B�:��	�΄3�?GŎ���C@��ٸzALS	#�<3����hS���F�b�M`�y\/���׼�"����Ezq������r�}I�X�m��"m��r�T�]�F&��秵�ޅk�0ν�!�U���~���� ��V�,.�(�O�\z��O����w?�O?��>�w���C3��X��0�7~�+��#��D,2�E�-hm�#-ϝ� י�6�Q�="������Z���<��+��5�/���/[>��o8����w���q?0�����Xݫ|� T'�vz�p�-� ~gEQ�[׍�^���C�X�^Jwm��"���6`:oݛ�����u ���o^^~���X���3ƾ����'��'���o�(I>Y7].�Wtv��RP>�eW��y���nާ��:O��e�M>W�r ��e���1r��])W"C�:���`���/E��^���eI����/����gk2��0x�A�Ҏ�9ZRdE��x�
 _����kR*�H�h�]��b9���D��#�r^�"��@�zHÝ*|�E[*A@,Ƥ��0�"���X�0Ԩ����/1�=�-�&dxF$�h#>���|�.-���C�y�[@�b���'y4�}��-fE��:���L�kM�������A~����.�����bo�x�Xe��_jF܇��ѦM��2� l@y��)}��Z[[�q���ϭ3e��t��|�6��K�*c=�P��ߦ&MO��QL�<����"�������H�\̩�J�{{��_~I���������Á��S!�����2al�� ��l'N+��X
������:%���y϶��s4�Y��G�y�mV�6�2J֧EH`� K�W  I Űc}��(晶��z@\�y�ȃ&�i�]���C�!�3�x�������|,��"����YD�Z��m�v��5t	|�9�����nܸ�c�����9hS\�� �\�!��\�������+ |EjB��HF�XRd�V~$c�������$N��^fA}:?+��}R� �Cz�#�!-Lᾮܜ�I���#����r#B�k?����?�۷��e~?����f�h����)܄|t�+�$��z�HG���}
�\��\�`5x����9f���^Kzݐ� |��yG�YZ���=m��7��'��{�_+�u���"��B�-�R��
 H
��ڂ#�swS�KŠW�z�Xs\�� -5�Y �Ixe";��8G����й���)��vm}-�f�5����oK�`a��R��c�j�+<T}�Qh�gڳԯzO���kk��G����Z+KJ�6�,cA�2����[z��[ʥ7o����k���Ξ��5
��_����J|K�'(1��XW��f_��# R,��/��%�_r�v��y��pux��׵�^�M�H�#��Z-�u\�'��bu5�.+��')g�L�Q��J����|n�M~�]�Ӡ8�U��` ��ݛ�$� F�X��~�6���]黩S��Z��P���?�ca��;[
�	��6���wߡ�w�V�m>{:�j��& X�N�pEݤ�P�\ =���8�d��`��X��� s�n
Q��3�s�
��^�,k�Ӝ�����N�{�nМ6.XFX�( `_��m ��]ip�+mi�I �+dOj8وl�5���[�� 5A#ڰ��Y�����Y���� �4�������끶��!��y�wLAR���6��LsY�v+լz��/SԪ�L� ei7#� ٣.���"�Lۨb�2ʨ����\/��Ѷ�� Y�O�s�����}�X�%]������IƉ(W���`���C��@M ���?W���e���sO�]di��{@���~i=�Õ�MM���p�����c��. ���y\h(��ꛢg�n��J��|�c�R��r�n.`8fs��!�I@��H�aO�b��	8�ަU�Ir#�V�^���!(ί�}���F�i>V,&����`�7�Ν;E��:9�L�-Wk����Sr|9�\�Z_L�9�1���]���2����ׯ�6�w����W��EL�?� T��1'��*/�vҷ�� u����2�$Bf��47���m�L>�q��2p�$i��/�����!�Sfaւs�� ������=�pqW{�QJIe�ۏ��3mXg����\����8��ZK���;�_i������ڿ�����Y����/����P�ʸ ��h��u�j�?_��Gm���J�	�\������U"ٟ��Z�`#�ۯ�k��</
�X�1����_�2�l��h8���\Ĥz]����[�LY��SkF_�,�֨��ҳ�ZI���GzBINJ
L-�BP�$I�!IT�߉�7�+sf��x4�u���\�����͘�)x���aEbN�*�Я�o�$�uEv&����y�F�/��b�b���u��s�V-T;� ��Q��<�벮��m'���6������J���mO���Ig0�tS����&"���)`H��� �F�M<�\K�b�=5��.k��
��[M���2e뀏>,��-!&(mg�L8���[l �P�͸ۉ%�HO��R�$�M������q�_ kkw�^r��p���F%5����~��s�b�F�`����n(>�"3*d�q��j�+{�,�a8Y��Ά�h�ln�k����̉�u�w��s�F斮Ӡ.�Y�˶Gb%��h��=��O��Ki��[p�~�[|K�V�'�N���!D���9S��Ϊ�ʆwsc�4��a��'O #�D#�� 0�?���m6���߿���|���gr �]�/�nܳX�΋��� ��e$�����e���|�5ZӂV,W�!ÿk�$�����H�b�8�9(� ���ۧU���
(�şt�/��֑#�P"��,�qьG��[+:��l�>�Cp�aAM暅��qM���h�=��d]�lTqj�=aa�FI��X7�Ҹ�:[r,i�{�$��¬5@� ���B���hcK�	��~T%P��D�ؼ�Q?(�*��>�f��v��o\��h.E9]����`�O�ߒ˶b�P��;r�����R��k
 ����֦�=3���EZ�����\�{�|���#*�^��&��/�g�EѤ}�X��[@��Ɓ���2Q�٢��,�Qd�֦v'I�d�c��u{�@Cu4�5�4���R'�8��q�2��)Y�[ ��hS�\��C%k�>&}%c6�^��|\P���<)�k�d��빾>w���9�]e�
ܜ���o��o|/r �|ٲ�F8�g�d5�����y�H�(�O�� �,�m���q��BK	���?o0G��L|���r��ڵ-'���0c��pDb���^AǴ�Jpt|�2&����zn�������U�ǻ,�jʌך��H�_�*Uhծ�Iݣ��;���N�2���ҋ�7�[՟����-���Iv��֖�z}���1�!�xA�do)ބ�����N�@i�����(.nb��| �&|��`-����,�7u���v�OU7ŹVki��^�,�D�'�-&P_�R�{�y�s���VeՅrцw=���YfI)I���l<�Ⱥe\�d- R��euť6*ո���K*SU~5�kw� ���Qx��i��k���N��/ky@����L�����&��|o��3�
ei�ղT��I�<
kOeIRW���K& ir[[��������&�o��:Y��;��&�]�o�F1�4s�jw��q g��-�|�6_om|'(.[-�����aж��9)�$T�eK�x�({�E"_���u�6�R
�����+)����'�o�5��h�#:��%� � `H���U��}�����G+T�,�;��+� do5ʇ9�]kA�+ �X*,Q�ڢ�-Z��g	�e���K,�y�N��Yyf2Xе�kt���t��t�ƍ�x(}�{�}2E:WN�g��r{��>|@/�?�	EIH#����j�ݿ�O ���[���es^�i�5K�)�Н�t����S[�2oKʲ&}�
�yM~[�I�0�F�%AրQP/�mM����)���M�0�7���%�	=�C��j�!��g*8����{��;��>>j�BԹ�_=��F�X	c�/�%�X��U)
 b��2�|ĹҼulp&tY��(6O��k���Ih�J	3�ur^}�qK�ys�(�v��23[@g_"�v#���+�x�)�U�<�\�P�������Ǘp�流'���Pc��ڰފ@!��؃4��x�~����-�.�[��v��]�Ƀ��"H��ǻ�	P�I*�� �T�V��4�)�s.�kN��	��>�c& ]�U�MH��C�Mz���_I[7�����`������x�TZD)o!�>Ԫ�l��a�.���y,�R�c:P��>����W�(�1�����\��SIA�
>G�uM+�����3�-R?m��1���L��K�f|$�b~������@�,[@�U\"d�C/�㋿�q�X��=�6�n��Ѕ��.Ah��KĴe�Q8ΒdCG#�W��ߢ䵷�nnl�[�ߢ{�>���SΫ���M�јzfvO�W�I=� �𚣽�#~�X����%	{K���G������Ѝ�ޡ��c��~L�0U�� |�zw/&�+p��@PQ���aP �x�ҍoݮm���x\[J8���h͋3�Q��6��O:κ�\N,��GJ�E��x����u�[XF5������N�p���Vj��`-F�Bo��8a����h��C�,��i(��f�r���RB�	��qS��$�)��G@Qh��첀�.���
v���y̿�|J�`m��/kU�v��� ��6*.m��]%�����jب���ɮ��f�iQ:ť5,c�W�.�����'P�ZxDY�^��"�z��n��݃F�*��j?�?�����?�,�j� $�:j]I<�"�P ��S�>���0�ٳG��s؛\I��B�!p*<�LlOÀ}F���i�!��ra��`��ѕ�~bC/�Qyp5%j��|�֨�#�v~�eX#�����=3j�\s��Db����.�� �6��,��<V�6�k�r���Lc� 5�iW��%:v�~���a_/"<#��E0ɗ,u��Ms*��R��1���[[{��h4JW��%�Dg!�{70o�G�zt@0��g��`� �޽���N?��g���ӗ�t��P��7�
�7{}l�Ys*���5�q�&���������|C��OXF�3�2Mܻ�iwoD�_9U����Y"���*���O��aK��� ʝO�h<��=��On�S��m�6������[���I�^�хb�.2k�������J9����c$eOi�pL/���:SO���6Z9�	�dy,a|M��0Sw��{p��ƨ�M�şJ,�Ya�5��"���V/��"�J�>�	�Ab��7i�{����'��|%���cI���@̋ʣ�/YR㺪�pu����
{S-���9��Ҳ@\�eh,�ta(��)D��-��V�h�-)G���^i���+�gJ1M u/
D����Ӭ���A�T�eg�Y��<�J�E`��(�*ͥ\ߗ��l�K~��_Y{/���"� t��&݇Z�=+��ג[�v,V^���tC$�n�"��x�OZ^`�� ��g�}F?��O�{���n'x?
HS���OZc'���8 0"��,M��߮��T��a/.@/��=,f�4"K=:�bp^,�����ݼ��@-B�:^'���@!!��:�	��Nm��`�������M���r��h�Gw����5�&�v����O��}�|��ʥٯc����W�~˖^Cp�ؠ��Kz��<y��1���IH��'��d[~K���Ղ�Ʉ����Y��pL�B��z�_�Դ�{Hx�Ɔ��O]�L��g� 8�Y	� m���7uo���ܢe\y�����txt��֗�G��ď�����Tb�9�t�9۾H X֢��[�����D���� �Y�e�7�<��j�V��% ����M9~��2NlHм�/���2yD��}*�o,J��X�m����冚�[&>@�W���,
�:0���q�X�h=��U������(3+D7�I��q�XB��@��G�aBv.G]��q��-8�^��Q	�.��h����ˌ���p�|@o���Wo�� XJ啞�I�fA�o�����石�4�_-�n9@�����s%�AJZ����[�良�2T�J*����6^@��&-N)�_Y ��X`�G7�4��䎎h�-�[[���I7��Ӻ���	���!��i����.^����v_���xB="w��L-�|��~�K_�uHFޙ�������Nh�]�7���b{ρ�}:v@ʷYpݒ�#��6>�*�2%�S��Dem�	�`R�=�Mp/YTA�4I(	��f��Gz����#����!FH��bU�<@��Űrc����v�i��� Dӥ�d��ĕ�����=�U���w	1������2�y�)������� 26�r��l�3n�ME�/����X�W&Sy���V	h& ~����?˭�TݸI�8��-����J6�@��LqZ'Y�mE1�sį��X@n���\_[�-�f,Ȅf�G��6����x��EzC,Q2!�C^���ιC~%��\�,�E p�� ��Ҽu �[�OB����/8� �֭[�[�k��I�!��<��͛l���m��H<@�!e.,��H�c]�r��l�噛ܥI��]rr�fa'��b�֒n��	M'#�66����No�ڢ�uD��0s��po�+���&��ޅ��`JGG���������3� vm��s���"q��A
��d+����"0V��su��iLc҂���:l��Y�&h�O�	d��Q�L�"��c�<3�Q��06���ǋ��Px�h{��w��vM�ʿ�����9"�Fѐ���{,g�GS�S<��۱^��9�u �ϗ@�nt���u�d6]v۩�����~����.�S4�-E!>�_o�{��g�+n�J�/
�P�H�xϭ���8�@��I9��������s�ZU�[:�hc�eb�MX{�}��;�!��̛ʹ��a
���eP�e�yw�SK�X~���#G�'�A|�gZ	��Z_�ԴW�� ���Hz��}�k�+��ߗa]���p�4MW@��H����湢��J��ӻ��+����osÎ����8��G"-�5:ER	�u�@�q�XE�'|$���W-c��`���Q����+�2���],�H��l������TN2��L�T[c��#@��v0�[��p�@�a�歭��QҼ�B�<L<7�8-λ��yB�^H�m�A񒃾/o�� ����X�O���zj���7��@sv��b7�E�Pk̂�T1�X����Ra�q��&�Y31�.���,���C�{<�Ǯ���c��`�QAAMK��R�M�:h�H�{�Z���=�~h��5�|����Tڳյ�k���sk�2$���x���g�;
g5��[0��y �דp�/��.���.ƕ�cpC�ϔ�ˢr�/�bmu���reh;���-D>�2�"a�Gf�!:�r\�K�N���h͠��(׎���
JJ�d�P���rA�Rn ����ި�n�yMl�/2�ݢ�U�g��b5�,��s���pe.�
<�s;� ���� _j� ��X����\������H�����l�m��ދ�dem�?�����Z���9��5���*��/ �J�� r�ui��-~�Ɵ�����v���%�4_��oٔ�0�H���T���9������}wm�@\"����窿� �[��IbErYup�"�.{��~�T����
;
�3栗��)U�
��˚�ݐsT`{Mx��h���V�E'30��k�b��MU�n�s�Ό�[	iRN��IO��rQE�	�z�ERZD��d����6� Hqڑm\�<��-GW���q;���.�!+㘶�[�JLfQW�+�N�,�5��s<�9��=]n߳U�v���E\���T9��g�+�{%�q��n�V����dm�aN���&&�)��l\���8�C����ϧ�r��,���V�	�$G1�Tl�c�a�5�q�_w�q����5S?D��ǒ���}2	16��8�,J�r�ٰ���Y�p���Q�&���`���,�Di�u޾�\<Ѻ�Ǵ%�9�s�<M���f!��Wy��_,����|~��]�gUZ kwfg6�%Y��w�|���<��E-�:p�@��v���K^�B'N�t^4�
��F���./��Ԟ�.�bBaq�y�f�Ȭ��z?�L��@H�:k�k���ݧ�����w_��A�Z�t�z�j�?����t��-z��w�t�v�� �4������1@4^aPy��x�'8/{}v�RniK�A�S�SNԑM
�$��Ca1
u��]�:&��u�1�(7�� u�QnJ�c�����k�hK)�,�ߖ�xAM�p4�A�\_J>7mi�R���˶����W��$�\�P�S��MI@cT/��E�VE�1K��I�mIj0�L}E��< <���	"�,��E�����x���^�X�����k�� ���>-Rr��^�mm���:�ߐ1 %N�gj�a��㽾�y ���X��2�˰��ځC(V�a�v٨�M��" ����1W�y@b���*�����(n�1e�4�I^6z��6p�-Vװ����գ`
��&g:�; ||<�-.GG#�R0�\X�Ŀ��`i�~�����pc�P<��)�J�p0O����+���R�]�����A� k�Uc0�� �]���������=J�k��s	�I��w���r\<*�R)�
{pۀi�@�nIg��(���y�U̗����_�6�z~��R�}�:���li�ր��vr�Rh����_�أ��^����$*��A2"Cpe������5�8n�ֵu�Аߟe��@�
 ��ܹ5'����������L�@%H/$	������Q�������G�1êDz0-`K��:#k� �
SO��"��%4�k���A�K�)��-�O�o�hcc脭M�v��6Q?����Q����ð[< rt<���}7�&�����V"��Mݳ�g���o�>t����۠���rח�eJ��y�X��יJ�U4�]}��W�W��3�{�Y@;�z���L�<�j�ܸF��6�u�]�6��!f'bA@�:e0Lbq�9t��j�Lu��O�������|��YX��0H�Rl��gD�4_&N4�z��Qa�~��q�j�Vy���5���7��{��߽E�7�Ɂ���o2�{㼫�i�͸��=pyH/����o��
cVf������sjuU�� [4 �zY�-�4y�=u_��j��)���횦 ����V(m]�眖��r�Ů{z��忒g�>w�/����t~�2ڮi �,��w>7��"Ts=Խm
�e(��%P[��́U�ua�׍V�։BI3(Z�O����ߵuh�hĩh�������5"�c�m�`w2�h$���֦o��h�>��c��Z�SA;�߈�]�F�w�n������J����s a��ې���� ���3�=���O_г�����3�,�[����LsX�9��}/u��h����Mz���t����gy�8	wyQ��%DQ�)�����i/^��Ç�\���`�!�.E{Y�1�|>c/0G�E4#0y��:Zʥ�T�E�{ e �_�`�ө
���4��㚜S�8X�\[YmǺ΁.Z?+*YC�q�;�׷苟}F���C�}{�6���t�>G�3
`���|�F�鎘�`��9��O������s����oh���G~߇UJT
 ���1�v�n
M��%,��|I��f<ѱ�qkktmk�>��}��_��>x��'Gn�� �N��Q�nV�|5tx����1����;�m�ww���tm�S�I��IJ��#�Ģ���]��V�b��~D��$ѱ<(�#!^2 �|ztY�`������$�sb���u�`j����.�OW��໢�|=/y�����e�v��6kn�b޽%*=[�X�Qgm�͕1�XzK���I��s��sĺ��WU
̣�,_m�����μ|��:yǔ&L�"������\XQ+<{�,��v�7�yǁ�5z��uZ_2���^#<	��ǎ��ݠ��ڢ���S\0���z<}%������AEם����w����9��gYH1���Aw� �!�Vy�9�)!@�&={qH�S��egw��Ga�7q 
����<5S>2M�wd�Q����H�����qr7��t��5������Oߥ[o��n�����=afv�F046'���	
���}��	=�M>����7G �^���[+��j*Y�=Nf�ߨ��L��K`�޶
���.����������*�(��<a�2Ϊ��1I�.[��;o���C�s��6�;w� ��	�������V�p���x ���`�&����uw�"/`�ح�G��cE1��K�X�7Q
/�
߸�4��~���b^س�s��ݿw�>��-��VZG0�uؒԬ�^��ֈ[��t�k�!|cMƴ�/����%����FA�a��L�
.�f�"�9H�����~�&���z�E}�$�
�e���a�9���/ �V���k�*F�+:}j㷹�O�����Z#[�L��z��L]c\ϋ�zپ�c�U:W��:��1߉fe��2}�"��EȻ�:�=o���}�O�Z�x�&=��[:	�I��|�Mz��x���ӳgO�����&�;����Kfn�5h���r�_�u�ό����Mtxt�{��G#f@W&�COFN����!A������K�(���9u�>��.}�������}���B5r�z�5-L��6.g���}�!��A�ߡ��}z��%��3�k��Im�D
�Z��^�4��ݚ4��̙
6��s�FE��7h㵵å��olxa�{o��}�:7it��@����z���BxNȂ�w�cp}ߠ�cK�^�����A�/���,zQ#��C�����O+f��63� _^a�ċՒVù&V(wZd}�r����Zg!w	�'�N������h�.��x_@iZ���cVC�>�=�Ͼ��'n���^Y�r����f�Ϸ�C�)��c��e���q��a߯��9��@���eh�����XS����`_��=��}����=wν+M��}���h�S���f����z���ĵ��8�k�GWxw�yM�#~7A �	F�����k|�+Bf�hNVⴲ%�GT$�o��
��$�Y��D?��ɓ'���K'����:�n���.�N ��{�wIA{R ��ans '/R�!"��ITz�U��s��Z�;l�w�zh�e�T��uV����./�YY��m����L�wZ�[�T(���;:����@,���� ߾}��z�-��Gg�����#z�������N��.��}��7�}7��a ᾵5��W �/_�����ޥ=�wݱ����=�f�X�a��+T���u����� ��4��t�e=�� �cKS�	������Ox8����3��:���h�d��O�r��z4��M��I�N�2�N}ן��}��}{��}k��!`�Xt�[`Xd�~te�z���ѧkC�6���B~��������k#�(�~��[��`g�͡�<��{ l� 2���"M�:c���]u�V�c��a�@�8X�rW�.!�m]j���6aEG�os	x�<��.�w�g��B��2h��XX;'���)[�:�,�eXr���8q�0�~G����)���cˎ(��z��خش��4�;@
�eex�0�U��!٩��t�U���j@Ac�>n���` x3p��T���1���j�Kϯ��㠕Qio���+:ӫd�kTZ��1�>R����ƣ�V�U�R}��\�<�8��)����;��ox����`MW �դ6 �)_���*<^�A^�2�C� ��{�.ݺu+�L�c��-[wm��>~|�uM���� X'� ;�Z��s�Y��ӳWq㴙��c(+�D$.v�_�΃9�p��74��_�|�@�1Gk~��!���҇��ѯ~�K���G���'3#8��^�Qb{g�<��}ғgOigo���]�Ϟ���!��Ş��y��[��E��Em|��wG�G4����BZ��Ĩ}�o�9U�e�}��Ak���?pB��;wL���HeX;��"�~��U� V��%�#/�ښ����X����N 8�d��	N�+���#�0�ɀ��w���}���	���9�։Kʇ3� �`4�^�]���oio�67��6� ���I���6XRв�,r�{֋��~��Ս7��T�J�Qc?���^	X�;�_�"���j�^X��� `Xiǜ����h�|Dk��5��0�1��װ�D6l�a[��>!���l��U��!w��8�}���**i	�u5�Qzm����W*��Ha��u���S�PxQ�U߿�o�o���]�',�L������+�J�>�3���#y4�c\w(��R���KU��wl�p��YBJd���Z�����Jۂ ?AX��_�B���o����l��.��bN~��#=_�@_^��� ��(�ݥD�ycx ֊ �	�s�����B��?�y/]�Vr�B����3e�TKgA� �
% ��ش7U{����L������z0쁰g�X��� �-�Z?��C'����e,���n�"��ԝ���������A�ό�����������u��Tx�~��u���1p~��1���>qN��Zp�@^�����+��YX�d
-�U,�P�JI`��S�����,����&��) /!�Rm�+pbM9��i�/��o��OJ7,�pvd��<d���;�{�Y�ou},&�j����y��r�+䪄d	���?(C��QMg�q�Թ<�⚇Eu���O�8 ���Q`��i��ţ�c�������/ʴk׶{!�������gLX�L�z}�y����e�t�"��|�����h�sТn�R۞�V9��_��<J�x�5:^�գ�>r�t��aN�Q^?��ƍ�.3�0�ъj�^��ҋV_��DQ)�yE���+�y�d>��Ӡ�����	�P�2�������<C9lm��Z榭����Ԏ��y�̉�k��z���Rm5
��W@��Vr�D�I�QAy56�"�$�7��Id&j^�縍�w�+���<��+
A������#v��%{���VhX���ԟ;	 )�ˮ<��FK+q\TZ�4?��m ��\zF�2�e-�������:�vK�,�h�v��W��r��[<����70g���ƫJm�Ӳ������Z���{yf�yO�H�nF�|�������Vd��V�GY4)(��\}%7]�����3 ���Oy��cJ���{z����/�&#�Ql��Պ�I�.����tG �~G'Arb���g `�O�1��&ɚi�@R�I4�[����&޻��+��MÞ#��pO�W$&�1;�������=r ���PM��'c��=�nb�$�h&�'�X�D���B��6bz��VآU�y��>��OI��S�}�c��VfWbo�lz7��-�
� ���T�ΓԂx���[�"E������4i^G�i��A˻% �*������[+��c=���%����kQ4�t�UP)vA*�)��~���jik|�u��	�7��w�*~��fUՌ��&"��~X��G�E:��1(���~y��Kh�]r�M[��)'��R�c��z����	���q����<䆽�Xa�6�$��V{h�SE.󝼲5xI�\%(�E�c���:�
��������P>![0ѷh���C(�����q�ܿu�����\	����>�y�k�{2��ǵ�τ𩌚}�䦮�� p�,Vޣ���˖�c�КxҊ�.�f>���e�L֟F;��h��2�\�Wq	��e-���cn�����M_��	���O�gz��Y�7UofN��|,�ϯ�gh%*����w��}��׌K�� ƥ>zr���1xG�_�^) �)X�ɻ2AP��HV>���｡��`��� �:<��c97-��&g���54��t~��[�|z�\X�x�|3H�{�>*3/�l�s�S�B��	�Y��"��rU~��"���B�����s���~�c_/��� ���7icO@U�k��u9�[b���(I@I�`+��`Wg���g���� 颢]̐�Q�H�W��d�j�͛.��� /X�L�g����ޓП>*)�U�h`B��r�������<�(�<C�
�N!(]��t�Н9*�)��b�9c�4�������9�����^y	�1��Xc$6�t:F��eU3(��#�Y,�K ����>�3_9~�͚�)�
9]`�`u��M�)]3+��5ք1����<��-7P�5�Ϟ�|��)�����&~^�QQ)�z�D���W(0c�I��!r<%� �E�DUC#�KP�(RE�D!z1�Y�+��Y���jU2�"��c}�Z��O��(U�����j��g�$��x�苳v��c/�����4�k���|��o�A ������Y�/��R"��]��_&j�rѼ)O$�ͣ��|~柘1�e�	 �Azn��z^An�AF>��� �g)K���4��+�����߻��{��޺�Iׯ�hs{b ҰϑYy��5�~�A�GSz�t�^����5�ĕd|��Z[�+6b�����r���c�����y߯����>��n\� ���A�t��/��� ��O����غ;�R�D�Zi0ȵ���ܰ�4����X��N���_7VP�J��<$ G�ƓD�ט �dK@�MTC-���:H��Y,�u�����l�-��E���t�)y���ٿ[��\��	y�ќMzeI7���M�P�� /�R����C%Ͽ�L,X��Z\��3�?A+�<C�M�CQ��e��ka�����E`�r�X^W�R~D���.�H[�䣃��6i�s�f�[�$>�Q�J�U%X/!�sV�h
�� VM�\j��ű 0�� Xe���R����`�ژuѱ?B@.ig#���-�L���ע<��I�)5]R��e7�7-�PC�gX!��uC�0)c�Dz�� R+]�y�y~_}^��*Y���G�=���N
��{���D���MI�����w)
/�B��J| T�v�qLTߗ{~�C��G/^�9�1 ȼ�H�����m����h�.�揸���v�e� �>���ڤ7o�ѵ͚�4,�6�_X�j���?�9�������1MUj��������ҋ���{z����$*4�a��-@�d<�oC��5��v���z��ݖ8��+��k�Òߋd�phC�`�Z��W�Y	2V|�����,�ܺ��2��M;N�bN��zr���<hX����R�g�����o+e��m�'	K�^����^m2z���cCх�|_������
��<� q�\Wްn������,�\o�����z���ٲ4��5W@�GU<X��+0�Y�JV�y���.�hq��iM|X��2����w	Hr���{З�~�v�k���b�����S��*��-H֝���%�O���q��X�_̮�$�!��#l�<� W�RԯiohCy���M�&��ƽ�6d��D�R.k˳�(}Az]�� p���ξ3�-`֯�2\*e��^%b+|>����d�K�揭|�V�.ʕg��6�_��<��7��O��e猾�4�Ĝ��~����5����wY�p�8�ݐ5�� �!KH�_�%�0�I���\\�TL��c���-��{D1�V�e��Z��������i�`c��7�ҝ�䭍hЯ���Q$�`�7�3��1���bh�hD���Em2�5i�B�߫�� ����0@z��`5�8~px�x�ߛ��5,��/��Y���:�X8H�͛7��kt����M�s�Ǟ�TO�u�`��EK����)��҂b�pv���j7k��<i75�)4͔��-?�ݕM!)�R��˹�^�dK��1
�����܈�.�"�۩��z	��C| �/���>��c^�@�������ݺ��`\�ӟx�R���8=�݊)�^��`z���
�iԮ�>�~��Ik�5P0���%��Wj�˔�unQ!`�k��@��l)A9Vܞ��NF:3�	je"��fs-�0��،�Q9F4��¶�|�/�e��Ē-��J�%*�Զߧ��+Z����R.\Vp�-���Q\����?�9� /�����_��=� 'D/2d�qH�Q��g|d������?����qRƞfJ�K�۵�|V.�le���s xП����z�l�o�#o������BAnMm �� ���;���G�>m����0`EGCӁ�oXe��> �x��׷����7��;o�����t��8���r����5��֛tp�CZ�X�m'���0� ����#��*�G�\��$8��4�ga6y!0d۴B��!�,f� �c��)�N��Ϙ=��Z�}��1q��+�4���]/
����?JV���a�������Ν;�����0�+ ,!� �7R������iL ����{�4�ZlA9`�`z8&��y��@����E�H'%�0ɏu��v��:=��O�6�.j�O��,m��5��x�Z�s��VΨ����B+aKe�5̷#E�(�1�����%��%��o�	�Z#��y����xq�I4e!?�w�9��ac���#@�Og���gmhX�{5��@��L���{iL�c���=z�%�z[��)���wP���F��"�k��i~�(����)�h*�Ӹ�|���E��i�U���kI��9�sm�+���_�'�ِ���k��+ڭ�l��� �"W�\�Q��ɴ
0�T XhF����������QX{����1�כґ��WtXzT#U@5�h��i�FD��|��G0lI�r��@��@�Ā���~ƹ<���� a��{�!�w�}��w���w�q��&ܽ�m3 �z�����c�#��ޣ�o�b�������C��/_�����a��=�p>B .��%�Ε�OE�^-��4?�iPA��^�8���g�Ϗ���ƬU����|Ap�k�_��=����a
��b��H<T�F�«5�:�֞Q�W��e��)�p���ŹI�x&�� � �LJ��H�����������+�:k�{���v�D:ߩ���^��-�O\P�;ja�U�	P蕿K�*Ņ޽>������C�X��v�/s��>���v��i��*x�H��Z����*�����\�4O�˽R��Q����o.�p�Cq���^����[
����}2���Y~���IƱN�İ�j��&Q��=�������׸I�=�zQʁ���2wOB%˜���� n�\qX�O!k�V�.3NJʠ��']ʮ|��B�_����_������y����8��
_�y~�d``�:x��-q?���+-�U�����D+/��N`dC���z�V̑CnA�,���|�g��9�KE>2.����4����(� �@h;��W�<km�p:B ~,߿�>�w�676�=����m�|F�A��꡾p��(�T��C��۷ߠoܠ��NA��[�U�We~�\���aO�I[�d�-�ό�5[z[��i.8��+ؙ���]�x�Q��\ �Ϛ)J������8�k�A˞���ߜW�N%we�E�ߡw� �g��S֮>�l�r�ˀ�=�Ķ��r�H[!5��n��B:7���o���0<00��i#��E���a�fb=�{����c��D�`�VЋ���룒ƨ-/b�EM���=�%Kx�N��etk�еJI�M���ʹ>fM�����pKEb]lٲaC�wx������9PH'^2ZxUY�2�Ȇ�Ed��ޖ-�������J5��Z��*��=����cF�6��z���eymS�t��E�}�{cY�8��t�d��k�3����_���D_����V ��(L�!__�g�e�ByM:��zyw�]Xp�����?�o�fO0(�E���㘗rpL������x��{����_~�� x�/C� �/'��w+����{��-u@�ߡF�G��k��g�g��?�?04n}�v
�=��R�����Çcp�C�KV���4��;o�ݻ�; |���/��5%p���Z<�xz����ڐn�z��}x߁�-Z�X�ͭ͸����ƓiR�`a�?8-�99�aP�U��3EU0�@�?���5�Kz�D�C!I�v��J e�L��nK�܆�o
e���z��*J�?Bߋ����_i�gϧ�����.�W5��P6���&�E��W'L:�ҩD��KS� �y����I���o���1��-X��,�b1���8'�G�@K0�%"ʅwͻ�K�7�JC�"��aO�y�@wQ�����,o��� ^�oQ ���
Qru����4�ϝ+hk�A!ŵQt�ރX!e�o�j ���t���n^�:��6�c����6�a��r)m4S��VZ �᯿ת����I������4U�$�K$�p<�j�}�6K�x��(�)m�Ep��(�*��6�S~��oR'�����:'�%:�ܻ�П+�.�z�H[���0V�璀b����˽�}�[��s�~̠��=���� ����������?2���Xo�Q�W� � �r��?��?qL��?�����/ɜ��T��o�K��d"S ,�"���7��:ȑf��m�=K)"A��o�v�Qk�=�4�¤H��HL���:���7���[�<�������nӳg?��^ �~S�`�ڧ�wp_tt�����w�������'
E�S���[>2tвG5��Z!}���gF��� ��
]#����2rI�Y�E:���?�_�jL;s�L!�Pn��&�H�[4@8E,LyEj����bp�������/��$]I=ki��G�tyZ$|C�Z�-�n�kX9w��=��:Y�P��x�h ��iJ~ADև+��]��A��EQ��)��v���wh��~����.:oD��v0���WL���f�b��J�c����rF�ؼ�P���_���͆d<�g���4��#ߪUk�-t�g�ҳq��+���G�c@]��� `���D�=����s�+9 ^K���<_��E�����V���z�>�1�g0x`�,hP޼q�����O��Թu~
�y�J�W���I���	9���E+�xE�*n�ڋJӢJ�Ӣ�2HAA:�m���ׯѝ��0��<� V�
�o��-Lh'�����0/��O���y�J����6m/�6}�"Pŋ��]�>����V4��I,� �đ"�8#�[���'�#!7���8ѻi&���&�	�R�?��Fh�6������l�fTO�V|�7Pz>�k]�9`Vs��l(,�#7O'�����D
&|x�%�R-J3�xkc+4u�Ji����'aZ�����^#:OY�[�Np�����Ewg:�k��(c���^<Y�'!gpN��s�,#�KY7�,(�L�b�~����z`�G)0��F�\�,W�����Bک���y���:�}���7���Q�B)
te�����Q��vҊL:��5��E,�g�8���o�:)�'�u~��"սm���n�׊��4O��-m4��a^�]��Gˇ~H�|�	[�����9p���=���	�J4X��'��=�/ �V(a��Aj@ b#O�U�g����m+��Ef�^d�f���Ǟ�����A�ݦ�y����ӵ7�Y�0�t �D���1�s �A���&c�&=��}w~�|hWl���A����5 �Ʊ�W`
�f �b('d��Tq� �B-�B:�m����^�;[����{o�r�{�92��a��OkdzCZ۸N7n�Ak�C�J,���	�ge�U�p[����åW���l����3U�m�x���UG���DI��쩾��v���ytq�Z��	{���]�����\|pL`Z:��( ��>R��[`䂪����x�O�S��i�ϒ�{��m��w�i���܉��5I��6����`��m1[C3�ϙ�bik�������Y�]j���7,I3���?b��t�`-'����<�(��Η�/2~�]��{���8�=~��o����G}��&5��u���&ުk˕��d$c��]�'(0�}˥X*��8��m-����9�<;�EHmwe��w��!����(�V�K��#h��Uρ_Kc�����]v�o����=Zs@�v�Z���'D�C�9�ka����4:v�y:r����;�����|N��	�P+	�*���K`�`o0ܣ��=u�Q��� ~�7駟L��۴1��z2>r��82WǪ��Y�j��~o����s=:���p�F.�8�j��
@��;��S^�]] �7�����������9����D�W(��fCT���+:)�=�r�@@U��X�^�@�����A��"���b�\���Y3/nS�% ��6���\���Q�v����Y�2�	��/�!����S\�#U�ա�*B�e>�g�S�J��7	�eO�@W��sgM��r�޶�Si����c��"����|��o��oy�$��-��Z'��
 _��S� W�/x�g�ƐmA4�ȭ�g�O����v�"V`W<��q��n�k�}$h�����tipN�΋��[[���yxhi{gB��@�p�/���p{��ݽ1��ܽ��am;|�8accCc//�2DL�uB6|�uǡ5��(�N����PX�oܸ��ݸ�s�:>�w �����w��&ZwB��{ߊ��'tp(�xՀ�}�Gn^��8X��۬������k��:Z��HH?�67lm�c���d�-�~�YuhE�fXC'�A�m���D�ԡ��d,���
�ٲ��w�^��x���>#��i��{�ԧ
n�&Z�/�Hyv�n�h�B�~T�.#��v? �/�
���^U@s�:	�o��T%wȠƘ���ш����8�{\�}꼋�|��Yh��Y����sIm���8���ךG+J�ޘ�w����fv����^�f���Ȏ��H���F��E�i`�6���6wD�}U���N,�H9�H�]cċM�E&OB��P�9�\��Q}}SӬV�Ӹƨ���m�<���tO~~ 0��b%�����>_|���r!@� �X�چt}):��t�OFEo)��x���4��3D/F�B9����+>yV�E�nױ.w�/K�_	��u��~p��,���e�q�� `P��Jǌ����iL�D������F�0��Ood��St�������?ۧ�/0t�:�h�	SiP4�LlK�t$@��/9�3\^��8������k�w'��$��O���#��k4 &N��������ģфF���k8o�Ǯ�:Т�'���-��{�Z��a�<X�b*"�k���� X�����}ܐ�=��U���"c��ZK�.փ�x�3zJ$u��Mm�� ���diS �A����7t�����cQ�tK|��~���k�c%���@;]����z��\ϻ~�9_��퉋����ȯ4>oj��3q�������g�kuX���ȹu��TkX���D�q>��.�Kݮg	���=o��<_��]�X��)8(G	���?B��#�n_����K5�,pgw��^<��R+ �-�A�$٫�ߡ�<�l\��r��*���+x(�������o��r(����X�d
�Ѡ��X�U|�/�6ėF+cRW&���v�.k�''��".�zL�%���9�?7�"Y���a� (���/�� �zԽ1���%��W�=�u!����xz_/���7ady�������<I�+�_��3-�&��ȶ�;dN���0~~ȍ�p��W_}ņ���4�^I��~/��Y����I�A� �ց� 0C�+i�?���5��1����6���]�7��;�Į��
��Z��1�r,jx����C�e8�9-��z� �u�HJY��˴w��>��d߁ZL$��SX�}.`o�uy/����x���1�j��%h�:�?��vy
B��h� Є6� j9��\�Vl��FY>�[^x�V^XW�v��1��8g/M� k
���⤮�V.�����My!k4_���k@8޶���għZ�'��&$�V���ܧ����I G�,��Lhw��r�^U�*�����5E-ߒ^��u�JjN�ѐd
�V %$`��@@�W&�_�8�A�"��(��&�?ud#�cxt�6��O�VIS�z�1.
y��
��t- ��L�;䢂RɅ//���5ϊ�f�c�����	��c���^������M"�!�v����������	���2���1.fxv���s3*Q�c�K�2-��=P���7�ヽip�+{�H�٠����-(�k�����l}�Y��%8�v�g�d��B5x���*3c�F���uƿ^&\��$�:r��+�� k.����[���kk��
��>~��J�@)CK����/m�W�/]0�cW[�u��E��-���DP(|� 3*;���u�ǇJ 8?�]��tP0�z#��;��J�3�z��v�<�wC K(HK�[��Ze=y5 0H@D�D[n���u��QM�cz�:��kDEh��bwg������w5���L4�w"P�ojq]��=C+��Њ��ѱX���籇 a
��`��7y�����ݷ�ѧ>�V�
P�.���G��^絵-7(������ֿ�OY ��-½M��~��N�̫�k�c��1G�� 8��L+.�C��N�#b���c�
��,°�s���^꽖�e@G�V<� d�6���/�ϟ-K�-b���4�22^�W:������i�c��=o�5��kb� b� Vyc�X�}y� �ؚ�m�\�{�}��<�r����i*�_}�_�LX+K�>?m %�Ư�J�$%~�N'!�o�] ��o��F���N/��˭ݓ`i���*��i~��~f@fo8�\��z�=�ZH���E��"@`�
��l�i^��J"��?X���֒���r<�7�;��c!z�VNǴ���4��ZP��96��9 ����
�%�2�-����8���h�8������o���"�m����~-����#������Co��AQ��߻����31�F�;��2�l%eI��Y򊀶v;=��ܭ�����B?[?S��8~���}��=C&��bs�b�:aV���fNJ��@�]P�0`����ȅ0��P�w�Xi�]�����J��bH�9���k��'?�	[r?��S�p�W?�� �A� ���?�ßp��8�f%/��>�ӫ�A��O��"�d\�Ѥ�����=rs 	q����r]��u�c0f��W�l�\�,�`�` `���>�</�e2���z���y�6���)��w>��V�J���
�d�S�{p����,;r�8Y�R�����k]���hJ�?ڡ���tm�r8ȵ�����$ �\�|��x{W30n�m9�[У�;��Ea�{�EH���Yi�s!(��}"����(!���6W}�0����{f/U�%�WF=�6�km�4�;[ \�w������ۧn�[�����J����!�&�	�����M�І-�?z��ۈʡE^j��r�C�xd���y ����xQX���	^4,�[al2�8���Q�%H�MuE�M �DA%�N�I�����(���:�k��iX�K�E�\�:,#p� �	��hh����A�OO*ƈ�F�!+h��ٯA�5�x����à�3��p�az`��=ן�|�R��Լ�w�k��H���5<j�:b+�ᑥ�#⠜�r����b[��u����4�=:��h������Z�RRR�.�����g7熍�1�z#�b�E���x/���XҮ���}m^�_t~����m�k려t��+�C���`I�ŪU���.u)$r�(2�%r=r<�#�!�����9z9�?�R/Mm�[Xj����{��c�c�ϛ_8�.�U�?yL���o���R/_��)d��d���^) ,���%&ԣ�7-,�3M���'0�k,��Hr�����ڡ�O�:�����a��w	������o�z���7�_w��h}�3\t���7~�����TSn���r����c���OB��>�\_�n [z�|�~��?����>�,�0�^�`D`iȞUP&x��`��!�N��m7Av�	XA�ɝ�.t��$!j��;��@4��6�� SKQxт�Y��D���}z����b��mmT4z|��G�zGKb�U����p�&���=}�O/������9�^�[ �F�V�5���j�P��W�Lqo9�3,���������%W�*�KRVU~-�*�ofN5� ��7���<(N+�/IgBs�6�P��4DP�#Þ�%!��x�]o�Y�E������t=8����ȭ+}��T��{��� ػ�� �'�٣�۩;3��ۇP�9.�x�����4��6�����ш��&��� ��[��������PTJU�bK��z�	�N9�'g ��Wx����:��2�}z��|��ϕ$5��Fa�:xy(Ս:�'����_*�C,k���6?��uY�}��߸G����FD�|���e���KZ�I,�j}��[���*,�`��R��Ӣ�C�횮�1��|����K~?| �u@�6��%�;�`~���[���f%������+����X��]���7���d�.Pr�bQ<G�&��Y��V�Ǐ�� 27o�����T�*.�� �o b,���{�r- 4��������k7����;�G��w�v�#����W���9��5 �>����r8;�vȖ��(�M���i���� h�O���F^8+����m��h�v�$���A z�b�}ӎ[8�������((&T�F{L( L^9��o����񈅹��:�.��ה�k��=֩p�?�:�gz�G�����;��uE����/�W����5�����9�
�IV��a�#��!��i���\���UK��K�rr�!Y��@���b�`s'ݚ��g�W����TRո���/���JǢ��a8P���)�4,������1 �J\g��]WW`w��Xě�@m ����#��������Mwk�tf�%���W�
lzk _�GO����:BnM�clcv�D6W�����;$��U��U&o�!������Rͷ�.���h�s�N�mT�3����<:�:�b+/,� �� �Y>�\�ï�˽_@2��2>> �=�a��\�W-��ů\>�I0�` X���܇�pP|���lQF�b�=��ye �'����NVb��b�<_Kȷ	G^v���p��}(��Ggc�`Q�����,�<�8�A�,�v�$�:i:HG���Y�$�q.�Y[wϾ�� ���P&��5Ӌ^$����,3�Az�i�%�� 0f�^k͸�y�GzFEfU�����Tu��៯��(���Ф`��,0=ު9��9�����1��]�r :X�E�.�ϒ�#����OVC�=���n�n�d�@�|�B/a��BX��@�k��A0��hL����X+Z��y�֛�/C�PQ��1�7�Y��M(��O���ʋ�Zp줎�x��7
}�Y�9�J�q�>�Lř���'��+����s�0K�3s��a����81>я�(9K�����[n��X���9�k�/b��r]E�p#�_ϩ���`I�/�[������6���W�@��{(T���鋯�:aЃ!(t++k	x����kx�GG3z���ִ)+V���ǚ*uy{#�>{����+V�0��]`�{��k�={���z� ,-oJ9 �=*zV�z�C�o�=��QxY��7���5���ƕ
/gx%���4UxƲ�#J��2�љ`�ha��Z�o�� ����6 C��29��A]�/R�^�b��}:��y��`-w��9��j��. - Zp
,Ȓ�������b �6���Lx� � ���1�I�+�`y�#>X,�؏�q>H��5Z��@^�n�$�Oу;Bm�昪
�Â x1]�ص	�� /$�L��Mu
������|���8�$NZÛ��"�'J��'��Gg<b��(�@��t6a���O2eI���.�gx�0ˊ�PQ�B��EF��N׹(ϏΦo��ʆ$�,���0��.���(أ��w~NsB>��P�P���e�`�8��p�%�B7�띆�K��OE>*\��Y[D�H�`��va>�]��tK*;���ɷ�_�˗7){����JQd�&�0��J �=��{�XS��#��4�&�p��'�N��]���:��K;��=�2����.�8�?�q�3?c_T^)����
��P�"�d�2�_���5�"�.��X�����X͟V�1�ޛ�m�u�:�T�b!�<=��Ȇq �q��R�sm��nR
r��	���rL���Y��8ǭ�+�-�r� X�-X��!��Y&q�����: ��M�u_��W _]�E�/ ���c�`@���?&��᪌��5�2@��v�ݬ��E����t�n�s�F[��R ޵QFR����_�KS/��	��5?�{����E�>q&C��[a:������+��^&�Q�-6$Z��մ!��`]XDa� u��-�A�;_���90�_r-[��IK���F�>y�0�����͝�?	pՃ\�0ۑ+I�0S�ؒc"�G����s�<oa/���+̀��J�"��9��)�A�V-qEju��.�m�u�MV�O��\�����5]n�Y�:4S��x/�;�О�O��x[N@�W��s'�������V_	����A�X�K�<��&u��<����͇<�,����l�8�'�����vI����) ���+�P|�GSʁ�O֬��&<go�y���]�]b�%�2+TȀ�*Ʊ�M]�=���Da%!j�&m=��ꚮ����6��8����J�^�{
�W��<-��z@������9G�7��2����Z_~�%�C�Qp�g[E� x��Ojd!���ӧ<0�ď}��l��K�E09Hk�e�hf�j#5 �`S��"�xa������l���X �HTrs�A�>���'��B�N�m���"Xk|�>��@"�7x�'�)d���4 �P�Qނ�k�ok:��AЏ"�U�ks����>�7�$��_3N(��(�f����^A>��h��pY_"&��� ��+������ >�A��am�L	?�����b/1p����m��XBWjQ�ev|͜7x{�ŌF#K�#�Q@��2dq����Q��P^���sv�"��Dm+C\�S� K��գ�Z jX�l3I��`錺r��6w��}�9N�n����H�C�E�$�ʲP�^%c��E����x�Ⴖ��Y6Χu������ �D�-K�?/���L�[��M���Y�!� �q]a��2�=��I�|�A�a!}k}�e����AFY�})�f��� ��i5 ޟ��V7G�+sT��R&w�A��=�����a���ʠĵ�ˠ9'r��׵�M�>F�ժ!����E�I�W�������'}o�?NCm� ��cG[P�3	V��9��ζ�Ѳ�1�{��������\�Upp��O§�.�6�(��P aQ���d����u@�5 ^EJ�2g����ʌ�p���tJ
��0fB(��.,�|�0!�o���_�EL�!���vΉF��N���V� ǳ9gx�}�AA7nm��;�hks���9��X,`��'��Q+2Is\1>�Y���tA�w�igw����;6�g�⮻׋��ծN���w!ê�kPX� ��_���w�����^?�Mc�69��-&4�hk%�t����KW!�j,�*v0�@`!�]��_d���b�`�1|f{���ͬ͞��Tt�XF'��X�ڻ�oLf�����R\�+�Xx�"���Xy�v2��oYB ��`ا���t�	� �-�쫬�NtGR��`���X�3�M5w�l:s�񐎎i:AB��R'�q�l��[!9R!��z��#^$�F�ӂQj5�}�#H����P:N��o��H
����,���S�h���ٵ%2�O�M�G"�<#cf_#F��{��Q�F��p�\���c���Oj�Y��V\s��ڠ����c��K��X�<��ay=-�K������|����C�~����ߘWX�u�|/UԵjE}��޿���A��R�6!�?��bi&�6����x�a[U=�e�B� ���H�2�R�}����u��jiR#8��f��@iQ��y�=Lr���s���X�@H�ji��Th4�vmn�e5m�U�L�W�1�hH��"�M)�. N�~9C�np{�����+��/~A}��AK}d��� ��u5���Ju����H�$��N?^�$ya����$�joo�ӥI&OZl=ǰk�2�b@`ʹ�EN[��-���Kp��޼A}�.=xp�F��"N!��+ϩ� \߷bC#���8���E1p x��������}��M8i?�0�f��h���|n��*��q������m�ogE;Dxi�N��#&lHw�ܢw߹E�w�n�@����^Q���Lr�|T�~d\-�>�F7�����=}���������K�Cu����p���X��8�_��-�
�� � ~���hh��Û�g<r��=����w�Э��`��eR�"c�2W xAXf?x#�RxBSPĻ@-ꝝ=�}Լ~��G����9{;�2Vp7�rj����ۑ3�箙�,�,�]V������J�a��3ׂ��Q4D���|���֋&�'61HCm6 ^[[Re��%���Ed����m�2�/�nr 8��X�b	����F\+��d7�+�K�M3�����b�:��Z,l���{r���Ғ����ZG�i�aV�o�=>t�T�G�T��kb�	#�@k�%���&1�<����:ߴ�'�4u&��P@���^vϥv��y6�^a�y���i���5r�I\ŵ,���Ɨ��x�)��:|�
a�k�W?O:648�g��%�����a�Cd�x`�FТ�/��s�9��q�d��� KH�V����t\�z�k |I(���I�ķ�R7!Bo珃U���Vܣ��V����*'�,tΧ�qP�w �&������.��r���_5���B��'�1k]K�~��]�	��-z��'�A9���1Mf�X�	����� ��NM
��Ex[u��y]w�N%�I��4�ԩHī l�4� X��9 r�~����g?}�����DH$�/�!Sj8'$n	�y2�W�qe���4���>����g�����٫��QZ��Mc�Nn#��w`^f�$	���d�z��(T�m������?�=zا�hC�w�m���|e�L_&ͻ�s`�؟��~"��'�)���f��y��^	�ɜ������}N_>yN�|ח�� �P��r}����.XD�=s	�ͳ&-8
?�X��m��ߛ�7YkP���K.\�9�b kQ_(�PsX*b�-mA�uƬ|ۭAomI��)�~�UV%�����Ϡ����Ͳ��
 7�\A[D1ַ�(��2om�$��l��F��[��mj%�jY�6̑*�n��c29rs��!1>����alf��D[[�9(*�B�5�
J0o�&���{���#�T٭�g�`\%�2L�+��(���E���/�>���;���oR de�phQ�\��=�VqO�\2�ęΧl�Æ�郵[�vPh��.�t�~*�]��B%9,��P�J�(q3��<�mY�S�y��Md_��r�y���MQA�B1*�چ9����{»C��_��_�/�Kv�FX����߱�����\	���������q��$Xܣ���Jgy���v��]5�  N_����$���t���ex���V�����b�]>Wb�{}��a��y�k�o��b�Q�8��cvݿ�I�=�M�n4�;��˴��Ր��_Z����x�Ly��}��mn8fV���Ը��������S�?
m�>JK���)��$�Vw��-˃,$lm������޻�蝇�4�s�q��P���+[Mz,42 ��ht�f�nn���4��S�&Z~Z�6t%��npM�B��`N	�<�g�%Nx��A1�7
�����7K���ss�G��P��Cp�\O*,�W�U�Jp����-�U=�q��	�n9�m�捑�|Eov�qp��0�*̂|�2ڏkw�W�Rj��vYLr�o�X���*8Y�5���s� �L�����v=_- ?|�+~)�ԢD�����G�y �!~�p-���|rpُ�.�ajU�����y��k��Ͼ��^l�0	8h��J��0!���7�����h�7A�Y_�" _�U�o���>�?����N�zM�A���"|�ƇlMC��Fz��/$m4�$��m}�3�z���JF��m���sk%��*&R�`�[�	 ��+��:�Y,wF�	�� .� ���O�_���2�: 2g��:�,Hǧ�C]�A�72�p������������v�w�7���˿��@¸����	�>���{�����뉢C���E,�8n�o�t�QH�Қ���MM�R�]C��9��t� �KD�6A�M;4�����>��O�_A��a�K�}���� /��h�����7�N8�����X�����P�4����A�N���-�y \�	��ݠT�WM����C�Fˮؘh��G^���"��m� aO&��8����Յ��A�Q]ڏ�CȌ���O'X���ń����H�>��֖���j� xz0��d�-�!��$m��m(Q�����_=�X<�	2��������xY.��3f��VB�]��N'pO�;!g���d<����]��޽����"�B1���W�lmܦw��ߏ�ޯ>����^��a���µ�W �	ev*��ѝ^���$TE�� � W�����h����}(�W��
� �D�)=�{��L�/�ߌp����Ju�)X��Eˑ��[�=3���c\)5��s�S�RvI� ��z���AQ�9���Ic���OT&e���DW����C��J����k�$@F@H,{ � (;;;���o�_]�S,����t�c��"�4i+%� @$.� X� ��Ac}Y�<��e%�t������w��������O?���ƖX�e��e�>���L�LW���R�oCEh=��6�۷�$�-X������! ���wc�n0j-�,��l�*<��)8��⯎�G�K7�$5
�X�\���9 E�C��zl��mSgG�Q��>6�	��8��6:��@��G�ULj����~�V.j������z<o�yMM��R�$ X~��:�s���e|ĿI�U��V��9�x��0s�s��w`�Ti�k q��8�n.|b��
~��C�g�� S�s��"_3�0���m� �bK���V9XJGՔ������,��;d0�90E|��ϧ^�Ʈ����/�.�9ڢ;wnР }������Y�5<וi�[��gO:�P��i�n�uS�Ϲ���6��i���k��Й"���|˳�P�*��3|,[�H��Rk�P�+�;��{>�ൊݟ��vP�O@t�Df�T{-�LX�: 8�'K�^C,�;q�ٚ�7���S Xmb9�M�!����tB���Bw��łQ^	���r��=9�����
j���$c����w<�lcKbgźM�5+�A��Qvl_���Z_3�m�%M��̏Ģ*m���C{��za�� k��zŢ+.� ����`�qV�y���$ý ��6��`���S�{Y(ǋ�/�;�y��zޤ��������xoR����?��ݞ����3b|?��3��}��ATp����˼���P�΅�mj<�}rpJ�V�q��dt�
u�*�b᪊��]����>������O~�&�m�M��y�ecY(��q����9d��h6���<�_����TH�u�<��*h�q�.�l�9�r�TN�, �H�z�,�l��e�����d+����J�%��Ě������R~��O�â���<D�R���,[�{n��[x�� n��� <R���� ����f!��k���6�ӱ�\m�(���5[��5n����N(�; ZR�L�p(FG�"�ߦ�9�~u����S�ލ��рn߾��������0C%��l�w�S��*:b���}���p�������^�6�������"R?U�bJfL�6^���I�����g?�>��667���Q1��X����m��:	Vm���Rh�'k� `|���0핰��ۣ��`�]����K�#��P���K�����{,��j���5S��60���=z��9��?��+N�'c�/�|�]3�J����W1����'-���2B��p���{���P����a����A-�G L��,m:ɼ� sO��-�`���[\X���
��oxy��J5�{��OqM֮�97�6(��A������-�1P�ݻw�>|ȵe��6�?:�5�/�f|�F�L[�;iŲ_�) ���<rH"i)W������c9W�y��rm}����_q ,���������b��[�kh�AkS׀n"A�ˏ �~*�6Sz��}������??�;�o����cc*J�K~p�
�	 ��Y!���XL�-�`��w�p�єb��uZ��c�`A)M�^��( X=?f
+�>�I����o�z�i���j�d����̷�����zQ��
�l�Ӧ��l�Ɣ�?1�O�����x�l��o�J��y��?|��g�^yL�B(�w!%����q��d��k����Lw�����௼v��RxO�5/�Gsg��m�<, ����*X�\�p� �[�&3Ko�L��o��.\�*v�o@��G�f�p~���ݠa���%{�XV�qK8�ќ˻�4��w���������Lð�ʠ�UCg�zr
�Uʻ��۳���Y��-��b��xp�J�}����r]��l�  W�6)��X�,!&��N~U�'i��S[ؼ���2�Q�b��Y$���!��ݪ]��_�všyNYu������M�d�]	>zH�ѐ�~�5�|���7�,be�tKb�ɵ!v��C7I�k��_g*�˂^���㴊WԀ�&�z��qŊ��K�����ۼ(t9�u��EP�]_�ETE��rc�:x
"y�� �ڥYܒ�) XS[_vy� ��b��	~��4�)��h�ݻw�;-x��'��2۞[:y�� ���eM�"���9�7��X{�����Sxo?8�����_ΓB��~�+���b&���P�AŨƨ�d��Z����_^x��'c^m�U:�;�H����,h����w�u�Ϊ:>r���;a��5{!�b�[�b�0 6V���6Ǔ#��D]^�1*��ӅE�����'ӲXDB�^N�U��*��Y��(�B��j���m^y�\�Kt��� ��6H���S�e�D�1-{ûf��D�M.��-��P�����{�"���G�����Ms,����>�x-hQmɯ�A�4��Q�R��T,3^C?_8f���f���v7�i��s�
�v��x��������m�v+��N��h�̊H,�7?�1�h~���#�	�p�0�UT�X���dL���>=}�KO������� �>_�����>m�i��}��������^Y7��(X9�x�.+�s{�����ή�޸��.4�ՂպB�y
��RQ�(�Gؑ�ڎ��C8�������=������ڳ��Wl+ ��.WI�-��w����q�����Z>h^�4j�柹�V���~���-n;Oa� 旎���x��Bd�F.(�����}��oҍ��	z��44>;�����@3�rh!�)��˘J?D�T�����<P]Z%"�������`�R�8��/6���y�oT�K9%���� H>{�����kNJ��9���*\W1�u�b��W�����Fm��9b	�{��	n���@`m|�w8�0�����)p�~x�����9%���Z�3����q@��u�#�3b�a��� �OX�E���X,�P|��(?ڔ�Y�R�� 8�����5O[>i?-���E��(7��Y6$�
i����
�!`|���n��!�ڭ!� XY_GVbku��9S�	4��"θD�#X�X(	� �+hhM��>�4�cq(���O�OuO�œ]�ǫ�Ҋ��֝�Z�f��W����b�͞�>Њ���(���,�t�q��|��F	��7����G|Lb��>�KNEwU\��V-H�_?�t���P���;+��B�I��/���gO�n�z<ί�;��IC� ���ZޕO����K���"x���Ƈ3���g{�����9>V��#�G,��{t����������ܿ����,S�#\��7�t�F������<^�H!��i)g^E��v�u�ۦp��Zn �@������mh� Zm�0��e>E�E:՛^�M�|�ڹ�_N	b΢��DS�ṫ���,� lq�E�[�dB\v9���~m��/��._��}�{p�<P��]�wb�U�����k�`����?��_j�캬W��>c� X��
�9����uE	��I� ^�]�`�c�.nш�����RZ����$��X��O�7��@���$��6k�_j��HJ�.R��
>���dg��z���e9������������&�u(H%�J
���>����Ĵ|M�26){t� pp�4���eAkdt�� �T��:/k�OC��+H��+İ?`���q[\ϯ�8�����}w.j����Ν������g9���8��I�T��1u���
p#�5�Z	8�e"�
a>�jA<M�B��	�I�Ô��b�KJ�������0�l�C�p�e<H�W]�8>k��l����F�Yq������EQ�[(;bDȅ�����������C�o�L�:�'��Dl������=��M���1�0NnXU�U��f7���΀�6or��t@��#>e:��]%�1�q n�VY��f#��Xh ���zl?��DQ��Z�����D�<�i,	�=N�|�mɒ�ckBV�BbMg,(��Ht���V�H6(�J���j�S�Kj���ME�����T]�=���m$�Y��8u��U��',?&n�����:I}Uo�DD�� ����_�kEb:���石��} I�0y�8d�"cTS�Vf�r���é�{�u �x~�ӟ�E<��:� �
:oe�0��B���݉5_bmu�Ĳ�z
�� �%�ЧO��-��1����MLn��K=�������_��_�2.�w�}�����/��r)X�{R������!�`�JZ�c�.9nk���E2� gȴ|�܂�h�,�
�ʂ�ax��;j1�ˁwo���<���(�99���D\��6�ˮ��E��mt��˺�é��#,2'�S�%�38b��;�7���&"-*����<x�
��	i���WiB��E[���P#�/!�-�=(����c6s��ڱ�ټ��	���S�WN1}�������kt�����#�ۆ�fh,e��2<[��R����`&
;3$� ?--�;׾kt�*��k� ���&�W���s*2ɵl{�*A��%q�d��n��5�l�k �qu�`J�J-��9ks�7Y��=�#ײ&�ݨq��Q�*�M����ù�6ݸ�U�X$s?7��7�(����'O�����$��c{C|�(�NC��`�C�W` £A�ςgPB<����񱋦.tޔ���%<��ko�{S���Y8�����O���g�(��}��|��3�� t16�� �q]�����1^�6��~Ex�q�����v�CFI)���jƩU�6��[XNK�M�R�[����u�f�o%�J_[nH�р�+o� >c�v�@{Ƅ,����y%A�DB ���`F,p�*y�x�ZXЖ�N�n����������Es9n벒~��S>6*g�M۰�գ A��=_�qv��n(2�1��1�ץl�Ow)0���W�L3���E�"��g������~�F2�����;q�@��z:�eᖠ
)���� Q�e�8w�,j��ВO�k�"!� �\\3C	�����^�7/�����6/�iZe�ls���i=G�\��ծ��`|Z ����ymm��h|��{(�«�&?�%;���k�C�� h��"�#
�ӑ����C������ԇ�m�}8���Ut���ٸf��2�m ������ ��ӧ\���+�u776}X�b�|���ۣ�`E4�h�����a��3��W��,�?��O����g��dK�|	o��}�����seP�|<m�ʱ9J]���K�?��?�%V^X}�eY�{y��@=��x�0)�<����x���2Kևf��������/��%w�-c��Ԣ��s����0�@K ��!(͉��(����� ��f�mm: ���! 02�Vֳ���s<�hx�66�P�w˵b�a��_=�0:�X+�ʁ���>Q���ª~��B�Ő��b��\t-u�Ϩ�s׫�%'��<�o9�[�Zˮ��Yа����6wZ{�'���A�d�qz�T�,��:����R'�B�4,t���a�ʞ�.���l���p�n��a���G}2����|">#eSD9C2��G\Nو��ŕ��(ghK�rZ��J:�e�i�i�yV���1���>�|9��$�A�ey�.���'�>�����f��Ӓ+�4�i[��T7��k��Kr��0�r��.���8���1����eBi� ���E�m�'� l������4��#�T��K��8�1�f�=��
�������p�ƻ�K��K�EZ.K�)���Pl���Y�)W 3),bŲ!��5tI�|�8�{}�ڥ���/?�q�I/��(�.{��OHL��d���g߲�
�9$�`MU`<�ux�f�>��sz����p��?#�3kgl]����[�����;�4�(B'����1�`-B��B�v�K�^Akt��K�p�X�"闋bD�rE����&�4�5��eZK������(���h�mbٓ�^�/������v�[D����c�&�M�mX��܇K�Cx�+�*[p���E��!����VIwn�o��ˑ;�y��xX�+�ܲ>���0.��ft8��0a��Rl�w.��s�)���2�q���m����
����[�����%�[��kH��.E�C�t�,2�s�w��rɞ��J�T,�EHX'���1>������G��2$I*#��mƳ�����{&ԡ��gdy����/� �����.�\P2�
!.�� ���C�cY����aՆA	���`<����F���mҙ{�d(}Fvq/{��U���R�A��~Ÿ��3��O@�s��)I�$St[O�.% ^~� TY�-u"��Em�0ۦ`ߔ���rC���� ֔�g*�Ѡ��YM5�)IJwLNhA��N�1d��އG���J�%kz/L�"Q�>gW]pAx�<xl�I��s�y�����QQ���w�d�i�	��:h��(I���m̙e�o���y�O86��ii�w]���S7�mj�廵2!m�ɚ���ڈn�@��N�kq�h;jcj+��MxwV�������\hƊ^uj�������=G���ٽ��O�Fb�	6_�������ά	!�"�z���Ɛ>�I����9��8o�c�43�@�w{D�o��;#���
5�ty�$�����͘>�O���%��,�EzE��\���%�ő��ڑ���vm}�tzL�9W��r�v�j��Y:�ֵ�ȻH߉�������o`  ��IDATD/���,���⢟k	��K����oq�)B��by<e�i(�,s2�؏��� C�c��@A�ܗ�4���/Z#�{�۳X~S	OC�^� ��;E��>
'�K�Ѡ�5��O�5I�j��t�_�9ɖZ�&��!H�Ǩ�Zs~�9�Y>S���)I|�1( �g�_v�址m�۔�v��2|/ ΁ߦ�M�9���YDg'x����ў��#�>5Z�W��.H��h9	C���I��C���X8��`�Ec6�6���G��c$}A]Lb�+� ��ݾ�>����:�8kj�gB�Q��_Ȉ������y��=t��i��{a9u�_!^��~�BL!�0�8�����YW�*���Uي�y��r�5�D��m�����@8��3B�B������~���0�� /6�J��A��������2T[�k˯�%ձ������D�ҩ�����,�*�g���~��q@�r�P�OXYg`�){4���[����?�φn��wo�~�Ǐ6���';��hv-��n����o��wn��}l�_����1z���m�wm�=p{���6���.�'�J��`I.�k:>���QL_��߰��묝)�kf+^�ޛ
s���%����c���Iu��g�7�R^h�=+�%�4��*ebt{�����c��^��V�>�6c��������3gci��R '�~��"/�)FV�+=N���S�Sjx�Y[+NH9%�����)2#��׿f�9��8F,k�1o�eT�~m�K�r�j^���^R�X2Y㹥��d?��	��4���#���I/ޓ�"��uP�5#7�5[x��)Y�U�=��;��h��oU�cip�`ٲ�N.���P�i�8ֺ��j����(h�dR¤�I)Z)�F� ~��(?{��,+��ݣ��_R�����=z�>���cm@�E���?W�` T-���p��u6���iwo��UYu=`���������<(��0�_k`'�!�h��B�&�X�t��r%n�9k�j�C�(�b��}fN�\=�@srIS�B��E%wP��dk�fx�jHz�����`�uͫJKj�KH&���g-i������L����,��+J�8YT�-|	� 8c.���hT�� FCǇ
����`�5ʇ�>ݺ���;����m�`��Xz�F�8AV��X �����w�ͦ=��;p<��'�m��Ka|��?��4��)'���c�V�%�[��q�����VФ��U�Q���z��;�kNpO�\74֙�k��3��\�T��h�u?�
ZM:lH�NDK�j���E"��-���ci��#E�Ӿ��9��~Q�J[�����V_��"�C� tq[���
p\�1⸤8)��3�yAp�7p��DY��\�>*�]��:t"��Z��ȍ���s[ێ���$��K���[J �E���;[��ڼ5�\�Pt�l]�2
�����p�,�ep��~+���z����f}ԓ��I��	鿱�; /&)�ǡ04
س�j�}��M���8@��{��'?��� Ȭ:�8�b��n�x|Ě.���Ǝ	loӋ�;��g�}��O*�
z���f�˖Tq�K���2��B�k�s9k�U�V�s@��u��I��i`��,&�D54mLD='�^�S0rZPu�ޑQ!�s(���O�����y~%�� a�{�"(�a�5}�R�7��}���&P*��r����7̎��*�j�X���!ݽ3s�j�\v8����dρ_h�g~��r&g�B�W���lЍ��4[�ioB�^�g�?s�������JǇ�	����VYhץ@�)<sVf�).��V�a���Lj`�Ҙ�%��r�2t�%-�z_�eA�}��)0�T+ݵV���W������
B6Z<�V	����#����|�Qc�x�XpqO�y�'�����LH]�B���ӵ�q>d���Έt,;�#�XaxB,��~��,k��
���>�2mǠ���%)����j���3�û�s���s~�����zg�� �f���-|��.=��/�+y�j+C<�� ��X\�������:��֌��0�4�S\4$�8�-�1I1�0�����4&&�*�����	u���=\8`�����焻�yi������9�g?Ҿc~��6��8&���}�ZZ;���k��s��3`a�����dhE�n��nA0�z�|8���7�>a�ﶙC�M�c[��;3N^���A�9$��F_ J~[E��M��w�2�j#Q��fW�
{yo!�ҿ�"⟦U��F��g��e�k#�&�A息�D�8�Sl:�2u��GE)֞�+f F����ŵ-ݺ	@��0�8�<�p�0ő;�->�5�
��4Cw����ٝ��xN�~���|��]g�-�XѶ��I'���{>/:+˨P�����ڍWi����N~���f��I�焰U ":N�sΓ.�����%M��d����5�6��7f}�������
��s΂���C�D	X;Q�퀵n�RZ
�&>�$��H�/K��uH��yr.H�C���.ޗxn�_$�}�t� 8g|J����w�i��*Z����3�oi���$m ,�|��~�ҍ-7�o���V������mC6�\"	To��aE/_�ӛ�3����%�	X��,��>�����~�����$n
�t2�I����|`�{���|M���a�q�����b��"� ��=���?������񌦓ͦ��/8q1�AW�����4�r;_X�����u=$������$�Z�+N���S��6��/3#�'�U��m&'C�u:���_�X'�u��Xz�Ow�E�BI�x[�7 c%^�-�xoo���kW�=�4�]}��S�ƨ���]u������mA)	%��9^\�>>!P� ��XfÍ�+�x�ⷊ�%�m�mC,� /� +}v}><�@�K�~����W�C_~�������M��S�9�܄��ב���.`�&��+"D�M:n��^���Z�q2�Sg�a�wC���� �e>��{�� �/�ð
(��c@ �$ɵ/øYEx~���J������#�5�A9 �W��$]�\�����>9] �X��Yo�- 9aikT����t��ݺ�#x4 �
B|? .G\c0(��vH/_Ru ?�9�ӠPò�&��|z��Ĥ ��pE�	f�	�4�ֳo�9�A�yw����hwo�K$���h�C�ˢ𭞹}��{���K���_|�1x�@{��
�E��

\�yY���u]'}���%���4,�ņۆl��e�X`�!�K�sQT��o�/�Q4,�6�Ge���{�W��r��խn֙���b�?n�#Y��K��X�X���:�@�h|��oN4ǖ�fr��}���8�n���.�|u��ސ��������� �!�JK[������3�^�E
X~1gʞakpQX�6�������,i>CfIx�ҫ��۾�������|儺W�ܢ��|'����4]��(����#@�P�����Kr�UWma�.�9���C�V3}���$�Y$��ێ��-�����Q���\�b�$�Ok^6����(�|F��{͍CZ�?��.�Uo�7^ȗϞ=��Pv�_ ]i�</�
K��B�$I��^vwh��!	�p+	��� ��<ߋ/X	���q��!��M�{},�M������:i>~�}q���K��"�>#��?�tkk@�߹M�l���R�7g�"X���
�ኻ9u y8��c%��M,M�8�@�N��iN9'0�1�y�������a�ű �qqf��ͻ~�[�X�zp��43D� ���՗()�u676�`��2��6�Nh�B�U ��z��o��P���r�n�����S��ay�~q)z�T�ռ�������׷ܻ�h��!=u.@|�L)2{q��k?h#.xK'�E8E�ݧ�xK|�]*1��{���k��»��;���̻�I`,�T��S�s �yӝw�zU��[�=�]����U'+B��>�2�Ø0��v���!�ۯ���y��k���@���Cbj~"�_�?��:�̙o�Z�E�^ o&�����
{-X�ЩM&��=␎o��������/vhg�5�}(kz\�gd�G��]^��v���uy��.���)`M�* ,1�m�9��=��׀ʄuu��� �p����m���"}O�%u���c]�Ǧ��5���N��q�O�xe�� "O]��֒h�L$ ��>��s����!�� �!�Ub�!g�"�O �Om)�0��)c+U]&��[��x���g)�4g��w�c����_l��o/�~J!�-ߵ��n�{[{s��$��ŗ�}ma��Х�Y7�z''����sR����߽9�A9�,	\i6�칿L�O~>��8��|��
+Z��)�'a���������T����--��MP�b��B9l����c��y@�i����I��z+l5�Ǔ�^����%��`����\r�XZ' ��`*朥Y^Mii�Qҳ���1�Ù�X�Z𨭧��\ن��]k�N���q���QT�D���@�t2	8^g������MA+��"!ZE�Sz����<}�~1;t�&~^yw��o�z�0�
�DR�^߸q`�ʶ�s�J��<�Ԕk:w��l�Ӵ.8��N7-3�xR�K@/B���Sz�?�O>��>��sv{����{oh��* `�(�42�Lf����D+|�_o	^�z�+1 WHҲ���z�j�^�|㶗�����]ks���p��a�ge��'>_z`�,)t����V	�]V��� ���vY*4hN�����y+�$J���� �w�W��J��o
����:�暷��}-l�W�d�M=��8OK㎯]��W�b�/��6���ij��T��fO���_Ȕ � u�=%�Sx�d����k�D �Ӗ.g�;O���T�<@��=��� <3 0\�%ɬ(��L���o`-�R������o;ɳ�y�Ǽ-J�O�\��6�k����Ϧ㪋g��֘{-�}ip����m�pT8���<�U�P9�i���ݠ���g���*�mH�S�|�dPcB-I~al@�����ҍߎG`8������~�� L`d��lt��_|�}��	k�^M^Ep�ς�ʝ᭿pu-C�M�^�Ё����A~ptH�;~P�lѠ"��2����lF��fB��������10E�͌����2�BY��A�F���3�/���v�h�n҃�k��a>�{휲��U��s�I�׫s}~D���}o�4\B	V�z�w���EA�_�v��ͩ8�=��}��m��xB/_!&�K�����~��K�c����m�(d�4u���pFO�y���x�L�]:m�Ҏ��'�Z�j��8��b�
��[)�+.���%������4��	ѷ/��'/�=q��s�M~���]����T�lH� ^.~q��{e�����8v �Y�o9��i�bޙ��<������딛�����֦4�O��w�5M�]B���ݖ�T𲢥l����KW�� �	�cNp���k����-C���������~�B�"*�E�Ϥ�9T������3�pc:-5������� ��eA����,URH�ݳ&���a�D���~��l�a�d ߻����e�`�b�1@Q���������y�_�k�/څ���pe��1��!K���[�#�y������9�õ����_��G=�.���I}=>��]���x[nۮ�����M�Z X�����oE%@-,���Sw(��r�v�R.� L�c���p	���ш��Ʃ��	B�I�T�b��
m�2�����p0҂�>�Q��M���-fJ��J����Kr�M�M�q�6ݹ{�ݡ��)�&�g( ����3�]p2��f��%���w`��R�����_� �" ��c:s�d�r��L��7���ER���c����~:
�M��y�+�^�u��ڤLf� ՉvM]��hB;;{<����oؒfx�^�e�u����jA\Cz׍������Q�����u;~=�E*$G�S8_F�	�Xͻ|��>g~��R2[�t4u��!ὃC���d� [��/�㇃��̈Ǘ�& {,x�*�<�c߈ цǄ�W�9���P�H��χ]�@��yҒ򄚠��{�p�ʪ�޿�{�γ��1r\j����je�;W�r}<��+]�r�H��8_jOR�YX����.4JNh�@>��q���[��?�zY�S��$���ڏ��(����Ȕ 1`%�  �TɁ|ȑ>�*9�l���ٍX�µ����$yv�xN��E3~�/6��d8�w��8^�b���R���ϗ�w�1��y�E9�Vn�6�):�iw���:}�FmJ�u����T[	D"3�$[�<��!�����b 9P�$�(���$����tb�d��3�-b4����{ _LXLHLf�c�}��L�ѐ�y�ݻw����%[SD��a޽x6�u�n9����4w fk�&�n�:&�K;��7�0x�E�[b+��-�������{�9��Vv�	��OV:������aMi:����v)����*ꨭ��5�&�ޜpV��U�ՙѤ�`-4��e7��ȿ���x�z������`��z��nB+sD�1Qc���8����#���H�J�/�&c܊ �{�!#8'��q��x�vE�r̗�\֏y��W'p9�C��E��� �E�Ja!<n\�&؁9�@�4�b�õ��'�+����|jJ-[�[NH:I�T��IM]��5���Q
`�ʩ%0���ɜ�e��Zo�S'[J�CyhY<�EK?��QGp���͋�/^��~z�
.|�n�y�B�H٠�Zy�DX����1 ��_XBa����u��y�����k��ׄ��ѣG���w\_���v^@N�#lRU�L����n�⺭���tk �A� �u ��5@}� �<�O�C��wȳ�@$o�ry���|p���4�w�k�[ڷW
 'S�PxF���/�iNJ��/���8�f^O �g#8a �i�&�� �$(F�&⮛�HRF�	z�m���~� u����f�5-fc��"4}N�9 {px�O|ׁg�۷n������g�����0�v��Ig�������K��9�m�h����`����*���
Y\��m.��n6&(z;�j��oYZ��'_:Ъc���:�[a�Y�Xov������?GGS:O�ئ�a�>�ӿy ���ʻ���{bl�$M<?Vt��6�K����j����$&$�+�\d%�V�p:��J�NU�&�Ե����-6��d6=x��+�f Wv��ǉ�L�|9��	 ���Ut=צԲ���i}�.g1H-���CX\X���b���T�ͭc�Xs���.�w@�*�EH�K��浄���������d>WB]�<��Zo�N���C� ���(Ʋ�"
  (������EU��J�h��<]@.Chܖ�Z��gƦ���צ$BI}`�i��M�g�><�3���:Oj���+J�u="Re�EQ�J�FW
 {
���~[�q9����ؔP�������>��U����q�&��V:�H&.&!j�!==��نI-.���'��|�qÏ�{�zN��~���|��q ���i�o�z���"	�Ё�>x���]z��K[��s�^�z���4��v�h�
���+桜ʀ�� � ׬��uy�RqE�1%��(0�6��u)S�(�(E�f$
çd:��11fڂ���o�:].e�	��V��xEE�j��-����U��.�x�/,�Xo���T�7��K�x\�F�	őc�-��EPƇ�.^^��PՃ]_ne��_�g�O'4�,����pG�}�.�RLy��l�wm�)�0Ǖ�OUU���çg�Lp����ySwoå�B�E!_]�ː�!�
]әSS@���k:{���4۫����Z�Nٚ�識�Z��sw����:iPp�
�	dG��a�\VZ��X�$�
���L
a�KmR+`^Ar�$���m��7�8glxf��@��}A�'~GA6�,.�(�$J��\Og@�.RX$_5�R 8�x��p�r �"�q�#'e�!��x�gr �������@��1����N$ u1 @����"!��mç���J<r�h~����;��<z���q������+�{�M;��R8s'��������`���}@w���[�is0���fn�'�[�"�~��\�^�O�|2�I�Ϯ�w����%��s҂�*\���I, L ���F#:Y��H��h�Q���"��{u�U��'i�(��;�-ߥX��ɀ�ƻ4� g������>��D�OQ|����.�G �����bJv>ew�;�_x@k!D�},0־�$��+W�9a8�o�/�e��� ��:�|O qkk%�.���}�F%vjy����k��f]G�=���Z����v�v�V�u��Z:�\Hm��ے������|�s���ߛ�i�����o�5�� �~�� wv�Y���0s���9��)ȍ��	�@�|'q��G���E��k+-΢(��d���,��VZ�}�`�7�UNK����\����א2� �z�"��<Xڼ7΋�£�Rvi[��m�9�2 �ٖ��׃VN�d�U�Ґ-K�X� f<X� ��m�P؁Md�xf�<-�ә�`L@���ӟ��~����pY�(����W��<e�c�� M��}I�~��z����`�snv�	�'���D��wާ[nb���x�'=���1,���Tk��yc�hOr�		Ьς�aQ���q�����ڍ9#G&X��`lm5q�� s���c�����	�7MA^bO�#U��B��{��D�2@��4s���Y�
�1��/�g൶��ϡ�����l����m��Zx�U�1 L?�|�9$!�j����J<�$���x���ݻ/������w��ir�B�l�=���2�9~8��·����ܵ�!f��ܹ3��PqJ7P��M�&z�����vp�.u�m�z�j���S!V�mo�v}�.�~`�T}ϓ�d���K�b���Y��\V��䷋���w�y�����ơiI�t9F@�: C���)��ϰ��&e|�"�8ח�*�`\ {{Ǘ
Kp�k������ ���2p��8h#�(%w��'��K_�xN;xfIF+����<�hK�70���� ��xf�P��=��V}��H�x_ ,E�[� ����d<���7��ь67 �zl��q_�qz,��j�:;�1���E�X�M',�l"�8�Ѫ$I4Y��ЮIZvh���	ȵ�H�I,`4�AYѨo��:��ä�d��I�
/�����o�X\�:/�P?��=��@y�h&W�.�F@p}��t�A9X��B��L��7���������k ����|MBB����}����w������̍�J�4�q��� *˫F� ��_NG��{��>����W��s�.�E�l�_��쳺��޽K=�g��i�7@%�[y������L�O�~�9��,���&dm��|/>>��5Q5'�ANP]�lWǗ�Y�-u�&�Ϳk�������k�/�^�����{7�7q<B566�4����
.
�Qρ06E9UZ�[�m c<�"���	~3O���HζG��t8��Ԁ����֜״>u��hK���\�.9����6�ں���6	��~�� N�u܆��mr��9���������E�°u~�̙]O��WC�j�c�����;�k�[�Ԩ���ZR�gۘi���ƭT�ȑ��	C
 �v�=��� �ÃC�s9C4H�� T*�Ցm�|w��BR���_������t��ͥ2Si���S��tVh�� ���d�|�Z��y�uxH*�^ �J�6�L鱬�e���,�8��u@����M 5���	TP�� �d��=�R{���a� 0�';�oi�Lg0/���t�����
�Flk����F!�C �^$&�u����ʙ�%^�c?��C�	���A��ۿ�Ѡg���-�����}X��1�`���;��Bs���l�\�Q2����n�s.���Pv����T �`5�4�E#�I��4�%1�,�Vb�������vv���;w��{��chP@x���'lkw`Ǭ�67�q���m�F�*�)�<x ��CO p ��z\��WU�ٷ�q�"C7"hN W>��h�����I5 nvw�M�f�������
��܍I���c��:Aײ�;�W���R�lS�A�YW��J#�e��1����A��dLx��C?����<#�w�����j��e!N�Lc��0�<s�Q�%�X|�����=����2G��}��5rsnĮi�V��U���^��3�cXIT�Bl-�@����[g� �Λ}�۟:\��;���O�����z��eYX�%\��^�����tvd�+�0$�J�%�E]�㪿�~ρ�Ԓ�*X��9����u	w�6��Y<���1x�糽���m�K{�p���D	���NJ�מy٭X�[�ri�l���냏ԕ<��	����W��/�B ��3v��(%|p�I p����"��7���`�Y����)+��,��*��U����Z��-	� JA��}����5l����5@I�0H�L�0�����E�rⅥ����s��)7�u���P�ą\��i�PZo��q:�RET�{��� X��j Jn0`�9[^�>b ��h�����N�
1�>�(�����̝ 5w`��8`���a92�<6��6wL6/��p�5Wz �q;���̧��]c�A�?~��I���
<�Д�ā1\ſ7]W�r�7�3n���M{V$�Ae��	I�F���C2&�E�.~��gl	�^>��s5 ~� jÁ�p��	p?���	a^,�E���/�R(�Fl1�,]"��,�e��p�-�W(�ʻ�v����c�qa�~!9p}���ۯ�i2�n�*;y�V��۲t�Yf!�S�h�ny������?C�]�:��f���&���	�W��в��J	��iR��Sb�x�/g�m9������ߣ�w,�����hc�����Y���B`�������U�4���� �aVP�''�ݢ�����^��u�А>��}��s��> ��Ap,l�H�t�����δ�
[�`�F9!M߿�8�{��-� �ϗ�n䮟>G�s��1��c��{��g����.Z�YV��g����V�N�A��O&�����rYc� ���j��R��'�g�g��*
+%���]��_��@dq/ƽ`��ۏ�l�<9 ��N�q�Rb��׸7�.ؒ��M� �����������bU_�}(���ߟ�&m���A�����Q(Y�����<^�����6���K:֗���� ������'g�:ķp�v<�қ�*Q��<��(F@�� TUAsl�67�+h�����L�[SP7�,y BP=�
~��_r,0@+�	��`���W<��� � �����>7�������l�s�1
��{�����{�QigwFo��T����LN�:�'��E��Mt��aH��T���=4�����;}��O����l)XG;�/���z���.ď�}�.4Z��X��#���h����4�(��s��xC,HGG����s�����w�z	���a|��]�i��B��y�"�kǍ��P�@��R�,�O	+#�R3÷�}ͳE|uK+��,x�P��޽&A�zE� f��ZҲ�u�Lm��}�/���f�>��=�WQϠ���~ߚ�mL����\����S�W���7��sB�s�Wh�˳��7o�N(q๿E�ߡ����~�������_�ŗϸ�]H�� ��3]�qH���ڦ"Pi��..��`��J͜�ZQ��XdWY_s��ka��v��Wlc
Hs�w=Cڞ���Br.��m�x$�jSZ��]J�?ʁ���RT�N��s-�e���ڦ��}��!��E
xo=�T�N0�:+3�8�i�� Py>��\x�B!�2���O������"��Y`yF���������i�JD�yf��cG�$<�q�]�K��=�9b�ZGF?	i��n��D˧�<���*T�`=�:�� ��Bɐ�e2�q ĺ	�8��e��¼w�\0@�۳O��IsR-����酧��[��&Iv9�:CÄ�&/M'3`y��-���Lg>�����D�1�U5c�(^�)-Ao7�-h����\Ɇ��/�-��q���^|Պ�����{�#�_�������d��+d��If�d��*��t���n���I^ˉ����$Lb��2��"����-b6� O&c�������/_����.�`�U^?V ���C���=d���满�	=_f ��!zZ$���9�O^����9��&��k��o~O�7k�B�JL-����rss�.ܸ\L�"	�bή� �8�,zl�_��b����L�u�-=�К�0����9��H��u�`��&�p�zK�{�	e��y�ڵ���sw}.�d1���6ڵ2�Z�*b=�>qQL�wX��aZ��b�sr��ͅx��b�߫�vS	�M�6�+��khu�� ��V2{vV��]�����16�����s��$Z p�2"7V��(�� �� DR��b0$ i����_�0 �H�hk��Fh��5�:ɻ��� ������[sV���穨J��) �^^�J�6>����5��f}?ݶt��V�7��
 `Չ�v/tI�r�_[�pvh��Ć���_x9!��/��3�m�JGi�$�M���"���dB0�<��W�bp�\L<X&�Q���m��'���o�`�GwoÝw�@��x�]{{� �8��?xC�Eρ�;.������T[~����1�4����"���_�[�K��<�d�cx umk��	e�h�C׿\�m�g����]�(�~E=���{�K���˪d�Jo-��)�1��:����l�=��j�����]ӗ�<�*��9��&�f�����f@p�P+��6�}rjdMb����!��MܪK[g����h^%t�3���NKM�w �#�Mvi|��
��٠��r�=�j�zdBp���ʯ��fn^B���2b�������`S�y+��yŔ��'���&���oV����q��`������6�y���<	<	��1�,H\� ��U(�T��m`*|�����oi)�N�{�Z˼���YwS �hW���i�\9ު�I�΂�r$g��[g)���*�q����2P�kA�gmH��١�[܃P�myӖ�U�E�:�b��� �F#�� �z��%	 F_��x6<#��R�)�9����x[�R_§�w`l�M�n\��u�Q�Ա�z�׼ @�L��  J�}��!�Td�H^0��Ja.�@`!��k��S[�M��A�ϴ�+&���d��Ϙ�Ϟ=#)ƍI.q=����3 X�� < Mt�7a��p���p� �M�-ߦt�_p�c���zCI�d�Kf:��٧�-5�����,x��Z�,��L�Ȅ�g	}E,B�-\��PBR0[����V�*<��5`��9_מ�D�tB![�ocH���i�5W� 0���B��TU�ӛ��u�(+�ف��4C4z�߯i=��7�p��-����|�E������x�v���u� �ێ܆��^��;�>[q��9������"�3 ��՛�C��s�6j�#1���mh��;��Zϯ-2�O��{ ��=zx�f�N8;��=����%�\���5�&m5�n�"�b�Bb�X� ��ڛ9ˉ��k�����*��1m��v��N۾�x�
��,K]��ܷ�s��*��y��]�4��|U2� �K(� ؆�Ds�1�6V�9z�J&�y�hKZzip'�1�I,�8OJ�B6�.����z�g��&�s��'���X6(���{�F>FM^"�ʛ�w�x��Z ��/~��O����ϟ��H�����Վ+�A	��.�����V�Bp?��K,zӗ7T�O5�����bA(����K/~�$�@����ѣG<�	C�\Ľ��'4�i0�t@v��n�s/߻w�a%)�` z}�b�x�u<t�yH7o�=f@���� ��ik��N@Kt&@'$���[x�"3R�w/�mL;�m����h4t�ޏ��2X($yD��,|�u?˽l(��As��Ƴ�\>F�ONb������#����po�v���E�K��e�=C@{N��u�y��JQ=���3�+�cŃ%@��n��θ.p�1�NP�P�usc<]p���/��W��9v ����PL�F=z�����m�����+Y�+s�����痮�j�
'$���������O;o�����9^�h�x�tM�'�<E�Ԕ�^�&����2v�����믿fA��B]BjΪ�v���J}���e"g����f���i_�u��*��#�"�߳�?��g$�F��ƿ���b�_z:s�p�(��XgM�q
�|��3 3����M���}R� ���7,� $h��Vܔe���N��MI��ªp���\%���2d�:oK�ϲ|��.�3⺸'����Uʪ��yzj4�b��5w�pK��M����? ���>���?��?��c��]�C�$^Dȏ������駟��,����6�X+��b �jˤ��2C5�9�F�`^��9+Q�S�w�_�I�[ѭB�:c�A�WL2��߰������6=���`w8	֛�#����v����� ȪZQ`Y0����1�	�+���
�mo�"v���҃P���d��Uqڵ��҂��n�0�!eQ��d�ELO����Â�ݭm�{���|�p����_���ZHQ�5F��lT�$��c߹_������kn����C��򓤛J�r��['mk�Ӽ���� {ҫ�)��t���֡�Z��KOU?sB��9����7Vg7~�
�*�Hېx�ߨ��X��ѷ�w���=��ٞ����S���U�`:�����{}�6�\Z0�-LWa^������I����x�>��F��]J��M�eps;)i$��]���=�.�/��"d�?�����s�>����,�����M�V�޹����}i{��_���s�g����ڒ-���uǦ^����r��<�ڜ�c��[���#��p���U(}������ǅ�cI��`����I]\Ȍ\&�ڨ�O�P��Y�V)ud�`~K�/�7]�kA=eX��?�<�}"�׀�+	=�B�/x
x�<�$�J��Y`1���6�k��B�o���4�P���=�!Q���3�;��"���9�����{�g�g��������Y�YH)P�`�`�A��M�d��+�X��� �I�s�/5��J�6��M�0�����Ms��sM2�Ⅱ|,�p� �Z�?�����sr��!O�<��ј�_�8���نQ؈�����a>s�0N�ƶc2n�,���* ���P���]��Z �y��A��T9�x��\8�@{A��|lx�ʆ,��g�k�7ઝ�DQ�;W,\�g(�;�f���ص����ņ�J��Z��NU�v��XG�hmN��qkN�׈j"���ߣt�Ң2��T����2��X������]hJ��ۺ��F�����krns���L�9 �52�LU���	�b_U��P�hw����z�m{�whhZ���w��+N��:�}���׻t�<6n҃����f%��Ex
��W ��*|��MO6�p^��GI�x_�5�-�T�Y
Xr-#����9-P� ���l	�R����=�_ �s�N�pma��Ӥ'��Z�ڡ���8���w�����O��n��@pW�׍�ӂ�s���Frr����Ӷ{g�省��}�h%��<�F�(�"lU��
���KQSѦ����ߍ�� ��v�$�]*�I��:�~=/u�q)> u����o�%�3�0���I��.u��-��j�O{b�%x0%�)
����f�
��� Ck���V��c�����!B�$��Ⴧ���}�>���L�l`��7�α/���?�L�Xs0�G��h]�Om�v p�R�c��4�j�`�i����`�yMB���A�IML�x������I�e�	 #.����=�� �b���w��5,AxU�������������{��1��H'ٖ������W�%Ҥ�c��w�q�o?�]�B0awf�i���,�ѡPOE�6�U=<4��fC�'�'��������g�Pu�x	-��[�gS1�嘂־���m�Ne��>T�M�B��LK�A�6g�6�1-�����lJ[(�S%�	PY��P6�0�4PU(^�߹��Ὑ޷Jj��ylލ�Y�Yt��8��z��W�� K[�?�uEnߟ��4&�
z�f@o��4�[�v	��9�z��e���ɀ^�9�;{��ݹ�%�L9q[ �TY�)����=w���Db���s�����6�I���hM��JW	|A����6��NCC���N�u��O?e��
������y���x�y
�tӾ�P���tH�۶�Eu�&�Z�C�N��!4%$�i��'��3�Ƕ�&�3}��H+�m<ǐ~Φ�Oϧz������EFm��.5ߴ�t�yF|�9��X7�i��
�H����4�VH)u$ɼĲWZ)u$@H�^��Y�mZ�  ���.Щ�t�{_&5���J�*�DQ&Ϗ��G\�D�ܵ&&3�	�TI�� �Q��J91���G�H�
�gS˴L>���f���a�N�p�e��Z0�\h.�:��E��3��g>#pF%,�cz�G����X&�B���4�����U�����A5�ù/Ff����Ib���~�� E�&M;Ủcz3ͨ2��|��ɂ%,�q9� �	��3�x����鋔g\:�.b9ν�^��T�Z=]� �ܴ�ث�,Mu��9�U�A��"F\���#����$�.ꄢy
���~�O-�9>u|�
�w8�k��ب6a= ����������iwg�[ �J)�����Ь��pI��1x���"���_��E{��l�<���I�e�E���Zz�^ik�,�US��;���KnMP����` �v��S�@�V�#<`��o]TY��|[�Q�VP��X?��sUي5��i�6/����C�u$�s ��rK0�h����W�1@�X~�j,e�����xԥ5�WM�n�~ sR�4�\�H�ڰ. ���!)ߨ�斵}��A�.��0�?��9�z��i���O�/ź��])���"B6������c����_���o��$A�(�6�L=_:n( n�͝:5l���*�f��3F�--o���@�%"i�APyq3$9x<�C�y7��?NY�X�*K�	�K�pJK�ϝ�t1Ғ�i����4�њM�>�_aQ�Zs%XD-62�e	���X���d�n$&�0\���A]{�Q�]T+~���-��bZ1�-ރK�_t���.O`���Ҭ�� �
� \�>c�g ��Ge>c:^l���N�y%>�k�R�
����P�;k|�nquy� =)B飰F�~�
F��FK�<�̗�;��V���8b�j���R�L���e��<��6�y��=���1��u��
,�u�/uw���Qjq���y����|Sˠ|k��_ ׁ��]���7�P4��H�>��0릺��D�W|���8T9�c�TBA�>�l���~�l�J�M��, ���
 ����|�~o��X' �v6�k���(��:�|���9�8 �{�<(C����O.�H{1ס\E�5�^����3�?����jݔ�KӍ�"����o�_�.�d��4kZ(A�Ab�^bA�$���F����B�g��JLb��j��Ĕ�֬��v���x� �^Ft������q�T1-Ƞ�!F%��(3g�-U��亾R�La8r)��3Ԏ�dc��|b���3Ro��1f����m�g�^�h��Pٖ����J�c�JI�����ҕR�zÜ�)�v��gB>�ߐ�*'���8@+1�,L(G�n���ii0и���n�Qa��[�����I�?�G��3.� �MP�� Í�`oQvK�^�9����	X�N�Ox�/����C�"�^L��
�A�Y�5�n�o���-ˀL,^�����w�<u^�%2-@ ,ָXv�@R'��7�", ��$P���=Z�.�M�*���]��c�x�y�����~Yʋ��`�2�f�������+��)����qrD��?�3��k�����k��������
�-�q��H��n ^5���U�뛩���',��v�6�SW'���+���*��(�Qn��
��6����3�۲o5��`ͱ��@$.ːXLD�����|	$,.��N�î�y'�l���j��rH�%�,$	<����7w�m'��E�p\�y�KhZ�sr��j�;ʊ{J�k)õZ�R�!Z0��}�
�L�j�+_��t�@d�^!gԜ���0� �x��鼵ѥ�v�u��P�{���	u=���.��ߦw�hw�k��(_�� ��66�~�s�R����14�Dg�!7��	Қ������	L�R�t^z=(�
�?�\�+�FXfI�RkXZ�ޖ�>��k,c��c�(-\Vv���=	�	r��,����c�$�M���wqE���@b	�e$�ؤ�h��G�>(�`����X��RpsY�)��^vΧל������v�-ᷔQmK��\<�+0,���g�kH���=�o��P��#	�a������ϰ�C!�ϛ��mt� ���63�e)���>}!i��-�Čل)�@*�s��J��-�ԭl7곕�_��Ub$q�9.R�$��OH4���[�n�$������1�\�q��>�!��qC����]�wi©��8d!f[�GM��%���]�E{<:F�u�h�^B/S�7y�	3y��[�TSZ�m��^Κ�� �6�a��nql�s�wg��ԣ��m���W�Oh8*|VzSЖ[��n��vig������p�*�c�+������m%'�B��-�؞�c:9;�kh��
�}wݢ����VC��%.����A��W��KZ"��� ���
��[��u�`=톫�# X���"��}���,�����ʎ����bnL�m�3[^X�?�+�.z�*�I�8?����=�t�
�H)�Zi���̆w��l�{pj��*+���k.,��o������c��a�e����g�LԜ�iU�*���u{�4�媯�ג��Z�dU&T�b�_b��D��#@i[�!s���g�}F��/��Q- .�xO�XKI,Xy����;�ߟ��=�pq����k���q�i1�aщ�ЛR��C��?��I'�9U�l �Yp��$P��"`X��6��S�lm}��	��7�����`�H�&f�E�]�A��Lk���t_F@��d� ����v����q±�W�v{~3%$�b�kڱ��/ ���rW;�n}� cb�5��צ>�,�~t��ߍl�僜`yF�����[z���\׮�M��YZs��%�I�ⴊ�i~�s���~���{�=2�Vi5�� �,fK���}٭!dy�6w ���G <�6X�w�{n�m���e��^NǧH�a�������p��{�C�86����38�o���E�uėn�u�,����+z��z/X�)���wcr_	i�)�r�u �K=zD<��$���}Ͳ ˵��� �	L	��g�g��k�@�,��wL��V����}��?����>NM�jKec��As�'}�Y�!�ˤZ_M�_C	���E��"4*wM\h�UQ[��n��K���+|!������{��o�ėP�}�&�o��q���;HB:e�dJVo�������K���Gv}F�$�+`�I�/���pyF�/_�]^��bT����\��= &KK�ss;�
xDӋL�Sk_k.�6��ez��Je[��:����/jۺ�LF�a���Ip��g��Q���	B���h�^�6�������X���o���?g7,&�UH�mG��Q[��� �@����٦���nllz-*�C���Z�������m�%'�SYd��I|��vh�-��C
��؟�k��j�������v�4��W_�����;.o��/�a���,�o��4�]F9�Z)����X����9��L.��|�Q��_�-��v�(s3o�za���+�z��@ �:�fp���6�=��pw�����[�76`1�����7��Q�a�] l������9�[Гg��������G~AY�	�<�W3��5)��/6�_8x`�AI?�s�p9�������\F�o���
[D��G�� �y�����&�ۓZlS ��u,�l����?���]�V���b��f��X���|E�J���~--3�40����U�/��Z�I�ba��~��_��<-յ��\%IokZ�u��US��/����5�u�d�O=H���8�%@
X{a����~G��կX�xa��Hr��?������+���\�Y�J� �tn��6?���/���.O>jb4���D�f��&K�	�;���
.7'�"Ԝ�y%���!�?�*����u�dp� ���[o�k`9��ߪ�&��pE�+6,�$���K��eQ�ǀ���=X<�61�p�2��"tm�֘��GN��iYi��~F�}R-|�][��>k�/��q�D��J �� .�	�.�;�|��>�I<�b
d�K��י�Xm����r���Ҽ�WG`פ�����X'���^�ݲ���x	!\ �ww��Ջ���ľ�[Ʈ�NV�w2=���������q�^�X˝�6��� �9iVf�5Jo��:<���^�7�>��~��;w��Wr}A��d�.��SZ��x���!	M ~q,�ؠ��p#Bd��q��2Bb��Y`��\�,�վy@�?�d믷q�5�M1�iY�x���,��[�Y���/mH-Jm�L�z���9d��Vx�|N�[T�$��E�m�� �/B��[C�.���[2�X���5Y �����"�z�
h�L�˒�bm��M�Wj>����$�_lPt�� ��kvy�u}!�$,�pu�q�RZO,��G:�]�{���� �D�T���7�ޝ�N�x��67<�BbC2
�>�`8� |*'�鰠	�?����^�zI�Go}}`�3)/�2n�5H��.�0����+��_���RL]^"���)2F��zK���F,�{��ӣGp�ދBPƉ�:,,�n�ƾ,��˚��03 �I� ��=���g��W�ϟq|nQL�r!7J 7�]^ɋ�Y^��8܆������|��M7��Y�o�VE���:����2��˳eϑ>�6�y�x��	:��>v�xB^��+�;j��ɩ�ahw�d��=�;�Z�. 4 ,8e8��ݤ��Aݬ�֜q�wD?����������۟��󷴻�еͰX|�t~�T��
e�����'V`ª�wzz���"��K�#��M�Ԁ�<$���\O'�i��e�oMb��-(�kЦV�Y�P������O�6kNs�((lWoIL�<���O�8��TB�Eȿ?�vy��+c�&hEq^=��Sc��	��T��k� ���kW������6d��~��1����BĆ
8��(Y���2Oq��7�nǼ����_F��<���:Ӽ��w�Y�e�I0�c<���෿�-˪ �P���C��
s�'��������������s����P�|�1�JF�&�����[ ɐĬ]5�V`�6{t������_~����v@��K���#�&df \���O���&[ON ~�������#_�����5������nk1��1�� ��� ٖ�d�41��HC��ڸ��M��s�׻[B Ł_��9��[d�n�39w�gG@0I��h
=*� x�)�����/,?�}<����au��f,�p*���rtc�駟�}�^遗M��nb����tK���~�W>��Y$^>L �w2q�gP������Yѓg}�v��-9�����Uڽ�
�Vddn����� ٢�Po8���6ŕ��k+�tY5q�������۟���=y����6�p<M	k�S�zK�*=�v�6�-h��� ؀���^�(S+�y�ɲ�vMN�>A�L/k��g�j:g!��^)�m��΍��9��vɽ[��ݦ��ڬb�I}6��y��U[w�Q#���h�	����B��)�%� p�%�Wdtpк� }������*)]CMkJd���.�WY�9��m1����3������f��A1~�q ���|%)b|����o���M��|�}�Q$V_�!!J>��y�Ƀ�D� �v9�iMsQ��.��p)�Ȼb௻w���F�w_�?��?���<����	��`�	w B��rr�<�t@n�]��	}�������n{F��|g!�4\�|���4��t77{,8�K���K����/�6-y�{Iy�
�ّ-����!3�	��Ҟ�[�z���^r���>��0 ����\ЖY]ȗjlZ`I�;h��J���M�R1�h#��յ]� ��*�%C��,�e�O&'�$B�;�����������g��j{�m�=NvŖ[C���e4��V�y���\�U��{��%5��lȱ������'�ӓ���k:����v�y��u٭���6�yIx���,�� Т^#�Ԇ-�>W��&�,����
�:[��g$�NjE��k�m��<�xѶ���V��䝹��Hr����Cm��6��j�?�M�D�gi����k�+9��֮�%���uW�m���^C:�X�z\&I�`U˯�j�A�'6YSW$<���P����:��:-�B��4 �sS�w�$�{�Ϙ���k��E��=��x�Z�A�k/�����˾O�����yOO$���'��0���Z�|?�ƿ�bO���;L)�f輮= �s~;�TM������.�<7E'��NL�nR|�����nB�@���Pú�8&���,���b�6�5��2]N3v���������b��d�_�`&�޾:���]���U���&\���8>	[���� T�c�>���@�s$�kƈ|m����k���(��K%٤OӾ�=����Fi|� �x ��6zX����H۴�eӞ�w����J�3�����Z�>8s 3��o���o~v/�hk�� �۶7X9SZ� 	��$b��������Bt��y5'E@ HGtt4�7o�����������)���{���5���29��{c�n�<Z������X�M>%��,���,���aYJ��"Vɶ����v5��6+���e=����c���U�I���ݫ��k�^��_�*��l����W��|N]Q5Ѐ�*��OĽY�_ G�"�L@$���r<x�$=Պ�����媺L�K1�k��lS8���B`����_��3�<��Y�A�j�ʌICN��ң�r��"eP�|ƹ�#�@6h�/��F�Zr��t���Z�Ey�Sئ�
��]2��_�f�;O
�7`�=�'�Xu���&�0�뭥��l6���^�p�]9�V����ǖ����Yr�WN�,�b�����j`K?ū����=�g���:Ī ɮ@M�>��_�̰B�j1V�^��bc���:ѵ6�s�����%���[M�l[����K����ۨ�Z'˰�M��Q�\e�W�.�߻�w���M����~[�w���E5n7��R�;�}`�E���s�^�ٞ9�|a��ѐ���)��/߆�ݺ��>D#��Z��TL|V{ΡG���"U��k����Uw4,_�����	���1&��Y�ym�W(�|'��I��
�zb5>�]�$+���|�Y�R�m�p�fqm;O�+1��I���}R����gM-ߩ���Z҅ΛF�~�,�~����;\'����I���g�5�~8i�g�
7<IY����~^���Ε��<�R��e���bC{$9@xx� J�`<�gP�IX�&�Iʗ�\�ު�Y4�� �;	��eח��r�c�Z�����Ή� |%�[��\����Y�;� �j,��A�.���A���7�|�Y��m�y �v����v�w 'O��ob5��d�%��&���<C[h�R1�u-���j���?�o��(�b��²���u ��Yְu8S4g2�����7�	<��-+J17G����mѝ�{���q�q,�cU'�Ī�M�M �wߒNNQ��3�L�5�u�}��][A��MuC��U�#<.^����� Π53qy`m9�	/��(�PbC���Ck��E�f�^g�>����ފ\�*i����l�`"{�[����	Ӻ�,��3U�M��K~A�~}��pH7�l��%\�/$]��m�5�s�������-�����r<�+:9�����ŋͯ'�f`>��s[�<��T�L�N�P��A�#۽_��㑥�ȫ��=�.�{�H-~4��k�I�A�7~L/�4`kHʯ����6�.U���gY����K�D��z�5S����Jy��%�MʁYV�����d�>^��ݼmj�������R��������`ų�����5̔��sו�^��1�Z�KJ_���b���wc$��S��uST���/� E,s؏�O�e�E��M�`���$>��(�R7m�h��oq�뢀����F�Lfy���Di)sh/�"X��7��-����+�ۿ�[s1fڛӘ*��+�2��9y��ޔe]���=8Л�o�����m^b� %7�v �"�AIfB�&V�`||��g82
ų��rrӬ����H���]%�
�D��b�o�[p�g�ݗ�d{y���l��u�����	��qIZJ�6
��Zo��I���}��_��>����r=�r2��dz��e���A��]$��������۟�ǟ�9A��#�u�5Lz]�:��/�Tc&U��O�Sm��E,�|L�U@8ܿ����G�
��`U�6�6�I�=�/�E�Ld��>^�U�]
LtE��Ib�ţ�ߧ?|@�~�����n܆n�
6Z��[��N�/�-M�{1駟��_��5�������l���4Βw�<˙ f[z���/ɻ�_���.'��ݖuz�s���m,�v���e���0�㐍�J�"�G��,}�2��(�,X�	��K��r�C��%A�F1�2�����$=�i$���7�ˢ���Q�ɗ��)�_Ĳ��Ʀs�}b	�Iw��Z���i]S}��Ԃ�g�I�����E͕t�e��Ԥh�[(�K���tX��(-��!ǀ��6��n����ڱ��$T�ȱ��hU��U��q�XC �Hx���	n�hc�p�� �G}�.� и� P�Xȅ�k���ϽHh�$/ų�� ��)]g��&�X���-=w]c�˲��Pj�ڋ�� ����ͺ޻-����6�9qio��\��o7��1��	 ��#ʕ��l�:-k� `P�A�΄�b���R�y���<��iF��n�����-7Q�E��@h��`���I�Ƒ��V0��`��:(ed��' �H~5 Ԭ��HF��`@�&U�ܣҍ�Q=�RB;g������&}���w_|H[n_���m�|/�Nd�H�_@�~����d4�w���#:e-���X�@f����EHӯ!��0�i�m<F\�EK�`ù�S@)�H�b-�����h�e��m��bs�G���Ч=���O���m�O�ry L���֖*�Y���{4g��̀�����Cv���^����$���T��E��������sV��˃��r]`�����O��V(�u�<9Y��R� �� �M�W,�����5�����L���+=�e�	�z����ޜ�$���䉲2�4��>���
�M��Y\z�y���4:� �-MBo�n�u�6�<���,��Z�VAS�hC��Y�D!�z�ͣ��3�O�L�5����ky��5�uBAh�.@z��uVU��_ɚ�^Xp�� Ed��۳�7]
J�E�<`F�ד����|�v����y�I�/�S,���q�T=����|6��u[�}����$������:�PE��³�6�L���s+xװ唢G�r�%�G7 +26����^4�6*�mV}��Nt��_��FA  h�yXAc��[��hŐLB���|b�]�: ���L�����|�!���w�=vL�5��!�B߈��nb�(p���d����ݨ%1����t%@�,����ڤ�ݜ�w����^H���5G� �2'o� ޤ��6�,���6�DG[2�4����eJtϼ�.t����f���o�{�w����n�ܘ�C7:��`��Kt��� �eRȸlw������=�c��̧/��|�����r�οj���Ţ_0 ��K7.y,���P[\�'B&n����E?TrFh�.Ў[� ��Of'�^�K�����_��oǄ�����r>��\���[�'��qx(�$���4��y�Y��|5"PzLJ�%��� c�M�9��-����5�&hκ�" ~5���#�U�yY���m����4.�"mI��Ys�����08�}b)	 ؘ��GF�ѰvTy.�r�Xȏ�#�T�!��V=~��CV^Xm�
�En���Jǘ�f='�B?*��3`��xfM~����"sD� 6\�gQ8���S��|HH��y5ڥ��)�	ٜQ���8A���(oDI�Zrm��=eYI�����y��c ��0w$�Z��n��u�ɀ)]p`L,�|��?��?	�ZI~x�pn��Iu�q�ևA8��x�(���k��}���t@��^�&W�x���M�� ����{�u�P&d�[�+?���!=z�A[۝𼾤O���E-���OnR��gi�gi��>�N�����Lご5:  �/6a�AM>��F���u �*aw���Ii�I\(E��xp�eY~1���)m������SE���:�����>����4j֍)��2�`5�� x���8�M8��<��] �	��)�����9��I��-��˪�Hx%�Z�/�⒆2C���B[��� ⺅�K!��rZ��RV`x�@�̛�;��B�m��X���+{��q&��cu�� 4��4ͳ���* �d5I�܋X��/�״�ǔ1S��Ei��6Y�u���.
l�ܥ���-�%ʹϷ N$�؛^2A� ��xvz-pb�\�8`|� �c�X~��J��Z��	 # �� 8b	�cC��8��ɵ9��d�����R�\w����N�����N+��:��=�����#4�mJ�&�6 �Η�pHG���=ט�� ���E�Fo  V��L�oDC��̸>�U~gӺ��@�am�b:XBm(���b���[I�?�g�}�5�P; Y��ݻK;�;txtȃ��i0�{���3��pf8�8�/K�I4���=���w��?(h��5p �A�0����X� w �@{7�7�\��c��S�$zp� X@��79�q�$� #��e�}|��	�P7u��c5GXY	�%���L�Q�����Il�r�n{Z�@�������v}m�'�譛�FJJ b�-8�v_e���wsiԥ�1�Q����z��Mq��
�j놊�.�6�D3����v�L��X�ύ.b�M� �����Z#$����G;�cK�'%[y�_g���[c���z�v96��<���Ǩu|K�tK��nb���7���,.c���p���cXJQUg^_5�k+@�t@P���ea��1��+���q��`"�Ǩ��½p��g�I�4��ɻ햲=h��[�M����Hb�A\}���(*���?��������}]2�f�I�5�:�=%���w���Vo� � ����w��oƙ�ѹ���&d6�!�h0x(�.�����
N����5�()�� �<'�QZ.q�����C�L����>�^����MBF:N��d{k�1�mnv9�Ù�K1�d/��l��I����w�iɮ�$[�|�8j�P�k��[[2��3�	�&����"S�~+�y��}��tݿ��_@{�Z�p�硚����Sm��_}�r�h{\;C�Z���$�����uF#�^��Ț�$ad [�[�l��.�?ΫR	��U��́�ujNOh���iɖޝ�=�w�� �L�;��vr���]�� q�m��|��p�zC�.��٠�#�M�0#q/P��c�;�u䙰����L�jj��ļκ�U�@kJ�&+�2�Y�Ev�s��W-��s7nr��q��J�K��E�'P�6�.�T��ςP����V8"�j��l� �v���&�� 1 �<�*I,������W��mk��f�K��s�؋%X�u䦼1}NX���KXڹ�@Yqs ��*/���8��q���T2e��~vxA]����0���E$sN�զpJ�N��uC p�Z�	��8!.w��H�q�9�(2�l&*ڐt4FV䂆��%2�����}�cK�`;����<~�``p�'kV�`a������	[0&Řc�������ѣO�K����ho�=o�A�g���+M��&���qO�����'�)}?xlc�T�`;��{��1����Xp�擸��{@e�{�jb?�2�Rw~.ՙ��7t�U�C���Tߗ�i�/���J�j��׻�Z�1�jSPf��H,����������Q4/ې��n,EYL^�*�l��d�q�W&��n�'��x�G���x�1mnthˁ�ݝ-�{g�ܿ�%�c$l	r�?�u�x�}x֞:�{��A�hh������Ջ���Y��a��7/�-�����ܒPhM5�)pM]����,��@�r �N�~��p���}fyI鶧�5y&��.����M.�m�!eZt�E��6�ʬkL�Qp�t�D2e��``��k��a+e�wV�����'��']j�+@   D[]�9����<�u  ���>}�����*�1^������ip�k����gC�� n\+u��wm�Y@Y�}��5�lø�ݻ@�\
$�e�����넷������d��T!�&���V��e^2�7�w��[<9��= N�w�� �|�\E;�4nwy㚐�4��m���hs�=\���
:<�����1hԍ6�h2V�R��ֶ%�H�;/���D����3��D8r��ի�a�ֶܽ����P��ǔ���3G܃�BX[2���Ӂ߸�5��C�4�m������T=����Hi���ƾ[<���t��g�Rb�E=�1���X��>S�-��ݟ�aT��:�cM[�]���ҫ���?�0-+��a�L����
�,<B���1%-�u=�dMӜ眻�g�1%����A0�Ɨ�4x�o�V���3f�@gA�{��/����񳜶�z�� �]���o�2�b^i�Ll�oWY�7,"�m0��ۣ}:=#�=���M��v�������W���=�Kf�+�����yyjr[�\�9�Y@c�y)�ՠw�w�e�д=�y��終�]�	H/��mC�X5�f!6M������)���z�D%�i���(;��W6�2C��*-x՞p�9ݯ�I�p�H�<yH�Utٵ/�
��/dP\����r]�U��h�uILXd��\K �љ���*����s}�3[ԝl.`�^���:yV����j����������3���Ӧ{h�T���Պ�4��y0µ���֏1��A>Y��v�>��!=��I�H �-�l���m8F�1�}��F�W\�rD�uhR�����5��$"��D�-<�`0.,b��~����_��|��7t68���7o��w�}���}���7��z��ik�.��a�Ha�����0N<���/���^��^��ӳ3��������v�mE	�6��DJ�\�Ui(S��	�y`e&_�Dʑ�ڔ�]D`k�
*�~�[E{�}�e�,�-gP�3��|n��٪�M ؓ��<����1;�oT�8����
���7�Wr��F��zq̳^����mI�\6��6��qp��E{1=F�����&�˯AG�lP�3�xs�����g�W�Q���4�qBK�p�2lc��}����t߶z��Gؖ�����}��/�:��3����BO��r�j�9F�S.�Ib�d��W�E��M����k.e�u�606{~6����Y��w�y$�O�`�Y�!}N
lfY@�S����4%ù(��dmE���L"4�����J����x�0R��3�x/����P���u�b�z� �0�� Q�zR"I NZ#u%�l � ْ��յX+�M�����>Cӽe��v ��0,ψ;�g�g���X��:b�n��_�,@��g�ai?xi�3�{~����MX��巊�h���ȭ�o���fS��s�~i��Ԃ<K��'m�� �@�� ��ͭ�9�w����v��5�N6��|�$::��>G'�y�h����p����bIb1����b.`Fp#�ɂE�"�A��k����7��>{�������x��>���tz�l�r �������)=y�����w��9��Ӂ�c�X+��I�v<y�Y?	C�1k�%��_�hM��g�&W���x�����g[��6@훅e��$=��7�[W���S�����q�2�1V]D���L�|8'�~ө�!�j��49�|�_�,�m�w�����zn��5�PDnn�7hgc�M�3�̙��S7!h��p���.�̸�.�S.��f���C{ p�J����o��69�,���L�q<���HC/_�kMH#��L��rA}ԍ����T(iR�ůI�Y��m׺Lj��utJ-"M}��.���60�"ٖ�)�Qb�k,�kʖd>.2���aI��Ƥ�����V��=`��Ŀ�ݺia�B�,,�����q� ��Bִ.�(�:��8r*�'��V��'T�dV��&��tde�)�,6I��눋r�2L߯i�K[��?��!�����1ں}i6i;^6]G+-�%~��9�Z�徚Z-����;� ���/�ᚧ]ԫ���e+DǠ�؍��ϼU���	��26S���hdIÈ(0]d�ca�}�J\8�Ȥ���wh��	�38{)j�N�\������#ǐN�uâ>fI����'2E?w���?�w�?��/^�`8a��D�&$e1�@���$K��P�3���8â���6���F��L�����L���Z�SI�\=&�U_�F�+ �Ґ�!���p�¾z�vK#�C���E4�U��;HHC�(�4��쵃�g��-��P��h:~n"�@i;T�m<qG�J�Y�k	���&X���Tǧs�h���G����p�k��������}A{���?��];��yR���$��[�.4OX�% i�H����j.����|V�ڋ�Y`T� A�:߽����-� �th��<�1�}���H�������U2�z�9�8��c�I", R�	� C꺨r�,�Xb%TW��}��_�:�R�M�/2��L~�!�ưHchH�5ZJ@�8j����wڢ(�n\}�}�k�<+��M$Z�s�u�&��n)� <E���!��?��v섯��~K!S1K~��ٽ�l���8�_Sr|�e��]�+�E�/E�T���`�H���`��E{��ɘ��NN㑏� 7MJ��ފ[���nY(��H�u�5���
���ck	m< ��l�_#"1h��x�k�|���T�&�<o�5����ԭ��	_i
3*{w�Z�ż�!�3�Ǆ_�4U"!}��3�)\�}SHwy@��\W��V�����m9"[ �����W*�-�9dM���tt\�� <�9QV����zݒ]�;��-�(���dn�W:~X8�;��~ϻD��}����7Np;>AB���O� #����~��iZ�
�(]D�zQ 8ςz�w^��M��zu���DI�Z �E��E��y 8�"�Y�fQ��/���N��t!�%(�����������ldG��a,.zPk���J�!X~a�E�#�Bm�M۶��j���F[�>�Ulx^�R�W\�e�W�n3��a�xf)�$q����{UF�ykk�:��(P�Y ���وQ��2�����Y���[j���J���N��@�1 ��y��yP���[��J4wؠe�bF�M�p�SY��Z����<�dE���Mα(Y'c���Xbd+L|��]7�1�wY�h�a���U�K�^Ʋ_,�MK|���b4��"����:��؊]�c��I~���V)}K�v�\/�7�v|��9���Q2M7�\c�濣\V~�x��9��ŮqK�$\�o��+AG{3dA�#�E!鄎��9�'��!f���6�X:9��'���7t�z�V`�"�;���ӧ�w6o���;]��2\�:�X��v�n�b)��
�,!˪ɷiw{�>x����Cz��	F�.g��r���ܘ��-��y(��&I�$yH�ۀ$�<�3Þ�ݪ�M����I���/�XkԾg'�m���IXfa����-�-���2*n��B.dU B#� ��sa�q�9"�%Xg�!?�x���v�Mh#涶����!�"��m���� �}�+ĕ{U��Y ����ޝ�W��Y��>&��*I/�M�[�u�ŨR  e8n�-��jg81���ך}s�`A���okn6Xh⪂E�0�X�bp�o��
�4 ���f�{�S�,��\�x���Vh2/�f��.������F��$`V��&dc�k�FA��gվ�[�Y�&4����`�'-v��8;���f���U ���WA�,�u�~r�0�d`m��7i8VNv�׿%M���xjVވ��M�Ąa�q٭���w(�&�ǜ�����#���!=��5�90�e ���=:<>��<q�m�(t�6~��l��53��	��=ߤ��.=��;���a��xZx	���4��<����E�ggѢ�tV��&��l�� _���s�i%[�ڼ��V�Y�d]�>�,�weȓR; Q2)/"?�' ������nψ5�u%��M�N�k��&i�l��
YZ����4��w��do�^X�aEǽ�L��lR8��Q�k��Xd\�YS/��k-�U@7�l{H�k��Ҁ����'��M"�	�M�@2��`�{��S��i*ж�y/LFkʰ��
��#1ȕm�5�o8��5]�����x���rx^XT��>����j��}������P�|]�4w����u��(~j�}�8�E)�g��5m`�ģ;P�5����2o#��ƋU���н��@�|��һJmnb����!��k��|��X�T�ˤyC�C��������c:x;��ߕ�<��Ё�3��Ft�N��wwh 8�\��͔��b���~c7W��FC��}�7�q������Yy�bV�[�Y4�,*]d�#6nvL�Rz�Xrۮ%;�Q
�Ēw�}m���� �PW Խ�<��DH)E����B�D����x���1w zq�$g����W\���9-�u�L U<�$�B�qｐ�s][|u\Q�@�����
�_<�$�Ze]쫤U(�4n��l�ŋ�ӆ�z��c7 ���j�ۆ��&��2 6"[`2�e�&8H9�OƂ`�`H��2�󠹪�w��0X�M4Z ���ǋnXh�0���E�N�{&䀰�pF�E���w�ޣ͍M�j9��B���Oa��v������чQ���X8��s�%���ژ�m��0ܩ}��
0���D��^МQ,7R��+�ؾH۵�mW3�k���W�'��o�0�[�h�:h~c�r�n�r񖐖GomU<���5��$	��e:��T�67�� ���\��� ��
5��N��ئT���'[i��v_D�l�!�%��i<�u�9b߾A�h�z��#d�/
X�'49����S�w�K;���,Dy���5�ц�<h˄s9B�id����c��gDU�c薮�V	 V~�؋�m�����B��{��+���L�@�xQ�rQt���"��>i��>;�����&YudMY���;D����7�BCn|��ǳ�j;K��} �Mٞq=�@) �ɭ�2I�
�"�1,�b	���/1�m��m ` a ~��ծ��x��i�ʃt�m:����x�e̕���Yt� 0����2Sq��wYw��,;~���Ā�u� �:����I��y��$�.Z%r
@�#C�1�F�=��,�����փ���/���?�(���p����[��@"����^�x�و�(���G0?p�ߣ� ��чn��P��`��np��������������Ξcno��d@/�?���/��>+�xx��<̽�uN&����@�eLr�c�`mh.�O�dಝ#�X&�u�t���Q�K�������οF�r6��L�j�������>�5�n>B~�QA��6&� dᕐ��8���ׄ� ʭl�[�/h�szi�ןٽVΟp�u��+�k�v�j.��0������k���M5O�Z�������n��쐛_�	���BG~�g>�I��n�OJ �[�k0o}!��7o��ͮ���w��N�)%F�z��=^�4t��	F�>��ߡ�-�҆���@V�b�R{��Z��M��f����e��<�*\������[,w�)�����Y��U�&���M}3��ۨ�n�xm9��2FJ��-�$)է?F[�.=� � {�}�� 0(��:T:^8�S���� � ���w�wJ�!�q^Tyr�5��/�����O���D��\�x[J�<'�/2M�/�Q��i������S鸟�^���i=�6�֪�sQ^�n���0 l����(�-`Y꘎��b�r_�(��ǲ�붜�9y��Y~�(���/Q%Z�n�5827-,NSρ���m�Z����"�����,	���~���������{ߧ�-vy~����glY��ꋘ_d� �Vo0rb�}@�?��S�dz��9�b�-��,1���>pd��=&%(�߭r=�~��+�΄���K���4�Z�7�~y4�>M�,�JhVb�K�V�u�� �|�/��* áepU*ˤKL�
Y�}m���q��y=��%��}�<���_���q>م/j�	\�FW똢�J��TY�+ \x�+��V�2N��,�T�H�j�\f%�[��lˊ�jW|c���.����$�Y��o!��ҥ�:��+�Y�%��V)�6�e��f[�:)-0睷�B���ۂ_g?�_#�c~S�S58�f>�rPS�e:��Sb�O���Sbd�����Y��eQ�1���޹�ےiG:V�� ��"q�h�W�ɖ\w�Ƕ�ٵE��m�� ���i��ӉhA�a��m[ɘ7�:-�|R*K�R��U�MQ����stQ�ps ���+�;A�)�JU �lH������4��t��OY����{t�ތ��
::�sKOث������v���vQ�eV[,F0���cD��"D#s������Baac��B|��]����6=�����NO�iwo��< `L �/P;q��h8rm�>�����@w�G�_p(�*�?SL��;l�-#O����e)p`6�Do�����g��:dcX��EІ��\m�ߘ�r�$����R��础Q�iE�{2�� X�-��2��͏3��pI>������iCx�����kN=g�RM~R؀L����)��C2�ۂ'��C9�@˥Obh���m��ݲ��x�f��$��U�J���.o����|zr�AD��� G�-(���	i��^ZV�Z�jp]�ͭ�泶�4�<o�6�Ϛ���l�E-���~��'���ӧ� ��|�'�/r��7|�Ě���'�O�mV��"��.Kϟ?gk�X�lE6��/�fCFX��̡����&пN�ĺb�%�-Tb�sJ_����2GfY�uK>/�'{�� �b] F�.�҃���t ��7C֏6 �l�� X4np�s�n4&~'n��q<Z	k��ո�	B`��N���$�?cl�}8�6��vrrJ?��=}���л���@����<���`�EvT��lm���=���~�/���.�e��Kr��[d����޽T|�u�m�~� 6ܚ-gk��4�1�Wl/b�1Q��#A�[�})��!{� �Џ��xbKO����6գ]h
p;.��4h��UB��v���!�^�unud��`5󻣡Դ6H�7�	++Jn�W%���>&?��Dt�q[�.b���������F��Qk>x
��3��_ѕ�U�[k�嘝�ݎ^���:4B�b�������t������&�n�Y)�K���oR��
9�.#�wRftxt�
ΣK����A��~����	Z��ⲴN�E�e\�W!l6Y�g��<�iwL�Kn�L�tJ�N���}s޹.dI �ԉUV;$DE(�(3�
 � �����E5Uzh�qU���tL0�
Џ熜�O����7��� �p� ��-��{�Rh�I�f�wBնԳL���B5�SϺ�U)H���`S	� v��.q~�{6���+h�FU`򥒴-�]w ��N�
��48C\�c
[����,w����*A16v�!l4��ֽuw�'>�<k~�6��~�� v�h����b!h48�÷/���� �B�#X�����[�ۮU�4;F��Z;p�܁��ދ��u���>#�.�>S6 s�o�D$ؒ�8 ��r�/���;�O0Ɩ[׿��}�b�
�E�T���EIƓǒ(�g���#3PI�"2�׎h狟� ���;&�^�nHM���d=7$�u��N:)'!�;ɸLt)��M�b,B��2Yv	�aqg�[Z�b�p���3�hsϳ^��CP����
R/��=�!	Tɬ�9퓶��L�5���m��;�q|m�e���t�-{�}z�ߧ�w6ho�� ���5��ڗl+�k���U�u���k���S�Yz{H�ϟ�kD'��Z�W/���-��R+K���c��hQ��E��K�W7��S+�E ���|���(�q�8����a%޻0�G�O Hq�����I����`<,� ���%ɗxH�"I,�xVX��爅�2�{)�t%d�?�����0O��\�pSp�-��lM%���:_{ \뮠y �##	`ѵtx<��Ċ���%�7�[��ə��;�{.�"��O�
�B��]�� j�����LX���gAR���=:9>���*����/pe1�m��������Νm��Ga `���m)�(m�r �t��.m���u:3�/����/o�s�(��c���lq�rm�n���Ϝ傥RQ�:��W"�ݩ���elK�1�հ^"M oT`��P%�<!1�� ��	�u&^C6��4r�W�z(�2ԉ�;���~�P:�{�����S��y(���(6�q�"�&�q��q�罨$��N�����!j�!���z��<2~Y��Ǎ��2zp�f𮭮�{�j?.&��d4��v�j�#y�&=��C�;���q x��}R�R���B��ˇ#r���~;����	�q�X��n�<�� ��ZG�ݬ�Gs]���rpMb� ��݋�h���ː7�{���6�G_�~WfX5��UO��q�s$H�r��@f��R"K��)(�N`����x<���(�o a���� z~a�F_@6_W�g�<`}7�e�&�\c��<6A	�f�m�~Y$<d���� �S�T1~5���VA�II7� �_Ƙ1}��˖1Ԇ�Дqr����|�BL�Ů���❏�� l�8�nt��&fH�py�A��??��Ϟ���!�I^�0��v��o�?���h��C�ۖ;�8����	��d|�:�s�	���m����#���VXt�*��_�>F�����lQ��G���F�ޘ�y3�A�M�`1,6 ��7�7��y�:} �>�F[[9����Ւ�E��@ຓ�`�+����~�Z��\�PǍk�rdޝ�+�(�`����W��Ľ���M�;r�e�(�C�һI�D�)�+�1�:��$�5|R<��,6 ]�X�9�+n�䎿��t��ߤ��۶�����;�:��ۢ���:�����f�-½��t2	1�� �փ��_C�mr6ГgtxX�]�{��-����-�� ���MȜ�� �Zk�M�3�͠�h0w�{,#�_f|��O�4A }��9BXBa~������ɘ�қ�\\S�,w�E�����K3��M��p�~��%�y��z������ů���:�P���-h��b��<��y�ݶg��}����� `�,���(���w��1�{4d�'L��p�r��`޵�gC."Ε07����~j���	��� ]1��wc�G���q��%[����l��?z���~���l0 .���&(c"d�u�sk�cfX���Y8�;a ʱ�l9�p��3TU�EN.6��������l�z2Y�A��1��4�T&���cȮm��	��~~��	�C��pҭ�anX<�s�2-�L�1�~{�sʠ�%�����MCtr2�/N��i8S1>q�kH��Uq{�ٹ�}���`�r��Θ��T����c�&���w徥�"5�mþ��&�5�oe���Ҡ����\��I�b	��s8d�.u��ק���mz��Ր� yPvr�^��l�{�H�fB��F����v���9�9���4紽�!�oc�V�--GM�W�|]_V�&Co]��"}1 JV�E(�+��E���OFC�`�Uu���k���m�I{�	�r�� ��]&qN۾Y��y}�H\u����&��"�^��d%�k���O.u����c=�V`���]��\_�|���lJ�1�W{�Gݮ7*IE�C'W��;�]!N����I���[��ѬqiZQ���O>N�`��dXB�9����IS�y�y p%�3H-� ��8h\��[+ 9���l�$%_��>3n��yΐX�b������X����k ��r��O�Ԡ��68��a����6*<0]XwaI��	_��zNH��͘�7�  x�?A��4etd�Ў8ĻK��r�����3>a*�C`)>88���������sݕK��J����҄�4F���lw9��xH??}�>kL�S�kZ�[
�o�n5�`�[z�e���UB])G�ş����쬠'O߸1E����r�8�Ag��j�/���0,!�� �♼�1��o���q��<���n!��Qͭ��lY����.��Y� ��dw�II����q�Ke�5`�m�kR㖥�q@�S?�}'�l�l҃w���è�0�N^P'+o/���4w%G�Xy��W�����l���S��W�髯�з�=uB�}��$�J�2w���:WM��N�M���a<<�:�E@�"V�e�]���+�k�ߥ�u;�y�B;lN�D.��8�-sD+Q�2�:��ދ �Y
���� �	)e���y�Ӡ���_~�%[|���?2F�Ux#"����?�c��9Uj�����.m�dQ�xU�$��AVh���������ǤW:��,���_���E<&���ʒEp�iR�Քv*��M��� ��
В�At�
Ԇ�=l�@l�FDn��#[=����� �Y1`:� ��M���#��x���`x�b S����{hّ�� �܏B��o@ەqi#?A�,�12���>��` ���ak��q<��."_m��������^��V��F , ]�u�̬����xR�`8���3M
�_��Tڴ�Z��^J��j)�l��ʊ*�������pp��}LG ��pQq;9�Pu�����6��pƊ�(DNܜ;:>����-�>� �%��f%� _RJ$(�J�qv��SK�S��.u;p��1�w�����޾�]��
�r ���0c&���������s4�X�w���?���#}���~{D��A��#_�PӔ���Cb��A5\�I�]��m�)��w�,�<� ���u��E��M ]ߦ��E�)���;�&pK�n�ҵ�
���M�˝�6��_��G��$~B��@ ��(}��5,�+l�J_kpu�T�f�g��VN�{^�I���/J#-�u��]��K�|��vV��"�&��r����2L����7 {�4�5kc�r͓ߧ�����]|�c�-r�d7M<�/aݳּ�@qo�P�������'���O���9m8���g �8������ctܢ7'kI��K�;w����!Mə�J�舳m���m���� �Gq8Z�(%|#}���e���}�e'4�g�6��\�K��ɬ��&�)�\Β=�Է0�s V'�##�� +�^�ުϞ[&���j�Hq� �;��j@���͕��(*�����JI+���xE	�qQR�ɳC:9zK{�=����,�YI�"wshH@��z��1�yhT�J�ș���Ƈ� ��h�:�'O^�w�?��?��zK�'C���t�|o��b�~L���=7������!\���7��CdXE.�o]�����6Y�I5X�~��_r����z�ڢڕ����/���b�5p�20Yh���5O�L�#�J�qU4kL0/~���r�?��l}��1g~������D��n��g��eD�eΈK7<�~�u�����_����_Q�]���F�vL:?����MAfM9Eͯ�u+�v,B� �by+�D�GU�Iӄ���0�|��k���ba�� ~��r4����1�E�"�O�-�c ����7���k<A�+˾��QəT3�a{f
.�ı;�wk	h �;���l�R~�b2�G��Kñ��=O�9٨�o9[�بk�]�\d®�b[����բ�7A�r~����ڂ��8�q��=�=7���*��L�j��x��Y��	๵��MP2U%AZL����N������ų� ��dV�;}�{��)�)�0�y=�WIpR/������''#z��-���}�������������m�{�k���#ņ�l�o��r�P:a�K�d��
kp�}Sh] x�cf���Ƌ��9��W���wzv�ݣM*�P��o�L-HM�%oik������?e�`�5J���F���EܾS���}��쮊�>v1? 
A/^�`E	ܢ��p��Lк��,��IM�	2ޢ@A�/�V��y�7�_d{�k�̷��}�)}�t=/���9�n���em�pSC������= f7� R�V�HE���&Z))Jo�%�HZ�*�f�e#0.������.[`�6��a0��Q
�N�������C��٢?���}BR�L�$Y.��fg���[�:�����'4{g�#���!�Lq�L��2��d�IĞ+�`�Bk0\)!�~�w��DLWC���\�Ҷ���\��
����7�k�};�0�Pj����U2��	������F4�E�*i��j3��:���L"������������!%p���L��C�_�_���0�P,���ȟ#�)���NN�rvvLg��z(���y����-e�|�����K8Y{;�%$������߳5	581F�QU �E��,jǃv��ϋ�k���/Q��񊢜�O���'��g�jX�Y]IoR�j���$�5#]'x��u�Y�z�jj�5nr'mk��:�rzL|N[?O�c$e� r��_3�ꫯ�D6$ʂu�wwv��؉e�d�_��[���x��*)<�Jd�Fۥ&0,� �O��*M�话�bٽ5]�>i����`���$ x��UKj$���H�"�([Y��|k���ZA�2<+Ҧ-��m���nA�b\�������ƨle{��+�<���n�	�#�-'��H�����x��Į�����	�[[=��ܡ>�^��-6��*S9A�� ��6
9a}��n�Z�H��j���*�[L�V-�U,�ȨiEd��O+�l���coo�K_����a���,S��������3?iy�K�Dn���&|%��6��||n]j��wgÂ^�:�~zIcǳ xʑ�~nz�jP����c�:���j�f\���s��/�����.o=���� �c�Ÿ`��}�x��^�R����2+\!tB���� q�\ ^�����T������~_����Ì�%�tpF�����|�����o��}�v0V�R;�eW��g���6C�Nݬ5к.�
+�O�Ch�'<8`hA��� o�78,N�1\�gI��b�E����+�I����Hv�/ܞ�A��Ƞ�S"��?>Q�̲��؅��H<9j�&k����@���`VAߪ�SZ\-�Ձ���4
�@�:I�gQ�CKb-�?um �6Z��o�/?�%H ݗ�^8�z���.d^e �~�x��S�h�E]d���up\�X`y��?�wO�yvT2����Ѓ����G���;���@ʉ�p��z�'�)�fwH/�z�K�!��g/������h���=C��2@���ǭ��+���a�d.r�i�v0������g����~��]����k�n!��[���$e5��qOq,7אkRҫWo�ۿ=}��n�]%�C��=�Ƶb��[�7��EF�g%&���9�>S�Z��R��8cvk(Ɩ�Q������o��y֥��M���\Xx�--K��Z��c��
,0"X꘱��v����e
�u��i�3�ZcV�Y��J66	�M\2�'F7Zi�H���㤭�MB�n_[������9���=_�5�I��%d����xS�g1��.J���	C.�e����>}���X��K4��w�����N���J�(���r|g0dO)
 C�ǟ|��� |��
��ŝX�S�ɕ�����)A��P¬u��c�:��ۼp��P�G7 �_ ��4'��L�43��3�&H~�&��������"�z᫩^l��\?��Y��̂��d��G����*�S�d�F,�	)h'�a���˱�b�wT��sZw��-�m�j�mѯ>{�~��{��ݣn� ��J�L ��GDe�-��N����Y�I/^�!`D��'4Md�vǨw�Q�m�[z��[ӕ$P���9*J�u��jy��o<�K�?7��{���G�����ݻ����&X��zV�>9���f9�A�N�&�����g/����d8�f��kL��@kk��j�Xc�wP���[> �`䄓���MI���U��t˭�-QI����X�'��Tׄb[6l��.��{�ߺ���똺�
�P+�>Ǉ�$5�#(��O�M���cy+��Y(��eߖ���z�e�y���T~��cb?��;�z��|b���^}���:��<g0 n�]����g?׬�pm�I��� `M�6�ߪs�,�r^�`�P����k1жr	��b���{f�%��zż�����.1���b#v�O�,�qM]�Mó5Ygy �c���:F�h;��'�l�����{��=����+n�xQ�iwg�2UɶYt�A]
������7>��1Sה�oS�\�>j���5�Q,�0�^�-f��W1lP&����l[�������ד��ue��4=eFT�!�&Hp���z��bP���:O��Eh�s�2`q(j
�ntL�
hi�%���Y\?��C��/?��{=�w`a<q@jD�Ղ���-� x���e��e�-�غG?<yCo���[���������@���¯.�%H��_AED�����5C\�-͹u<~��w����N���; ����/>����u�>psaH�2C"�X��֭��FI
5�7(�n90c�x�b��s�+��V�̇�?��
{V�w�������Ǩ��eN�.�㺑�V''����TP�X_���C))����%�F�I�`��a���	m�Uo���]��-�\1x4>s@��ˀY;���a
��R�|Y�Zj���)%ܸ��#�Zu](h�e^�x�IF�7%W-(��+���S̺=�J�
b�F>�#s8��"
_2�g�����YR��!Q�~�^Z>�g��s�����Ia��V��YYa��I�zD�.���2�2ښP	������H6�P�/r�~[�z���V�����c�1S �*จ����E�#�4Hj|��Œd�j�"�]H�"bp��O0 #&�`��"6�`˨'P��{S2�6@��US��~b �֒�5�'6�ed�}�������ލ��V�{�k꾐6��7��<�Ux��<G
)�R3�i�o�  ����d6N�J��L�L?�P�ش�$�� ^��z��Q�,��&�Vx��rJ]d�!&�4�fQ�f�[�$�S|��dW����ޝ�����iL�5�����J	���֙��fga8[u�.���Ag�-��٠��DXZӱ��t\Ш��!T�5u%��본R'lu��}��d�:��8�w�����҃�>�w׽���	N7�0�2�
��!N̋�ˇp+͝�y:���es��k�e�-sbV'�L&���V�Dkp �60%o��Q�XS�Xm(G��
��z��9W�ѥ}�(�S*pސ�e��;q�T���@�PwxR�8���A��������%MmZ�4i�y��f�Ž�;��SPb�l�y�'��p(r�!�>^��q��q�o(g���YPfg����U�[@K[<[�j�dʵ�z�+E0�T`(��L�*�+[�?����j�Go�/��M�O�1���k*��36��閾�g�G����Y�I�㢊��v���U�_�ʻȹ��%�O Zl(e���s�t8K4x�Y�&Љ߱u8?������Qkc�n��2j��}��=Xs%�@.�+nܨ�0�I�1m���B�1���B/���0I���q�4P�It� ���y0Ǔ��1�H�Q����6
�c��o�1�D������p>�D+�:��@,�5���7���F�d.w�MU�[j��v��>�_|f����g�slϳ{�-�[�R���{.Lb� @I2��͛W+�2I$�@�b�;4l%IVf8,e�!�tu�����uP�Ҝ8�@Z� kG�`6������a�^����0�|2�0��E]���< ��s/0��YN��[yd�^��䟛'����!e�_���3�\Q�������IZ�(i$Rf!��Sj�;t}5���D�������Ҝf�w���ϖ)�z��f���)S) B�oKtLP�m�L�c�G�r��j�3�Dk�tk7k����s7��q�M,�y��*b�P�%Y_KS+@kb�`�\��a;*�'HK���3h�N,͈W�x��.}h��&�l���3�3����xR$�$�����ʽu�Yk?$X�OѦ�Nb�;L2͡QY�=!9&͢$
����<xU�o��h�wq���*�KŖ����}�"�_���:�k�}���3�UW��9���L���k*b�aF|0�a}���6�0�(6X^���,��5��	�V[�b�w� � ��[��/��q���R�l�D���8W��p�|o��������0��f�;,O[��h���L�g��|�V�~�Pl���^��ϵ�b��2�q��Ρ!����3Sҁ�5��Fpf �x�L���$R�2� l^k.,���G�+�P�2�O�r\p>�d7D��t�gB�@垧�ϵz*�V�u�}��0\:o�w��012'낪�1��1�m��e�[K����'�x$a ̂��fv{ד��@��n�ty��{")��i���͈iU��̋�up)=:�����I�� �s��r�D��ziJ����2C�&y
��q4�]���;���4���ݩ��7�(5�%6�SV#"o�`˳��;T;&B����Dj!�Y�B@�a�0�.��8���0s���S���V���pP���G�<'�s�)1����&yكCV8U�iu{���j�����l��*%F�_� �:��� 8T��Y��s��2*�V_�Y����� ɦ`�@���]�3 �$���	�o������B�|=��b |����P�	V_���-�ϺO��m�E�_z۶�����	R��i��M�u �&� ��WTvѠ|i4I�&��۝�#U?���Ą��� <���I�P�ץn��sĆ�c
z]��$�N[�Y�s�E6�J�	���`�N7ak3�┬f.6�R/�U���H"���ۢM�2���u���0
��Kċ�X(N;�8���b/M>��`�i�l��ځ����M{ Z%�*gA��Y��J(�lV�����`pm�Á:]�ȖOJ��w�LS�@C@
㌑a�������1�슕�|^R$.�Ѫ�`l,�q�_|G��g(e�E�y}�k�(I�5�B�X@LhU+�ܯXCB����Oh�`Ϭ�vU�<�$3 97�0�p�և�ت
�w��FV �l���	/�.�Yb�AA�B����-ʀ�f	ϛpgYg�W��z�/��b��J��+���k
x������_rR)���hl ���x����H�!���&l�%@@_�gc��`X �d�_&��m ��/r^ ��T	��u�MT�Gw�� �K�m��
Y���7�ثu�]#��X~���e�D����t�aF�J�}Q{�N3�,d�z*�xe�p�xedK@�E%e��X�s߲1N������ o�t���}J-�O]3{�KSO5T���d\��f�D��;�ڍ�+�DFҠ�Hy���u��m�<+�n�s�Wl�?77��c'A��C�������x|�B����7�[6.I�:��+/e��Ѫ��[���h�}��?�,����z�V!�e�)�)��HS�� ���*��o����Ҁ�+N%
@-�N���,�;�<S���y�H(H���*����u�޽c�rL��~�C*7sT#%���v�wۖX~s.#Q[����^�zG��fψ�S^j�) �y�_�����z$�����1|ƫPP�G�[�Zn�����Y�7�a��샼)��X\� ��4@�X�%>7,I%�J"�;���;+4�/ 8���ko8���l#-3��\��c����G�x�KJ�;��ſ(���P���HVBi��\���0���W�}�e�[�Z���L&�c9�N/���7\Vi���F�8��3H�8a_��sa"�LX ��:r�@p�\����R�5�j��jĿ�l���-���*N6��8*O�uNi�o�.>��&l6OM�qv��V��=�vt�)�*С�\u�-M�%K�n ����tĖ ��8�����ryq�5�R��ƪ�mı�;�Y߿w�!���5��W�����x��ym=�:�$J9+h�b]R4\�~s$����g������n��CPi�{����a(˺��X���h����<zH�����������/�va�S�SCMX�$�.ْb9u�wkm�q��{��ŋw�?���G�~��Y���*����s���\5[Ū�:�Ⱥ,�M@����Ն*]�+W��w�(@��D ]7��$B�mVD����g�&x.,���`���s��Ŋ��_�b�/ڕ�\�lKj�b���Sa[B�����D[ <��U�g��v� �j *�Ql� �Hx�n���+g�X4�%O���u����5Y�1�]/d>x��(;sE�g�v���������Wt��	p�
���%����>�>  �=��9f���,0� ��`��s�-��&ɚ8F�.���Ӕg>����%T��xs�j�W��>���j��3��q��V�<�����^��i%ֲ��B�Z�����V����Ǻt�T�'��VP;B��4���B�Ds����]���TK3���fؿ�\��ʡ"�k���f�0;�XX~�߻ǂRX��`߀�#.���$Nȷw4/���²�po�G�~�����>��><6�ɡ.�e\�י䮜�W�j�=5,(��׀A�����џ��-uvlg�i����A�p<����unK:x�Ckܯ���f~�чO��	}��N)�1 �������
���3uQ�� ܾ��3;|L�G��o��g?v�66(�Xr��s�������^��6}��۸K�����o�;g�{xn��
�F�=�c�^Zwϡ�w��e)�D�n�`A�� �H�r��x� �}]�E�"%� ��n��xS]�=0�yl�ռҢ�ƪ�� ��� �<.�U���wU�ζ����&� ���TU>��)@�p��0{ZE��^�K��!p�	}��/X{V�LYf�|uyI?��#o�~�l������׿�{�o��7F�ۣϟ�hxA{.W++'�P.�gwV\�֎@¾a*}�w�#�|�^F#���!'�h5k��9"�R�G.됒T��[��Ė��X�&��y�\?M�(��m�I�vs+*Yؗ��L Y	���b��?����O-�p�+�'�p��GC��LHY ����V��6��:S1CHi����X�F?�寠����8^]��h�y�J��i����kU�x��4z�`�����K��-ڂc�����aX%�"��!b�X����0+(��
�$�ɯ�=؛�^+ԕ�^�'��b��[Cs~�Q'AN
g��-�!-�E^`A�s����X!�����|�3�����P���YK/������GfU�*w@ݺ>[p���'��!���Mf8��u�V�����?*@�<(Cݮ�h�����vBt]�XH��QS,cqǜ5�!�X�ڸ�����G��l�N�VgE��fX�y ��C��zS��:��:�0˰8W;�OI	K�ͦ���
=������m�Vϯ{����i����(k(�uP�x*[bm�4k�8b+F�,l���i���{�wyyE/_��^�O�=�OP���c�{�&�K�F]:9�������9/�c [,��=� e�d�\�N�_�5� �&�yG�M|"�.ӈ	��Sg�M�>lh]bܖr�_��*��m��7˄)��Q�UտX���E����������^�����ɵ�@�n�j�KD3οU)�j�����N� ���߹�h��� Z��p���
*��9[y�\{��w���;�����_�lGn��(�K�Ֆ�U1(	���GY<��I�=�n
�1eɥi䚔���uq}]y{�� <�5��rNT�tq�#��%PA���K΅����"q�$�Qg��w���	]�c�:� >c ������/��9�JI�3����Uv�Z�(/�#���K�T��*^�"�ͬw���s��m�cӵ�΍�S��Uu�"�ʊ.�.�@q��4��;e�k���!�|��ZW�8AXS?������'A�ƛ�P��}����|�}��q�s 84�W�Z1	d81��?�B^E�#�ly��_9������9��^b[r���^��S��8+����'=��b4�Zs��)̔z�}����bD��חX_����KVP<[�1A��n�s�r1)V@'q1��W"���hM��b��Ǽ�UP㚩�O�]�t�ڕ��3��EX��h�a�b����V�W/_1D}�O>��>|D���v��M;�adaٯ(�g�/`�pJS�[9��ܤ���A^e�Y �\� �+ G���P݄C|����wC^�Sue�0��_��}LlB�!ʺAۊ�"#�9g!������(�T,��KM�=���/h�9B�Ë�L�i! ܰ�NH��lS;�Ь�'n���Z� �>q�*���*�;o{w�Bp9^IX��Sj媐���>��<}��m$�-�����68[�UM�\�򑁥3���QSbӐ=O�|�|p?����w�M2��bX`����� e% �Et��RF���-:AR����9ʄ$$�<�۔uS��$��X؊b�"��d��Fb5	h�0!���퓬}���w\l�n�&$
�`nh���㋿���BB�� ��HH����g���u!�e/�7r)��=뢗������2���s�P���*iG�"Ɓ9�i.�7rې-���Ԃ_�H\��Z��yi�m�gP&
�I�o9���PWw:tߕհ��iE; �Y�a��Of��; �_�e�ǺL"��M0�Dν�`鎰q�k���Z�� ���y��^��"�tU�kK��nS�U.��{x+�m�Yۦ��@�]"�!�-%�[��$s��y�qU����u��m������)����X�藲�6�r�~[r��/ܪ�w]� r%9 z=���wkp����āPRl�����~������#��f���t@�� x<� x��S�+��*"����rHf�e% xS�nh�Ф��5}9':����ǡD�~��;��;���TM����ڹ&�����u���X�ӎ~6įt��o�.�<q��vJ5Xbb�� ɭ������$Ί�3��
��o�[�W��_���P���[���o8� xr�-#o/+�+�sf�v}��`f��\U �5�V`s�F����h����_)$��(�HZ�s@ּ�m�¿�(��;q���@6q�H��Kr7hv��>�sǂ~���>�[��(��m�Y�w�c�s�h��m�RB[��(��sGw�D����n.J��J���6� �Yn�U}X��f�2 \v��F�h+ V��	�^�np<�2(,T�`]�KνS�GM����&d�}&=�9�@'֍'m��/���pNb6�b�&��B#��n��nT�Ą3E�y��Irŉ�b�r\��r-`�1�6�IS�?(�D»`Ӵ�2��������|Mȩ��� ��uT��J;$;hYl���"�D���Y>&��0�����-�(`�3݇g`��/�����MbR^<�^������c��"Ǜ1�Q�%J ���FO>|�`���7����J��]�>��Ԫ�"8Tשq����9������hB��s�=�A0s!-��9B��J�))ɖ��_ϱ�8�� 0�=5W.Z;Y����
l7h��W�}ӮU'�(�Y#�\���,��}�����۶P,�7	�U׏�ϲ2N+8槦~0�2|�r�VnU"����?��U��]������P�_E"�0Yج�$�c�S:_��2F[�u��㬉�@���/���V��hb� ��{U���!�:�.��,ic��n.3���j�}�}���"����~��]\^Qm-*��|}���<efu�EX0#x�!-���.��� �d�ᗟ��Ɩ;�E�y+��҄k@6����]U�V�e�򾺅k1���Ɛ��p��Iu7��^����W�L^_�=v�*�`��L9WĤ��A��CA����T�.�|���(��_�����~�;�Y�2�B�f�.��U���O>|̙�����`�E[�,�f���HDhɿ?�w����F�ӟ��O?q΃��K�^K�݌_���	�7��U>w%���l,���9��r�%ڮ���it3y
�P��]�8��� ����deEb���'��u[�\~�KPHm�U�s���
 �
�Ѿ8�v����
~ς���ٙ�Nϡ.�c�k�6jc1��b���FX�����/"� ����Ҳ������-b��" �H\iy!�6è���*�2i�)8w#hN=hv�"k�[5�X9�ǔ����<��*��t��5K2�4����q�+X|��(.Ѱ\����KN��χK%��P�(g��.�eK+�ն�`u8��c����+�e��ּ(k�5q�@w˨�=�eX���(a�.��	2��k���K2����˓��[;�PG"��`f t���Ŭ�zjA��oŽ�����GG����{�*5�y?�$�R_�l�+��d�v�Ӕ���<�g��B��F?u�V�Ϧڻ��9goOF����^A?�@h��h����H ��G�t")cyx��y/,��$+<W��`p��og�r|�P�^6պHCaxf��K#D�`AaKp�� 0��=�e䞛�ݻ���v��x�-H>G[���V.�S�xE5�쇎X_��Y�c�'�
Ϊ��$e��������9k�|���S��y�c��<��ߠ�Du�N��Tʹ`�|�=�m�][�ʸ�: ��F�1u ��ϫ�?�������I��MXC�2s��Ǝ��Hjãc���k��|Tx��D�c����u��>?[������Y���%
�=&�z)uS$��AO�h� 7ː�jBÑ�p�S�; ��ɴ+��.hb��i ����l-Aq����#�=��?��A/�6X�ESē��[� �N�K��ʀ\2�pSFf����u;�/G�l�E�ϠX%�/�VS���}W���@[������M��vͫ�f�c��a�(�����X�5Ş[�Q��Ƽ?I+�/OM��~y=�$�d�����0ُ6n�=�T$��AR>�R�٪Č�ɧ;�9D���A*p3�4 0�)h��ͶJ�yh��('��Ż�[^���A�j�_��SכQ�:=[a���"��Q7�Q���% ,�6��[����4�mI�>�`i���ؚ7�����7������CnL����������<�)���oc�E ���h��Q"�*����ocEq�$F)9Ŋ��Zq�[�!��Ex�qB䪯�ՉU�t�^Ѧ�B���K2Ҏ����ˊ�"Jֽ#�{�W�/�g�ܾ+�*^��;�����{3�r�5 e���j'j��}���=��wO	r
)��&�|O,{_d-Ilj���j���S��V~�� �N�]�VѶ�/K�V��޽{�<�իW,�cF)��Eu��.��~�sμ��&B���FM�n�� ��~����oy.��C޹��Zp,��Y��Y^��č1��3��v^(���o ��I&�qm=dD�wԥ����H�������ܮR3���̤��6���J�����f,+��N@�@�^>��S�CP�&�c��oX��>g�Ƌ��b��P�w4�� S��yl=m<A/5�������X�~x���}�%}�fB���ľg�e'q.,6@�`���M�����y�,6++����q�S�����)7�ۀ���/��4�ź	���B��Aܹ`]:�E��Ͱ�rlu���{���*"��HX��f)
μ�1�<���c�������5[����7�S�1����m����JQ�BW>����o���+0��C�'"K	�&����cIb�^�yC�|�+�l��d�$���U����?���)�^�� ���a���$M }�rP�Ūg[����kM�y7�Nn�����x��{��S�Dq��8U�~�k.���
���t���k����)z��ߓW|���j�_��ၾ)QV%d�<����/��:S��b��� �s����Z��\���)��ceS��3}q��ye�����Y�}4�I�a�%V������$<�R���`q�m��V9������9l���~��^1���Af���B��O�7ϖz�m�m�{}�]���t28���YHa� �{��=~xHǇ��0#B��2 � ߣ��#ҫ7�f�)�_�m�(��H\L�\�BX\������Ç��G��_�.�O�>e�`$�AM`� ��s|���_]���9�^�(�tm���:��M��պ#k���|��ńz��<��v�h���-�*�f@�M�"mTܮyD(�$)j��uO	;����
(�<��>;�*-�(E��-Y�%=�;6p�35�L�������
/;���l'��U(�Y������j�M���(�O��L��dځd	H;�(�8�{�@�N�������&�k�I�KVI�������{8�) ��ӟil 샇��V6� 0,�ӟ�m�5�W l��P�\�]�����4�Exyn�Rd�ŎZ���j�k=,w�KB����P2������Ҙ��H;e�۴v�cp]Z��:,�h|�^�35ecy% κz-��x��{�_���* ����{|iHW�B<��2���ʽyQ�Z������B�A��X�:��E�^6uK7�'�Ű����������}c�H�ug����o���Q����:�-���o ����X!� ؀��{���>$�� �1�n�!�.% � E�`m}�>��k�x2���ؽ�X,�?߭9K����"�,���J!jX����<������;!����ޏ4�tt��f�c����(�4�~�]�d��>��̂�3(H�4��i�P_F<0�6�����g$�z*IY��l'=4��-��1B�T*�-�Y �m���kpj6����k��1l��=ɧ��, �<��Ii�M���1H��3?2۞<�c��a��%�cw<���$5ǥ�v���C��4l�� g�6P���S�۬yk���۞?��j
a���(vU�a��b;=;5Z�B�aP��%�.��yϟ?g-w�J�tO���E�
����䫻n�6�C3���@U���T�YX0=��5:/ �&�%ڋ�b�rZ�V�%-��;�W�������;GTV3���Y{�q]�k��[c��Z�+�Z�,,�V�7)���&�m?(m��ش�Tx6� ��y�ɓ'�tx��1��>�e��tagM�s�ɏ�$�u?7Q���<y-����/V#)#�[�n�C�oӓmZ��mѵ�fd�;=��-���8����G�o��h�@��IǀJl���?����n�ˎY�eWuH������Z2�+B�_RE���������#�<�Mr��nH� ����%׭���W��F�7o��g?һ��۳�tr�1�{���#�z�o�mj㙑��WU�W�С�/�3s��K\���w������ͫ���2�����X��N�ꚦ�t���N�?��#E��MW�x��}D�]K[EC�w���������O(��8�����l+�_�j��|�7N�XC��a�{D�̑ξ���q��1+`J�u%j���k @pb@0�o�f7���}����OlYlc)��ӯP(a
�w<eW�x�w�q�Ȣ��?n���gP�/Y�AP���X���6	tw�]����f�R��>
���X+��)�=��X���W,���^�����3b���V�� �G�����ik�R��^�߮��@2>�p�n ��E����~V�w|0 Fb� ���G�����KP#�M^8��7i�_�sO�<��D�_�������q�xF�Q�-�g�{^�6�뛦-����[hN����x۝P����A_9>�\R'���6v,U=�R�v�]J'9ͳh�Ce������*��I�*$�J� �Z?�'Ȁzf qj��D�_�x���.��M'g=�������(�G4'l�V�3Q�i�[���R�Y��^=Fo_��޽}n�+��b%���a��V�"��c4�����!e#�,C2\3�1�<����E�V�F��ۿ�צ�W׈s���Va������bc3�Ɲ�;A2�:k�ף��.2��G�vGfƜ}���s�#[�D����)k�r����:������Ke��T�D	���z{���sx���s��'�ܼg�/�ҡk3�����*�5�����6B -�y۸/��mܐcᩭU_�We�����+�=ZL~w�j���'�t���N�쀤_m���+s��-R`/m�����ehO$��t�qh�RA��)uYS�E�`��a�A��R1��z���W��,���������������+�"U���PB�m?�/�<��ށ��!oe�m���2 �G�h<�q���w�~G����J����b<@ŋjT�IQG<V-5fMܵ�h��?m�hK[�'�d�$뽛�l�Z�8s1������9a�V2�L'|�l�����mY�0���<���RW3!����g/I`�ؐn/_}���|��S:7 �����B����Cn��n�sq>2���&�)d��I�:{�lkݱ����r}N��]�itqM?=e �+���G���@'���l���`�w�{I���� ����s�.(3�[˺�',�M�,�Z[ws$�N�=��{�6�9e��,�u 8�w3̳"�ԭ��O�r������;���|E��=�7����rO�~&�'�a�ν[��~�<���Pӫ�g���_Х����i�1X!�`�0��*.:�t~�Z@���}u.�M�!����j�o���U � ��d���mȵ��Y�V�r	
-�}���c��9���mW�w��q?~���Q�)e��0��}�+��=>���ؐSohQ��1k�L�>l%,IWk=o88V��b�"���a;��=+�"ʪ�W��[,��� N�'���a&��C�
@��b��x�&�W�
�?ȃH����#���JY���i���g#�<ýn�py�wd}F�[[i�^)��g�^Yo�9��ݨTk��ΟuOU�r[��(��ӭ� k"�ޥ8<,��O�������)�.�c��dc��k���������ך�8c7g06�8!��=5����%�ׯ� |Nd�2��6IQ62m\��s8�t�Sw�3���pB����iu͝��gCs-�o���+3�3�#��\�1/��]<4L�������_gHtMP_�ڴk1@�����.e�P�������sB/�4�녋�,^�4�Ƭڶ[%|ܦ�'�G3cdp��%ǡ�����ڌňH��bK�,j���m&�Wiw� �NO����s3���6S8� ~E����;/ n�?s�p�&���ʻ���}Ui�}g�E0��8�M���:\�b�M|���K{���}��6	�M����~.�����EK��i_��Ǹn>���\THVŹ��Jy<M���
~��-�Y�Pk5i�6-;��O$�]��駦�i�#�k��5���5Y\�O�^���[|�e8ʂ�:kp[��E�	�}�����!C4���_��`�y�Y������`Zm�׮��U�Q(1P�T2>�|���/�VƱ��뜛�5B������
���}�Rh���ux'�kC[��"��#Y,��7�b��!&@�1K�������`�n��i��Sn�"e�b��������z���g�9B�UX`����]��x<�{Y�m҇N
@�'�j�9b3{���\;0�I�l+٦.�U�-���і���@-a�!Fv�/^����P{�B�럘�Pn0�D2WJ|W���{F���f��4-�6w��*�����M�t����'t5����S3����O/9�֭;k^�X� +I���kV��]��?��[�o��L!c�6����O2
Iu�z��1�j�-�?�%Ƌ��^�^���y��y��XT�ްO�+�M��^
�Y���2�v�-(���B�jͭ��z�s�Vvs����@�rߕW2'��I�d}�5�ޘ[�u���c-��<�NG��.�>E>T�!�Ķ��D�ν�)��-w#꘼����-��I����	�����{%0L��Ӯ�����}q�jl��xF0��N,@0J�	�$.��λ� W)cD��"��0�=��K{�J�E���n�o+����[�I�d2s����r\��m�:vY�z�b�#V���o f��[X��͂,X�r%x\ZR�Y#�l���յEk6�3ܖ�Q����X�x���t���#>ׂL$�bwU��*z����^π�	����uڹ =[��,�c:tx�O�fKQJV7��'�+�	���p�<8D�`���&ߘ �:���E��]��<ӵ=�o���gc��J�,����q���z<���=�MO�E��iQ�{ �h
+D mh2��|tI��z<�����i ,㛻?R�3�;���\@�!�� E����'�|�-�ɘ�0�Y�����Ґ�϶�ݠ�}�2ob���r~�wݢ�tN۾�m�+�4���yw�6%|jU���YY��>�[�9��K�`	��6�b�('	O��K�����OA� �r�S�sK [S��E����Q6�B���d���W�����j�=Nւ�=`���]�E8�?m�Z�����:R��;�C�#
���� K��]��� �_��F�v���1�5�1|�
<��IX�^Wd��*��0.�)T��P���l���{ ��,Ynm �D�S�Һ��0��`�3 ���0�\����4��Jz�қ30v�S��R�j��4��K�l�=X��m����}��ܣǏ��� ������tv~�n�U"qV�><���G����3^a.d��`�+sC��t������0��p�.�4�$�x� �),~(_���ޣU'��b�h� �!y �H�ζ}���Uц��C��qn!��os���R���L�.�,�n��� ��EY��M� o�תX%���J�NZ�UH���iG;Z/�j(ZY�Bn�=��8F������`�3�v��׹.�N��=v�P��Nok�T�v�b���	�Ӗ�bIO"0����,�n�� �P<~���M���<;қ�4E8��N�
�UQ�u^�*��A�Pu����e�;��Ŝ�l���#HR��� ����_�U�����3��t���&p��GWQ3����gJ��7�]�* ,k!,����+�e�C��}�.�(�,�Z� #�	,�(g���JB�]Fbk��ǺE3��4.TmH^[���7������Q����]�~�K����!�e�{B�?8��~Bg���̹%w�ü2�~j@̐�R�6�g��z�i�S��<���K~�~R��
�c̔����SǼ�H�o�/���"�����O��S �{f u�'ty=���1'�b|;���uS�Q'���G��C���~o���f>u8S����5X,|�� d]��������mƂ���,��6R��g��u�,>����:,$��6�w��Um9��~�: /,$H�0 ��O���=�U����q_)�!��<^,��
֤%���-��B��=��*O�����U��V�9���-1礜�*T|�w^ _��M�y<P��Y<(`KǪ�c��A�@. `��Ѳ�	�g��4p\m�^��n?���0{w]r���T͝U�W! .�-k��d�ߣ�����on�_��S���׺����m 4�
�-������&:;�^�KG=��!���E`�O���湸���|D����;nb�ؔ݃q�����
���~�\�
/���V������DC6@�㘫�+z�������t|��S���O8IVw�؀��i��@2�<{o�ҥ��:��-��	���#����������l���sB���n�(�b�B����ѓtr�o@p�	�2�y 쟋�Wy7�bҲ���i�G���)�{F�gׁv^��x�(���us�W>��=�~�G��Ѓ{G�����Й!żR����".4�_�`!�Ge�2�!�*�_�9������8�E����,׺u�Ԧ>m�����!��%_��v̚�e�5>����J��̜Z���B�]J�_t���ж�R�� 8� �z�������e����*Û���D���C�?�hk�*�(��o3-��^%-,� W<62��d)��Ba���� �ue����p٦���u��Y�y�" ,d�bLd1���:�7��u��k 0�;#��f�+$i+�����و^������%��I�����'��%|�k���s����M�uqy���ɓ���������w�^�� u:��w�2 �
p)���:��t�St��н�}:0���Ib>~.o޾r@���������
@�� �/���>��!죞��و�K�f�!ZAe�s�Y�ɤӧ7�(��G��8���xi��&Hd���m�3��59[~�?��?{B���#��2�#����Z?�.�\B+sM&���d�M�A:=��go8I �]�*�(�]��^�x�hG����go�}�^���|�u��Sx.�.�E���p�&�sUr`�<0k���U��W^�jRżz=��E�b˄�������YG��K��^�xx�[���3#��?�B�)6�"1��Jji��6�y�{��F����-�~XVEun�m�K��b��@�v��� 8fE{(�9�����^G>�1�a)ȸRh���I��:������h;Ƕ
 3sG��j1�*̙��2z���[�,z�vA�w�}��Cp}��\\<O�5�]մUk���ٛ;N����sbX�PZe�޽{��]�9[�x<◬�����=~t�ɪ��s�:�Mǚ]Uq��l�
若�t� gl�>�S��GX�R� e�T�>
�������\Oq��o~����?��Cd��M�H��]�n��e����$��:=J{����)'"���z��W�V����OK�f�x���@�w����\y��}���>����W��c#pe���X�������o5��K������]\����3/��g�^ޠS�����.�P�����Ў�:� �Y~����������#��u|7�C� �&���x�t���ڧn�ʬ�}B�VIxV����eo��߽��y n����ާ����PT_��rb�K�*��zl�5I������䄘��]�9I����n�܄}*t�^���u�iĴ����k]4o�B@&ٷ� �]���v�^�s�m�(2l\i"͚��}Z帇.�x�]�����j�Ē݆bECR�c���I����:BU�c`��5 غh�[���x ���PF�AFgX0�V4�E/��9��8q%� �|f�P��ZE�o3I�2<	2�u���ЀƇf"v8�=ҩÚ�ec��m��(��%,(���'g4�I��A�̹枲�/Jh�]�ǔ�Ylj���sooL@/��B� ���>}���A�0��������>�F��MR��e{�R��{|=$���3��S=Y�� u��~�̺:>.�'�} �
N��Bsj��H��c�"���}�x�>�� `3�!��"a� �{�汛 ����q� ����<W�*U���{[+Ǫ�p�u�6Ӭ�K�!nG��S��Xr-_rq9���/��{�ߌ��aC��M8���w�V��=a�q���iVz����Y7-�,w�	>��?z�����&��b�4�6q�=13�}u=�����~�ѐ=���S�* ҄CS,�%z���/l�*Y�.e?^;>�j��3��T��MV���X���n�w�i�i$�+/�P����uYR묄m��n]񠛢���H&�������R�2��Բ�F/H���2�3s2e��}�ձ�rOM�PF����i�N�|��j�)!m�4�\��W��)��A.Q�(��$gX��r��rjk�r�bWI���7X��l%wT<��h}�	�+�Á���yq�w�O��_~I���_3 �%�/�}��w���c3Qw22 ��3>��)��;�3��A/��#��24����ed��A����:�(3@8��Jܞ����,R�{3@Y��G�S��zi�0��32M�9c/�X������MܜUBcX��NL6�.��p��\��Ugel&\1�
c&����'Ǵ�| ���B���k�PD8变�A?e:�����Ni4xE���ޛ�����_҅�U(�RH.a\�90�j6#��
�����>oY����VP��������E(��"�>7MwE`��,�[�?�\f:\����?1�"w� a���jОo[�i����r�^�xO�~zG���\�-e}r������׈mԑ�-_��7����kz������G����^[��j*TT�o�]X7h�
ӫW����)�/��.��";jq�����R�*���սǡp_��^X�g���y��������"����ȗ���XG\�:i�Ko�)&�9��^cU�	ᗢ(»��p�v	������;�F��kK�:ㄲ~r�wq{ 09�+�`��ؗz�?qI%�IA͑vՃZ�
��bW� �/~%�f�b�t1��|��ă�)����1�Gw�w$�:pu~-��9���c�י�ў�=D����,�HX�h?I	Jн��ioĵx'ڂ�<w�����0��9ԅ�"iR>�2�Ź�̵�Vr��`�B"H능l�erIŸ,�d�l�p����&�/�Hrzw�-��?����.M+��Mb\��Ӽз�Tq*�k-(vL�<v��̀a�ز����)xd�%��N�bhl�<�Z��06,��o�t&�'��TŤ������u��u���q'��!��!������ꊞ>��N��ɢC[y��G��t�I=o�u&a��4����޾���`�������m��g(�=�M�?��	�����)�,G�{�}G��r��E0$�4�����!�_9a0P�;�G�M7��,Kn�����ڂݢ��u
.�H&���#Ń����:�Ўv�s�Py�܁
40��u��];��������p���}��-���W� ������y�k�Y���+ϼ�?v�w�P"��=8�	��G���40�/_����`��$Xo߾��� }g �QbF��O��#�{�<Z(w��k�}Bz?5����M�YBW[�K�SK;+��RN�ȝ�w�VCN44�@s=�B��ʣ@����H p�w���$_�8���6�q@X4�v�m0��pU�-f����Z��#�;<��8(�
Y	�#����LX١H�o�ح�b\���.;��ݤ��N<��/� &��������_���&a%�R(e��p`@  �S����W�������g0�5����xO|guYOJ�t 5�	�,�)�6���Fd{
�[�t[kh�[o��Z0W="��u�~��lL@�X����. �e����Z7�˝<V Ϻ�M�a��_��~HO�<����Z~��.�j�Q�-7��kn+�#�$3m ���M q��g�PJ1�<��y-��H�]�_��4a��R�k�p8�7o^����e�o^����>�{����E<�Y[RB�w`���-\l���]��gwo� S���9@� '�mY0$.Ѕ]����ef�����7E����'E��XE�C�Vjx��Y�9�*g���o����b���9?�[���*?ܸ{+�ݧ:��,�;�%t�~������JnT�]& �u��i��-&���[N����uǬ�I��fTȋ�j��W�8�p�iN y~1�6��=���e��������9X7�"�F��=�X����:7�6<n-�JB�� � ��_p�(�O�'I�ns�Ͷt ����5�
 �.��ߛ��b�xP<~����]E��7q��*�kr��[f~,�\� S�	^�wb"�V�ׯ^���K%�%(J,�F��p4��ْ����i��nJI�7�?b��g �ht���3d�bW�:�����d�C�@4��W�;߉׋���ovG;�юn���(rH��+�]8I9:�8 mLq>�ػ	9rV'�a@0�7/���M�G�� ��y�¯,��xl�Wo����l���z���z�p~޸0�-,�Q 0�j����X�do+��9�[ �7I��Bu1�M1�7Ia� ���]IVl�:v%F��&+k@�{Fu}[�Q.l �=�F� *���}=0@���LPhr�1[M���v��Ui�Rjq���+��^�$˸�����F�!�(���ʝ��{C~;tq51`:1��\ܳ�V	&�p�E������fZ�k���tIXrF��g��0�^`&i}�onGk��y3ˢ�֭U���#�\ ������[�Ni���a-D�Ԛg�}�y%|�T(�aI眚�m؂R��U.��j\��Wr:M���%z}�-���[��渀�8���g[���b�Jt�̍ Qm'Ɖ%-��@�������[ߎ��?�Y���֍�{��\Y�k��HRkbU��e���ۺ@��� �=������.ϼ�%���A��l��̾PV����J ���jxA�~��N߽���uSd=��y��ڻ)��\�I0��=�ܣ�{��	�����t��JӼIp�4KE1��������GE�\�õ�0GeA�-?��n���h~
����_|�M�5�� �-��������*&�_0���H�N��r�
sbum��yVW���Ԗ^����s�pK�G�3Q�+;�ں�$9���b���`�X!@kզe�eig^��-���W�Ǳ��^\U�Kq��p��;@2�
��
�&�>�緝3[�A�"���f틘��Q���ZSm#^���6�D�t�Xdy�6� ��y�h4����N�.(��{L���p'  ��IDATǏ��C��Nґ��y�$Wh	BT�K��u�Вv9˳�O������\���AY�����Q�7]���q�&�[53���Yi����-�&�Uoem�+��y��X��\-j�����_�ƶSs�:jc�X�B�X­���yc�Ib �̒���ַX��u?zK��Y��B�<��~F���R��[K�}qk����$�oTJ�}V_ge���
�����ϱVۨ���S�/�D[�x\�ܡ�Ϭ'��m��Y�x�`�E����H��U�Mx�� ��m�a�v�{h⿷Q^�I�b�+��1���Y x�,T$lO��K9^���;|Sq���͋�[M�.��ו-��O�� E)�P5�*l[��8Q+��6���2���K������>�꫿���������	�<��4\���˖�VF��s;�w��b@Ϟ�2���&/�p2[O/�Aܨ`�Ĺ8Q�\���K����UJ�q(Y�o� �ex�i0)؊�������z��{�W+�G�_"ĕ�y�b��?�/�(���Y�l�y���,�|�"�-���(�k]���>��-s���f(�֕	ߥ�&h�4�Y����~Z*�J�~ ���Ǝ9�Y�mRx.qu�[M�[�['�J�J��L,����E�m��֌�����T
�����!+F���)�g-�R�۳2L��g�׊��Q4�[��mg�k�M_�����SP�zg��F7M�W���{"�����W,�U�a8Dݽ��Iӳ_$i�"���ph��Dcmn4lm��n^�m�D+Bhжv����EH����v[�����������s���h�HO?�ý#�6����Aq΁H@���9�����Wf{�ɸ����F��YS��a�HD�PE&�D�s{5</�S����z��y����Q7���8���r�^�� �����g�j�CʲP(�i7~�T,Uq`H��{K������`~�]e10��ء���k�<ks����Պ�6B������}@Z[���������]��m$s���A8�v�p��g��h1P���5V
��pY�"@z"s��;�$-Td-�Ee%�v���{*:��A<�oۜ������C�+fU<c��"�?���eh�mnr<o�\Z��@]�xS� ��#��� ��WT��� p���siR,T��X�z� ��b� ���k�i��8�d�G�F(,�X��qF��C��W3�M��(p]3/�Ρ8���g?>��������s��O���Ȁ̜}�t�>A��y7\v�N��)6�~��5����a���޼}c'��iY�m���i�ȁߔ3J{!{��n�"]����,���r�P���;��:P`��⚷.jkl��'����=+���c�Em�/_2_A��* ��7u�*:�⁩�]e���ZP%��e����mGm)\���y�n��*q6�q����(	EY�˒f�,`�).�c�?�K��[�ifx��֝�R�����C�C�_�ue��q�s)T ��^�K��0�%��(���uΫe�6�ߛ�C(��*?/ ���<���0T#망i��8�h�����/U�4�^u��� u�u��~��M731C�E���p
�f>�_�[��������hL��\��\�£���f�kr�= ���5��h0�7��3 ���~���b�����ٹ@�j	����h!���� �����VZ;2�͚��c��tcL�1��@`�k?s��������H�q�X��g�
�謁[U�[��Pݩ��n�c�_3Ӿ���:�aa��;=��T���r��}<x��k�I��*�:�Np�@a[j�%�VO�9�ixm�
��M `Vc]��|����5̆B��-��<Z�7j[�݇'U�#�& 0�׺������n�=��wMO~��'#ߜ���& <o��Zy�𖝷��u�G15�����NHm���O(����}�'>|X
�e%Q0���s �RԽ7M�}^�4���)���%�I0�uM�@�pPӵ�s��Е���6�`K�\�: �;�1E��ޞ�� �w���� ��(6-�Wd��XJ�CKzz~����Vz21�S��d��q� X�k���Bn;r���%���b�m�'�^�('��K���O�d��S;U��q@����*)�����8&����C�5+���9������;��B`�������|�_� ~���k�����{[U�H�6vG�������I+���#v��^1��4���W�����X�3(���{���������%����n��VgM�KW��M���p��@v���@�|��|X��X�*u�Zո����}�V�uS�۷�3�pH���,J�=y�~��_�o�[:88(��u�e�K,�uJ;к� ��ĬZ�����\g�w�R�PE��������S,�3m�s��l{J�i2���<��sU�g��q��0� �`l��CDEr+P��Yk�+��;@ �������&�I��H����,�s�����|^�As���T+������:��xp����t�pd��lܜ4���L���2mZU
l������7�kps �
�/ܠ��*^3��5}ެNE�Z���_����zA�*yf��i��mh��ol�-�U5?D�X�[x�,�i��&����Rc�,�����@Q����@V�ťN�����oD�������a ~��-Tf���3/����_�M󰛼~���V�~�Yz?c�o�2�<�Z(ѡ8��W���n�{.�6�.e`ڌ��U�j���s���F1_7�Mc�n������J���k묘�{��!�$a�z����%�
^(����،�i�G	>��5Ā������o��69�pd���;�S嬚�z������*uu�u�ݩg�m]�B;��p�%@��To�2QbR��.���
'� &���J��ط�{��oW2l�7*Z��ơ	c�[����!2n��5�뀁l���Y�f�6�8n��_��Գ���ΰX���O�
�@p��m�\5���B����;n�:o��5=n����Aoӵ7fѬ�����m����x̪�1�(淔�A~�%�<�]d]�y�W� >˒�*�q ���e�R5�U�1�Φגp������C~w&�J�p�F���f��rL՜3S7�GxݦR�~_������iX�P�&U�w��EQ5H�#o�m��Ş��bm��h���.�~����EK�G]��~�k��"8�'�r�]�	w`y��;��������B��)>�������XrV���:��x#�	��9	�]��cE��`�f�_�y ����6w�O��U����Q�f�<���&T��U7�/aM��\�L�E���e��X#v�+�])�8�S7Y��LҙqF;5�ϱ�T��*�em?T�E��Yc�hz�\���v�X��nD`/�7��w��,��h�[ъ�[<�1��V1� V	��VA�{�d�j��Ze�����zm�c^�gS8��� �ȷ��m��(i��%�?��± ���=���- ��7똦k	@�n�m�`X�X%�st�w�c��so˚Y�����[�����=����6Ƈ*t^�$/U᨝���]�5mH�r�P�[�q,M� �'kqe�*E_%(zbL!��c޶Z 	���OB���0���jH2s?}�K���vm��ɤ�����u9�6-�ߖq���c.eA��Yk�l��$+�0�@Q�纶
 ��$��}!�5������뢝�a�� �1nI�>�j1�u�t��><��23�,B����]sl���bP+sBs�,^h�$��I�3s���wb�ʏL&yq!�	:�����.��w^f�����-���z�>7[{�`�j�h�mT)!wT�Z��x��Ti�!�߿���%����P�|Jf-z�*���@�
8�@]-"��=wV"��1 �1��1��$C���}�By��dW�P\5WB@Y���ϯ*iP[�y3��~����d�>�}���y ze�*�	n��dU�W����3�����%4eJ�������RMB���y�^�|�)V�#Y��;	Z�dm���݆l��ӂm
0�<_�/�[٢V��GV��zN6��A0XXlSJd�ݣ�c�q��������0�S,�|��Zٖ��sMin�p��1��.��ɕB�_zn��a��]+�Ǌ� q���Y��f�v��٠)d��Y�K�S���* Tk�os�C͆��Jʹ{�lm���wHj2�D��Ma���r�,ܿm,�,�p�7`Y%�fׁ7ܣv�w��	9���r��y,�8u�eX��|��7�P��-���j���?+��P�����d&_|�ǇC��E.�Z�`5'#l�u x��R��-� ^�|1\���2�B������͢eyH[�t|l�E+n{n"y���x.���c�}�|?�:vS��Z7��-���SB���0�J����)��N��p���U�͢� ���*ECx?��(e���A٦�涓��[��Gg0fq��%�R.�1^�^�G�������I��B��9�_>�\n�e�MFe��i ��l�l}Ӷ����pZ�]n��v~�&+B0c�����Et8�5�	�EL�v �I�܂�ec+pf�@K.�|Y�ۅo}q��.��'+.:=�����wߌ�1e`n��z����צ�#so���V+~Ia|z<f�މy�|vX����P:~�VI;�z3t�o�6]�!�룏>�,�O�>e@Z�I�9R��U��y~����Z�w��E���I$��'��?���ߺc�E.�tw�q!X�w�8W�h�1(�cߤ�	=>@Un�!�C�o8o /�ਲ���P��;��
Ae��MS�Q�4���1U�6�pn�Q�^n����(w���>���'��k�e�ç��h&[׀����D��c�;$E+�B% 3j��W�I ��qF��]_O����J�j;���Q�by�)�X�JpQ�`~!��ú,�x k��J\9�� _��26��-��eb��6kxʥ��+/�-ψ|�8>Týe��.�s:7�76���:	[��Ô�Yb�k���I��\���n�N7�~_��@��Մ�v�n�}��:��&h��ϙf=��f1]�� �=R\&߼yÙq��zs�c�v�9KX�9G�$s	��o�=�s�`<g�Z��C�,�;�D�]kA��F�u[(6�.� `m޿MX��='�?Ck��<F�u���MQx��gP����X�[�Z�1�l�Ҝ�L7���s�h���=-�&t��vhA���:5��K�W9=~J�^��=��wYî��Jܱ�%�C��M�������z��./�jO�$SΝ��F��Y�V�<��bY��XSW�o��pc��t�7� �6�{��i�A��`������i"�րh�N�n��_����,�E�);c�����޼��~|KW�#.L_3�A8ш6c0@;2�0q��3}+�gJ`P�?����Wo��s�H2C�{7;.�zZ��/~m�����fS��,�.�2QR���~������-K; |{H�)ܞ�������!t��U�g���`	���ց�*+c��M[���-��*iY���R��v�i�x����]0o��/w���C ���k�{���x�'(L�ؖ:�wb�m��=g��я�MR��7(���)[ߟ��^���+��X�4��D�Q�$�,f�­��ߧ��=��5��]��0
�}���ko�O���^b�u�Zpϋ�w��tl�S��g��M���X�\0s���� �o�����9߷��;�����XDߟ^�ӧoL�:>��;d���Նa��93L;�~%�b�Ŗ�p��Gc���kz��-]_�=���x�2Դ����P O09?;�/^�4�m\o/�//���vs{>�y�u����]�!�ߴ��j|Wu�M��?�7� �:�$%��̺�.15��Z7I�/J! � Fȅ�x0����*Y�&(V����}�V�����P�*��*�3KIS'ޱ[�: � �!�V�/�`B��;=nT��/����n�#{�})���,���Wtq~i�ĈO�����Ⱥg�ܵ$˵dHՌ��y%��?7�}_�x�>3���Sz��=g���v:|���i'�=KE@�,�T�d^���^���=�hx5�W�^��������Ol�3%��=s�{W�
�bov;G��<ewja�Ht����������h�i�xց�P+/�����$~P~[m^�yH����vJF�Щ�Y
]�b�����L�2g)8�=�H���.���u��*˛p_�B��/��O?��>�����]���ut�<�(�nz�����������z���3Ύ.�-��Ibº��{�����:����yМ�{��oU!HU�)�?P���� ��6G����ͅb��_������� ���zzv�`�V��E�-����K���4�״c��:=�(r�֪�M���yV�l����Z�E�#� O\",�����y��	=6���� �ܞ*m)'l �ggb	μ��]�����X��;7J� �.XR��YS�����Ƒ#�߽���f���
��ǋn�����B�����7ߊ
z3-��w��.�ߛM�;��b�d�oW_3ֶ޺��w�`[��p�d3��z�,��s	5�X� �n�l9�m�:jZ�b��GY6��(q��Z&WI��f����/��EI��u � �����})� �s���:��V�_�ة���Z���Z�C �^7��l ���|��3���8M�"#��_��RNmI;+j��Q�j<g�U��ڲ^/� �eB�U�
E�x�r����Y�����b�]�Wj�����������0��6�$��F�]rμ,�ߩ�Q���=y�1����2% U\��舾��+z��	����5zC�ܰaAz��C�h��rO��^�z��?y�s|q�dX��e�����t��ý��aZAp����]�d�ơ��n����Du��/9�j;H�=_\ ����Qae��P(����vSv�fK�� Pl����&�md�WYX��h������&��,��i�g7 �oq|��"����,A��AƖ�E�����Z�W�F�ժʽs`[��C�9K���������_���` _�֨Rf���3����u���%�l���pS�8"1����yyI���o�o��������y�Y�DYX�����jp���^����y�si�o!��]�5���w���K&����	�W:��U�ɂ� �ժ���7ES/�mcq��"��;�@1 ��{'��ч�2�z��-�{���{X�rj��p@����W�ىV�K0v��eJX`�n�1���B��my`�U�i�lo�U��sPT¨x��+-h){�E�c�~�ZE	5��S3~�Q*ϟE;�U�g�u�νK�~��t�ˮv�i_���B�[��J�ֈM���}oj<�ʚ�/���CI$ ��\Y��&� 8H�J�x�UܓXA��
`���~� @�`�&U}�����mr��kĥC�L�q}��1ˊx������4���ch���o��^�&���I�U��,Y�����uZH���\g�wdI	�5�Ȇ�b(�#ߝ��JQ�0n�:�ؒ���K�,�`�"Zf���$Z�_���V�����Bs|r�e>��S�����5����z�����z�q�\C�҃�9>��'� �������Y��&����BS�{��8�ݵGÌ:���]��8�5 �:�p�q�k�G�=H�q;�_i �|��n��I
�;�CTrꄍy�\�H��x∰㳀Ҏn+U�P[�j)kk\V��&p�J0�(��2�����_X~?��s���'���K������na|�r��̖|X�%~��L��F�ڂE\\�1��@r�@�k�I�W�.�y>8>,��U����!�S��L�ձ.�d��;��3��.�9W��-	�X� 0��<|�Ȁ���B��6��-��ն=cm�t���4�Xp�����|h���'�Ё����w���O쾂$��
�� ���/�+����&+1� 6@3���ѱ��@�R�˲��O��$W6${`�?��]�/����H$����	(=e��V��ZAgZ{wtH�P�za��uߧ��{~�Z�∙׍�AN�L\���*�1���n��K���Nhn�碖�M �y����*�6�^�u1h���An���x����_��^p��,��߿=$�S� #0�`b�Q�r.b���B�Z��t�qjZI;K��ֻ��:m����=�P#���Cl貪,P.9P��Z\�W�M띠eR���S@�ï���&2-������~qR$�0���l�F{ ��Ȟ�����GvW���g�'oY�Eϴ��Ȣ��_�yX� x�����>���o�QH.[�" �����K�K5G0Տ>��ƣ1}sy����KևܝW���&�o�<���3�����m�J�-�?;Z��\awtר��U��0�c�ߦ�6J��+E�_�_K�~\�}JL�����T��;��r
̒z�g)�'¨��aM�*gh��3�7�S|�6�o;��'�~��߲��'P�yD����{슽J࿣Փ�s�cp�Ki+�7���l�2����,����Y��-��~�֤���}�	��J_���;�^�b�������f���ό(�AR���[i^�_ ��"���i��� ���
 �o��{������������꼷ק��� ���c�$6���Iܺ]�H|�^��is�X�a�M8���������+z���(�[z�D% \��ϥ��VW&E��{�|x��Ѳn�;�&
]g,���Oa���vf<AJ���.xn�y�L8�}>�\��γ�NQV���E��q��??)��J��.8�E��܌e'�P�,G6l&��*r�����V�rK�r?���I�{$����#���X�b�K�3ps���_|�{qUex��9�&����7������w�"��e#��l���4P�y���Y[��O��u�_�s��<��; ��'�a���@H�q��r�i)�m�m@�7o�����O���Q
�+��Teͫ���B�C��"
����P��pa�:;;�L~peN;=����s ����?<���}fb6���Hm\����j�YjA��p�-g�I;4��9]�]���5V����r������n����u'��\i��[�G���jG*(s��F.�C��>|@�^��F8C��ꛏ�ْ��j[Z��P$5h
�R_�};Z�T�T��>ծY3�^ ���%��=80�{�OG��v��Y?6㋱5[��mB�̭��Q>��uy�mr��y����C�禸Ū}U�:�/�������0�m��O�ϰ�?��(�VdV$�Bi$l���yu�y#�M�ݿ8�x�1M�{Q��6�e��?�P�����Ք�JŻ� ��Iv�J�*.��o�z������Ir�������gR\D�2%�a������G8a?�[��H�����3�w�^��s��j魪�󐘪FaI �{�=9�
��K.� �p7���D^p{��/>��98��|��Q�E��D&-�h�8�nc��"�����O���.j'�7��9��R��4�B9�A'D�0�e�=�����|�և�d7�w��I�f��c,��F���)�'���-��y��wNF쬓>�bk_���މܡ���o�s"�,lI?���w>�Py���K�"�9E�*J0_T�z�K�u@��>'�kwz�ht�{�A�z��cZM��#��y!,��1=GD�ӝ�0ƄG�o!,�9�<7*��S���-WPg�H�<-��]ZZ�9����m����P�ݥz�M�5%��բ�w:~_�:1�Ћ �#lRd���O[7.	N�F׀��! �H�����.��0��T���Z�/�d|�Ȭ���?d�0���+m��dfNVh�zF�N�����CY�i\��	K��8���hrs�Z(�$�)˜�<�k���b�O(��xK�)���%���~E�8$�YÕ,d�jO�z]�y��k�N��g�P�q��vL�7%��x/�������p�����,W��0�2,?�gV��^	�qH�}\��6���n�.L^�W)$�_��$X�S��xaT�ۉL��,�X���']"�]\������b�Er�V���m��Y���yE�攐V�\�a� �c�
���}ܣ��c���7���.�{�GA�Z� ���%u}}>�-��|2𪼣��܂n%4t�4�V���_!���]5o�KZY����E��v��hcc�����W�07�v��b6kuzt\k��w��ó7������S�ޢ���c!�,���)�`9��1�1�1�B�X�ָI,QI�XP6  � �����Ob����,]��i��4b.rδ�x��,�&�XM��[[[���͛7���Y�>��m�,�<J�c>gI���zw�K���I�ҷ�	�D��;��!5��a/�a� ΋�,C��|��P�7VMJ�.81�]5����o��H�8��gV�.���4�w�8�~�/�%ߟ`n�:-\T(KӠ��g��i��������$4��je�X�ȸ�|9Ő��/�Viks�>ܤ�?�O��2�����#/�s%��j�C!���^������@�W��ue��w����J�0pȉg��޸�W�I@�s�^��������c�����=��p�R�Օ%���=}���Ѫ�ime��%*@�C�t��Mj�v/��z�6�ha�����B�D��#��6���*�����1̀�m�gq�,�n��x�9�H�d�;,,���lz��$�iqK#<繞�6��[$s�D@e�=q#6����;-�<�	��u�s����mރ�x,�3AiH!���\�I}o�K��#L~IWQ��3r��'�}>��E��n� p[��� FH��x)�Dj�-x���F���O�}��/)�S�Z����]~K�sY.t-x���^������z��K��W����>�f�5��.��ϹlǏ�W�(��o�u؎�� _x���t)�$��muZTZ����e���=��_��>x�I�����2���{��{��9=*�Z�*�\Z���5E����֏���^з߾��V�r�yJ6�R�s���Zx>�/�:b�4�ָ�t�;��$@r�발^Ҭ�0T��Q�"Dp� x��in��9o*�b���,f���V~$	v���;���u���/z�d�8��N�o��U?khrO�Y�a�M����K~�&��4�q����H��ۡ��
��Z��~�C?��>}�t���<�^���=Y�eϡ�"�AB�k5\��*%�Ε��X�vxt�Hw��vO�	�M׈=6��Q�4�[;BÉ��:$�S}U*���2O>ݡ�?yğPXx^Gm����n5�|�|!�n뎧��#^�X.��/SY�	/�1R�Q�~�tQ=����Y�;R'���=8���nR򛌙�֯��u��n��#������uD���bI�3�Ns>OS<\���{���s���GK�-0��Gw7�{��kqQӐ[�bD�3$X�FhȤH	Y�������=���J��������<�+]��M�����)���8���1�0�c��Q�����yZ\����e:>����s�p�u��A.�zjg�.��'F	b��;Sя�#V,�?�B��Rɣ��yz�p���?���ޣ��K��	���ڦ�[�z�Ķ}�E�]*�=ʗr�sr�Ej���=z�pQ}ާz�\@�^�)�~s��0�i`�߃iӤ���srSI�I��k�1��0,y��H�� �x����������y�������vܝ��68^x����W�N��F���<�o�ѣ�������5�΁�6��Q����]j4�tR;����$X��r�DKT.u�1[�d#k����裏w�Pթ٬Q�7���9J����
�0�4�E:D��#h\&N�]��e��\U��N�Uo��S�U�n��}��#�3�x7j-��Z�HvV�C��"-,T���0<��|���"磏����P�����j_g`�M#���@�M+�$��h�A���xY$۴j��ٲmĿʒ<g�߲��m�1���5iM�*d%rKU@����4����$�_�}��,%�viq�� [XXXXX�hh��o�Y��9`�lu~�?�O��>mm-Q��)�Z��GtZo���	�����Et��X�x�R1G++����"�%b��n��WD������"I�{'Q��?�L�B� @�g��HB�V�<+&<������T)�у[���&���.��sۊMtYKǛw�o���N�f��kC�TZ]�҃���	<_�$��=�Bޣ�O6�	���:>9�V�A�)�O����$8IFMw^Y/�Fvk]k��I���M�L��1j%�E�<���$��V��f�qO8�D-���:��_�}�Z�۠�ɲ]rl�Ƌ��H��n��Y�u�� �98F,��ЪYXL��4ƶ����L���OP�,� G���HQ����igg��˼���iw�ޣ���y����1���jS��;*<Ev�ҪH�nHk�W�B]�T���2��A������En�`�P�-�B�����;��,��r��˻p/�dX>[�+eW�i��_�rV�"������:�����	�~�ϟ����kw��p�S��awy(D��(_�U�M�|�VW�����H�<Ϳ�*�6�$J�GV��w#�z�[�b\*$N>��	�5I�e�%!�f�"�o���q�d�Ba|��i��,����%�9�HLq�����T��u�O�R��'ˆe��,���&���	����tC����&|�l
\��"�?4@~���VZÏ2r/ժ�������l`��{EEr;��wD/^���GtZ�)��9�3,�ݎO��>���tzܢ��"�ꘊt�l)�>>-/����<�)��}a%��gd���l
��СK�?���a&,,��^*��P���
�wo�-���qg���i��W���~�j(%�J�+�%ɭ���Mj�߰|���
����3��E�qN�^�R�}=�l
�z�nvC^2��_����_&9����U���l6�^�S�V�?OOO9�B,��$�&	��I�\���^P�,d��w����8�A;�<����g�:��(+�U�a��%�?�]��/M~Vl��v�
,�S���gaq�a�'��D�:qU�����8��XB�<-���|�B�\W����"�=:8�Ӯ"GGGmjuHm�S�c�H��Hr�ۡf�ͱ�+�Uud�.k:
>�-���R֚������N���q��{1e��	��]�K?�\�
�s������-/��N�z����$��j���	���I�G�^�<E,\�H>��.�j�[u��]�٩����U]E44�-� ��/-Ϋm	!⎴i�\��!������{3��z�@j�dB�gL��YӲ�Rc
�����7ʰ��e����R��/����){��;0��I����N�lǰ��Z G����tO�'�*��R�I0>��^b۴}�]�$
�ˀ%�w75Ө�Y	��Q�vm	��7_pX@,�
Jx,)�Q	��Ԅ�d-%\���F�bB9���%u�\t\�Ndu�E١�i��&����
-��\��+QU�#��6"d��i�~�A�.��m��J���2;G�b�
��z���hw��T����I�<���g�����%ĺ%��P�[>�R�Z`2\(�T_lF|0H0��ݵ�_8��mW� � r˥��>)r��:�<�AGGGtpp@���꽡�q7e.��H*H,�u+�h�&��dL�Xq���[���O^�c����
�����ښ���*���ɼf�O�d��2]���\F%��'t2�:���ٗ,}�v�i��j�u�)� [XXXXX� D��W���A����x�� Q�Յ%'T$�G�f���Y
"G���t��QA\i�c���~HME��j�^W'X�� ���Z4��(���Z�[9�v�YC������s9���͌>F�+R��������F٣��={a�/R�!ӳ�����܂�Bk���A��[��i:�Cy�c�:dq1��i6���
���$� �X@zy�z!�x��+� FB~e1	�i�L#� �B������v��f��Y��k,��˴���V�d\�){ӈ���*�;��`������2s��4K־�p�
zK�-,,,,,f������~(� ̥��0ȵ9sA
�LёЉ2H(��9�����Vbw�6૯�Y�
�T2E�9*+�X��Q$�BP6bB�N̖�M��O��|��䗉��#��ž���]�� 1İ�C�T�kE�= tl�"���-�-�[�a]�yX��N�Nc����J,�@��NL�	k�۷o���������B	�+,� �fL��k�H�X`�R(ۛ���D���_�[m~W�wE�������A�<x@���lFے� �<�E�U@��]fR3����nn�Ӵ�&�̓m�Β`�%�7ӈ���%T�T�j1�p��������Bl'�]�&ð��t�Z��r1a��͸�v����ι�����5�S�i�Eĉ	sh$�	���}VmG�y�3j;���p %E�K+!���֫~v#!Փ}v��e�s5�f2���m|��LmG�҈E��L�����߰�b9>>f����{^`q�v �pA��Wbp�sOV�ai�I��6��Gbkp���a�LK.X��T�oKKKܾd|p�}�E\%>�6���0�n�*�W��\�u�$� [XX�h��X�:��,�����7l�I��2�Z\��8Q��AwJ&�qvT���Z	������X,!�o�ʥ<Anw{�� ѕ��shGZ%szj=J*�pY���yv��q��S�ݥ��^��-��/Z("���wW�ZxA�dtT�u�=�Ǻ����g��IX���gjpi�R��]�{"���$�+�2ຊde��~V䨮�E��-Td1�H��M�����DSX�����3����EzA(����	�P�<�7�֛�=�l�]���✕J�:�� ���m+B\W�����g��W�^q\�G�h}}=��j�=f�f��K��1,N�&�ù ě �+I��1ɰ��\c|\5��-,�	��d���E"q�MB����5ٞ��ꉊ"��plj�i1Y鸬���s��l�i9g�I�����E��-,]&��'�	(�w9;42�*rsx�V$�C������kA2�R۫}�W	�p7Tx�ʉ�P�q=Ez;t|R�����ދ3<��P#�J�����G��ћ���K��֫�D_	���"*::��>l�>����ܐk���y���r�����Z@�u�"����C�*e�ʴ�T�����2̈́9�Hr��j|�NZ�\Y���xg?�e��>K��,�%�G��ERe	�aڃj|^E"�a�<���j��E �� ��+���"'��4�Œlʴ����q�MM�X�M�%[���XsuH�&��(����C�o�`��|��%��΂Bع�74	֐�Tf�rQ�4S��Ŵ�K�4�K�ĉg=���MWk����˸��;*�[-��SHxZ���7F���t�2?��6��Q���C�l��01�%'���#q$j�)-{T����� �[Hj�RK�j�mj6{�+�就O�J���hKqo�������(�Wi�?�`�]���z�Vת��T�x�[d��(�A��:T� �w
1!h/����"n�]KY`��(ɭ�i���>�}�H{{G��\�b!��"����b^�W�j�������ȋ��1(��nR�������,���
+9�૟�^Im���a��U�v|��[��C
��)L�ڌs�)D7�{r[�x^Ϙ� K���� �F���B��:�x���;������b����$U��Q��Þ�d��%���3F�� ����?��O���kz��!ݿ����y�TJLs��ذv_5��<㌵a$XH�9��xn!��2C!���b|e`\B)/|G�;�k����CFү�`�;��w,.�L��tG�/�f��'=�hғ�ht��m�y�։-����?NQ�G���� /H��p�f�g�wBG�T)�T�)�V"��Y_]����v�
9�ڊ�t@����cda�L[��jY��Hz�r�l�yo���jZ�L\���и�0�Wv���8�Y'��g{���J<>n��a������<m�{T(X)Q*�hcc���m�I�6t���@���X(�=E~ѿK*K���=�8�Qh�}���@�b�H~C�0L�00��d�!��ϴm'9�E=<F�ݞ9��Ź��T �� �>��c&� �o޼ab��AA~�UY�h<��:��5øۤ��,,1�b���R�	�_\#�OH���_�"5���s�U�/d�J�|�Ҿ��R�gE�7s?��^#1���{����@غ��R���J������6),����u0_�����uc\��(��qRk�I��8�}���YL�k�PKM~݈��M�ۊ̞֚���;�XSDvmK�
�zm�MO	)y�\%@��z�����1��r����9ZSDu~�)���W1�v���#z�z�v����l&��DM8fK����,��a�3~���FD��A#)U���i�޽?�{���nm*�R�E������WT�Uiw��HO�]�q�R���j�V�ʴ��@ˋv)����z������{�������hRI��q���B~Lk��e.�?���×/_2��V:���8rL�q��[�uciy��#����"�R��O>�k��Ȫ[;H?]�;iXl�v%�0��q��s������=��g?��O��w�<�ܧ)R �O�=�9��~��_�5�aݿ��g	���ŭ@��}��Q�qc�e�%��8m��U�dv�y��LL[���[�:1�9�<�(��{_�~O+�E��Y�JqQѧ����7����bF+9j���B�J���"ǋ,<w�m%#lN�@�z��;z���N�`!��W���Պ���0��E-~׆��D}��&+��h��՛=Zߨ����*U�G�O��E��E>D�T����[��U����B��KT��T��C�`��%EvCz�z�~��-�W�{|tL�v�~Io����;�d\� ��X�޽{G/���7o�0!Ar+$���N���1q]��F��.���{.�$���^��5�qĵ[H�y<�.}�eX���O�D��F���!�e\~�~(!@~?��s��/~�J���f`�l���㸯�k��?��î�`�� M��`���{�	H�I �yI�!B�(�h�Ԛgq%�1Fݫa�b\Q5��V�a6���9�E��:��r|n�Ӊ�^�~�Hn@�����%%*�"�dש���ZZ�S���c#^�H�9���o���*ѷ߾�����]��5� 7Z���pŧ[�t^�N㡐�I]��Xr�ӭ)����sDk�T(�huyA_�V���iS��P1_���y
�\�;r��̩~���ㅊ0{��%5f�wH�ß���zF����V���9"ļ�b*H*6M���A�`����ݞ_��~{��",q�+��5���gi���}nn�>��C��� Ê����/�`+1`��N�3�z�,�0�<�q�)�� 9bcc������~��_�g�}������Cl/�.i9.�_~�%����-+g׍�`�%x����K��������|I�����Q�޴]�.��,��f�I\�Le�i�9�	Y1Y�
�0I�j7�ȃ��$�ǃ��-6кw�t�<��z�0W������-%�^P��E�C�)�ł���ds�Y*���@�K��Mz��}��z�r�j� hl��$8"�Q���4��XIq��1��'�8/�7��3J!��S�E���~A��<ݢ��2'3sT��.�Y.x9$�&_	���TK�ا ̓�����>}��W�՟�ӳ���ZS�{6^[
��1�[L�xM��P$����l�Z\X���U��W�J��q��B���$���B��1YY򴻻�����Sܽ��Tׅ������ڑ���Ǖ��f�[X?��c�������7��7�0y��$��`gg'V��z|��W<~��0� ����Zlaaq� �A褮�hy��9-\� �#�pI]Ƥ�vd��/Q@a�{��(|��&Y��쑒�s�-�E�f�Kq�G\7j�*�t�D���Qk�o�Ύ"���Y�Xp��)��j?</ X����[����Nӡ��N9zI�������`��k���
�N�����:�͞`}#`�J��0���3\�߽ߧ��N����O�ɣ�X_��{�~���FxG�����ct\u�<�~{@�����o_гW{�x�������!���Т�$�3އ ! �H*��<x@�+�� �bI�$���w鴈�0�wfb�	�p�G&h(wq�H�B��ӧOy>�V,���������˸�,7h1.@&��-������?��?�����-�f=�4��n�e�0N�? �p�	�LXlaaq+ /wLtpÁ�^�X/ZG�X�E�/B~L2�@��F}C�`�z9���q̘/��{�c#	
& ����ݨ�a1BW-X��B����f]��'��M���'��_	�8��i�C��{����.׹��\�㺱�R�K��::�4F�4Ԑ=����~�~|�GR����iw��j�]r�[�-��.y�t��f���Wp�7���}����^|at���=�C�k���zv��!���q�=X�����+Q)��v�]��5r��.'3kԑ�K{�-�����_�H�^����Sjt�'6�3��E/�{�����/\��.A�(�KlQŰX �0�_�"qT�P2��O2|G�2�1\3����m!+H�(˯i.��ܘ���dF�X�8C�����6x��'#��<���qpl�}!���$F]⁓��f,�$������ /F�|�م�/OyiW�a�q�o�`�aB�I����MQM�����+�mI�0'ץM@�[�I� A�%��Mr��u��SQ<&����3�p��jztrL��9�zw@��Uiss�v��hmm�����\괚������j(怾U��ͻ#��J�lR��UdW=_�&�~D~i��������x'y�}���뛦�;køt�u�q�c�l�\�
5�߼9��{O[�Kto{U=�sT�x��"񙣈�����C������o���7tttB�Z���;������	s~ ����C̉ �D�J�e������|1�R�E��q����&n�&����	� ��	���M,�P`[��b�,�d^�e�!�$^7i~f��X��P�`aE�ZyL�͓�&1RȽ�w�MIZ&���[A�O��|5	,�����)^� s[[ۜ�/NsB�&6?�m��d�O����8זԢc2�=�4N�ӈo�y��YWm�Crn��4d�I|O��Ɔ���XӚ"�'�}:<<�����[�ݽ&����|U�n�����o��S�Fo�*���?R�q"�f$���_!�F�/�_�Q$GH�yQ7�O�!E��P�T;��Qd]�}�Nk!�������q�vw봼Z�J5Ϯ����Tߵ�=E�YzsH�~xM�o��?1V|W���z!Y<�w�${z���`y7���BQ��(~Y��T\^�{s��2IF��-e�ǵ�@~q����k�Y��`����#�M�U�D�YSo*�b�ǩ�kBƀ��H��$���yb�-����5H��&1�	&I��0)�u�웶�$n��&�߳�zH;�X�ۈ�K�V� r;��.���5�{JXn) ��p�@��� 1�]j�:Ԭ7���.��7V,�����T\M������uB��ɒQ�N>`Aw������z��R�wpB�b�rW{D]�W�?�B�[=j7:�P��Wbae�����[p{�!� �s	�/b�a�\T$dP����rAR:$X�T�Nk�L�٘�T�B�	�#ܾa������ c�p?�  ��q8�E�D�kk��Lv��ګ<�U� ���\/��k�d3�O�aIhy"=.,����5��N�_F�|^�ud��e���}������c��6�g��<��s�e����h(a�͛���wyW�-���yN��+8�D��}�n���`E���9�b�JhXգ��X`�Ƴ%^-.�iaٝO�mʝ4U��#xJ��LwQQm�T���C����=8R�Y	�Nv���ɚ�	0\|���j�Z����;IZ��a)��X ^#dp�Hr��5]n��-�mXz�d��R�����>��s"ȹ*�/��u!�L^�<в����C	���u��eQ�o�g��s�kz����vK�-,,��]"�.UI���,/[H��d��Fww����l�_&FR�&
5h+[w��aM�B��|A��v;��T�D��ñ�A��Ll�5��4�W�Ĳ��m1mI7��j�IW�V:���qC��s�w�����+B��S�G��Æ�Cm�a�bA��"�~W�at
��^�K�g��@f���7qi;$���O�	�<���Ʈ� ˰�#����M39SR�*�Lf<0ڏ�I ��$�"M�n�g��"�g{{�I?0�Y[[���I7뫞��K�`޳�p�$y�I�q��'>��{(��~��Σ��� ��c�%umYך%wYlaaq'0�iV;L$ݻ&9�uYW�|�y�q�}�ݏ�i����_��hB�."�.� m=t8����ؕ�yvcV�r(���8�0E���T�}j�<;gۓ�N���t=F�F�0J�F]�:������؎��8�U�� ��G�P�{����3���I0�#��@o��\Ga�Dr',��"�!���sIX����u � � ΀$�������uåȗd��'U�]Zr_H	$\7ܦA���Ʉ������q����.�H.��Es�)������VR��Uu�������Na�qL�y�뼎aʃa�ֱ��J0�2G_�	/j�B�@�P�6�C@�":�"ʆ�J����:y&K��!�A��%IE��HM�-��-&Ǩ��j�I��J2vVV}%����!u?��(��E�3�T�6�-ܡ�9�_��u�_���2���	�gXqA�|��S���%X,����c�� 6:i��f�b!��H�/X|A\�n �D�'!��<R! ��@��{��a86��I=y��V����1��6�{=��/~����Oc���`(e=7N�	�1�V2=�ܶ͑����-�����dY~'(�������^Ƶ�Z0��{ϋ� Jp���Zq}��'���2i&N#Ѡ��Q��U��*B��M�	c���0�'��8���U߉L�,��*�]Եn"�b����k~d#�+���8p}� �=���	��5o�D~KC1;���̀�ͭèP�.e�`�р�N_I%��������*f�b��B��|�ii�"E��hZ����䔎�����>�&�tK���,$M�I�Z}��L�vww�ހxIR0��c7�oY���(/%J�A�csNֿ���w�Jx�|��-���a`����_�� [XXX\�B0�Ƅ<��[���Ÿ���4b�.�\��љ��)X|g����u4)������ͽp�#W���Z������L��9L���C�U�?�X����^g�v��w� {z�/ٴ���� p�y��Y��t�vD�H/�ݥH�e��fE��Q�p>[��bR�A_!bƿb���N�����pZܧXDA����H0H,��$Q�!	��B*�賕��2��_�:���o^3q�Z��:�t�d]�8�ǒ��c�a��5A��m�ݻ�Ǔ��Ik�m�0�&�w��{�o��o�|qc���wr��<
d|�"d�7��M���Td��Ӕ2iפ����������
pn�7a�u+�^����D���e��ڬ���ԍ�>S�����^tL���Ǝ!D� �};XU7��ۗ�Y$�@�����a�,�BR�*&����G���X�=GȀ���D� �ޜ�
���$V7�ʨ�D@}7TύK.n�~�C�([��X�����У�#& ��I�[q��Jz$c���H-] �d�was_��^Ƴe���K�����$k5�}%�����7�iK�q���A����^�w������e|b�a~��W���B���/��ĕ'c��6��R�����ٳA�1�6S��o,����S���5�B�$���p}7��.�"�%�眈X�ni�7'�S$l;�۳�-z|j��B�c�A�n	�Y�	���P"�i�-�N�
�a��7pm�ub���w��Xz�-���p��=�=���{�y�Aj!_ /�K.��}��0ݎa)�g@H��c ۍ;��/gC.�L�/١�R*5Y�ڬfl�y`�_��������(�@�^��U�"%�;�:�+	�p� �8&>/;Ǭb���ץmg�T(�_�o ���}ܗ�,��k�gI�&{d���j��v:@��b��k��%�1�w獹���;7���7��nF	biq[�˙!Y�j!!8V��[�����ˬI���(�xׅY�N�/��B��*ǿn����"#��-�y��Hh�+:���%MȈ����?�.IjŅp�Z�� �P��J$-����%\�ay�����$J'�"��������D�*�B��M�}��Z������2[��8�$�y�qϐ}�e�ngg�	�8�/~7;��F)�gF��ߍ�1�AQ�Q������(��/}e`�-}�ɲ��@_`|�_����#�r,�������!�Ҁ�x+|7���^�@��Y����}�a�3rD6	�X>��r������å��!�u�DX@�ś``K���eC,c��;���;0H��+�S9rR���[����
,�B�/�%،%˯i��x	�F��;_����d��ظ^\�k��S��T(H[�,�&1L.i�i�JZ��>A��
T?BQ�E��L��կ�ѣGL�)�ח��[}Ŝ�w$����M����	���Hk�y�%��i�^��}ʹlB`� �����$�����!���sb����a
�l�c��a����1�`ȉmڤ����<���Ӽ��y�HX%����a�3�;0H0�EA��zL��$�3!��>Ǚ��c�T�Kb4�^�ey�$�W%�Vn�Wb���wqq�Jꚛ�f�g˸���P*�����>N,�܋q��7	Y�=cVc� )��?�����K����J�4 �5ݦ�r[���T�Թl�K�-,,,���~]HӼߖ�%��_�&���-���ǏYx���kOb/�R8����,�������p�c������g�#��.���I@�%Ȗ.�Ą�q,	�*���I�4�7K���̍JV%�Հ��7��hkkS��9v��9��`�ɔ$�V� MY)���;�ї_p��{m�(�M�_��W�8�m�'Ex��d�;�7X론@��������>��C�jXqя�C����.�a`L� ����[��C�u��s�,����0'�8Ki��G&�ih9_�JQ�^�)HL�q5��&�qڑ��,���]�P����6`�-���x� ��3h�>9���d���}5���42���qp�k<���,�B���_�����B�eC�B=�
ɯ v�=<d��N�k��Q-�O�U�3�k4�0�����oK9�52.!�Ūb#�~��YD�SP��&9�&ے6I;p�G�s��x����d{���1��p86�.�/�+f�=�,���&d|J21(�>��3V�~��'�w���o��bd���?��O��7ߜI�(��P�`�aLz�k��`�[L�����Dт_f������ �n�{��uRA��$��0�Jbd
9öK;�e@�\O�]�}�Y��Р����)�̙�Ģ#�Ô��m��Y7Y�8�OpV^��˃u��$G����Z� �����jq-֣�øL��xS� ����<�+�,!�x�A@0 3sr�s�M#�b�y�ҊOXB�l�X/
7�6�$]�@G����9�G=b)uR�$�1s\Ɯ.��$
E����R�'k��Tɐu�7�Be�����G��O�c�_��_� ?}��6G�������c; ���7)�4g�:';F�`�[������/N�Y¦E�/��6��d�4'P�8�D�Ap#:�x���9�C`�.����6Y�L���*Z�0� 'a	��0���(��g�b|�Y���y圃�U�7�	B.N�%�X�`���j�Sd]N��Xc��@�q1ρLH&�4ϠqHbRqhBb2AA@��
H�d�B�(Q�J[�D|��'�=>���+�����ƹA�d۬p�� mٕ�*�1>��<���ӐTH΂��E �vpO���_�`�K�C����oNd���K�Z|��A��)n��2۬bp������V /G!�p��D	�"�ъO����,L���ɑE�s�"�&����fq�L9��0M�	T��H2�ۈ�=��q�b������D5����ǽ-�$����>[�o�G��N��H���V��GO��	�љ��T[\6�P�=_�H��ȯ��|�F=���Wb;1���s��B%��9^L�d�UZ��S,���
�UV�[_L�4ڏym1��\��p��/����������������wϞ=���f�g�7C�̸s�%2���B�$�y�����`�[�d� �}��_�Bg!���	ׄ���H��ysH�( t`�ֆQ�w�˞��
����^wyֵ�Ũ֦�)�+��EL�	�X��x���u`��.�F�b�b�	p�O���gϛe��[
��g��
���J����x�$Dq���-�A��/���|�yB2�� 62� �r�m`��wq+N{%�0�k�jR�c�z��=/�7���<0���ޚ%���S0f�y���������k�;����x�8n�S��l��5�w���I�rK�%�wx	b}��9��΃� �@R!�`��	t��X��Z���
��wh����I�!�`��0iǿmVaS����1gDq�#^g�hjaW�̸g��Ҭ�����f�3ޒʈ���atv�887�]MV�;��A4�p�X^����ea{�>K(�OW��M
����a�iۊ�R�v@(�.р�mB�,H"��8��c�"$��d�/���E
�I����B�-�\w��S���9�M퓜"���r;t3极g:���~�Cqg��XI�駟�Ç9Xb�Y���׌���fޖ�;���ya	���ŭ�$�0-��btqJ��D,���0��`&�I&z��d9��cda��<�{p1�@ۣ[ֿ��ǌ�2�����l�X�)	�(&<gy�1,�&-��i��翏�'�.��@�Eq�X\�O�Su��}�Hh���6�E���G�}fƟ��D��w�3�������/e�@���v�ϡ�?e���Q2���	$a��K�+��U2�K�!l���X�����!m�[@�G�21�s�y\�%~r�1�b���1����y*0f������B-F3?�8��Z�-,,�,�/��`q��S��2,���#ߓ	5�`N$f�ͬY���oo"�A�ɪb)�"'�W��iirԷ�Q��0�[���r&���4?�:2�"S���=���,��,���A��� !\Y�� ��Hcb���1�_S��Ǧ�gsD��m���M6"%�x��{�� }�H�[q^9���-Dgww�?Q'X\a���Lђ�_|��8,� NB�d޺��;�_Lu!�漒�cL��w"ݍ�!�}�x_�=�������\)�,P�K�4�W�f�����e1 ��'缷� [XX���0���YOu�^{�B��	����� �Q`�'Y�a��`��6��|[�j�@�!�\X��}�j"��4����H�W!����|Z�_�h���)��'�L�}.s������S��ef�_�y-��#���~�;b�&ۨ7��j*��d��0�~���b,8�b�k� ���8�u���5Xm��$/�6=�YJ��x/���Vd�D�y]�_S�*1���ĻA�!�{�V/��]<�ĕ[��4I�+,8,�R���Š��Zg�n5uL�;��5��A�T,\��>y��<�C ,��?��yZ[_����g��R'}����-�W,�R�B*�*%I���y��`�[��L�Ү}}1�q�p�kېS\��b&�H�q��"�ȧh�e9��פ��U�q�}��g	&a	��&��g+p��������[�xOׅ�%I?�]Pu-��w�o��cY[���B���igg�c�vvvXs/�!@Y�gK�E��8dc�
���=ƵOz�X��{���������[%��+�a(ѷ �.$�rB�������3n�ߡ��b�/��N+P���.����`3����'��e�͊�1,�b�5ߥ����I���|J�d]@02�Ģ�bѕv�� CX0f�.�g���]����K�=�XS,��!;�=M#i�����O����7���?�o�K������/����?�����JEMQA�,��S�!�
Y��������� ¦�'M�8p?�A��	K�-,,n�K"1�U�	��q���b�Il�ۥ��N���_�P��
���'���He)z�Ȳ�-l ���<G	��x1����Q��J���1�sen��|���W�W�����HS��Źf�~�	�i�8�h:�9�~�3a�y�QrD��,�� �]�]iLd��U�Ǚc�0/�Ͱ��57���ﮐ�0ryNy��1���Ϧ��1w�e���ǅ~�w�$�plXyQ� ��$H2;�w)g˞$E�E�@�d��dh\��e�� �x�{�Z���~�j+pֺqϛ��I2q�$��`�G~�嗴y@"���sX�Ņ��kl#�І�s}��v�K(�7K�-,,,��j|�a
$7��k"�mp4À��w1Xu�	}[$��K�D=��)�Y~}�L�AD�u&�p @;F8F��Y��'O�����s�Њ��P��K�u�ǵ�
	�
��,Y�&���b2�<���K��؆B���{��;o�:��>��r	�T`��j���̷ ���x��0to�;�b�XDc���� ��V#6X�7#�q"��L�e*r�A~e|��]�ö���x�ɺ��}�	F�����Ax�[ʷbQǈK�e����a�+%�����8������c!!-n���a`b�_d��I�4�k���cE�AFx3%���z�1��EI9�.�@vss�8{��κnuR�$�M����L7h!�p)��DD2�j!���R�K$��(F���x!���Hc���x����b�q$|F
�~������Ըum���'��9���t	��kȌ�n�%Z,����@~A|�
�M�x�"�B����!5�+E�t[0����]�"^���������k�dX�%���-����!d9�I����H◄%��
���0������zlY�u}���AVzj=,~�H莄6! ¨��Uۄc;p|N���9T(إl��;�-����ѷ�~K7E�0m��ybzǅX�`�EX����&nd7]����e,��Tq����d�W'Z�<	���(�sH:��� �j`�jL���� ;�[tp-�g��RW�YC��BaK0�x�> ~���ĂA92�#V�$��U�gLr+$L,�W�a{V�vߓ�?+�뤞3`Zq�]_��kHB�L���mzo�x��́"���!�7� [XXXXX�0�,8��	0�o.��T.�9�#��1�p�Ip�)�{jQ�8P�H�*���L�(�ol ��u���	L���"�����d�g���4Am��j�w���g�S��a6Rv�PHR�H,Y��F�_X}5�\�W�>{�8C��"6p{��~O�N�Eݎcݐ��]�x�Zq\y��3����zv�$�RfO�|Bd����$㻉iY~�m�J�5�1F�~����dn�~[XX�Օ��(��>ˊ��-� ���Xɱq�1b	��������B2�J""�cE~*��(bR*Run��T)����F�Z��kM:>:a���I�Z�@����Q-'4l����E�[#�� Jr��\�X�<��6��1�]4;m���i�_����B���/B�%�D�Y�]�bG��N-�d}��/���-.�q��iw��l���)�*rszܠV��׊���:���&¤V�i�,ERֳ%�<��	�����X�:���,�¦�q�u�:�Ѽ&I�'�Mi˰<iǺ-�~�X��W��ol��/�Kz���8�[�7�{���1��?�@���o8��_���̨Xlaaaaa1#/��I�e��H�+�V��󴲲LK�UZP�dii�V���
��6m:>����<�����ϖ"ŧ�T�Xɡ�4���*,V�(Rd�6l�jyFnh�&�\ZF��8��q�Өui�ӴFO�l�c
����oa���}����ha��{9�3��;_=*�ha	
��OyZ^�н{+��2O%NZC�V�Vk��uJj�6�����:��m���Q$�]�%^�;>���s1n<�Y��\?$�syH�_X|At��Q�X�w�.��b}�#)im�+�$HZ*�}׌97ݝ=��MZte�[;�0>��g�������3ʃ����wI4�7����C���ի8�e�`���D�!�A ���#�"���]�O?z@�o��ڒ"(sT�+*��J�	l��Rm&�''���0q@�~��޾�%:�S����8L���4S$��y�đR���FBb��w��(��4c��,�Ib�w��,QRҵP,��1"!��兂ER�-<W�1ENrn��_���}��z�p�6���*�|�@e_o�j�t贆L�uz�{J��������C:�?UD��c�%�p�<+ҧ��)�"y�s������,Y��^��w�����ﳕX6r]�IZj.�|'�m&���s�}J5���<�e���ӂ�,Ͽ�կ�Tj�B�k.\�2n��n��"6�ѣG��g�Q�T�~����ʊ(U.�
l	�������a�u.��D�o�챛���"&k�ӟ>��W�`Yf�[,zTȻ�Ϲl��G	�yE�+�l�J(i}uQ	9�}�^�+�rH��Om?�$�8
]�lYb�K�?"$J�'���W8<��8�}�:��>h~?Ld+ͼ)��3b�c�T�)�[���9z�p��ⳇ�����U�Zɑ��� ���c#s�����Q�����%�ؘ�ťU(���;u�CE���K-��$x�x,KHD�"�B��ViZ���j���"�:#9ǌ+"��X � �(����)y���y�&����)j�k2]yC���3���d���(����~��ܗ(c���_s]r���K��`T �����<�A�	�f��4��n	������Ō@��;\U}�T�.-/U�ɣ-���?��O�hm�L�,qM�;��o���hWi�Eb7G9E���Z������5�����L��S�%)�>:.T'�
�[g��.��шz�Wc�׮�H�+p�(aա�j���_�/>}B?�pK}qɓ�v(�k��a��:��dWuA
j\�Z]�յ���TD�u$�v��R��r�qr,;���-!�6&��O�+�2&�i!�9RR�c�7����Wc�|X	Q�`�R��7��b�,��Kq욫�d.�v~H�$�"�X�� ���"	����?r�������	0�� ���={F��ɖ�O�2�Fp>o�4K�-,,,�0�i�{�܉�5�ۯI�ol�c~������G;��'�������"ݠz�M~�M���,�(�.UO=�Q3b���$Y��\���lw�=j6��kK;7���0�F���F"����Ud��dW ���"<w~���M���{����уe���������pVq���xj�p|_��H4jw٩��C򵞯�r��#&lA�x�n�'�[V�=~=Y��16�H�E��R*�AP@f��V_$�+�j��/��4��j$I��KkZ���f��uɾK�b��� H�w�}G?��#�A����Ĳ`��W����a�y(P@��r.�ò��o,�����c6aX\5�{�|��35I{-�9���D?��1}��{�����S���͠M�Ma��%���(�t���C�n�|ERzy_�.y��L]��Ӈla>>�Q���BvUu��jl�i���
��w�F���:�;Ɨ�L�m�-�Ͼ�����=�i��٣v���ScF�z�)��Km1�v��"Ep;�tZ��r���UZ])җ?��J���o��	��7[�\�b�3��m&j��f��� �pw���X�k ,��e�i�>�>A�Ar@�p��W�_��X,�I�y]�I�qN(u`�L�˺��p���&�L\�1&Ч��w�WQ|ȵ�]��2K�4�(F@��\��IR�:��,�������zJ�&�0����˄Q�m�IBYp)�b9���yE����u���D�R��o�ߛ��v؊w堇}N9�V>��C�]�S7a���T̗9~������K����k@��Ť*g�OcHM;��"������z9Nu�:��|��hkc�~��}�x�*e�:רԨ������ԉ��+�xp����/��(���<�˥*=|��^�|��Q����Z�"�6�R��Q��(�{��䙸�(�d�$:B,/�X�Lʂ���4��O��8p����_'�5	�X5�df�v����;���s�$s���%cQ����މ�Y�J0Ʊl+ߓ�%��41V��ߖ [XXXXX\)�(��3��cnI��	f�e^��h�R�յ��Bɣ�
pCUD�o*�X�@{*�!�[J�h�8O'8�o>�qX�CEP�^�:]��|HKU���J<ݡ�z��s��IT)�L4�;3��Œ�ل$LB����8�)����H[[+���Dˋ괏��Q���J<{�,���u�z5�:QyW�\H����c.T��&g�.�K��Z��>�+�T����n�!��13&�$3�8OR�,�VJ�p�;��q@z�	���>��g&�@pa)�$S���Hc|�8������;��Kb��ܲ�ka�Ji^k�f��t�1ۢ� DA�CI����a�kQ8���Va�i?r���M46S8ͯ�� ��q�m������M��o�ڹo����0	�&����$�S.�����%X�N�(���F����|��9���p�n�񕊸ֺ���P�JX����5���	�W��")y�7��P�~W$(�������
�yB/^(�{��;�l-�z���9BLA$�4�3޳x�s���a�*���"$�o��X*���"�߅9��n�:���\ۜ�9\��j5�T;nQ�4�v����95+syZ^��r�@�_�}¶:6\��4Wqhks�66����{k�o��v�ܕ�X�w(&B�b&ֵ��y��<�	����)�=�o����_����_,� �b��X\`�t�",.���u^��1�c\���x�}4�u���m!�IHb4����B��mƷcA�"�1Π1���C�f� �C��Y�)������$��V�maqa3�Cr��Vdq1���{�?���c�h�P*�@g�E�!E��઼En)��I������� ��F�޾�ӟ�ݥ�ݚ<97�&Z_����tO�iX�9% � +��n��iE����vy���~�8亱ڂ���� 1��I�@��1I�u���;N���%��j�D�n)7��mm�����A�:�,��+�5O-5NN���m�^<;��ݦ"�=�K������&m���Pʫ1D\��B$f��q��|5O�乜�\�P��9���X�+luW��$q� ��N-B6���%�����:ȭi�aY__�Oq�6�}�1�:���G,� <�!E6i\��ں�޹�P�!�,ԓ\g��8�X���Z@Г.�YƵ,���a�Kg��|������_b�eQ�`<w�}Fl����cK6�Ur���]�!�Nc�I��u���"�P��8�%laq�`����Z��B��4�����+8�;*5�/�hii��@�� E�ɘ�\�a���I�����ջSE�O�	�r�[��2U��+穘G�_�%$�Z��啶���{��P�ة:4���wg{K	3���W�X�2�X����ƿMi�������3ﯸnr]ΕU��ڊ		�[�"b
L�wV���{�����F����\F�U�	�O��!��C�۫S���,�jw}�J�*�Jd�(��Ϋ�WrL�+���6G�FȊ��XĢiqҿ�G � �_X_A$@�8��0���i��\ # ���������Rn�o�f`lb_������9p��Z��H�������@ܕq=�>�O�m*�%Y�8��q�ež�/ܻ��=Vf �J����hIo ��������/���������M��=l��94��14f� �Y'L���\o.�^�	��cI�����m�lo$"b�w$���Tԟ��Ď���,�X���L�^���;U�B	�A��1`�a��.��ר:����"��.�c���`��T��Ǐ��W�t��#�0��bHH��mphm}�>��#P d��%�/b-��>��1�%�w������K� �3Ǎs��6�*��[������1�j� 9�B�����<���-j��������iБ"�o�*���J���"�G��K3�R*V9������=�n��Գ�w�a&��U��u�3I0B"
�a.�,��48�<�_����\R�i)Ss�p޻w��``|�ju��ފ��I���;s
��7�1�=�!yύ�Z{�w�"�����7�p�=x��676iggG�QB��(.X�c��>`K0��:�_}��z���pQ%�`�00�X�c<�2	�����Oj��<�F������
�����`sa��P�'{&��r��A����n��fG�_]��^N���w�p�i�%ڜ�(��%�r='JDS�C�.��j��Y��Q�e�6�׸�g����CM��t!ϴ�Bx��T���`Y*�TA�A+���^mn-�bU�f�AAg �OT�U��V��p-t\���l�uCj)RPk����.��ؽI�0�rJF+���`[`Wh(t&u#��H�@`UA���T�>�Y��y7�Y$�ܖA
Ar@D����\�7rǾ(�@bA�9.���:_+�/%��Z�Z�N��&�^�����BRq�v�j������k'Cᶦ�`(��~2]�M�$��I������^�|��� ��`��s���2L����Ƀ�Zk7	�1��0������h�D�$D:y~��ow]p�:�Xsɰ�
�����(v���mơaQ�w_()g��{�j���#E�����o�u(_�S���s���K��R$����l1�0	d��q��&�cd��<��G9��y�=��8q /���y�!;y�ᅰ����I�(��Dq�� C�-'*��z"�r>�������Ȼ⪛̧c���{?+�����25H�X~A~777����t5���r-���Qg�	��qr%cߋ�T	o`�n��&d�*p��a����w������=zD���g��H������^�xA����I��=���4N��!�$1S0@��~��K�w��%��vۈQ�6B4H n�d���d7Y�baaaqܦ�w��r_ͺ��xԱB'"N?)�Ry�tTJ��-p|o��{:�Xm[ȫ��t� .y�
�SD���(��G�߼WBnKq̱�y��/�ԩXB}NE��3q\�Y�C��9΅i��jϸ�K8�$0=Q�+�ׯU���!�����7���95~�2Q�iY�	0\���Z[V�1�b7�"�*���j}�Z�J��5���l�����o��Xծ�Q�����=4I?�� i/�E�5%���f�5�=A��X\��ŻD,�8�X�/�$Yk �s�oi��|�.	�.:~�H%�׸��Sk��;����p���]�q��&NZ���������G�8���9l�N\�mB��$˜dyX�)��2,�0@;!����"܂����,,,,,,F#�;��ƾʘ0�y�	��J�@V�Օ*�O�tz�$n�=��cK����Y���e�S$��!ы�r9(q�S�qJ�?ۣ_�������&?�r��;�����Gmnm�Ww�b8q�.@R��ߌ�'凫�W�����۷oY�����%�"ŀQ�W�~�woU��O���:�-T�[��<��7��V�55���j"Cn��J��Ksml,("��Hr�ݝ��-q��*j|����Pܤ�ú��N	�'-�ȫ����@J�H6hȽ X��$4�t��:n��j��[|�b�Y�)1�BXL��eXb���z �K�*��ݻwl���ގ�b�{ܬ6�m�/H�%�bt��s�����+���?�!�@�7oZ���q �%�=��6�����[V�]N{�g���p�;����f�/�G&��@`�M��m��K�q��Ջ������$�c���oh�u;M����2��v�����
������w�	ޥ��zƢ��4�^kRo>ON��V��a+\����b�����n�h��q�^�X�������"�sT(���
f@�����o9�؜қ������o���4��F{����!5�y�851gax�����"�����*!��?}��=ףb����*!�I��񱜣��Oy5��B�-^p�^^�Pk��ĵ\*R�𵔋m�q��V��j��5*e��������F�N�m�	CDW���ȁV����$i��dr,dhȹI�`"�kG�5c4�lJ]^��Y�8�eX~�ז�Y'��b	�uR'8��%ϑ$��D�%��G�9I����Y��,w%�	�
�q!���ًq������S�?iD�l�8�fN6ά%�h��]B�4��������7>�R
7G4Q�y �8�b!���*mln�f�������z��v�v���8��Ȱ�q̌vL7�b��6?�׉�Wi�]���A�h'�%Z�}���i���"2�\^#��S�U���%�̻�G}_%�V�Z;�2���� W�eZ^*���Ժ.�x��{*_�b�Ljs:>m��Q��h�~.
B�<´�U�8��x.�\��V	+b	�K�Th�N#-�.1��:��,��9���NP�#El%W����Rcc��\ZQ�H�<n��'��,���
5��xv��A.�"�r�܊PwC�c�I��^PPcʥZJ�� �Z����N��b4D�Ƴ�K(�!dc��0�@�q ��f����"�˼$��ߐ��)	���Z���fV��I�#�o�Z��A�Ԕ=U��q@Z�p�R'X�M~�*�q=�,��u6mO�Z�s5��9Ic��Vf�_�̱4��w��E#.������'��wx����1˚��7j&� - �VT<\|fAmh$���S�$���^\��.� ��_�ܨ�;\.�#�C⏲�}���8��F{���j�8��y_ҳ2���a'��B��.��ىNɿxWs��]�X)ғ{�2?��+0yI��HHp��P��s^&=^���J9���:˴A�+(R���޼=���t��Ȓ���9`�.s�V�	⦅dV��&��!-Lj��z��"l�A��
\�?�і�0j��������3��I�/�����R1���B�����c���ڑ����1�ƕ�����h*b��X���\Ǔ[B�q�V�!aI��\X�`�Y8��ɌN�[s<��@Ɩ:����ʌO3�3͚z��k¬�"�����VX��$��z&���{��"S�)oS��X9C��gD��$-�I�հ���ыj:����@����K�n_�5�l��<�� '�/2qQ �O�<�Se���'��� ��j~LԒ�J�:K��E��EK�1 �bZ� ��޾��}��!��9^�~Iϟ?�g�~P/��h�֢�K���[XXXXX�')�D��N�d7�%���yɡ��}|�6�(��K��kr�+$��r� T.�dHO�.gwF�_.���|����:D{u���oԼ�ڞ'$�Z��q�q����!Iܳ�t/]q�b�Jh_@]D�*�����z�
��E����J����P�Q��%O�ٜ��E�C�����!�m=?T7��Y^�D�7������w~E���R�XgX�1��y���i�Y��� �
Y���+�$��2�)��2�n�� � � "���*cܥ��&!��.�Qg�A��&��X��^�#%9��g�Ϳ�8������}�H�%۲-[�,Ŏ����f�!p��I�c'�ĉ�ؒ-k#)����}f����q��=0 f���p���U��U��+B�/�c�&t����>*Te%�+����[�������m��?�����jרt  �j���B��e�=������DfB~�h��\�ef<�&�7���0�����FN�<i�^4s�P��p!N����g�1�9f:'O�
�Ã�e�we�6�L@���a���
��PCGYhЃ�����Z�#�ǖ��}���p��;��;.^8�ϟ"�F����Y��V���h�H��*R#Ͷ̌�����l�}o1|�����wí[w⽺�5]�%�`x�^N��� m�ג�R_U=C\|`�����<h�:����f�s��ͯ���N�����u2��0��oul^��|F��JC��D����d��E�5:�o͇{�V��qn���V��	�q.'9��<����4��nġ�8� �Uuy���H��~� @E{��a����ߐ$)X�"B�R�_]�%~��׀CG���Jp��oj0�oU��؎C�͜�t�=�	sܧ��}��O<�A����|�IK�~�@��� �ҧ�P�l�`%�>���Uh{[��t��%���]��������R�v��K�.��/^�/_OǶ}�����hI�777�f�	�L�������PCqʴ�4���Q���*f�춳<�Q���"S�	7o/�?�wݴ�?�����K�Ck.2�հ�Y�=���ʍKMc7c�� ���E@ȅ��։�tg9�����,|��RX|@T�Pj�s#Y����	�A��*S�*�B���t�|��00C���\괻a)ί�̇�o�����{�é�($�E`�/_��(��bs,Gǹ���:��?�T��;�^W�|�اᛯ���[���7���T��̠e�0 �=��3�� L�[ZOo1��7|6�7��F,<>K�S��\|� ��*�b�I{� w�0}Sz��'ԛ�>��o4�(��gY�j��9�t6P�9�wѳ�P&ؤ��=� 2P����_̞ya����љoۑ>�_u��,l3n9�Բ,_��l@�H$��g�?u�����{p�7m0!��/c��ݽ�������_�F�PC��*��aiz������aֶb� �M��i�K���,.ŉ��-Uͅs����)�E��@�ެ��{�X��Ό��v�N��YX�Lo�w��"\�䛰x%ln��}�S��vK�N8� ��0�e��v(���p�ݲ�Gh�-�tw�Kq~}z�f��sfnv!l�_
��]'����x.d3��8wL�lP�&�d.γ����Z
�?�>��p��7��"��sKD����a�K
�����>�������	�oi~��{��"����J[�>��?[��ﬀ,8@��c�[�S%x> ���/VC�<ȾKQ����W��h��1arp�N��7ߴ��	H�~�3������U�#	nn�{�ws��"H��"f:����{cc+<�,���f\��[{^~����'�k��jR����6ܿww��٫|�-b��A-v���dn�rC�R�.�a�B&�>�p��v���X� �]$���"����_O=y6���3�m�~5~Z�_�E4ޭ��G�0~6vb��GW>]�:|tW#��,bt�������kއ!W�I�x��c���)��,�7���֦=K%�g�g#�R_~y'��l���/=~�ʷ��^�@(ί��7g��C��n�_�I���`=�q��'���D0��8�n/���u�?�	��-ea�ߣ���	6k�`Q"��l�7�MeE�<`Ds
���|iG���0��c�/��>�% �WF�+0�GFP%>
����w�*�� Y�.S���ԛ�ˇ]�����
,��ms,^�B;k�"�kѝ�h&�HY���7�'l��歛q!����۬@:H[f�l�<��iJf Ya�D�[���|�B(�&qׄ�����o��Շ��͛� ��<��ַ���S�^�w½�wM��94m�&fѓ�9z�qƛ��� ���H�Xc�`��$*[5�� m�u@U���ԙ��;?Ȝ�����:��oc��A�nh��e�AP?����2�T����<]v�΃�a�>�]�uݭkJV�>c��i�r�E^�$ ��f���%��q�̄��#�w
M�l8v|����LCf�fum+,?\7����_�
W�~>��V���aq)2�E���e��~���v�/�\����_s�g�z��G��V \���=��s���(�jNvh��@W�&���sp�K��Z�6��φ��ZZވ@�L8s�X�[���\0~.3��mJ����~W"�>��v��ӯ�ܺ�-��c=lls+�7=�l[�t����d�}�-�)�s~L|�O��k!|6�� ����oV�#���k?����T>�u�>��R�Nc h���] ���. .�v1}�����]����S�;����v��x�q�����*W��|?�|���˥�r�Mc���Z��\�@d�̣z=�x�RJ�����g���,���f����^E�87˄nY�^�:�i�0sn�Oa������Ʀ�E[gnbV�L��SL���ݻ�B�z-���xy.Y8��-�;o���ջ����N���L��A�h�W�<�[�슠�r��M��B�f)!���������U/D��J�|��T2�ϧ�"m�����SO�=À��6#zT��7R4��`kG��Uh�fa/>N�lp�AUfj����(�9R}\�T�5�`)*-�����6`����㏝O\:�p&��p:�<q<�n�E������_
�n�_}}'ܻA��e[��ڙ��.fCVX[Y,A�\���
��U�1l�΋�����l�2�d��y���1ﴏ�@1�s���L������ u)Ι_|D@������8�;.<N@�q~aR�5kue-�[��+���oE�`р��j��o�5�-ow%\�	$��f��7�/|�3����o���\�l���sJ	
o��K/��?��Oe:#i�8�`Ww�Љ�f� @��z�	T�t8(�Z�zO�t�	�E)ȼ1c���1����mJ.��x���zg[����P� ��q�]ū���W����5����0/ Ί��OX�N�ꙧ��/��~�i�p��y���O�~��7f�\2_
 ��M�%�Y8�����s̃c�ܽ��s�`�ba��i�����}�7�G�xkc}���nw��̄��s�ҩ�֖�/����p��-����Vv]��CT��M~"
 |������^t��h��ۃC���2,$W�^5�^���'��9�OО[�;��Ӥ��Jy%	gzO�K��B/)��~rήۓ`�����S}���KDU�d�I���?�~/uC�!/��������ԯͣ����Ԟ��0���h�9꧁�v��雛��Q����m���k��nG��T�������3��Ӗ�`.�H���m5(��=���x� "Y��`D����JOW��,��}9T�u;�6��n>U	,��~�� �����$ �/J��U^\<�PFa.�Ұ�-�!�X]��եp�n	wN�on/����s�φ�'O���WW#�X6��͛q~�[ҝ����B��w����j�F�'��9*n@��B0,̠����W�Ay�Ѡ��B�P�g�G�>�E���p ��8���}�׃���71�P���+�_U���W�6��q���@c��0����;�D��Jp9��� �&����$,R)�`�A>'�K1��������/��",.=�/f�r��K�s߆�]�@Ul�D� ˼�o�yf 8�H݈�w-� ERp���(N��7-�9���9�|_��6��ǟ|b/��(�x\�|�ڋt����6!,�^)�C�$��o��f��믛F^9�<��d��c��
Hخ\�R�<k^�
��	<'f���9�T�EJ��=%��T�6�}�`�8�~2�Z�;ux���S!��cn��瓦^6�J��FBy�=IS�_m�� A`^�h@������b:�Z_Ou*���8�U5�x9�T�<�֏y�24B�&bs���n��a`���{�m���,��ҶeJ�oD��~�US�;�Z�h
�g��.2b�/�L	�\j/�E`/��������:�� ��<�T�0�����U��\�ϫG�GϏԪ����j���N�i��[(���V؊{"s̔��[ox����X v���������z�g�r�i�����[��=7)��Q�C?�v�_J�TP�h~q�d��(z{�σ`�*��T�`�3��$�:</>j��X�@c� g��7�(s�s�ԉ����6� `W>�(|���᫯��<��b�,;��63��df�l+!���N� x�������|�(i[��M��[�6�WVV-���&".-/��+k�<(VfZk�w �7��2��z�����K�L��g7L����oF��[�J����Dl��/�X���{@�"�7c����&�ȞM�L\ӐGpKY���'s@����S6iQ-�Wl��Q �X
Pοt�C�0܁9��,����:$~��?�>�D�Ky�ܴ�z�xp��|����Q���F�c�h \��ohHsD �g'�>C�ڮ���?�h�<�@�wH��Q��e]2M���3TMQ��ud�c��-�Y���xd�vx��N�i���]��-�+d.�5��3oqQG�}��ѮWQ?06l�άq@w���Az�0�|���w�M�4�)����N���v[����ʅÞ)���^ssEBC�Gz��sȲ���5�7�v,�>������QH���p��N��������0F��ڝv8
��n��b*��U블��#W�qh�@j܏g�F^Ѹu_/��pGy~c� ���R����h`�d�����k�ڵ�|.[ٙ"�\ml��R�f^��1����bN��o�`�r��*��T�)�(effrS��t�J'\�x��un߾nߺ���M|!r��.0��Ͳ��V4�Hӟy����<�ͅp6����C�0[p�ܮlb_ ��" x��J��c��� RQ�5�50��Nc!�����ήa����o�9~kRS�/�0p�DNZ^�5���P?��a�0E,Z�����ߜ7K�X?�����O-���}S���k�Y{x!�˃���n������:8���1�fE7bY����|�S>�W�����M�v�G"R��CU�4���I_��w=�)���on��Ih������&�N��c�������O�oC�k���h�)�M�spa��ҵB����:͞��[l��J���m��xغ�O�� ����q;�$�Pp/�7\�؟>��S�?[��H3o���9�����0>���%Y��;$X-�l��
a'{�x�����cG�~}�v��c� ��������˗V���=�3��;L�����p�	4{��.���s��Ħ�}��Q�����ݤ|�kP�>�����������icn3r3NB�c6l����'�� 4�"�w���8��"sv2;]2������ڝNaz]��z&�Y���ge�`@-u�O̢ݎ�����F�6	�댜vk��ob;NG��N�EM���<�8��3v����D�K�v��Ab��9TN��*?�9ƳZ��^~	���}�w�z`0$E�D�x����_�gO=r�)�,  �s��x��a�x���B\�K�<���7�e ; �K]������m@E�}�~�����N�
6!����gl�S��?-��i'Ϝ�x�<'��-��@��9,/Id����7/���.p-���G����O�d́�iT�a���֝ӷ���꯺J��`�c-C�"�&sQ�	���z�

�ۭ;�t��� a=�ӬW 1��c�����K�J �2�ψ6j� %H���d�W��＄��2�,��Uħ(:tZ�4RU@ZxW�Ci~�?���^�p�|��W���a�jG��s𬠹�Y���4�T?+<`�a�~9O�l\�!䀪���1�.H/@��x��'��[�M�he
�L��y���4\�� � /�^����lnfS �`�Yf�x��/g��f8n���*3��fz~nޮ9�p,������Ր�5�L�e��
�ߛ$׾>�q=����3Ϛ���E�-�H��?�J��� X���䅏JȒf��2i���0H�p�a���{�g���m �/��X��C��\a�N,ܴU��f�^��p )/=�x�(K{�����o�mL��˗�-��Ch;/RC�Q�+��ғ\]>3��Ht��zE��X��#�sH��h�F�y7���F}���a�pz�xGٸdꤼ��0A��1<����(h_�;�z
tE�W*��9��:>�s�+���k�����Z�Z[��y�$�����HמR����s��`����:%�@��>����}i/�o���:.y(i� �Q'��� �V�+�37X���+5��l��q���\�ۮ�κ_��V����n~g��P��~����C��&�[��7��t�P�� �Ax�ŧk�z��q��X��N�?�`f�>�d8~�x�����0�
?�e��%��S��sy�'���[�h��!ڧ�4���4<GFmn��ooT��yV+���jmkO�]�Ў��W��IE �N0� ^^~A��f�~-�td)�Gr�=}ټ�(��ؓ/Q*��z�#�N&�&�E�^��@P�Lm4�"�q��k6T$vj38/ĺi��\+8�|=������Jgڤd�2����d�@}��|�r�M"uh<d����i���
���?����475���y6X L�85_����,xEZe��0-�s�u�û�toiZ�i�a��M��ܕu��n4U_iO6Xk۝�jj|�~&ƻ���5���~!	�������xv�?����?4t T�i��}6YBqL��	�I|���f�Ӗ�Y�T��k�����#�`�g���J*����Q���Wh.��A�r)]$cN�/s�D1�Y�y�!M0�:���>0^�í��F�1k��Ν���`Kh~���,�_E ��%y�A�f�E |.~Κf@�'�[�G�6��"B�̭fH�4Wh�
 I����8��Q��S��c��>�ԁ����R| [��-��_g3saye5\�q��	3��\����b���>A@&���ib���:n���z;5� ���;Tņ��?�X1��G��~`��,F�C(�K#Se$��##�c\�	6�aQ�)�fZ��^=m�JU�L��1i���* L�d.$�k懂gq^J�@�L(�6�����O]����Ґ���M1�֏����:R��(`zRH5Y���^�})5���Y��s��K�AY�@�H��9����� �~�n�W+�{�ظ��k?��|N�����w�j�y���%K5bx4��B��QPQ����*?pOi[��DJ���<�q���7��>B��e����GG}	�J�4�7U��	A�z��+!�^*�=��@��\/J)��(��}{3 �o  s��%^�{q22![ɀ��p�ef�H�,�LЭ"�U�[�Vj��ϔ�V9(s�ϳ����������\s��B{����0��l���a�c����-�<��gN���Ç�a��xlib'ny-�_���Nw�ie)e+�=L���u[T1�(���6N�ۖ��(�H#�� G 0�RGnMp���>��t����r�OQ�4�-��J[+4�� *%u(0��G��	�4���@m�]��H�b���nۆF��)�M�(�^�j5� XmN%��"`��3*���q�6�uRLB�����1���9_`GCCC�Ǫ"�/$P"�gx |C���~�W?Sw�ai�{���[�g§�o����*�*��n�\G�(����#V�XL��q�W���H�YQ���s+}��<�*hX+��G�����!<��c�����r��$���<~�I�*c��v8ؠ)�sKf�YV���f��G�*�eE���ϵ�Pk&7�6�!>������{�y5�ݭ��<�fƴ�D9\]yA�M��⥋��o�'�Ҥ���zmI��\_n��u��K�B���?ڷ4��/_�2H�X���b��v�k�Xl��ř�Ma��y�-i�� \H���	@S�R�r�ׅZnA�r�u���y��H�8/9�Ѵ���u�.�����8l(��vG{5��F�k_���y7�5�o�Y��Y��4�Б�AJ��C|�Dk�xT�G	�4C�+�n�Yo���5=o�q|}0�-��O���OYG�O�B�J@;jF�à�{(�\��/�SY��� m:o� �W��6��K��Ҷ�y!�˄��w��g�@6�j,�Q|�H[��(�&<������0.A�>�K������c��V��L{W���Uڛ�je�uu-�_K��K �	/a�q���Mo�&��� Шh˘C���[)��HR^Q���k�<a�Sc�(0�����q_ +�����Hϖ�M˱���`+77k����	#�PdA>��V��A�4��ӴHP'���j���U����<�+Ja��o$>J)i|����zh/�H)U"�TQ�/����R�(�
� ���cT��]�!�8�:����4�S�@p�z#�g��B���j��'��_ק׌Jc�2C���d���ɋ$ `��Ec&���L��DD���Uٶ�A	�J�OܪUh|�- �(���bȊz<�e���i�	��py� �R �� �`[���A���E�����Y{��7 xsC��&�<0էg����	�����M'�'�P��?W�j��V����d���M���`9�v���_�vb�B]��gnm��Nԭh� X}+b��!h~+�5�����p����b&��g���iX� �n��r�WG�
�_#-�H��eP�PC�4��7�PC�K�T�"�;��Z((��- I>�����U`j?j��4Z���?		�*�$��w4xFx7�鳟4�{���8��tW�i�Z���o� 8D���ʏ2��$|u~�H������@�TG�+�B�V� �=����'������!$���i0�Bl�\l����"�}nݾ���l��HS���F,�;eS�I�
��e5M�K&	����N������^
���G,8�O> T�1�8E��"%Z>),��q���N����=�_��*����jC��s��"�T���k)��5A�8����0:e�i/�)6��4��Mk���	��l&�GK㬍�Y�j��G����5�wjƷ�aH<��^�T|�u����G�[��Ah�:S�T3�R��%K�K� ��%��(Ç�����~��6OyC�i��K�T��돋v�v��hFN�r�N<d��YK�±�'�����S���<�0]o9�c9il�@�*�I�k�	�}Z�
�U>����0��'��~,��I��.���t� O8z+�]�)|���n:�`*u�<�T��5�&�(�4�Kbi�T�!'���)��,L���/�8 �ܟ ,� K�/=~s?]|T� �]:/3cF�D=,~�=�̇{��{qO�}���,s�k1�� ����x��fB�`��eQ�e�����&$��E4<�N����鴑��PCG��i�i��g�>�HR�����@�Fs��^�^���k�P�z����;5e�Fni��盹{<��i+W��L�!�9�Bڍ�M�z��v�lx���*�����Ώ���`|i��H�m�]7,�.�1�	�;��=}�ES6�S(�S2�����u�W�i~�<�Qi���F�n�g�	7��ӧb�N��zcm%��l(r�����X )5ͅ�/G oѣ��Yy�Ю~��e�+�\���L�Yx �\�oI�D2mFbH@-XҌr/́aPu��݌u�B�����4��R酤�[D�ib���y}��"*~�KE�&�V��BȦ��l��,�Ь��j�I��$�W@6��c�K~4͂�PC�C�����R�2�xzf���M�����O��\τV�e�z� t�l�����ǰם����ޔ�Oۗ���.mKU`��R ����m�&��1'�O	'������hh��9�3�(=�,��G�^�/J	�# ��?� ����wXaf�>���(�-���g�4"/�0�P�,^0k?\���6�7x�:�̑}�:+��YSzi� � m�+@Z �^�\�R���{��9{�ڀ̍���կ�*����7�,�W���"t7/g�f���i��l�<�����؇m l1�⢁��M�,�����ؗ�&��.���~�@��XRFA~�LdXL � ?@'��_��	�HG��
T� o4�\C}���Ĕ���E ,��_}���S^9z�.��q�
��*J�A��Q������k̂/_�6Y�ʴp.M8e8���W�W�#Ə1����j=���1��3�nJ���I{eR0��{�*Tl$��H�Ӳ�VE�AJ-"_��"���SR���Ҽ�>莮���:o��BR���:�yҴ��lç� ��ڢ�h\��M���(�ڧE>��_��U5�{׎����X� �)4������pi�0fa����Z%P������l��������AJ9.bRzJ��y�:��o�G�3��][7����r�\�N�e��s��y�'J ._ߪ�&O�z���$Q���� _�ߞsP���5��<�?V�nmmf�.BZȣ+(�$9�&�E�e�h,�T�-�mwܒ�� �_$˳�Za�.�1@���fy�-8Ҽ�)����h�0}���E~�*��Z7���dA �]�r�6��%�8��h#�ٯ�xu��O)X���M@� 0�Q�dKmԔU�d�C���K:���[H}���9(?a��.�����k)�sֵ�����
`3?�H��
8��LY�jkl�85t�T�-Ɠ*��ꤱ��7M�O�
� �4Rպ�:��UH�`¼�J (��)�JϧD\)�����*_�ܪ��u���U�_��ٗ�u��Օ��[�ח��������vO{!{�S�<e>�ۑY�ź�eª��T�G�ƹVd�wˁ��=yT%p�|�}N�e�GYE ���(�3x+}Lc[d�tAU��ҏ3�̃t�[��������h{�V�b�����.�i����n��Q��� ϴf4*ɶ��;�C�0� _)ŦRh�������v�-v���\���C���U��<Zu�\n�1��zq����O��I����!=h櫊I�X�8&mA�Ű
@o�h����6Y12��$_Y�=W��o<�&�flSNRHI��z�e����P2�ԧr��͢ꙙ�ĐO������i�t��Bu �(P�0&��_,���{K	a^���??����L���+��^S����M�B�O����T���ԁfπ���%a�0����k`����0U�[_��H��1�#ͻ����&	;�����ߞ;{�7��7n\������{����E��a ���߶qW��Qm��#�7�sbޙb������{�����)�%se)����܎�!�X
�8oeR����"5�]��tN։�����7t�4I��x�@��X_�@H���P)�m��Y��mS��7K̘��^�����7)T��Q�����t�e����5���Fn~;g���lR�O6-|U�㞪$�P� ��*��@�4����$�b��&��PB��O��9�ۓJ,�-&̛2�
�ƺ��AUڟ�JuڴA4M ���Sh����o}�[�K�赱��0���|��'��Q�W�
Oc��g��W�G/,p��Q�R!`���2�D�Ʒ����R�;�)�^�����u�W]���
�륽E����؀,���>� ��=K �F�> ���c�DXH���7�(s�*fGC�.��殄S��b�0���V%�6�fJ]!$���<�	5�4`X Xy|�R�P�A2yN߷�*)��� �$���IeZ��K��^�g�V��A�x����}h��� ;���e_,$V7��o�&h�(]�����*-�(���OSڦ:� � ��}�yi������e�(�����&M��P=2�J��Q�D�	��Ѵ�A����G�L�#�z���w��E���s�~�� ��s !R������]��m�zMo���m�g"lY 
�t�y�_	-}�*�&�L��<m�/��=��_T���u�u��W�ӷ] 7=��y���?���K/�d�����`��h������ݕy<< ��W^�߸1d�УM�H¬T0�L�-�N������ʲ��p��B�
Tڣ���I�]��wI��GeW+ &��F1�MKr��3) �ےN3�f����vU6����[�Wk��{��# �������v� Z, s�3�@��M1q�1a���R	���15�*�{�0�UR��>��0}�w΃c�SkAUTg�H�$Ȑ	u?��^��<��d�'�9*TB��4H�c�i����P̿�G�xN�@A��Z���� .k?�� M�'� � �d�3F�e�SNPiu�U���W��(U�4�bj����[��(�
d�^c9�O˺G����s�:唗����)��>�O*P�[A�I��<ɥ�������EP�V��#m�4fҎ)�<�L���o���@j���/�k\��s��R(���9�u��[�J�{T)�;K���z:g�{���,��A�5O��[U�b������^u�L'����Ѵ��i�OG+�����"�D{EPl	 f���`�Zy���fP#����v.e��6V��d�������az���~�Z��7�|s��xX�Y���c'i]J��G�BҌ��(}��g<�ߘ|��B׫�t��me�Q>��R��&�v��z-����H�߆�(��N
i��{<�ͻ�B�al�"v�4��|���G��ʻVe��R�8�����µk�l�� �h���o���&�h�^/�
PBS8R�%�C�~�iva|�O ݔe?d�k��=�kI�'�c�l���k�g��!��J#D��?� �! m������&�����?`O����ąF�����9D]�����}���P?�S�稏���16�ør/��O�ύ6q�~��V�k�~���N{%R�>(�^�$~���λ��K=����<�<��'U�^Teu�Z��ǫL�Ӳ����[�L�Տ_����X0�j�0S8�����
@Z��Z��v���:/�-|X��<�P7h��⭏Rk�ˊsEE&Yk���K�[L7��D�-r�f���[�5`�3���l�jm�� �݃���%]X �dax`Ҁ#���N��������()z*ٓD�c���/o��Ny�1oIs��Ϩ�ޔF��o0��6𷀷�.�~!R��S����M���:?��ق|P�t��ϯ�ݑK�3E�].֥~���x�1)e��̴�������M���*PѴ�vUL��� ��~h�V�����/�˗/ ������φ�^{;�+] ���L�������[��=X߸/� t\��:@9 Xk6Srx��?��e�K=�<?�]��Z��r&߀Ni2!�X���. ;��k��R��^��w<�KY�i7�E��Ƴ�HX �/2��G_W�[�u�!�`������f�ٓ9O��E�s$`���Q�O/#�q���������12a��\y���h� -˦S{T���Pux�x~�������ޣ���`��^ŉ�� O���js��lU]����c[є�_���P������u��QU~��v�4vh66��935:7�cq� 7�]��-�]���Ι�±�PP=r�$R�V\����Zc]��vB�L#��_���/���"Uӎv{��mfV̢�n�s�,_�o&�u��o|S�r���6��b|������eP�1����"�����񀑠<~c�^��h�Ny��(���_�U��0���E|�aW�a>�d+�7�F���Q����
��q�)���c�p�\K91�O�yj�_�_��ʉ9�@xR�i�t���W��, �Gq�G�L�e�2SF��+틟�{�VPk�\�9 �A&��X� [h^�������{c���'� �%�-��W�*��� ?������G[� ��5h��D��׿����> 8~���k�*�,�c�|>^φ��~sb=�5�V�O L9�?�o���Ԙ��M�(�,7ډ��O���!�/~��ꫯ�P/s�y�:P�ޅ�Yi�h3�po�g�!�ô�g?��=o�/�����8ךA�{)�������2���~�(�Cs\Yt^�uHkL{����J�}~���>hN���~�㣙�Ϫ��'�e������Ve�������*o���a��7U�n���My�\�s���(_�xp��kN�H�� �S�"�X.�͵հ��δ�X���l�˞�$i��3c���C]:ۖz�\��h����)&bȵ����l٧��ogÒp���ڷ�� \0�mr{�1\KK�;�y�4�����C���x� ^2�jYP�c�1��_O�'>00 ����ƍƁ����Iyy�a�؄�^6x��V��<6���J��Ǻ�7������C�}` b�o�6sF�v+��B��p�&�P�W�y�J���K�0�S?6��?
�ARj1�Whmdnx� Ш4�x�2�BZ�.��B 㨽gU߶%�v�?��� [��/���qY� �)�xr���J���i88K@m,��`�����D��k�ӝ������ �h�\�� ��}h�b]��h�8�i�`y@5�2.;Ʋ�S7mdWNz冧4��K&��Ͻ� Ŝ��6��?2sfݑ�T�B�1�8'�e���̶�0>�5���3��Y*͌�	`嫭5�P�V�c�OcT�4�=I�����z@�-��2~����{P�a�My%RU�������~<�~Zߴ\���(k��l�60[�(��-���h��V�y��>��q�}��y�R�-�%�f���t;}I��ߘ?g�-5���&Z�M���B+ݱf�Y
 �>��>�  >c�"�,��[ے�����/6�l �l�J P��ϛ�
 C<K�K�=c��0�A�5H����?����l�0
�B6}�E�� ,J�C��_����H��C�x�Y�?������uQ7�z��@�i/{�q����p���p����&�Q��3f�{�Ǝka��#�&~�w��(�	�t�0����u�#��A^��o�O��m��נx ����-����>0.`Dy�OhhD�W�(��)Q�Y��+��*  ���5�2���x�R@){�)ZQ̧y7)�f��r@&�&���z+��o�c|�������'?)ͼ9�� (�Ⱥ��[o��8�Z��:�)2�Ѿ�������}���k �� Z���_� ��~���,���oƓ�$lFH��Ii��SEו���%�����0�Q�̟��jP���>�Ni��Q�T�W5�0����C�X�0��8�iKL��sk�_�w].<s�I�꜄������N���,������POz�[��fcج���	l�JtM�j&OD�����͇�����5_��x?��� "R��*�zZ�ͺ�=\y��V��7�M��1nD3-3^[ˣ-�ϛ�m�����h��;n"��*|Bs���FM%��K����U�Λ@{0�M�|�L$ۀD�C6b��Ɓ{0������(���
���a���g�\Q �������0�<������/��	������}/^�T��1)��Xri('_3EѤ�*�~����'��*s���C~,e��;�R�QhT�a�L"�u�	����(�ӘxR+A�Y�X�|yEǇ�~��Ǭ� Y@1k��yZ����u�}�zX� 6e���=�?���oXåe����������`�����`�� �5 _��j3}���q�^?�D��q��z��T����ԬH(��$k"��a�j����2Ș�D�.��w�dɪJ��< I^�d�9j���]���J{ף�Kx0Y#�\Se£�/�{��wR��=��+���_�K�<8X�5��<�I�wNY6<�uڹFu{"����*E�a3����,�	��_�#�le�Z���57�vHV�E+�>3��Ԁ6��j��e W�~;*b�\T���y�Rn&���bo��l�(��6�>u�4� �Z�ٰ��Ih0NJ�ܪ^&���Gy��ݛ9�eS&R� B���1L�U�t�-�3���Q@Z�������s�р��9�&�50JbrDԭ�bP�G�9�6�4�WL|�d1���|2�F
CDY�,��DY1p��>�5�ϙ��5{��H�"����!����P����SAe�fT�u�����J�O;�>d�Aĺ�&���� q�۬o�N� ��c����6��>e͕_�w�Q;��P������~+���oh#�0Zk̪Y{�����G���������f `ˇ5������RNѕ�"��@k|�4��~��P������|Iq����5�_8ƽ� �b���ʋ�tO�-W#	�鏴�Ǌ,^���t�B�f?���/<�����4M��%�'z�Y�����R�A�g���u�T�@��@�`R��b^����@�r،�������� w��0�婓��Pَf��\�)Z�)�l�;gA�R��rm�]ȶ}�)\F|."@Az���r�%4�->��F��֔�*���Xd
l�E�pŴǶyLU�Q����K�،e>��ތ��"�1.a28��ʩ���4 21��,Q�L~�����2���n,>b�ĸ�� ̢D;�ʟ�r0)lZ��qF	�φƵ�_i���L��s&6L���<R%�h�ѩ
�YB44<M�\|�,+��ѳ>f�.���>�6�^!,D8���Eެ/��H��K��U{�אx��L�u�4�])�um�c���+����̶ۛe0(�v��g�6ˮ̗@�ۛfQmP0*�'Վ{�k���̲w�E�yH�˷�i_� ��Of̲�JcO(@��&����@P��R����ν�@u~�����F�יs�8<We�@q#޸��#	\S-�U���Jϱ�$��V{,�n���[8�k�0�F�z���P(b]ķnX���onZ8�sg�[�,@�i���L�縧X��,�hu;�	�p�e��L!�4�]����nn�lm��F	�9�|g��_�mZ+�2���ie4�'N��<�IƗ��|l66�m�'�v�d%��eB�Y!�Rj�Hfl΀D6nv�i)�&�H���{��U;Ɔ .�a��4�{�a.�T�S�F��ސ�[ѣeJ�q>Y�� (lF��2������V�M�wiP$���)'&cB���D^e��?Xc�1OS(5 xw�k���Q��h��i��I�Q}�<	�ؓ_|�%[�X��b�AC (�Y�\Y������G������;��o=\�4W�4��6���i�d��u��Y$`G�)����˿�0Rf��	0��-2k�O����W(�L��a��̨%��}�c������|lK`�F�{��"x*
5��ߗ}Bu�|s4��/�y�E�.��y~�|��J�K�.�q��Y�A/9Oy�joU��q̻i���6��_'- �AB(	9�_pC�Gz�f֎�����ٲ����y_eA�Ӑ��� �~/�0�C'�K��_؂�؅� �9@+M�U���ӰP��?��R8;;��&q]Y]����ƅ�1�L�V�*)q!o!���M�# nfI,W�r�����kŴ�wm� ���r�eI��av�S�!_�x)�8~2|��Ǧ����v��ת�Ir�J�Δ�Yux�~I�e>��.�\�}���͘�^�EB���R�(Ӓ�f���F�p�-s"��0)�����X�\�ƴ��Rɼ��0=ژc����U�c�ʷC�m�n�%7����e&�0(�4����oL�mNz���;h���}a�>�����"pS͚źL0�'�:IY�#V0�K�a~a��.�@��N*-��+�Ts�����z`���4����0�Ei��˗�{,�����b����k��0�+R4�`]V�ż�Z����0m�M����$P���;/Ǆ�ᩴ�2���^%W������� ��8�RH�U�X�@Y|4��R�G.H���\�S9}*�Sdiŷ�k�Fi���u�WyA��S��}��N�Z1����t{m$��߲r`��@�a�� �f�J+�:s�A��I�O�������[�|�c]@�B
8��,%�*���G���a^�Af0��2[��^�j���~�3�`>7�;q��_vȺ��Aj���3i���09s:|����R	f���|n���M�M�?s3L�-3�6s�rc^0�qn��@�&B��K�A�����?(c�l幊-�w���Bd .<.>~1�?��u~�ŗ���?+��N2���K��#��ԬJ���|m���m[БXr��bL�V���4`Z�qi�����4K
�1� ꆁ�m�	s�h����M]0������Ac���)m��vlV0�֋h��F�h2��^�PKC�B9���,���{>�b�7J%��?�g�9)4̻��+e�X�X��s�z����Ȼy ��(-?\��Εn#I��\�ND|�e����R���',@��� ���b=pk11#X�z�u��@)�=9����eγ� ����Us��#���U����B�a �4�/^~�4▎��gm_@;N����E������ DP1����\�ܽS樗���?��]#`χ�|��f/3k�8��5�'���V��=FY.�����S���S��cau!������*�;I�~t�p�{0����L,�B�>k��\�̄3Y�g|w�i)B>�%oߟ�aM�>�W'X��z��Z(�kW�ZT|�ZY z+�G��w��3��Qǳ����w��́�(}��� ����P]悋O�FXZ0}]J�O���T��B��ܟ-�fU�3�<�!��R��v�9�2�[n��&X]�H�ka�LR�[7o�M�E�F+<�����53�N���ؖ'�z*<q�	���b�ρ��6�I�����-��PN�^�&�� 3�<_Na#���!��``�e���WR}6j�|dc�QN�t�#�aÀa����#�I�|Θ�<���CiҜ��S�>��=��m;��C>n�S�,ƃ���	�+r?&w�i��w��G�&�Y��ﷷpN�8�E����~�-,y`����������!�?��(�:��Li�$@�N3ý{/�<s3~�-Mm���(/�\�u�  �V�-� c��#� ��CQ���������ʏ�gi�]\h��J�Wy����iZ��~�=�
�W�Xj>�/�\��~�>(!�YYY5�k�$n�*ӲɧZAi�R�)�3m����h� T��G1����J�j�O����6�I�U\s�v��Q6�e�i�E���أf0�,�7��OyjՒ��&}�'�?���@=-/�Py�YKY'��Z�z���I�i�]i��KC{���Q��R�7��� Ky�PD|tB�� �0�@t�0y~��g���&�v��!�A�6�V�x��b��D�k��ہ�: �bR��.� YT��_�;qS�O�GL�67l���L�b�y��<�,}������凥��4�ZZ�d����&Н�H��5�#r$���\DS���)=c�tD0l�,�00;�%L	��b��P����vq�e�VQ�i�L��8�����,t*]�4�>ȉ���f�6�h���~�G�OM�ZE�fq�~iI��@�� ��/�Y� ��j���z!
��^��@��V@T��2� �< K`�}Wn"��h<YW)˚'/eٟ�;��<�(��(����o<iR�0K����J����k�����/�3�-�6u3�0��Y�j�Gv��|vi���ǣ= ����7�'��~������Qz%���wߵ�������ܲ63ތ)u+���_���������3܏{+�#�@ ���3R�#Ɛ�@{i�2HÏ���xM$ϝ>�|:�DU{�>���]��[b�������E ��#<QP�T�^�{�m8,�v� WYC�Ǚ�K!Ļ����C4�Z�<jh2hV�78���db
s��^*i�x�Y�y�ʫǆ�$����⾵��7#��td��t����ͦ��
0��_m���̙h�w-�b����:>��M��2.��؎�·�"`c�e�1������I%���MM节=9"[3��-��Ȥ����~�L��{%GA�X(ߢ7�CB9������;��l���a� �Y H��$�J@��7�TA)�"6����H����,t��Ń�GߨK�M`Z�&c�3j���J�J@�o�,֣��\1F�uʯ�\�:) ��9�KZ�FM��ҷQ/�:up^y�������f�D�!�*�Y��*O:m����5� ���JK'Ɵ�Is�`����[��O�$�fo�^w������C�KyrEj�6ߔa����3��~(0"���3\�~�v�?2�����t�̳��ɺ|%>W����>����n���gθ+�bvp��p��c.����Ҙ
�x�"wԅ����n,����y��p��ⷆ5��q�t�g��Kϥ���/Zcy����Q�X�~���k��w�����vS��Ѭ+���(�m���!�
��e#b� � I�%Wp!^|�VfV�b��}'ߤ����=N�E���3a+\��%nw�h� �V�lY+�Z�@ �f����a\��/>�o��h�Z{i�6O�V�1�����mx�L�i�a6A���ݗI�t�b<XTl��4�NøC�V�L	/�N�Śg��+������*�}/6Yk�+<��䌺���%����4�0
�<�b������X�Xx���!��:����t8&�+iH���?��K�?S0 bA��9��F�~Kk�e�m���F�:L�sb�ߏ��q���NHk<��r��7V�PB_�F�y-�͊�̇kY[Y�)Ϛ�y�`~��-����Y���e���`�F��q4��;��/[	Z?��s��^�Zf��Z������ʾ���~l)����Ң*p�L�\���TH҄s-�И
��7�%��m��2���XC�E_�s�����
��ߊXMJ)��2�V{���o�</I��7��o�����0�[Ϥ?�nw2���������ϖ��5�o�-�)H�L
�{�Q�Yi|�	�������v����TH�d�$@��o 	&�����#�V�wd��@TJ� ��	�s����8#�@�n�__�膞�t�	��my�_6��++��TL�ܜ������ܬ�z�ȍ���OY�b�ĢE�}0�ߔw�����ӗا�cĦ@�����K6�8�[`O9'�93V��ubب��n~[��8�����hf`�%�%I6�B<�a�0��ˌO�DD��RF��y�lD2�c���R1����	LCb68F��L�4>�[C5�Ш���)C�\�&{M��!L-���Z�8�(�s/�
��6��+�1�HK��S��,����k�k(�p�#��)o��/u�J�R+���?i�|�x_&�h,56��=����3��2a��!�E�#���v9m#�y��<����q` O�W5�Y�����4�5U媞�AP��l�`���b��C)��sx���4�$���@��T*o��Z%|�;*--'��4�G�vɥ��S�_`{N0�f0L�z  pA�K�A �[o�eF� ���n�vmm�̛��s`s�OF r�4�P���Ǘy5[l��*ۆ�Sa��3�����X�e���6 y���qc�S3������]�>���rrk#W&�X`���x K2�}a�m� �庻w��z1J jRG+�ĨG�gb~�L`��!̀7�V^^�����)�__;Ȧ�*僤�fWD��u�A�L�r+r}cACL�E��lP�M�\D��H���	���wC5�P?�NT�P��C҆z��M*����T��[�=�N3P�f��M�R7�>>��'X!���~V��5�u��������>i�o��}�[�H�����0�-�Y��b?�$�D�*��Ǒ�z~@{�w� �[����j�^2�U0.H�e�Pu�zŬ���z�;ݧj������ΫA{hjb{�J	/��Ǽ�D�rBi�|�Q}F'�LT5~�}H�*��ID�B������Q�aR��Q�Y . �p+�5l.�8��fE���F'��;���(�+ ���@���Q� %�����35^��a���M䕕�eT�|s��~Ñ�p(�_����7��k�ac-nF[�,�P�W"�l�,NX�ċf���ϗ�<ׯ�(�;�MdRI/ς� ���@uk-�e��K����R�.&F�k��|�lG~���)2�EO�dic�>1"�u��J)���z��N=uc.m骾��6�Pd��14����0;�����4��'?5mP��+6W�pT1>5�PC)�i��u�}w�aJAsi����Q�ֵ'B���^C��������7�Q�)��!Sb ��uu_	m���{��*�I���{�<[�%�{Vm� %�L�<��}�NÜ��@���/�]�|9_��V��!���[�Ҡjn���jF�gŽ{��L��P������[K���-x�tcZ@p?�k��uV ep�n�g^�V'5H&��>���'}�UQ��f�03�
'��`O0�WV�&�:]�xq˿{�V4A~���>?�яL������4#��3��flM7���CKQd����b3�r�R���Gs���[�z���V��Ri!
e��� K���b;� ���?7����ؚ�2S���w�匟2���"-���ԋz��Ď�$!׸���4����B+ļ$�^{���M)*�%��e�� "���[���K�u�k"�q��M���PCU����cR���o�<�O*����N��y���]�&�K��UZO}�eуŰu=w�!��I��Q@�y�l���xm�tA��f?�תm~d*�#j+E�@���|�aN5��=���U�J������u��g�_<�����߻���a�;�}8}���������݂߆��	pD�P�JU^_�a��fy����y^���U���5�b�~e&��Y���a6���N���Ϙ%0`sk5��t���m l%�7?lhz!�m%�&O�/_��e&��Re�41���jbk>��0/|ɺ\���[������؜�=��F�{��	kק�+��ϤS�Le{�Tǀy�g�zFyY�~ԁN�H������G5�yJ{^E��i�j�����~��3�0��
�4X���%�}@,���j��yҫ4l��ۻ�C�u����I8��g�����7�C3�-�d��5��~�
Ifݲ��g���3���.�^K����ǫ��0Ӫ�� �������q�~Tw���>�R���^�e��x���k�~S%�	E��
��^��R ����*�j�U	��sn�`����Xc����6��i��jๅ�~O�sΘI1��Yk��z��	�F�����F��Q ��㸴o�Ҳ�uBwo/v�[d9��m�����8ϖ�'�-��.��ȿ����=����w�t6G��f5�Ҟ�j��i�*�T��Δ�`9졀4�P��쵊�,����9�v"� 
��z��p�[��ha˥֣>�N���Ǳ���[�A���q?VN^��(��S�-�zʕ��r��-c�ƃ5	���\|�e�!�ԔaN�*AB?^g��~h��iЪ@pJ� �a���u���AP�g5��oXm]��O^�!ˋ:E4čw̏��Ke$�k�f���c�����Õ��p-�έ�NVD�9�E�fp3���,���I�A1�в�������L����7��N��y4���z�n!��;����?Ν=�z�Ik��4���js~��Y\j�����ꄌ��AA�H����/��0��=V9d�;33kq�׎� I9�㎄kBi�i|o�N�G��9�Z�x�C�9�9��J!TE�]�߇��H<��|�;��@,�P��I>f�;�X#��W�^��*����}��e&�����q�d@�@� mx��O��ǃ�	z:v�Ώâ:mo���7�"4�a@��4�G��0�������3�-�X^>�{��UD����	������n�c��f+�a׊�u��;��my�PT����)���D�����o����za�ė �Ŧ���#3�����͇��|8}�T���
�=�\ܰ_�@Zlp�<T�{6�ILw��o�Pm���:z�}`��1������3�Y���%i��������o���<��q-q9^{�5���W�*���	��CÚ��ӟh$�
���^w����)��W -�D�L0G�Ɣ�N �nK�����/��/L(@=���+�p�ޜ�Ԋ�E}�B��S.���������o�<B�m�/�c��;�SY������iz)�CM����A�]�P�̇�c��*F@����Y���(���?b���l�ǎ���M`e3�[����\H�-��2i�4ؔd&�q AE���Ħ�Fw'n�l��X:#">wG�s�`\�	���?s洙3!?7�'�x2<v�m�Hu�D{V�` &V�LY��6�PCY�ZE>�cXR}�{�3a-VT쟞(�^Gl�o�� 0@S&�*烼h߃i@�;��/�8��3 �}\�{�ա��~�S'�n��y�/�IJ}a.���>�r4�[���N�	d�~J��S�1� \�����L��ƕ��O�0����kL��ďU�9�nLw�+�w�TJu�דBch���_}�	�xɿ�~��y���%�~Q�ߠ��}��s��][��s��\<�b>g�6����|�\i�[�q���6�ƞ?xlJ�Æ!,̏�|#�����D?��Y�u�VX]Y���@(�[�ۥK��g�y6<��������.��Hn�*R�( ���PC5�PC�E)h`���J R��ĸ�o�3��b�HCC��/���"�X`p���VR��.���4G6so�c>��'"� �p��e��� �(�@�����)��Zc�>2N [��=��n���)��R�G���t��'?1�����4�N��ԡ4{����4������~�y�*�;%m�-�������ws ?h���6�7U�����^%�Ư<ӣ4'��u{����)��<[�3����;f",���t7��Q��	.��:Q��Y����:?���mv�&���ֈΝ�4GP+k��ٙRBN.��}�Qϝ;k��#>�9������f��WR�F��PC5��AҠ`+u����0Ȭ�kzr�0�_���ow(,� 8i��OK�Ҙގ{�R�K}4h�T"ܦ^@�r�s_�R?|�cV@.~����`x�%��/.)�(CL�,��꒩4}1˯��teJM9�CS͸�l�����%�̼�(1�G�N}����V��80V܏2�9<���h�j#�Y��_��\�8�KY����~
�ŵ���naQ��N�/t�| ���Vi���0y�A���h���
���ݯL�mnl�|��M�X�B���HcY�;�X#yS�˪����x�\{�]u3�[�
`�-�y���m`+��b\��7��Ι�8i�Pm**ʤ�V�Zm�����w�|����y�g���FX]_�_����o���[J�07g��'����a~n�z���\��7o����Ek����N���PC5��tRU0�~����\��(�w� <
������t҄(e�\��{,`�am���?6p%�,&��d����>�{�4�"�f�/��/���	���
+0E�Ve����sf '�_�J�u��o�-��s,p����,c2��4u0n�ï��$�=��s�4�|3f�b����h���s�������+��b��/����ߴ팁�͸�����7�4�/�5�o��o >.[Ќ}�y�O�%�ꭷ�2�� �����a���l� [)�;W�Ʃ�
�� 0��kT�1�A?����:�!4�Y{?aG�{&�U��Ӂ>�!�w�eŵ;���U}����5 �Չ�w%<�� ����`q)���d(�q������2A$�eAGb��HH�ؘ-����irٰ�GP�&��"�eAǿ'�.`w~a�6o>s�o|���g���WL��80�b��ַj`wӷA�4�PC�#֬?�KU ��T���}.?4�2���J#�-�8h�@����7 񇯾~��kv��tnv��`|^l�:@#����k��W�VS>�2����U����d�/ ��B�ds~��(χ������X��JY���`���vb��Pw[�.��G@R�D͸1.���\܏c��1�[�z�+�� �.��@��sN��9�\�r��N�ѯ����q�E�n��Y8c�]��i��_k\8F|k�X��n��e�ќ��i�Q���h���=h�?;�|U)5G�G��Uȳ�粭�fHn��K��{��.���W�7lw���~����CȢ�7�6���;n�hu��B|?�����<�&�X��尶�f��h��ef�P?>l
��U'}o���j��âA����${ �F��� F�\���� 	�$S^�F�޲/�m�������R�&� �x܋_}�U3�U�f�`����\n� =�-��1����8/�'k�% `O��m C�	 r-��>pϿ��_[��ޟ힌}&�3u�S��8}҄E�%}�	7��>L�I?_}�U���o�m�w��駞�gE�e���| �h�	"��t�J�RT1&�Wi�Ȩ����w�!���_�����_��ԺS� � |��N��(�4��0��Jô;�pp��k����N:VW���=�=r�ir͗�B��D��0.�];G��� �7��
�S)-%�ީ\C�q�}�F��pl!��H�ɸɠ�&��I��" n� �G>>�>ʓ���j���K�j����?��:pe�c��r� p .��0Ƭ�]����}�g�	sjZ������ 0c��)#J�c�m�4�����f����]21�CY��8���~ �+]	�>�fm���U>�+81�9������-MSdkƛv�'�z� o�F�|>׮]�z�<{&�O�8  4�p���o,�H!E���q�|����pP��1�(C��;�bͽ��<	)����-���w핆�!�t�j���̓|��5��xՙ2��n�.�z(*~2���N�k��Y'�~��Y��@
�7�4�8@v���0w.lEʙ?Ӭ�8�I�1 �noٷ����ߝ����>�Y�n���jhڈ=Kf��>��fej,����B(�G���*���~����π(��`�쟀5��:hYeq�v
i� o/G�����M�:Z/�mx@0�L���=� �?2��{�n��4�n��_4�~�ͤ������_�e2n��rK3 0�R�0�)��ז~r��b�eƬh�f2�0ocɽq��<��o����'����c,��g~�ԝqT�kᙸ?��#�����_Ǻ���O�OC=�Tg�~����B����&����[���'�n^�ɽ˧����骝�Qu�S� Ե��'�̩�7=s���pl�;m���Bu��PC5��R?? ���� J�,e���!  �IDAT̢����h��>�ZN��J)D�@��8�J��	6��̝"�� �"SWQ���Ahv���? �k� M�/m3����|p }��u��� ���G���A�c�HP�0��H�XM����M�Y�^-�I̴�2h����3e����YPFf�E��|䋌% ���,ῂ�i.�`����AP��
�q��PC��2��L��`�uu�4�l_� c�KI9�66Ͽ��U������<����w��Q~��u�E�0��b��v�����.zaC5�PC&��"��	���2�D`�{�O�SVl�]�RT���囿�V����P�d6��� �>~�Ō�z�nL�
?�a5��|�-�L> `�Ž��	`���ꏲ?p�	M��.;�p	@����=>�	�2h \E�&�5m��<�&��*�p�sn�==8LǊz�h�9Ǹ��g?��*�q��HW+=wX)��mx��:��A�5@�zJ�=�����N렴G���4H���7E�4�e��t��%�nQ��O�̳m��B�k��}
�v����͂�PC5��$Qʘx�|��)���tH�Ж�(��H���O�4_D�F�HY��4��)� 20g	�3��@- �(�� �� �O�������$��G3��[��d�y?�YM5��Ø�F��8�6�'`������]j�1]��7�ch���Lkl}��p󼩋��4��dk.��N�4s]�F�nn���UB ��@�z��àa�+k�Љ�*�pؖ��Ώ:�t��Y���Tp�v����s�i��2f��s�)�}�\��H�ӹ��ӡW��k�ݾݤ����au�9w�ē�'���j��G��1�J%��4�R�N^J�k��I[�r�.�k�]J�B��A�/L�僋9/>�
��v�����>+3`i:˲��7>�\@-ZL����6��`O�����-hG�R(16�c"~��eӔRV�9L����Ɵ߀V�#%>��m�����M5��_x���:����!��:��k��`����<c�&���<4� ����q`�0��+�6�O�+���p�����c?��P�����m�9�|�BԴ�橡��IB�J�Ls=�kn����L�}�<�.�y*�L׿A{֤?�Y!����ܡ�d�K}.�:�:��dq���П�'gTC5�PC��۟<�j����9~Ugi~\׵i��<L  %__�� W�0��כ�iH����a�f��A�0���G4�hYi3 �>��Їo0�]���h��~b��1�G�����~���-�@V� Üۑm�d�s�h��+W��~�h��� |���0?��t�f��m�����y
OQ�eV-M1D�D�~.��v��_��,-�Va��o~��7�W��{�lO1��	&ҶslҨj,����/ì�CVTk=Rw�׽�����*K
���N��N}w�S�֟�F�����O��O��5�PC54I$�h��_ԃ+o����:M��6�o�Z@$������mK�� a����*PV�D%��A�����`)Z���U��!So4��NLv� 8� T� �T�7��	L����
>EYR��������_}��qf6�<���_c!�����&$ྀi�,�����63�hv����,5��w�)�4h�|�M+�13��vB���5�A��ԓ�pOߨ�����>��{"�`\���d`���S��=��U��a�,�iW�L�z��&��������+9�4�|u�	t�3�|���z�׍��$��Oz�Q� ��Z~�ԟ������F�=�Ƣ��{>VY� ߆j���&��O���� Wh�  K�V����QcEEV�ZL�e���l7ڔ��Ἦ�oʥ�
���ި_fЊ�|��+{����v)]"m �c�˵���E�`����h�ѐʗ�_�/��#��|����r`я ���[�~��Vn�L�}��	h&��s��ZJ���8��<`٢bL�rSo����})C��y�eY-�G�O�
����3Zf�9~��)r5�P*'�t�����Rsh1�iJ�~��Ͼ�B�T3>
�9 M��:�0��6�4ցD��L?���GS)LcA�.��{+���ö}T��s?��Np�¼8��awט�A��n���j��#H�z����+|t�JX� ��8��Y�~��߆?������(e�v�� L�դ.�����(��믿n Kit<0���o�m���y��q\ZW4��zV��#mZ�w�}�4�|3�m��2�b�8�5 \چf��'�2�`L,�x2��X ,�/��}�@���� ���[6>�\�� � �RZg/l��Ҫ<�i�m�X���p�{P��?��i�y~�Ѧ]��o�� az>����@0�)������J�?0Ɯ�~��_�!}��Ai����Lz�Ao�S{��Ak������O���9L�bb?��b��L��XJ($A��m�R���]l�4 �Q�m l�K�Z4*��Q�� R9e�w7���9ݗ���`s*5�PC5��"�� V d'o�0��T>p �Y/ @p�,�	�& H���O+���߷k�K4�R�S�| � [@���GхhP@�Vy��bt\{�����{x���9Ni+}���;��q,
�e[N��S=���d3��Y�	�ݝ��U�3�$>������rl���T���?� ���GX߮�%��7iؠ0w�xژ�iW�")�篾^o�a������)m�7�}�O:�[����Z,�9妞:2���Ro&.����+�-2O��s,�u\�/_���Tq-��V;~/��V���<F�q�r?J����K'|�N{�����T���\��J�s�^&Ș(#6�֋���D�h0`Ho�I����7=��:kp�8s���e�n	v8�c>4��꤭��*���|j��a�|'!
:�I���@�'�b�]�$c���-d�Q
.+.�d����<y�������ԁoɣ�`e�"���� �i)���`Ȣ��(+����������$ے��?�48W�l��4�Z�8+Е�9R;���c?$WQ���R�֜����q.��i�r��_�H{<��qhI$��$��ڂsR��H� KK@Yi���Z|o��b�̱�m�v��쓿�K� O��cI̥���z8u/��t5CR�cε��<O<?���5ZC�%�t�%_�R�y���>�C��tC0��]���vU�B/YG7�����f�BՐv�H��b�]�u_4��}H-�����}���p8%T��ioO��%_B��$�v{��%�g� 	D	�e-����es��`�$K$�	���\γ��L���0K�U`([o�g�vP���t�v�ѵ�H��U��`2�|+E�V4mg�>u|l�9��%/�Lن5�v���3���;�rJ*i�)b��� �j�>@Y&/��ݛ����<]3[�����}M�|��1�5��NC����:~L��C�S&@���XX��I<�&� �l��&�T��Z�9��)���R:��O�NF�Ha��Wב��p�H~���"�D��,��dtE���kB�W��~׫ؑ�o���:�n�SF_����[�Y�I�YwR���4���/�����;/���t�� ���ׁS���_�e '&������Ur%��U9��H~�#���}��9Ɂ	<��ZX���gh�)h;x��9�n��ה"i[2hIo�d���1�@N�B���>}J^�y"��)\Ȯ�9s�RU�h�:�^�ۺ��BxT;�|.?W�]���ہ� i��k o��ƶi�Ө�3���T�ڍ_�ݣ�)U�#�0��'1�,�s���{�l��f��|r��L�ɍDd9������'�p��W9�(�!�)�UEcԑ����D���H�o�n݄�冭����I�ߪ�>]�]׫p��J|I��o���:�b�V�lo�<�!EQ�Db�i��	�Tz�_|�'���������9��PZ�����"`׎�|(4�R�.V6�AC��
?S,��+Js�1��T}NŔ�lL�8�]�ӡt�)bovȹ��Ү�]ژ��Xݙ`��b������
CёK��c�}*l�����\�c����"�.��9^�k����&�����@���M���[��z�R��\!bg����A}J�����zS}�U����&����6������6���DH��&6s �R���os���#�I�b�p����]��͆�-[_��ꞯ������p8�"J3�֒)	����_W��Z"����pƶ���	���BL*Ц�g�<����^�A�������7��vM(�d�ԇ6�I�K�+��֢��0;OA�9������1L���?t��E� �8��ÒI�8�<�ۜ�(��@�-%�c��������,�2ܮo���N�7�wm�\/jZ1l�!HA�	=�3�d�mg��)n�HiBb�K���;�lw�L�c��wש!�f��Y9���ܰ�LX�U �H),�|����7F��|�J���wH�({�X��y��I,s��ka�n�Xq/RW&]P���k~b>��n+�t8��)��CǔT��ؔ�wC}�`��RH��D���8�l�I?�aCF�)�ũ���u�ό[�"�ŕ��ݱ�]�txM8����,�}�	,�_,�$�#|�6���i0�7�.�Y���nKb�u�����.VӒ��/Xd�ZZ�m��%�>��yc/`���p�m��Xn)��k@d%s�yC����0f��%����R�}�[9��^��7��~Π:���Ѱڀ8�{�����A� ����@�B�K�J��SQ*�M7'��,��������+�S����>�s���YPV�XWAM�� �U�&ØY
�߿�u�w&^��R��+dy���w�`�p�AS��O�h�;�ײpy��D8�c:���nZ���U�}?o���|Y���x-(���9��R8�(c���_�vJ��!���%�<��Ti\vq��b_f�H��S�fV���,��)���O	������:[s�D����|����Oѡ?|�P��L��=� k�>����Y��Y*@j���o�?ï��v��$(�e���)���i�7N�ɉ��SE8G��S�ޤ�ݩvݗ�ty���;���x~Ysm@I�D�E:?g*ݷ�)�?����FjM�����{ж�UU?�«�&M����d�S��v+'�����o?^���Λ��Y���ʦ����@Ǘ,�Ia���I ˩��q�f���0L(T����>>�U���~�zD�<��&2|�|��.ܮ߅��*�x��Xh��[�����K�~�!33�jD���'~�$�tK���{�%	Y}��r8��%�F Mӿ�w�o6����8�r���}ɐ`V̐%G�`��eY�A���k>�<���e�	��DTǩ��gѵ����(��ͯ�;cX����0�"�mL�mQhK3e�/�V�6���
o��?�=�VK+    IEND�B`�PK
     mdZ��<�`T  `T  /   images/69c28b0d-a0ad-46f0-a190-03e6ecfe42fd.png�PNG

   IHDR   d   5   �0N  0�iCCPICC Profile  x��||eE���6�G��y�]�$�{�R�f�IvC�]�%�l�l#[`�H�"Mw�J�"�T�"H�&E@`��3w�N�]������@��79�Μ�=��{I���挪&��y����L��ǞՕ^IF�u����X�����#�Ox���{�%��H3������;sp�@�4,¯X0��Q����- �~��{?G?K�0��g9z�xǓӛ8���V�)�V]20}�n�$���^�0IV�O���Ṡ=a`ͻʅ��;s�̙I�*$�̚�x��ci̹���A��$c�Z�?<+I����{�\�FЭ�m����%�����<���L�Ze)cͩlf���:��լ�y��C[7MV2M��4�9�5�kʴ\����Ӕغxx��6���Y��"��t%,I��]�*��,iƫĿ,1h�HZ��x�*��&��;�%��I�8S�ׄQ�u ���M��{���K�<@u�ǵ�1c�%m��&���_��^[�/X:<4k��j4m��>o��Dғ�,�6�~{��ǆ/<�����{Hl;�$i����6�Q�\�`��}yl���d���䶶H<os
�R�^�e���vLrjr^�<�6�-y y2y5��a���D�.{7�pfõ5�6j�Q٨�u٨'FWF�0z���F?3f�1�c����M��{�������J�4o�ߎ�x����<q���X�UN�����U��j�w�ֲ�-��կZc�5�Ys�5���'k��k�θu�Xw�uo^�{�W�?�~��6��l��F�o��&c6�vә�m�ك�[m�b����R��~?�-��f�׶�f����ŗ_�撦��;�֫������fױ���`9G�g�.;mۮ�������p���|�̖�&������4~�;��~��]�w���ִ�Zw]�}i���'̘��5���s�7.��ߞ�w�^o����3�ۇ�:b���6�7<�w�6�Ȃ��wZx��K�?p�����!�~w�CO9|�#N;j���=f±W�k�?z�~'�;��S[O{��#Ϝx�o���ܕ�[~A������{~���/�����g-WO��랺�7���C���֭o_�w~���w�u�=�w��>���G����d��G<��s�<?��/��ʌ�����oLzkǷŻ_������p�G>�+V�~����>��kWrQ�aCo�u�6u��7F����5敱�[w܍+�3�:��o����q�������k^���k߾΃��y����x�57�������MO����_}�1��&4Ml�b����Z��q_>{�˚nn����W^H��>�b�\S��76���m��j�ݶ��C��{}mA��Nk�x�umw��ؔ�v~��cw٤Cv�:u��.����Wz�O�r�λ����=~��/���7_�֊�u�ڪ����͜3�p�f}g��C?������s�܇�=;�����p�EM��[��{8�t�A�|�!˿s�w�;����;b�#�G���|o�cf���#����x�'.��U']{�/N��ԫN���K���r�yg�u�i���Gǝ{�y���\���2|���ɂ��]����.�t�V��uE�\��U�|�Օkֹv������冎w����C7/��!�}�I��s�%w\��_���>|�ӿ{��7�~�����}����O���~辇��í�\��������'���'>����������n���]��U_���F�<�o+��ګ������׶}�o.}�^����<��'����m?��Ã����n���c��_���a��Fm2��Q���Yc�{ĸM�ݱ҂�ی���wU��rƪ'�v�ꧭq��W�u�������/���Fo�ކ[m��ƻm���'n�|�;�O~�/����Ħ-v�r�V{m��ˇmsJӏ�^��+���gϱW���ߪA�dV�kl��W7�n���-;N�ڷ[�O:����?n�f��Nyt����٥���ίN흶���]/뾻��cfL�m��{�q���o��[��{���x�l�m���}�f-�}���^���s��Լ�$��1��B��m�nKfpЁ�/=�퐇���w�=l��7;��v�nG����}�ǝ��K����[N�������ϝ���/���鯟���>�ݳ�;��s>�ч�~p��x�G~��A��$�|�����m�.���/?񊣮<���v��O���k.����n����w�#7>yӳ�|�����[>�������z��l������~W��߾gֽs�s�������>t��G��GN|��?���鏟�������>���9�f�_vyv�粿6>��c_x�����ˏ���Wn{����������eo,󊷮���8�����{o�k�k}8���Ώg~BH�#�Q�Z���>�ר�G�ї�i�_{Ӹ]ǽ����g���ʯV~�ʕ�^��٫��ƅk^�ֵk߶���>����_��FS7^���޴�3��_ܲq�/�3ሉ�mq�m���o�n�6͓j�}e����v6�D\-oU��G�3�o۾�ݘ���a��k-3'�z����~�ӟ���>���b:v�\:�G�n�z�{t�����f��Ż�f���\�͍�%�=�o�^�������|p��}�����7�>�o�9��m��������?|���-[��%���_?(9x�C&|G������X~��G=~�k�4��q�/�o9����0p�ܓ�r𩇜���;��}�1g{�������=�S�?��.�鏯���~�=���O,���G.��e?���+N��ȫ��Q??���9��s���/.���n��������7��WO��̭�����o���?�͊;G�n�]��W�g�{W�o�}�����������w<rˣ7���]���O\����<��ӟ>���<s�_�x���������^<�3^��o��r��w������X��-�����o���a��޲���]���g���Go}��O>\�p�����$��W�x�+v|;i��v�A���b��$+���O��ϕM�i_J	{�?�d�3�9V�qi��=8�?b��}oJ�2<88�?pm�|�A+6i����4�����c߲$�UW����Q��5���3�%����e��@����o����	���u}��_�{������ہٓ��z�7^�34<�W��M��(��y�Q4~���	�Q�x��׳�
�Q�uo�w4�)_������������=�� ����3�	���1��ch[��������1�����;%}�y��H{)��P�8|�/G�C�9����c~B*���~-~9������8�$^6f��(SX���t�{opPk=�#?�w�J�u,M[��I2�,�;�ڒ�I;�lż��[�{.r#���F�m0!�OݚZ�O��c!zP�1��1�g�i`7m��A����Ջ3��įyJ-#w��	�x���a�i1ֱ�>˝8�A �!���2l�¦�]IS���Gq��k��m�')ᘉ144�d�2#ѹj�g\������I�$�d������I�3�)������V��Io18�ªF�.����S}H�K�y��o�9 �fH�#���a�_�-=z���;u�e��O?f��>��/�����ygo;�V���䶞�����i��Ɩ�YK�̩����{����y����Y������U���3xn��X���>�}j�Ȯ3�.��Xi�nk�m�\m��_T��_Ze���m��V2Wh��3�[��Z;Zzz����{�:Z�h���O����7��������nZgWߔ�=�6�9������cZw_w[W��{ʤ>���JoK���޾��=���;ۦ�Vwo�Z4Xʪ���9�K���7U[�ϙ?ܹx�~C�����׻GW�ݩ��g�j��i��ˤ����v�7k�ĉ��t���v�t��:�wBjS�s,��ur'�6ZQSYfLZ��&�f,�f��eJYf+S�uw�t���6��wZ�}Y�V�h�i��h��6��czo_+&u���O���5���}RG�g�Lj�I�A{tt�AD]��v��=��%���gW��{�ͭX���@(IԪ�8�E�3�-�$�i��fj�ƫ��fV�o�쩲ZVc���N���Xi�:�t�ʴI=m�3ڠ?��Y�t:�8���ul��so���v�7��?wwC��i-m��܎���Z<s�ҫ66�xz:�M��ySWKo��}=m�NoñT�u��w��/�0��6KþHE+S�wNj���Fvjo��S�^ē[z[�v�����tvu8� M�v�Nq���d����=ܿ{:!��=b���ޞj��9*�;�O	ae-�ˑ�5m���v-�kZ5��A�xժ���U�j\�TU��p>�?�'�y�ʈ�3�,�"���&��*����jF()����(�?�)�+�*��헱�`����if������Wߏ��폣#,R���Tl�s}?�j"���^���6j�BK%KK:[���3!,�X�#��Tq]�FhL�;t�<�2ص�0�B�1�T�*SȨ訲��;�U��4g�E� WX*/Q��Q�,�R�V���W�&��Q��]���L���t�����Q��>2Yr�E�@ڌ����h�N�c��d����SS�IH+��"}͠yZU2]r#w��dF�1C�R�V2�C�;5nG�%��P��:�D�l4��b#�e���؄�n!ӌ����Y��~�a"-#���N��L��RCH���L��t�	bK�;2iXfhaIYa�jk&�L�� �*s���-Պ˨�e8$zTPB��dF�\2Nrˬ��W�p��=Q�ϐ\a3Hڱ�
Ù�֌c�'0�`��X-�7X-�<����i5�S=�jLm.�GB	�rH˰5�u��J�*\�N�8b�0�e5�H��'OE���8t�tC+�b�P`�2�_G�@��K��h�(��@�Lׄ��'�a,ܶ��H�Y�K����O|tZB(,�Y����Y��5t)K��p,�|4��`�2�DX�ܱ�����9����`�$�J��s'��fp'4rYc�l��@P����AjI�X'��TX��1�f�`Ka�i�q�Daͬ�U�ۚ��:"#���+2xr���`2�G���VO��+�|�G�N���q�
�Bp�N��zlL���R(-�Xr�U����=Z��z�R+;��C��x(�+lj��� 6KDHN���RؐU�����#�o��?B\�� 6��`�h]i	3ѩ��ㇲ< 8T��p*]G�L��
����3tU�FZY	A��*�����*@*!)����3�5�!�#�8y���P���#���4��G�Q��a��m���@��4�O�b�Va��La4�j	�%�����sKR��"2���I3�	�	djA@a�z8bBZ����R5l#-#0��� ��=[M�� �O�������:� �}!��'U����H��	�K#SY��&AJ��BG8.V�r�����3@�)�E��n�H�g���#H������r)&N
mD��M��:B�#f�VaVP=�� 8�
,� X��zB���S�,I�Le�uոF�u��E�J�82,Ug�Ȋ4U#�~c3 +��%� ���R-�#С4-!�aN��W��lM"��w�u�~�	!g	�}!: ؊ʪ	�%ͬ'4�6|��3򪁓����΁�HR�z#�;9�0&D�j 2,��0#�'��0n�V
@2�ei�:
Gk�_Gg�wZ�0�0�=��
�����H����`�kI88x�;����TI��:x_B.�����U�.�"T^Aza�X�)�1r��ʔdqFV�+Ek袁����%�Ṋ`�@��$�P��dP"�iI�St$?�p�Q��a��`�8���"kD2��?	���SV���=�w�_��Ffjd:d���*�����:B1�&�H��]«�E�ˎ�H��ړ�E�p5h~1Q}G�S$q������!���ܪ�����B�p
���	/	к$�ǁ@	��q@�̳Ba���e,�qF>�.��!�Np.�X����9�T���I��������8���!� $mG@��b��8���j`�@�
pP�=��)+�ē��QPG%a	J@&,��(L��F�C`^[�R!#Ќ��Đ����`�1��3��-t�Ȓ�����.P��I��&CA>�pTI�u `:Npy���RE�-f�n����3$��"��rW$A�&-�jJ�gGNF��� P�N!Q�[�b�{kT.%E�y�������|�: "r�EsJua�*�����\�h�C��22Eq���\|E�d��*r8GFi�zd�by����T 02��4P <��a,� {՟?#�,.��Ud1CE*XŎМ���*!j�����LUt��XU�1.��~� �
(oɬ��K ]�K��H�R��=�T1J�B�)q�Q �F�{4�k�Qj +ǖ�Ǣ� -l��9������diY�)�F���3�`=�*ziV�3.�TQ%OQ~&U^�L���#+q��ڦ%o�H.�z�H��%�5*\*rzF�Ukx�	 �z��U8�`�Zr�H�r[���^ZVE.V6�����P�.=$���eu�'BO@.�:�		]GO�8�9�*�q犒?�����r�)*��e��'��APM�<��*|���֖G�ZJ8d���K9׬	�W��rr�
�X��^�x
NZ✰s�YVO�=	;�dp�]�ӦH_ѓ��B c
�M���x����D����ʰ��PM�Rg�%���Lu
	!.#�4��l�49�R@�#k��=���Gғk���G�7z��Q��8O�8eje^����}������i1�xA+�Pe�)X6��� lܧ�Q6�ٙBl��Cќ��g�L)U>� �*���@���2	�!�ecJ$YZ���SaY�T1B�
�rA��Q�R�F��+�Ѳ0���9�L��)��t�ʞJ�U��K�&���\�0�.0Q�3T����*~�*2T�}�����zO�oJ5*�P�`9�T%^3j2K	�T�2N�mI��.�Q%�8H6lH��@v�D�dkJ�eѓ������Ch��AO[�5�*�'$�(y�礷�4�)�6�Y�$��-�	E7h$�?Nn����5�|W�'���d%ޤhAb��@��p�F���	�l���'M�w�0����<��HL�x�(!���t(��t
cq	���SD��s�OHN������9hp��FGM�T����ܺ!�AHka %=�j���z�Y.[�|�{6�~f��ڗj�
�H/a̤�$\��en��IپѮ�! ��
As�2�OX�QퟜeJ�#���Sde���*����<�*דe��dd{�$-!0|�����ؚ�j�Y��d��WKuGX��tr���F�y��>��EX�9���K�U�r�h+d�q�j������x��e�:�!�zF\,���V�P��9u	֌��!mQAO)X6�>�'�iJz�}R�����@�	���@o�-�#�	�j�m��(�i���2㊚��@J���G �8�Jz�-�Ee)��'U�8�s"�K�$+�Y�jP;�R���H����%�6�*l���)k��<|YA�)E��-zRI�%�B0Տ�t*�S�X?bvʌ{�.�ӤU�C�T%=��a`��ӣ�|NI��,�Cq�4g���m������)�'�-%������yM�Z����$W ��gĜ�QO�!!U�:�	��=��s�|�XV��0uT&U��_R\�G���)�г�F�	�A���aD�L0唝C�/�秽	��<x��E$���D����j�� PL�,�E$�&J�D��0 My֌�"��E�h��,�*d����X.�;Iݜ��J��k�i�a70��\�T�6��>MY��	 <�D���!�/���e!�Є����=���{f�t���'l�c�.
��I��,$�G�P}O���hr+&�~Nn��n`����i��פP�f�b����jt}O*	�L�,^���ԓЛ%��I�� N ��P������ ����e�� �p�L�*t�����N\240����=�����z�����^�$6,7\�d����V���0�{�=V�g�YW��Ɉ��-���Y�y �K�U���dPt1D4�;`����DO�讑�HXmޝ��5{�������?wh��>&��x|��������G^���*K.I��K�t��������4�:dP����H���H�#T ��{�JIǫ�S~%y������ h�/��\+]��ܓ\�Z�R��x)���"���D��c�����U�hϵ*:u�I���"x#^�������i(�ʽ���v{c:��C�-F��Z�I�����YF����7C�ܓP>'(�6�KK��V���rNbk������(�V	hH�ؙ�� xG���'vҩ'3����>�@J�xuJ��]�ͰObe~9�N<W�M�|6hDrR�r#����f�5�(=i��$N �t�HQ�o���M^�j�#�*_��õc/�A��)����O.(���� H3?��t�x���4�<	8�G���+�$\���f�̌_�R���r�p�9�?BA�7�F�T9^�2g�)��'�Hs��HL���8A�� ��ۚ零,גe䋤��61��taF伂�3g�������ʜ��o�z��V�F�7+�n��.3s���K��]�|�J��Ѝ�8�;��q�/RYDG�QE/�u*�Z5L�g��t�Ϗ ���,7͜���'��Z�x����r�.+`�ĩ�n��Q� !�UH&o<��7'�4�U�+��kԊ���@�T��eF�����^+h5�!�;^���{�X�C��C��� 9�ίݑ���@�4��u��Y�9��+H/�&�nq�2�	�ȯu�d1��+9�M�l=7�)xh�T8��M���>a
E*���b����
�IhWn�E��j$S���o�.�K�+��X�R��
 ��"e4���ר���?�"��I8O��+DՉ�Aa��'�:�zI%d����ݞ�ys��[--���^ؓ�Y�\�D/H�DR������b?~0I�ϓ����C�k%���Q��y)�z^���!E�Γ�%�$t�xYD+oR�@f�P{�y�!?�%��t{*'c��%g�[�t ��n e�������O�I�dA�G�xe~A�Z�~0Lt�H�����ێpL���T��*��y��`B~9V�`�y|b���<�E�k/��כ�je.�y�Yo���qs��j��
I3�I���y������g��z}`)=%�y�������R��/a�[-��� )� S���]�k�>�_/�f�	@f��Y�0T�5�T��@�ԯA���,�K�t�5�<���;o��̸�6��Ht��r��Z�]�Ԇn�3^s(�Z�(Ȭhu�s^�_���w� Y���cO��10	�)�[�)�7r~0�% D ������A-��)��L=��0��n\x���@�5�)>µ$bk �6d��Y0�	r�y8R�\�<bFK�ޜ�U�[`F�@:�8�!����pR{�����GÌ���	�H�<o�a�h8X�d�4>��aA��y���*����!�����F6�*�y�0ٗ�cH���Z���a�n�$O�g1�����P�D�j����Ѓ��7���"��{$a����6b��-0���2�;fȨr����cz��@fao@�1M+��9�[�V+�z#��6��b����O���0ئ��	2�L�4�g���0�KY��GHNI��[�0o/�p��yxeP6La�#$���pł#��@	£�z1��}��ȴ��ĆxН�a8%�~�Ȕñ 'h?n�0nһ�i�:Sx�2��@r;�!R#�a8��c */I�a=o�a����Mʤ�k�ƹ����0�),�f���խ�Kg޽�.����<��X�v�#� o&<o�a�~�
��o=)�q#���r  ����E�"<�'2����rވa�kK�Dz?)�=��@Hʻ
J�6-��T�⁴<�J�x,"�p�Ap
>fa�J�q#�4Ͳ�aCʺ=�ټ|#�����D��*#�F{���2�w
 U87Z�_o�0�|����7S�,�mHD5U<�Z�CNJ���a���y^)����SE�04���
�~�>:�y��a�=�,�l�y��H�b�<����d�tg�������^��0��>���a��� ��ԍ+-�����މ	XH�T ��ވa�+B7��@B�r9Ȉa�o� �ӤB�����g�ܬ�,t���(1t@z�����Ւ
��>Ȉa��ZRp�*S���1�D����o��/��LF��5`p�������`��JŞ�м"��T;��rO���@d�0�����
#�u�[`	�*�*�I+�<VFC�-�@��W�,�Sd{��^s�C9o�a0�I�$G�y��?��a(���i�f� ��a$!.H�2�|<>��H�_A�*0�1�:���'Dw��"�A���R��{�,#���)yH+�a>���H�.���9I�L��"b��0.`uX}�Ï1ZC�����=�����:tCLR��T~àU��
�WF��v1�A5`�q%|R�HJ��,��4-�v�y3r
8���W�o�a��PI�,ر�F��e�I�:S)���Ak���2:�"��-0Z�<�D�g��sSà�����������yC�}_cR��>���|MAE��>H(`�i�k*b���_Ae�O�gY�&�"��O��@���1���BE��)x�R��ރS�������x��OY�:ӾN�"�Q���p�W�l<o�aEw/>D@�;�U��8*bEy��K�t1�x#�Q��^ri�~�=o�a,(���8��vz=�F�~�!�T��G��y��Tg����0
��?'��Ǩ�6#��v��/����/߈aa]0�B���X1�,0hHj�*b���^��@�P�R�`��0h܊���a�~�O��\�n��>1��9��t9�y��(k���7S*6{���е��`�' ���#��pm~o`��`0�sH1�Ί���{Aj�uRGC��Ҥޤ1��8UGC����T�����a4}7U`p1'��up1r���K�ky����g:b�|*��^$�uC~� /1Lx�����g:b�qo�#�q)�;�h�>^5�i�b�3���a�^�Oa)�
$�g�7bL!y �GP�i��-bL�|��y� H���1�PޭhE�<I�sވah
xU��Q��c1C�FS�ɏ��w�1�~R�TC�1KG�)����ݐ�r���a�<��C87#��/t�0T����i±y��#��!�j��?��M�wL�0�>���[�U�L�0hUAa(��Wf�^J��0huO�2Q��U��(B𴆊$���+ӷ�x]7�P�wx����t'�-0�zC7��0��y1�f��>��I+<^7�P��;�$�{�D��"��V$���SP�e1�c�Fp�H��&b�
�4�
�M�P���-b�J_7d��|�Dcx�쀀����j=~�à5�����p ��^'M�0��K����㐉*lP�d��&b�߇�TW�����>U�ݕ�a��W.�u���;��F�1 ���&b0J�@NH��xC���� �I��}��Dc�{����k�����DCu�`8�Ӡ}�a�
*�=�F�c|��D���zhv:�q�0����w����R�ve#�!��^+��QXl�-0dX:�V�[�AFxc�1e�!y T�9[��)|�l҄q��ue1��/��l�O����xa#�J�>�b���EK�Ҭ�-0�ʐgY��#?�Kp���06sϸs�4�4��h#���4l��C�|l������\�#97�y��A$�BH�y��t���җ���s�P?e>^f���}/,�y?��S��>Y��
Q����-0��Jc�P��;��[l�0�A�0�^�2��8��X�ҍ��B��7�I1��YAH#U�Fj#���c���.Hӕ�-0�h��?�q���ECu��7v�����ك�MgA|���6b��p���0N*�-bk�2=�N8Һ�Q�[`K���y+?�Y6��.Z���k��պ�3^�N��� V�Q(&�[   	pHYs  %  %IR$�   �eXIfII*     (           >       F   i�    N       %     %      �    �  �       ��    x       ASCII   Screenshot�M_  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:exif="http://ns.adobe.com/exif/1.0/">
         <exif:PixelYDimension>512</exif:PixelYDimension>
         <exif:PixelXDimension>960</exif:PixelXDimension>
         <exif:UserComment>Screenshot</exif:UserComment>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
ǃۥ   �IDATx��\	��U�������N'ݝ����$��%�T�PAk(PK�-���*GgpFf�aTD0��R�Ț�HBBHgOw:I��}{���~����~M`�)o��{�/��{��{�����t�jAAAzǆ�?4�@��?s�O�q�L&������gn�5m��sz^?��\O$�=��'��s�����'�d>�,[(��q�`08��T*�u]���7�5�\�iӦy���~������v�y��H��o��cǎy�幻��۶���aT����:�7���32����B,Zt�0<<�M.�����B�4�a||\��|QQ������&�_p�8u�֮]�s�Ρ���V���ӧ166���y�B*((�&ǃ����b�ܹ�7'����̙3q��Y���L��=uuuH$(/+GWW�ܯ
�O���Ba�K�,�/~�����X�����8�u�%��<_|�E���t�r�-&�������X�j�b�;~����:000`�J����h�՘={zzz�x2g� %�%�D"����A�2������
��ىy�������R\\,DUWWcŊX�f-��(JJJ�
���F�I�����w�Ʒ��-���/��1x��سg�����BۓO>�O�Ә:u*����V棖��de�
�t�9sFh��-ƶ��bW�&���ϗy���k��1�u����bp�����A$�%Z�~z{�L�~<x�xVD�Rs��t������.�;v������o߾]����::�+��If����d������,J�O�8���n
��¢B$I��7�o�^^^.�w��Q��_�r%v���Y�g\�O�ʃ��5u��]�VN���������t�2�y�
Lݪx���h�$?֮�(g!���'6b���¤X,!D�#j	�U�PɳQ0����B��5�~��{��7�0 f��0_شɋ#�4�v1T�_���b]�,��@ȇ�Hf���f>�hѢ��E+����ɜC���3�I�x�7���o��}ٱL,��~�i<��S2�
���=���1}L�>M0c�����w?-�9��۷�6�#���a%�&N�
���@o�!�5kֈ[���a���v��!<���^?�
�鋷.ǚ�����#�UH�"�6P�]���˖���_�y5��)�<�G[F�hQFΚ5K�e�T@��D��~i����^l��|&wnڟ}�rh �gWw�0�q���C�'MP��9Gc�L�c�1��|�����$�82�~�҉�����8z�o,�Au���}�1�ܼ/n����l�^g���sB>�Q�WlX��Wcxh.������\���<H�@���ac|���%�M���O��Mz���?�;���:�o�Az����^v��98AL�x�`�21_2�Ea{M >d܅������%̇�����Ţ���9?0��m��ju6>�㩩(4�DM��ѓ��`��-�1�z>g�����|�U����V�k<"p8p� ֭[' C��O�{f�9���L��z��p+
�!	����� ��j�+�� v����iB�=p�]�Hl]��Ʉi�Rg#57��=ބ������Y[/y�e>4e7B�~�A?��CQqQM�'�'��ߌKD�!l����e�����'�4��1Do��tu���0r1I�Dk�$ɴu"�,��D�	w[�3��8�������g3�9^\Җ��+)�$7^���j�#O��X4�W^yE܊���DP�Y�h�J��W0��?Մ���G��GQ?�$��>.��Ȑ�pl2��n�(��/��b�m{Q���I������g��>p��xv�sު �߶�!�D7v�u71u�E�	��� �}f1z;�����+;�m�^�$U�S�Px^�~s��6���8��_��|doV��x��ۆ̴
�ߧL�2!�رǞ��6�5Q8Y9K3���.K&Ƨ,��@f�W^yeTd#�$𪫮��ի=A�.����w�ox(���a��x�h�)�j�qT��y�nm�֝X�0uxk�Q?'f���p�Hu��b6�}�jj��~饗T7W�`��{߇@\8:�}@����MO�>]a��Y�Ї��,��j���^"����D�H�d�?���Ϳ��[(()����j\{�����;���M����@�$�ј�$�!�.o��$�	���gz����r���}�>��	�ߧ@��[a����aU�֥��+�����	��=�h�|���Io۶M�}�Oki�n�L��n�,�ZQ��61LǾ}���+�r�q=<�`��9�t���g���Ͽtܸ��Qie������f�l�N��xOn~e��{o��������"��djM���a�9S+\M�!n��������:}&ۧ��2Cx�͹-;�0����$�����K3�XZU)�z�j�#��`�5xm7��
J#0q-�I�;����������E��V?���*[ vF��$��lү55>K7<{��,����v���7�|���^{�*�4!p�<���b��u8��chinFc�l�r�mR�y�Gp��1���0~��lz�}����y�����ؔx���s;�9���m7>y*��ق���Rn�ð�x@���JG����g����΄�j���L$CI�&�.�<�Q�y]-��U����ddkk�7�,���aDg���2�g|�'>T�Ջ��68��Mg\&�(**1�A��N(O���_�a:�����i-��)���4ݢ���u�E���U��ш���7���������K�d�bè�$�Z8t�gH �[5���<����YT����0BE4U�5m޼Y\�M�*���>�g���?x��	�5
�Z�9�4��
�8��X���S���R��B��y ��Bg�����m)�2�DabZ�@�����B=�Z��r�W���tP�k!�ģ\e��Ć���a���鐱���L�wcZ(@0��?M2�:��Q�d2��!�Ak1چ�E�[��Cx�u�|i��&~D�lncc�T��W����:?4�f�$)�9L�>f�*�xѪ��:{����A'02r���
��+82�%��船WQ�O|�1��]�V���ۢ�Q(�'7��W3�)���D��p7ݰ���w8�w���9�d�����֋p�g�=h�Ap�
���qY���s!_Y%_ˮ�ϒ��?��e�ҥh6�^�ڕ�����D]��x����)Y(�Z��������O������ѣC8��i�D�9iz&�=���MN���	�Qa��hYKK~����t��	|��_�*)�w�}76n�(��I"Wm���U�n����\47\Y�����P�3$`bJe!n�v
���[�;bY�$�{衇�*�]�,�'j>��(���W��9?��3f���s3
�Ѯx����]1|�.,,BIq�x'�+*�|6,���Ѥ%S����-T��HG��8ۑt+K����p�����t)�U�뮻��C�7���m�M�������w�2ֈ�����%2�䔸=�&g��3�
�y8N6x��i�̪�瞬dӶ^�z��/�Kɛ�)�!,f�&�E��kL��}n�#�.g|'O�0�tA[)��vva_S�1�"�E����G�벺����sg0v\��U��
r��/�aI�Uq�^6��B$}��qajV�i�!t0��CO��_?_���1����[-4��'���{�0ٸ9èT,%
���EN��FX�_~���ҩ���^�ü�LVz���+,Z�w�!K�t���Pҭ>�K���v�'Lf]��݌�?3k��၍�����8��_"a3����z���a����x�s�Kq̣���>��0��|y��jkV֠w����b�fWP�ۿ`�&�ch$h�(7HPs��#���#�0^N�4#L&���$Q"ذsZ�����ȑ#�b[��\�T��4�ֵ��I��	�@�gE���q��A.���z�_� ��J�V 2A�h�P���w)I��C�?�k�p8��hJ��0����_�F��S�LpO���'��3#�_�'�܀Ϧ�{�ĚL�D��Йֺ��9FV��n��׿�)z2a%3S�uq&�� �n*7��A�����yo�C�0C\�<��pg���d��
J=`�?5�<�����ȏ�Zc����1��V�U� ��jԚ�b��Z��Ԏ�~�d�ɀ�����Xh�./jb��~sc�=F�����������z�~^}yJ���>+��ɡ��s��t����A�;��.� &|DQ��h�册�~�S�c�/���EA�~�\����L�k�|� ��g;��A��tF]f|H����Sb�)�L�O���n���T����Mt���w�Y��;ObŲ
������qB)##O�%h6�Zh uv�I/K�ۆZ��6d�.����)�Ux-F�����m�7�p����g����>	�H�ןk?'~�qf�aNãC��KJ��4::&��
�`c�%h�њ��Rc=�dB�0�/�pK�0\!����^�JJ)e��#+��s��.�ӏk �ul�_׿m�1�p�A2��y�X*$��d>!���&�~�j-I�9��<\zx���y�5*:�

!ܪ3ݸ����ը�*���[\�4�(śMq=�!(�{�FFG$δwv���u�g`Պy��*t�'���w�=�&�PW����ńŅ��CG����:䷪�'M��8��\."S��u*b��r��r�eV)��ta����(K�ٛ�E��йE���s\O���1�SW0j��ͻ��
���
}�~�C��q���X��m�a8�.JN�.�*����k����p�T������q?k]TCI��_X�w�b���9�����:��ɂ�z]ݚ����)縟nq5 ���,*�y;��B�����˲�|��Mt)x�@���4� ��8�p7��
� _�C�a��``8᭮�;���D�f��İ�`m�,􅔇�leW?�	��0Q=�$��(��BH������7mͬRj��u��.�~�[˱Q�pc�l.P �y5]�bX���a��6��/����|��	!�q�&�������P\Tl�Q㦆�?`���O�+@W��(�C�q��7�����{������v�Y�b�����.:�Z���>�J���7��R�͠�8&�W?>;'��5z<�bF���T&�Ln4�;J�/����{Yjb�A!��dǱ\T�����gcf~W;S�}c���X�`�� ?�O�������c�O��٘p���a/�Vg՗�럛�ç�x�E���p��ϙC,a�i���쐉S�:k�pA��Q��Z����s���5�h�4<��0v�9!A�Bi�U����B�����@���m%l��t��R��;x�Q�Z�ޟ�a�1[8y�.]�B�$q���A*0�a�L[���r3�^t����BrkYNV��o�1}�22��J�2���xg�0�U �W�������gP^��I����o���:��颕�0�%�ĺ ^�c�����8K`Jy��G�ĤD��x���Z}�L�����Ʀt���J?F���ߟ�8��A���-��W[m���<�C7UZRlbKe=�����F?5�p{J�ƽ��dI����}Q<��۸���*Jw����\w�u^ �&Zf�ݶm+�y��n�N 2�d��C��	�c�Ḟs�'�n��w�G����4�.���,�s�8�N.���z����Qok+���~�Nى��L\�˦=�=h:zw�25U�8�Vn��
/�������[)����-6�2��߸��Z}x�u���K�)N����g>3�w(r�阬�{�}F���?�?bd8&�e� H�r����K`�aI��1��pu�����}k���t1��ϵ�|�� m��\�;����}�̕5�-[���L�a��1�;f�׃�=dLޏ��s�2D�����0��EgV�R�,7���1]��p�1�z�-Y�L��i�,�	���^P�d�7+_H[
�C�Ns�.������`6c��>����ڴ�7p��QL�H�/����EU'Gv�!�֮�h1ty��{�m�F�r;�%Z�����@��\����Ĝ��8r����S**+0��5�S�t���m+�I�����	3Q�a�=�0FW�l�L�L��D5�@�홥]�Vyy&�I�	\dY�P'U	2���
����'v�wz��\�Z	�����༘�0��*�D��.��2Cv�[;�;��2/�c]]�x|�⻙��zo_�r���i�S��|)�!�&>Y˝����\����]d���'w��$�N�\��jD�lX���ß�nŉS��{iu�b����$�Ӛ��d2����5�=���&���݌�P����\�k��]�r�2X��Xt�$2̜���D�=��u�o+��N��F�BR�]�,<��|�te<A��M���%8�ҎO^���2�TvE�M_lUz�5�բi�\	d�P��V�/�B�8�<H���B ��|V������G�[��o�N}���x���N�v�\V8�v��v̩�!o8�%.K_�ɥ�F��ݹ�$>�f.��q��˘ݝ��M'_a ���5v2�������3W��n��c�f����4��O~2��%Sw�A-�9�ϵw�S���r�iQ =�����v���P��m��$aB��/ǖm-�ދ�&�9��Ս�.Y!cI��Ὄ����9s�d=k�>;w�\�2�	�2'�.@F�g&Lk�K��E�k�S���a�Aw�eř<)h�`bd����\�9
��4r��M+�Zۢ�[Jm:����N�6�f�'�i�s�҉.ۚ	|�ߔzЦM�$;�ݘ���ԭS���Bg� �_���#j�b�e�=���mݺC�@UV�^������0������"x�J��qE-?��#¤P�wJ&l%�A�n��ß�t���O��/6���^sw��׾x	�^X�M/��L9v��#�J�IZn���p�J̚Q��ol���r<���ز��DJ-�ګ��n-$�����I���R*@����o6O Z��E�L��ƹ����$�o�w��f-��V[��rsn	-*`������uwP*���`;��Z�0p|���"���uxu�)d튱�����b�DI��m�c�Q�T��3��(.'O�����6/��Aj��Vgr��	܂����|B^+�	�p�wr�������Rs�,��F�c��+�ڧ�8�]�
R�౧�����W�P]��ġ�G
��X�*S\ar'b^~m'b�3�|�4<�����s{|��eI�Ua��w
��,_�<�*�Α	1��]�*O �;���7|��-D_?^~�%	�'�����ӟ��<��vQ�Q jv4a4n {/+!3�;'��z�|��E�s�M7�������jr�L&?p��׏��;�z��O�8��豱QÜ~<�\7�eHIUY�i�Ej���M��_6RQi��B�+�޸)���̟ہ���̑������)(,.ü��y{7�G��\����~W$K���}�{T�i~:�����Oh7M���.q��VBەil��W\!Ȍ飢�.���y�slT�uk�I6� �iz�INS˥�(J�N�#MJ/w6�T*�,��B�;�m}G1��$�{����1���Ƞ���~1�ܷ~��^���08aN�hAw�s�C�y�k$����~�-7�V��G�{}�Z�	ҷ�)��;��Z�����uj{�&Ҭp��7�K�;睫L��%��ubt��O��\�56:&u����6��B�S��`~�d9I��uх�Tb���n���2��i��{?�V�m�v��ǅ�wj+ĭ6Q�����y*�
VH���R6���0w��+Ԗ�T����d����`͌rY:}���seͯ��[�� O�z��c�&������K���K-��ӟӨ,��[�V�@�A��c�֭���JB�`�b�M�ƠOxLKџmR���*�'1ߞ� ���\a;�LpxpTV�r�0E=�{�D�v>5�s�_�AWIw�_m���jt���񂮖`�ej:��+����m�W����O	�� &�|ހ��H�tj"�D����E��v��������v>�z��e�7���ͽN(J�P+�
i^x���J��gP���&?}����8����,��/�ʽv�9�j��!�4O�t��X*u��T    IEND�B`�PK
     mdZ?�>�oH  oH  /   images/a038ca8d-f9eb-4e93-ad0b-b831193aa106.png�PNG

   IHDR   �  c   ��T   	pHYs  �  ��+   tEXtSoftware Adobe ImageReadyq�e<  G�IDATx��{�W}篌�-͐�_�K<aF�	�!���2��,�v��?vON<J��s��X!�c�l��q�g7ɑΆ�eA4�+a$LV^�0Y4��H`$�&X�H[�����.UU���n�����>��3�]Su?������BCi
C�
C�
C�
C��Da^���|y�!�3���̙�D_L�0�h�\�}�)!
(!
(!
(!
��,_�<|R����G�4%���wB��Ȉq+!��!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!DAi�Y����s���fj�H�U����?�[�I"���ĉfd�n�u�CH��R0::j-H��V�q�&���!YQJa֬2;w�2���aj�UnHV�R�͛7�� �f�����*�rH�A�ƍ͞={!�RJa�=j�l�b����W<�	@H+�R����wlxx8hÌ��mڴ1xmY�c3��QJa4�w��t4|pl��J��۷oG�t ���B�����n2�c3��BH3�^�c�vs�u�����B�t�0�f�،t �-344� ��#�v ��7m��o��1� � ���:�>��]��F�(a����%1��u�������k���Q�[��aZ��ߐ����pWؽ��{fH�t�0 ]�2���h�Ha ��H �!�:V���AL�gi��T�fvQ�0-F����{��F(�0(�)4��1Eƾ}�3�I�����ne�(���<�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�((�0X�k,W�����`���^n�����tQ٧�F��w�����4<e3��Hye��A
�ym�U�STJ��H�&�^�ϲm�h�wM��a�>\d���Y̝����-C4��`����300h6l.|�TXap�$�t�fɒ�ٯKj^?|���׉��ƾ�X���ā ���U@rn��ǎ�cǏ��V�j������{�k$����WD
'
����cEY�x�Y�r�Y��>Od�G�O��2�'&̾}����7���`����6.�b��P��K���ua�}����̓�
��Zs�e����|�>�!H��#x@lzU��z#�<�DB-e��s�����n[{!��j��A��c����G��`���_ֽep^e�i�װ�D�8P��<�,`������W�B�4�f����3\!�A���\u^���ݾH� ���3\\��S���}�RfwI1G%�jխ�E��s�h$2�Z�H�;|��L�~�����T>U�*#$���'N��wܑ�v� �=�]��c�\ǲh����e������Nmq>Q��(6"F\[�R�����Ê�DqTFG�N������ka�dA-�SSS�,aڶh�yx��c�1Y��󊨂��L��N��hHm���5\��=掠2�h��lz�f�#����]ԏ��������@�{�/����mՂdK���
����Ƶ_ B���$�o��!���c�S��p^}�Ka$��M�o�H�v���ip�����J�mHIҰ�)�4��u�/��v� K��Eژ	���8��V�/������эtD�A��}�N4 �Z*�o?d��A:pq1��{ר���~9�_nQ�?��9eօo)�W��X��4�ѮJW ��,�!M\\���Eͽ|�oS3���WT��^�z�w�=���
�<I}���+a��H~����P���g�\�z� �G׮�^\H_�\��z�m�4���Z �!*�����Ho�MvqjY "Ktl'N��SB R'�<�I헃&N��Ge
�{lڴ���aO�@Z�G��YY�5��]m�`ִoQ�>�(�Y�׸�KҨ�H- ���}� �B�b/DC�Z�E����pa}�Վ.��^���g�~�Ad�y�{�(�����=yD��d8�mAZ&m�jC���Θ�LT�m�$��i���0h� ��!��B�))dyQ��R�+5qq}Ǝ.�o�8�$�_*�aZm'-���@>e�4ۍ'�̥c���
� �'"�T������~Y�Q\$A�A{n�-�\�[�� �@~
cL��r��f #e��c��,@jTI�PP�=1���X�����~�o-���e�޶c��EeAdA�1�,e�~��0�yͪ I�D���~ �=��k��|�J�ŋg��"ұ��SY��+$¤�3�v����&E������JԾ�ㅱW�5a^��+���RX�2�Ğ��}:v~���t�f��2&s��I�n�.�+�d]([�6rg��ƶ_&�m�vE499a�Mۅ�/lVS6�]�w�4_��d9�(����Ʈ�a�9�^�ViT|��:@��I�%��0�Iۅ��x��W+�M=Y0QRd�ws�'����t���va��*=:ǎ�&�,�'n��"ei���K�=d�^��.LV ��Ŭ,>w�,��v�,�]X;r��"�Mj��2��G�����`������e� n�k#��x�!�/�r���#wV2ǵ_��Ο���=W}���m��������c��Ap�ȑ�s�=�n����č�n�0�D��,B�j�i�"��ݗ#�2�B���l��}���Oaj
ױ�{,ɷ}�EF��l&�n��*#� ��mYM��>nDL�3.���}��0>�R��}��v�l'��L���r�Q\�%���QЙ ,�d�/��""̾���u��-Q|�ȝ� ���
��t�&���[�va��kn������|�ap�"n���j���w��s�tl`��NpÕ�u�s���pR�%���6�����1^�����>�{�y��b��pK�������\T�>�hZ�cmf�\R���t~�>�>�i)x!���"j3H �iB�S|�ܫ!��o����$@t�l�$ĥ^����yEe���;ʠ���|��e��"~ ������Hw�6�D3V���~q4�����0 ��ls�s�P��&�g�9668��-[��ۇ T@v�n�����t~�ϫW &A�*�5�*&q�c�7��U�%
�Vx��<��-Z�PaOJ�\L��u���z%�IB�t3c�%�d��RD��I`����a� ��w_C�/.�r1FvO�%��y�N�g�C�櫸�(�󃋊�ݲD/*z����jj�Wl�d��z�1���Q��^�}�>�08a�D�b�'����7AVYV�qϞ=��T,
j�;�W{��&n�%���r�y�yD/�C����t�2��,0����pe��!ݕ�Hصkׇ��D�4q�,��K�`����y�V���b�-�Dp�R�1M(�,�Ȯ��pO�I����Ep�~�t8�v_�0_�%�0@�A��=���V�8눃����]s��)M�e�-��Kz���E�[�֮�]<n�Xk����-(R%�0 '�СC�^��5��h�ɚ�-��8I� �f�.P��H�Еo�Z������A���Ks��ej�=�QY�r^!�F6��� Bf,�8����k�gw�=Ԭq���'��~��,(����G��h@΅�̬v:?�+"���DJ�C�蒷)�0
.v,F��l�k��,:�#���f�E���k�����W�Ư(�������]���?�h8��^�Y�xͶǎUV�YT�I m�miw�b�F��x^'���nwق8����ֆ�۞Q 
ҕ�f����|8�����Һ�'챴�o�K�S7��PHa��(0.9��R\l�^"((x���+A��U�|`�<��%�k��X�^����*���ސk�&Ƀ���.�wc���'��k��G�:��w�[����Oi��""����X��XB\@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ�fdd$|҉0�����@-�[o6o�m����y�^`.��#����W<^y�<s�ET�y�K��x\p�)��y��k����r�gf�9=sּ4sμt�\�\g����_<sּ8y|��f��>��a0����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������8��_=h=?P�����I#���xײ�߿��K���/�2׿�/|� x�淾͐l�0J���o�S�N�'�9i��ߟ<i���Q�T�Ț�@ڟ����1W��'���@��]����u��g�q(L(�O�����
��ȃ��c��ϝ�sH���;�fKC����sr>/Dx�[�"�?�o�_�QX1�Q<����
� ��P7�{�y�[ V��d:N�/���"H�H<�����=�kQ�:-�Z�5 EU�ٚ�4O�D�����2G��	��/|���R:<��?������i�Dᅩ�V����%�#*R�_[��P����]Ha$�<����@/"�L���u�}
!�"���_�<�"h��kY��mo��%�; �ߞO��� ������x'ҭ�|��(I�k.�}�o}�*�Ox!�����t� �<����w��E�Aۄ�;�-�;I�N��a��?F���4.wa�r�fAź��	�:��䝲�"�������O���>FBZE�;�4��C1�y��W_y���u*��?<j�T(!.@Թ���>�կ�ܶ�w�/����>ω0��O��?���{�����/~>|,��uf��������4�rA����0?{���g����/�ϞgOiǟ����;~�\:���ο7�>�!��5Wg��-s�GO��O~�<��݆�xṓ����>�[���C��4-�S�|�L}�3��2��΁�*|�aɻ���l4���w6�>ja~:�������O|�R4�s�����}�4���?P��Z��=b):ߛ�Z�x���N/���.~��)��SBPBPBP�6���g�������qC��i��˗�_������o�>�&2��.9z������~?99iN�89�|�z��O�� FE��\����>9	���hU*F�t(L@o/
[o����5�lD��$JA&<�X�N�	���fY�nCt"S\�B�<xLLT�v�F��W<�)�>8���(A��KT*aD��c#GNH�444T}���Z�vQ���A�ש��OZ?��J��fI�x���URήԿq�\$�+�_my��
%���"�Zz��\.�]��B_s��;V��my�W����\,����@��;�b
�0�pk�'{0�^+��V�|-��k[�����V�Z�(�
�k�cػwoC��/����� ��Ep!$U�X��@���\7|U�f:V�wh������By�Nx6��0R�Tҭ�R-�8�7��( O�#�?���1-\{�G�{llo�Y>\϶	cK"��Q¥�Rr����(�x�"I��20��P;�N�p�GGG��m���]I��.�4��Q�.�NB�L��'�i�ҳ����ۃ�\�ٹs�ɓ\�Am2<<�Pý���9O"l����D�-[��m�m�Fs)+΄�����^�C��Zu6RaJ���-�����
v�G�n׮]��Q���B7pR!P>�~��!�1T��<ߺuK��4.��3�l޼���K��+��c�����IB����I�A�C��U�iI�M���i���h"��>u���@(�sӥ*!�l�|W(z�Z)�M	��B4��.�Y8�l��vR���Um!MC���4RV��qU	ca*���7���Q���t"���T�����y�f\�Q�҈����V���R4��G:�S��� �a<$�"B\cw �@�zѦ�0l��N@���Ëɗ�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�������==���p��b"�
��-���54%LWWw��E�1�������ܭ������ �Չ�"�k�N��4%B���)�֢����n�c�Z
C����"� �X�Cmt�dB|Gv�n�����+��7B4`�fQ�.A���h�0�h`#c�.ύ���J��Bh�暄�����]S�A->��I,z�()
vW26�Ey��TV�00v�vC��`8��%ۍ��59JS�8 9�F�� �v����G A�Ҳ��x��W���M���2Dm>HH^`�err�����`S�Ӵ0gv����G�����e����.�.9N�!>c��m��\:Z��s�0-#~�T��h��ݒ0L�H�ӱf�^lZ�E�i�{*L��}�ea����2-M���pL�x�=���td�j���!�Q�����1��0�|i�e�[F| :X��$�L���-�A"U#���Jhe��&����/_V�Ȇ0�UeH���/�ʂ̄A~(�p�0��L����L��)� �ĖE��gAf ���F�1I����,��t1r�!>`��c�#+2�e�^&��{tRY�y�ؽLڅ����e9U+��ae��2
C�v:Lv��\D[�f�&�Yj�٥c��0&b�'�_�]3/sa$g�4�\u'N����ɰC������Cڂ��pa{z5!.A�n���l	3
�p^���)����0 �Hx����0�9v6�����L.��+o[&�q��΄�g;��]�\��:M��PF\�v2�B�A�E00�K�N\��L`�c(qI�p*��S�٩�-v�慎8�R��[�7=:]}�r�yJ&������e�܄���\��d����Y��
�d�ե��3A����������)qI^��!��M�gOqA�R2��{���$_��twwU��]�dE^����0�{c���\��:pNq���t�yJ�c�)��MBZ%a\��0蹐�v-�,ɳK�"�=�t��ICHV䝱�Ԇ��)���0�dE��/�%�6��C�Ln�d�bH�Ԏ��:���#�b�+�X�+aqA;�(r]�]FٵLZ%�)1Bn k��qE^7&2%#DAn��.{�)i{�q����	�{��K\ߚ,�&%[�f��'h�oܸ����b�5�<�܄�����-;yϟ�����!~�s/e���5R��l�y楋��'gf�ks&������~�%(�0ga�\t�!~23/�ESx�#��a|�)ǵ)�03/3�cfΕ�ڴe���dg���҅�(e$lÔ�\G��Lg���K�㢔�3%�4�I�΢�m~o����+���/�0�F���䪔Fπ0�0�Ba<�dg苷�aJ�3���4�W(�g��~�R����VsIׂ����j�䕯}�y��_/|�%�kg~���ُ~l~����k��H�_�5�VvsQ~�mo1^wM��������k�1�����%�b�Ht��w�SG`�z�k��~`|f��/�yn�
jǙs��>���_}����_�|���x�y���9��%*"]���_c����ɿ���3��aLn�����]9�0�(�gg���ް���k�����}��_3?�淪���~�\yCE��_�]r��ξ/a�Qbo|�b��vg�"$pYS^u�s9d�������n����0�gN=g��w���o=a�>��\Ȃ����w�O��o�hôc��df���|�ܹ�\}ƅ�\l�y�M��@���1/<��y�D9���~ȼ��~8�~���g~�;��8m|�E�i�6*%&h_8z�6��ϸ��Ef�ŗ��3���9��3�-~w�_7׾��{t�u�'�e�~�y�{+�� �+���\��M��W���<h=3�=��c������d�Qi�8J��6L�]}�k��,����	�����o���n���G�f�UW��=�������P m���w���,1�^��_}��˩S�3��H�y����Ϧd�>�+���������M����di����p��N���%�a;��?7?���B1^�`����7�?� H	�[��L|����;K�Z�<7a��\�RFGQ���K��3^1A��_8y���8��g̥�_^y� E�}��T�X�z�㗿lΜ��A4{��;|~��_����0��.nJ�#7a�F��U
ݶa�
���X�`N�炚������� C�^=nt$��t�6z��Ϙg����WU�4H�~��S&k��y�qհ#��s�aw[#�l�3Ά)��{�}�y:H�N������0��fƸ���W�:�,r��#�L�a�����>�l��F�����[�ϳ��sI[�0..�6�9ㄚ6����IP���/��˛����޳����ӗ��3�����8��=۱�}[R2{򬨤dn�S&�1�/���ʠ-3?(��~�/\uUx�?�=m����Nzߙ��h� �q-Q�R2GƮ�]}����=�~���L��W�m�dy�ŗ��y<�ۗf#�\�8�x�g����8��![��%��1mI�\�S.#����N�q��41i�{[%U}��%(��U��/�gi��ib�)��N�0��^+�:oy�e��%;�np�}��l�Sϝ2���?�׿�M�� ���7����#��;���
�/8����g�_���;����ߌ���J��'`�"��AKPi����3ƚ|��3��G�+���\|�Ŧ�oR���c�ߜN����K�M���\}����;}�����G��x�:nD��c��'��sN�G�q�5yO��E���jk5��d�u��l�3nR�W͎�?�7��W���������_0��bsE �o|�*�ԓO����*�.�9��,WC�@�p=�O��sҚ=�c?c�^ZoZ+��6v���qM��Epچ1V���ߠK�5W�6
ҩ�}�S�]+V����_4�}��G8��?|:�,��B	3�q�������<�5n�]��4f����w�g�9�0�q�f�F@����φQ��o�3�"M��{��ߘ�Og�c�7ckQ�a��E��a�B���A����z����(O"<=+ë�F=�/�6�O�lC���i��{���C�p����z��(m�0ُ�sa�֔�g��/���8�6�H���0E�eOY�0n��Q����"��Rt$�0��1�����0�0g)���8��P�d�%*���g��\{��10S����Z\oE�\{=2Wc0���%i�)�}祽��S������9k���Mooo����bJ���e�k\Vf==��
YM����!%��>w�O����@�l�q|i��H�<11Y\a�J�a��u��WO�Sa�J�@���YW3�H���._.'a:��}�6aa|e�qef�/�sʜ
c�c�&]
������w�'�6V�������>ʝ���Ka������0��n��g���)�G�ʘ3>~�X�ز 4��R���k17�'��7g�Ԯ���ڕ08��\�q���yl�F�)�Ν��~�}���w1�KJ�G���b/���<��#��:44���;f�5�O�M!��\���$O��f�ìp"Lm:��B�#�+Y����
�a`��,ˉ���٥L�	*�9a����������t6ftt4|��`v���>g:F�A���x����i/�c��^�T���_�~!�!ڎ�R��{k�1�_H�@C_�1{����۳y�L���1��R���k+=�Y�gaƪ��~!�M)���0�,X��SbH���ٛ���̄aw2��f5M&3a������!��`���^k��,ap@vw2����e�e^c�DY�O�Y3Tӽ�*�c�_��"����[�A�V*�����c�0�/Ц�(�ʽ��D�1��߰g/�:�߲0Lǈ�HE.����e-	�t�"�P+iYK�0#E�)���e-	�k�-�1�/�Х�i�n3c2MK�� �%��������A̦��m��B�':�)�������FR����[��)a��pv2)
CCk���FB۶����M	�������L����v�/�0ب�^�@HQ��{�r�ja��h��Y���A%��-��p��H��2Z��c/�����Se44-���!�����*���`Lƾ߿Q�c/y�WX��糽��C�)��|d�n�n��,ܔ0)�tB���6 n��4��]�	)#���ja0���IY�v5%L����s*!��!D�!D�!D�!D�!DA�������ׯ<��!�0����������������������������������������������������������������������������4�ѣG�������4'N���Yoo����1}}}M��%'N��1��(P�A�3{��5������5k��7����l�����ٺu�!��0u�(t���Kb3=}4�[< 
f�{��ڵ����Ea�¤���q㦦D��ъ7����}�v�i�޽c�������uhhȐt(L�ׯ7;w�r��(�������8M����6���_)L}(L.eP�#ڸ�����0:2�YA��0��5R�ИG[��.��1C�����"��ԑ��3tP$wR��m�(�2u�0(�h���H�mc�
kl�P�	iV��5�4Y������;������P�bil޼9x����!�A�ݶ�V�J��!j��n��4���:"i6��CafAAI�Qڱc{�	���C�̍7ޘ��DYԤ� ҿ8a ��P�Y��!Z-D(�{��17�pc��!z�*�\k$�������qQ���t(����$��(d�4,R�uIr���*L�؋�ޘy�e��O�J!K�%�������׫�i#�vG���`�0l�'CaLzAEM�%�7�3��nVP�m��sF&�ƥel�'CaL�0(P.ry�o�g� 7;��<	�cQ��26���xa��M�|.p5�,m�)X�kI°�O���#i�����D���j�cd@�IJ���?������T��r3؉��.�"���D��]��L�0l��O�c#c��W��I�h���/	D�w��Carm���k��h(�i�6� %E(6�k�0932rw�Ϛ�.�m:	�]�N�0l��Bar�ޔ�F
w洱���1������R����(��L�I�.�q$Țtk�sP��شiS�lh�1k���w4��I����&P�Һ}]�)�i�F��=��Ѥ�6�+P�@�u��oL�Mf͐]��^�H�*��
��z�`���ޱ��~�T�z �$	���0�@j�{�Ӑ��!m�����I�d8��q@#i
g+_ԛ
�,iSe���0�����Y�hK���R�%-K�^����0����������:.m�L�7�)LF�V���Y���ې��-$M�Nn�S�hdi٬dA�6���-ՈPiSe:��OaZ@�z��aQV���i�(��yZ_Lǚ$���ŒPE��4I��xU��$P��Y��[���� i!�!�c,����$��E��Y�U�*��F	�i���{�<��iK���۲Z�(P����w��ÒH[`�] -�0�<dK�F���ŷ��\�(P�:hz����j<m�=�ۆ�U����0)���8�z��~�3{�6����;�i�
�@��@��^tq]X��֤vgwR���Ш,.z��%��!���㐛ђ��;��OabhD=aq$m�*4s�X3�M���?�����z���	�#�w4���M�t����0�%덳��ץ���A^����6!�S�f\�z�(�)�'o܊�.A�?m/�Nh�S�Y6nܘ:O��K��\�v[�0����0�20���@�
�.��	�g:&�m�:��OaL��X�dr�I#Ȩ}�]� �tL�Z�i�a����� �L��2�lUn�#3�"R���1���eo�w�0���oim��}��Q!lZ�D��/LZM�.�$����I�~2�̍��F���z�z�>�7U�̍���7ꥈ�L�l�Şv�em�w�0��hi��C:&��'����ha�X%2O|:V��A�'N&����$�)H+��IP�`��N���!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!DA.���K_2/��!E'Sa.��&��c������0�d*����b��k?{�!��[o5��L�yE ��?��/�Ħ�~�J���V����=��[^��[��/�>�������L��`�s�u�;bif�z������"�y��l0��_gO����s����g�
�HFHQ�\����g?�ۉ�3��Sa��`����n2��zs�M��|^�]}��qccc5�-_�,6e�?�����{roo����ٕ{���_�^2��)���w񾲕]�} 6{�~*��]�{�;!c�!�7�ծm�I:N��!A��?��[�@B�3�Y����?�ש�·q��}Q@w��^-��ׯ?o��N��7o��^�́V��5qoG����O׼�֭[����5�罹����eݺ���I���Z�
����/�Ǯ?�~cZg�0Ҹ?�Gw'�g͂ha0D�J^��W�Zȩ��v�-� �]�!]WWw�s�6n��f�����wx߸����'�0�9�\B�f�4Y^�����s�"�G�BNjv�8Y���F�Gt���5��}aAJ��Ie�ɓ'OT?�ZTD��۷i�t���Q	!Q�褽8�0�����q��>�-l���]��0"��{,ڠ�K����0�.��m��s�����D�h4���e˖��qR��m.���_�r�n�X��n�jZ���_�}\�	Q+��� ����K�ӏ=�j�6/}�	s�j�\�@��6��3���P���u�N�v�	��u�ְ# e%�lՍ��?�6[�4�if�
��S(�Rp���eO���55m�E����-��T�+{ll�i�-�?�*xm08�����蓦N�L_*��rz?�((�x\wݢ��#E�4�÷�_�.d�m�q�_FG���F���̍	��dL'k��O��� fGoR��A���C��'I�0�챒F>c;҆�`�WSB����Ԟ=��;���ς�
I��{aP��9��y����R� Ht�u�7Ҁ߼�2��!C�=�HWo�z"e���{qĽ?��Dà��o�{���0��6{]��C����ٵkg����V@Ã�K)�I�tH[��G@�ÂJ��� ���-�fH��B�>h�t��5�uJ/�4h�'���(!!YAaQ@aQ�S�9�F�ʳ�0}�sҩ0%#D�!D�!D�!D�Z��Ţ�����k2�C-�4�)�,�b��Z�d�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�aN�8a&''����ݦ�����t�@��������W������1˗/)��G���sz��H%dW@��]������˗�?+�f׮]f�޽�cL�w��x��A���A�að���1�����hU�$*��x�{�@�5k����`)�g�����?�eg��,��?v�;~<�w�>($x �l�|W���@�322��9��۸qS�(��,�0i����ҥ�1�/6�-
�.�}���92e�LM�Ç����9j�+���c�vS��SOT8K�,	����!�*�c�*���c��቉����糨�N���֭�I.��2s�m�;���������W)��շ�������}�@���g]wݢ�"o/tو;��-+�T>K�
(����������5�8�����,R;�P� 7^�~}���nݺ�fepQ@��H�v���{���j�A틋�g�C�,�YD�KvǈT@�EDh���O�;��B��������t�F\XԂ6��D��c�a�֬0�{߿d[(̽��Wm�@�o��P9	T>;w�y��P+�ā���;���J3z��Ո��oŊ��֭[��А�B���qP[�WjFH��n�͂�x���a��Q.����V��sz߽�dr���g����_��	 �Ie�4���m_ذ���3�e���
O:j.m�2Y]|&|����"U��,8���n�ϼX���f�{�cn�v���@����Z�^X�qQF^G�3��B�?[�U�V�C��M��jx��\e�z�{�}��tuu����#�
#��B\-Q F4�$��Qi���Zuki|PT��Ϗ��k׮��!uo����[aP�H�$�KΎ�D���E���J��������r����-���zo�~��L�4�?~���� ��DI��hR�p���a7r(G�����Tj_ϊJ���jG ��1���M��X* �����Jp�}����h(|"DZ�]|pw���p�^���荓T����R1{P2�j'2������}���Ɩ%�l :�[�6��p���Oz=+��LjEJ<|��b�bHU]w�*HdR	�<l߾���W� �؍R����e�"^w!���2# i������b�b���v!�xǝ�Gy��$_��W�l�6Z}����O�&h�q�9b���,	?��\����\`�c	��1���^[	�e��������&v�Y9;]W�D���T�v��w2�8�1;��ܲre�|��ز�c]���b��n�&ȁ�G^�:��
}�!�ΩLJ-B���m����1/f x#�݋�����q�D
	���NQ��[��or�#:OP�d�(�A�����$U��ؤ�w�R[��,q��Ť�(�\`�	�O;���2X��H��<x0��Q
#��9$J�ٮ`f�#�i�/��Wt��(�����i�.���0�A�]�D�ζ� Fԫ_1�Mu� P�5�Y /�GF�}��^c�"'���� Pca����T
&��~�V�s*�BD��()&�d�셊H��vo�o(���]چ8��T�_�,j��(�&w���GeL�h"�W,lh�6~�(,=i�T>Z(�������2 ��apN�=��a��iM��e�ymד2}�}aQ�q�"E��7�jA��X��j�F���#7~ͭ��$�q����/�^イ6�˩�@z�@;sn�pU�S.�,�(.}��H����3��k;�mw��&�gl��EŅjά���+��Fv���Lk[�F�*��w�J�{O�^:ہPJ+H�2�'e�L��l�����*�XM=�$}��,R���R�e�&kf���Voo��$�P��(�}}��}����Y�����������dQ�h��4̈�N�iY��2�yE�)�}]Lc���2��$�����RB��)`��v�0v��>AY��(..R��2�'���pO�^"�5ӆ�6��z�@�E���RBy?,;+����v�0�"A��Ǜi�ed9)�>�v�DVsN��2it�	�H��^ ;%L{?�3�]�pҲ^)i�%��vtl��4�h�ɗSG�8�[ t]����R����Ik�ǽ���m>��^�';�Y�IQ&n��Y�P���+63���]bw7��@2ݦQ����rn��R�A��Z��(�դL�R2;��=���r�:0;�3N���}Г���'D���|���b\��j��ko�v��;�TҲ}��´�~��@���d�X�xqux�r?�I�F�kR敹TL�U�Q��fw�,��&O�Aa�m�耧-������7� �?"K�ZO,n���I��e��5��'�i�ǃ):8>��hg�-�a){z���J4,S����E�I�oeR�=����b@䕕c\.�%�4vti�xQ�'G�2(ԭ�G�(�Y�����b-��n�"�����`�%A�����(��+2��^8)��r�hdCM���v�i�9ǃ�JQ&�{W�������u@�ٲek��
�l*�}�e4�2!3�5��c��tU�h%�9t��7d�R@z�ܳ����D�]��j\�hQ��T��}����Y��d��`eF_�.Q����j_�� "�T@8������Ka N����nf�L�fY���%K����hw-�|�yT@8Ni���1P�K' �o* o����N��GRz�P�g)M�\��I�QYP}X�p��M!����~��Ѻ�ݲ�p˾&�`&�[��Y�n��X�}u69N�8���`dD�Ǵ!9��4G�iK�K*A;�`�w��;�y-�Jp�1��f���A�ҝA�`w�qu{�nI��&\�mj*׍�Q�6�,�W@��AZ��iZ]8.�Ȫ'H�EnÅݲeK�d����rL���2E� �m��y���B ��ԑp�b�Ռ��Z�rK�ڦ{�D�w�Y)�g�` ���)C��4�6m�nb%i'mo�|&�
i[P�Qǁ��/Ӊ�Qa�\dL�Ao�DԎ���[Xx[;0g�X���0�2���ر���v�H����`��w��D�me�1��`\�-
(�9-�0jx�p�^�[���#����/�⊚��lp1���h����Vq
>ϧ�LYS <Rm��E�}���M��Ѐ?.�tb"��s�U�H]Ha �|�v�i����Ǭ�_-����0U(j[E�D���Y�s��;7!"G#k1�(hw��VA�A#�Ta��!�En�B���8�k���-����ϕ�����L�d*�4+[�0G�N�,v]�#�&x��D�V�8�h0� [��\�{�D�u�sY�i�̔)B�F�(�M/2�Ǯ�{#�N9ץ���cy�UJ��������������α�������[L(ĭЄD)�0Qp�?ne�m�pR\J-��X�n=�ɌR�j��N��dKi�A*&9`	!�����Y��V���ު4HͰ�YQ'�RZa z�$�H � �PZa�ZLt�:t <��!CH��VYZ	��ɲ�X��˼�%qKi�d�kD�����i�����2�bF�ٸqc��!Z:B�)2+VTVlĸ�Y΅����rD�f:ı��c�X��i:�-��l�D򣣄9�`��3����  ���'<� ��pÍ�s���@�#���^b`lf�~
C�ӑ� 4����V7J�$��c�A�e˖�fժU���2�ԣc��݃�W#$���	�����' ���zt�0����@H/@��];kv[&$�R	��bY!F;���@����t���]}��q��G��!�5��������������jap+/o�%�
#!
(!
(!
(!
(!
���9�����!�
#!
(!
(!
(!
�?2�p7�O��    IEND�B`�PK
     mdZ-s;�.@  .@  /   images/3e0a96b2-ef1c-4fb2-8b57-d71cbe1f3744.png�PNG

   IHDR   d  �   {㓊   	pHYs  �  ��+   tEXtSoftware Adobe ImageReadyq�e<  ?�IDATx��]|T�����%Xpww�P��k�-VhKi�����-E��+$� �5	��~s�p$'�rw����~	ɻ�}�������8�����8:J^Ԁ��(�g�A\�ŕM\1$��8&�{�F�gq�$��$��� �u�ƨ�����'4BU8&�iBBb��ŅZ�jEY�f��)�l	��>|��\����D3�J��&LO%K�$	��o�~��D?7(�0K���I�~��5,y���Bc� $!*�$De�����A�2؝��w�ҙ3g�L�Ҕ/_��~F��B�<�`��$���رC,��R�:ui׮���!00�Z�jM�ƍ�#F�D2׀F�Hǎ�y��ӠA���h(uj7rr��S��Dttyxd�-Z����e�R<�@�����ݻm۶�F�M���I�0�N��P�4v��ׯ���P�֭I"1�MxGD`��f=��w�Q�X��s�|�H6B�=vpp�3�S�z��_fҀ�I�m$�yS�n]��>}:ϒ̙3�Y���7G�E[��C3g�fojI�R��ܹs?����K�#2���QQQ�h@��[��W�rw��NH�ҥiȐ!�+�?}�4�=;U�X�$��;!ժU��J�*E�'�7��[e�����A�2$!AAAt��-�q�:=~����r�|��S���(}�����������u��={�?C�r���k'Dt�v%d����h�":r�(ݾ}K����+����p�"Ըqcvϗ+W�R�/_��+WҶm�����P^��}<�Ҧ��v6�.]�P���������K�}7R��Vʘ1#ըQ����M9rx�������/�ӝ;w� �?�����eǏGy�����駟~�A��Ǿ��}x-C�t��)�+�ءC{��`!M�4�~��W�޽;���<sl��x�b<x��LM�4�lٲ�v-�u+vU�X�>jӚnݺM�6o�e˖��ݻ鯿���ў8t���ً�h���}���@�������=��瘹9s�	����;w.mݺ����O���6m�M	��p�СT�l91CFq�I��Q�b
����t�K/���3}�Q[&�]�vd�_��:w�L��Yi��S�*�y�`�����6��_��ݺ�Lz���ԩ�[�u�֡�&N�-ZВ%��cǎ6k�����f2jT��b'���P�����$��m�<y*��f͚�W_⫫�A�DgU![��Ǉ�v��bq����5<��v����Ey��Ϟ;����͍�T����7��7ԣGOV�5kִI�lB�8��V�Ǐz"��Y��ɉ�h��ԪeKjժ%?~�BBCQ�Կ� :x��ͬ��O�
�eȐ��M�,:2W"2 ���W�R���Y^��G��c�39r�)S&Q���g���8�3g���6!dܸ����+���o�������2uծ]�ڶ�����;�:d0=|����bp��Ѷh&�R����/?�,�����o�!�o� O��q�7��:�k1:����K#�h<do�M����m����=Mk֬�N�GŽ����[4����j�P�<u�څE	�����K<�p��T�Vm�3g��)��0���ݣ߅���]�f�dDFFҍ�שv�b`<DD
1g��}�)իWcd޼yb��K�i)�&dݺ�<�?���[#�p����S���^z��.��q�G�^V�'B�9p m߾�MMk�a���������o �ѣ�!Hə#�EG(��iӦI4�a1�Y�v�H{���0�X�N��E�����F��Ȝ<e�0%�%�(-Q��P��h�xQk	A;===��x�1`�B��+t���?+Z���xVQ��bE��[�rC�YS�d�6%�@F،?{??��эɘo� ��A��^�'���ׯ)M�4Ij'b�ѱ�*Ud��9w��5*R�0�����~�ڵ5:��N��x��l��M�%KJ*�"�ɓ@�(�lM�֑1m�1�ܙ�'N
2���G�B�8z>888Ʉ�8�s�v^��a���`uqq�6�~��ܽ{�X�<H9B�={*�leʔ�h�dl<��~A��>M?�g�Xɛ"p#�Ӛ��}$BȜ%3�c@[=zD�K�;w����Ư?�msww�؁/^�5����c�/�����5~�k��3e�Q�
�M��x�MB��<�#  ���,����Z�"S�<!:}�!ka!X`���b�z��d�ΝG�wS�xf��݋jժ����b��CёT@o���%戽*�X�hz���D�9c��XXf8Z�u�5���`�\�Jߔ�}?g�\z)�ߍ����3f�WJ:�<�7�d�LI"^���/f�)@�ݺu��6i",� �(���J^H
�2`Z��K��;}�+wLy�<�#fF��KB���ʕ�C #b�S�No����T��Bw��xV�N� �"��m��G���֣���sXW�߅(���öm�Ұa_�YY^�G o��B4r���D ����1�ϨM�.��6m��gϲ#0����Q�]�Qۏ̊+|�.�'ξX�	�Y�ɓ'ӊ��lٲ��Jnܸqcً�20�^�x��*S�,թS��f�����jժ<���b^��L~!fw�B7����byx�`稵���-XOp �3�9f�h�ǧN�n1 ����K��7h���lvZ��A	(��V��0�6��C蹦͚�>H�l�L��]]]韭[Y�M�8�j`o�A��8�$�C�֮fk&�d�����K���獟O>��l��7�ԩ�ٓ'&�}u��Lٳ��]�ٺ2��0��+�g$[�&����v&�8O�<���©k�.T�F^,)^3d�=F��r4k�,�%@���Au�֣aÿ�ӧ�k����X�A�\�F�z�4�?@���aÿa}�g�M��&m�َ!�x~A
Bh�4m̾ 4�ޘ,��b|��%-�k)�W��dt��Q�X1Z�r��}�����i���5f� *U�$o���Ĳ��Oډ�ALaf��6lX�֕�`�=ulm�ݻ�w�0�7o�"�VG��eX#�A�Gu
;�ǎ#o�t�Z �oߞfϞ͇D��C;���K��=���C:v��.\�@y��a��ډ�=8t�f�-� lu���ݻx���Ů��e*(�z,$�I��3ׄ��Ɉ}�ҥ�RVЧ�v�� �I����a=�fͦ'O��f�c���]B�`V?~��^�Ц�7�ŝ�8t��Ĕ>����<t��޽�ܹSL��X8�?���}�5klhٲ%կ_�]$�	�=��)�D�M����{t��eڱc'��	��7�B�qn{�^�F.b��U6.L��u:/���h��q!�X}�P�\6	`P�d�X&��7' �p�R~xJ�I�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2$��֜�0C��D�����h:q��S*I(#a	4�>af��9�А��,a_*ӑ�'(��䚚j�Gy�􎱔�Ցһ8PZ�W�=�z��| y��ء�	���
�����X
���h�>D�=�g���݉HIL����#�.K�K��,α���I\��Q|�$��n�h��]�_�.���o���M��aA�:<�^��Ux4��K|Itb�J��0jeEGEPTd8E�GG:ES�PB����E�Nv D�~"	�"B)fID��CqE��#�1v�O��*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2HBTI�������g�}�u9a��ط���/6��ߨ�!�N��������5P V�nTd��Q��S���Q��g'��t�H������rvr$�
�#1_���1���X���b� �F�8* �yt4QDX8����Ӡ z��=z���<���'�48X|}L���'�S4�+z����L�lL Hrtr"w�l���FY�d�L���5[v�r��K3f"WWJ��J��vhI2�y��HBD�9h4\3��IC����WH��ҍk�����tC����`
W��h�����f�qpp$W�T�*eɚ�����*X�.��W�(M�4�N=�I��̢d�Iv#D�#�فЧ/�?�;�oҹ�'��9q����01�o�u�&��m"FXX(����Ā��;�TLH*Y����Q�
�(O����Ip)�e,d/1gӷ�Ғ�����t��m:s�8?z���{�n�w]��U���x���;�tz����<f1y���,u��<��W�JUkԦ
��R���)uj�7�ǆ����Q,䵳E�^���%:rp/=��Ο��Œ�΀�0�!)6&���YB�/��k���Y裲�+R����zͺT�H1J��-��(�gN�Aw2	B��Eҵ+~�s�f:�{;�?w�+�h���)ou`of��6:��`��{�rK��ʔ�H���FM[R�B����L��LNR���ظ:��
�đ?�G�����	�C����pHV��`��y���
q|��_���"�iˏ�^���3WN%�a�����x���dX&���t��c�o�:ڽ}3ݹ�_\C�_L��I�����K�'[��ФEjҺ�*�]Hd��˼�h��XJ�$��K:tt��Mg�VJ��C$����@]4g&-�c>U�V���J%�6 �ԙ�!*\kK��utv���t`�:�cݺ���%���,b}��`�RT�u*U�9gέ]�@��h�������t'�?"���W.Ѝi�R��S�V�)��S��1\X2<�����K"l]?=�M�L ''geuupPo|J�Zk�X[��S]�[��x���Q��R�r��iӊUqjJ�.�X�8�W]�zxx�{\�r1���w�~��ի�A/_��ׯq�����ה#HVBu~�t�c�f�B�s����gAʓ'eɒ%�����3!nnn�M8)Aȋ/9�(D,Z�>}Jw�ޥ7nP@�5�DO�<�gϞ%x��#�\�+!�������E���%KR���(�����.�j����+_�Yƀ�Ȥܾ}�Μ9C�Ν��ׯ���'~�w��h�g[���he����#�+F�+W�:uꐗW1ʙ3'�x%�%T��q__��Q�R,�L���������,��Tb��
\ho�ƍ���;�I ���Ct��a���癤��}sV�/���]�\�rT�fjР�*U����g�����Ǐ����G���{����w��}�� ���#����9�
DFF��U��VD�&M&G��E|MKٳg�#�ʕ[��\�-[vq�����l�K�OOO�@ܭ[��t��A��������$[�$�?�@ܴiS*]�T|G� 1 9��v�j����(���<�3�7ns%�$ 3��Rb��M���Vƌ�@�LD�bE�P�B���k�Y��jժ�___ڱc�޽�N�>MϟkuPRg�r�b,^R��_�j�ZԦMjݺ7\X8����ʕ�,�/^�?y@��3��a�����$#�\���>��*��2eJ�[\|_�ʖ-�׈#x�m޼����o:v�X�̱��=�/� _۶mK�:u�W�\!ooo:y�$�:�/ݼy��P��F�}����$��:w�,-[��j���RŊ�J��L̗_~�����
Z�n]�|�8�B�H3^�;�B��mݺ5�P�j��>>�h�ܹt���T�4}�b����!� �ѣ�|;�C�g�x��FK�:��^�zԫWO2d0?~�V�\ɳG�W�-�D�h� ʛ7�k׎��oN�8I'��: 88H���!�W�k���ߏ�ϟO�2e&~AP]j߾=u�֍�m���@�	���n_8o޼T�Z5^�ݹsWL����ߘ���n�
	;f.�+��*U�r>��9r�%���'z��ŕ;�СC�z�j��wA���A�]�~�/��#��\\\ؓ�#%��a�C\�R�����P�=|��C?�!�ِ�ε���D�B�2HBTI�� 	Q$!*�$De������(!��s��}uBZ�7�V�p�dʔ�␛���ۨ�)��<T�D� 6 a�$��ڵk������# ���c����S���7n,�o߁�Z
��?�K�|�	{y�:u�oF�HR�(��ٳ{��G�$~��w�8���8�6m����pJ���7t��I"m�/�6��D�`Zb�_�Я_?钷!����۷ؠB\�Y��Q��?�!b��ٳT�B���,YBE�᨝u��&[E�s��"�-I�m�Р}��Ӱa_	�e88� !��ݠA}Z�z�92Q<���@�#��:t�@���7x��ub`ԣG��jժEI�tŊT�JU*]����Q�722�5j$|ڲ�I��@P���g觟~���@�=��«#�B&��hp�����LB�-L�gb	��B��A�R�'6�����hS0�Ӏ��uȾ}�$!I�X> ��\��YB
.�G�����_���8~��J�7oa�^����Z�jӟ��Q���������)^��콊͚ܰ5�3�ӹs�$!3�ĉT�R%ʐ!������pB�ଈ�r�$"�G��A����I!,f�9��FEP
�*C���(�9�^����L>��sʰw�^6u��+)&+�q���	*I�2��/�P�p���:ń.\��8q��6mB�q��-�L?�����(&�qv=%��ƍ����)]�PL�#�T9z�(��0�;DB$Ȝ9'P
��A*V�@k׮�����~��i���+U),"3S�Ν;�3�~,R�y�T
��;�.\�H6$	�x��1�i�Ʋ��E���}\�|�$L)�?~D^^��W���d�)׮]'	Ӏ� �,��1����~HH��Dd"����,�ń,X����'	1�۷��73f[�	�O&88�	���0��3f̠�宏$����)a��u����ń �$�l6��5�Iq�ZL\&PV8pb�m��7Q'4dn;^^=���bBt���<1OJ�eVFm��|�7�P��YPڽ�lY#���і�bB㋀���FdL���N��7e礚
8Z
g���7���{������#�
IIqe1!�h�����qr������!\l�ݥC�Q���E�df�����w,�6�})�@�G
qO+�ĕK}7�,^8,"B���콺B NN�d),&���-u\*X�ЈFE;����'�	� �����������(g葰�pR��:i�yw�x
s��}H%9ոr�%�@g��Q�:qE�����tkȖ�c��G�@�� y�x�G%3D˄�с+@kMe�2[X6ptu�'E���i���u��#f��J	�&Pp�r�Y�j�&?K���S��M���C���}&�,��B<߽tir/S�\�wK������Yzv�F��u�S!�DV�[�A�g1CBŢ��ԛ�.I��J��磨�n
�cnDBt::�g����t)zt�=�p��g�,@۷�;>����7"6�
�.����`��p�螋�����T��#GE��}X\=uS/ι���FDF�&����X����\�JRfAƹ����7��o�^�\�Q���������r�("4�\�:�	��{D���UN�жp�����mRY�$YY�Af~\��1Y �����H1����~����](k��t�?ݾrU��7f)2I���LE�Q�R���Ejצ��7)[���6�<}F�v����h��6\���
�ϓ�'�bB�	��+�V:�ݤ
��1Q��3D;��ߏ����F�3��s�@G�@d���P̌�ŊQ�X;���N�D������LӦ��j:�i��F��h��f	25X
�	�'�� R����aq	������?'!��ԢW¢��Mx��%/� G����� tJ��;��LW(K�\)~mr��3DW���;#uHAz*Ka1!�z��y{R	@HXl���#1��{tp��>T\�&�gZ��H�LrME��s	��(L�Tnb�M�#"���bvG�8VXu�QBDƊ�iu������
�']����-�3J��z͗�h���Xmݚ�X����+"+�3�&;@t��

�L�����o��:N�Ly�ғ�O�uxE����1ڿAڿǄĚ�h��,*�]�v��H\�`1!�i�+���t�:/kVdň{R���h/���A�"�:���sT�I��U���]"�n-Q�e̞��=��\\]㞭�hf�n�ĘY��-Ju����E�K"O,&ǳPgDi�5DV8��X�3$�S#1fpL���%E�F
��w��R��@�e����{�����=^��̗�r��q���)����E1�� :,F�����	�k����#,��A�"�` ە�7�c��4�B�C��I� �8B�߼u�^@΋1���rL����y��%���s�ݾ{���,EK��>��o����"#=��9!�������g���Ř�kKE��_�|a�b��������+�/����c��&��mڰ>.����:�i�-9����p�������>,�l�)f�A����ַ%��s��z�kL�����ܹ��W\��R$���N�$+'����XR�v��	��ELsGh��u0p�F���z�X�*pq`��|G'K�̼4�@K`!��(�ӬY3şa���]o�aӂk��(0�P\?�����)�i���Cf�!����� ���s�%�����%�+������b1�o2�w�gI�L���鯿���!BV�9{�#�1-%@8LΜ��S�NB+�CQ+P��a�R�xU�"(�:e�d.�j'B�1J���q׮���ɑbb�]F����䘷�*ų�f������8��bB��Eh�-T����'O���U�һ�`צW����F8�ܳgE�QL��q�W��J?�E��~���������s�G�Q�X�!��(!e�����VLȥK��.*F+�0�׹��>��Ϗƍo��B��)S��订��	9x��h��,D� � �������-���ș2mF:���G(��B&Z��!���=�ݻOтZ!�������ߏ$	� ��˫W�V�G���aa�,%,G��Mh	�u�Ș����������� �>,M�����>L5j԰�D���Y�[�n��ݻ���,!Ȉv��-�:u
I$	BM�ݻwQpp�Ɉ����RjT�^�$��v���_-��45i���}F	����;vr�E��%��ʕ+���"9 Ę7�(!p��9s��
��=IX�ȅ�ڹsǵYTXR��@+W��L�2S���I�zt�ؑ֯_�����?4H؃3�\�4iB�s�&	�Q�^]���^���i�ABi��7oޤY�f��m �o�-i���F�Gqe��G,�����ЩSGZ�x1���HD��ϟ?�`��{4��oÚ,ʔ)#���K�»�%KV���N��!���{R)T�j))	t�Q�=�3!�`�����E����n��E�����sĈw{�Б�0X������f)[p��]����U��YY�&M"�=��ȋ�3�~������2:C��o=b��Ya���el�`qbD�:���YS�Z�0@�ҥK���#�cDCyu���l�=��������0Zk	�!*ʰ�Qu"��ظڭggJ�P��y���{�y�|r�P�$�ea@O�P��[LHlxI��D|�_�h���3�/K�2HBTI�� 	Q$!*�$De�����A�2���B0�����ӯƀ����v��Ln��E'N������|H��踬Y�Rɒ%�]���n�:N ��o�~|�����|T����&����E0���Dg�����4g�\j޼9M�6��Ɣ����v횷~���]�vU\|>9�
BP���҅��b��م��!.,,,����X�u�?t��yڴi#�Q��+W�W������\�xQ�|�	VR��~�>{��.]����B�
����,���Z��3w���$���5�!!��Ι/_^:y�!cɒ�$!�X�j��=V��;i�D!�F�u�.���Y��?@��(f�9&)��	�����'�}���h��C��0%T-����x{{�W�5j��l���ۗO.]��Æ�i�С\��0׮]��ڬYS>|y��5�]�v���)J���gH�7�OeyT0��/_�$^�z��1�,���q���ըQ#V�u��fB <x�*�{����f팥ԩ��IYb��ٳq�+RV` ��1B֬Y�	1��ib�}���x�^� ,T-�=E	)Q��;wV��L���� ���d�f)u0:�A6��[��ϡ[�fMNr��E�?�_|��`��7.K�}���PW��3V�d׮]�:`q�x�v������[�h΄���wC�_�ݲ�:�F�+uK��S��+H�wp��X��5k�A�2eʳ����g͚�A�Z�F(�����N�ӫC�~EϞA�h�H�g��3x/�-���W�	KiW�P��>>G���W��}p�*�w�8a�8�?n�M_|�ѕ�ƍ�C��V�Z&�>�O>��	�3��8Ȣ,��N�2���+WƓQ�~;v���!���B�X�R�*�*U��͛7���ǳ��{����� �\$0_ud`q�4ƒq?~����1�+�ڵk��)w�;�mR�&�p�n�9i�2*��{Sg�̑�@�`��M�s��q�hX���)��UK��]�vc������kЪU+M�]y��	m۶-�ڳ��ƍ3z��F�ƌ�В�s�(M�kK��$L���:�:2Z�nMK�,1[&k��7��+y�ლ.4�7u��+2x#%�X$7TG�o��F_��}@����>�O��:ӨQk�h��J��qߛ�]��`��a���2i��d7:租&�7�|���/_�	  �3{��Im۶�lԦ��D�S�N�cǎ���o��g����P!:2�g�c(C��4g����ʓ0#Ջϙ�T�����?��+*���gϘ��Y�>��� �?��ȓ'/;�,ɳ��ʆ�{<�]P���5�#GN�f �^���ɩ�S�T��[lJiϴ,�)F��3�BT�?�g��8���4h@˗/�� �[r+�'d̘1�T}�b.��0J��k-#�����sҦM��Nl��c& �+V��pA�N�h�����.���}�H���+\� �V��\%�P�^=*R�(]��R�^�$�rOQB�u�J���'�ٳۢg�⏷w>�Ӊ+d Mj"��6mZs��<(wÆ%�rO1B`��:�/oM��W�^q�n�
.��Z�6Ĉ͘�s|��ՋP�t��;,��B
���[�:\��ׂ�U��A�JŌ�*�S��=�^�я?N 59'�HL	���%�6$!*�$De�����A�2HBTI�� 	Q�@�L`fO(#$. �!��+�W./�����7����$��"BR5jD�W�"��#�^��\*U$�Z�݇���}� c߾}�Iչs*Uʲ�&j�"B\��#�jU)���S��/(ݗ���G�c�l�2���-a��q,�#��	�"#���!�r�Õ�m\C�X�j����d���{O�FtJ��~���=)
�b�=���&Ы�ȹ�9�OOi[�&���xK5m�4t��mފ�z5����9�Bt���G���Ç8��ѣ���;X�!Czʚ՝�����9<<��W_}���ABu5p��\�oذ�����i���{����@�����g@��P@�T�b��V���~�V���e^�'=5��}|�e�<��{�(6,�\ �\��f Β� �̙3i޼yԽ{�Dl�6oނ�=�����ׯsڌ��~����K�ʕ�R��Ǐ�|'gΜ� 8��S� o��tT����y   !��Az9ciR.��io1���r��i���=!�s��e�7�n�B!k�Q��e�y����Bՙ8�0P�� J�a�1�8|��p޻!���A��ܹs83��e?>a�T��=G��9�G�l���ĉ���-ƚ�lD��[�vD�^�v%�x�b$u��)���(����u�gH�"E(X��c�ե����q�F�㮈���Q�5cƌ�?6��(�<PHt�m�V�%:r��o8�Q�Ç��ѣy� ѡ��ڡe��$���a�c���b�G	�U^yj����ŋ9��˗��Qc�i�3Z��abԎ��ݯ__��}��	�G�+��b *���1U��W�jժ��ݻ9,G����у 1�x>���¢jŊ�2��3�h�b����,�aS�Iv:q�x��1zq�J
������ � 芄7:�g����������Ʈ];��Brc'q�5�ݗ�fq�U�F}��a��>�6m����Q:2 C�>�Ϡ�p�/0Q�����o���C���5Ya�4�� ���<"�z��0�[�55 �k*C'�����@�;	{Bc���Q� fcE�%�,CC��`C���-[�+c�A$l�rtm�u����d�4x�����F���ޕP�#�-�2HBTI�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De����N�p|ge�jb؝��/_r^�����G�q�|d%͖͝���a�:u(cƌ�R�I/TF8y�$8E;q ��)��W���${�n���2��-X���v�O��
�����f�ʧh�hٲ�4k�,ʗ/?�@5]y�� �d#�ĪU���/ڙ+gN��8`z�ߟ���GS�N!�|,ǻA�=`B0����џ�͍�L^Ŋ�k*>Ά�c�?G"�/҆��AѥK���MM�6%{Ჿ�>�F�%f�+jР>���[�iF�9f0�6b����;i����F�;%5��1؜�s�۷�x�4��/y4�#E�J�.%�UX��8��9sf&�V͚,.f���hђ�� N��H�e˸z���Q11Xte���_{���,�VV�(��ƨ�6W�|d��y���qn[���lڴ�>��3W&�|@�nݢ&���I��`#N��^����Ƒ�q�'РA��� �[g�{��� ���C�{��c�螮���W1�1}-Y�����1c���R�r���r}�H��4u�$.ō��k}����B�"AL����M\Jw��c����èQ��A�u�ֵU3iܸ�L��!C�k�.L�%�(uIp�>�Ř���1��MAg���'�dX&!!��X̌���*�w0�8�3g5iҘG�����$�����ԻO?<xת�E�`T�A}�V�Z��܉;7)g(u�a;�gܺy��@������	!۶m��,C��Ž� �|T�ӓv��I�:v�U:rԇ�5m³��9s�AB����{	����D��pw���TWU���a����Q�c��5��=NnB�̙C�=XG藨C��_f�J͛5�Y�4����1�!k�Q��U����O�����BI���4�1r��,Gb�HB�CM9r�.]:��?��)����V�r@(]ԺUK^_�0�~���&O�ܜ	%�ׯ���jԨ_��@��V-[�T!|}�sꦤb=gr���麀uL�����8˲Y��\_̌�q�'����ϸ���Bf/\��5jȲv��T�J����ʔ-#LOW!�'���#��PaQa�q��)�
�j�^y(P�ʔ.�bR�3��A���Ãʕ+˙�@�5�>�&eﰐB�fC���h�"��=�ݻ���Fa_�t��%�N��es��%�*��:7�������А	��Y[��i�S���G��B\�|9�[��*&L�%��O��M�#&� C�O3��o#W�HL*�&/��XٚMM�4�5LH�F��6W��C~���w�
���j��t��9J�&�贼< J/N�j���ă��8}���?�ݷ��	�d�|"&�S�x9:��5w���w��(E	�´e�Y���A¡Ç��[f($��YP��x�BX-�g`%��t��΋��ժV��\�.���BY�L�E�U�re0s�n�3�2�rݺ�1SF�,X�ʔ)�3I�����{����jB��7e��v�V�J�z��U�V�aEn�<��u�MI5)u��a�a=]y�Q}��U������u��nڰAj�Q�w!� ���5kų�)��1��!���Aw�|`I�Մ`�?S/�e��,A�_(�F���h��3gN�:{'x�����d��t
�0a�#�l̊���(����ؑxM̠?�\�톨�^)S��k�N,S1m�m>ǎ��3F?�WR`5!eʔeg^ &�1`� �k���i��-TU�X&�v�>}z$�/H�+'��E'�m�BT%0h�>A0 �{����	�Hw��$�)Q����v�<�:u�;�ˢ�XMHYa���Ģ�a�&���F�?��C�N���4a�A����9v\,S	����P�Xܽ{��l�j��+k Vfp�ڵ��h�+W�O�/�,ĳ
���x�&M�Z�j5!�έ[��E���SҞF�u�Y��Ӷ�;h�Q�ѳ����>yK!r1Gam����̊)lU;۷�@��2�W�={�P\���{�g��~+��=�wv�"������տvG/]�\t�踺�Ɲ�XD���b��F�9c�v��;a^�^����_|au�U������+����OJ>}��F�sbq�D,xkȇo)lB,�����ɓ٬��J߅��K��o��HcF��\p��UnK!��T�(�J�k�n���Z`��7VtZm�5�7?~�Ɂc:_���~g���ߓ-`���t��j?�
�J��,��0fIժUh�[X�_�`�"��@
Տ=�}M�&M�Uِ@�elx�޽z�,���20;
1�}�v~&6�l�ЪU+�>iC��Q��g7;�H(�"�+�#H7��7_�R�.�����^���j�%!���֭��F��ϰє�դ�SЁ�^�M��[�w�΄�
6��`˖�Աc'A�h^o���-�ַ`�TQf+w��m۶��c�qrH/aN"�R��ST@�����ѥ����/�`��v���S�cp�w��y__���9t��i�@@�-��l�7o^ڽ{��������l�ԫW����7^.T����5�B^��c�_�~\֌���7o.�ֿ�n��݇jլAͅ�՗�=9�83�i<���k�u�6@�,aQ�����m�K:�Uz���S{�����斚Wƺ� u?�E4i҄f��3[C������ΝK���BD$���Enž���)@M��8	4/��強%������q�t8��#�u����ਃK;o),�&L�@Ç�ӧO�ѣ>\���1�K�.C�J�U�X^���d�텘�J�Z����Y��2HBTI�� 	Q$!*C��e����?��@k֬�J;�\�Б,��×/_Ƈc�.���!��%�Ē�d"9,�֬YÑ�����WB�5�d"D�n��.�o�����H�dS��9�vA |�
��HB�5���r��|(2Yނ
�
�i�h��p�>�V�XA�}7�v��A�Gaz[!Y�!�%��b[�yN�#��Rdaح[7>�>v�8�嗟����"=�2e�d�W�>�\��*�j-Rlhb���qG$�H�u��0�������{#��]��YQHB����A�t��]����&�H&BL���G�ϻ
iި��A�2HBTI��`�����I%LØ�(�OArH>V�@~�G�%,�3�pUCHDn����cǐ�}���=��'�T�,1t����D��!���p��ɇx��OΝ�F)
&$:��������h�\l    IEND�B`�PK
     mdZ�.��� � /   images/ac27922a-fd15-40ea-8551-3be3f9cd5316.png�PNG

   IHDR  v  �   K,�  0�iCCPICC Profile  x��||eE���6�ѫt���H�w� �l6,�d7$٥X��lv7��l��.  ]�4\�R��4������I���̝�x����/�}�Mδ3�|Ϲ�^��3��¹��I2o����I�{�wu�W���o��$��,Z���Ց�'�~��ǒz}���J��~֛9�h I�W,��K����/$�~♱���%z�ѳ=zeǓӛ:���V�)�V[:0}��$���^�(IV�O����y����\�w�@w漙3�d5H$�=wɼ!��И���>'I���xv���=�:c�\�GЭ�m���������:���L�^e)cͩlf���:��������C�6MT2M��4�9�5�kʴ\����Ӕкdx��v��{Y��"��t%,I��ݓ*��,iƫĿgZM:��d"^�If'��|�'C�@�m҄v��5azHf&�k�%5�R��BP���q-`�%g)F��I���ןŃ,����͞���M����5��$$�͹�^����OĶ��r?��μ0Iڶ ㎱�|�$W<�$�\���$Yc�$��m �ۜ¯�:����������\�\�ܖ<�<���|аj��a��7��pm�C��ZcT6j�CF]6�ѕ�;��o���ό�pL���<1v��3�^1����#�=���+�_�+o��Ze�*�Y�
��Xyՙ��q����Z�e�[��k\��Vk���Zk}o�O����9x�q랾�V�ݼ~���lp�6��U�m����xݍ��d�M�lz�f37�p��8����䋷5���-W������j`��~m�k����[}���.n�ӼSm��{_�Kzov��� �s�t=�t�)�w}u���qh��w>�kg�\6���G'�c��'m�k[��׏�풎�:ߚ�QW��K�/�y~����q͞+�������'��3��;�2�Yl��sާq�ṿ�����>=�ˢk��_z�.;�u>�kr�ak~�u��[s���vܣ'�{⸓.<����O?��g���Y�t�%�w^��Oλ���-��+/?���?k�z�k>���q�~9��]o�����x�7O�y�]��s�}'>pȃxd�/|��O6=}�3>���_���ޯL��n���Ƅ�v~[����}������bE�W��h��(�v%&6�6\7j�Q��zc�L���1��=p�z�n\i��Օ_^���9���a���1k��օk_����>�ޟ�m��7\k���ɞ�.�������՗�/}a˦�-[M�z�6˶=��gmwY����������A�,�R��M��q�m�������Խ���-l9|©�M����]��Ү�|}�n�v���'ϛr\�����J��S����s�<j����o<��W���o�����0c�@�̹��f�?�;s���>�{����=4��o.�dx�E�,nZ���������e�<�3��;7}��C�=���W=�z�8j���<z�1K�=��?8�ǟ��\u�'���kO����O������'g�{�g�z�~t�9G�{�y���K~��'��w�~/���.���	�ms��W4\����_���G_]�f�k7�n�_��[n�q���9t�_|�Q��x�ٷ_|�տ��o����w>����z��w���������?���{���{��?��������;��>q��{r�S3�����gv�v����ϯ�¸G�4��[��_]���4����S�xs�['���|�w?��&�o�����}t��ϭ������{4�0j�QG�zg����������m6�����\��%������Ʃk���k߼�=�>�ދ�������6�����	�_���'��֗�m�����v�z�6ӷ]��C�;����?���{�ǳ�ث�m�oՠW2��5���[��r���'��-&�z���]��o'=������V��b�W'�NY�u��u�����1���1q��{��i߸��֟����������fN�54{ɜ#�N���}��{���濾0�o��-��mK�X:g�8nٹ^u�m?�������숶#�8j���?��cN9���_zܵ��r��?x�ħOz���Oy��WO{���~�����Y����><�s?8���?�����B�8�������o����.;���8��î:�g�����Ϻ��k���_�q�}7<r�7=�˗n�ǯ޾��n�ܱ�7��ֿ����w�w����{f�;���������?x�C�<|��}�GO�㩏����O����?y�SK�����g��e�gwz.�k���0���_��KϾ����~�W�����q�k�__��%o^��5�����y���`�������㙟��H~���0�ἆ�GMu�h5��1�c~2��co����W:o�i�l�ʫ�߭z�j�~�g�y�Z��}�:��{�zO���V@����Mnz�f7m�Lu��n��K��<|��[ݸ�Cۼ���ۭ״]��_�'=8;���/W�[�=�Q������0f�uw���ZG��	��:�_��Io��������=:�M�є[����3�w�ԁiG�qў��빽W|s�o�oO�=���3f\1p��������9�ɾ���l^���t-��o�����x��_.��?����A���w�w�~HߡK;��K����Ǐz��c�;v���Z��<a��8�%'t���~�CO?�G�q��ǜu�����sN<����8��~��~rÅ�_t������t�#�����]~��_y�U���ȟs��לr������]�7�x�Mw������'ny���o{��7�x���fŝ�7��ݫݳڽ��7���~�������;������Ǯ~��'.��EO���iO�磟9�/�?{�s�����x�{/���/���K_���;���?����o����o���޷�y��wO{o��n|������~壷>��'� rX4��< �8>I&�+�jŊ��N��]e��X���I�J����b�s�_�dʗ�D�^��$��t`��r\�su����cV�M������M/�v�*�N��d�?��ν+�ܷ<IF`��'�utT=`M�?���iI2p�{�94��V��@���uK�j�^	ϯ���������v`�dc����ߍW��U!pS�0�0{��_�+p|zT/^'��L��g�Ex���F�6����?ݿ_�ߟ��S����|=���+����;���^���h;s�{�
L�K҇���������%������2p�8d��-u�~8$�������}�[�@�K��I�ecv��2�E	iN�g��Z�� �A�[W��c	h��b�O�9�f��)�ՖLN�1f+���b�s��oD6Bm�	�|��Ԃ|��Ѓ����?N�iG2�nP�n�^��	Υ~�C�S�h��|�Mh��\�cMK��}��Y������'�aӈ6}�J��d�>�����\�$Нh�>I	�L����$å�Ɉ�U�?�2��ԇ�M%�'�&�4��O}H"Ȝ�O��$��?�ҥNzK�9��V�0�tY$�@%��C_�ϛ�~�9 �6C��h��c���o��Ѓm�ܩ�/�/}�1���|�w��Ŝ��;{�y�Z�T&���v�w�N�6��^6wn���Ќ���C�W{��g.���^\�?k�����2��}R�䖑]g-Z8<�?��������6���ӿ��ٿ��L5��K��d�:Ј�������v���T'��tu���X�i�<���ob{g_Oo[�$1ܔή�I�m{m�sjGo{cǔ�jc��	}�Í�ޖ�Im�}�{z��v�M�6���=�x�:�U'b�s��u/h��.��`�s��}�B3V����w��6��Kw[Ϯ���S>�	-=m}��o�X����jk��n�ȻuL��&c�X\_��NVm����̘�jmMp�XZ�R[˔��4V&O��l�h߻mb_���4�6����X��>�mJ_��޾V0L�n�m�2��kJOO���6�T�І�����胈����Bo{*�K���ͩ6��T�[��ՁP��U[q��gV�Z<'H�Ty��l�W��Ϭ�'���Se����͝8�����6yb�ܕ)zں��A2˳>�THqBGK�n�B;�G��6����o����l��Z�Xٵ��7��x��}_�Wml���tN�һ������]�z�v�چc�6N��m�{_8a��5e2��}��V&O���݇�����1�����'�����B��[�i���pJA�������u5ɾ=ݿ{��vB�{�=m�=�L�sT2�v����Z&4�#�dk�Sa%�Z�״jT-���U5�Së�ո0�����|��OV���g�"X�E�1+MZQUvSߏՌPR`M5��Q�)SVWtU���/c5�,SUY��pK�	&S!*&J��%3�GGX8��S��ظ��~R�D&9��(-m�*��J��t,�,u�gBXj��GF+�⺒�И�?v4�yVe�k�a�c��d#T��Q�Qe5w��"�i�0��2��T^�b���Yn���2)-��M���(;��1���"���L1[5�$�}d��������יѴ���(Q�T�1�����*V(3E��A�d��8F�4V�Ɍ�c��:�d��wj܎>K@����u^� �h���F,˔��g	�	�&B2�II)�
���DZF����f������D�љ�)��ĖZwdҰ����X��L�-�z6)T�Å[�)�Q��pH���� �ɌT�&d��Y-���:S#�z��!�&�f��c��3���VO` �rͱZ�o�Z�yjmN!�0jR�z�՘4�\b��6�*�ak�����$U�,�*+p��aF�jR��	N��\#�q� �V*���he���5�2)�r#`��=PY����	I�]O��X�m	��b�ؗ�}a	Ο�贄PX2�P9U#�ġk�R�
[�X6�hN;�#�feʉ�ڹcq�O>�s��#��I����N>'��N*h��,�B=��$�!�Ԓ|)�Nji��n�c&ͬ'���(�p�b�Y��*�5o�uDF��Wd��֑��d4#����� mWp�ďȝ
Rc��0h������ؘ�QW3�0PZ���P�
���{������V0v�c���P�GW�4��)X6l�,��.�9X��
�!�
�9�[G����9~��;l�(HѺ�f�S-S�e�)!x p�
6.!j�T����(��?����g�(�����"��U���6U�TBR�
�#�g�k�C�GX�)q�>@9�(^{^G�PEi���p��A3�6��[=� �i�������a��hH��K"�:�+���疤
5�)Ed@%@�f�0�Ԃ��@�pĄ�2�+8#�j�FZF`|!Nj{���6�8Z���7VuA��BpO%N�W�)��J���F��* M(��JI��p\���mf��RZ�@�H�X�V+1�_G��Y/!��R2L�,ڈ
,E���u�$G��¬�z8;�pxX�2�����$M#,�(nY�$����q1����% �T��qdX���i�F(%�:��f@V
SK:@& {��ZJG�CiZB?&9��ٚD�68����#��B���Bt *��U-
K�YOh�m�f�U'U�ۑ�`�F�wrHaL�>��@dX*2-�aF
VO�&a���dH�Ҍt�֎��0Π��a�a�{p+`W�ϑX=��4�גpp��wX�EE���!&: u�"$\�%,��(]�5D�����ı S�c� ��)����W2�>��E$geK2��[��4�I��L�ɠD�ӒL��H~�4�L
���<p0L�_�+Dֈdڥ~��5���e{���*e����8t�đ�U4���u�b2M^�B9%��W-�=:��Q��:H�'���j*��b�����H�#+ ��'C2���U}GA����#�t�^
�uI���(B�(��(��g��z�-�'�X*2�|]8aC���
$\챾#�#<�Qsʩ0�Ó|3b��%eq UC�AHڎ�,EŔ�q�9��!�������{8VSVȉ'�����J���LX*/Q�(.8C�����<�BF�E�!GqQ���cF�f$�.Z芑%E��! ]�<���QM��|ᨒ�#� �t��
�����[�*d�xc=�g >H�E���H�tMZ,Ք�1�����Fy�&B�V1��Y��%�֨\J���nIu'�i=��u D�����Uj5:f%�@�`�P=red.��paι���� eU�:p���:��d��/�� `d��i�@x6+�XZA��?F$Y\80��2b��T���9e��UB�����P=^���c\*��8xPޒY!]� �V��Ǒ
��"�{��b��2:S��& �!�:�hH�(�� V�-q�EGAZ�H�sN
7I�V�Ҳ�S4��"'g�z
"�U�Ҭ�g\,"��J���L��|�
I�GV�Z?�MK�F�\�5�r���K|kT�T��|�����@��%�5�pF�.��\��\GU����\�l8;CU$��'\zH�=���EO���\Ru&���qFs�U���%�=����� ST=�j�EONY���*ydEU ��1Z�-�:~��6p�)%��r�YL�d���b��e������9a�Գ��{6v������M���'+�& 08���34�=y��D	Q��a�������K(=E��B\Flir���irƥ�lG֔�{"IǏ�'�Hwa��o�T%�&@oq��q��ʼ8_M��%3�ۃ�b��V�9��&S�l*+�AظO��lJ�3��L=��9mI��R�|"	@LU"CY)���be
0@CN�ƔH��
��²��b�p����"�p�1V�5�e*` -�s��6N�SF5錕=��� ߗRM2/��:`=\`��g$�p<B9-U�Ud�J��%^3�SQ��rߔjT��D�r�J�f�d�v-�Ne�ڒ1]�5�JPq�lؐl54����֔@ˢ'U2*i#OE?
��dX����k�U02.:OH�Q�N%�IoyiS�l��xIFu[x�n�>H\�����)*�k*�"�PO%��J�Iт�)�r5Fኍ�)�`ٜ�)z!*N�*�@aX)=yL鑘(�&QBS�Pw���fS������ğ��fya3��ss"��<y�����%'8Nk�uC@���� Jz�����?���\����l6��T�'�/����^II��i��lѓ�}�]	XC@N���e./����?9˔�G:Lm1���\A�	T>���y�U�'�,�����9HZB`,�r)I��5	5԰�
���5��ꎰ.W��*�ɍ��e)|�I��)0r I=%�������V�5�
�R9^I��=� uTCr��X0C���2Ms��}Cڢ��R�l�}�O�Ӕ���27�M����C��
[�oG����U�YQ�Ӑ��e�5�Q��<5ݏ �q�!���[f%�6��R�EO�$=p��D��IVҳ �
�vT� �ߑP)�[�K�m�	T�b�S�`gy����S�[��(�
hKF�`��=�Td��~����]ʧI����Jz��39��T_�G����2Y��>i�,/=��J�?�GOS�ocO*`[Jv32q����0�Q��I�  F�ψ9=n��JCB�4u,.Уz"C��j��V�a�L�F����B�\3�S�+�g�%��
�8��È��`�);��)^��O{��y�f��H�4^�%D�J;��pY��H�M�,�a ��E*3����jUYRU�kK�\:w��9���.U�����n``�0���m��}���7R 0x�D����C�C_�!e�BX�	˥{% R���(��2Oغ� �]�/��'�YHH�С��p?Tc��VL*���0����H?�!��j#�I�:�r?�8!������TN�tY�4ܕ�'�7-J�1�r{� �	��T==�AX��7�DQAf�f�,.�U�&��݁�8�th`�SWa{�/�_����{����IlXn��ɪ��ͫ6/v�a�g�=V�g�YW�geD��A�̬�<��e��]e2(�"��0q��o��Mt�HS$�6�I�뚳`��9��v�74wY�__2�```Ѣ�js����;?�ʒK���$]�l�� �_�C",��wDh�<���<�"��H��D�R��j��_IC�@�='-=�p$ ����G�9�JW!$�$�����9^
�<祼H��'���+��+F�k=�s��N]x�*o�H� ވ��l�G�fb�Eʠr�5��ޘ���P+B����v��k��f�/B+���m����I
�������3z���ؚ�e�x9�;��U�.v�$< ���E����t���%.��&�;^�ң{�j3�X�_��Ǖt�%��@��������`q�"���D�%JO�=��"/R�[q��wS�׹�H��׫��p�����|��@�E�v�����mz9@���f5]x ^'�|Ct�)O���o��
'	�jp��'3�å"?��,\�@N�P��?��,U��8��d
'�I&�\�8��r0Ny�1��9�滩,�ǵd�"���ML��6]�9� �� t�!�,�2'9�����,y�U����J���9��̜�g�rx�,_��t�&t�0��"oE��T�Q�nT��y�J�V��'9���#��7�M3g�:0�Ia��`��>�\��
�'q*�wp�=@�o���Oj��	8Mq������b$�7�6Ua�r��w�r����
Z�n�������;Ƽ��3��*�&@Ϋ�kw$>F %�,#p��z��CΠ �
���	C�[�L�A�&�k9YL���F�kS?[F�M�@
Z3�"w�y�5~C��D�B�J�*�F�á�@�Bxڕ�fF�"��T 9�ۤ�����2��To��H�H��5�5*'j��9��vs�ӯA�
Qu��AP�n�I�ΰ^R�� ��@��2A��s��4�VKK�$����e��(�*�KR-�Tj�&�!D�؏LR��$�x��ZI��rT�x^���W�r�A���$|�'	;^�
T:�Y1�^y^l��u	g�ݞ�I�X�y�Y�V�(H�@��%��r@�t�0Y��:^�_��V��1�i��-�#Ӧs2�ao��29o.r��_�&�r�X�0�8�{� ���������Z�{�d��&¼�~�F孚y��B��Lr���x���=#��`�^XJO�s^�a<�da0(��,�K��V˼�2Hʟ<���z�r�Z�O�׋��{��z1nM ��2�,�k��'0,���9]~$O��y��[e!3���$]/��䭖{W2�����ʹV�!
2+Zݵ��W��W'>�]&H���ؓ��CLE�@
�V@f��܃x���bo�&�lP�p�p
a� S��0����tC(�a�a�χp���HƼ��s�{��d΀&�/���y �7'j����Ѽ"�N&�������>܂�ޤ)8y;��0c�pƆ~B+R.�[`��B?Y ��<b�APpl�s1���=o�a��Er������j1G���ұ/���-b��f��@f�YDé �=)�7�Z�x�0� Æ�����)���a�IX$=��;���y�������2�\y�0��޻6�Y�Ф��FC�
�t����
�ވa��`�ظ1����-0���z�.�#���-0�R������S��1ś���,�&l^��@�S��I3<o�0\��H�4D��h��EC�e,92m�'�!t'bNɢ_$2�p,�	ڏ1���nd���T�����72���d��H�"bN#����K>CX�[`,=�q�2i�ڸq�/�-0u
˱Y!>xu�y#��ҙw�����0���j��]�H&ț	�[`���/�[O�b܈a��� H���Af����#d����7b���!��O
�~�=E�0�򮂒��MD�<o�a��x -�>��a�r����YX�~܈a M�,|ؐ�nOb6/߈a�C�>$��@���@�ў��0�L�H΍��1�@?��f�͔.Kz�@M���Ё���-b!�}�W�,����T1�롄���߅���x��`9iX/BO8�)�y��`9,���0�=E�0�>� |*���,"��夁�:����-"b,�8 �� u�JK9o�a�j�wb4H!�7b,Ǌ��*�P�\2b���:��4��c<o�a��Y87+-ݴ�>JF��.0d�}��Bb�2bh���ܧ�T��DF#�9�p ���˽?�� a�6������A�*X`�R�'!4/��a(��Ɠ<�51�$������t]��F®�n��r��<��Ðv�4����:����Ǟ ��_�\�P@�[`L�|R,�Qz^x<��"b�� u��4�!bI�KR{�L5��d�0��W�ƣ
Ƃ>D���"�*�	ѝe���a�Cli��q�+ˈa$}J�Ҋ�k��!e�0���ab��FN�7�����6�XVF����F���%��7=BϾ~&#�A��ӂ��&�_C�0h�:t����ч��]D�)DP~\@	�T�0��n��e8M��y�Ì�$���U*�[`���TB>v�"�Q�|�{R���T�=o�a��F*�̇E�H�y�Vnϼ/Q�ٴ��T�0he>o!?ώ��Cy��P}�ט��O�h0_SP�(Ƭ
XC�nZ�Z��F�z�WPY�S�Y�����a�Ӻ:�,xp�|�P�(d
^�0����v{�"��G7^a�S־N����Ӫ�a�(­"�����[`E�݋��|��9��FQ���F���+]�'ވae��W�\��_k�[`
��#����^�"�Q���t;'U���(�C��C>�x�-0��7����C@A�1j�͈a�]���w�{#En��7bE�A���t�<VE-�R����.�WE~'�6ԮT�0X���ڇ��k+:b�_� *W�[�OG�<-�nE�8'5]�d���0�� ���͔���6u�0t- 2X�	�����a4\���G L�RG��"i#�^�Zy���P�g�4�7i�<N���n�ã8F��E��:bM�M�C�I�|\G�� ���Z�`0��F#�
��b�	}ݐ_C�0�KLgc0����|ܛ����p\��N�0��Wx���̯!b��AXJ���Y��SH��}ZG�s�S(_/:c�? (��EG�)�w+Z��O��7b�B^jxT��FG�P��Tm�#h�ĝ�F�)���$�ЪC���`
냰F��}7d�ܯ!b�B%4���H��1��~�F�p�pl��00EȻ����}d��1��O9����yhU��!1ZUP�x����-0ZC�ӤL�y��>�<��"I�-���m!^�M�0���'x ]��yC����(��m�DC�Y��oy�
��M�0���=���.�h���a��	Cw;��Gx�EC�ث����:�����-��y1T��{�����A*_�6�^<;  �!��Z�_o�0h�<8���>@q��I11��R>䧀�8d"��
��c����!�2�ա�`"��O�zwep���Kco�0�����v��1��� ЇR�a9����-}l1D>B��}_c2��a头�Z�a�?3�P�#�4h"��;&b0��
9A����_s4À!����g1��-{���ᢔ�]وa�!��
�}y�N���Vz����rL�g�B �sΖx#��n
0�4a\c|]�Fc��B7��u?>^؈a����-�p�ҭ4�y��2�Y���������-0���3�!�)�-ڈa(5������)[l�0t@,08�H΍`#�A	�R`��-}������6~�(��F���Y�0�|��Kxޏ+�T�z#��OVa�B��>�yc��&T������1}�0LA����+9���0��t#0�P��~�F�)lV�R�H���ڈal��X�� ��t�y<Z(�~\�&Cn�P�!��ħ�o�a,}� t�Y��1��.9܁��m>���
{����LO�����l����C����~�
�Oz�������`�Zlh�.�����$�?N�Qh*�   	pHYs  %  %IR$�   �eXIfII*     (           >       F   i�    N       %     %      �    v  �    �  ��    x       ASCII   Screenshot�Ē6  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:exif="http://ns.adobe.com/exif/1.0/">
         <exif:PixelYDimension>1190</exif:PixelYDimension>
         <exif:PixelXDimension>1142</exif:PixelXDimension>
         <exif:UserComment>Screenshot</exif:UserComment>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
�QM  ��IDATx��i�۸�- )�d������C����V���*W��QI�a����i���t�.UfJ	�@Ď�>����H)�X^1
1ʛ�r�0�0����.P�m�Ϟ2��q���@�8����XN���];�_9�^Ҽr���k���é��n��������@_~H�g��_�Yk���;�}3��+}Ѵ;���gi��~���q���Z�Ξ#����T�)M���!+]Wee)���L���T�4�h�]�Գ��Y^��_��Ǘ�Z	�E*3�s��������z|=���\����z���z|=�_�3G��״1;�jk�8u��7��@��@OJ���2MS*�nq���@�|>�8N�o� �;� {>�� 9[TL":�?������e��S��6;TR���Q�����b�Cy�s�U���Q#[�wb����u{�������z|=��b�_����d��O�YN��k�����:�_�/=���]f�;ڋ#d�տ캋˝:ψ������!��)��G���o$6���~y/v�E��DS�(t��9=3+>C���o��@�o�Y3�:e&���E��3�����G#U/���EmZ���),o�6>���(s��q$����KF�d���D-�7�{�]9w��G&:9�������qN��_������k�۟}���?4�w~<�)?������Ѻ�_�K���~s������xCk��m�Nԅ��i�fh�7��6�����ᑞvO�rb��Ⓐ�[�R�1�޺� �N >K;�OR$ .�ia�*
w�GO����I�-4?�9��ܠM�(As�_�|���ay��#��te��y�$����ݏ@�95��b���s��D����"�+���?�7?	�S�߉+�̦�Sn�'�zъs��3-y�|a+�����N���?��L�? -��.0���:R�����XF�����q'?/o���c䗟�;�+_���x.��;���m_��Y�z����:�;R�E���$AW"!��_Y�F���@ρ~��+�����Ġ�۷o�՛����^�S��"�/Q[�%��i3�(f�$�B��"_l�@Vh�A;O����nM;�&Ҧ���O[I��0o��liΘ0R&��PO��H�y���߼�N�~�r3Y�)�_��:�_���.��,v�u��jvݶ��o�;q��x�9Q�9��){v�;NO���
Td�">�suu2	�gl2��.��ѭ����Z�4g�R���|�jĭ�_���>�뗘�	a�W�����Veb�N��l+�l�Y���~�V]=,]�^�wUf_r��@O�u����s�n�����`��L��f:h�~�x�)�[��*4��[=�%�/����!��:5�V�����qYϬ���^{Ƀ�9Nm�o~�_*ek���=l�ˀ.���"���/R&o�"���7˧7p'����VF1�����|]~���	0�r<�n�k����s�N�����n�QgC�%��EЗ}|D�L�w#d_֗��B�Z��t�TO��K�Mrr9:{���U�̹������zN�w{~**��fN�~����-8 �M�1��>L�������������_cف��/?з?|G�'f��ͳ?��{��.������Q>��Q�����C.�\�a��K[{����� ��� k�Vп�{�VƏ��94��m,}p�������TZ`'4�����:m�Gv�~����I���l����G�l� E��M9������:~�i���]�m̤��
H�`�Nmd`l2��Y\}��=[,TVpO��4��t��p��,?�i��%kk��R�^�8�B��
�Y�g��P��~���ܖҷH#D�o|��nYCS��H����?���o)X��s�˵�H���,��X��׃^SV�h��2�v&����8Yi�@�V4�:֎өp���s��,,Kmh���/9��͇v�Dy�9X8�� �g}�|�Y�r�,y�}���z��ڍY�B�����Y9u���g�����2��޶��p��V��_�F�%��s ���G^y�D�|6x�r8����xǝ����3��Z�k\'#t�9�_�'��0���ֽ��If�P�NUm�g6yv˗��{yHɯ����ֿ5�L!��O�wr4��֌��HɈ�z��"������ƶp["/M����:D�i����̗s�7��o�h��|��<�3����r��D��cŲV ��j�f?�-��,��|��֑��r��ϸ-����=�M��3���~�/ڛ�/Ν�P��ܓ4�H�C���X%K�8�C]O����^�l?q��g�=����w����s�+��!M�־�g��IbQk�y�s-��nG?���ۿ�+�:���A	i6���}�yU�+�B
=��7
�G�Y%�)�T�aG��2N�pR���OvO���	��쪄����q�a�u�1�2���>옓^�>�8r� �i��vo�J�s
�I�`*v�O������p��
�*[��Gd`g��N�J ]nF�ױ��l�;uƖ��&{��Dp�P�U�]�ZvJ�>B�6�߷h[���~ό� �1r�0gv�'`*�������k�d�,).�u�߃��@ M�y�Bpg �� v�7@�������W�G��(�C�_�E��|�T&��e��s�[t�d���N}�Q��l�̶;�TsMSq���|:��I���X��N�:��Ͼhϱ�ߨ�V�7����3�Չv�`�1����������ͽ+[��Ǭ�����2	m��'@���8;w��N;����(�qGu^Ο5��V��+�n��3��'~�'���J焏����۟_rs5(��^�v����;�q�s��_z���y�����=^����oǬ�^�ŧ�0v������߮R�����mU�aE�>��^�e�i�Gk�i�|�[���|�|���r>�/<Vl�����<\������]��O�b�+���Y�����1���G33Ȑ�?[A�.R��/|F�ά��_z���3���Mۢ���JǪo�)���ϐ	Ԑ��k'��e,�8��No��D�-� �S�B@�X��&�9��8o����S�/��������Ͽ�����J���|uE���-Ma����ô�Ŷ�}P�"��c�HV#��d)S`��q�t�� ����KqP��@R�t�	�@y�!�#OdiIY�#/<o�,]��RKS���#�ɚ�u��g@F@�n>���ʠ�Cc���%�=KM��q��}Ų��/���=�O)x����"M�\ǀ������;���_}' u�{e0,�P�-�tA��nJz*r�v��M |�R��w{���e�� 9�n�_���iG��bF�@�S�73���Mv��s�������Zs������~�����[z���� �2�ڭ�O��&��H;�.G1x;�έ�,�6-8�Rt�y�U���\���0;o1�g�Td�:a��T?7�F-���/�i�XP�{/W��z;;B��5�揣bh2>�u�X1f�N09?�L^kN��8��9w����Zɮ��^�\E�P �� ���
<g2����6~q��[��+��/�ʜ:~��f�K��Ԇ���6�9c�<��%y�Z;Z}|����#��cs�Sv���cp�X>͙/7��lq�Lw�VۺY��#�Y�f�Qc��ǚ�y����W���'?�������9;��3�dtmUx�FN~?���l����z�[/���N-j�Î�{��_na���%��%-[_xW[sjM~�)�����A��GL�5��¢҉�?j{ӟt���?�X�D�K����w·ުb�W���i�
��Ak�f���F���%�ā���\��ٶ&�����Uk��	�T�Xy���������_�J����LO z��2]Q�2�A��S��"�2;��^r��5a��(sA&v�'u&u���N�FN%�,%N���)4J�Oq��@���qi}D�"qħ���HM�n���3�_)��X��-���2�Rn��q�����>b9��W\�x	�����}c�p�����"�$����r�	��?���y-m'
m_n�ty	Ġ�o����>�y`�<><�ݧO�	�@�1���5;��x�� cd�T�t�g���ot�V��?Z�W���W�^�w�}����o�}�X�(IM���P]ܜU�ꘛYeP2�#�XO�`N\{*��<�1�ͥ��)v������h�SS�&�zW�����eu�P>����y�f�G���>Q���\��P9-�{,H��m}ƐKg��<����ԩ���V�vk!�ӮAZmy�G���D�1��Fs��}헖5]���k�V+g|�q����}�G��km֬�(��s��R����+Y崥����U�|6[�3-��x����c֜�����Rc�z��������V�@�|�Q;�ܽ�{y\(��I�axA��um8���5���`:�AN��B|��s����ܧ��SZ�W;GՒ6�K��F+��^t�ٱ2���꧉��c�����f﮶�(�`�|1d�Ӵ�ؿ����u���q=u�����
'�L���x��+�|=o���|�l<�.��tn���zf���[��yS�E�?)��;�P�3��1��u�J�[H�K���m��M�Cӡ�,����j��V׮�\N<\�۷v��o+���m��e�:���\�x_���`ɖD".��OƬN���*�Ç�"�Þ>�}�_��~��g�ɹ8���3���\������2�r%Z/���a�߹��3&7��E�;��^R�zI�P#{�W�b����08MM1!_X+��VtY���](��1�Iҿ&g�x�+['l�[�k-L�� >�j�0(:eR$ Pcb��,������b�5�b��H �P�f�.NS2q�g����MrTЯ�6Ny�8��`	c�iz����:H����p��~G�wt�����ǧ��O���v�x��I���3��
o����hcJg,Kà�4|Z`L!�0	��c�����[VSL5Ye��S]F-P2�oSM��XY
�uR��U���s�7O�R�;���Z���㶋��o
�`�]!Wf�lĦ���ѱ�  V��։�%�4\肌���Bi�!���6��������~�V.�=7��T���[���跴���Zv�2��^����$8�T �(
��ٕ�z�}�|G�bma�����|aԺ`��y�oQA{�=���������������חZ=+��W8��H�L�Y�[�����6<K^H:�</����4l��({P�Rfa[؍�Ƹ<٭�x�|	Y|ֺ��d�>�Gs��Seϻ�V�w�y�M�S�e@����^���\W��+W��ё���w~�	z<�|��Ҋ�n_�m��j-��g��>��������r��
���G�!�?��k_/������s=��/�e{̕�aZ{���k�`�y��,.sVJ���;U?tɰ�;�R�`uAhΙ}��y������b��y+rc���X,Zy���h���ߺgZ��g4eif�< �z�玵���͉�,�LZ�^�x�}n19uT]kvB{�ls�,�YA�6�D�g�d@�75�Y�+�����[�t�+k֏�.��R����-��_Z���<���X$�~��PF�(�n1�i�SNI�Sw���#��������~��g���#�������� ������@Gj�p!��t�ԯ1ܗ�`;*Y�Ȍ c�p�e�Hq��.X��5^..�tq��Z9H��p��t��cvo�>�,�1�l`�nC�F���A����6��8K^Uу�5�W̞�k������$�7�	���u�A��=�P���: c��2vex�P�	�%UH�%Y������'�H�V?x��'I�饞�E�|�B�@PS�����D����~���[fq?O2����>��<�j�aW9�S�p-�-~B��V���@� � lw0��]܄�$ŵ��|a%��0O�ږ�]�uq��v8���(�w��4pZ�\;�Lu��U.j�[��5�&�e��oeR�i?u����n"��j)x��,Ȥ}��B�=����^3^z�{���lg��e��y_0V�Z����i��9q��૜.����S�`yY���Z&`�ty���)�y���^[~.
;/R��ٓEW���쥅Y�2�����q���cCō˙�]�{����C�{�wtX �l'�k��Z���p��}��̨�;6�d]��ҙ�3<�j𬥫�\����������To��|���':��]�<��s�^ʬ+�4R�զ�Z}ޗ���Qn���=�֠�z3���S��6�B�g�kݬ�p��o�s$/O�� �/�bX���;�o�<���o��Ds�7����U=(c��ѸG��Ղhכ��NuԊ�a�s+���l�'�������<\O,<�}y�5ۂ��ٸ<y�v
�	i���#<�I>sF^;'�a��5�lA��r��Sz�2�7ذ���8K��e��ln->w;��r��w�D���Go.�ɋ���ԥ��l������k6�O�.���ٯ&\8ye��w�1�o��������\�7�0[4��a�r,�j=UdmP��?ھ8��^~��ԇh���ꖮ^��5hX|�?�̉�Áf�;G�;fs�)<��d��������V���O��?ч��ӧ[��?r�8�`o���̦����������==2K�o���5��~ Kl&N��Ǣ�l�sE44U��߃��w\���p��]��ʻw������;n��eq¯.��P��NPz/��{�Ce8� �F6�a�8)h�����I������AvkJ��]`��W;b~.NIJ���o�&�fө�݉W�J�Z=�r��9�	� ��5k)HYe#�J"�+b8f��M��V@&�E��$q�ў��+z��� ��M����{z(���/?�m����{�i�'+���E
�fg?i�cN�3hS&w��0�c���uj-��L�`#>{zzb ����;(���n_�����>�}7,O�o��}S���o��w߾�:T�E���/�wquE�2�;�%����CW���b`�w�3V����B�L�h����n-�s�s������B���M��*�}����2�b�en��k��ќk�Jk �;lZpa���N��u���Ū7*8����S���pqq���'�o�z3���굙q�N�;��43��;�K����uU�!��ϭ&�	`'0���*�}�ᨲ�����������E�"�k�K�Z{��{�k��yK#�h�����~G��Rp8n��]ۻ�Ÿh��i�����hS�}���;����ȔZ+���f�nr��z��k���16,i ��}�����>�IYtߥu(�YHg�@���0mm��it^�Iɬ$]�M�q f�/�[��.��T�vTs�.B�a���߲-�m�`1W52���~���g�]`��&�r�<�ڑ��g��1��ئ_���&L��6���]2o]�m���vImmj��V��1v��]Q8������8�O�7ϱiZy�+?'��W������Cti]��]fO��z>���w�х�o9��(�L�L,���1��h{����LF�f�G���p�x���=y���s�\��ٲ����~h���K���y������H�^Y�e�N����k����ǩ�z���̛fk�k�8�a9Ϲo������0��/ܱ5폙�jכݢ�Ĳ�
��X���"q�Q���덙�^��!�DC�ԡ�F��I�TlW�㧟����##��)�k8�Jͩ%��)@ A�+�O HH3L⶧v�6�8�`4`�$8��NVhiT��=�����`(��vC��p�l��-����������D����@��"��.A�UJ+�,b�c�)����gG{pD�ʹϙ`�l�l�9��V&	�b�	� ����:a\$��\*m�ì�Iw�¶����ʃ�-�lM2۲!��ߜW��x2��C�=��	SǷo�p�c����{z��=����"78���:�"�ff�ع� LMZ�IR�ď��C�h� �Œ�����Y��Q�sK���<3��0d�N{���@	'9uA�eb@ �nرㄔ9���'z:�h��`�a| � ��3g�Leq��ئ-�o�g����,M���<9�$���13�XIj���ϡS�0�neO�8d��]��bKw�Gz(�)ם�L1SU�霐�����s��Z�h�IeU����i�� �1j��uǼfYm����M�5+:���饪7e'>��'c㘒W�+7�6f�D��A�퇹2�X�G
c��Ⱥm=��A�7�g�*�Vk�f�︉����㽞ǔ��&������$O�[^��A�f|L<��E�y+���0FMim�04.��j{G���rV����9�-��wl�
66���Z��`�L֠}a�W7�_Tw���Kͳ����@,� 0��!K��>F��/��w�7�7����N�I"�������(`if�Ik��U��Ec�ɳ?|�.úa�dsZ&���9����s�I��,2N �0�[�e>ƍ�r=>}��	�R�'�^�\n��Qk��LK��S	��
��|0;��r+s�ǚ��4hes��fps}&w&����T<�)r��7
6gj�y֎s>D;?Vϫ3c�Y�9�Ⱦ��>����L�*�0����9�H���[Wꑖ��խ���sm��s�5���o|͂��z�t�z�u�O��f�s;�Ls�-L7ry��ب���m�(DHm;��K\�j��ï��r[u����h',�H�^U]jWTY6����ѭ*��JҜ:g��������ek��/���n播���������Y/S��(���tS�ǃ� �E���Hb�x�qwՄ��S���).E� fNtu�uI���/�C;nگ��_��f�Y�����8�ѹ-�mS��Z�2��ytT�9x���q�S�����:iiʡ'��Yx.�t����Yӊ`S�3X�YQ����㫇���?��AfS4�`�(kj�Qfy��ص� ��H�kJ���Izv-]_[�M��ʺZC���!,�OV�4���4���mi�w�"��י�u=;Z�n,%?�/Ũ�� �=r��3g�XK1�Q�W�y�l���{�/?ᤏ�����F ]������KF�e�`�������+׺�����t+uPR�|�s۬8.;�wX[e{����0R�#G��bC�`�`�$��T���b��#t��6H�1�C�|Y�v�.F�Й�� h&64��P��^�k:����"�w�� �����S�t`�wf�d����P�l|��,�q�ԑI���0�>�f!uȸ="�l�[;a������gfR���s�HQ����8��"')���o^������������o���G�<�����`��h��Dݖǳ�����W,,q�t�t�Mκ��\<;{z_������v���%��*^��
}�>R_����Ӂ���������yu}ÌK�{<<Jے</���,mO�ڈ�X�t�$elTP
)j,?�VV,oHH�cP�RR�9䎀2�r�{�Y?
{��� V��a����#}���k�Srp�v��H�ֆ��v6V9:u�!d��4��\�5���q�,e-1X�̤��X�W��<����Y��4K	�=&ٍ��=����El�HZ��c��|������w/L�hw�DO�E��wQ�����]V7�YFV>W��؄RS���"��̷P�%C^{qX�WE���&��-�&�7�G����:Ό���Eg�)S}�r���j\��f�[1��F� �Q��:V�_�hm�������4/�Z(����ɀ9>�3`��D�̻I٪�E��x����H^on9�!Ӽ�Ņ�L�H-�]S��$@|R����3�j�l4�/�%����y {�Σ�Z=}�/�~�m��e�T��r�SN�tL���ZR�ǀ|�� o�e�|ܼ��ׯ^�� ����ݖ���Fu���A�ֹ��3y{�F8x��,g���}��;f��==p*jҹ��`�k�0U�"hu���{��Pk0J��j���g���ɀ��G6Φ��������p���e������E)g�v�v���[�*�5��4��:Q�%�w�X̜�LY�~rѨ�|o�BƎ���I� ��]�i�X�ϯD���u����<�1�`󏉃0��ص5��\��&;5�V�����*�A&�O]�`�o��:nVU��f�A��v8����x�]M3^Œ��y�,`�Z�uv����l�l)���p,�5���K=�o��=�88T� mL�E�G�_<_����H[O+�v�ǰ`u�z�A�����c���Z�����ـ�S��$�CDr&.%A�+4��0{�|�q�ne�`�b�c�?��J �i&���9�1�͘��mw������)�>�z�Q�Ci��y@He�m��\�5nz�`�'��e�y]�����鹴qH(��0���<V�;0nõ��[�v�\���:+;\Z�c)y�/��d%�N��F�=?/��U�̠1���.z=�r�F6��4�&j����/��Жڱ@���M�q�L�jM�`�X��e��Ǐd��
� HFV��J��<�ne�9���8
�gs�Դ�]�b�&�U�WW:t!�b�b>�w���!��Q�����z>�Ú��"���n�y�s�<``��b$��6j�8�����90kg􅝋07E��0�t���T�^Ҕx�92��#�v>�PşO\D8��ߓ�}�
J��00��Ż�p"�F8���� ˾��sy����
�x�r�(8a� <�6�Ԫ��N��$)" �FDJc�ȠMl��>�ݗ���F�}=�"����Z����Pe͐un	��i](:� "��� `���>�H�_����,�Gr���I͎�mOO����#�����P�41�O���;��$0Gjj ���XdZ@&O��Iis�zz��[�Gfހ&���x�/@��9���.������5��ߗ���;U}��,�f�b<g`u?j��!꛶��Ib|rq��:�h$�ZP`�����%lL�ˁ�W���9 ������֨�%(16Z���MiY���%x�0c��[�0�Eո4C��ʞP�+sg�\N�r�zCn�b#�Ψ�`�fP`����e�!ek�r߃�g�Br����ߥV��||m7[	N��|��'��b��3#��#�D�o����;��H갳΂a�ˢ�]��v�e" t�®p��� �:��9M�DYskqfMR�V誃 ^���!�~�/�o�Y���P���;��|��uk�⤠N����E���Qr3Yl��qp'���zw��fό�%���xbgB/�nk*�����aQ���e�D����^Swٙ'��8"f4C?`���Te��MGT x�`g�mQXi?Ї�������:��[گ����c�D
������t�t���6�z��|�޽{G�򂬂��ӏ?������H�~1 ֬�9Wpǘ`Og� ��9=��Q���7���aǀ�;��y� ���p�A����]M{�D�;	܌n���q�������r>V�S�Fj
0g� 5�g�kzz��K�k���)C�:����I����f�Z�qN8X�ΰ1�m����M4�w�=X�;3V��a!W�#oE�k���f�k�Hn[��vC�+�Y^�Ӂ��nk����`�ؑS�kR/y\������-i��9'a��rۦ����%��P�YY�&����#���8�S�?�w#��;_>�Ͱu�p��l/���~�����,�қ��7���#]�6i�kM�6�äv}Ե�������<����S�"_�Zy�uI�g����:�T}�\7r�̎�$�~X��E���<u`�j��p�a��l��Օ��� ��k��ۍ���'�������)d�P��~�O�	6fU�fu�]�,v�ϽvuA�=\���*h�V�ʟؾ؉�� ��ehX��(-��p]�򫏛�]pk�g���La�����GC�lV�U�rcI��6�`"�=�MNY�q��[ۋ<"��Y����,���O�+�=f�e���@�,䝗�^ �����˰�� pp-^�����Ʌ�	�
��h�B^:T����,=:�t����u�Æ{P�&GW�0���9�yx�ݓ8��~p�K�$`_p}��;�LeҦ�H���������;hj�3�.;�� #�h��ʂ�^;V�uSV�����A�) rU��77�D�,Q�ҁP����A�%Gl;e�h�QI��]�t
D]n f(e�hJ��7d�kۈF^L�����lh��L��fA�t����T�
R���5 :X��}�XO�>*��Uh���Ru٘�t<VO�'��"��� �j�	�=9����?ч��O�|.�����>��Ik��Q�'�9!�ˍsM��-�4 W:��o]!g0���������<�塡
s��Z�Y�W� ;�w��<�"�~��8�����5W�E�;��T�\)�5��s#�-��e>��h ��"G��Ag�V�~XJ��`޲g�q�Fޑxǫ���^��P@ ��ʾ��9��:����f!���-��LՈ��$.�w�k�6+ul�-��ro�X�bλ��Cy0��,*�V��b����$��+$5���Q�
*6{�)���0�.rY��TC"���`E֝��p��F�# ���`6N���� ;Y�GV�7��"����
VK�K{'��Ӷ\�8��a*������.z���V��1x��Q	�)GC��Vktg�V�W�o�IY~&]TX��ń�A����z!�P�0�á���V���g����r</�"��sYЎ���S|�F7������9���D2`����{<#�`�s3�y�C�+�a�a�(.1��r�`c�WC��2]�P���⊮�W��)p˔nv��,�``R�ݩ�Ij�2_��,���8��ϕ��{���ARJƤ��T�G)�������8��1��i�;t�w�K�~�k<�_�]��������K���u:V�'�huG��a���\l���- ٕ9�Pּ!���c/�f�S�&�/�/&)�E�cd9��c3fB�[7ҭ}��l�j�:��	+�c�@X1��Ѯ �����u��,wzN�8��N~.@|u�2�n��a�Ƭ�*���U�n2R�34M�=�>�R[g̞-��qTPǞ�d�&^{��$,mI_��]�{,s�aW~�h_~�?��w�39(:e��(��*�Ҥ%��_�%����_~����{�����9��� �/Ԟ��RRP�s�_Im�i2p��,���f�9r&��%v�`�+�i,��ztm�]�w#D~ߤ�Zӽ�шc+����Phd��;��ߙ-����V��&�o���8�>����~ks>+�X�̨���BV�b�`��5V�������c��Cm'_+a1���O*���i��}*:��-)׿��.6�%5��9��?g�����dS�뛷�����t�LL���&��f���z���ʥ�w0@a�d�$e]�1��v�Y����Yum-s Ĉ
��]��)Y��n�&����`�r�
��<V�ׁ��{�
/�7���p2 �YW����P�N����Hn��@�������X/�S� ��Ħا7W��rs��a�$�GY �9��%<�Ι�����[�Tk�ڦE�����cM�]eAkf��?p��	e)��s�.D
d<x뙥���w�,�R����\V���ٹ�G?��E�rH�@�EFc]`�}��7G�
�4&KAPg�F�����W���Š�ldùd���ǖ�rߤ.��$X�t�(^X���,�+#�����8$g_�ns�@G0Iu��a8֠�#�)./br͠��7�Y����p!b��Y/m� o/Qp�+�ոNV�@��(���'K�!*3�^c�D���U���11:�8�)*�z宒���L:�m,���1�Xa�����8�����k�����t��#���Ot��F+�{�z�兒 ��BC�;W?g�T���ן���Q�H�)�X��Wc��^o��h���~����b��X��̐넢�5� ,N�S��]ܨ6�}q|~��+}{�-}z�T>'B8e��
X@�_ʾ	�;LV��<r'?Iz��[)v�E?������91�d��u��X���ؙ�	,�`�ĭ��$<� 12aHL^��8Sln10WAjύ*~UyZ�AR5d�cc�ud�'����i�dqŀ����(��	�+�1nc�Ҿ�:  ��3�|�d�P�چzUܭ��&x}&�d��i��t�����²3�}!]<Ѯ�:+2/\�'H�_'��iF��$�$ ^'��0�Q8�F>r��\]�Y4��K�;��*+!�s T4=���P4j��3Z���&3D��s ���6P0&cb�ܰ�`�gk������R��r�c��Ffk$�;��x{y<'V擑n�It��c���5q�O
���#�2٥N�+*�kZ
�q�5��a�u�|wձ�0�1O������ǇG����Ij�d[Ô��FOۇ��d�.��s�������:�����v ����W�\�	�p�5PH���Fu�侖�ˌ8X������6^��.fM���uZ||{]ֳ���4r:M�Ɖ���aڋ(��E^649�`��'�)I��O0V���#��L�;_��3��@�����<���B����A�Gڝ��*��7��L�|ΝugX�@������-ʩs<�)�5 ��uˠ�<-l9�,U�
���X�-;��W�� �4����f}�FY��� ��qv�k�2 ;�oV�6�ɿ1����6�PO
�@/__Q8�w^���iX���@��fܒ���H��RsMt@���C� �Q�ʾ�W����(*��(L5{�zm�9���D�[ 3GS�U�v���[=W���,��#j�rФ��g̲��w.�l��@����3�Y���vj���`�٭����K�#��̌ź���/�gV����$^��8P��cpgD�A��'�i�!K	[]C�~4� A��A�˛�v�������-u�C�M� �ͥvr��-Ҧ�+��nG��K�N_7UY�ۻ-���v/�,Hd�����Z������Ù���c)ҩ�e��sMͩ�Ӏ�9�� ����OZ�>iMB2`��[�/e{ؓ��N*�g:�]�7�Qu�  ��`�����?p��(�ծ���e��P����O��s���o4���N'�'��g��^J�$lRD���n; ��p���o���woY>�n�9+��c&I��H2#e�F� ��� La�dޠ%�_�I�P�� aO%;��=�:Xr��2c�b��zz䔪���>~��l��!��w:�ºrJ\���Q
x��j�h[ky���������#�"�"�$L!.~���#�s��6�e�PA��)���Q��NF����n�/ޱ(Ȫ���]�v�3��E��U��$.�̹�=���\��VE��ˀ'����ȯ1EةV7E�T��.�`�;X��چ�1�\e�PR�&0��x����D�s�3W��ȶ��]Yt��%3�6��� oz�k���ʽ^�~�������������_x�����.���3ey���~S����8�Jh�`OD�x1�7OU�l���@$~^�Ӑ[�!x��5:�+"�l4t:��	��vɶ��W�� �~��H>�B��� 8Gpؐ��P�2�3f��]͓��|Y�L���M^��j�T(ƀZ(U�:�%Db�gM+���4�7��G�`��:����9�Z��A�ܼVt�/���w���N�x�Q*�����S-X��Sb��־��%T\��b�����*���`��:
�pt	M �q(��fĘ����n��^\�2q��1���'!)��n ��	QA]lC��X��ʜuW<C:I��Jt��P�����?�S�%@8	cӌ)Q+�1w��_F_����O ��6�px�4��M��� �>-�r��N5K�k"�}M}���3*'K?��T����S#�3�GУ0�d��hua�Bs|y=�Ygk���?Y�,+�D�Pi+��k�N@��4� L^#I1RV�tX�\ҿl�%���l}5rT�I�|k
�yYF�^�\vj4�F魯�{Q��W77����w�G����������%��\��䩐i�D�`K�?q�+n=p���$ͥ�,���e髞����C��5 �WlG�]Թ;1K
�kC,�.S��0�LY�I�X�\S!�N����Ѣ^�$i��n ��k�L��TS[z9h�+�\r�E?��;�Bh�E�c|�{�մ3R�����򮐥ד��(�4�|�륁'zߣ;�%�X#��)�=��HҗY�;�Lb�E�vE다�μ&����K�����a��Z��v�1�����(V>������Y���i�A@�	�5�Rd����e{�(�2�_�fh�����&+9p��'��R�	�bۈ����֞5���Qf��!'e��\Q .j='��!?��GT��4�����#Gs�<�^c2�'��į9�4K��5�Rg�����U/�w�=�9�5D�f��9���-Ӡ� �����S�*��p���x0��� r���n|x�Ѵ����kE�5�r���na7O̜���%B�ź�6�U�*��q?p�:k����ƀc�E��l��2��`�ČђD[a����-ܞ]N6I�Jm�j_-�n�7��z�2OL܌�i�.�� �	rw����Z�R��A"y�V4@�.�m_Y���}@tz��,7��]ca��V)X v �!� n�5����8���<��#2��G��ܾ���Zw1xY�NA����4��e�.�ߓ�ϗWR;%h���ݷl�y��� �qI�ŷZ��Yϓ ������JV��^]�����nd�^k7��<7}ޜ8z���ſY�s���)W���������my�I(��R;�P'+#UX"w�/ BE��¡E�'D/{��\k��U�(�P�6u���~�R�4J���EI�Dbyq$'����>�qN^�41QH�_�m���l�o���z<P*pe�I�5Ml���}�U�R[F��f�O�9K�qv��KA��*I��E��=�tNe�@y�@��2U��{[��)Tt�;$!մ)LM��*�
m�v%M}B��,�E��Q}E�c
�Qq:���S/�tuqE?��=}z������ӧ_?r�&���l�ʹ]
Z�9��6�>�|�6��e5�`�#�4y��s��h��9��y���8������TgG�ׂ�Nϡ���_!��l/%uT����Sm��SQl]��[���I�F̚�ZP���M��i^c�"_Vi(spT��g�v%z�pJ�, U��-���$*�i��kҝc�p0�qc�AYeW��Ċ̻��N�K��8	�ʍ.����D��N'".�]�"�^vgSۆ�S \p$���;�(u^���i��1�bv6U��S?�����ncY��@a����Ő:0Zs�$mG^cVJ�x�<��$��(/���{�QS���9���8�i2c����"�G���g��E":M��[��2JLz��`c]���/�2e�/c��'a�q݅��.Gװ��KjA%�V֞O&��$qr� Nj`�>�\�6K�S`g�4�_�2s:��4q*C�eD(In7~
�M���GM#�~��ϓ��X.Z�:��"�M��81u��S{��F��r4��^NH#(���g#��휩��N2;o��|�Zj쀭�5g�޻�F�G8�
��F.����Z����N�(�	�ˑ���#�m =HAմ����� 3��4�xp�'�4�DYJ��e���4Y�~v�a�87$���D�e'amP�y}J��aMj<��v��d#��O���а��eg���:��J�sݎ�qo�?�~���ؙi'[w&���F1*3h�g��s4�co�A��kL0хJ+c����.�����4�C��,Q��"8�R��FX��5m��E��� $@_^ѻ�0^�qh��Y�w��d}�g�ϫ6uj��rG2\JV"A�%h����e���DJ�OQֆ��N�1���
n�X���U��6�k�p��r�{�cr������U�&�yn`nj�4�X�1��3OfSqY����1X[�N�Td=�`2��jq<�`)�*������<X:C�C�*C�|)�����#���y�N�9+�3��^ء��y� w`G (	DD��h��;�O���9���VC2{�Hi�Ǉ�Fi1�*�c6�����I���F��=�⚮������^��6˫�u84�����G���u���^���ik�#�$�~�è	���J&�ڛ����H�+k:�z�Z�s؜$��G��z�&# A��함�9��r�P��u.Z�,�!�={�j�L^���Ì�K����vR��Bd!!e�Д}�<�@����L��݈��.� <��Ll��Ћ��	Q��+:��A�+iJw{K��LŮA v�P1z���l�ՙ�ѯ�} ��&u���D2r�<r��&Ny�]���ou�?p��8�hr'B"�jPDFM��9���b�!*���7En(`ృӢ�oe�uv|ǁZ8=0�:��w�A��7���u19�P��@��0PX0E��Z:
x>u�m'he��ь�ח��[)>�Ŗ�H+�����T�@AS�}��W��
kZ�F��l�EsN��,8b,�w����b����5��_�B�Þ>}�Ȍ-+����j�z-�9�#�a�i;dc��l�x,�)�kmڢ��aS[g�v@d�j��T#�o�*���V��OS菘?OO���Î.�/�w߈�� �	�Yv �ܸ��PQ�A�\Vj_ttX�EĔ�_h�\P Ȩ�N�(�:�Yv��-�%*�O�K�U%���=��a*���U�J�͑�g#כXA�6ẍ����Z��q<��Xj��d
�^�X}� )��n����J߷(��yI1�pҔ�&J���t�W"��悿I#-���5�!d�V�Q���.) ��%2���M���q��}YD�aT=H�������[�w8
 ��-V�Ol�+;ۣ͝�N���.���e�A�n���w"˨͐�I&^6��2+t�j�O-J�:X�����$:E��I��k}(�sk�C[�S�/�9����q��w�w�P�9#��g�S��Qj��a�iSӮ�׹�Yeg���h%�C�g���`�j�*��Њ�����!�@�=3<E7mb� ��ݖy�6�ל>;sX򼡏����6��t��Z�i������a�;�����s���$gRR547�f�ቝ�޼y� l��GG�j�I`-d��Ԁ�-M]�V��S�y�RsL접�e��6RD�b�1.I�s$�e7p]��Ŋ�r,���Y�Ep�,����?�Փ�s=j���F��s��qp����c�ʂ�"Z��&D�z6gs(��֎`�3�a<�]����N�q��k}��w���$k�6�9Hļs`g��σ;�a�~	��է6
v� px�X�@�����Qv�,����}����<�m���H��M�r�o�0` =�f�6p@�yĉY��m�D��U���4����N����n�`��T��vE+H�r����eװ�ҟ�.�޺vz}9;O����`�F� �ɚ���ӘM��$]����8��MCOΖ�58�z/O���Y��4��j�'c��|���m(�z߮IM_X��<��}mS}kfo[i�f�e~$�K�"{d������8� :~DwQt۝�];�n�
�hە)�5�x�N�0emn���wV��g��3R��������$����߅/ׅՖZ��+zë��}��4q��:����)@�v�$�c��a�;�d���0� {��5�煭eƨ���.����k��rn�9Ȯj+���q'�#�,VF�23:�GQ��`-� ~�0�|�@\��m8;fC�>Ѿ�T�O����G�]�k����M������ݞ��#�Q�鍵<���.�ڿ��GMTdm�6����❎�?�@A&̡���=�]/O�iĻ���W�t:W����9�NV��e�����l��
mLL?>���ݕ�t(Nưg��t��[�t&IbCQWE�m���X4�/�jTO���m�����Q�F����K���*N���}��j�3eh�B����(���^A�^�HK����kõw��(��eψ
����X����V���^���� #O���sM��м�yy��a/��Z��0!�42F�ђ�8~���U��r���.V�4uK��f��ѷGec'H(o��v��+��-����5o�L��%̆QXI�ns�Jݖ^_��۷���ׯ�a��2�s���t܌n�>�mͭ j���R�iY��F�����UY2��GvP'�����&UR�2m�J�h{-/��N�ċ���<&eH2:"=e髇�;��������}��m�WR�<R�D�.1�����ʈ<w�	����W��";.������*�{@�y:v�GL7Qk(�	{e�A��<�¥��� �(��E���Q�̀��`�oѪ��+:Ȃ[YUP:��ĻMh=����E͡�L��^�|1͟���w*#$� �j����2J6�F��j�D%:��V�E�t]X�К��x�s�-�5�t�"���Ւc�-Bd�a���4TYni"���
H8zN2�DZ�[�®g��I�)9x�Q���h��A�V�=�����pjn�`1�Ln��]�R�:�bp�Ǡ�u�&D@wW ��7��Nc�,���QtCATت�i�&�-PeQ��cjl:��-������;�l*5�en�8b�E?O��Ȉ�Z'W��s�.���vuB���˾uxY�9� ���b�2/x��
FL�S��N����v�R���)S2�^��g�$��&K�J� +:�/)T�)9u�P#t�.+�O5��>�}��J0�d�&	�l�A��@��0�4���59�Я�̈'_����Z�����賾WVM�D�;y�t�%�=}F��׈�ak�U$�v�U���9���l&��g�-s['T>��$
6i�0I		�G�Ȁ�������;2�z��#ŷ����6���z��I�J�:� �j���k�\wg@fJ�2��s����Aa^�8 �э:��:?l'����-Z��˰�#�x�:��`Z$.�85)� ���w�&�� [�J��Xx�Q���x[�r	���������^d�e��&�l@8���[W�Ɋ��=��x���1��,X7[ɀ&�Xڦ �
X&�T���FF�'wM
O^��"�k�������l_��BS�==ĂL3M��X��f,Zz!��M���=��B���!i���Xph`_�j�
����`�re�}Su�Q��f]�g  $�Si����Þ^=Ao�m�>�Z"Y 쟑�(��L׵,a�H�	�ڟ��=o�JjMܫ����Nd7��b�ZDA�9�Rv�53N3�+4zG^�a���4&2�LmqW�sr{B �F����g߷5!�e��h Yޟ=ә�A�` /��$ �Si�����A�����V���Zf>�(��y~��������3��(�B��atg�NȌX����-��f�)qRey��=eL�"��@H��9�k'>xS�	BM3씫TDaGߗ{�gr�x���{���X7޽yGݥ�D�ߢ6}�pZ�4&L&Y=S�%�>H���!�ػ�;��cP�0���ST�Fw�)���l�o{a��#è�������^�S�[�#=��q,d� ��< �|
�p�V1�����qn�Y�'�mO� e	/\WcT��c��c�*ޅa&B#��f��B�g��X5eؔv �C~�D����J�C	�����!x����� ��
DC��$J�ɻ_!k{Iץ��}��x����o�n�Ht�(��=S��6�DI�IIW԰uH�1$�pO��kq��Wěۅ�hߖ���+��.Q�c!tܤ�=�?"��Q�A��I"�d�*��dS�pT攡�����ƭ���q�.+�P���q4T?+=|�]]��6��Du��jʗ�X���yZ��S������_�����nC�F?��8p�8�pb�v��W�D�-Ң�?I0����K�@����Ũ�;b�X&Q<5h��_�2]�\w�[�'�(R>��N�z� "e��Vg=+�#)}`�,F�0�(XVC00U[������AG����.��>�Hȩ��-$꧋VNj��؅Z@V���W(z%n�q��H� 6Nc��z[q�F+�>�嶃E�Pj�A�q�I�|��>��k}�n�$�UR��fP{�91V�H�G.���}9�srʨ����PkS��aEy���c��=5�)Г}�!n���:��������X�4eT�w�k�y�B�F4:��pڧd��,A)�U︁��<bg7i�	�:�>aN�XC� +#�<�Q�vN��]�i�x�Ac�q�=�r�&�IĘ�I��KzY�/k�x=�ʚa�m�I�Y��"�qC�4_�if�h�)�9\d7E|�8z�s��IY*��IR45��R��A�v��a�Z�n����0F`N�{"_��-�8j�H�����-m����c�c5['�ӂ�,3A@�<�β]�̱A��0y��W�k�-s��	���	Ym��q�8z�o����(�%(K��90(U��Z�`v��u!�1ƒ8���Y/������N}a�4�\m�s_�]�?YM4c�f-�-��]x�ζ�֠��ú@���,)dO�A��&��sٜ.���:X����f�g�ȹy��8�S���,��k%&u
��g1ָ� :;`nr���sgq %E���j�Ш�ox���U�vaf�F�-HQ���UT�M�ѱ�
#�����bs3�G�^�r���H� ͵F$�.�8(w���)�{��.��,���� �	��S�b(�$�N��zj�6�"UV6�)|v1�r�8q*�e�=�,��:��ʖ�H^��o�Y�]���P���}̟m6�9�,�������9X��s/t�~e0ٕ7(`�Mߧ��d���\6��n�bh����g����l`j�q�0��8�з8����^�[����D����Nك�F̀_�ų�=�Br�+a;�_����7�G��,�H\�S�E��+��bLjۺ4w�����AH�>G�������<y��@�$
��2!�K�~w���Z���arФ����	f��nn�p�h�J$gjX��@�����U�K�V$���P����V��9��^A}�^qD.K|��w��O'�����@���C���X?g��=f�>v�+MP;���T�OY�I���E{�����F"�v�N��]W����W]�Ķ&2+�������w�Y 6������	��;���2c��R�8~�9�!��rL|�~��j!IZ&5 �\K�H�`Jw=EG����A�;��=���==��٩��+ K�n9H�+�в"�Z�E��0`��~�!�iȌ��@_m�đ�h��bcW%�0�ۂ�ȷ��"ԝҙ�� υ������W(6|Y�}�h����[M
g�(|dE�玶
ؖ�����>w�)�)�A�g%������RH�>VnFY�r*��['��P�/�$��X�XH;- '�mFz��:�t�m��<��PI2�q>y�I)�ڨ�Q#7�����0G٭��=x�ȤE_�ܼ�	pw���;a'�`cy��8j�p��Ri�"Cm�c��1��s1����ܾ�*��}]��=�!ֺ���[�F�Z��{I�C{RY�t�I�/��m�^����O?2�0�.���0���m�)�md9AOA��(N���Ar�IA	���^���I��\UQPavH��)��?+!���z[��txb;H���������4reo�G>7��1PC���4w�M�X$+�Q!N��2��`�P�K�"�ta7�>k�)�f�a$��s��`ՙ�Hz'���3N�Ÿ�1�-��V]�ED�lR��[���+mzx[�GP��ߎ�z:��x8����)%I�u���t�PRQē����E�H��C8�A���m�%�L���L�*� ՙ*K��h$ou|��f	5"]S�Ԁ�:�k�ǌ�@�97jŷ�N�N����j�_,
� ����^��
���B�5=BU��]�Fr��tb@�f����G� w�a8���<�b�嚨�����Hkvw���5��d�Y>{Y?x(�I�f�T٢/��M�3��WAv`���NuQ�����}5&3�tǦ��I&ݫ�7�Q( ��L�lGND�����^�
C��=���[��4��W��>��6�G&ST6�H�Y�%e
쿲�H��s*1{��E��7�n"I1�
L�VoG��ߐ:Ids)8��0!�����^�,4F\V�S�b_Y`�,N���At�u�c��!Fw5-D~�>�� �&���Z�P����5 a�|���"�2��d�49*������H0��
䘔�4U϶��䦶V	��@V椥Fo4}��ώ��*�Y����uP �1���E���rՋʦ
���	��y�փԺI���=��@��ƃ9`��%��9i)x�2��tw\c��z@�2	�M?�c�l��7H�MY ��*��z�S94l_�9�W�k����`��>0�K��!;}��L�l�a;i5N��=�}}��%��v���H�����?*�0�g�_���,(�8�N�\����em��M���2 cGUk*��m)�Ȱ�I��'�<���a�e;s����w�p����A�$�11��e����57��?��*����mm���5	�J�=����uR��υ%4��0v:5Є�~��H�&��2��`(�[.6�Wy=� J���>������3q�����趡�2��4U9��o��c�K���5@؎�5�)�MԶ-7�Я�T�icoj��z��g��;�)��`7
��5}�:��� f�D�d��;l�����5�P��4�,'M��>��~P�s����>�����u��}`�X�,AK�S����3ٺ�eZT����8FKr��^V}P�����>���営�=��C-5f/"hV^WŎ�tD�@b�%]��,Hy|$�-2z{����|qE���c�~YЍuln���#�
�A�Fa�˂�ZO�� ;O�X�8�jl��vTT��Q�i��*E7̚�p������\2�cYh����*�q�
�\�<����0�|e�hŖF1� ]9j
���A w 
�"�Tz�aB�3S 7��ݿvl���WF�������R�[�8;��7|Htab`���Z\jbC���袒�@j�0��D�3W՗hVH�8_V�
��D.ψ��0��Л�+ �ݠa@���1)�"��k��j�W��Y�Б��I���S�2Sѡ�>�}��R���b�,�ɢ �B�Pt��㔴N��O���T��:��Dk�ٌ��A�w5����?l]�C��3�����5PP�{/Qf(',T���c��-r{6�y{=N���%�y���ٙ�1`W\ =K۳���\Mu5�qw���F�Y� �e��dS#{IR�c@� ?QT/��4
�gES̷�E�S��G����&�Ze��a �GmI��ym�����I�[HZh�g�s#&�M�-T,�k�ZF��)�?0�h �F�b6�Fx��u��J�$Fܘ�}aE>�����\3��sp�1�4;:$z(�;��\Ly�%�fR��"��$ѥ/:9��Q�e�������+S �ya����tA"{�&yG.˽.��a��O�\�e�����4��f7"��d�X]PI楥Yn60�3���&fV�3�N����}A��+ %��A�-8�`QO�]fI���:���3{#�u��[�ɲ�K/�5
���փc02K����k^C���1 �9�T�N���˴�7�
�>9���5��Z���ըlZ�Eg���SvCP ���IҲb-i�P"K�2�Sz6�T�>�K�2v���f!���ҫׯug������d�����Z����� ;����8��Ng�����*�+u��%,��� ѧ�kr�U&JA�+�悿��8�s�ZvJ_碸}Mٱ� ��o	�d٩*�W�N�:$��p��S�`�:���)�'�OA��,f]g@��d���L�lizY��e�7�P�cʞ*!�Xl�	5���>2F�w��ڿ9T۔�i'�Zn�ڭ�������{.��c}�;3G��2�.�, C<�g�����fqt�����m~��Nq�s���L���t����-���� �S�#q�Z����%^Y����;u�����i�ֿI� ���R�e,�W�ۦ^��7����qګ-(;�����9��ϑu�h���Pg�S�&GµΗ ;�o�bu�\^��x�Gc�Pk�37tLx�/m3v =��^u���k�s��S;�K^��@3�bhJ	�ʢ��=�����%��O�T�&5���[Al������Cع����{v#LV�7�� l͝Aܫ:X�Vn�s�������®+�;0��ݏlF�N켋Z��hl#R����n�M>�iH�[���FY�֪`��]�y��݈5ۏC�6wi�U<�[�0�7}�i����JT0���}R&���U�WuR�vJ�4��%�5NL��Tз\������ݬ��{��Z���)I��wc�: �3x@,@�����6�ȠΤL�>H���AC����������c�vR�vk	���3����2S,X���Y�J�PB� �� �i�tN�IO�}�ۏ�����;邃���m^�/ۛoʼV0Z�  ��aG��GֵO����9y�<ن��� ��'�9(Y�[�raJ(1�q2z��G��x��C�<���JG���.�&�#퇅������f��Z�
��^vy��z⁻,NטB	����)yuu͝����\\�Vwp��=P�)&���"�i�K�1��w���N���m����'��al�ϊ�c�1�Ô�������Rf�7\�d��f��(xc�M�w��^��:Y:���q�[qt���J�qZ��#�_ ��g@tUr�rC�t׍�z��L'IWQg�Ph��	ŕ������p������gL�@�D4���?�O����'نNו��ZG-��-Uj6�Dy���.��"�f8�>�`�Y���"���/�$:��'�qТ���H1_^�q�l	l���	�kK���	ѐ�~�~�~uMW������@V�J�ם�ڨ{�)�N�Է�I�67�K)�/H�����t�=ck�wv x��,���SP����7q��G�b����)h�^pc�z���"�#X�%*�4<7R�hǫ�g�-��G7��/�}k~���E��������"�B�GÒ5���85`��ܰ����k	��6ߡF|�Z'��`u.�u���B!U�?KC'��5K�rg��:�1��>���;�d^ń�L�&�w \T#�S
���Rc�ԩ'���v�`b�T�f�~�_̡
�l�3��`K�#�uk`�C�bAϮ�u*o�K��ۘZY����n�de;h~����eN�
j�yB5�P�H�d��Q���78���iL�Ѵ�;MK����Tȧ29�V�K�DP�d@���6K��B@2KOa*�!뮉=�.�%L.V�G�#-��e"^��R�)p�æ5�XEk�y�ة ��;x���~��č�\�,�� �^����kz����4jSx4�E�yb�5e9]Z`g�\pDq�t6aEJ�?�#=�/v�4��N�uq�b�U��<���zo�o��|^�ƲAw�$XJ0v=�fV��SUEY1kJ�E��|��A�v��9��������Ѯѹ��Q�5֩ �@Y��Y
ґEa���X��o�r�܈xKZ���={*y�>��-MîQ��!�_y=�kveѻ��9Km��=��:Jd`��9x: 6��9�N������;]��ּ��!࠮�Uyi��V��  �ِ�a�h��e�e2ޖ� �/,�HΌ�׽�;��-
aX�n3���V�"�[��Es�nB��A
�N*����+���;Q����'Y'Em3ɳ�GM���9Tٜ s,�O:�I�qM�r*n��K�i�{��U�;[�dNLMmBaǬ�o M4P�ar�S:�(�Ф�n����o���|����o�Ωl��L���'������t�Q�F��Iv�m'�\��#�WA����	#o�nz��UYd$ !�w���~Ie&��ʺ�����4�צ�)S��~ֺ���n?l����e)��l�����&�qI�h&���*J���ܙy������{g��v۲$��Z �˳DT���U��* �ˉ',I�䷯�b��3TdR��g��S�z�Y��Î5���󚉼,�w�س؏ |f�ti��x����sY�G".��aW��ȓ�*�ɡ#��	��դ��gu��,����<���`�IWO�Sb��_nE���O��[�ϖ(���X������=��wf���7S�іi���k�0����Y�<�gG]>]W3���/��Sc��_>�ْ���]<y���������p�F���Z�C*�xL/ vj ��W`]pR��C����9�7:�A ѝ��	#��>ʺ(��S:�A=��@X:\����9�^�ݕ�$�t�fw�^�=[0�Ƅb�C��)�6=��9-@>�Q��G�F5tn(i��s�A0È�"�w��i������	��h��p����gV�ϫl!�~O;��dV6>"�Q+K^�H����/phP�ƵGk��'��O�	�^9�/I'�e� ^�h&`�tb�`��S�:��"M�h&b�g�p�/��o��o��-�����41�K�ժ�d6D 8n!�]C��=�q���?���	��Z��ܜ�~�g�ݙ����ai��b��-+V`5���-D���1US���>u��r����&]�\뚺�j�v7��>*`\ݏ�n��o���/����׭,2TV���L`��(7m���g��� ���1�����Fn;�]aOs'���V0.�.@N���3� *��@u��I�*Kh���EBQRc#QCǢ����bdk�7���~�P�:��Ц`���_�	�"���www�����5���o�^X�$�V���������c�G�@$��zeLԊ׳���k��޶4�����Yv�8�!�
��{S{��n���W�0�JLF��H�� �e5G��30�‵^z���K�5�-��dn�Dp<h�bv`l�+���t:�i�M�u^i�*� �k��y��/D�Y��i`�tK"Z�n� W`��/���ϱ�dB\�����V�����:e]���'�C^@+>�.�GNj{Y�^����R���Z���Τ_��MB�f*��;_����i0�.�o�ر]�"�+���j��jh��*a���4e���_`�mA�h���LkBw�����*]^\ؙ�ka��R���ц���3�;}QA=�,
SVP�6�B���d��>;8yV"�6�N�&���>���TDP(�b�ҏ
`�8�V��!��i)�L�y� ���^bA��;Y!$�LJ߂�e
O����	]��ذ��+E�I���8'�NY�g�3%p��n��b�r��b���t��Z�u(���˭��l�%��'p$�Mw��TαWFiP��S+g�vb�c��v������r$`j�9�]� ���Wq�;�q�=_��A{!�Ӿ[�qvv�G��*w������
(H��[��R.� �b����Te�^C��u=ˍ)6y��&y{�̼��%��T�.L���/?�������Qs���^���ͥMaSyd^��$}��m�GRjE4U�Kzk�n��H��kf��t2�0�>�9/�Z�ů�#���`�ڀ�v�����}���h�[�	����8 L�Yŝ��@�`��C���[��5L,�Of`4�&�MZ�K�P�����v��1R}:x��'���8l�q:s�v���ӱ=�ٹao����b�0�xB~
 ~�����n`�Gk%�*j��Gn͔>1�6��-v����f���9��T�G>s
��گFa#�@�	MK��[K���d�oJjb���w�5K����MTg溙9`j`�� ��q�7@�Ӕ�R�LT`'C�{n�n���;�����c:֜��������:����hR���VZUX7�%	Ɯ'1�����{k��X�������Z\7�j���{]��r������}���!�Qڵð�$_��Ϣ^*$_��Sc��d��%О��R'�*������ק	�A�vW���KHT�o��yf��A����-Ph@�%�6��������ӎ�6���^_�̰� ��F��6o��O_�B"b,"�@�U z����O{����٦�f����g/<6����X�Yq"��J(Z(�}��A;�,F��7�2�*�E�h�m�и�t�#G8��`#[/Eoz�D�����C�	�jM���)�(8�o	l��I&[j���h�"@#��u�Ń�P*�x1�}�D;_O��G�W���Z��I�m�&�\]^3Y����������y�k�w��+3�N�z���(�,��J<5m��5#i��Ϸ{Ġ��8�ʼA����K+�(N�R�85�*E/�q��	Ǌ�rH��ld�=^%�7MѦ���:�e9�E��H}��i@���_�3�+��;11kN(�s�1P�0�V���,D�7�(>�"�e5��N^GN�~�e[����is�Cv���3;���j���Dqe]�	����Z�At#�#�SJk&O�e��'u�W�F��h`/bTd��+P��yj�>�j��X�2o0O�Hp�m%�Ț'o`��J�xEjDRk%X2S>�ڨ���Ǫ�TN�O�� ��itNh(�P�7����ө�}\LD������Y���i 
&l��$/i}&'��<�s M$81�NΓ���Vؠ�3�q��4�˼0,"���WWl�������C������=3~�r,��RɊ��dm���<Zз#c(�G�W0��^ b�\ �ONQq`�t�vMx{�Hx$��Ym�4��}�������b�q:�r5�� ��H�����B�^y]+[} t��M)���-y��<|��v��e����cI����4�nn)��+�5�L��ξb������5��j�*�����d* )x6��53�>����[Xy��c��K�l0!"_i�ҟE3ۉ��5����8���n�0�(���	�Onx�:';*��Ӧ�7V�Y/�T�4��Y,I@/����1��g�=� � �1��]��Xe��M�sn�L�y9��1�q��sjB��3�eq�{cό���������֝ca�_��X��	����	���mfx��M�kk��)�/u���,��k���悾S� ���Z�q��1m�V�7��8m Y�O�3�P\��9�<#&����Ж޹�L�1`�{����`t �����lź�y���#
�������8�6w.��/5���S	�ph@o��r�d8��m5�� ´�Ľ�b#���v%L���ۑ�[��'���|����4����#6"�Ϻ[�X�����q\?��Pk jO��#W�{ ��Fs�"vDČn'��a+JnZ�e�Q��	�:R�rn��1�����jS��X�����1��b%��Fᶸ]������K �cB��3��6Q�\dk�#���q��t۞���� q^��n��k}I~��0l���1˼z�����C�/����A�i�.To�6c�Sr�'�1ڻ���vaZ�Ij��(lE�0��3g��遌k�:G!X���m����ް]���%���_ү���,���Y�΄�V�&���q���4`'Y^��3)NQ*X�|�yL��wRl���L���%m�D��ag�4�e�hQ��S�ǈ�z���a6��}z��I�0H����ʹ��V�����鯿�-���D�.�/����?�HD�	�m=D��E/36��i�i_,Сp2�bDg��c^� 75�'���>]__��<�B3U�a��ǯ�!>q4*�q��+�@���Am"u�^�H�侸�9��cj4A��4jb2V����2�s��?������Վ/	���� ���z?��>�6�]����Ǘ�T��Ғ�N�~�����QV�;�
g;3�����:A�4����(�٬�Y����uz=�Us��_�KP�~��tDϱ�r{�ʆ�نY��bѺd��딜�)ID��
Ѩ��qX8�#ع�\������¯�>�Ͽ}b���2u4�lJK+�'��1E,F��0�0]8��Ϫﭸo�V��}�N��6�a�|c%OEѥ��*�s������9��b�Rq �iT��g��1�q>��� g�Z~�	��]*��U������d�$�L�� vT-;�;CE��6�����h8���S��Gu����(��z������v��ͩ93���za[T����j
���3+��=
1��:�J�f�X�	���"� ђ�IȾ��l�Y \�TPLG/��w�D���3�\�=̙Tz�1��ɂ�bA�S�y/�m��#�����Ős?X����<&ᴖ*�ZNmJY
��鮞ž�{��&uM��vv[��Pљ�������1�����w�u�=������+�����\�X����&1�����`hh_o �;!Yx�dGNo�A���u�m��'.�䐨f6����-�lQڥ(?79蟬g��#�=u� �W�c"��M�� S�v�-���|�v�[��!���L���qb��942QT�ه8Q����'ګ�w�Jc`�1X�ګ�5<�S�-��þ�A��3F^�ܰ�Fd��/�(e�M#(%F�M�#f&F�����u���X@�"�Ԫ�A|�$�v��"@~�:2�����Q]o�#+@(�q��[��9T��gr.z�
�`" ��':i.Ņ�Q�/���V3�r1�{^�k������H:�`\#��h�� ^,�P<�.7�����.7-��7L����,1�O쟰a��W�	�<i)4�WS�$-L��j�\��p�N6����C�k֙�DO$��8�)Bl�ؘ4��0�G���bC��U@���S4�P�R��"�����&MZ��V;Pa�';5}��A?����	��{YK��,I)>cyi,�5�l�d�_A��&��^�!b<��ס؅�G0��([S){o`O��MYץߪ��B���;2;`�P�}~x��rqцr�'�X%��ja
P���b�1p��d�!.z��H��H�F�د �F]�@�h;ĳ���0�u�&����o��d�-f��úF�jd/Zp��dP��kݦ��܏*:�.��Z�����dT�������`��Q*�ZOF�)S�^�g���snSV�C�lR�eKt�N|)���E��u�T�ҔF�.ȩ����{4�8��k�\9����-��=�)� z�|��r֞�>��!@n�5���?g�|H $�((�wAP�M��lS|��M�F(�I?/�>�$[��jo������L)4<��?�� ���|�g�VJ2�=C~�<�)��kE>p�Q��"w���vw�xi��Ko��7 ��g�B�Й��+���ݻ;J���bo����������^�Ц�ߵ��S A�?�?�f���Scp=�����NG�@A��
�~�k0�z8^�F��¶�X�케P������N]D�;�F-�:��3U������s6�;X���P�o� � x��j0_���ɋc³(q�a=��_4�]�8Z9�LJ�t���1��]�0Me����\�C=T>>?�N���g���������G3���L�G8(& ؤ����<`��]s����՗���?��$â�R��+�	9*
Lp=�g��NF3�~���dY�;�T|�@�]��V=�N���42u]c��tx����=<�Y����ݻn~�7p�� ���ȡ$���
��Y�l0���AC�瀴� ������&�W�q�X���:���������k}�s��L�c"��N�**��]�#����nNV;��F��oE��Clc/��G|��Is�_Z1lNN*jk�a�B'Z�,�Öd�מ�]��V�L��������<�nF	Woi\)�V��N�˨P|���=8�hRKPd+�k�ޭ})���E����A�tP�	h|�������p�xl������3���,����Y� 6�ל����Jb��ҜG�ԓ��Р@P�����pf�F;.��:U� �ȑn��7jK��Y����곸�^�*���6�^�r*��R%��䖮��#�Ͳl'����!�Ȱ�4�p���./g ;��5��B�%��D�c���g𰏳��� O��h��*gZ7AW&��*���Lc�̭Bc����a��P7�-��^P��+g
6ObgP�a���`�� w�jLt$dHd�Y�������gd\�%َ��0�e��UL�x�l���N��e8��mX�;A�4�@�#Eg1��h��zk�ud�B����:���i�sD,CJQ��6�)��8Ϝ�%N:�)���sI�.oS��Kp��v��O���`�$On�~jh��+���#�L�?��<��u�Kc댬���*�@������]$p����[$��E�E-UJ�Q�\�/���ݱ��3��y�V�5��.l�Y�� \��,�-)�vK�Z��-t��m3Ӕ�T�	[�^��JXb%��F�3��|�JI��`��a�s�
}� j��V����vh>ЗN��uwn'�
Tc���E!Ai�_1�1�5jљ�]Au��-,���h�)��]�ɬ�ی�� ����Lc��p����&�&�Z㡖��t��Q�:��V$Z���C�oqb>��d���bE ��4yӒ�4 1�4�jY�x�X��$��g0"B  � 1����	�Y�-lj�`<�f�p�����F\ª��z��F�wd���@5(Qc+r��y,���������%
W��%5�g���knW��V-��Ņ ��f�s8 �/�	ZǶ��[9ᗢ��1��	F�����>Vj)�-eтi�f �H�� �8D�'�}�Z���������e�@I ��Q�s�jퟓ
R�
͕���W�=^����׿11M���jim{����Se"$}��J_���}�q_�K�s� ��d�?�b������0���.0w�ӆ��"��
Ѣ�X�Il�#�*"���Խ-!h��ǱG�\�Eۯ��C�j/���.�R.4���8��Sj�k�>[��G�b��Shx�D?Xb��C&��Vw �L߻`��y8~���&�5 I�H�NNO��v�k�8�`��M,��.��(zt��
�nC��e����駿��}���������L��-
wkf�7�X�E?Z��]byD;i�߄̉ڔ�ޣrH~� 3	(KD���G�B�y�`�B;^����F;����F�.j��E�����ƾ��~|~J_�?�9^_i:��b�Bkr��7�w���T7}����/��xx�f^�6��LU%-���E�`�������F%W���-����#U�a��|�̖���'�� 1�}��;�/���֑R�@؛�,Tɹ��I����(�^^�ơC��7�� `u�{2S��!~��������b��0���VT�%�� �#���u���$�W�Є&O�R>���Z���M�d�Voru\ �B�$`B
��� &��Kp���E�p"G�ki����z=�غ�!_�y}��՗G�}ȡ�)9m��"�SC�����nL����)@�g�(!�ІSQ��M['�U �Q��v] ;a���+8��5�0�M��8a"B¥HD^O{���
���MF�����z+l�)0sQA_�DT�;?#R�fg�8�>$K��f��JpjtR��uEr��>Pm�SkmX���C�$0�vtd�q��x�>�����*J<SA+�����>�Hhi!�o���hPr�[L�,���T$��[tn���@��F���u��sy�g�Ǎ�G�U�f��[�Z��cҴ��m�)��AeE�`9��A��UGJs��g.U� v��m�,��3���Jg�˄:6�J��rw��S����(v�RU�T��� �W|�R�$��ͦU?<Aq]��*F�7�������i\Zf�.�,�,�}h��7-8�Pi��r]k'��[ׂsRe˹�m]���@��I{�U\z���B� >���38��S�
�HKn�dF��\��z�q�h��Вcͩ4��U�hX�q:���5�����3�;��)��X����;��H��. � ����:c�RiFR�v�иR<B�q��qT�O,��[u?�'Z�x�G.�-$X'�tRrnu��v��ܦ#�Ib��G��B~!&&�����b��t�9ڿF���.�u�u����AQ�yl����̟�$B����g��h�ĵow��V0�������h���~X�B�Pg0�fz�_�κ&��naI,
t�BvSh"���>�a��y17k-	"´%�j���NS�� wrV��69�	��e-D�- ��dVm��v��WǱ%�Ѻ/ݓ��@F�����V���Y41�|��ZdvJ�����X4֥al�K+~� x�q��溸(�^�w�h�A%�ٛŴ#�c+�ĸ��Uz�ج˶���;yӺ��|��l!�f�B���`���~!��/%�-A ;�ߧ�?~'��� ٨�8�8���X�sI����m9�j>$���'�@��Mb���zS�������uM{� ��t�+M놢
�t@Ӵ��5{3-���C�_���gŌ���О��6�_3�q]܏lq�܊��W�~���g�V*O���lW{�Zj��,2��.����y�%-�L��|#�`vn6׋x,`�\ u�������F쏬��A[<�'�LQ��/��O��6��Wq}�߱ߣ��;|�{R#ʽ'{�'(�ؙ��G=�g����3����(�}������f�����D���~-��� Iw� ����m��߹��������/~�oy]���Ί�ː�h ���G�Ɔ���+�*cЀ!PX�] `��O���������_���%���/�\�����L��b;�7��������-��_KZ�;WNY� \���D��	�g�O==?�Gt=ߤ�����#6Vx�<9�q<[��x[�Yxى�_������)=�<�v0tRqX�ϼh�u��9��n�P��aѿ�Y�و$`�H$�
��80P�WV��m�����L�� ��F�X��O?�H�M�l����yP�|0q��F4LT�kRC� �n��[�!��b8u�i�jlb=�ނb�XD�mf���=�hm�V�pB��H�!ZZ�� A2z�
�ӕ5�A���?0�V��}wun��A������s����Rڀc:���[_���\ �5Ri�>29ҼL��	u��b�nn��j���c8�tzR�;�L����@�P0`����ST�Sd $��sZ@�8�+@o������W��J����6�'9(~?w���	^݂�κ��{���S�&���$_t�.�M���bZ���h7�ZϞ���4]��a��vf� I��Fi,+�^5:xZ�$/.4��w��H;O�
*�z�h��w���]V"�zˎ�����`^�e���J� �m^X �߱�Z�3D�D���8�N`�A��Y�Bx6G��2�'��73�R;��~��Č�p��LR2�ܚz`��wP&Q\��k�MjE+9��uLJVc�gd����ZG�����+��jo�:�ޜ����!Q}�iU��}"�*Q��x[k��6���=�J��u��7��*��^$� EZ%z����"
q� S�CZ{*�g Μ�IP���ߎ:����k�7��K�����e�������"�>�,�Q�1��1}�3�5?�hZ���4���/dCY%f�P,���61��Ǫ�`ّ�������t�`df'%�`�N#�9Y%E���朶UuB��z?�D+H��G;w�c.�Z8���F���5�	S��O�1�lk�H�Ͼ�=G����]5pM��I  ��8���	�G�t]��iI&ܚ�4��R,�g�u��7+�e��2y�$��yn�-6�I&|�L��m��#C�|^@�U�E-�g��/:% �|��	�Q����:�qB��299�W��������XK�^ܦ��[����h�,,_�܃��wÕ�Eо��4H��>N-���q+'l��8�`�}���
9���լӡ�Ad�/d�R�K�<��#�%�>�ڟoZsʢa�v��v陬E��?�,.���F͞>�K����0�V�d �%�������(����|�=&�����|}�c�=��d`��& ����dSp^�(9pɁ)�d �,�Ͻ��5}��S�|�����:h�Acҳ%Օ�3�t�`�P�e�!&��}���Yر`vlKޠ˷$3��R�����������5���5뇞O�4��.�'��Z=��&�l���IH�I�l2</����1��v[Ǵ̵��L,���l�=�7�V$Y��@pgk�m@������;;��5য়M�)Z�CX���n��⵴3@�F.宍�q��yO��$��خ3(��z3r�T.�^�3�X�)YFgM�/�C��nÎ1Lo�6��fH�F�zIn!��ýY�,JV.�4���C;���&����VY���k��9���6 ��.�уy�,֓���P������ς�K�>��>~Lۋz����_�������5���`/�����u��.�s��5�"�g_͗5�������Q�����l�݆��a�%Q]־��2�|.mc\!Tۤ�~�DR�q��ww�|��sx��^� z&)A�A�*��J�9]hn:ɨMCpg�d�DNdր6t ��A��-��W�P�ݏ?��A�5�:��->���%�恽g�_�PY2h�i�(��m�i��Q{S�h8yMP����3X��^M�*�eO��uU߼�0�pHj�]T�U����4ʣe�T������(�����J�@���7N>XGt%�������ňS�p�pvЩiHu=/�1�7���ZzW�7�B���%}H��'2�ؖ�J6)����4� vP�{;`�-k�>��u����
��}���0�p������=�5*��֚I/ȹ��y_Z�djb��̐�yCT̮�w�XiD���2�H� �q�@�I).�3�`J�.W�w7�3�n�I4UP�W�РB7=;�C���PSh�>���6ѣ����"��T��}��C�m���q7X����@t3ή�j��,
��i�=%�$�&d�Ԛ������"41"Hursv�C��n+aY�Hu&@�U�+eV����K���t��8/Im<����@NY�g�+����*X1�-��*c��.��{7z���f��#��op
A�/P��l�3Þ�͞fW�Y9om��y����x�)���m
���}Oܓ�@���]�O���2��ζ�U�=a��hS�U��DZ �D�Eg���"�	p����>&,ֵ˪2�8GA��ﳿܔ�
���tBp?�qZ�Ɂ5ڲ~��0T�j��{��������#���E�&V�m��mi������4�\5$�b�{V��9�e��!|{���Xe�=G
���q�~|�����b��h�������o�����[��\
6�*�f�gG��"pԛ)��LT��.��D�6/w�Y�_�lύYA�Z���1�ef��:�!�1@Lf�t4�k����b���� �ɜ�]�(3�s�5[1��d��¼�;�gŜ�q�d��Lsv�=yS�Ń�ya�H;�}q�k�WK�[��r�¦�A1Xf%�N$
O~8+xmXE�xB�}��f#v`h�P#� `���*��J�]\X�s`��+��0[��Ojr3�3m�D��� ul�V��V��ΊQ��ȐN��1M�u.)
f����4�쥳����z���d&]��@�Ś��#�o�>MK��/��y��ѩ�g5xr[�-Ov��ky5\
�}��=����sz~y�$ϫ|S�t˶G��fc�	
�������n�W�=�E����=�,�8��Cb�q=κBN�MT��$��q�cK܋�s���='�.�8S�l���:o[T���vD~���M`�pߞ	���hhp r
_�Κ�bs%��ͩ�Z(�[��
s囗�������C{���"m��̚��`��.��A�_v[��v��<���r�qfɜ[��#���asxgv�X�~2k��-o�N�~��s��
�X��i^ƊGn '�hq�>t��s����yl�L/�����f607t��9/��{K�Cpb<9+?L�˨�Fy�χh{�M���v}�)���`�WE��b�b�0�gv]����m����O���Z��c���WNU�, =�\8FN6s�M�җ�5-� <�c��"��q���c
�wr���πY���tqY��z�n�n�ͻ�V� ��i��~���� �ћ�Z��z�8F|��(�_jl�aK��|��ܜ���恆-�`H���-�T���N���)��'���Jrsv`����6J���S3Mg�H�v�<�"��k�Rn7��������¹/�%=L%�h{�F�,�N�C�q�u�%罚~0��JHv�}��#�.��فa�e�ّ��3� p4��:5҆�S�V'/�f����r�V@�������/ڗDCYføFYcJFT������A���J��4Lu��.������vH�RFu/���w� (^s/-�� ��z������n���fuⴶ����},�9�,=�P��R��f���ZC/����,"�bBY����F�H�)wqu����
0��+�2ILW"٥&i�V�� )� ��g�]���\OY���\S���d�xh�>{�M�nާ+ ������<?������t;��&� �D�K�I�>��`�BZ)����Y�a{/�j0�ݻw�Ç����ӧO��G�N�um�˳E݁'�5&������(�v�
0�m��g����N(��*	����~��,$y8.N�z眞�Z�['C'5PG�Ԓ��띫C��H{BaR-�A�w;Q�r��2rv�������B�W;ia����5[��=����/���w�����ov�Z!�$:x�jl�(�J��{�����v�ypz��T�bx���Y@�,vZ-�\WW��C@��qT���Z��:�x0����S�T��k�T����K?�XAqy�SX��䉆�7�M
P���	�_^K/���tn���Ӏ�>/Z6����Nۭ&����A�876.�<���6���Txޗ|L�9��|��v|�a���1Df�v�R��>ҙz��u�ّ������g��)�������d��-�^�����k�����o8aI���6c$��Q��A���&Y��&W\�(�	k�QZ�z[���8������couy2�!V�[tq-��>���`[�g�作��aP[�oIG��w����C�I W�8C���I`#*���L�:ŔV��~�;8#;@ީ[ ߲�[<�6j7?H/2c*�� �8���SN�,jY�X�E0ͱѣZ~��4L���\l��$��BŊ���|4B�t!�;�$�9L�[7��5XR<4�D�9㾫׏b�M��ٽ[O(r@�� ��3�N�%���>R�Cj���
>�Zb@cJ԰��^Q�������t��ҲT�V-ڎl�Z 3�g�U-�S�$qǄ�L�}}o����:|ysŮ��ŗf��k�K�۩5/ڵh�r2J��Ù{S{Ԣ�Lɒݙ / ���lRn�b�&#&@��l�U�N�p�k����ԫ��߭~6`$�����Y�l�p]�=����i��,���,0�?�-��d]��}�M��\%��5�Bd���I߰u��,�9E��t��F��|�b?f�g����yy��5y�^$�1N	1J~;�ALk�Ms�>�8����<d�=�3`�k�� ��l=���]�f;�n��Ĉ� ��'��q�K��^Ņ�fj�q
��Q���
�f�W�Bi]g�}3�&�f;+�9D��hR���*��$���"[����J�+�h�j��ڃ����AS����I�.ߥ���k��Ͽ�_��3ul9ā����$$�;r�B\No?Hm���^�����V�y6绀=����}k��7K^��Cz|zN�Ϗ����ÿ�8�y��A��R�g�$R�7f�wf�u2����D�]�8\�N�������.��|s��+P���:8��*�Z�լ�hPuLo��Ue!-�N΋����^�t��g�� #�}�&�h�hF�s�����J*Ř6W�^4H�!��3�ѠŔ�^?I�FS	S<�]l.��h':w[�و|��u�#����� vb\7)ޝ��� ��^Mx9�}���6Z!��M �W�R�2��p���}L5Z�.ڑ֕���?pJ n��i� �+�S>���m*�)����a컠c�o��d����m.����!\�����Z;1�'ZR�}@��+��9 �m�ޞ�����$fT�'5{jZ�_��t�#3L,�<�>y�UUEA5������+h���%�w�s�Gv�*�Ty�,�r�dH������Ң�@I�o��߂;��,� wJ�.�����斏���3{̧9��������1�]��3�y��3(ԫ��������d�5&cB��)�[���_?���@�Ě��grt�K��`A��l�M���ـ�*���:��������G:�P���T�OGA�Q�<��`m��~�X�G�>8�]X+��+x���(#e����K
��N����\v�W�w��~�u=��rn�U�~�{��A5�2��2|}��o�?�[��᷽�ٙ�ws� q�V�9�	I�Ep���̇��/�d������8b�݋I�n�&*��}h�����w�H���V�?��Z[�`�M��.k�x���$]�}��w?�O5�9פJX��3)N86��L�2��.�T��4���Zs�a{cn��vqq�Dq@���Y5�'7xf �О��r�:0�D&P�I;.І���� �(&^5f�7�p������Z"�h��D]��h�L� ��i.�����˲�%��g�ɧ���G�/� u�a�d�4��rxyM��=��kn��g�aSTCC���CZ��8grE�����C��Ъ ��L�� y
&c��&���S�j�۴V����!��XP ����@[�����y��L���"��e���(>i�����f�;����F�JO�:%C��/�Hl� �uy�ʝ@�*�G#&�D�M:mN�i�G:�W_�����0��${Zc�n�sM�$�W� 71���/��I��pɢ� �̈́C�+@��B·cҿ�m�~-���;ш剏�A�� qJ���k�+�o������ۋ�%f�hl�V����Uӌ�ІLX��A��U�]�߾wl�����������f��M)b�$&����X	:p�����c#�i	�C�������;�.��ǆ�~�6������]|��B��vp� ���k�P�3� �hj�V"�e�L�L����m�Y �u!���N�}�Bs]A�s�W��V��?��{����_���7��>�XC��6Һo�a����s64#�ޭ�]�B�<[Kά�v9��
��'0�����A72��[f���l����O�o�Dӣ�溮����:��8���&�=����|�kY��@o�+ҳ,m"�~��-Cm�N�?x�a�pg`�"�3�ݮ�E�y*9@�Y!��WW��7|YD��"_��)�mӁ͍3�-��8b�k
� ۟���k!��5��L�Y����oš �R�-6s�]���i��6��������?���}W�!}��5���������[z��(fV����=����Q�')�+l&�¯���Ⱍ&u,����O�O�m�҅�r![[�2ϯ/:�z��F�K�2����8I�"�Q��Y97��2�@�1��=���t���N�0G��F��l�4��kq�	�(OJ��#H.����� �XO1��)��9�y̢Ÿ�h��}3.+8�lv��B�:���D��G�்}��3�U(��R8|1`p���i%d��:��ϫ��KD��U	�m:Qg��|�:p��Ytܨ��,6�΂lG_rl
ЕN�[�\|�Fz�P�A��
Ed���H��R-�bY9�,���H���j�|��=��\PT1�rb�����싄��Ĉbu�ISW(:�m}(�B�	
���eﾥ�}{�׽���Es�-��́�
�J��
�SG���7��[�tz��qv��5mC��^}��r���F����SB�'Ө�qKG_�
��˛tw��t`�=߿и���͆L�w7��{}����0 Q:��y�d{�3���C����k�dTA&�?��A�}�[U v^�.��7�~Ga���t�#_����oTuBk� �'7zK���>����]aЂ �/d�\P�����ӯ����+�Ӧ�X���!1�=)�ACZ����^ZpO�nT�GM*�~�����\_�?��=���D�c��jP5�H@	�f\��������>k>{��<����͋�(�=�<�k����I��"�J��D!�_�P��t�[�XU��F�{����@`Ȧ�B.kj���Suȟ��^ꞛm�h��l'+���Ȃ}�$E�!�	Gb�
0��á�pw�.���cp�Ps<���9H�s�W��_7���a��R_:>g }޼�/��k�) (��/�[���2�$��U'�{]�u8�lE&��� D�b��nG�?*���cOJ�DH�p�8�3P�Y�}�k$(�,�I�<���4Zv�!�;n�
�������~u
s���g�綮�K��&�����c}�����-����8�)���7_-O� D�4�Ys�{z��B��R怑J���|���Q����������t������n�$�*Îj̳XT�6D�ͮţyD<��䥂���Zm�#�Cn@�~c�� ��06�
�D5��A�v�k�~J��GN��M�v\�s�9�f�ݦ��b�Iw�6#ݛ�^j��1���p3�~K�djz#��a�����ҳ��@+�&�� ��}��iqI�H/T��w���_~�[y�����n�[�E&�u� ����|wM&hcD�c����W"6B�:ه�r�-���-��X��U\�uZKߛ$�@f 8d%���1�y�����b*��!k"+�'I�j��\q�[l�5Bk)��ͥ]��g��xV`y����#�1��5A�^���b��-������#l&ۀ�uXX��-_��'��\t�?���*�T���ʀ@�D�Y1q��}�^�gOh�~�Z�g6�/c1۪�g���:��z�, �c�;�����E���͜�k����ڳG���/�֊�8X�a2K�_�b�	����X�QL=��1'��+&TN��k�<��6^͎���U@���~�M�]��)���HK��T�=���C=?H���Ū��چ�
��cЎ�1����ȅ������K�\jg��[�韭��熘׻�x�p'�����1�D�HPl�D��;�cy����%����l?n�$�mª�&wm�b�u�h�Zj\l�"����5H��w��V	LM0�l��3i OL�s*��h-z��9n��E���� �w (/�(!���i�������n�5D�e�.-�r,K~�ъ��^b�4��5�b��Z _�Vg:-qv�}GNN�����o��)=<��{�����(]��f�VЎ������C&_x���3�w��;��:�<oo���5h�ru�t�����ΫC_Z���z3���<�TG6LuPn�F��f`dRMC���Hs���E�������ݣ'���!����VI��h��pᧈ��(i�ṉv9X2]�nCw/�@����zU$�p�c ;�#"����k9DZ��/N����J��
膖؅�3u	�0��jB��4����!2��.fX<���D0����©���J<F���������T�R���u'�+�:�-�od�w�-W�Z�k���v��>��3�W��m���"�蕶��@��K��̕ ����$�(��4]��uh^��uM [�N4�Y��g'�[s@?FRzsq-���;��>��@���G��
�MT�޿�@�H���C���K꟞���L��;�M�`<6W��֩s ���;3.f��e�����N 
��Uа�k���P��Ġ����Qo�Ǐ�mM��n��kU$��aL��^� d���^�Y�Ƞ������	����=������5d�	~����?����fu]���˨p���M7�3Щ��#��	RO���=��BT?Ikg��΃&"P�����2`l�p[���u/�~�'���-��$KEc9Ϲ��S�ڸ[�d�n|U��]�Մ-Y�/���Q����%=�?R���h�e�j�Ʀ�ޓ�zk��Ms�z.eje9G<�]]+L{s���:X��Mx�������3xyyN�T�@��A��m�p���rp�����&�YϞf���������9�D�BX���M�Ǥ.[\�!��[V`�끩%��������d�vy�v׫tuu��n��̶be�$`q�0�@�-�)D��[�أ��,[ӫx �jW�%�'T�ono��U��*�H�KV��^���
Q8Ii���m��C3�o�yk=������� PI��I��з�Y�D"��_Q�Mi��q�������T5�	PU�S�Lz F�xT߃��xJd�{&٠x��)��%ș��}��<ͭ=w�=!� �&���Y$3�)���?�){
��*ƺ�V�k?,m�Ib��x**� �|�:K�g���i�.(�邭���J.)����4���X��=�̎�����&59���v�-X}���{�4s 2��_���#�<�� �`ˋA� ������ ��ڛ[�ʑ<�ր�5�/��:���$�-��`o����Ϊ��a���d�Μ�	���JaaP4��Xz�1���<299�^9���F�?!���ń��mzLT��@{c��&����*����X5���!aۨ5,EՎtfl�W0d��c-ɔ��g>=�m��k����%�,��.\�:��:$�;>#L&D�R.�}���1�����1I����H\+���}�/����gY����c�\
&�/�	��W��JG�B6��"��Qa��ZM�^����F���x$4�h��	;�go&�Â��mk���9Ϩ���9���j�f��% Xb̲��e2���e���-�0��?��^{xn�*���}�"P';l#�[����^q���{	�hrg]e�%|.f��ɐ��!6��1�;\tg�mv�Z�?	���F۬�}$�[v��D���红���mZ&�
�p��-�v�b_�s����+��<�}Le&�k�Z����Ʌ^�����{�� pw�N��/�s:���ކ�LMS/�F0�������+_pr o�4�ڇ���ߧ�z�`'�~�#��￤_~�9���o�͢��>��ܝ��iO-L�7~=�HZb�8��{"Vq`=piٳ\2��n�:2<0	@tNlm�'�fy�Ĭ���d&p��ޫ�J�0��(���9��6����������A���� $�����4��Zag���d�(�B���5���"0 )�� �Ɛt8O���mXg��쿾�l�ݬJY�5{�7�?Y�]=l����������}��:�4��T���Ac������ἧFAc��N��u-�p=�A�@�?��
�M�?�fL�y�L�6��O�T}���J�^�Ά$��%kq�]�:�S�/_���`�^�Z.x�t%��j	��b�̚B�Z ]le��]��s�mݢe�u3al�SAs�sVIn�{^ �X���y���Y_�L^�9�1�t�xs���OP�^SZ��t��Ag�=���|yI���˻T^皸^�>Qd%��@F����
&{����4�����	̺jx^�\h�M9�Xxi,��w�􍒐��� 0����Uq����o��;wt�p���i��DUcF��٦����|J�|��D�����z2��kB����c��lH���C�:�4�Ҹ�Nh��o;3�����o�Ƞ@`�����s���������w?�ۋ��X��O`-��BE��E�I't�%��x�)t�2H����f[�"�R�Q:+�>�U�[M1Q�1��H�t���̾��0�ZM��L)�:1��a � �	A�̽��1�,oT�{�*��(K�I��2 ��m��9�x�Lb�r�ճD�J݉<�6��Ǩd� *�HJpF�/u?��s?LԘ�~��J߿����T����nȞ�lˆ�	 ���L��aO�;\�Y���mw]�t�]�˾���*����S������:�%ж��{�>A+p2#�:˪�J+hV�sQ���G5,6�p�ܤ�,����Aṓ_>�&&��&��i�L�`�}4+���z��k�	�Im$xV�6�����bJ�Y��.R�(XZ���.��/��U�<۶��:�Nn�x��T��3֛�!���ŵ-�����n�q$��-Mj�D4������˚<���}+�b;�g�Ҟ�5	2�SA���7t�'��]�
1�#���`S>kN����D1��h�����э��`��s��T��bՖ�N.`6J7�E���[pan8�`׆����m��!�@,�v|�;��?s����b��
�`� �����k8���Q}��s�hϿ�Y1&����v�&L_���2���D�V��
��������y���%}��j�Qf���b �����f$�2���O?�����<k�I�������7f���u�u@�Q1�� _v2�|����Vp�{�|{{��g��X��2EK�.�}ݒ����T��C�=���a����i�``:L޿O���1Uz���&|}�Iۻ��C=��������Yŷ��u`�)Z��ӳb��X����JLT��h`������?������.���3���أXS�X7�8g��ߥ������O[�ڛ�Z��bH�5���~��_����5k��N�ؑՅ?��FT���GkwQ�����I��N�#�b%*z��s+�����(B�|Dg��Mb�ҶɌ�����(�O����7�pz�dd�b�!^ F5��y.dQK
9!~���Of�E|������w�
T�1x�b��dHFK:LZ>���qw}����o�_�|!��������	��(
m%������C}�|�����f!sYO�,�����`2s}�����j�6c�ݱw��d�8����yh71��VAi��<�1~�s^�;��N���ٹ,Ty�9�S=s�.��,aݨ�7����n���Ù	ʢ�6�_��a�H����4�h��c�8Th34���3�u��7�y?��ߥ������篏����������×��^y�P���v޷AQ`��Ȓ�/y]ľ̯��������=�J��_���B+/�^������K�I��(�?��t��C���y� �귝Ϟ�*��H]���5
n�>����8�����b:��.�D]u��邳&W]Zɒ1f} ;�*�8�u���Z	�Z�x	݊��ɇ�4������Q�25Z��I}�#
g
})p�Z 	��O�]*��&�:K%0����J��NY����U&���t�o��W����@���� ��%-#�ףl��h)��T�~	:bi@�܂���>�I_ڦO0֪��@<s09r�B�*�=ք���Cz��Ҿ��ՙB^��SD��Â�TX\?���_۰4x���i�Q�1�b�J�*X�^�x�i	�C���[��S�.E��)�4H��N�w��3A��_��P��)�ѝ 8\mX���<e��c���N>���t��H55x�.�'{���r���xz=ӹ ��{C����3`S����A��d�)(Hx���'ڱ�=d;K	 *c_��tz>�׻W~6��罔��[BJ��|L�sM�$:�$M�=��{��T���%�b�7��Q��׺F�HX��z��>
��Ѐ�V���s:�`�GqS�ۚ�'$��)?դ��$@<Sa��`��I �"�P�M~�~"m{d���c(�b1�h���)�4��Ao��Z�$�%#�1��>�Y��	P#����S0$JL��-ΛRswvv��
>M��O�|�5���A�1��$@I�x�8���(7QҬ1��|���&ι4H�s�d�J�NC���VF�\��z}>� ���)=ݿ��y�s��o=�\��[� h�y�L�:�\0<���۬��)��㢻HU�yR�k���://��`�M5(�o:j=�>� 6  G�~�Q��X��LG����V�dc���AUU�3a?�`o�]��|�_��zH�#Y�0��p�V�&k3�<��0�R���MnI���� ����@��P��A�q���H�c:�(M$ �e�Q�n	lV���OM`�"a��Cg�dQ�M�5�1!����A竘����O�����[�[�W�N� gVY12�r�A���(��a�DN��S����,�:���ٻ�ڻ���^��y��6[ �i��7)�9N�Mr���QI=���f3� ��P~����N��W��Ek��E�0�b�[3���`@��uS����]v�$b]7h�i`���1��8tq Z�G�������=�Oƞ`T�$����Hr�%�}& �X}���=���\�������B�k����w%,��0�,?���~��W
�S:%���"��X8��{��Aۚ�raw���Hb
H;[�M ;*`����9G��"9T��5/`�n�5�	��#q �������^���@����cʇ���>�E��o��.�J0f���{%�u�q�U]���t]�����V�n� a�;�_�Kr�p],2���g�c��\^��g�ڟ�[���u�>H�����S��&hP�
���z�3�������{��l�ʃ�W(�|����}�_?�������ׯ����|w}�r��DĴ��}כ-�/��6W�Qx�o`��5��'9��쩓l��v � 0�P�FO�t|6�_$3��Y�!��4�Ŋ��51��~��T�����ųQ�otk�]���-wM�E��i�%�wB*l�s �:k�E<D��%�;ǜn�z����N@]"��Sz�������Y�-=ms�Z����]����}=�_������V�_[�� �ysq�,���2�8�=��[|f;�G�l�o��0kX��,���3R��Hߠ�i>iD;��ӨhI$�+	����������"S�N��b֋���̘o��I�W�_^�=I����=��(f�9I��O�8E���Y�������_����s����_�>�[�>�̓X��2��b҉L����=�ߐr�▗;��@���u����k���];��NK������s�LJ���!��^�~��Cb�F-��L���bǳ_i�/�����������7���!5}�X%��v�Ľ��- A71f� ���Y�A���ܦ\��^�p�G�S1x0IE�x-`���ab��hH �ÈD{֟|����s6�*���#��@DȮ�,`I5)��i�3>12����!�M��$���$��+������g5�������N�јj��X1]��J��k�[��k��4�)ħg	ƆpǠ���� � ��̔7����6���+�������7���hU� �"�Qޡׂ�H������dE��[���Z5�bOX��������F����5��&�ʣ���/�������n٫k��i�<�.�ջ_#�{��
%��ֿ�e�v��ðs7�{�Wo]� ��Lt�W���m��k$��{�H�lK O�6�6b���Sb�ዦP�mb�bRI�N���G
���񏖃.�_ߤ/�>1�c��C��&.��|J�?vu�"�^ӗ�>30{zy�A���`� pLG@E����]8����c�5��u�B��}z���`u��s����@��5�sΣ��5�,��[�-�eJ�R���3p<[�4�#~ς�J&�n� �b�p��;1G�k�6!
M�y_O�-0�+z��NP�x\�r��V r�(�I��k����#D���y}�Ԃ)�g��wyY�~җ�gP�}��^����O|�5��<�Ȫ:Ч���s�x�P�~$@  z���?|J�U_�t�tzw��3�G�ά�}���U��v��ާ�ᑠ�}�[hY=>�4e��+(��������+YH�~p������w�s��BM��@��|�j0)�=A8���n��#���0�P/ۚ�\<�<�}S ���E��si� \�:������dI�$R� �J����W6P���U�Ɍ��:�����yy�j۪ء���&a��{�bZ�xЧ���J�N�2�G�����1��l7��4���I����m1s$�j�B{��������¶�vN��������)��ט0t<�=@=Z���[�c����X;�0�:�ѵ=[�:&ol5�u��P�l�3ȗv��pv1g$ �2YD�˹�Ѻ@\��@k�p�O�:��sJv�mbM��`mjo18-≯,Y�x�@Ƙz ��O{�`|A�	���������������l
�Lp�Ж��~���zKѪ�4}�����x�nI�!`�
y�$``=�݂B�'&�(꠰��?����t���ʢ� ��_��v�5K�$��l�E���$�v��ˑ	1��gO`�z�{��� �=`Dҍ�E�����Xj|X�˶����u}�p��^�+'�.�*x������T�U}~î�ի�A�����=_P���,�V��ԉ+��5=�ߧ/|6�f�{' suI�v	'�a�������紿��i���W�~�����/O��[I٩Sa!qZ���^7�-d��[~�z,�q?Џc�v��c���ٮu�ޞ����R�ԳHV�z|\�1/���6�}Xn�Z�v�4ZOel{Lm8ː�`j�[B�����y�pk���A����H�ŰF�u9�4e
��{�:���I�|�Zs+�!fH;���Q���?ʹ1l�/�Bܗ��*�r���=/$�e㳇�^��Z�$p��B��Cc}QxAK)��}Hq�YhR�]�W� &0Y/#����\��YX�d���^z	�r=p�`;C�`*b�b?��5� �?E��ߔ� @�Y/i �ڬI�d�
,�?����3�@8j���:�O<�>Gk0Z��,0���?>����O�����\\��G����&�[���8 �u�-N�3]�cBb��#>��'s����_�@8�I�Qt6 ������c����؊�����r�e:Z�o���aV�JoiI�khU�YR}Z�7�J ���{���v2���@���g����(/$�� u�-`³3;31(K��cn�DT�j�����J�k����A���(�����63��F�qn�M��k~�aȖ�P'��JhV[��o!��,��&�u��沢m���+j��!ɺ�,NX�P��.�2���YDq�=z䧂$����y1Y�|V�D_x�!FzK�m:f\g�z�r�ъ�}���(Z�-���-Gf�ԃ�DVO��+�)/�jݶ�Ғ̉	�4��M�K��e�'UKc�ic��PN�Ͼ��`�?�]rp�=������q�P�Î�E��t�Xk�����~�=R/@j�
j�4�\�9������	Q6OA!�jͩޣ#9=I�Vӈ�8��1�t�_�m�m��C�o����H}׀��B;�}�y/'��s����j0�𔞯�C]#P������=�� n�]�	��{&άNccY�Σ=���/�2�!"a@"��r����R�a�@
kO�&� l90b�΢ꮌM�����bo����Uq���f��#K+�Y�
V�m�8�},���\��~��5�n��S�c#�KB9�b��@��\o`��>O}��Zz��#L��
i����؃%GO�P%�^Y�O_i��,Q�=���C��[̗aO���t��ӄ���'F��q��}�h�X{���{�8�O<�3'yy]Ou/ ��7� �u�J=�����aL�_$x����g �I6+6�О)n�lm�(�_ŬA�:[ �?�$n���jB�;�5�ȡ}ä	��m�hrD�	f��E`tӧ��	}r�$�7��?��%0k�19Ymm5s/�� Q�z�9^��kc�D�'�'����R"�j^o�`^�+������+�`I~������ϖ���a0"��sW�o��.ڇ�.��uj�Y�|��-�����%h��b �^��p4;�e�Zv<s�A��X7�/���e�Ӱ���4�;��	�`g�v���l��(���8o�/��/���ت�(�i8�����}�W8C'�6m
�
�cri�h�>�7'~^|���v>=s�6�������0![#���	$��*�1 �cք�m� �@`(�5������Ȅ�Е���f��}O��Z���q�T�n���9��rV��@B�8)���
�g";���(�bL�
�PF��_t����}��ǽ�
̃�c&3*YFA햲��9�D�T����的�o���>Lտ��r/�,f$����I���j7,~�Ng�5(��D§�� �PDPG����/���O����,���+�;l0D�� ��
��]�����IBڿ��Gv.��O���?~�����Em\���yD���	@��X�)���c�׵��D�D��j���dC���H�I����qf�̄�. �|��� �W�E��n���J+Z�[nu�{��O�X�8f�C�v2��ϧ�1� ��r�3
N�8"b;9�/�&��;�5:r�TK�� &���0P�}p�߼���St��pO�#���uo\<ѧ�aL�K�t�S��{�>�٨~��Z���v�b��9����2����Ƥ�$�E#}��tO-�h�4�B|<� � ��S�:a���u#��|<� ��^�i��\"��Ǿ=�z���j8z��&b��	T�� �[�j� /��˱�m���Y�h ��;۫���|>��_��s���w���8��-�z�����D��W20[�?�|l���V�rY��#�Z�����*�`d�,���+ks8�=e��6�.7��_�������=��q�DJ7W#۝�=9�A=Q��]M����bL��Ul�g_C(�*T�vSʱ81O��x鮭�4����"�G���(6�4����v/c���?uvZL��K��(��DP�u"!x��T����אIr@��qP����5e�}��D���U얶��^���D��E�̡Ǝ* ��e��Y��u�.��]'`m���_��{�I�`$pݺ�TO��=���₹� �h�+�H5��inAb��u�t��r���>4��AH�{�� a��	$�w�u�\��V�ՊyA��Ab�p�(�8J����*ǣ�!���ܙ;/T�������IL��`�ꆹ%�l3�D�T�>����nץ�݅ŶK���ڃ��n�:T��U[�c�HV�Ƈ�JM`�C�eB^?�������� ��|J�����Ve�iYE�����,Ɗ��1B4�DE�{H�!�/���j�(*5�TuI���ͅh�1�78+<;Tj�m/�s��I"�m=B��PI����g�!ORQ�]�z��y��^*a��,��$�w�&���U�⤹'5X�h�=�<��IgŎJ����pn�@5i4of�xlvL��J�Y5�'u�C�����>D��\3'!��M�ݶ��pY��5ɪ�/IwNW�ّ�l������ �t½S0Q��=߃�PT��ځD����M�#Ir$AU5s2�̪ݙ�������ꞝ�#3#2H��������x�3�$�t�C@ c$���<�^_<eX�uX�L퐗������pИ7 K�Q����铦�w�z=��jY���V~}��0`^<W�����\� �i��/���Z6����Ҵ])9�V���/P��|X�K�d�J�,6X5~(��kZ�rȋ�Q��v���֍�Zϊq�vXo2�}�H�j���]s��J\�<�gi?�E�%��2��N���8����K�ue7>�UQ����+9��5W+�O��&:�C�nz���7������:;⴪#U_,y�N~�����A��׻g�Xz?#��Gz�f�2��ܹ�x9����v�l���1��?kq���sN�0XF+�15	8 8��dS����L)7�y�(t��R4ӻZ �2��u쐑k P؄�U�Xǚ���K�����j��8��U'P��������_Y������E�w�m�_��oQ�r�?�?���oǗ�E��.|i
Nuۻ����,�I����,>%�A���Z`>١��_$ �UTA���, �pWhfЫ�������Q~��ˡ;A������}g����M����O��/�_��/��?��`I�`(*_����ͺ�i9�Z��l�
2��$�GQqC�������k�������+,E�`
y����$<9~C��@�̧d�J[	����\�����A�gā�_d�_�������)>}T[R�W����?�l��Z�1-�|ڊZ��K��?��v Ԭ�"|{E9��Q�2��n����?�U��w:u]��SϒC�|E��~���|�/]C�EKc�+�2�}��B�GЎ�g�1�Ͼ�gu�Y�0��1���6�[{3���ݿ���������c�X+oZ~����]�Q�w %㩙��*l�`��_�<�������Zf)Y�,A*tsK�26��_����
�����7P��jz#�ŹOAZ� ��Z��pG����؈�����#����2�H����m�����ކl������Y����Y����l /��5��K�r��q�?7��j�4%�OO�`g/��� �_M�oǿ����v�o�w��o�˱�h��G�/�|�7��7�������tQ�74:|�[�g�O=޵U����Ѳܵ+���v�Ky�`�f�����z����O?�����W���5ᅁ!v���_;�)��D�k���8V�-`9�ݗ�!NUciWj��Uwv7.:�%M�]��cA
q1L)q�v�s�9o�NQ�uA{��F�	�������K��g(|ޢ 2�a�Y@5D`��u&nD�Yu���Ŕ���H���.+>��#Y=ڱ�1\��s֒+��$��4^�����i��N�L@u� �X$��y,ꯠ܎�۶��Bi�BЭ�#ߝW��S �+#�
m����%i!K��83H�-��Jׇϯ վ���N,p8g���z��0q��b��Ȑ�Zf�tQw�X��}!k�zU���L૆�����n`�o���Q)�S�k`	�r��Fa�D�6���+)�8l�����ߩ1X���Z�?}�	N��D�\6��e[vc�at|I���8pq�T��~�è�����p�nc2>���+I:���������$p$����Mmi�I�p;TKQ%���m?�UA�q�(1_5G����JM��t��lk�õ,��Z����Z�$JI��p�xh�;�Z_�t3�j�ÝDE���L�̗՝:*�ͺ�8o㪝�޺E댸�x��x�j�&���j�V�3#o��u�����ן#&���h_I �h�5-3ݬ�����d�����XVJ����8���}��:�it�*�/u��"EW8H!�o���8>L�}�v��_�����-Q/��\��.��/���Ҋ֤T���/�oW�6ȹ4B%�q +�h�'>:*:�4'��k�O� ��	�˥*y���������Ý3�Y��Z�JV�:OX�b�(0�]:�f�h�"�z鐑 ���K& ����$���͡�I@��'n��n�r�q5S)����Tj	G���#�2�]�Z��٭{��1����?��1��Ba�M�猔��r�g[�#�4@Źa�ɥ���ȏ��{,�H����_���{vv�2��0ے��{�D�=�[���9o��2�HK�eV���a��e����4}_K���yL��h�K��� �d�=�-�������� ���6�|�/��ܾ����ģFh��,I��8&R�+���^q(%h󻔾	��Dp+����ǥ;�?{d��.����P/�8� ��W��^6V�O�}D����ݲu���z��` �g��:\=���9��i�vd�M3|��	[뚙l;�BF��-^_YT_�o��&V޷�Z�˺�ǿ���;�3�t��	~��Q�uѬс�co�!�2��5'��U@h�ND���ק�p�o���+��Y�U��F܏ݼ���Z��0%xG@�ۆ�kY@";��Cd��(��*��2F�>e��M���Rcp�gw���'���m�}����C��D�Y�ʪ���!)�[4��UJ�>X���y6������4J:[�W�T����Mcj����M������s��Ro��sO@��$g ۃ��t����o�3�H%@��ߊ�L�2�(���>�c�J	ZC_ky���q�|ҍ�ve���cl�߻Wf��M�x�� i��C/hw��|� 6i?Q��g6��x�n�Ț�1�F"ن�}��W �{�6�2�����ڵ����rJ*�+7��l��U<�l����_Ͽ��3|<^�䙬��LJ��J�׷C��$���b�r����TH��l�}��@}{Hg0CY�d�����'`��`���xCs�1|�Zb��U".��X�X��5�qA0������0�*z�S�8	d)����<#��	�N�R �qu��-�,t��1�Js��@$��B�/& ��K�0��#����QT.4�LDԫ;�\��1c/��}�HgZ��:�l���l�+�ʹ�)�2�e�K\-�X�u�<�u��|�Q�؄��~�Bm��n�B�)y�B-��1��)n����&y�o�s�X�=���o}����o�l�5��)aj `�S3\��`օ��0d]�@�	yQ6F�v��#��53	݉�©!���V�`� �2-p08�����ڱ.�(Xܰ�L����u} !��"%U �m��P�M-�+�
�Bz�цm��c�4����cKj��%0�4Rkş��]/d�h���I��yʽ�͝/����Ĝ�`�I�5r�4���S��@+fUh�^5r_��͹O����K
�4�n��O������0ڕ���bk��o�Ų���A_�V��;5$��/�/����rD`ȱ�
C����(S�."2(����ϝ}/�Ì<��7��g�B/�o��o/Vˎ�*� ���7o���OΦ=���}AG�m����50�ice�A	���X\�C���
�M�~{3�޽;���rwwP�-n���<�:
}x�����j�A���,S��n};:q�@�_��|Ǘ�h��~ԹT'��:�_�/���IkeĞ!���A��6�L�,�
n�� {2[3�t��_�����<t�T [��* �uqGQ�=9�e H:.�*9g�ڞK}Zv7�#���sp�l"�Wf4k��j��V���4a�[ �cn�-6��`��d�a��`{U8�ù�*Ʈ�S뼎�D�:s� "�LE��C0�Z��DG���K22����3�����5{T:$jS��ZҝJ��H�w�\�zg6fߩ'wspYⳘIɀ]�ݻ�`t�ݭ�$��d)հ���n��\���W-(�/)���^	;z�. F� 022^YC�eQΘ�\r���>���'�����a��{4 �ڣĘʷ�b6˖���#��~ѕ�y���c��\�Y�`�π�@�a�V�ܿ��$�
ξY���{�p���gۻ�J��30��꙲"K.t��Rj�&;�wZ�xxa78��w#�=�����\�z��?�w7а���}��"��۪>���F�F$�hZ��< T��'�~��I	��Н�����Q�R��?�-CIJU�*��2_���%�qA��f)�W*���|E�Id�3���5�v���<�+ió� �7���e�b?�$z?�������&�d(�Am�Z7-�ы�;vY�[��/,is	�h^�1;7�]	|Jy�7��d���?jG(�RB�M �ޒ~ߐ)�|S�G����'(�(�͎������w�7)R|�P�VM���ic����yh'm�s�].-e2�,5}+k�&���w�O�R���nh A���)�ʠ��@�����&l���;H��Ŧ�VZ5��h7��b����!o��H!����ϗq#�]'�A��@�|0(:�.ܓ�swX!���(B��e��c�@�׽:�'��0"0a�TF�O�n��1閙�^�\���<Q�y&BK�1+ƴ�1��p	��\�g�������0�K�4��Rbi�##\`��y4 _��k�����c�S�Jɇ�Ơ���RtR�������-IsD�NR*h*�1Kn��~W�q{��r���?�[��oϺ�pg�w]�vz�"��Ȗ$ڔ�\�2�:�mN֘�o�^Ed8��!�,!��2�lџU����:���f�L������ݻu�y��9�TxXh�#u�����Q�pc�.$ �h2)}�v�t�7��1}�ֶ�)ŵp伃�}ޞ��jP���F�az�=�i���SR�8��Y��Ş�F'�Z�x#R:�Tt���i�:f�E:��b����*+D���ޗM���tE�u5�uR�����y�2 [Ԏ3�� vd.��~��*Ț���?���x�+�;��	Q�:`�k"��Z�^+��.�JD��ī�,�օ����|�����������#�����NI�k�h4�WZ��l�ɬ�ܻ!^a�I����ޯ��;C^��Z��[�P��n�,���|-��L@������ﴡ1FP
yMN׎4s/%��j�
�������@I)F�"rpJ�T�B��B`8���V�ؽ��Y�Z
�%pO��<[�2�FK޴y�ejj{��aL����ڥ��>�]fVDy�g(0�~���C��~�<��3�Ϭ�s�� ��3���� �U�X�����۰�X@[�@��c�{Wݭ��~D�~\GÀ���{�s��
#h|1xo�je�t�X�4A��Ќ!W�E25/�ڝ�e�N�ґK2ᮟ��U�,���?�vȆ[��~T���Od�i�re�D5>�3%zg�	�)�Ct$t�0X@���7 �T��h�(M��
��*�ѱ�[&S���8�gޤk��g �7~��ef��YT���侀:��p`*�c��z9>���u]K9x�(��cG�(�N��>�i;19ǭ]u�n���+e⶛O� �~|��ݽ��)����Z��X����!�
]��1_�q'dV�!�RK��	گ;�t�� ��V�����=%��Z�nb��-t e0����U,',ty�š_[����Ց����@�Z��)���t��p"	8а.u���e_Ϻ�����W����R�������3�~  �vY��� 2J��2�F�۔��ܞ����ʉ���C�3����
�!����[�������"�}{��:~C����Tb3�7 �� ���t�]3�c<��;��v� �Ң^6���l��Ӹ�6/�3� �ĘuZ�Q��)��˵\W��,sfN�%>�~�W�˭Ilf��W�X�4��y��ً�-�x<��v�;*n�?%��M�ce[7{83�u��0n�D�B2����H�M�Fy:&�I��ɤK����u���1�H����hwD�R�S<�d�e��|�iH�t�
U��L�l�W#.�M1�;ht�)�j��_HP`�3����a�	���TI���!��I�_��j6��*����["I;�Q���h>��1�)`�Q�T�F6X}�U#��\U{�K�����aA�?������LO@�/%��M�z�1t����_��f����
RV��� ��gT��K��y��b�ST-��6�&��k-j�s(��F�����E2'YpQ��@	��}��i��C�u.F���7%h�bה�>|,t?5��/ ��R�2%.��p�����8D\/|���P�Y� 5h�-�}X�OH�MZ�Y��#mǼVʽ�h�|*�`�!��	��֍��7lg�o����J��@�])����S�Z&��k�K!����*OAO�I�;?|�r�7!曋�v��噮�n�/����<Փ���6� �%?#��� =��wY>h9,ú0,����h��e�2��X_\�*�e�(��p�,�;���@��suXKa��^�Q��e)�X/F K��4v�]�kl�_�pv�+�dJ���ܳXdٳ��ֽ�ԍ�Jcex� ��a��c	�I����KBT=v8�����Ή�^����FXw�+�3�#uK���ED5�Գ3瓀[�]�������� :�+����������O!t�����v��w%�&w�Cd��r�YJ�%λ�*����AFm 䢧���\���$P��Xo�c�a(���%=��(��W3e� �l�u�\Щ�A����vC��\C��/[���g��eK@o�� �mNeO�\�=c�;�I������#����u}��k�:fcGݬ1�f"��J�Q��;��ռ���:��m+U�}v\O�:d�dfl���!]�~�� ����C%e�j�/k�K*�ִKJ-��İ��̉9����8�	+2�Qr�|mR�'p��^������+4����qm����TGz��RФ6�����Bf�ud����)��:���f�%�Z@��ʱ�o��� ����f�����@�:�kd�2ք�����ޮ����a>�#�0�Z3/�ŁV��x-K����2`��;���Y����^��Y�k�VZ���i��f��r�I�;�jn��W��#ň��X��t~����5`��׬rbP���E	�q^MW�t��R����h��voj�r��
@3J����C^�:����{��q/ݵBap�JV)�b�c��we,{�#�k����A��ј�z6�cg�*����m�ow m4�u�����F��!@Wa�
�ix��0W��1�O~j�أו�&�yMm�D���C���ORv��QKӝ��ۏ6)���_дi�e�-�uj�pJ�q�=�^b]��5��Y��e	�H �Tfa�ng�$t8�;Tjt�A�����h��Cm|�������	
���/E�� �����m#��E�;ُu%;�4&�мCy��<�C-v��X ���TdpLY�jbxd^D~ֶjCy4��Zk�&�|�rr��q�-=9,E��Q8��5��R�q��z�q�ǚM��.�}��'��^E�w �M�ڹ����aem�B�L7���Fa�OS��9��J���µZ�όt:����;���������3:�G��Hur���YV�9:Lpm�w_�K�ԭ3�I�l)��G�vDXe�V�O�@�ݪ3 ��9�ivH�.�}d��qTC����1�o��ҠG=��L1,�i�D�mLY��D��#���$K��	����q��Sc�^}hu�2";HQ�z��#E燎�([:��8����b����:8�2�u�)����KP�'����Sɭ��T���בb�����a�l>���Y(��-�m%��Gfci��[!?�q���{)a�����;͛g�шH��2O5��TC�HH�*_�Bm�-d��w�a�E��0]�V3VYb�ĊR.#�,>>�F��5܈3�Y&<˶G�rłl/7���ԝ�6�־�d|X��RDJ����Tj�Z��f�[��n��V'n���T�JXܸΑX����3@ d{AV�Ӟ����3�vtGT�V��a@�������{Ɂ�YGР���	$!�y-f�l�ݝ#u̥���do����fK��  ��IDATB�h7�3�#�&{D�F�Row��` �Z	L�ܛ�H1(�3Y��cM�$�4�@�p@'�ߘ)A��<�p����lB������T�;8l��r�ws�\����GСY` (U�IV�e��/�G&�$�|�p| xP@~YpmGǯW������|@x����oI�`�-�q�O#�v�C��"薮)�����v'C4ku7�w�Q���[�)ϒ�P�ګu�Q���W�/!nU��D��y�j�# �1�V���#�*d� �4=�F3	ԊE��%�/��	�1�$)7/c6�^�� �Q��v�������~���-�L�ˢ���Fxy4���e���fp�Xhk,=2�E�.ЭN-�ҙnN4��vf�n�/��
�H��p��;_۶ȸ-���3�ٛ�"r;KE �����Lp<�m�v���	%r��&`��[{�k�c�wr�h,�xq�L9j(��FIgf=^!�
�s�� cr�����s�1e��+��7���@Vy�UA����~����:KRl�^%]�5�É�v��Z��_ ԑ�
��]�͸���Z�V�'h#�E��z�ѡc�su7�s���\c�ٺ�<_��U�]-�9������?K�5��'��Лt�R�gw�	9�)��!���vb"M�s�m�2�Ӯ l͒/���9�g�����gu���I7�f^�t����4@3�Uؑ�Tw�����:l�]!���4.�=��JA��d!�M7�v�H9���X�D���^����2?-����;�}���J��p�7�Ԯ
d�̓7N?����<�ϵ̫"1���"��Z�������<�qW�^����T�&'��0�nx�)�D6�$jC�B�t��9QO��ѓ��szG�pL9 ��TO�K(p������U��>X���q�4��P��3��V�7%�Q#U�G�R����[��ųb4ʧ�4M���2x������s^Ǖ6{z����4��>|7���`��{�2r���>JqG+ύFr���܄՘>�)���E�<nހ��'�$k ;.`Kt#���9ݏ�Q��_���͓/�HE�A9͇ޝ��V�Q�э�{�"�v��{l�(r��ef|7�� @w�����4#��@A#�It�Y/T�;J�tKY�ϖe>��٭$��v�r�7e;�>ұQ)9P<6��.8���K+U,�%n����3�b�h$J6�f8H���L��s�)�*��҃���o�f�6YnT#��Q+�{,�*ƃ�<���U�$ﱗ����Ʀ��Z �:�Ȓ�������j}��R4u���b��͆J�ʣ�L�X�C�����Q7 
�ę�F!�r��u����H�'�6�M�,���R�E'f�r�dy|o*�x)@�4����u��T���ݞ��'�֛��"��@.��5��л�lw8��"��v>B��[�����g�u���XJu���1,F�mE��fv3���t@���O�����O�,��Ѳ��V>�:�4[��x���b�J"���Ֆ�m� #��x�v_{�E��$5Un�l�L�zih������7#'��4sK���n��<Kdm
ƘU�y��KNC��(�T.́�������������,�ʺI슬-��L���2af�>���1�>��p%8�
d�SM�����f9�e�B���,�2w�+�C�XX^�q�sL�0uw�ְ�����<L\źpn�Tn;��Ze0C����p���<��� kW�ܫ��$����(˴���8μWx�	�t�����E��aݺ�O�]_�=���I�Y*�Y� ڰ,�\I����`�h%:B���Y���G���Y�B�L�A~͒�l:Vi��Xnс��%2�.�[p���g��Wm. ����]�tl���YW������&#P�=��̻X��O~o��Q=�sVՃ�����F�|�^�)�k���U��aYG�!���������/�����Q��nVf#a��E��YH�7�n×x�Q@ �.3JaW�i�&[���02��,�+e�oRmyF,��7�G���#6�ty}�|+/��T��CG倗�����V58�i���O�0�:В2.v%�8>+��������C�јᩳ���J�<L���[*�,T7�������
uQ��K<O~����>t>��]|���%�EQ�,@���~��5D�ꈛ",PKat�#	!���;�iTsX��>��Tt���T�҈c� ��`O�R��{`g��.;��g<�Y����+̕�V���Ш�J��.kS�f�d)�`���O�֤Ek^a.ʧ܊�ȹ�Rb���K�:�rv�����3���>�Ʀ=ˢ ֻ�V���eT�2�-b��HąP�)BhNh8u*k{�1���L����%���$phҫ�5�P�,:�x���S��<;֑ӛs��=��d�a�m`&.]#�سBԢ�6�6Ԑ)�#�X|��N������/FDT�"�W;9�!�(�ϢY>¯#d9�o�áh/�W�f�.�Q�gL���a#&�
�]�#F�y��:�3�h0/�����γ:��c�E�� ����;?C
�#�S�;���`K��R�Ϙ��b�xy��	�l@�\P: �������-�_x�aC���w�}����X�V�����h26�Z��ع�#" R�~ɥ��W^}y�p�L"�3�o�ǜ�/�3���főc�k�Q�`���|�9� Z�(��ÀO�!8��s@{Ϝ�5�l.��
u@��r���c�����tZ�����z��<F��0��l��>||Ja���ϫ;��޵�9c瓖.~��Is��3�V�hC����� �񔋂��4��vFI2���St��9��[��p�q�DPHxb��9f�"�F�QU�c�`p-�C�����T+�뵆��u��/2�ɕQ��﹘�u9�BZ|��r�}[��"�������s}�Ļc�:�A�v��6��Lή#ɺv없t�᤾lβJ������ι��:��8JA�&PQ�-כ�Q��A�o27���;Q�U�f-��߃�ܞ��M��2���`70�#��-����cThP^��p��3�甄�{|)XA�cD)�@�jdvjJzqRk��'D]��>�r1�EK}�U�F `��YS.��3��a����Z�~7-e����d�ت��ߒ��rs`g$yҐ�sYsV������u=�Wd�� ��k	Γbo ��(Q����;���e��$O�P��p;4ٯ�I�p;K�Z�֏4�I�e�$����a:��i5J�^������틎Cg���<zz${���w����G٤�~�Q�}b�\�ё�<�YVp����U���o�u�W���1zt��W��v��Ǜ�^4 ^貸�B����u�j�g#4[Ʀu���Bhw�W��U���Wo%��r,��v�u(���@V�P{:㭸!�":�(hC���ĉ�k�V��g���' �y�+���և����N@v��*p��y��,��{�F��Ш����L�E]_�Pl�>���3�$̲)� ݳ���	��Tr$�y,+�I�����~g �wf�w��F$�i�����vkYY�L%jeT	^R�����ޔ��R�t����6|���_�sd�&{6^}�k�#~��i����]�%^_��um�r�:9�G����a�0B�a���NŸ@����H&*�G� �8�悳g�ˇA���9��c�d=`�^���:߭|���x�	�y�5��b-_.����,ƒ:Q`��).��\,<]��>�4��t�X��*g)-��|����+�sn����߾����)(uq�~��'��ʗ�k�,{A���KM����s M�OTC�������o�L��{j��������HF@e)��묗�h���%�Dg����@�Xs�q/�B`�\U�V���2���<5Q\�2T����|�2Ǹ-L��X�`��ˮ�l��/>6hh�r�L��na�O������X[kNT.)�h�JpPRd�����O� uf�ls��t`��a�@��i����6ȶs��;��!��#�93)6����;e�;�����0�E	a;>�+�Wd� ���R�g%>l��&̈ag��u�.�y������؏����jiu��"c���\�TF��`U�5}2��r���c%��ܚ�����TW���O
�p͙#c]�v8�W���#��ʭ�4;�2\^߮�MKN���Jvݒ�,N�4�,��\V�H�oeN����sd^�#��-��邲V����L"��`P�\Z?}��	�$�OO;�Pp�@��� ����R�EA��\�dKp�K_�e�9Bs0こv��D���ki>��Ǿ�Q������d��"���Z����]$H]m��2�o<|?J`�/�^߳�.E�д����_U����l�~�ߐ{��TҴѲ-��L��e��HN6�"Bά� ?s��QG�>���� �Qֱ�r�'������ܧ	�h��v��Z�V��\��C��V�$�n��q���-�c�5�g��ߜq�!ëO�{�n�����#ѓ��!%M�>~Ա��4`�[��Pg]x���A�.�k�����6�P����-G9�q /V��8!�������ܨM9�qC��.lx`�T7d����S�s*'N7m�%��k�M*ӽwɦ�|v?��y?�ښ��m��I��I0E�k�_�yx���a�
��o_~+��#�� !�L���nC߇eC��H��N��{��y/��Yok�f�����ZF,|B/������YW+s�� ����e�&j��&�m�W�.��q�-^r,�XYw��_Y֣��t)S�U�8�CcR+�1J5�)�I6v�KH�nf��1�h�	r�.����_�3��:C�A���.��|���xq��rZ�����A<'�G�L�����|�ѹ�;m�t�����}�.*�0x�r�pf�y�ts =@\���Ϛ��J"� 5�~je.�R�/��~|��S5�Oi�5�xF�p\��CZ�	�,F�4������!!qM��x >���i׫~N��B6������7{�>�9�؛��
�'��G	I��p��	��n7/����%st��h�<��XJd��V��>` H)#��ĵp��$�����
g��"9$\K��{Z��^��Kߌ������_���1ui�|�� �I�<������g[`�(�'�'��!<��[���G�e�0����gakT�ᮐ��?�����Or���_��A��)���ު���=u*(��dJ�@��/JHn@DEɣ�~�(v`�v�_�#�G�J̗g��{yS  ��㡑@d��u��5���}���wfqt�c D��o��ʲ��������Ny��9�d��.x.��d���Ȏ�!�\W%��0�#�
��Ğ=�0��h�KvNX�6���"KQ����-��:��Kr���p���Pȱz�����_�_,��dtn�(ՉM�u%��R��%)�gsڼ��K�̫4yҺ��mZ���`@��ƃ-��"�C��s���v�A�Lyհ�w7\�z�z&FD�c��yx�P�],����a��$KV��Q�4\��e�b�۫� 7fm�Wp����<7};:����J㋷�e{��bݐ$��	D�����ZF�<-��_��W�� ���V���]�ȑC��n�D�t\ع  �uFߘᾬ^�EN`���܁|��~8�2�7��i�=do8���7�n�T�52g��Nf��]P>\ ��yN� �/�je����O�Ѕ��lcq}t=��r�t^M�E�$������w�*>�:�}p�$����4�5�Mb%4#4g@z]mmMWӂ}ΌB)+��I���-^�gvy��|Vv@�w[��7d��n�g�-��Z�C��}d���AH��\�O��\>��j�/8���V|��`���1�E�xvn �������-�>�xw�^��p`��N�4}(AA_V&4B>V8���l��o��6 �Ú�h���m2p���3hEPX�C@�:]�1u�|����	�!k�Y-��J������{�؁>���;Rgə��ܑ{�9�}(�����k������u}E�u�sy�A���^��@��<�a�O�3�K���ޓN��7 b��(j&Z�WY(�h�V����M�)� ǱoC��j�������4���ϴ]�i�妓�KvqP  :���)2;���U��+��
���u�Y�>-��@��B��_�FѧW��x���Ƥǅ}��sL�xk�~d9�Pt�i��s��Ѱ'�� n���)�l�8��,��Y���X���@lњe9e��	5,Aw�J��������L�H��F��)����5���tT9��d_.������J�LBB�J�ϟ˟~�Y���0r�[ޕQ�z2���`���?Ca̛=a�ud|�K|�F����}�w�0�ȍ"Y�����l��Lc1v3����,�X%��p��m��dIk����� X�k�釰g=%ʠ̡B��Y���үw��w{edc����N!��*wt<� j�Z7�nqp%RZA#�c
���m�(	��4[o�y�U�F��k)��=����ǟ����O?�����?}�����n�ܵ��ou�P�Q���U�ݢ,��~�x~v��5��1�z����e����փ��IY�|�8؂4���KdZ�c�O�W#�O7���d�9'6O$n��G��{�R�.Je�C���T�uF�}#��݊����d����H8 Ι&������Æ��_ʹ�,�� ���%Y��5�`�Z�@�$K ��b�k����y�������a��%Fx��i)s�H�ϙk��h���6�C�׈�]5U�����~/!���R� W�_{�(2�9��%X�J�%����*��e��+:Pʏ4�4�)������dxTϓ�ӡ]<�b<u��ʎ0�m���Iѣyq��"�}����x�<����ȸ�Ns�u�Ne`�F�n�� �b<e����R�*�mp�
�Ȳ�T���/������?��r ��e�?}Bv��I҉����b�>�t��#��;�yϪ�>	��\�[l�����~�]��_�^���S4� wօ`TK<j���ٕ�(%�cmk\̱%/�e%��F��,Iܫx���z�^ Ug�:��w�R���L�Y`�E��R�j�]�����Tۖvd�؁21�iꠃօ�~!�]��{��`<֐d�|� ��2��(rO3k�ȉDε�g��z��s�I�wؾ[�w���1��`�a��Q����L54�XX���ͳ������F,ۗ�o��I�m[��Q��}U�kF�b����R��`U(OcFx���]�z\�M RF��ր5��<sT㯔��Vw=�V��< YX����F�[����6�~�{���s<t�)t���,��٩3@A9½0�̅�{oQ���m�j ���x�k�&�/���$]+e-k������?�� �G�u�|�L����NuРL�j���E0���2�屘�B~��z|��7x:(�n�z){t=t�r��}�����|��� ���\��Ö��:k����b.p���B)V2sE��#/�rB�|�ϓL��ﻟ��g2�TJ�wg����hr�ږ���>e�{Ӝ\��@�������Rrau���:���-:�w7Y���0���l0�v=Zc����}"Z2��<j�GÖFml�h�1� bO�ӝ$w:�8�?�L�� �V��l�@b!�sv�wݡ���Ѓ;��Ţt"���'%���1'�)�� ��u?����F����`������hͻ#��5K�z؁!�_����+/��DM�iq"nLnةX�K���w��Jẳ�NE&��!|U8�)�|J��=9JT�Iq�
���<�ז�0��@rM)�xW��˵��n(�qR�u��:p~W8-+�	F	0\�����?)�#�rqn���?%�D;���^5Q9<�d���y�{��_��"�f����ā�N������R�tpY詄�'�x?4���9i��Z���L��w*zqٓA�_��S�_q����ª�>D$� ��$���� vt-�S28n��̔Tn�k�kGD�׸w�ߕ�N��3a�G�+�{1u�I%$k��|7�h�K���B�ջ1c���#�\km�|�T���Q2ڗ����꼑�w5b�G��Ó��Ky]�2�<D�s;�y�"��Q�E���|D��b��:�@.��&3Kޞ9���:�!ڲx�,[���S֑�ٕ̹ڸ�}��N��Ӎob� ľ��.ՙ�,B=��/�̑B���8��,��C�e�n��C�Y/ʨ-�qE��k���!��:stMϐt��2�l�Ş��Ju���	�5"χ���yZ�5��<����)���g�!��sAf���Xƌͷt����N�V4G^�\�o�!!:섧g�g:�����[7  ��g5,� ̆{�w��$nA8�� ^9��XFD����l5�M�m��fdi	��'�!3b��>Ic��֝��I���
w�]g�l�$��k��ޢĳ����r����v+ˇ�?�"13��>�D��v��������5�l��je�UݹNY�z`Qͫ������<�<!��l2U�)�� $�N��>��D��h�p�������i0h��ݷƉX��FZƫ|�=�,35�����_I��D�|9�td��P�A�����۩��w��2Ӹ��&�h�>xm��y�,v��<�c�?t�uۢ���i=��t˶��t�+˦�P|-K�o����:7�g`�|��?:�%�!���G����B��yM2^�)�[��V���?�û�Á�;M(ގ�_[��Qܸc)WS駷ԁ�xF��M@�Y�f�"�1�c�â`�WJ�]=!)>`
�
�s=�X���>�T�lF�8�v��?/���t�{r�����R`0�0-��.=�JE�FR������R�E:�P����-�� ��)tӍ�x�5���'�7��Z�[��$��vى'��5_dZ7h�LϺҮ�B�`� G�D�l��N����3���Q3y�*����.�=��ih(#3`�D��H,��}t�E[=
W"��}-	��!nh��ix�	Wd1�T�~N���97��Y�yn9*��U�9v�yF�j��u8��\,���pY�O�62)���)ћ)��Ԛ�򵟣��nҖ~�2qA�L/�ގ���s\v�,/>0ަz���Q��σ�����6g;��L�԰���b	��;�]o����`4� M���/����wdph�m���pgB�	�=i7&Q�BZ�p4��ϟ?����FvSv5dEʲ�|�ES��Y����EV5)�G����:(0�U��e��������p�`K�M�u��t��,�}��WO���(W�P.×U ?(�Y�~�9_pO��{ c��5�	%� o�)A�0��fhDg���V��J� >���M����<�U��G�%�{ԕ�\����'J���-���1v���?�O��S�5��7��7�5�3�<Y���}�=+X��Ɓ����dKY���\�S�� �8��l�O��tqc�2Md�:� ü���mu�rv��垖}����!�^ǻ�����M�Ew�=f�N��;4�1�1��k���`��vw��q�h����bc�.̬�u��1��߷���A}+�A��õ�Q���|6u�������ó�;���N�:� ��> �N�FݱL�:Bf�ht?���nZbaeӗ���3�����%Y�V^_?��l0fO���� !�;\7gD���sY-M��ЅƂ
v�C��:x
�.c!�B[�(���<�*���A3GTo����;�� L:?�-(�m�D�i�8�f>,��p�"�_�Zp�xɈ�\�S>�z&׍)�B.�.�G0߷�F����8���UŰ�MUN!��r�}ލ�O�������A���.%�%m��dh�!��ߧ�Y�����1d7E�.zN3�$�z[2��ǒ�8��T�Cg]�����.��%fn�wi��D��;hsk>�r�46z@�mP��m?2(*�������L�ݴ�t��<O�u���7����|�����E�|�t����>u�X�հ�\����>8;�ҾV9�2�i�.{ZZ��`�k�*/W�:�Us��3I9�u�]�` MY:Ph ƥ23�8خ�]W�2�㙭��|Y�a'/D��9!�/�z���k���|_�#-lR�>�q�����4<p&�`N�Y����C%%�Y uhN��|��iء�5��ɺ{Y�9�ۓrM����&ƕ��φR9��l��1�{���������������+[;q���H������(Q�v9n��xQj==r����&�o���gi���2;���%I�K-�xU�O|p��4p�����z���狾�'��p��
��t�{���ΐoґ����[��: ��>�4�7B%@DwLkn5F`{O��7�i��ȏ�.%�����R�	9��㳻�ڬ�ֈX��)�&�����S��8F��E���,1���p���VKcp?�1³�3�9ƶи�q�Ǖ���5�t
H�u���7^�9Կ��l�����@�p�8��F�4B���|s:�ר\
���N2y�ǖ^��B��<#LC�����"��/S6�"�ekzS\�-���W|�d��p2]��[��u%�5����ߵ%��;��
��V��Ĳ/�����G�{�F��&��ܙ�Z�2K�>�/��Ǥ`��<�y��ٛt9������攉qb��1����Y
�q��y�hKJ�܃9�}��A����Z�K�$q��֜B���g��>� �u}�U�q�-��A]�뫤�1��pG���d��h��� �(ݓ��~��S^�����rc��p�\��3v�^�N��S����mr*�|��Ϳg1�o���#���n�,�3<B�_��1ʽ��v�5��vCuL�!���� W{�@w��ώ��H ��<=��ޱ��\4]Pk�Jf�� B��ӳ�B�~����бV�h�_�i��H2ypo`�fD��s�20�~�\.�G�����D�����2�}l�b�W�݌�s��Z�U�ׯ_�˷�8��Y�Ì^�H�	�#��8qW�r�,bu�� 9V�<gq]���ɾ����OeX4��FJ��+���'����mnd�#2P��i�u�����3}��`F������(A�n�W�4Jv0���}���y{�ayY�X��������P�a���w<��7�9+#�<ۚkKIvI*�d�B �����j��E��̣�nA&'��$J����u+��c���tP(�嵔R�M����J׊�B-�1�4�2sFd$��dW��l�G�'��?-(�C&� \��$/ 艹&� @��d�!K,w��1q�k��֛ ������u0�����@y�fN���uՃc 4�=�x�ة�[��#B~�G;	�Ҟ��J��怎�A��D����Ջڞ����=*����*c�Hn�������w��2o��4�7#�g����9e��]�f�i��՚�h��j`�eK0�R�݊^�=[$ZD ��S��q(W}����܍��{������02?�K��3�&��cJ*�vl�,
QN�P��а��͈`��h��-7(9t��`�N�?��o���}�[D��V��?�^8�d�E�B�z�k�Bc�{�Y��n��!���{aT��)��&9�lq$29�1������?R
͑� V�A��3�8٘e��#��G�Qh�GF�
E��q��ʬq&�0�>m�l�f�<��T5��eB!ɨ�*j*(�� 0���Q�G,a���I	��A�6��Ry%�o��B��R��/?oF��d�1�X�sFĮoPSL�J8qg����۬�~�ّ ���c�A������>t}Vw��A�� �^��ٵ(�u/���GY�e@亡��R���o������:B4��o-������6F��;ѓ!C�Z��T	�$�����5����x�0�Y�L�ļ�X��0�CLo�c$�5#䢏�5dJ��QƷ�2��{���,�#v^N@`Gu�>=����5P
")�7�� �=>,�$����;���c�g����ߗ��{���b��)��M2����m�^̨,�~9���ΊrW�3����MO��(��}�#����k�C�9�=!n�Y���s�7^y^�#�2��w��錸�|��]���쵗����~���2����<~����{�A,��������	������`��%C�H�/�%J��"@ȗ/_4�k�,;�e��"^�Rl?(  �o�'�y"��s�s�Q���9yG������ϣ��H�':<]��:y�`D����"���Gp���ޝ���x�����U����W��kǡFRi��JT�/_r"��K�X��Y���H�$�iOٳk`o�Ȃ�St(9��!��;�_X���<��r� ����Fζ%�P��^s�9�ޱYl����J�e>o[D�� ;Az�.�D9����(Ϙ�%ٌ������}`(?�hpB�G���hh���̪XP.��_X?��v87Q�K}!m��x)i.�֦r�����X���Xw�c�
;-JV�g�|�X+�#z�E�+e���uo�5�Ƙ��n��I��@W��Q:�c��d��cU�m_�'E)�tn�V�@W>F��:�y+;ng��e-C�M�ͦJ̮ٶ����?����w1��~�k �5ԕ��(i�u7���H	 �{�?Z�?�-���y���$ v�Z܎��ݮIA9�����&v����s�R�؝xľ��͞��C>`��8G�T�ȱ�`�e-���h�C���S�,
/�}m�ýIZ��4�E�^U\�,�w=_��a�=-u$�>��Qh�W߀��,�$�������:����Q�Ϝ�r>�3�s�o�����NB�W��"���r+Y��1�H�oLS���:Ot��}��]Mi�� J|���#@'�����-�0���p�t�����y��c&Es.�a5�� ;k�q��;v�xԻ߱3t��O�cG,-:��,��ġ.�g�����#���՝�I�:Xԙ��GV���%�,#��I`筗������1�v̎�y�F��4����=?Y�z��}H6\g"�Y{�uqP�H'櫓(t��,rI$D��(O��@yw B)� F��a!���i���r���(]Ire0�#9X�UBn�Ӝ�3c�d�;��'Ǎ��3��e~n�.9sgLN\z���θK^�����pL���2��v~�{G�l����b��}��]��>YR�Gd:j�Л�y�����N9���er��@<֩�a��k�=`��ٙ�;�徤����5Ցa5�!�P������3�h�d���|p��|��xv�9ٰ��!?g6Y&8���m�{yh�����CyT�X�	�����Հh)��L��1��ø�������H��@ ��T3�%�(m/�wl]R@�>O�!�Xk:�~Z7�t&T�i*Ƚ�r;�|,bf��k�V��"�┅���{��nK&GӂLȦ�i�8����\�e��w5L&�:`ˠ�a�q
]`�Ѽd���i����܁n��Q��[���BgY8 $�M�l7�]�ª5*�}�s���� ��o{�[;>O%���M��Icp���7�?(���s���z�A��gE����R�W����<QӚsU���l~vY����\����6e��iK�z�7��e�|��#�� �����]��;1hL�߶̀{f�g\R������ˌyr2����O�G~O�[�hq\Hֽ��3	��6��R�����2��^���yo��@P�����;��C��?� r�F�aӲ��7�L�90`�$bk3�!�sʽw{���	>]��Q�Q�(61ྃ��LB�S�hz�l�=��0=s]z	����1+�h ���6���#��U���:��oh�Sl��]��$�h�sl���	����g�'���B3u������R��C�_k�z����1��p5�kD'XH��:�).��ջ?�S�[%��8���S�64��~l����>�vg��Ji�����'`���22�W��T|��+P���=��n��)��y��|�Pvt�;pQP�\�(�{G-��h�p��L�Z��w'�3��^0`$ndY:�����:h>�C��?��{�N��T��%���Ì�.�~>��<��
g��:����M�eI<M��kh�G������Y���X����'����q	`�IMa��AC�)5��~a(�=I�+/�m$�˿��%�D������o�_�y��T~��g�"T3��@��2(�aCP$�?�}�g�0"��q>�$���������h|)9���5SL��� q��!>F R�N"c �5~�nhM]�ZD,�Yu�3׌�,������ҘWZ0�����ѭ�y�����ע�'"V2�7���5j-}%�Q���$��*��c��t��c��]����?�Y����kF��A'�H���N�SN�ٙ��<�38op��Z �5��]}tf_�q���^Cd����Tm���^`����9GpI���݌� �;�����P�b/4a6�fڌ|+��6[t�[��NBc�6��2�kr��;/נ��ɺ�<��445���g#�6�QD�YU��˥Xt�	�lr�����������q-ܧ�T�>��5{g�o"B'�m�<�a��?�Y�~��'���ݑ"z_}����&���D��Y1���\a.P_Z���=S�d��yl~�Nڶ��x3�oϟכ�+����@ei��<A� �-�8���w�� ��Hot�y��{p�Ö�^�]�4�-�K����V�Nr<�Q��O-�f��{L�we���2_�^�-��:���	�T��o��a��s
�VC6M���іla��8����l��jAFt-tؙ!�v*lS��[b^�����Ͻ�Jf2�9�Qj�.8W���Qk$ċ�xW��L.�F	���N c)(L�1��PpU2��� ~>?��wp��zʄýW�iF��	�y�P�T���|v�]�t�
N�]e�eD�*3�� y ��WUn\Nw ��6h�U�����w��6b.���{_��f�~�p萏��%������� z���2<��K3��L�<g/sN���ܒy%k��jd�ή���L�m&�d���q8aVL��lY;�8�u��4���C7�U˯SWi���1fن��HPg�YC��Bh%:>�o��:��@�ޑ7�KP�,=�3k��#7�tn���8m���2��Λ$� �P#2nF�f�����<@"_<;%E����A�l� ��~܆;���2�4���o,�Y��#YKr�D��kT�B�+�}�qdI�גC7�s�~̟/�v��R��gC�;���ݦx}y���e���Sp_��C�{u��Q�R�J1]�\�����8��TGi�q�w���4���m��i�����5�3�q*w�1RB���f�1��ِ����R����'h�_��@ZL���O�� %y!�b�n&�g��Gr�l���&�q��h��,r��U�$�Ӫ����~���1��֔+k���Gw����zk�F?�����w�'���c��s�<���
�|[7r��R��d<��ڤq� e��\ߐ�ۣp��c�;�iq~v��(_��~yǥ{�f�;:�tb����!W�D�WFΈmH��kD��z�|]lwr�y����;#�v��ja�d�V"��M��'�???u�ɴ����o�&��ψ ��APfo�x�эK;ࠜ��+���o�⽆Y8~�-$�w�Y"�Zoݣ��e h�]���(�+f�����`�[�V���fap���<N�=�xFPV�!Jf�-�;\�tZ��6eI�Ӛ��d�.v�^ �!v"�g>�cj{��Y�~�v7y����, �l��[���ME�~�cf��{��P�d|W���:���h4��hu��?r����o�w?�=�Y����1u>'�	����n�pt�ZdzV��8rm�Ϫ���x������,v刦<���:d�#��+i�=1;�^:n�v�ߤs��.���)��(���:�H�^�6�l�!5��;@]���:�G>�;�{���j�O'y�]�sRcd��w��" �׊ҪE�_3u7��C�Ȳ�l�hZAy��j�^���X��ߓ�G ~�w�2٧����s2"xo�4|[f�U`�,q�낂�Iƍ6-����K2�rB��q����ǎ�bY�`)�o��N*���a� �$v�<��P�¹�)(T%���j51�Faxr�Fd�P��ĺ<i��W����n� � ��|~�x�Ch2��-���P�a�s�E�b���L��:��?�0pT�q2�Ec=��;�E�[�WW)�Kx>����͍��]��Y� ��6X��1�\I��pG��_::�����pT<�+�-(e(ipNJ%~�����xO$� ����C+�d�P[�'c3Gn��F��~oߟ3�gV��L��H��N�������_�s������������G<��/��R݀�S����m	%���q��+� �%;K]zp#ѐ�.C��Z�$1:��!� ;5L�T�;�9�.s$�O󞣎��Zz��р>���xTh��hp�:qA���F܏st���s��4iq��7+�rY�Z����I�F�'�gC�����׻�xþNa�1��k7;��s$=<*n�Ěw��RI��?���lN���<�Zβ��.v��\w� i̬<]�ƛ�$''���^^RҺ��Wc�X?�}���ѱ����c�K�̳�W<9A��䵜�����H����G����?s�����v�u���@��r���{�#m�^���Mqʉ�?4-0 ���.�v�-[i��:�:F� �9  .-84��=���<{�)+ӊ�{����X�2JO���J��1@F6��Z2��Y	�y^l��7�+�/�4��^�$Y��J&��M_i5�]���➀��o�.(-���u���t�.e8`;���~#���&�z���F�)f�c[��m�2 �=9Υ�� "|��t��iǵ��q!��{G�86��{�n�3&� ~�����lGS9sTh0Ƞ�p�;J|6d"��0�!�I���4U�r�W��jk���MyK����&�l��g��6�-��V��б�B���r}�SK���{�Ah��#lX��̲zt�^��ߒ�"�ɞ��`�u�Z��x���������Ѧ>-(l��Ӡ8YFcp�{G1�����?����w�/|�T�ܩ��
�	�.6�@f�F Z���^�t�����m��s�������q��P��Y��[s}'gٽ��^���͆�q��=���J�;�B�,�Z�����	�^�ܖ!ߕ<7,Fr�����C�ϔ�45i��d�;�urR���Yjڡ%����7�ynԼAN�=��߯ghl���􈔍���g8����A�4��*�y�y�b&ɜ]��pt	L58*4��+?>��:�߳����ya �\ȷ�?�m;�.Ʃ�����)՗F6��b��Fl����P �F`�j�&�T`Y�t8�n ���K���]��[N��|�u���;:��/�է2����Ns�H�LQ^���8��&�g�+��������|/���������;wcw7�����s�7k���\�b���$�2@ȉ��b�V=ʧ���8f�35c�Tv\�,�,X�c7C��nӚ��l���>��R�$��`N�N�w?����1#���; 3Jq~��h����V�&��Qv״�N�{�ڠ̆J�-�`�O2|`.�w����i=�a����sD9����4�ô��W�Z�-����	�`���������%yc������ ��ts6H��6�.�{�[��0H�a6��G�pD�q�l$oX�LJ���#2�Pj���"{I�<�9�wdY��c��f��gy��(�?k�<g3��YpM۞A��kI�B����ě8�^���|gp'���KG�vC'�ŲH�\BǩY<�r)�ۂL��q�
�~��o�ʗ��Ϗ���D���s�x�yH��O��~�A�5V�+Q���qX��7s'���r�z�<�\��ۚg6��l%�9�����lok#�Qr��*�A�z��]�ap���
���鶚G�]W7R�(���ɡ�. ��}���E�q�W�;><o�ϰ�F��%њ�{�'s�k�kR�����<�[���~m�:�<�R(�d����:��l��:�<X��uO��@0�$#@>��r�F�������
�k��қ�?�dX1����{����:<�����{�H׾x������l�Tؘ�{���tב�}�^B�0+��$�-oߝ�4�{!Qk�Q��9�w���Z��2���I�Z��/�
�}>U�S�(ԬO��{�[��*�Y��<�fi�/��g��#�k�)Q!t��X��C����AS$��ʸ2p!Z�|�����U��z����X����`��\�X���4��{-/�x��y�[Z|�M�o1��С��Ps���a��0	�0����"Yh���n�[[Vd%�isQp@��d��%������W�-�,��s��ʶ��,�*%���5��w���CѬ�O����;��f���!919U��4�=�W)�Z>7�J�膥�9z�--꺳Ie(O{:��١���ͧ$��:4�!\}]����R:�r��î��r���?#��5tջV(q�1���:����~��wv�f��9G��?��3a��N��)�l ���:�k~��_��|�iw&�Εs^��VV4l�E6"s��K��m�@.H�l���ꙷ}vV�F7��[��
&PL���|�n����y���e��;V��{#GA�!��S��x�1�}A��<�vc�?\�/R\1�|p�Ȃ9�����ߐ%3�<�s�|����D�9�+�yK�.)rJ��<�����9RN��L������R�( ����#?ǷR��1sA>#��f\-!M�޴�m���\ ^�I]`���˺T!���sB��²*koM}V)��J�:4�Pk�tcm��;&��p��c��|��vz���S�������KN�N: �A�v�8']�X!��L�3�]��bv.�8UdM�y/��(`x��N�U����zE��d�'Y��g���b}��9A��%����V����(堏�%�����-��2e��pZ�YZ/L=��V��v�����N~��1�t~'8��$�+�à�0T����v�X�Y�,)r���2D�t���l+�;��7���C�X����������m��o���(<;܆�>�h
S	`�&Y{~���a�{������")7��6��%	Q���N}�6|�ߝ#E��G6��1^�@ף5D��=2���R�d�=�u�)�%��po����|ri�.=��L*-����[K���N I��C��s�&�֙�78�I��o�Ȥ�C��/ܸ9��Vq擝����w��`K��~�6��ωLF�@o��E>��|�qH�c�.�<|O�Ǣ�ƍ���ks�cd��gq�Fտ��ySHC�C�+�Bw^M]��֬:d���cBt���(�̀0�e��vb��z�ef��k�d�G���B�2���ڪ)t��T�!� �T;Gs^|z���<�A��)��'���+!X[�S�������+�b�h�M���~4��Po�2NƏ.�Y`�]���3rPK^�f���	d�2�/:�A�����җ=d#f$f$JM��q��ʯrC�ߪG49���̀ �9��Y�=�ާ��Go��r^7&Ӛ;�YDnx��7Ki����h��`��Wx6�����˹�ܞA�Z]�Ώ��V �Aj�h�;G(`��+�;� ��X�Ս�G��|ǹ�0�5%���W��0;��z2�ɣ��X�����]�����;;3�����o�{��Dr���X|OVgޢ$4�@��e��-9�s��u��ή�46\^*�٠���'��	E����O҉E��(��
�������%�u΃v+$f�r����1�3�X�غ���_��}t��X�lȲc>�ñI�<��x|��L�q?�Qf�b��s=r/�:s�w�_��J�u����H��C�d�;�L���s�-����̡ƲFv����Fo���44�&���?�/�)c�vED���ޙ�w�P"���e�in9�����|R��E'����NX}�R��N#/�@��Xk��e5�b��C���)�,5J��W�YRٹ�e;ǧP姯t�T�d����]�om�Т���/M��f�YV�Ԟ��w�@��y����2!6Aិ�q����c�����=9��v�)�O.��?��"�F��A?��}����	k�;����Γ���EHU��� ̀�}�w���2I������n�Y#��YY�T�ׂ���u������͹�;�������zM��rN���7WLn2�Č:/,�-j3��@FZ�R+,���L}aOqz��n��v�_ǃ?f�Gf�r Y��ڰ��<��w:���Z�Jh����>�&���#�o���Lf�t1P��A`�LE���A���Qƻ�2�����z�l����ߖej�d���K709�D�	g��x�&X�Ao�@V6f�Em�݉�C�:�Nmd2�A[��^��H�@~ĕ7�C�{	\�Q�3��������𮊴�af���8���LO��!d�襢��ٌ������w明�8�%#4ؓ񟄉w~�x��&pE]�[�#)�F�<�쬉�=Ό�먅\1�N��a`0R�����i��S�*M�y��']���3���?"̣����&��	^כư��İ��ߣ������ϝ���l��K����h�F��������Q�����j���rOٟ]��i�^+��p<���:��k�����"L��,�ѹ�����	~��G�<�uw�c]����q�4涼��7[�>==���Z��?F�#��7x�0�9v9�z�8g�=O�����OR,s� Aia�?�b<rz�\��%D�����y��{�ف�/?���QΆʽPx���K��!W�C]�k���\�ot�������|��T�.��+�,_oa�������k�e˰)��;�=�b��c +&�4�Y�ju�	����H�{@`��gr������gȀ����|��{� ��pn&����ap�v�s>q��،��=��8��N0��q�ϑ�aqG�]�&N�1&����d���R>�eU���}#V�����PYdv�l���ݑ�ɚ���-��ތ�gEG9��߶rZ���껻{��Z�����j�S���4�)4�۴5� ��U}Vw�X�g���5Ɵwt�t���y�s˼��׽�/�r��N�2��,r���1@Mu�ex�3쏸5�	%����w�.�pl%����D�q#�E%�R����;�w����ۮ�\%2.� �E�e�?�U�)Qd0��`C!Ww�Q�_ܜ� 붅O����d=�E$5�����RR_Ζ��:
j�<8 ��t,5���s>�Ӊ� R�u5"2�G�cZ=��.�zq��N�ŵ�䝇���$;�_Ҁ����jq,��������'(%".�����@�=�5�1`g�H�35����i�}Ǯ��,�����j���� ���U�Z������݉
���3����yh&�C�~�z���\k�M���;ON	��pJij��gjQx��QTtJW�رS��gAT��P�4�NR�a̓�ቇ�P����M`�T�exZ�*4f��&�J�kPԪp�#�q�S���w�}d�)���,�玡g�V1�A��eĠ�D(gT��M�է.�7�9[�7u��t�k<�]o(��Mk�$�t#q��]N�;#���B���P8�Q�޷����kB�g���Z���S�w�ɿ����=�%�j <L�U\�@o�d�����,Ģ`[`�;��=���*W>/��g~���<����j=���%{㥺Lq&?�P����oo�:�w�t��iN��0�d�[�l �V�AA�;u���{��E�DL������<nN[۠I�ș���>�{/q��9B������;.�_a��9�m�gY���_�̩�!��,�Y���{l�ʎ�"�_��F�-�-0B(���W�1�f�i���u 3�i���mz�
d8��[˳֖��[G6��a��լFMwO<i�Hf1�Iþ��/ڟ���U^M[�#0� ��3��NҌ,��6���s$��j*�Z-��M��_9���i�ɬN�ҭ^�iZ���5�/�S7�̱'��o+Z��)2����s}N�{:�h�5tr�R-���ڭ����B�ܛ7oK,����@��:k���}�%�Ȕ�)M[�ϣ��ʩ�d2dNά��u��L�	�fL��,h[O�8��ʒ?���/�z\���4xL�  �Ƶ�����"ؑ��֞����69M�ZJ����@�ܚ�ռ��L�]��XNJ�zV�St�{G��ɼ�{vY(��7.ۂ:�����uƯK�}뾇(�QA���%���ͯ%I~����}ҁ�� ���a	��?�j�^�R��p<�Ou���g��1�9hڑu$O�{RZ��ݬ����c*B��*H�M	[w�j���q���ů�!����J����|�ʰ�D��X��FE�&�h�Bk�/���6W��7p4�>�a��iCM�T���5i0CK0��\Hp��bx����)�B������t��2Ħ,�.�b���b�hz�4� �)_#�S� ؙѶ�B~�-��5�V�_:"�!��� ؚo���������������Y��z��E��_:)R?�'X������	��ѳ�B9.�,NX���c-6��q����p�r�m�I�� aP�~� ѓ�����������|Bx{qE��k���j*|?D�-(o��n	VC��<�?�d?G-ۻ��r}ڒ����7��Z�#~�C��˹<�`ڹv�F���g",~��a�4�� ����_�qY���;0�s�9�* r.0B��]	2��k嗃�V3Jÿ���B(�^���Pv������JO-�g ����^ߜ���3�|�y�k^�SV�5��Ao�(�"�!��-E*d#�Ak���?(挠���M+�j��=H���:Dݠ3"&���퀱�n��5rΩ^�v��p}��܋טDb��	)�[�y��A}��w3�g��GV� w�*C�	w��`��N6�H�H�D�0��E�-����� �)�V�!��ݦ�!�@(T���)�<�~��R����϶a5�?���[�Pt�R�>�麌�=bt��뤑R
玧 ������\xm�t-_���Y��=����(w _����>
�b/����ip�����IA�)uG$D�fY�o��A8~}q�5���{�e�z�lI:s.@��� ��ʑ�u�R<!����X�!T�ok
^���'A�C��{{ڻؔ�M#��E���=���Y=�ߝ7�0�wc�&���h0����u<�H�`�\d���|�6Y7���Lk����{�q�ׇR���H}��]������s�6h��"�x��.���|���MÅ;�� 
2S�g�?06�]\���ݍI�����MΘ7�W0NXg�xl���3��X1�.J��2Î1�k�'�s-)17D^P�Dj50�Ac�Z�ew��C�� �hQH���+��q�P��9L�_#���%�N
��*�ݵҺ������{�=c��5��/@'�X��-��]R��ܞ1���|g�W��T��x����L��.N�Js�
W{�X[}�6��W8+Û;[����F�� �f��8��B�9ͱ[w��H��Ϥ�rCm(�!�oݸ���� Ƙ�Z2ja�"_��v��[�(R�<�G]��F�q�d6�7V������X\�$�1e�Uɿ�ҶZ���q�O����Y{��H�fE�sݜ�zd]�?����D
��R�i09�)�+Y�B�CJ�����E�����0шL�9`q���H�z�rd�yU��;���ZOE�}Yh5���j�ke�ҕ%�y���V�ε�
����>aܪ{�����= P��N���ʳ� ��fkΡo]�>v�Pu*qy��S��@���c⫠W���A�u ۝gbLi|{� ���?q=D�3�$��:e?��3���@�0��[耺����>�����L@v��ޑ� �HQ�J�q������II���V��;�3��x�UAd��ٌe��lҶ��VVB��OK ��ec���:�zu=��������ى�W�K}�⃫Ra����u4B��%�t�
��������(W�י����ql�|Y~�,�d�b��J�U���N;R��K�s/J�L���e���DH^P���t��������9�0�W؆���7'L�]I��"ЌOx*i���}��TgF�ZQ��䠜�<c B�Iii�
��7BAw,/�3DLh[<��q�^Ra���nZl�$e�֐Hn��!+bY��@�0Fa:J4�(��B�gY�}��� X��H�%��|{{L��4gW����{&��#blkC�Z.c�Ӷ,���F�跭I�䍴�n:�2���ʙ�:G���j�hz�P��&�P���g���zӼA��_;:�3Mnl�n���9���}�r�(YgEo�x���������7Fؿ^���o�Ɛ�;�e�lEs4FVVvҿ�=�ể��=�[��(uo�v*�t��w�2ڕ�m`η o�;����,�����Y�	�e�ɔ9�.��{�c�w��E��x[k�dL%��_Z��������ci�.�g2�#{뷎-�����{rI�[�"����ԃdŔ���4�׎-`g�FW�ų4�����!
���ۿ��e����\vd ž����՞�6������m�噬�)��t��Ð�����)m�ѥ�E���W�Pg۸آ���h�_�5��u\�b�e�:J6����A� h�F���:��Rt��h�Ӳ~��M�*Q�?�}W�v����ctdY��T`x�{ṐB�}[yΗ��{d򮁓�X#@�g��vH�Oj|�ZP�U����H6Xz�vFV���%� Z�9㱥�X��bZ[�q�ZV�gg���@�Kf�6��֡6O�:JHT^1�h���U��$PP�GB׎Ț0$3(�w������]�����@g�y��'�@�R�?���߇�����Nk��o��^�6��	Y`��|�����v�ET�>��R���к�1��-��Ϛ1��w�0 	<T#�)1�{�:Z����W<���V0gw��� WU\4rZ�9m%=s��zIuY#����o5*��ÿ�p��`�#����ި�h���Vu��:��q�3�8J˜J�z�v�B+<MS⨔I���h�':	�iVWk��v{Kt����[�r�b?Z �@�����Ha"[���S��\/��M (B��yB�YPhPZz]t�!��H�ɍ�?(��0ۊbQ1��ZAuݚz%%���6[HB�em-$�h����PF̂���	xkȢ��4q?d(`�z�Q ��p%_K�.:7-�!��8�K�^ξ)�p��7`4����t1!kR�����c>T4���ht��
��9��� u�֞�8�aU��Q�3Z�U,�Ct���Ѻc��/.e�NWkE=?x-��]ti�
��0NJ�ߣ�!���:!��<��ͱ�r�:�(���h���-�)�����s��4�Sg�H/����;�K�?������ӝ ޶Vy�~Q^�=&�7F6ϋN-s�Zǟ4�؅���	��YZ����#��}���g��{�z0
�_��
��L��k�>���;��n
����ک�W�at��[��w��^K`%��4�x��c�C�{+�b����w��［��rN#K�*��:���8X�[j̾�h����k�8���{>rM�.�h��3p.���]Z�[|}�V��g�N�&_�jm�YQ�k��1��8?�H���J��� oÇL��{jz�|]	�&Ko���G����WJ�j������M[N�s�y������$���$m�W�艧(�;��|�����~ �aM�ހ���1�Ɠ�a�3��垽/Oi�!����ۢ�M�;�>F�뙗�/���0Z��Z�n��`>OR����?9[�.93�I�k)65����9�7u�#�c^�xΜԷ��Z�]9��^�PE�=@'_�xo ��3�ev����L	�{9zꮇ���m��Ə��,���yG��z��a	 �σg�%t���e���D:6�i��'Z$������8��s�>�R���f�K�(�m+�����8���4YT�Z��@����%��#sv��qP�d-jr8�5,P�Ϧ�6��\�->���M�8��\�����^!���~n��oZf���o Ґ}a��5���/LOx�d<&:)G� �ZSĬ5DB����$^OKy�u?��6?�5�
���?P�S|�������%z��s��,�P"͸K��8�]Bˑ��3�E��\��0�����>����Sl賶8�DGx$-����� ;Tqc!��L�S%�����v�r�~m���8�1N3#?_�;l|����ʴ	+(���bV+��Ǣz�#0"�[&Be����n1�-R��ul�Ka�C�+���B)_\���s���y��
bV��ʵ�08�ƙx}�P|a��|���7�)<XÄ�J/�\���KD�D��R0A�z�(37�1�+��eO����{���@��D���ӗ�
�+9+G�)��@hk�,�2(֮�`��__�i����.KŚ��]�b�8L�'$�d�`���g�\vES��-�!���13��LQ,��	�h�>�A�C$9{�0�����<-�m�Ϡo9��bأ��Ssťd�������`�G^���Ru�Q�lܻ���k��i8�A%Bx/�; g̳t����`�h)����}||����3}������"��@稑
�h���@Cn���]j��:{JO��E�����x��<�ƮU&�9�;[@��(�JQ��ǖ���Z�eШ[�8��A>�y_[��NE���5efO�Þy���ٺ�Ҩ��ޫ������|�*xO���~d٥�t\�;+�m�6�7ؙy�+�^_�d���R�PҕZ�����<�0a�7�5���CTF�5�<U�D!o�5f9<�E��s���pZ�t�<�m�,%MmJ����b�v�'���&���v�"��Ϛ�������#�	:H�q�H�^��e
j1��5�uB��%�nV�!�$eG�i� p�9��r͢�SG�Q�8�/ִk3�֥���wu�����LnSQ7���Fꢡ���;b��,��E��Q����ׅ@�τlgiq[ a���;�Jv���խ��~�kra	>�^��(��v��b����7�\��T�m�
�6&6��uu����st��9!h}�)���U"
R\���R}�]~���R\[BKɲ���k�NU�V��k�ku���pp��O�l��
y �$ϯ��>_-�=7\G��5)����G��:i)n��ﶗ���_Z��i�����C쑛J�ul��W�Zs����}���#Jtg�5C��������������_�t�_~UІ<p��-��W�48��(�3Z��	����"�+�CU�����5�l�I��w���֜����3͟A��礶ͬ?�����?��C���a���v3�;����ut��d���Ct�#V0
ʉnO����#}�� ���l����F7u��aes��%`��pw�]S����L�j���.��ȍ����u��5���ć\�\�����r�����<����D!��v��7�z^.�`y�y��xz�%gM��bƁ�{��'�J���#�Sx��\aa���a�-��("�_^T9�iU�I��g5 ���B���¿\,���ENS��qK�O�B�#1�ù�#r/� ��t���l�4. 	�egxέ1X�H^&4tM�j�6R\@�ʙdY T����ۣ�8~,������O�s����;m�3�KC�%J"R|�jN7؁�Prkva�K /�>��� � *�"��L�J�%Q�!hmg��޿��0��Ʒ�ޫ�N<.�8{�[�G�t)�%� ����V�'�c6�)3r�nd�C�7R�����|'G�5ya����v;m�޷:v c�k��3{&я��re����&����k�@d�,����E�1ɝF��M�kG��]��QR����\���|ͼX��b�Z�}�n�u&F���(��1���o�E
_��^��8J�Cw�������'�|m,1љ"`�+��U-�bOw���Z�CK�`WFn\W7D�xu{(�n/d��Y��Mm쬎d�CY,)}b1���a���(4�&��W��ϡ�C T6d�B�C�yW�x~����jn\ol��9�Ct3n_+4�:��o]m0�:��S�������ulJI�~>����u'�h7��(�/S"H{�%��\�J#"J� _������k�&�(�[g�<�M�v� +󛄕�%~W��6���]��7[��陮s3z���7�\��'$ZDٷ�K6�I� �t��:���k�֗��e>�ϕxf�(����l� ��އ�.��4��bV�f��ׁM���]@z*����l:����O�ǵc��o���En1������� ��ד�>�|��P�5���ٴl�����������^-aKH3�,'+*o�J�W�{t���A���t�����nԮ�(ԋ��4ը�8P�U�:��x>��3;Uo�ҡ�!��׋WfT�x���Ӊ>|�@�?���DqG�&]�;byh>�^mΏ�n�;��5m���N/�����NER�d��Tx��(�c�U	"�NN��9#X%�e�kfh�������D��˭!'i���F��31p��p7��?c��������C���Ǐ��>@�\q8 ߙL�������ؑ�󺰧��-��S��e$�	hT��# �x>����r���;�p�.�ͫE�pڅ(��籍����=�
�k�"��s$G�R�>z�i�q�}��}DZ�E��#Ns	ʕ��ٲ�  ��; $���NBv�aj
u4�������X��7����#+�Hq轂��9��T����C��	�I�ѣ�1�H5��Pc��fV�>�z��K?8R^�����J
�*�
�B��#ܛ�р�0#���l��M�}+������p�O`~c���ց1`~�iz�`)*�:}i���!BG���eQP/�<��1+����)�:�6E�֍��a ��8j螵�:O��4y;勺�L1����W�<�ҿ�:oo_���n�sbO��ϝ����<׀���������\� �l�-ǽ��In.�T�N����Cֈ�2�)�w�p�����O�kH��=UÀҮ!�Fm��%_��{��$R���{�q/qC��yMt��O�l�2�3)˵��
#=�K٢M}�ħ␕;i� ��	OL��y&�с)�7�Y>��&k:!����ъv/j�"�8�X�K���Ʈ��2gp���d��	�o	�>���b��_�h�u���c�&�u���e���Q+�-t�\ �5�7n�[5������(� ��t��a�b+�4���K�`�$Q�a�6!B��s�s��Qval��x�Ţt R�\+f��ދ��s�Lk��H�l��[(gx���*Ϗ�	MEli�����k١9��>��~8yZ���V;e�Z_�z���h��.'*�%��(�	^D7���57ﱡ������s���[��-ތ���Ӽ��i\O X�=���Qad�.^��o�'�}[�j�1wz��"�����E�;Ե��k��}����]��@��L��F¸�a������1�k���J���9�A�U����G�ᗗg�����nN7������#}���N�Ro�qNS�z�����O�f)��.���EU:Ot�9������?�&x�2��C���c�e~��@�'r�"�L�Z��>	�K�)2�����&��eE��:(ӿp�O=�x(�n6?��͍����.	�-�IO��A����bX9ŧü.ö�ҫ)����1&jOq/j�f���ʵ��Z�1�ZK�0=�KC�_�t�H8/ "0�T��hI\Rm���:+\�z�5D���eK7�%	\|��`t����3IAD
E
ㅇ�r���e����� �.��[��^�bF2js�R6��O����?{�zA9��A���j��9�^M|����g�j�똪)�=x��sk=3@�O���!j�d[��&��|7�9X��Bȷ���~%��gZ�|�`���Ҩ讼���`�喾8�����!<A�̯9Q���H�N�b#D_�t�{ܲQ� E��8qx��p�6s�ה�W �B�������Ք��i1��<�¼�����qǬ��b��W�W�G7I�>�:�gub��Oٛ�m�W~�e�z~�M8'�����f�M[�Lw�z����47"�S		i�F"ǔ���x�7g>�;@K��#�9TLzͤ�bK�����(�2_׀�v���� z��ׯL%1y�NN$y!�Ѐ���ǭ�0>2���g ��n�l@�[�i\ͼ�y��<]rm�����&ɶb4QKg������j���B��E�	M=�_u9N���z��Ƭ�����Z��YU8��1ս�VI��Z�ҹpn�A?�nm�K������%����H����}���$��1�� �!J>jVql�ez�9��8:@7jϦk���8 �9���&zP osH�B|�0hA���NX�K� �Ԥ�[K�3x�i��nl�}m�m|���qIo�st$�	�uEɇ�S �����/g��%
�~�^Y�R:��;�����)�	|X��}7�j�����ք����I��5����H�y��4uuwܦ4��
�I��)5�Y4Zɾ����x��ɏ)w�Y2^��0���If�3���FMV�{6}�>?Sy��E��sN#g=���������2��~�B�>���fR��uє�b:;w��bt7)�ȧ�,��]�!	�9�q8��Q�P�P���ۢ6(�`,^����tvҊ�l��r��'��q����':?��sSod�@/c�{2����NЬ��{-8:T�R�D�X.V�̈������!:Qٚ�?ɻ���Մ�l���H4D����y���e:�.),��kըKl�����i�t�AN*��	J�W�[u�>�u�&�����CZ�����~6��j`�O�U�传A)W�4M�0
Y�ctȑP�N(�y��?�ͼD����)j( 
��bLPK�ҟdD��e���z����N��Ɉh�,�y!m�;����&�e�p�<@�͊~����'�cJ;��)�`إ�^j���V���\�s$݂hO��~��ga
��c��Jh(,z2��n|������ysᆂ`K�:�n��]i�Vg�#o$:�8=f��������?o�n��N��"5r��R�Bc�=�»�Iç�F��<%�<�^u*�"�����\���5|C,�x�>�y��nd��?!7
�&,ݾ<��nV���̟9���!��˜2u���u�;�:9b^����e#������u�=ƥ?Yn�S;=��ۿ2���R�9`�צ4��tf#bљ�_0��=��-3�z}�-`���lݙ> ����"�s��Q`}�?���el6l�[��^1�\��?_�C#�L�3��� @�M���";|p]&�<��J�^��k��ۓK�k4��aD�e��w ;C5�vi���Q+������~���P'	�Q�<@'�o�Ts��c[�dt�k�Q����u�C)QO�?[O���ÀB��	i!� ���w`����uR���ꚴV��Ԗ觔H�ã
Z�%�{S�1R݋ir������5z��P���@er��,�t�fҪ�����/��H�5�% ���#d+�_߲x[���$�Y붆Mr�cvݬGd@�5�mDk��:	�����:z̩��ݽ��G��:Z)��Y���2O�����ut�Ь�d�'��lm��Zcǚ*4���?ԙLV������m�U~�US�&���i���h��J[B|>G��{���P���c��� `ݛ�}����o��/_���p}z=S���I������"�4��j��IѴ����C�]�{(�z��0��6���+v~��DD��F)���1R���5�}ww+ia\!�����ǃ��2���Gw>H~��	�#7X�z�&+=���0�<б�۷1�rI֦=�3Ȍ8�W�M���^1f��
�b򶊗��������>�s��� V5#�	�A05�4�HR6P��ES��:��y��6 ��=������W��D��T���3�~����C��g�`��QJ*|x��Q=�/)��t�R�p3x�B9<uV��=���CJ��[�R��Go���LV�ѯ�~
��R�����;��ol�@1	,��fľ��KP���a$,W/��~�c�2��`������[��	a�Z\ea`g��j�%Ӳ�����c|� 8G+"�>���
E�9/����G�u��ż5:^{,Q'.�^#����a��l����}���q��$�cﾣR��RG?�u����Gnz^=޸Q�;)�p�|��W��;��o�:1���K��D��L�|�ڼ��ϕ�ì8a��9R�tY����Kӂ��ڼ4w����p�]?�[��OE�`I ��\|`��\�����J�`yH�Rm�%?}t�w��M"�[�L�;&ھ���=��4�J���<���\\k�g���5X�����χ4-����{� �a5E���P6�	zI���G�G��{��o���]��Oq��l���'EϢ�i�G>���eS���9PYtw�;,��hp�l���g`��dL�܄�h��܇���ԅ������yQ���[N�b��koy�N�N�+Z<a*!�u�s�j����k�_������W{��6e�͢���mp�GN���s9������hP0&;F�z쁝X�寫cܐm�{��B/L�����obx^�����-7>];�|����Ƈ%"	'�@	�Nӯ4��b4=`��,�1�;�����R��֗z�wZ}y�,��br��A���lH��E�ř��BV ����/�`��=�N7R柿��~��W���+���]&���2�� ��2�R4��E����o4�;>���8�Ch������Il�
!����ռh�Q��Z�bfc|V�X�b0�~~}��>�D?~c�������я���R���_�h9��ݽ�G��GI�ωn��r�(⤛�l�(������T�S�T���!�6j��oSc����A��]`0�e�`�����h�!��	k����n��8q�\�_/�V+�3�w��9�,Y��S�F���zAg�F�P> �	��+\�i���?X�v@$w�J
|��G�L�Ǚ�;���3�#�����:����\<��<]��)mrPгa������0�������k������']�o4 f�92��I.<�E)PR�3��L�͊v�m�P�%���|��S	��N�v\1�D��9o��׎b�`?���U{�.4���P�x�Iw,cPR�풀6l�簐�ֹǨ��@+����F��QJ9p<���߾,�ޔ�f��烜�cݔ��Q�����I�3�˿r�~��k{ş��⋔t��{��U6�kx׎=C�%?\�n�v�h���d�<��Cҙ
 ������ �
�D!ګ�.��Wq>=�@��Pw4C�Ev �}W��ЫOw�p,�RVc��J�= ��h�c�S�ь 9#xDһ���������%��'J�*�sHA*ݒ���4�u�\�ۼޗ(^��2�����P�	�����z<8��)p=�r{�t��W��a��p��,ׁ��9ϝ�|l��ua�,�h:Z��p�.p�=7�|���f��j���(�x��d�D��
�@W�F��[�������F}�����/��y��L��Z?bT�E�'�[D@#����"���� �k�r"
�fy��)@���a�fh��� "QC�fjLW�o����M�Ͼ�p�z��E'ʲh��H�m�0 ��e��|fG`?��Gx{Ğ�s������#��^7v@g��Z6";�S�e]�D�(Sgj��4�	����-�-:`�1���(��I�����ge[N��{JǏιu�],Ú0���Sp��E�o�m���;�g���.���}�đ:_�_���/�pwG�����¥u)A��Z������"Q�������T�nE���,G����P��#}�P�-��Y��8Lo*l$ʄ���.���GA���飌���o�c��d�if�|>E�'� ��=y�0�qs�"N& U	� �dB�!?�ZJ:?��E�@�oјR��-�e��v��֬8**�+s����ەk��nN�:o��_��"����3�}��� 9\uŗ�z���zfP�D���)`��4�w/���0�T���/���[17("��M�A��V��$������.�/`;ZLV�]f-�b�ʇ4/��,���!�v��~���y�.���m\�<��!�����G��-Ƙ�3�>���Bٖ"��E��Rl����j,���)ed������KZ��J\��E&
c��3���vW��</ܡ��
zX�`�[o����Uݭ�8c��tnQ�P�롦N�N�Ѩ�U@�
�#�8�'����]İՈ���k�h{�J��ђHE���+�02n"�׶i�U�r�n��]���)^`oEK����^P����r��e�RϢ7�{��(���d�J�q�ź���3�4��mTbرyb�q��]߻N��+U����K�7�=x&��U��B������ F?O2��ۭ��B��WK���Ɂ~ib��;�9R J�o_/�7��0Dԩ��W�aw�s���� Z���e%z�<�h��_w"��<(��6���%�y/��-��P�/n�C��/.����-������U�D��QO��oD؏�ƞ��E�%����!�[�5��R*L'��_�~㖡-:���;"��͍�[�<���qR��;%�b�."
Һ%����T����լ���Wwi���GsFKR���&�z��U�����{���2�4�N�^۾�Zv���� �t� � ��e:I+n[�	����h������u�c�i�%�2 E�<z��N��1y{�&A؟�B<e,���1h��A�Җ:Ӽ�ӱ1߼��MG�����k��\����yK<V �Z}\���ߨ���";4�?�X�7���E����ӝ:L�e����>K��x�Ѭ�ڮ}���wӯ���ų9��3�/)���,��+ ��/	-$�?MQ�
� �F�;,��ιv�j!���*?����9hƧ��l�:�C7D���j�*?�}a�0�3إ������6�9��T�e',Q��,s�6������?���J�>}�r
<S�׋�����%pXW?�jç�64�OJ���+=���(�<������<��+>%��{���
ı��I^b�A�)'�Z�pj����g���A��E0dZ��.�8�!��\?��٘&�?i��E�������v:i�
�]3��V�#��9t�_��:�,
E۴m3ٌ�o�3�>Oc�MN�9Ĳ��z��Lg��|p-n}�����O���}^��y\E���n�n��˨T�x-�&rd�h�\�S��kT�|�ׂ�=���y>�}��,=�+ſe�z1d��`@HKK�i�p��
�	���nP����%��e��8i����*�W�[���P�H��Fs%O�t�Ä���r�4N>�=c �Py� p���lKxN���Ƶ@/:^�>@�Q�����P��2�׺� �m
X�m�\x�� x
�a(�5u�H�r�L����0j6 lh韾����A���Ww�8e��<�4JG���=��6��h׼��:Z"��D�)Vpf)2g���E)AY�j
�]ڞ��S;򹋴�yX�x�h�z�tw��+i�I}Xer����V��{��S��є��{�^1�/�3��	���l�Q��@�3�P�2���]7���^�@���"MӮ�]�Z.f��F]*��PW+�82xp�vj��A:N�s{c����WZ�e_���`{B͔�հB[W�+�hB4��⑾�M�l�d��q��e���EP0G=�<��.�`�U�KOy��l�w�at�a��jn�<�3�o��ƶ�ح=HZ+Д�|h�St �������&�*�S�}��Hϛ&����kc�GZ�T� S��N)U@�ɐA��������wi�
��Lon���Z�M��a��]�-�o�ܹ��c�WkP��-�E
�5�N�ŗgChX�0l�����;|�Coj�3�}��.P�G�Le��#���:��ɺ�w�.[�u�Uݘ��N���gk=dF��cs�a��yS;�kR\X����� ��ĕ��,�I1��D���-؍PaG@�!�eA�����A=S~���$�`��K+�����:�4�6���7@Ɩu��Ҩ��;��@�����t9�h�����8�_�~��:dU��Ѽ�g���X=X��5�("��(�y_6}�F&�v-t��G�NcvB��嚻�ۊԲ[�Xa�	�Jv��*㣃� 7����B�m�@-�>�����N��_��O���_��Gv��0�Fz������J�,GH=�=9_�e��3�wͯ��IlL8�PmB���*}0j�7����uĠ�v����E{z|tE��o������a��Er��kp�2!�҇E�9���r��fG��H�I�.iú7�s����wB��)L !z�K��pk�	a���[~��+�(�n�=|���=><[��؈:��Hg��
Q��$�Ӊ�:{E�Z�BM����`�PU�����h�㷢��Z��J��[��A�wp�
���������<���Q>f�d��1���O�h����.��e�x�<b�sڀP�+������f&�yW"E�y�߯�2��Ƽ#�L'	�{F5u
�F�%OR:�{o	����Aצu[մXqI�.�jt�7���}�<Rn4Q�#VŽs�%�,b�^�zƊ"�*x1����y�\s��NkM���y�A�.��) �3�Z����cJM
Ou�m9�v�m{��r��.�8��iR�;���w�T	w�=��}��4j�ޓ�ɏ&_��U�w>r��@1��1hj���d���O��eJ6��>��IÂ����<��"�|������b��4�� 4%@e�P�ns�IU�k)'��snJ�h�9�5��Bf�m���d��S��)��a��N#���rq0�d�]w��tos���X��5c
rW�A:�L�7κ��МG�P��]hu�>rdͯƫ�Ơ��6$�b�V�ڿH_��hg�&�n���Mp1�,
��D6�
;�(6J�]��&t[M���D�� ����r��s�����^��t=u��`Ǘ�~ѫ�u�e�l�AFn<��ⷑ������[p)��xXǟ'��^�0N�i�r�2�S���荗��w���W�)Xϣ�j�����j������uK�\όI2{KA����T�n5B��J�R������.KrY�v=����̆����p@��OX�X���KJ��{�]t��Y�D�PM��w��羚��-�5�������޲lm���u�/_��.�E<Z�D%�'��p/�1�2�P�3�u:@.+@��2������ynz��qyK�Q-�ҚQE�!�A�<�����\7��c��ӍG��-Ϳ|����N‖��,؁��"<�"��x�5 �y��xz�����Y�|y���֋����7?���;��#�N 2�)�=|�cő��ܷ����������>} L�C�yQ��n��y]�rk��~�'���o��/�����
~�����L�Zh�牋��J$�u�A����K`G7������?���*��Jo-�����@�x#���<=���g�V�0����:�V�����Qy��i�TP�h4�T7��#ze/o�=a��$k���J�':5k����I�QԘS��B!��Q��  Ž�Dn,��5#�#�6U��J�a4پ��oo����
u�90 xo�{W�n��&��EM��=ǸnM�k1���(�R�������P��ߚƔ�BA���4R�}<N�l\%	UxF�� 1�X�</��C�"r ���:3���/� �6k�8ZD�Ţ�T�o�T6�<d�	���k{n��-��+\�.��pM=�F��pÅ���דx�)��&c�{��K�� ������  �2] wV��9j��%z����qM�_; ւn0���㙘��g�cÙ�粒L����&���%�O�i*^K@�5mF�݋���.[E*v�F�,b�� �򓁝ķ�������a]a=~��{գ�f���H�A*�&(���wj����/,�T�W���<����>��:O����cwe��T׏TC���Am�|��k!�|���j�^� ��Ɍt	���p"��r��A�{��ED���W��,ŋ+_�絊�&k`GEW�w.�v?�Ϻ.O���>�*�������n,��w�΅Ȫ-b�1���,AJDg���5�:��h�bE�5� һ%j�4s@i��S��u����'���ݴ"R �
�^���@{�[�f���dp��R`vt�[h�P@)Qk9��*� etźqt��	m-^���,j�T�8|;���l��Q�>�^����HM6n6�83ߗ6���S/�X�9�H�tٍ�lŔ�7���� 8�,Ҹ�dLk$�ƌsq��p\.ge5O��J�DA#Z� �Ѻ�Idd%�DZra�������@��[��/���/���ׯ�������Yj�0�#�[u�ε��G��m���� ;�<>?I*��ݫ�
j����a�����1M]h�V��������FP*  0d���!�}��Mۜs!�ּ��YB��[����L�R���I��|ޗyr�����ժ�-y�c3�u���B	�gm��w�a(���imro��(�ń��f̏�O��?�.��]��]h�1�IyK��+������pun&�����{�/.�ը<xQ�\�}��5���"�T+-�x��"�
��9��A[-���C�O��5�u�=��0�����_`�����`
�w5XZ���y��m[Bc������n���{���^���~K���uIE�Vת��7�`�߰���5,<� v��{�~�+��,d�X_+, &3�/0�{A׌�PpZ���Ѿ�Ƌ�%	�^�v f���Y�>RN�o�<#݃�4����n���4�)���� }�A���
�.c��P������}K�q�~��ߟU��u c��l<:�Sv�0��dS���ޠ�Y�-i7QWb}4_����_uş)}�G���+��c�,��� �F�:t�P2�
�-y}qڱ�$��
+"+ꀆ �{��m��a<��kGTE��3�&/�::�w�,� �D�0r==u�و�����3��K� �xWk�'p;r#�~/x[�b���h�`i�z�m{�K�:����6��v��<juq���	I�T ;��V��묐#��c:�4}H���"Ա@$P�ȳ��^'k����\��^z���2\�E�]t<��[�U6N�G'�_��t��=ׇ��x�ܼ���2S��z2��V9Y?h�?^�t�?8�@3���.��D�"��#����Q��RiQG%���M� /D�#%�ԡ.�)t>]Iφ5 5�rt�<yIk5�L��n�C�jou���Q�r��7��^�kJ��8�M�+)r���q��O˶~�!�`��j�.����ųi��)�"�lݒ��$w\����,D�n�P4g��h����c	��8�~1��iX�����k�y t��)?��e����B�sZd�?5RiiU;����>��Y9������9�����E�$��I2�>���q��/�/4r�Xkr@՝̅^8���|bP�����=<=��óD�|��4�ں��	���d������j 
j�X��yc��E��Z��r�:�0Hp�u>^mqoN��#w8��b�{^�hTa��0X�-�X�|��B|Op����b���`H_|3�^2Ƶ���7�`Q$�|�/��ܽ@<V���^���2���3�<+Sz����_���Ơ*�$L��兰�5/<
����Y�LZ�ȥт��Z(S�h���sA ���w�L��K!��# g`��G�+S%�ͅ���,�I�o�&8#����: �Z���+���;T�aV�ڼ&�vVs�a�^3��Vz�X��LWOj�Nn'X�<�n����w�(��~;F�qnM���[�Yz>��ۜlF��0Y�v���#T�tn+0~��O���:���������D�7��<��
�B���qx�äc�vL���e�1:�jz"��u��g�~C�/%��c�U�\1q#p瀁���M�o�@݌�^h�׵�נ����i(�@̀��Cͼ��nG66��&��n(v�=��s�W�&(n����K���΋�f�k�����uc�y?�i+Et(�7����a�ΆS#$.����)�i�gk �G�Octb���U<��1@��~����Y�����{ʷ�>�8��}�� ��ڶ���E��E��'Z��=�~Ǖ���#������{�dʆ���ֿ��{t�+7�:B��;�yp�u��OO��*�׋>�2�����=-���k�J����k�B�(��?�E���H3��/���5�R:S"�c�CD>/���������zۊ��9�d��{�X�
L�sb� {�V�/g�ne���@c(^��/���Cv��#�kvj{ph�j�1I��fHDBkV�۞�͋��
�/A'�~@���V$d�]?e9����L�R���B�YX��l����ށ2~i���w{�hq���xv���/��"�W��1�u��9�Υ	��;9!ݵ̕Kg��������ӬP���{f`�TЄ��x���/V�M��:��tL
��C��ǳW�ݹ|u�D���X4���q�3G�Y�g�d�O�D�7Q�i�爩�t8��O��ᬡ��[)�wc�}���A�{�>����,���5w�HOl�?=����������9�E���:r��2��Jl���P��y� і?*����	"�����%�°��b �:�tuÅ0~%"07���@
�h�}"�� xK���\<�&��OCL�l��>��SHp.�1�5
��]5-�|<�F�7�d�xx�?��F����'AT��,��V��7�B7������bM��ٕ]>�=WU�`g������P�e�>�~�����C9mq�4˗����%E�3�mT{F_�(�؇t����Q�: 4Z��h]A\8�@@��)�H�K{޿�=�G6����*-f�]W�
�C�'[�3�A���٦��9��D���D�{��KYx^��)a�mk	��iV~�Ea���ɋ)b���X�@U6�9 ��  ��:<V+��߁��{��.Z��x�h1@x��co^\5�-"`ޣ�.)�
WN�z]ѥs�>���nԥS�>nd� �{�ުl���%y��h��\������h ZLC�(���{I֩��Y �ɬ��.C^��o1�<p����^r>�65��?��D�NLYټo�Od�S-�d}=W�ǣ���-m�^��r�sNBG�z5&����C���ۭ`,�/�M��x�癶6��b�� Ǟ���8�0���Z����4�;g��kP�aD�l#?m},�\=[�����hiE�2�+�WF���z�j9 )d���~���qU�k�4u$J���E��A�J(2ݦ�V{��i�v�`�$�^эՌ�(���e�A���KA�,Te��;���8�Pˣ�.����}^�J[`"�V�j�a@K�q+b��J:��SJ�
��=޺���cMK=X���K�!��GE=�C�DmJ�*QH��Hd��t/Q`:��D �G�5�I���3�q�<oбh{.� ׬Vx�a
�q�@�P�z�1�ҵ�$Kуŵ̞���ak�����C�#�u"� 24�*���lG�8�1먖믥�1��e���d��|jE)��T�I�Op��z /��d�����rͩv/ȅ�EW(Q+U�B�v\����tF�v���}���>�,����g�X\��s'+�1y � �_�y��*�Q���@��??���Ǘ'a0���v͑���`���`���JΖ��rv`�V���TB]C�)��ꌲ�a-F��!U�����\!�nđk,����0�y��y:�c�e�4B�q��T�9o�4M�d��)j��F�ǶʱM�x9[G��D\@��>��ǧg�������A��iz��3�{c����ΎDQ���V-n�+��dí�� d�wŪc�b�76�[�_���<�Nv��S�&hv=t�:Z=%5�`��3f ��5K���y�q7�̌�h�h�%<p��U"M4'~�Ȟ+xn�@���E�N���ε���`���E�����k2�Ɛ|]�Ѻ��3X�_�Q�1�0���6�?-���R��A�;L��pP�)]�� ���̙����-��O�A�D(�͊E�+�
�|.��Z��?��7?���b�����"��V%`�}+�1@��i;P�C�Q�l2�良��Wζ(( ���B, 8��F�E�|i1���)Gh�A�� vH���TP9���h�A���4&ґhE�3?m�ɸ�r�����4��ǴG��~/����!���`�f����L��X������>��~��f��v˩XV7�h[R�Ē�bYG���$�S�'���&z?D|Q��g��褵�Cm��(.��M"� ��"r�i
���������W�y��۬<w uk}w9��D��¦Q���"Z�����󒾛G.h� �؟����%o����H�BN&k{�.�/,kz�83J�$d�!�GyL�&J<E�'N��:�#������O!d�� J���R/�J���jH�`~��s���l@��ۗ��o��xG5^)0�kD�� סs����[�����tΒ�7��4"z�L����l����]2X��H���"=��h&�\;`�I�^Y�=?l�6�<ói��9�����jrG��hPC&{�c�}���;���m߯6DLCN���eU*�k�
[��w�f'�B�Z�I�dc�?A���V�?Q��̓��X���2'�� ����1�ɞh�?��)@��k��>Yo��h�C�<x����BW�6���O�a��Lr��-�a2!�%�����	M�^kS����7 *�i79���m���H����������d�g�M��;�a5yn�q��i|;�����χ�Rc�S����ڠ4G��������W���Wz8�ɳ�z1�E��=�0�,zeR$x��i�ٌ��:ZQ���ER���Q�3���)�2+� ��֌�����B��?�ﴍ�d�@�N�{����g��/��+���h�j�,�a�(�� ���U��Pr/�w�QbEW�� Tx�y�q4UN	'�+ziR�[����ȼ1���r�?��NOϜ��C����rh͋$N��s&���h�Eӵ�XS� E�4'�l�N+!�K��5e-,����y��m�G�`�C�A�	!�}~�a �iI�o�C�c�QEiy��WF`�$�}� x�T<#wt��
*�K��<������kLgO/�t~�D���F��;u3\�&Ez�h
�-�}��|q��aPgD���Ef�0 ն����	�rH)1%2�nB���=�2I�(�U�$`y���\��yѽ�� t������*�}���&c�A_L7�?y�qn-�;Ӥ(������u�C73����ǡ!���������hՎNL�M���Wبe��0����;���=v�n>���$��
&��T3_hN�K��`�(���Yn/�y�|\��T5�j(|��Uk26�c�
~(_��<�̣���.��_�0�䝏�נ`z:o��8%�/Dy��[)n�6f�ClW��˓$t`J�n�˷�y5��u�
x��e�r�6σ�t��dz6/'�w{s�� x9�\*}�́��W7�������&Wl�!Q]���L�7��L���<�(�T��=�%�iܥު�h~FΏw�⒮��~	s?��ze��,S���77�qBOj�����+1X� �Ģ8�*���D?~���u�翈#%�1��5;ϯw�ɲ)�M��R�>�A�	�t*B՟1R���];�/��d�B@�3Q��GP�Hp
�ޜ���d/�.r{���w���5�@;{��"�
@G����O$*|��?�^���G��D���.Am;�����ʳ��$����;�����ZD8����E 7�a���̺4�`O��Z8rL�\T�ӈ�b�>��V=�,�ً_��*��Z�QF�O���2�;P��#F�"s�m#Zh�C�����%�,>'�knغ^_]��G��䑶
����<XmQM�f^�Oy�JZ�l�(/���UW�i��#zK����9�_b/"�)0�	����8uz�����E	�w�MMd� 7S�=�Ӱo\n��`3���.Zp9R�T�r
!�4�Eb��y/�ʾb:�r�;��M$g}�N������`�8���i�xG�0PKǖ ���2�X�Y�� ��t0�~:�Ot���5���u��aD���Á�iB��v�@�f����s��ps�4g,0ʧb�J�.O�OЫ �~��H]�L�����,o�(#�.N�+LCg��{�[����lR;~t��"Mq�������=��Yi��Mҽ��ͤ�2�U�`6�s|Y�jv~K��G���@~�F|�FrGp�iUg�{_����܉�-t:�	�%�k�*��a�'�̡C>����<Ic��}����u�IM��M��h�"��s���K�1����kIVObȭ�i� � �f8ʏ�����0?0or>����~>�ޗ����勀; v8gs4`� 0,���O�o31$a/��e�\���pt}�����ZIQ{�̙���a��n�����0i��iп��;}g���
�1*H]Pb-F���9R-�@���UԔo�B�q��3}�蠥� ��c��(�ZF-<H5
j�2:y� ZH��[ c��
ӹW������0����E{Ɋ�V(��i��M���[�!��`Ъ�2�)M�`(e��U�;��>W�K�����Awʴ�����!$�߾�����$�y�b��#_/����^��<Z ���4�����%��e�.�xqR/��M����C��T�52��;5'V ����y.�/�I�0�S���ʳ�O����_��� y�f1�"���f�����QP�k�Z��r�DO	�?Z��0ņ���ү�%��R5�6ap/�4�Fr��9���<�>�������g5&CL�fNgF06�T�����T�AZ��Q��h�1m�9��ר���Z�_i�h.@��� ��@_Y�_oXS���-� �Q��ݾ�{��]�����+\���Rn���fg��I�q4}��&<o���0-J���Q�e�k�zd,���l<�9ezc#Q Y�v�ޚ(����5�0|�a}o'��u�h֝�z0f&�|ȭZ�Y���QD"�� �j~)��ށ�o���x�눒c��,�����_Q��XW<��n
G5��`%d&M��R��I~��W�E�皁����� ��/��,�/�Ic��U����������;&)Y�M/(9H�A��)|u����63p�<i�^*� ��W�1�������̏�;� '�)���
�{����`���F�� �����<�L#b����cd00L r;ީ ���=r��h'��?�p�G��8W=���|�M9?�����v���W�W?z�A���|I5k�����A�u?��7I�@�<��xUX�B�R�E�St&��<���2c�̪��T[/t���RT4��ysF5rY��;���)-
͊a:?O�#��tV����_�i��=����m0����k����r��:���q-`��KZSG��.��:X��>��� ��*��-?�ٚ���g#G�ʰ� �Я���`��d��i`c��S"�_Yc#�7�i�ծ�wQ'G�����z���~��q����fz?�zh-�������3m�ͺ�$ �����@�T�u>�;�ZԜ�wG� �lS�ns��@0��N�t��+�hN��Y&3�����0��,,[HŖQ~-)��C���k�`������71/6}X��y2��賶��XR	��s��I���������[��W��\cR��r�3@V���
,s��08�'Ys"d"0v@ � �NU�C�C{T[�!J~.�=�j>Yk�V�x歇*|�i^�?~��������������o��e����ۙ��̼�d�$-3C�أD�C%m��{�f�Q�:o�v�t��0?+gy���� �\D�T1��DC��w�D Xq�Z]Qr���a<��Ԫ7��t����+�G���a΂���At�2�n��Oi�G��^b���(a���xz+y�2�&JX��`�%N�|U�T5\<�2O�/�̰�r�K'Qf����g����=���2+���M@��:s����L��~w�Ra�Q!�I.��^���YP��v:��&F���`���O�C/�0�Ѣ(��mڭ��Nn��7��(��(ƀs�
�������
��0@��k3IF��0��gK
F@ף^p��Ϲ��k�X;��G�%�9,G��hn4��*�ų(�	MW��}pb��*�~ ��x��{�9]���E ��}��@���e�\L�7�Q�F+�P�����QbҎ� ���{�8�B���=�`H.,˗��3�}�������܃y�>VE[���z<�:X{S����1 �A[��=���AqDj'芺A�/���«b�K��%#�=TQ�G��!� {|�dJ� ad!�c(|����/�f�����I�!�'�~m�Ff����(�ՔQ�G3��*;B��9�
�RD�ɞ�t
��_���p���4��탼�C�5�Q�٪�P�h����(m6u��Pϯ�@�H�����#��Qg aղ���Š��|}8���A�s�g�WFTL�ⱔ�q@*K��K�ߓ�q�Ysr%�p�8fL�D�+���� ���4�'�c�8òzY��������$mn�Ϗt7D�qP�K<B�@'���`�;G��(�}G�ba�������E�_��xo销��$���3%Z+����歼��Y.�`0���@��.xL�\Gu�<�l+H�|�e`�?cz�1]pԊ����Hāb����gS�z����v<
��O���Y��Q���	�D�㧏�"s�;�F�ւ�e�ʕg12t������8˔���� K�톣Lt�׳��h�t?���b��J׊��m�-�yN�+S�h/-���R���hN���G7�l�s�5#ZO������|��ݍ�{<�I���%R4��p�
�#�O#$�L( @&I�>
��~�
���x?��IW	٭��m��AA���d��1RUDN��	��+��#�p��~F� �sD�����?]*@�i�?џ~��Yg�0��ٺ���H�im,P�8��W��!{�nG�_��J� B*���KMO�*V��xV�����5 =)gѠT|>5��O���,�k�Y��t@&M}��x�0}����F�
(��~��FXWD� ЃcN�v�=�%S�Qd�$run��\�Y�7г�`�H�{ZNQ;�5Y[�f�֮�eD,/yW`\2H����Ns
	�S gT������V����Q�=1_�9=�~�6~���� �V���?��o��?~�����L��6��atR��P�0�8 u$b":Ю��0�">���9jH�0?���	�C�^_dRxC0@�����p'�&���}99�\�p�z�� 5���X����㻄����+&T6�8�	Vڥs�<ٌ�&�="g¸��:��A}k�ï|IA���<�uT�� ߷)E�ʅs��"��a`��D��p�(� 
�<�_�~�����������'��5���IX�/�x��/ � �R=:��e�$7.��DcsV��S�?��-L��+�R�5��]!R	��9�j��@���^�ӅxF�v�<%����3ڸ��9�����+Op�^��%B! �^!���s��yS���_�tRpQ��j;�2�4��F]՟��2���*Y��ǥݬjr\?e��T�.�ş��ś�������~��H9<ITĝy0�G��;��Z�ĳ�m��t�cy�H���刲�y�h�퓅�?�r�2
�-�������sA��M$5 F�q҂Ԟr��/��v�M5r�17 ��C>�R �1�,���^@��i����\J�	6�*�C���f��s���*���pK�w,�5}��3�y6"��pb/���ރ���, \Y�v<�
W���9�=q��uC*L�~��y�xbo@a�_T�����镨n���҈��ݛ|enBY#�N���}?b�J��^E�Q����=��x���h��#"��[�7��!E�%]��r�����[��|�!�`��ю3�T�OF�������2*�p�He~ĺ�Aǖ������ɀ��(Mrgc�NЦAX'�%�4�i:�^���΢����p=�)�*�QRgY#:�I���8E� �U�툦v��{��:&��iZ\��7��mo���?�b@��)�4-�N���� w)hC��tբ� �k��)�[<�(sӔ*֕��2��f��ͧ�7-@�.�$ߋD�O��x����H�~�j)Y F�&���:�Zbou1��{�7;v�;�b0��E��\��Rz�����ynV�k�^�'!��u`�O������kǃ���l�|�mvX�3�t�f�	��˜�\���"%:{�7N�>Ƽk\�����ZM�Uv0Y����q}���9 ��&'�*�Xt��W(�]��P-u :���/_響�Sl@v~��\�����n�����+�����@\��4�ށ�U��/m\S 3�WMg�^Ŵ3�������� 0jeǘ���0�	B,@ Q�ޙ�r�gCI�Z�@�~_k�"C��q�Tް����'��c]��K��l�*sTo�5b��\l��# ��c�[SR���j�.Wݖ�R'�-p�_�i��(V�S�]>?�����S���`�
x��s�^)��ɝ(T�p���#O*�
�s������h@���f�??��h��|�F�����tŪ��R��o�C����<�:�;da)�A68�yr'svbcs�I1%�0-\Q�3B�y0&��s�!D^��"��HB\kR�h�83 N?�����ۿ�%�O_>�f���i~\���`�xð��Q�R�j�ΜOfOB�Y���)�
r���X��Lv�D,ߝ���u�*B�d��"��Y�|��pJ֟���s�������:J}��YaT!3^.�	Ĩ��V����� �tj(�-㳺4jn�n+�&�ɾo�Pz��M���F4%;m.�<�YQ~����s�W�S<� �2��VR�G�aC2N���޻?�r��1���5�FO�w��(��98�R�ɿ#EjY��v�8����0S�T��u�
�ݞ��ׯ�eރ���~V�pP	��k4�L$��/���<ވ�?�?��r����iy�C���|�xx��s��ۼ���s��,o��aVo�9�ny������� ��C�[�E���6���CP�(��袝�	J��Q@���"j�;1$eN�V	�ׄ�����֮�5%55o��T/��1��G���QODa�(�^,�b�sDx��u8YtCѨG�C(~��3p(0��@b�+�Z�<��A���i0;	���޺�a�d��S������ab_�����(�sd��h�c�����K:ũO�*	T�H[�a�| >B*@ަ��꣍Z2��;q�*S���5�ʿ3��+���q{YJ=��>(�V�t�s35����9�y�5� �Y]��!�1��i�zMgظ�z�>??z��@C��z԰1��~6(��<J�MW�n��l�F����	��m��K�/�⯖����fF�:4X�i��$y�u�6n�ghJ�����xP D����@<GɬH���ُ��^��3�q2�v#%�ف0Y�7�]�����W���*0 �F��|Q6�3kĘ�+���LۣE9��"_$���mr��_��tN�y��P�Wg�}���������Fd�.�Sv@_����hj ��f��A���+>EJ���h
�z�]�bN*�p�9��1j''��-�Rgf�7��Y�[L˄uV���AjsĠ���ZM#Yk�X�A�l)=�(�a�hx��z^Ⱥ���á���@�E�`}�S�u��Z���Z.�+�w�@�?��D���CAXuȰ��4���z�u��!i[:��Z�b�� �芄&�w���s�3��;ݽ�I���dO�S�A��������S0Ni4)5D�|�\����}y}��(t�mҢ��Ao�_�q�l��i���$9���_�a���&�2��NU�8�a)d�*��𠪒�=�sc<X8��ﵼ�JR����1�.:ܜ^�;���:9��8�dc	�*���ХJ�]QU�2�K��<��6�3�:��I�������%���zYB��zzm��g��'"~����\���OڛvIrI�f�Gfց�
�`����S����}l�`u��n뢢�fYr��̪�8��PS�Ns?B�{�I`�g4Z3�Ut�PX�N�8����Ŏ�6^��`t'k�����F��~g	&��~�C�ݏ�K�~�mz��9'�M~�$o!��ͧIU�L%Wr�����6M��a���x�h�KI���9�ߪ@��&�:;�f*����*�7˘�\]�0ߧ��қ�Ԏ��4��Y�CյIF��+p���la���sÈ�:�[Ƴ�n�S��԰og�v��;�NBu�4
i.u�� N5`d���a��	9�95��3�اϔ�.ꔪ0C��/l	M5��DL�����Y���$}�o�s\�瀝z-���R{��Vnlh����`�p9Gd�^�u��իe>����u�2�rR����Z�c��==�8t��\�ո������1�,���t�&c�\-ϕ����5���x�DN5Խi���)�:��w�g��N@�6�f{��il����π[9��f��*�{ճ؞˟H������~��lK�*�#Ǝ��Ce�u��2	�9����Vٟk�z��|�.L��C1Ř�����ŋ w̦u^�c����}[�6����/�v� 9��]#A�����S*]�4�6W��W�a�r�p|a�0��8�7v@ �)�C��k�F�j��iS�@NŒ)���g�?tN� /O����G�"h�'����1՝� ڹ5���S�M���>�����}?�>t���Gg�(�2�WJW�L����vJCٵX� �\*ƽ�sj��L�@�>����r�����Z�Q㡵���;2�lץ�g*'O3�G���phA�vYz ��#|��}�ϝ�Z�[�$�#5�O|����n��Iv*��y�Zzr�k)~�z��|��>Q�T'�)@���vl�t�᧮�d(2��5�nٕm����X?���E����z\����6F ?�A�ǒ���5:������sMJO�,�c�n�I2Hw ��o_;ؕ��Z��`^rv����i��:㎦Ss\��6{����[����x�9 &�}茕�P7��ˆ�W��v�8W�\.�>�l��ÁIi�Ddjm�1�پM�h���U�yk#����`�s����K�/����)��FL�܎G���~�G���6���1���	8M�+���6��lp�V�k�>�mc]�&�U�&0d�K���X6ػ�a�e���y^����e8L�4u�?Y�V����6��u���8��+�)�J�m�@����`G���>��n�h�:2]z�[�R�?J�ͮ���ǒὍ�����Q0E�����R�t�b���K��jCՙ��7j�q�
��k�I�UUn#GǸ\3�Oi�}N���bK��gu��֟q�aW�Zbf_�=VG��%j�"0��U�ӧ��ty{�>^}L�������˿��HĹ�ٹy��\+��k��ב����欒dND�8���(b�DK��:��B���  (���K(l������4��]]g��@�F��=��ि��e���J����O�o��F�g�:��y��.�x],ڹTUo,D�eϒ�0���P%���BG��$7�Q^��u,���������8�x\~��z�.��m]���i��~%"��缹 �<��Y�F'��� �=�BT�n��JP��w�;_��9^229�`doPb�k]��Q{�كc�p�?�OL��KJ��ԵJ�o>�-��]�����g_!Ǿ���#����z��a~������W9�-�Si�g=D��l����1t.�\X��O?�h +�8��*�G#�ף�o��9�kLk���������.PU���2��#K���9 ��7����)���Ӎ�
��2{fe?��}���@gs�"6#�i���jpSۍ�R��9kY&�
���}ks�B�bA\�� X�}�h�kȊl5�rԾ����)&�&�fJZ�Qէ+�&��l�I�h���.H�ϳj>ν�x����A�8�~a���>�X~#��,�f����,�ΰ�Z��>��ϼ_������Sf)X__�������?��Q �L��������d��Hoi3n�EN�5���7��A�(X9f���l�|Z�p�{�jϮ���/<|��:�906Yi���3G�M1��j8l��5?��I�9���A�%��~e����K�t^���@"���b��sw{k�>��Y�Fs"���ͲP���?Z�K3@���Q�I�+�}{?�Bg:ΖTϘ�$����Ȧ7��Ve=�F�G�����&�q���=0-�x#C�:ud���.�Z˿>�F������%c=~���kw2�m�\}�
G 1�5U evܙ�����=�w��Nq�Dio��}Ά²]�?���w��򱲣{���;���%�Kv|b�'�h����,g��5��� x������Y	-Xu2�9�#���݁$)���
^h�j�n�'	��y������8�k*��>�����/�����w˟��.�?D�G�E):?}}�@zr����t��n��ͩ	��S���ya6MA�gi6�\�ׄY�T�e��D[z�꒙Te��Z%e����=��#ќh�`K�\B�����;�u�Z��W߼fY�7���H�&�‱:�^��l�|�^��+��7�Ɠ�I�\Z���Y�I��iG���ɩ����N
�m�i��@x �c���E�ѡ�i��
�z�W 
g�}V�IW;���ju�d/؍��:cƵ��TFW}�~b'[�7Q;�	#_�ʟ�h�"�*%�d�$qѭF���s4��_�L���||2��[Ӎ~�_�8���[l�~Y;hݎ1x��������M�t}�>�,stw�n�oIA�r�j����]I���Ү,�)�����䢗(�J,���삅�����{rC�8@ֶ��w;�2�0V�~g�W�D�َ5�j��*��;���"�	_f���/�:V���_/����w���y�k�r	J5Q5�2���SSKۄ�g�w<xۼZ
`A��@n��ș���w�I�}��,�i��]t-©t�� ���{�dA,;��ϿJ/^�L� %@������[pR�5�2zkc	Q�6��!0f�]�=���̠̼0 q���5K�h��	ֲ�N�ϱ��J�Td��"�ŏ�B+�Ly�EۮT�!h�fu1���W@D�0����z�P,+ ) ��oL������顺�ōۦ {}�o��`�K�Ω��>�q�3/pG-��� �œ�����v0~��������@ڱȆ���t����rm�G�<� �1ţK���5A�[�~9���lA�e�=��i90�毮����hk�7�r�@�c� W�@*�,��$Shn���an�Ԛ�S���B��
&��GZ�u=A��p��fLs\Ñ� �c�Nf;ش�r3 b����\œ�Ҏ�4縆��Ԁ����++h �'�UO��\�D�������[���1�|���k��gk��uR~���<>eOV�i�ٗ��{��u�R�*������B�( �rpb$[�Ʉl_Yi�X8;k�i�v�9�2�Z<�?��Z��d�}�(�n�������bݶ��oa4u��69��x�a����	�e��5�2�fTf�lnw��um���OJ�ԟ��ų,����V�����=�f�L�~���S����Ծ��ZY�K$����g�	��z�g���� vb{J�9#�ׁ�/��N�j�ԉ+#/�{�}^�Cb�%�Q�x�v�d�3���-��I�]&bK����a,�P��Y&H|�[,+P)�u-����������ג�!�h$uN�c&do �n
|jmWPR��M=\dU밮��5�{'� e���0���c�'���<�����:<X�$��|���A@v��"�Y_�t��<�^|��Ϟ�^I���R��؅���|�
��Im�S�T�2��R�=���@D�u�1�P�ӧ��ȳ{�����?_�ίl���uάt��������&�{���җ��+*z?Wd�lN�b[�^˫�z:��a��Tϸ�$��v�Nv��݋��x��`j�e�M���|����� c}�q�ܶ�c˽��d�P��A�����w�5`�~���K<�,lKo'|����2�b^+��M(ʌ�^a��\��ߑk닌�`Њ��ѝ�!���ir&=� ��4�9C?4%5+ҽ��_��ޤ<z�u�#�T����|���n�46�����:�'�].�X��5�U��HI�^k��;^�ơ�����Ē�}%ͦ�LI1&*i4���XF��g>���>=�;��y}�M�w7� ع��2P�at�mj��XJ}n|�T�|�K�����"�>� ����'�Y:Dp[Â�7��α�F�%�Ԝ���4�gg�!�0��,�E�S)P^Gd��2*����qŗ�����Z��c��ރ�)���=���b6�s�"q��oonE�h}�} �Ϟ>5Pg��ϙ�Y�Ʊ�@����W��=�阅�I�7
o���j"�d�=�6��I^�i1vC�@%tGy8�rkn��i�m�L�S�)�J�3Y���u��и��!���Y:�����ňJ��DfܙͨHGH�Z��b�Дa�'�������(@]�=>��9��Q�]>o&������=��REM�@�g���8p��Y���y��=Y��Z��s��;�h��\�(E`\�'۬ݮ0D �\�L�2�̓��r���%��q�T�^%S��n��0��.2֍�D��8K_�xf�j�ǯ� ,:�97��\�U"�r`G�X�|w�Yt����/�8'*딃$g'�KVb�=��I����=k.������g������kh"ذ�u��䦰���t�R�N�*NQi�X�D>�T���y�v����e�΃��j���e�
�� ����d�N/,) *.��V���몳GP W&�����>�jpik�H?C��4n6A���p?�;\�N�S� ������/^|�`c`�P2v�)�ҜA��u����v����9����\w�X;�9�(�����kI��&Ce�uf��F S���P�����8��w�������=8SO��t SAP�����GX�������I��t\�N
�Yᯜ��Ja�&��,#�0y�hMK0QA_�iM�G��<zY5�Ucʲ�ɵ��ql�� ��a��ա�x���P����Y~��4[�5fb�@_��s�:k��9)^�;575��S,(��#V�Cwbn<H,�?I���j����h/8_���a� �X0�e4j�M�D1����)�ܳ�i��4{@Vm��gp�k/� "�g-��_b�1t`o@.`c6 �lp�_�4�K�}� )0����f}�#Vv;�OP�;^[uؼ鄿nJ����ɥ�ߦ�����u��b�Qحb׎`���bs� HW�;�p�ʹ8?���l�ӭLi�������ٰ8���
SöY;)����ϐ ��$%U �uWP�:��f�^�� n����(�j|Ź�h�X�]�y�#w�`��x���L����'E�g�ϵ�{�=M4P��6�T׶�XY�3�Ub��x����6�gb������ƭ�A���u�ĺ:}���%*��9����t�������]wfs��	�M([�J�'Ig�\�iR�:J`�}�⹑�>�;o7�NVx�bޖ`(I32�yn⌲�7�+�,~nF���XR&>Y�#����G#^�}����;�.�3�ޭV�fi��`��Lɩ�9�N�[�1̆a��a2d��VG���7����I��˓�5v͙!�NN�a��?���|/��;��U�
���j�0Kp�T�:��)�mt��t��$�@�΃�5,Q���ԝ��tH����O���'+���^ʫn͗�e�"�b�;$u�{1-;ox�5���9�n��T&GH�K�TAxpZr�'c��.7uD&�ѭ��73'��)l4V�z�ʲ�GA�IG�>Nvx�ѾCNԬT
���&�� #�?���� ��3;%����	  
����j�
�CNtm>~�d"i��P1��=i�)��>{�A�҈x�` �5j��ElP���á�.7��� �G `��-j����ⴽ\�f�dg��c��k���P��E%�)t���q�mG�:(<��+cFl`��҉�*@��!�R��m;WlLď��A���2�r�@��:=��m��p����i�2
|���9��v�Њ��U��H�$��<�����zXJYR�;}�0�Ss��w9����#2�F�B$��s�U���������v�K�8X�����mWk���s�u��ʰ��~�o����3ͅ�Q�����Y�R@AQ;f��jv����=����6���#`�m���^vN!�|��Q�� �븮��q�� 3]��.�F]_T�5ϵ��	��h^_�I�?�6ˀ����u�ꄥ}i�\�\��u�i|T�A'�f���a�����+.Swx[,�J���ޞ���I�)'�%B� �wc�a0��=� ��R�3�a��W��������,�oϒH+E�N��!ɾ������z�ǯ�35��\I�X�*vj�Y�؉�� cg���2���%N&R�Q��P�ϵ�-q�1M�6b�Z��Нh�QFnu�y}�_v
�n^aИ̺�-�*���.ꝕ���5%�D#��
��� �D��zP^�S^��Ȃ��e�^25Tpe�O�����c���?�~���Y5�m��d��(�1�\��>����^U��T3�t��:�-~MM���p���$n�f>�q�I숵�m��آ�5����gB�%���o�.���smo�-�삵�3:3�ae�/������T0�0U����z����渗�'���63Y�X[��#����X۽�a�>�<`t�E���d$%u�\튍e;���4��� A�n���Q�*G�y+�i�hA��	{�F[j5���9_|�'V����pK`'��/=���Uv�z/��n�@R���}�ڀ�K+y��K�/A�h��M��Η�uvnIW$F!l�a�>}�J�`���t[�l���]s�!=��P5p�i�p�����iN��}�K�9_r_�ff�s ��ݎ�N��7�BVs���K�*�����,K�,��f��)�rɺ�L��ot�S���{t�@�1"�{���o��Z�0 � �bY��^���7�>ʋK������{�vd��IM	� ĺ�K�-~-�P	Y	c]ߜ��ʶ�l&�5Վ�����k�N\x�<��@��=-��b��t1�+���}1t�6�i�/�/�a����`�����u\@N�o��?<� ��01��[�v;׵^�����`/]��T�Q%MJ�Lů����,w��c�9ޥ�%6���N������Թ��N��-k��po�;���Fپu�J�O]�\��j��|�xr5�j���*�hj<��y���ᐼ��3e41y����X D�~����o�������tuuI�-�#Q��j��0g���6�kJ �L����2j_[1 "ZHqQn�OB\�s/��qU�dA�T�%��� T�,��:,�e�����¸hzc�DƠ��3�d4��� #�l,�A��?i��ذ<0�&(��4���`m{���2�eL���<�	�sd�cd-�on���ｃ-;nJ
��r�9]^]��.@9�̄c�����+�[�%�?7oU]O1�@R��`'�M��f`�w�����������`4:"%6Wi�2(�I�{@�e�j�+2��Md'7��8k'��?{����� ����[�B�f�Xy�
TG���':�k�&�M( g�ŋ����`�\�c�T{wL�z%'���z8P�s-��ݕ.�bR2&�ҐT�-	v��.|��@�������`���Y;��y�)ɱ��E 	H�1�s�b~GwL@����Y:<�mܗ�@K����� �D����hJ�Rj�_s@/׏CRF�A/Ł��Bj��jW(�B����v+�;�p&m�:�o��2��#K�̙+b88��k���($�؜�A6 �p� ��K�}x�p�(��4 MYُ�_;Wu}������J��9񵍹�:��R�O�)���*	�8=�yh�n�;���g��4���qN�g��u�<F���Pw���4;���ʶ�%���o���~Ա��]M�A6���vpM��s�6�S4���,3l�k�����=�V͞L���X�o��Б𼮻~V��(��̃�kvԅ�G�7��Y��3wk��;+���8Ӯ��.[f0�%_O�ߒWK@��g���X�8�
#��f������O/Mk`�ƛn?7?���``�%�
u�NͬnX5Q�l>?�l?i��&����QϩY
E��¿��k��5��\k�)���.��;Q�
:���b�R��R��-1�v������e��4G�>���'/��lU�U��(ҭ�������=E�Ձ�ʰB�=f
�"12tV
��HI�M��/>�j��:6�+�v��E?WAz[�ʄ��J�6��������d@��4�G��r���w��vo0DI�:`U�6o�ހSq���mX�;5���+��R\�A7iy�g�w4`osm] 9�D��|�.tI�$�W��qv���>g��r��=��o�����X��*<��,����<�?X|�pk�5&c�[�]���a��Lm�W���hL�9��A{��8�V�����xD�-?�_+�F�0O�(� �r�jL�՟7�Vׂ9F�˿#i���W76�y]١d�� ����Z���W���d�f7��`d���kt]���������R7��?�$BR(ç|d(t�wq>�k�	-;::�vU[�g�c�:�V�d��@"l�Y+��C���۴��/�nzX��6}B�|s�nno��9��$�(q������(�~�&
��cGC[.7���d� ���>@�M���m�F.�݅�g��˗K���@�VQ-7 �׍{	
����d�5�Vep8 �����͵m@,06�� ����o���{v���0�}	t��3����*`���D�ܑ�Y��R1`�T�39u�a���1e\����2I:��rj&��Ƴ>�&����ի��A����:a��&D�\��y��k�U��}d�$��B�T<�����Զwι��4W����,Bh��!2�D�� WR���o������l��W�W��o�M:|*9�$�AW�7y�<9`�ZfE�)5;�NtJs鰊ѵ�o<`qy��ݰ_~x��<z��Ǧ�ԕ�T���\@w�V���e����C�9��e�w8�pr�ؑ@"�Ț9�W���H[�Z���	�Z��*��$E�,�I�����'2�>�TYc�1��3Omb-�I)����@�x�>��yEI��q&�����ޖ��cD����>�j�moPtT�U%�cλL+�ՔH5 ��@�L�3�Nz�<��]�)<I�U���z>�;��7�{���hܮ#�C`�~	g��Nk�l���&�oY��9�����嫗�6���؎pLܙƼ`.B0�a�sBO�ĵ�$%9����<3�\̕q#)7��U	 ׶����8Oa�� |�,���,?�a}\[h��qb�r]��k�C���ॗ��,^��lA��������M������)�O���ŏݳ9^FT|>��������J�<�}Oi�	 �3Ե�z�X[����ZN��/��P�D�҂	������oL�XɯlΪ��Y�!���g�읗G�����,�oPЗj��,j�PMN�W��:��0�k���<w?��&�C��vS+��3[��Р+ʜO�k���ד�������j�KI��ٚT��T��^6�
����Ϩ|2�*_,�Nsd	XxQ� ��Q��'k��@HkR��u�}�j	amnM�lo?h  �P$󜭺��'�VM��k髳�h?T��,6.x��PA��:֘����� oh�q~�78P��ɻ*�`o��/ U���&����zA�V�4Qޖ���[3�I	5%$�=����ƴk ��2Ϊ�<_�L�ݯ�{��W�)��.�9�qZ?}_�V�̪�5Q{,�s0�K���,��*�4�|��Y�D�栒Z�N��G���m6<��x�����c�'ƂJ��G �����{}�ce���} ;��,J�A08@^ņv�]�}t���&��l�*0d���V�q$�LÉ�9����.�[>"NN�\��A�=b���Y v�~�_���dʹ浪!fd�����_����6��y�^���u����}ւ9�X0=�MX�j�Lgi�����*C�k���������>=�cz���W���xo�W��;?�s�������R��G���ՠ[-"�S���p���@����!�,�$!;�
���7�����ű<><��>��oߦ�o~��{��u��n͐d������vQf`z#�V`Pv։��Sg'��ea#���.�=��%�5�Ń��J���j�(�#����jL ���=1v�h�%x}�"v̹��dLd����ɫ�h�&?���8?�|�"�C��o__�Alb�`��]D�"��<`^���4ç�կ�-�&��Z�Z0�*h	a���pk�e�������\3��\;�X�����/_X����3(K%0ƍ��_�3Y�hk=�[vALq����;��@	�	�&���$푹��d�����Eg�����rmvKr�k+�Ǟ���tW9�q���Yl��!����9�àu�a{X%�:�ɟ�3�1�ʴM~@P�	b�X��j h6���p��H$�o�i����7 �i�T�g}:[~��-�6�Y�E 
w�$�}j�Ҷq��V(�y ��3N���T��ܰ�R�۫�����\�uhZ.���g[� X�efI�����s��]���Y���P����_����b�މ�;&��cƲ)XupWQ69�%�Y��mg.*V��&�Sۓ�5e��8�ƪ6�I��<��CRv�C�)�f`!��)�}'�F˸���m 8�
����� #Iﾏ �fA��c���GW,�Cc{N_���^�X:\�'Ad���ē)K����u��6'v�ص��ù�Y�����,��5峷DO�rk�e�����҅i;-�|�����nƁ%{.8���w���5�Yq�ұ�`/�AGu_�R������6iX~���	
0N�3����#��� (?^Y��i^��X3�1�(SD�Kq�!EIt��g�29��ru�|s"�,PFg��\��bI(S,m��������'kYi*A�`
�T�2Ӧ����B�m��e8��I(G���X¹3jCX`\i3�y}�����L�VW��^�%Ř<�3(%�ѓ�s�/ݫ3a$%-�ʨU����ܞ��i��枒���R<G�5�bnD�Y��K��-��J�TB�{����:�L�Ey��?Y�76%4�.�d�e��;)������m�Z��5�Y�`4���a#7c��� `Gg`�ɖ؛%��uf�!G�m-ְ�b	v�,����
�W��l�.��٥2��+�����2)��)�G𩖖���;�n��e��qm�F\/S��~a�dR��Ǵ���f��ɂ�J�����fO��98�<��������F�_z+bI�̩
'�1p7:Wҁ��n��f)������+��lf��y }�)˼�$M-�޶P%Um������4b+�q׹�}D���:Ghݘ.+��ѯ��~��(����m�~�>F( C�|ϱ���s��Rן�ί)��,�`>�q�Kߝ�&.)IO��ʪ��Nr�ڂ��o��`��.�il×9�i�4��e�/�w���w��ð���1�1��#���7l.?���������V����h���gr�S�v�K�vC�f�b c0[���91B(�F��H�ɍ��6?D�����������޾���m����:Jl ����8U��3�A�K������޲Cy��@�SU��w]�B���rDB���@	Z:=������a�XǠ[˲4�R&0`��>�N��G�nOs�4YPys}k�tv~A����L
��0`�`@@.��C�BW�=��P߃խ�=�NA,�����V��.Y�� T��U`9�ά:>㉷��:kA"��gm���-؇TH��r
�T�@7NM,�\� H� ?V��PY�/g�Cɩޭ3����5`��P]�ilc�v.؉u�8����<�=x�a�4s[�So�j�WD��^�Ss(7Y��a���acG���B����<����/݈y�]B����}̬l�@8�ly �*}i�j��P�p&�<�Cd|%�&{Q����L�=���5�#��B;x��v�:���n���l�ƸK�E\���s4�|DP�ۆ^Ɋ�N�����R�e�:0��Q���JtG ��Ju��|T����u}usc�K���VwE��E���w��v�4�(���\�ʳ��ڛA%_~�BT\�c��~�� ��\D���X��X?Z�^�&J���ؕ	�&���|����Z1_ؐ��	�9}v���,΢D����� ��oN��Q�ա�������G0�5��g\�˄��3
�O.�D[�a�� �놰bܤT�4䀇S�>-�sX�g ��?�g���*�^o�^K1�}du�L5�{SG/^>�
�t5K�l���Bp������{-��� G_�0QJ�Ж(����!B{خ��h�v��Ӗl�5p���x���٪gϞ���q�{��>�}N~�Jl���䂜��b�`u���%�:���s�1��Go��~Yט~h^��^���Ň���CRI6&��i6R�>��J8���̻ud�����ǘ�����4�")�� �!ޫ1R`#��J'u�L�`�s8 _�T�1:;B���f��-@f��*�QI��u/x���=#����	Ȍ���GV��᫗bD�x�g�nY�wf?����m������D�c�P�C؅mQ�5�/b섦[���}�:�r�G��O���N[^.c�%Nj���V�����C�㉣�;��n�DZ�Y�q}^c��CR�����^�����;�踯8�U���^��C@�j=�3Xg�tKL;���KvL�'����Z�EY^գ����ɓ�v�i�A�^�1M`Х�j$�%��&�M�(�3-�B��u��.?x�}�;gZ���RL2�r U,c���l-맙I�8�ˬn�Y�c�V˟��kqY]	�669�V�����W����l���&�=2&�5/6p�cm�ݹ����*WQ  ��IDAT�i��^�P�a��j<�C$H���'=t8.��Pw����M���/�$�Z�b�"%���N�q�f;��xw�/.�{�mź�����&���@0Ag˂��9�sv��|�5"We�M9��#�,�n��&U�~�R��!*���ݳ|������a_�,�q�H��嗋�9u�G{����_Mo߽M��f�h�ڢ�L��pwϨU1#c���ܦO��]O�1[%�^_�u�Z�*�"g���AרJ!�� T:Y9�h�=T��z��l�v|w�;<$�+V:朹�ώ*�6.���ČK�,�Lkgr���Z�^�A�!��N��׍��f�,�/���O�˦�d&P�g��@��h�笙ơ���2F?|Lo޾�5�?�hB/��Ps�;Xk0��d1�	���r�p��Z��~?h[ Cx��g��C_��(m�lO�ͨ����G@�="��Z���ʁ�,.�[���S�O�Íh�]?�Ȟ�N�X3����B�ԅ*�oI4�ݕf�n"͝����e}�1Ilp!�p2Đ�=�[�&׀~����[ 5A��?�1�����l���q
s�ff	���S��92�-�CAGk�|�2��x�I�f̍��(	��=�K`��֜J���D��4�������7ߦw��pye���y�CF`a
0P�CAm�!��{�3sf�ڼt��h�5�6����:�'
Z �l�(������D-N�D'WG���~02����f:3��7�r���3'b:�[�;�����Hve�%�E;���H��D�ႝ��vˮ$8߰����?�>�����X0��ٰ`�4�mX���m��%W0�Y������j/�؏,�PEB�F�5U@���郾Ah�w�����
������c������ώ9:��0O|1��f B~H�����bſ�%�j���̛-Kl��eN��Ü��N�v5�bh�\O �/���X�C_�_��n��)�A�$�?٘�D�4N�����#2�[f�r�ЏB����~�.����F��]�����3/�;e��5���z���8g(�^�1	ǸDTbS���@�t4�X�Mz".�<M���Gz���%� l[2'v[?���R�_ �4�5#Ա�&lx�5H���|4�D���1�
���΁o���:���`P�B`����sv`ك �`(�һ�P��O��]�S�n�q����vr�c���`�h,qK�ᇟ�{/ϱ!�B0q��'�m�;{����� ����$�7|J[[��� �K�S�8�&��:��[�Ne]��? ey��#��t;���V��St�]◷oߧ7oޱ�����\��H_ƴ'����Mo��s -n�~fK��<�U�/$�4Ǧ�Asb�K��_��:�t��3�$�Ͻ�R��'�,�����Vv���5��S'9�F���^�2Qo��}������yc����~`�#.�B{kt_�jq��l��ʚ�>5{�����{׊�_B�e�d���:eŘ���P�1��!��߶.{JX̚�/�N�6�I	Ij�B��g���˫O�Xg?^g���lTd�َk��T���J�>J�Q�;������g�a��c�vUv�/�d��O9�c�� �
�$_�|вr��H���6�8�(5/��`�\,I,G���<�6(k&V> ��:.���{W_+�K2�I��㓀FD��Aő�o׀r�[�3�0���;�������M�N�b���(TP��8����A!M��j�7ˁ{<8+����k�� ߨL�-$м��u@��H*��&��eI������~d���AQ����Z��z7w��^e��i����l���`�g���E������/"�<��|�nf�T\�	ca#>f4�b�h]>�s��X#�G���3d'���̏?X`
���Ǐ��p��� c����N��, ����ȟ�<��T
�)�Y�]�0OV��O�rP�Kc��sg��Q�g��vv�	�a~Q'�U9�5�*���&�2�ฺ�quor`D�,��F)�=���`���H�f��T��W��s�s��%8�[\��
�l�,C�ܺe^�3�T�.'����nM��s��d���w�-�K��0>���0�T������e/���!�'	 � g� Ot�R�D�)�_$9�ş'�jvߑ��)�o��U�&a[�g)�˿o��B����cz��`��4zu�U`[�}|���ZL�Z8)ng]h��������i  V�6n��w�����>���x鏃��v�@0F�s� O����q��nDy= Ha�M�UL<0��Db뵁bʵc�4�"����~��H ����:89x��7��O?���}��W��(�)����h�_�>T`��i���O������k��-�N/����<KӢ����9��+�0�/W��g�m=�C�C m	���`L��,e��R��J�������~��f�5I"PN���=��ܔ���s���`�]&�����YS��ڵ����k��Y��P�+����!�x!3��v�bt�T��:yy�H�u�x�܋��>1��7��]�:׸ ��9�L����o_�zi,��v�{��~���TX�C6Rj�-��R���4kO�;���s�����.�ҾS)v$x�~�{W��y;�1��ݳ���4���<}�̴�.~��ɳ� ���)��{N �ou��dU�kg���d��T�1����ZoɁR��S��/#yҞk7��&�+أ�۟ޓ&�m7��K�-���I	�U�|�R�&&�z:���y,KCLT�z��5-8��ixB��M��]���S������B��K9|��lTF'���K�7�I����_:���������C��}��b���t��e�{��:'D����?�����e�]J����+��S Z_������x���|�Rv�P&(8O��U�b�D2B{�oϾ���E�EC$��j��%3I�ad�_`rr;/�{��Pܷc��R 7L���7�1ڛ��+��3�a��İ�w������˥�Se�e�ٙ�ē�������. >%0Kw��~����x�e��'	�oY�8�>-��GoL�>]^��
�Æ�G�x�~��B]/\;k�C���K*)�Jۉ-�HdQ������2�]0uh�,I�Wj LUO�^OcS��!�߰��cJ)ƽ�G��s��	P�S��_f"��,�prQ�Dg��J���,�����)�^��������=7��~w�sQ�S/�sx�R�2�]6�q��GG�;�)v���� �tq"�8$�X6eo|�z<���	83Y������ ˁx͖5v4@���k���-����I?}���>�(h��&��Hʔ�/�t8��w�1#P�c��ȩ�g+�#ό	�#*�l�������F2q��R���+�u�zHӑ�a/���Qb�>}��D�=�o-�� ����|�1Æ;R�Y��|��=�J|q�̭t2�Z��er|���5.�4r�/�>8�w�08���{�L���"6R=��'��-�<���x0{@/et_��� 7 ���j6_�>Q����G��{ԯ�zIa
gVm�� í��r+y[愢�t0ԝNדRk$�U����#��Y�3�t�;Ǳ
���]{ �ֆ�S݇,��a�а�D&I"睺&�Kt"Bk����C����́��?�x���[�[NW˾8�5l�l_;Es<0P�k~8z��v��J�.���]��,{��ǚѹ��w��tk�I��A>IB�f�v�	z������W�v�wV����+X��ѹ�ȳ5�h�\x/�ұ<����?R�,>�{����>�� c
?��<!3�A�ɩ��Okus�H�-i�X������u�x�[����8�p�|{w�N]�]\�:i������wލA�2��mVNNcr��Q�A�~�E��2GO�ɳ�<9���>�n�1��u���9j��Y��TT��L��s/�v��ɁT^Üe=Y�����G��kT�A%ɋ3�קO��7�����SӎZƕx[�g�&e� ��+4�Iu�%�{�9&m��2,U�q��.5��YO"�s�sS9�� i�<�gL</�j?���{�K
�.;�e
雨��ͳ�����X�/�RF�Ə[��מ��CƔ���`�X)ಾuvY��GڣvMM��֎@��,J��#�ϑ�)��-�W/_83���C�d�6PϨ���6[�k���7|o��=^����*�{��3���:3���1�q^�����g�ӓ��������{���f���w�ng��XY j�m�o2_�#P��=����)(U��N��:*d3���q���9�g�8C���O��(�ǼNH={��pJ���J��F`�"Ӗo0���-���s�5f>@_�KS�-X�+�5Jϝ��n��)������e�X�5�oI��0~����w��|݄�^�*S�5m-ؽA��2>�c�G*��h{y�	��!�=�o1\Ȱ�+}:6��~�@����΁����+���g��<�6��x��*-6������l�y��՝ ��8geAߩcTokx��F ��8�|FM"	4�������5
X��"ӳYqf�3gtV��4r{.�����wu���.�ߠ6�!v]x���f9��J�}�s��%�.׸�&C������[�>�k�Eb�Gt���:���Ͻ���~x�֮6�%��+��:�8��Ce
��B���!=��"��}_ԥ��V�7�\�7d% ����\�V����A�d� �`bխ�� W��o���Ey����������No<;��:��v1o���k�]��#������&ƥ��`�}��+��y9|zuȤ����$tؒ��&I�XŠ�T`�647	���<�v;�X�\��gg���؋�kN��Q��="y#�<~||(�ܥ$��\s�]�T��v=�8@fv�)��Ԯ�=����e��k3����ł���l��5AG8�g"+��j���>��Jxd7������M�́��uĲ`��1]_�����[˸�4j�ج�b�!��R�-�}[t,�:�.�:�^��9���vypoz�0��60�Ѕb<�N�d�Yvez���z;��F-趖�fYB�Z���+f����9��;�G�M�г�y4�l�N�����K��g��/��� �k�c	#� ����K@�&�y�6}���2o�;phن�۞�JW�91ϰh���Z��C�o��C�%�3��̛���uU4�΃It�R�x��jY�s�3(G� @"�=���M]_�����a���-'U"r2T���1��0�w+ӱZۇ�*�q����;�
�}�;���6�1b�{�@/Nד'g��W�L��x�ǑJ�q#<;�t��;�{�q6C)6w�0:8�.����J�ԃ}f������!�������b�6�tH�Vu�>T1oe,p��1�L���<�r ����t���ppW ��S�EP�������Ԣ�q!
c��?ǂV�x�*�9u m�^�j��@�ྦྷ>�����{��>����*����ua�o֣�ra����>}'E�l��w�7�Lƨ�l�@cDtߺg��h�b��n���t�	3:�g� 5�9o��ڮ� {���Y�2W�ĩ��>r֣����A�Z�&�U�>�F��GFR=���[qm"��%q��Ҟ,�6��ٳ��vc���gr�	�/N����,i����i�3Ւ�(����;}<�}r����99m�ܜW׮��Ҋ����h(������K����j��ŬZtc_Y�J@FP� K�*�,E�䁊٬irG������tԄ6ǖ��g�l��[P�3x���r�<{���7؊���ABG91�ـljS�:r��+s�2̑�����<�@
���н�Ei���(�%&���] 5��&�- �s�N����c����`�n9�.-�uk��;�Q���K���>~�����-�M�/dp2�m���,
H��Zk��!@�y����o�M _���]������A2�q��u��Q0�s�A&OwV�
;��p�9�o�7���ۀ���+K�6��,�*	�x��Aa��8Ƹ
�T� �L{2N�|��5���	�9X)m�*%b��e�<]�%�]�e2(*<G��{|�l�%e��oz��	�xמ���}��m��M;�5?د��a$���ڝ����ٺA�$���>���b�y�8X��t����+ oJ|?l�ŹVR<O�C1��c�qzȇT�ĺΫ����I]K�'H���Y��j�I�U�uF>��8��#��k�]�E v6���������~�����N?��C���W�?c��]-%�zޟ���J������	#�G� ����ZFgW�dN-��J�8��kN1���s�ܲ,��+�l!�1����[KnіB'r�����,�A�a/Q�=��" M�',�&g����Kj�����z�4A���,s�%-E��~��ߊc*Ct-Ey���A�I6@���M���� et����(�u�U��;뺯{����QC�R46�6gi���~�xiX]ף����/�����ɤMFiI��0��$��3���n�,+�V��H�؁���;x��p�fT�F����Jqg��2:�߽Ko޼���?��@�(��M�K�Q�L�3�c�x�8��|�u����bI���1��d��i�&D�팆�H`0k;�2{�͇�`���sn޿��~]�B���f�ׯ�^�Ə�R�h���*�9���yP���*�qF�;
McC��x����Ard~�'�ָN���^V�;��r�`�c�8Ⱥ����� ��K�tH��j0�-�Y�T�тPpin嬀��{)] |����8{vu<i��y�X���è hźSG|h1���6���ry��3D��u�n�f5��\���ńd5W�?oonaGX�����O�t����7���wFU��Ǝr��e]����	���s������`k�,�W���?���Ď,m��GLB\#��w˾���V۫�k�l��=�9�`A�]xq�p��@����������-���OLe�Fb�R����n�.�?g�)�3�)f�M-}�O�V�������w\C!% t��c^��w�>Fͯ�"���v0c����Сg�k�6���Jg��gw�FϬ��{w��8��0�51΂��+c��0�m�7�*|>�(����b$���l�1��k�Z�-���>�:���a�z:�
N�Z&���F��N���]_E�4�gR�)2�i�S�^�N�=uYf@��@6�(й�Ё�Ջ}z��"=��:����O���)l�[�X���t��W���;�G�`?$�^�S:UZ&ݣ}������j�yi����*b�%�L����&{�̦	\�U�(�H"���m-��{g5r����1(D	���Q_}�����;�ؤJގ�Nk���ۛ������v��qc����c�}{ˌ�;���3gG[�;�����./S������J|rm@�4\u�ۨ�E����|y��5M����'g�`�ހ��Y#��=6L���MùA���(yA���;�m,�MGѶҏ�2k�ѭ	Sr����1�(ҙ��3ź�Mb$�t��4`��$��8<HW�Z�7A�U陋j�f�3J4��y���GgM�KcR��L{������ٽ1<����K����1�������A��YO�-K��~�	���+_~� Q~$C���v�!����d�,\��K��YM"U�.�T>���,7�}�x��SB��R������|�k}���5p��r ���&�������?���b�w����Yy���C���$�lxx�M_�@͔���;3!i�S��b��<�Zҽ�փq�M	zp�/ؽLk̮��~��77�dmo_�9��1����՗�K������,�'�_��	X�L�s�ۈ�t6!��?�����?�1��H��C�X| ؾ�H����T\�U ���?��`A�$֓�d_m�����3vMy��W�D��8�~a��ٻK���kc4>{�d�\���߱�I?�o|'�& &��0Ɍ��S=|/������T*ı�[��>G�%`�����(	ml���E� O�n�����	A� �ؑ�/�v�=(�+���p���Qc6is��y��z�d�l�=���� X���̬,��~��3��FKM>��J�)�i�ff���Nn�(�u���}Z�R`]R����CmG�ҹ�D��n�Un#Z��8���Z��93�@Q�� �ҹ��	����k��.?ЕK�A���� 2�=���3��8`�[$Q"���X���	�!�<0���vb�����HLO�P4T�j���|B�(��8F���9 *�����]�_.N�WF�C �@�����W�#������'Z��S���G h��2j@$�zl,��W�vX���Ý1����C]?� ���*��b�ԯ���,@��W^+���ASJ�R��xڜ�(�	�x�P	`.1C� �+o��C�Y��$斵q�Nax���6i�P|��9.��%~�[E���  �7�m|t� ܼ|���q��)h`�R�iKU�g�#,�4l�£_���!ٟo��io]�,���!���gKp�Yё�l͍�.��T���"�1[�n6l�H6bE�(�0�H�����C��z���Cil�;=Y��j��c9�D�$x����=�|#��,�;z,��-ȫz))t����?��<]e���m՛�L�:oQ�����m��%��L��K�b�=���k;�t��a��֒���|�1J�����\;D	�~d�/�(Ig%ڎή�ұ닉sg���;IC��?-�E6JU��$}�Ԍ+Z����l�smb^�>R-�e�Hk!�xC�AG�h�	u=U�2c�ԝg������?���H�\\���k����n�\c[�5�Kf��ی3����r� 祉3;�2zJ���>J����K1�,��:`�^��㹵u''� N��I��(:��b;bg�NXP�L+�����`K`�����d�J�;�`&�]-jA*	k� g����s���kj���ͺ"�8�bO�����K��ҹTf�� ���<�^�)PA�&�����_2�w��'�������nc��^��E�D�,���ߡ/���p���� zo����D G�,��1�L�B������ܨK�l$6q��Wɷ֛�7�����l�t�r3Г͂�� %r`�r$P�=��u�Jӡ���	CG�������fZ�/_ڵ	�Ś�lj�F������/1�1�А,�{�i����'sn��1�t-�`g�m� �6I����)��,��1ְ�ydbyɘ�xn��j�i����f�&J �!��[�?���u4	��۬�!�{?�y}��Cz����`��R�.�t���s�Ͼx���6h8xr׌�6�])l�o>��Jj@�l�����O���8��/�Y�eW>z4��:x��|l���wf,�dp��~8�Y� ��w��i�(��9�Z�:dx-��W?��S���~4�K�$����˞v:5�i��ʏ��q�`�"���e���1ns��<�79Ј1Vy�!���ޒh��ɓ����Q�������v߿w�s{<���I�l���䇝9��ͦ���p,XN�{|G`�+.z�~�%ד9���l�^����óT�/�
.�A@M�n�Yv��e\���d;Ԙ"|a����RPjV۫<�s�6�H���;(����Ʈύ�?yxoMHIR&p� ^C���%n�*&MJ1}Jd��%J�ن�/؊���6=y���..��C�d�ΪH�;#m��:	)%�,�]dk���RAI�K�D��>1U{P�-�H�Ё�	ʧ�B V����-��w5����)��ɠ	Q0��,�:���I_�I�+d�^ާ���_C�#'m������^,��$}���Ȑ�#D������1{f}���ӆ9�9��IY]k��W�'� �����D��[7d���%�J�0g�D��8����wv�ܐZ�
���{�7��5uX5��U������X��&T�`��q�vʠl|R�;MX� �QӬl�j�M�*��6Pi֩f��r8y�����%��aL��_~�%���K���;(����W��7ޅ�������g�a��+:Dp
��$��£8<0�`�@��K���N�W�_0�+�FJ�
~�O��3��{F��2��4�R�E׺P�(�������P�$����ˮ{2zU�S�5U�	 ����㍗5iNRzf��Il�z_�� $��b�of�jw:85pb�V��`2jf+����F���s������g�/L��u��_�U�:o��ꢤԘ��\ ZU����!S�E�o�#vsW��d[=��p�`����r���Ӏj�\B6��K��XS��`�f� cG�|��rf�߃��0TKz܁�(P�����:j� H����]�NT��1��e����[�f��ƫ����H㬄�G�ͽ/�3U�������l/��J ��&Dg�h�N�)�l;첂8�f)!��wZ�䱋U?�ץb��}��>9T*o�t�>�S�3��֙+�����R�M16��z��}���|�o�ym��_��_��_���%�,�3�w�v�f^�в��(5�^�������~��(���O�Ie�6S��ap����2XK�u1�:�O���#����N��`�Pz�v&�	��@0 ����y�
d�X&v���������M��/������E�Ei��mL�h̠`LK�h�Yrq��۳�	H�~�ڪ+P� u+_8��τ����y�(���3c�Z�2h�-�$ L�Syk�9�ܘ��g���x�^��������Ջ������*m�LmH0�\��g���G��>??�w��=�}�g$���$%6,����g3�ə�[��.]�V����p�x���C��������Rv=]�-ש͉d�u���9/�r?6���ֹ6ͼC�to���IB,��%�7����=�;o�M��[ja���C�+pG�#u՚QW�3z7]��+�`�x�fxM�I�M�� ��&!$���z���L#ppc�����_z���s��(M������ ;&GJ|��������~P�ɓs~V�ErO�J�۾X.eX��0��'G^��x�^��:=_�,�(c7EB��/d��"`Թ�����FXW_��\���dw�yȫ_L�	�f��$ػ��m�aݍ�H��:ڛɸ�=z0���c)�}$]�����w�={X�K7t�.ZX=��J���e��ؽ1&�T]�^�Xx{�)RM��H�T+FuS�MÎl���ŵS���#ۙI��:Y��@ ��rMvm]� �#]��_�9��hХ�������r���\Vq?'��#3�-@���h��&��*F��t�o5�KT���8x�:��҂D�m��(�T�Z=kF!���>5P�,2uh$��<���Up1�`�$����p0G��a�!���_�j�Z�ZF��2����z��c�#5�W���Z}����$�=�H���L���E� ��̣��=�6� �Bu����2�qo�`���t8|~����$�0�O?�����[3���mz���k�|���	������s���
T*4�Z�t�xp%Tl�b���]_��p�"�z���xFA:�,i�;�&LN��;j�A__�ݎ���kZ��9N:��z��hB��1�5��A�:[|)�<dg!
��}��ʪ��5�p��U�kNL��=�J����0��ܙ�/��Ǐ��/�� f� P�qq؂���w�1%
�%X��,��nޮ޺w��3��}rL��w�Y� *�5���/�f��}��-�tg��9J.Ě���Lf��E�#�LAKb��a���1����D���2N� ��*�C)lT\d� {�H���<l٥�Qd�����@���\[��Ѣ�A'�P��|�8�!�'��k�Y�O8Jw���� �h�|�	� �X;�,����Z*���#�r'썷�#�rP<gB�;
L��0�W����{)��СIU�X���^m�%j�@�s��;��V������H�v�+{�s�} !c��[�Y�dҞ� ����.X�,j���\:uMBΌ���6+g��-���;/����tv������kD�%�������&�2�a0Nޟ}0�N �X,�8��%��)i�A8|k�+��]bT�g�'�B�{6/�٪���sR���TAr�p��v9�Ƽ�& ���&�yk%�`���`��׿����o��19�7F:� ^ŸS�O���)�.CG�_�=�Z0!��P��[�����~K���$JJF�=�1��i��H \L6삟�
@��`Oˤ�W�!�6��u�尫��5�oᶆ>ز&��쎉�)����3��#��14U��y#c�LU�	�q+_�����<W��ÁBĘcב��)�+%`,��w��b1Y��	�c5W�_�k��=�� Gh[t��Gp��)��G�d�w�4����w���Vq_�S��e+YŽ���"4��N{��H��v�����7����@�q�"�0��e�t��)�D��ߪs�e�7�g�]+@�vK_���A�lw��an鿳l����Vg/��3�F4\Y>��bt �u��!*fgP`Z���!�/��ծCw����l��{ŹZu���?U��������\��m��W8�F �Y9�s\�_��`�۟_��������n����'�����K����ww7��2mǡvJS繚���,�E��v�`��Z��;b&j��ѝyp�y�u?�� ga���S0��DF�\7�P�����T�&W�%��A��] =���mɮKF)%��f/}��Z����x?��T�1�n����m��b�,�܈o"��!��dS����z�^��b(���WnD����D��{T�������s� ����vI���G�k��~���(%U��K�`���D'�݊{�8�&7����8���>_ub=�� �ĕƟ��7��L:����RJ�����	U�)nk�¶�Y~�u�ϯ^�d��'O)��?�(�S�������*�H2����e�Ptӹ��2���e��/��?��?�
�m:��>1c� �:!�y}H��eQ�l�ʿ�z�X��o�Z�F8��9r����h8� �����*�yK��e���zwdco�n��r�&��lDPo�[��A��ݛec]�_��������W��㿧�����o���2F �pE�\��r�̠4st?A�Lq'�4�->k�U�>�h\�Sk����J���u_��)���1��2�<F��3�hbf�*�ЂblC����"��6�m�!��ü�����Qy��q�t��_�b"�@�!��<��b�M֫��ȝ!���f-2N��|̒��:zj�l��ZM�������ݲ���9_�В�E��Ɯ��`��7اطJ���@Yݭ�N�<�y45|IX�@��0ųo-���#�9�����X����th�Q���NA��,<8�ECkH{����<:�g�E8Z66��4&*qr֘ڛv�E%FFЪ=�J��z\C���H�m�@UYZ����@�ur��%l��R�4y�@6:��[�&܆�U`�3st���28�`(�$t�7��\�!�Z2���c怉�;����I_�Z0��)��+K�` D+Q2�Uw�l���6��͎�f���C͂�c��+�q�Ϥ�c���q��G�ܲ��(K������:�%����,3��5�!4ö`�,��4i�̱�1OF�6���Ȕ��]�wal�R�/�w�Nd^��2�&��;�QF�dB���(G�p��6F�b�P."�nL�_1�2�zs2#�����w��ӗ
�St�H~i�1`*V��cYk7y�Em�[��v�ݳ�
�o��iiWv���8�љ��0�6����������f3]��׿��J��P�Q��;XWE�!�F�_DW��]�#G6�:^��`s��ѽ��D���%�KP�ݱ&�cbTJ
I+��VHR�4 ����tz��m�n�6�u���L$;AN ��$��b�T���ޅ@1�Ŧ�Q���F��l�+�(���`��� nȒ��tƤ��2�����Y� �B�E��8�J�fF��Q� `w��bcm�n�nI���ֳ���"b	����|�s&me��ث8G���{��K$c�|6|N ��j&r�$�'��εB�)ş�����5 $��/��Z=Nϡ��}F�p���%ճ��k/�:�۾��J�[���/Ʉ�������{R$���H.���9kL+��8S�M,U_�˿I���5s6b<�sf% �е�`v�Ԃt$>F�ĵsn���x�����X< �������G׬C��]�e,a���V��=}h�ݽD���C/5�$1 �g��(�ƹ�E� �KW��*e^�b�At�Ο��O��?�d���aX�:�#���]�=8�#6e�c@����"&�.�a�F�@@�9 ��igv���	dJ�
`/ !0�����44j�т��v>0=y"���Ҩc,��(�k���&��t~5V��{v��z���GP�m-C%H�ٻ�h>\��v�;��x�X	kk��I��K��V��U�S�\����!���ܗ�s�w����Q�Ҥuh%"���z��	G$�;�{�}`�������ѓd�U��dm�Y{����{���Ha���~�W*ݠ�%�4!4�q�AFU�D��yiCnn�b8Yp���\�h^�d� �-����~�>a#H|��s{��Q�����Ū���0(�ά�]%�(�@P�~q0>|xo��n�N�݄��f�
^_���w:�6[:J�A����D�VY��kv5tP�q,�9�ùotH��-F�
|���}�T�@��9��� D��8_��e��X��^Z��������۟�O���6�w߽����wU�"X�Cg����+ ���IK�&�Ǘ��\����bC-�G��X����u&�Qv�ٲs����f��y��%s�0Ql�]k�r,�%?�Ч �@�@j[�(w�s#$����3 ��5��h�4��@V-G�S`�A.��]Q�i��??��X~`ۦ�C�WZU�I-[4::���xc&�eTlK�dq`P����sR��C~@��i�)�&Bh%��t��yp�R�%�']��s�Q,j�XMw3=%��#�y����:�/�98m��9 Bo>y&p<)��Ό������!�v�@���*s�%�p����\�(:<�H^�u�؂��@�|�,��iYM� �V&$4�R-�D泟�h��n,�T7e_d�̶�l�.W��*��?�����A�l1"�ɵ����:��=!�؆y����K��@�n�Q&d�{`�û��<*��f��c���GfY)��z�VC(�5-M��3M����΁�aC����Ͱ�v�dkN\X���@����l.��R;ߤ\;j	$10�gY�2�x~H����&�(���z�P���e��i�X����U����W��?Id	\N_~���e��r6o�Y���2��Ln��W�8'w�V�3����+01;�?���� �U��&��������]�z��M��h�8�۝��l(�w��/11��g]7^���1��͑\ɕ�%3�@��K7I���iͳ�M�_?`���=���܊����,����,~od�li�ޘ��UD�Ȉ{��?~N\G�Xc�AяY3.w����V�vm�N}�ʹ�}S /�7����#* \P �E`�m�&��Fݙc����;b7�n4vk,�>��+�oV��oWJ��Y|Ӳ~������>?_�tpq����*�?���@���݌TFB���d�Z��'���:m���:k��oS�8Y�&�f��!���	��,д�v�B�k���a��9�y�\]���kO���9�kc�����ES��U#)(k�^�����b�uX��}b�v�fS?�B��W�9��ste�?v^�d��D\7`� H����v��H��gs��3gtނ|s�x��,�\Ͼ/s��@s�#6 ��n4�@���6h������#d엽AU��:���=�:��9re�d}�d`;bj��xx����l�������n�)�����Z����+g��T2�^�i�Ҁ���t�4s���%i8B��� z���87$�S�bg��>���L��ö{��ԩ�l�l�T	H  >��`d�5���2#��	��ty��`m�����Hz��,����f��|tkx����&@�`�,��h0�qo/��	V&�l7� P#���U�c�=4�qHc�a�s7�'��L��;5
��M��7�u1�'���A����`�y�K�̂��/�94Z�f5�<�G+=2T&qIf�$�,���q��i�.���g�Q��%�1�ǀ[��/��]��(s�.΀�É�1��hN�u��]�1�0��g{7R��P��ѵ��� ��@�/���E>��9���Zw$	Ӣ�v� u�H����`��71x:}�A�6��b�8;�C�d(:k��>��*��<y�c$XX�8��V갆����T�"K'�	�*��B4#�ϓ�]/�
�Ea�� 1\��_vx�F]�p��24X����V�P���;8C�N7yP[Y`l�U��c����f�[�˗�4>z�}z������w��/>'�?D^b�;�8�m�"�l-İ�r')h��Qk�����4nSO���6�jy��uo.��a�/f4����TOώ�~��k\�0��낟B=Kx?<d����O�_ǂ$��Q$���q����m�$�F��pO��w�� 6w��ݜ��@��4h�}�A�p[�5�"^�!��̊E�]��8kPE1��dk{V�ժ� 2�\�B��r�~���-�M�y+ݜ�+�L�#$7���S-?�8���a��.�ҡk@��Eq0��F5ӕIv\��ȝ�T��p��31d��\`k}	�6�]��ϙ�x6ۭ�h�� R
�6u0±�1{��p�c���}��XTh��ѰFׄ��tq�� �И��{��A78�
&H�k��x��$�gK#q`y������:���6����N0b"!�/f�Pt��L��G�.z�%��֋�Z�r�dD{$��S�'$�7�2Z�4
���c:��Ͼ�kP�r�c\��(D�존���A}��c�J�O$������>,KS^ �0�@�e��+A&�f��P�XE��14�#�orx)֩q�r��)�, JLy�kΤ�qn� !��;���$'��֊&�(7(x3�B$�qd<vv�M=E��J�*IS"¡J���TI���G�n��tr� �`�T'�wd�RN�[ ��t�-�?��W�l����e2>���=G�T����H �v�1҅XE2�, �����__[��]W�K�O��(�5	b̕��7��(�Q�\J�ogp^ Z��2vϵ�*����j9Csc<1����9��/�R���N{��)������m�'����af��B^�_�4��o,.��_<��\�s��q���%�(`�|��C�`>����*��۵u��6ͣ��<�WQڒ5�sE�`:�:6�3��1s��~����tm��,[��^�x_ X������󺱖�8$0`����ާ��ҋ)g~���tv��*��-������J�� ��:���0�'��H���i֊��r3�������w���ȳc�F����|:��ve=��ki�d}����{m�V�l�+��,5G�2�����:{�È��e�X�t���3�<��p&Q?�q`,�^����k�}n��~�A�@?�Ҫ�W�V�����@Îc����F��$�ͣsz�/�
����.�K���[�"ƣ7���9�O�q\��w�-����fU��I�.�si�c~ >0wyu�޽KC��?=�>�5f��^��Ϣ����Ab�m�XGOz[7;>G� n�J8C����d���>' G`>�����^g8Z�6,��r\�~Q?�̾��M��(^�	F�����Ho�Ґ	6����u�)�S�ΐa����#��q?���V�Z>�F7Oڙ~�gg7rn-�uz��-�Ol�#.t�~Lμ~u���I���fPq`>�fI��^\�5����O�U�GS��������رv
Ñh��L}�n����a��.�a���5��b���a���@WQh�Xe��fn����d�i��:������>FcY�v�7D��<�cyf�p��.I�����K�;�IS�s ��� 2e��/��)��A��שp�s{: os|����5�v6���)ql3���@��ϟ�gO�R$V�������j�tx�=c��յ�L��&?Ĝ����C��HT��Җ}%�Y������W�,�	vC���!?G[S�X����xay�#�6��{��_]O��j?ݓw�ol��1�
����l���I�{�]r6M������sa9T�L��JlJw�uqC�ն�����	3)�k�72�V@����[��VP��>ˠ����=��cd��g��!2����Wf�gs���	(�E"��0LfR��q��`���h�����:��v��4����=� G�].GiL�}��`�A\��n%mԡ}T��+C�p �Fޞ��h7@+ �80qok*�A�E�	�}�ʫ�"��fq'���,6��ͺe�^���w����lm_�8  � @��&���������ŨܢPT;2�~|���}�c��a������$:|?���t �&�®a׎g:�:�z���W���\�fcbXW�|ѩ��!�+`L�Ҏ>�E��b�Z�J����2�}C'�]>�Pn-DN9�����p� �:J�	@�	��3jA� �z1x$*+���b����0A[��.%�{�{��F�� IN�n���#�'����_,M���C9��y�q���)'�<�.�i��kM.�����#*.r������1�:���*nR%��|�F�9LIFF23#>����G.����^�s�P�e3�`�+��
e����:{>�"*��:�a)���5$'���
�~����'��&Y�WvPX��ΚS٦�l��H�g��£�k�
5m?S��r%۱�6쎝W��`͑��aZ�r�`K�@-��0���Ӕ�.y���º#�Y+��6F|��I������9Z.͘͋:�wu|����'?8ƴ�cxlɕt��`���p����kW��56jT�W��<v�:b�y�^5`�"ojQ��q8���h�����y_8�1��Mf��M �|�ԥp����:c�x���o0~"O&c�GP0>Ao�`�IR"�!@L���f�JCgm�ˣ#_t�=p�b-{p
�lD��Ȍ瘲Y�q��ԉ?L��&G����b(���x=�)��	̰ͧ18�v���1�ȿ�wr�1�wocٜR���L�ShJ�� ��6�,��<��5�їv�Ȃ�Q��޶���9�vf�^s�p�q���`�����eP'��⺀6N�Z.����l/�n�
w3a^��Yq�}��#$>w������D���x��ē�4z��1ž��ќ�>h�5��|?�(&�:��6f ��p��:�֗=�:t��0��<�k��Ë��h���[M����t�S�k����R{�y_\�3�mBd_ڝ�����`�Ok`=r$�����CC7��K�� oԝY~��L�Ŝ�_ lp���k�v�&��r�{���7b���ŶS^#ʋ�+ƙ.�03V��6k��T�]jx-��q���{�-�(�]S6>�̼��w��U��`6�R�JF�]�/D�`!s���<�߀q�M������J���9}������v�)t--,%�Ҥ���yNV���9��:v���>�!�I�Y@�{�#R$��n߾cz���WX��!'����uT��3E���9�:Ϟ<����w$Z{;�l݉8�W��B$l�$9��5�@����LU�d:���h�(u7�&P<*bOE�C"���E��r;k���%���:Z�3ZK���xr��8F��V?�}�j*�_��D����O�o?��� ����3ޓ�)�RDn����'�q�Y��Կ���gGqH0��+�-L�k����R�u����Bj���O����`E-��E��-�����PU>�mM��ݴ��~����O�Q)w��P$㠽x_�M3� ��}�,�/i?��C M���,~2ؔC�v�Q܄X0�-<���k%��{��wR�[IN:w�
ԙ�`���ws�������Ƴg?�Ǐ��*}EvZg��%]2N��Ab�è$����&��)6k�D��܂p�He����M�����Xhq�*te���X�r���{�N~���U�z��bA��`���y�6/��*��M�i帖��ŋ�D~)��3Ι]�R���q��4N��硔�f�`���h�n�F��/Ա/�(���eqI��G��>�g�f*�a6dq�#���5���Y�)�NM�~Q@�������M��آϫ��H +}/&�Twx�j�-A��p��İ��k���G&Sx���*:�к��`(����`�"x9f����(���3-�1�:St0����(zr�Y��h�^�g[%�Q���U�y
1� �B$�e�{Q�_�77krS׳D'e��HY�gqs���,wv%�OuR��ǚ$����m(����8�~���+��e�Ry~y��T�(l���o�qϘ�@TѸn0��J����C�� ����1/�a uț�7��x�}T[�ut�ڛ�q�>�}{�"��Eb�ڎ��V�A`^z�1h.�!��
�N- t�6�Voy��7���<Vb�����H�gO�# ���ߧ,v���	�.z��y	�����(�ou�q�cQ��i��;7���d<x�R?�>���O��dT�^��b��<�_q���E���k�c*L� �c��l�<�R�~���.�D���|47��6�%��z���Z��nJ.#i��F&S��z�5��,*�� �'�бћrΧ5�.?ާu-��:4ʏpnc���Η���l���P�b�F��_�Yj���ű��ˀm��Н�y� ыN�a���/��n��J������S�&�v�Zk������>��Z��K���2���{�(F\8�VWy��=����`��Ï�_$�.���#�b�(�>Bᾲ�Π._[ͦ �hb;��u��c�m�c'P���'t �n�Zc�Q��I����9A���n���4�s3��3t==��O��A�Cb\�>Ľ[$��)&��D6t�:��k���[�4ۼ^�Y�ٍ�q,.H}��m�)j7�bd7��~��@x5��d�`�uudw�P�Azԥ�e�^��n#�Oe�.�&�F�|�IO�p�p�Q����Ɖ�|2��_�Ѷ�:)�W�>�%�0��(4�&+�g6
�h7us��`�"����cS+M�����>���`�S:�&��@��.6
ym7It4��O�v��H7������_Uyޙ��%��7VLz*7Yr�f��v�ԉ ����W�\X>dBU9��3�a[�|�E�da6%�?�sw*"�ݥ�����p!
�/�ʿO�?�<N|("q(��	�.�9��ЮQ4yN�
1��"���Lk�Hc�k��mZ���1S�o��iF�����H�bt͹IGu�y��r�4Uˢ&�19�Ү�z�pmV�{P0�x��R��Q�� )C �yv��6W�̡px�V�# hpx��M�k�(l�������ߥ[�o�g7���n��[7Q�]M��Mf0!N�ņu���g�βv"����W	e=�k��1\K�yW�`�(~{��#6J��_�<���fh�.�XS.�9�)��,�X��D81)\v������0��{3�'�'V�W����t���=Fv!�5�M��Yٞ�n�=��4�2HTQ�Q�Q�kw��4D��A=�� .��[�n���[�PuSl���_��'�^�Õb�S�w{�]2��@�"rRvX�8
5 �ҩ�=V��uG�;`R���\Գ�},�t#�V��5�D�63G�ܓ�{ral�:ӡ�+n��Q`+N�h�u!��/�~mb��D��~-��R�fkw֡J���⯮�T�*�0���]��kdM�W����^� /Fk���0%��$��ٔx^���R�����>N<brjm'j[��h�T�ץ3�q�2UvJ~��O{�c�L���`6�C��d
�E�]+�f��K��ґ-�"��%2�}�G�S̉�XkӁ�E�!-	%u�fC4�s��Y���qE�{��ľ�3�ė./�hm�����y�(a^�g���x�qGb�6zE%1qԏ3���ތ���j�`��]��B�gJ��C�g�*�[5�\ N
��� �>���Կ�G��9$Q� k��Wү*#�q�l.����`� ^ߞ� 
�#���c1@)��{��`��V�[9�\Z��c)�a��Y(8���K��}�
�t���Ֆ�8�_�:罻��������C:6�jX@��}6g��G7�u?��cY�(�.��d�r���J'1��~� �f��h45g�nOg���Q��/�&��������+k/���:"��+%���9Qh�pN�j�r:Ö;�s���`a�q�\ �x0F&��<?k_&u�	P����R+9a�Kp��F����v�5�3^��ˬ�9^K��5p�:�!y���iX���N?�+��ņ-6.w1U�ɿ�t�}&:��ȥ~����J�����~-���b<׮��!Y�]f�t}iN ��8�����Gn�`�h�JeMCT�F 8�G�8Vf�[���a
=�k:��Q7*��8����Q)��=�)͢��kǂY�35��������56��^/r�����LA��jWܧlhN?v���2��`��wb]9֙�2��Y�
y�A�8����1�ufV1W����Exy����AM� E�5ˑl�r1L�1����un�5f�c� S�9\���W?3��.=�1�3������(�0x���F<��Al>�$W���&~�.��w�?��qIwD��?��$=�����<�u��f��y�{U��Q�q$�D�V`ǅ���@���Z��jw-���.3��|�]zt��Mg�r�3��U�#V%OH� ]Cn���ٕR<?�X�QW�gF�s/���\~b��X&R�6~9Q����/:��r�eE��/�����ş5��p�#pC"L�o�pG�� ��9���P_qa�^�yϟ��8������~���8�iC��|c�.�(xsn��m&J���	Y����{'�Mf3ER Ll����j�ö��פu#����!�יn?���|��^���=n]ȱ�8�.}"0��@�7�Z"�8P������r`:�:�O�#1���,(�8$qm/��J��o�����/�gӿ{�(����t|�v*6���G#�}X��$t܌UZyq�ʵ=��#�9��9RR����7 \/�=+��<�*���Ųq>�{��JQd�06M5u��tjͬ�Nx�!R���� ����Ĳ�-�7D��e!�;���d����ϸ�ޅot��s�Ik"�:��W���-X\tx�s\���J!��H`*�8]TAA��0�%��cOW~)k7������ã�қ)!ȃ�F�ϧ{�sb ��%$�����c��-f�%@���T�weaJ4}8�����s}��0���n�|F���O�>#;��T ����翱Ed��@��2#��Cc�rw}��3s6�-��I���y/��_v7�#:�UO�z:���Wb��u�S0t���=�u�c����e�Wa��E
�B)X�xI�`3�ܟ�iW,\'g�������H>'J��vg:���K��=��Y��]m���M"UJ>�XO��;k� ږ������67y����ľ ��B�e/�� &��;2�v��xӶ�9���ta�|��ƨ�q��&^"�{u�6�9���O�{Lcl��6d֍���h�Z�H@��� �(�����$GԨ�w�R���p�f I��Ç	��`�_�PB��.��aWx.p�A�����w�S�*��u~9q�'|YT�h\����l�a���yiW�`��-���3s3�u ��1��i��}�5W��ةpMޯr&�s�~���,몼'�.�Ӧ��y��P0�(�>
��HP00�;��t|��p�!8���͍�S�ǿ#���g��o�Y, Q?!o�x����6hy��N$�#�o}�I�v^iGw���Sε��:1�^4.P��|��� ;c�p&���3
`�G�0��`Ű�`�VFR��rA1^B�[�.��ii٬V��Cu͕�Ͻ�6qWj��(ZBPX��{A~��	���7v�E�cM�`!��&�؎mn�%\Ϡwvd&�GZrCm@P,�a,�	:+�|f�\ c�BG璎���h����-C�
�}g](k�xyBe6(�4��{�UM�A��F���g��8��)p�@]��蓏?Ḟ�I�z�׼5ˆ����y��9Kh=ew9i8��L�{M��3�;�K�q�h�$��f�����k��H�Y��G��:�k�y�l���7�hi����hfe.����q��9rJ�tRC�z�f-�,hvW��2�29��0�٢�i�p�<7�@v���kƛcف� ��[��@�Io<l�H�[�H��1��LG��޻/k��~�s&F�%��������V>�Ji�_1Ɲ��I�.�ե���}8upu'��.7�b����v'��6f8��
YLC7��ӹ� �j"� �����s�g�Et�w4�<g�.��o�L�,ɆD�]+�Lh��<���ʏ1�͕�ԯ��j�.�%/��^�3_�ʝ���Ҏ��`�L� ����'ڇk_4����/n6א)�� ����}]�m��s(����F�؋�EUsގc�2�HLCw�g�������_�?!�8
�Ic�b��Ev;�h�̩���?<����c[.����R����do �+@�������Gߧ��V�n
�rA�.�`&D�M��Kji�+m�4&o���5�C�H����5����Bs�O,l�>�L���n
��AA�̓��b�F�w-
ӱ�����k��j�J�A.	KI������Sb�Ш>w��G��������_������%�����'�p�GN�fG����/)���kk���Wu���2]P�ף��(P 
s3����cU�]p$)R�G��
$0^�eP ��äo̟�g�1����f�"ī$6 n�:
	`�42�Qq�0ᝂJ ��*���q`]^�.J��'B3���x��P��u����١]��Y.�J�d"ȟ�)��m�}	F�MҮO�n9�]����{E��\_���?�=�y�-�"����a���ǄFQ���`�*϶.\|�!��Ԋ�p@E��9��+lྮ�[���C]�H٭�x���
!�.��ܻ�@ ,���41-g��c ��E����l�C��ή�<�w��H�����g�{��c��e<n,F����6ul�:�����*1@����$��z�꾡#�^�,&��δ�bl�`�Օ���Y �Ne���� b�$��at�Q���^0Ȥ�a%��E���C��?�U�PLh#�QA��'��h����cm�q��HJ֭�9��}Hڟɀ��8]�E�t ��jW*���慢��/e70i��N���Yן�U��}�G���`_k+~Wk�
�x���'ͣ?��|��4s�k��ms� ˘a/߀��>��)sQ��3��Y\�@���J�ŗ�}=�)�)�'��͐E_�	6K��~�/96G��=Pg��6�;F"~,,r-�>Ո�U��1&�2����j�1TzW_�`���霵6_����mS�P#ܕ�ݙu��1�z*�G��I���#��ğ;�AF7C�8��G?�Y�q^pP��ba:�eñ�F��X�*�5����"��Xc����`�`�G���o���9�M3(�5''�|x&�i� F ���8�| �Z�A!�2JVp��K3)G�k�Ҵ̷�u���R{k�i<����C�C�L�ul�8�8=3[rM����c� ��L��.�u�S��Z�q8�p@�7�,�k�{k��C�ʉ����@h�
2
���W�>V%g��,�¶K+#N��3���Xkm8���qQg �Y�n{1���|M�zp��k�8�����#F͜~�7���?�1�[���Ŗ�`����3��ݹ�m�ꜿF�>��/!�Qh��Դ�5P���#��l:b���=��i�Q�(*�0-����P콗��X0�si���۔��]Lk�g��bF��P,Y�m��T��s�9ʚc��Eg6���:jcg`L���QV4y��Y������r��3���:�!ߐ���F)�؉&PrM���gǘ\���X;�\2K
��Zg{i�!n��U��a*Q�C�-���7�$���b� Wp�;B',M��T�O���buu.$|��j�j5�Ƣ���~�YBi��p��+y����"�%&���Ԥ��a��\�=v�L:PN[K�|o����0B��!'41�z6�D����ov�����:9��ƒ��5P�l�T���ZhW3�s�i,q���j�NS��0�J7=��b��� VU����e��L�Щ�O�!�Ӓ2=�����'�>�t*�>!Gw������ߜ�FM��uz��E����7�~�������;��V���)�G�#��(��H9q'F�R	1��Ik<a��F�
�>M��$
iX�#��댍���@�lJ�!
��/���P�z]3�m<J"1��T�
�R2"��qtk5%8�� ����Um\��v�t�X�v�����"������nY��4%A7�uA^���P��~X����my.>��Z�D��Ak�1f�F��B���y��:5��5
{N��hg��r~�ҿ��k�XR.��j�����3��
�4��mtp̰
�D<�'<K\���D���'�(�9�t~l�K�N9�q�u)��JZg����p������= ]t�Ot3֜�?�����ҫ�Y�K_~��\��}	���#5B"�[f![q���s��}�����������Q$&��Tz�-���mS�.����t��@
6L|O*��#��8�0t�P��$K����QL�^�8=Nw�b���O?>y����?����&��?�S���Y����zhp��iD���"�&�����!�"h��)�� ��e��Q�a��o.FbF;����*�T����^��rb�:5�	��Sr��@$�Lb�,�R�g�&J*@[j/il�m������\S�G~V�۴ls|��X�`W����gb��		�?����Mu�'�O�/P�� k���S�s�[ƨ %�#nO��s��u�| ��� ��!?��N�e���X�ŉ��e�PE�r)�b}r�}���ߐ�v�$�E��������!ȉ���v=���_��l�uk�t��x���B7*- ���x���t������Oҗ_Լ�M�3��m��ه �/�1���> {"\��J�6���\�G+���}_��Z���EG* ��A� ����7����H�}�D�8�Dwr��{va2��b��h�}��G,��t�I�����;�?��L�7o��d $�`�H�r�ʅW��{\qȮwy��LhV�s���)�>���w~�������9��v=��\�	��"��3ŕW��H	�w��	�V�9�k��r�<ԅ��Eq��t�פ��#��dB�%u���)C�X:ЙS�j0��>yBGQ������Sdw��?[��5�:8���m񻤿A-��)�KaOa�E3L3�X4Ų�Q5�/^Wt�2��_7R#�E�%�ю�cz/^>'�͙z�ò���@�y y�Λ��YxW4�s��\�&����h�3P���?�_�=�8����(F��V�5��C���w23G}��jO����� ���Œ�H�����3%� ��[�Q���D�:2�j��7�} ����ӭ)F�}~����V��t�S r��ށ�5��޿{k7!���0�:��A��kRR=���C��<9б�=��m&BJ,�TpW��Dl�&|n��Ƶ����D�Cf(���E�Q�T���� �õS.p[�{��:tUkU���Z�s��Q�&�k!�g�Q+>v��s�ƍ��.�>�\�GÑ{��"&7�q.������Tw��{���ɧ�P 6�sX1G���U*#�`��y�i�����p#�#r�д��h�V����b�x�h�	�#���v��F�)	�����:WB�G�������k�� *@�Y͛|�iLQM�в��6a52ހ����8N���U����k�^�K�|B�9�t DJ�B�9���$ �f�x���Cf����9V��?��H�Ms��2v�ks�A���zZjԃ0Sfq��\���rZ�G�)Q��qRS;��`^>���;��8��	���ߟi���U v�'t�ְw���xQ0y���x�v6����X����^=��1�� ���|�b?�;�k͇�/W3j�r��li�W��:Y���>w��Q�*K�Uy�5>�p�������p]LI��`@@@Q��}�Q&,vnd��8İ�PԠ��⼮�o ՘OS�����˶����i3�2�uÀ�EJ��Ŵ�_���g�u��H���D�L�Q�H�E��O)'�}�������W��6��P�eu$�5����1j��Z����yG�o􆪽�Î�g��:Ul$��52������b�@]���5����;R�{��u������a�g���h��l��;q�o[9��s����r{S4c��(��s��D��a�� ��Ïى������2�2kg:�������?����H6���>X/��0(��6���E'G O���В�"g�vǏ��r���,�r�#�RG n�z�LA}����ל��h�����Uzu��]���~��ߥ���<��z:
t�;���C{ktRU����(?��KUN�n޼���[���A�"��2Ss������h���k8BMSFff'�����b�x.t!�f�m���OU���8c�g���,�R����K��lT�PAb��(��3�b�'�':K�����#&��R�;�#�.�ב�� ��*�89
=�8y/_�D:*5������\����yf�cv���(��	P !�[{�E{�����@�	I4�c�I����W�ئ*�>>Ⱦ�8�ր�����9���bh�\��?�>$S�?M���g�o~����cҫq�!3�.x �:���Y<es�W�<�`@�V��dn~����At���郏1��<��o�^("�c-
��)Y%��x��3������t��*;2?K��8S�1#A*
;�ӎ���e�2���(b�v��(OOX� �j����>����2�VN�}l�k$E������{�
ҒiؙW�?���͖������XД���q�_���4w���6r~n�{7Fs��N	
ӛ\�t\����Q!�}D}�!~X�ڡ7.���d�|+:��a�����]�g�n�� �U�L���h�� �P��V�c0e�����q�"�}(���t*T_p��54�u6�G>J��'�&!��X��[Ħ�UE8F��"�{�Q�+��+�'�-2x�s���/�]�H1���Z�u��J�xvn�p�3�!�v���q�w�V��'c�{�����dbM�������z<�J0�&h����q�`W�od��Vk~����6�e����
����46:Yv���pT�ä3+��L\8�en>@d�:��~�����6��x�C?rr�Cm�/ΙZڣC>;4������%��#o;Z�呎m뵭�W���� vQ
����I�����ޑ���O��B���t�a����V��fZ��@�n_����sl�gKq�?�5�R�&]��3��q�w
絙0�ܿVG&D�a�u�@���.k���ާ�Vc�������Ɩ����Aj�%^<FS�+@��W��q�n���`���i�,H)���d�G3q�Ԝ��E{I��	�z�r��vI#�U��a>�<�e�¸����1ǭ���M��K�6:�d=�*���<��}��wI�4�!�ʫ<��0Ū@��IX�C�ɦ4���F�'>����UZX�k	�ά$�Г�!TJ�4c����t�M���\o`�YZ���J��c!�y�D�[Z�i��@�)�l�.X�D�U�����o�I���nJ4Lo�a�i7}Ϭ+��Ӎ��	P$��ZY=
�����J�}$2x]4&�����Zh��ȍg������뿨��5����2���EE,'�Dj��N�k��b��ܫ��4
��?��\+��h9ZJSG��d@,��K��⺧�{}�٥��c`_����]?ptޜ�d-P���9HQ�{�4�N�2,r�ݤ:�\#K��h�9S	f��@��
C��,��{��r8��Cƿ7�:�K芮��D��L��(y{3��~�X�� ���,ݿw�����U��G7�	� �㖶��Ppu���������3�s��]��`�q��pSD�c-�k$�[RkO����0'���}Pu�ɉ<;�I#j�_���������c�q��i��8
$��`���`��UA�L�a��}�g�̗���˘4��h2ŵ�Jq�����2'.;�T�50z+Cgv["�s:ݏp����?����'O��)!�ŗ_��i]v;1���a�H �r DS�P�g�}p�n��=(��$wK����γ�d� ^���"ȷmv~`g=�4�!/f�n天�11��h�bNX�:;�����Э<rb*2;��h��m�+9-l�L�6$h��=�:�K��.����t$M�J����U�PUc�X�B�ի,bT��-��������tc g � N���Ik�u�;'�d�U;6t,ܫ��Uq��k��׳ִ���V3�����o�_t�����G��G9�d�-Eqe��0;>T�v�8s$�~jg��.nxH�60
w\?b��w�`Z��J#Zo߼cw�����}�(}��ߤ��������u�C8wj&)%�O%!�ʨ�(���FK̶�,atVQ��9xS�N��/��f�΁Ŭ9��tW�GwN������2�&����!�J$���g�7[coLg�)���!�йu�=�uTN���Kv�������x����9�@�<m��x��\lc�9��3�0�0{�s؀2���e����Յ�@>��W W`�����%x�F4!�4��¢��>�i�������|�L� �/O}��[M�.�i8� �b|�E����Æ9�v�^�l�]��!����(��Jt�z��SZ�>�S���3������� �P�`���X����P5uv;�����������?~L9�=x��F�����E��#9��{��Us�W"��AN��]��M��{@|�@9�����!�5����Py]�u.t#o�]�W��b�#���ì����*���("���M�b|P���;l��W�z�"�������O��a�qv�M��tQ�K~a��Ӿ���8����M�՚����z�ܲ�}�5�h;Fh*�;��,�m��"�؅@o��!��j�̮�nZ��b:ho�����حK�/y���z1@d�;%��#7�
v��Jj�m��
�y��֓�uak{j}t��5�Q����`~h�=�>1V=�,�@�(�s4A�_���ۛ����3���}5�@�S�)"k�r�S=_끚��X�����#0�@B�]�N�ձ A�%>`1�n����J�;:�ٯ�r���}��j  :�d�]�q9U{�X;nA[�ΖzK��k�d�d��JB�d&�%�gVU��(�=��d���B��N���8�P!�~��N}aY��ą��WK�$���S��:�q8�V����b�Ꙏ�0&0��12�5h�s,?U�>�L����-�h��9a�������/�,����ţ�r��N=*(�| ���U�.œqc}�N�E<{��N�n��?;��ϐ����j�D��W����9Ǚ���;Raႅ�ʫXBS��;��C][�s���F9%�౰u�7rh�a��{��3�M�N�ǋp��҉��"e�}�,���{[3!>�l�Cx���p����D���7�{�b	����M	8Nv I�0��U��T-��7�?���!��?�6��8��/��pN8D�4��M�$j<���ٛ�ܫ`>I0Y��'`v�s��<ĵs�1�0@A�ј�KvR����v&u_�q=�|���?�ZH����~_P���K�&�r����������
̥h	���TЋ�eg�;�����1��N���|��m���[ڭ[���sG�H�0��FǨա:�J��`��=-�)	ƨ��ϰ��Q	!
�����6ة���#�*�2��������-X|c��F[=�p���J�罞���~'i�}��	�)迿�d��{��g��>�)�O��� A�`�U���)�[�S�օw���1�
JWL��:i����މ�$�ܩ,�dh���8�`�,��%��4����L���7ƙ��FI�m�� ��)E9Qء3�࣏X�"~I�S�'��1���r!ӛ�/{�k��Y��>�_|���.��k�8��?�{�.�WSѡN�N�6����n�x����,�d28'j0���Y0x��;����q������o�s��#����l������Qm)���w��^nb�" ���=l��,M�?D
�R0p��3<+����Ϝ��(K,�~:�` ��a�U�,���~�����/6~�/���K9�J�5ڦ=2O��m.8�V^P�v5��js�b\���:����0��~���!
����x�{���+�|`��ȃ�q����d+;�қ�s�_#�u=�2�c�M4c�b���a�2J7nsE��!�W��/S����x���<}��9���V�|!�nܻ0m�?����RP�qT���jv�V��=�x�é�������n�:�vgS���A�I9)��d�,v�PX-M�/n3C�FWq�	0m������Y>�����##0?�Q"����Ƣ �F#��k	H�ۑk"�s��G��ǟ<L�0�g-��Ŕ.ݍ� ��=6
ѕ�/N*�j�!O��?<�����Ƭ��8����(�:�e��&́^}�#lT�rd�l���M�<���s�!;U��N��y��@ ��/����v���Ң�`��;�)��(��,NL_;!й���ʻ�Ő����2X��R�h����T���+,%�w�\�f��Գɵº����<�F_��.WFLfD��_�bۈid�R��l������QZQ��e+׳�m�gÆ	Xy� �h^ծA���&�C���˗�y� �T�8C;-\`(�)���{Wb��*yCܰp`���`�F<��A,� ���g�܀tD4�X�B�T�s��k�{Q߾}� N8���GG�).Cc�ƍW�޿�r�w)��mw~���xt̲F��3���!�9Ox��X�;�5��U�w���df�����n\?�l�W4�>��qy��=�ז�?�����Hf	��s��g?�R��	@�nSj8$��9��΂,c�??�>ͮ)ί|����m�;����p���b޽#��!V
g,7�Q��@��c��l�gQ�LA�̯o%�������W?��?�@M�o���D%SU{�to��`�bG*>x����w�2�� K�.�z&zj����B���ō �F����4�>���>u+���;'�2go��i��������p�,:&";�o&��ϧF�d,`ØL����i�	���ہ�C��>��E���5�*��NIƥ.���k��$^�"�&��զ��k�s-쬖������|����pm8�pl��P��ޢw8�G��s���E��Y�( 3���l$�=���0u�*JN.*	<cF#=�cQn9G���X���>[�l(�#P�"5Uo�Z�9�5�ek�unO����駟N����.�Y�\����������4�����.���7,.!\�^l-���ҁ7���0�O'���˥X>���F�uF�c���
��,��q��q�]S�W8�;��q�w�\o$t�g������ۦ��%�ų�����ǔYT�W�ww�-���R�o,|6�����Y�|/� J��;�}G�7�Tξ'����ω3��J�4;Ԙ(�ʵ)�:(zV�E���9�D�B���{�~0}�#�����ՠy���su�²�:�W��sGRFaj�P����T�M7��W ?>z@��|�nw��-�N�t��V���d+V��`�Ѫ�������[ٝ��Ϲ5X�Y�L,���<�*t�x���Q
}�����ي=��.ƑؠH���6wO%Lj��6wɰN_�|��`AAs'��������������p�W~��E$zȉ�\�Vy���!tMg�:h���k\tu@e�CW+i�-��Y عwF���HL��Ȣ���zx_��Oln���n�VC�}�ZI?go67t�b��m�l!�ϔz6~���i�;��p�C�&_d�F��3�EaǠ/��b*z�T��{�|bi��wa�:�]͹�S��0�����MJ���x�	s.0�/1/#�'<��[k�c^�<����n�鴸u |��2K���]�9�)��E�Q�fi�r�`�����e��B/���l��/�W[Y�~Ep����������}�f�Ջ��#3��|�݃5����Q?�����>���_�����W6�~`Q�bԥ�X�¹��~�<{�ZS���/?wt�O�aй)Z��p�_>��8�ء#�󜮣�#i�M�n���/���[�|�`�����S�DE-�X��k	{N��ฅ=&Q�}��X���(n��_�i4@����癍f�{�C�oʎ����]�k���Ad�OM�����&���%���NU�q�u���Ġ� �#��B��9�RZ)7*�g5F�56s����&9�i�C{������L��'X�8[�Ɉ�?������cӯA~[�檧\��i4ymFaky����`3��߇��"���F�y콗�Tʼ�gc�lS���� <��o~�i��Ӈ���{l,<�����N�~|6����O��RX�����e��dʱ1g���g�\x�L�Qک��+��1�	�Kǧ��f�h.��1� ���#��E�q�Ԕ�s�VB�j���7ģ���Y�UO�Yq2<��H�g10������tƪ�u"��$R��g?ԑ[���_el���Bi�{2Htp��	�6(ӌ��|�H��*[��*K�ǶA��k����s��?0�#~Oh�|���|��)���k'D���HV"���	��SB�׀����H�nj�d�PUt����Ʀ�p��$Z�]�PEPo,�3����+�=��(�bтO���=����%�]j	ICh	��ۣ)�MH,�D3M�TP�U)^�b�1H��t�n3��7�@�1k6һ�#����S�0��]2<"�cI�$w<[�}a�I�J�����D��!:���)�\(��.7b��ޠ������|cހU�/�����ZX���%�5�,�*�` �$�F�k�f
����&ճ�;�?���00M6�M��?�qL:?f��L4
	��cg����Ys�]3	�J���_��/�)	;�؏��k��zt�m9�C0���N�-���ښ")��x��	�<@�Hv��P�'	��f�
k�q';���������1�>� q�?z�׃�C�>:fru䆣ds��2�'�Kb�H�l,}����O����x��ȴOd��܅�+�ಅc auXD��� �J:��H��@�>���L��rC�#�G�29���T0 `�}G�?(f����t�&bim��jo�/_���
�[2���=W϶1o�nz�،C��Q7����0���p�����yŘ���״w�χ1)F)��� E��4�Atي3�αO�!�1�)h}�Y�qLlC�#W�}�E��U������� �3O�n{�D}kr8>΍�O�{$�uP�X��{��������϶d5��_�D)Eg.��c�s0���*}�f��+��&W���,\A%�-�>i��\�J�߇�tJk�&�1�"�����&#? 0M�q6ӏ�A�M���Q_�oc>*kͥo�d �c�m;/w��M~�Mz�d�����R��"�wZa��CM��⽁�gkK\9�f
HSkSc�<�A��`\/
Ъ<��$�����r�P&�i<
$0s�G)��3�����״���yu
v����T ¹py�X�xQ� IU�Ejc��`�T /�a�p����=�5�g-�(���_�>gW��/`�M<��cN���ȕC�R,�����6��Ѯ U�S���������i#9^��Ȗ���6
}���5fR�b*�Z.�q\Z0J��r���H�pU�a�κ���>p�h-�1�x��s����f���ɓ�\�d8Ng;��>��3m���u�:�w�aϢ9��6P�"��m<��|@ͼ�%�:1g����~�!j�D1��P�C������b�7����R�}�˺���Q��*�0�>����<9gca��_��rp�n h��J�s�Ese=��W��Ҩq*�4���fY���t���Ѱ�)���~5՜���
}�h����uޛ5��#�� }h�ɥO��X��ch�T{�Ҫ�[�@��q,���c�j��u4�Q3�n���x��z�V�oߝ3�{ ��2�<��9f�)�fd���z��Ca;�<���h���fS���VU��h`�V�d��cf���ȸI�rK�h�_.d������z��^P�\�O�"���8�F�=���Tq�ԈXS�q(a>�1�v�vR~Z�3jVNϩ[,��T�~�M�����`�v@� ԙ���|�e��(���b]�i����W����VX�C�R �,�٬�ݸ`}�"��6��t��������_����J$�t2�@ q���+y:mFPLQT@��A�=��"e��		/���#���q��&�9���I�E�:�=AO*���p`�5֓��lܶ�!�$�r��38��w���+�`7��;1����`���\�����v^��ͨb�@��͔0^L�kG�P$_�,:O	��w�f�쥞>ǤOO�be8rGJIV�[i<�֮'k��I(Y�b����!�}7mt��_����9���*6^J>���sǼ�ϯ}�z�n?$�ՏU9CE���2H`G���m�\P	1Od��G����W>�����]��#n�����;�,Eý��]��ߺ��S�F��v�X��'�������?���>Q@bE����`�56�t��&�E!��[������)����m=����Hd�I������b�&�H�6S�C<Pkc�B)NH���-�D:AT���-_@4r�*�,pz:lL��7���"��C$��R�X�:�]�&���;�{
�z,�ۗ _}��t@aO� D��:;�܉���*k6���30�loc�#���GϾ[D?�sV�4����P* �[�9~�"#ƞ �f����HEU���ą�����)����㴞����Ӓfe�3XxU�� ��N	�}K]9$waK-���p�d!�?���X��1\�Q���7|>��@3vz�v0{I�ȺiL9?��X���Xo��4�^�f7�E�ON�l�ޠ-���k��h�ݺ(���
�NL2$��}�q�� GaZ����F�����������A=��L@J��8{�+��1�;�z:N��z44nXe��1j���ֱ�����<�ͽ]��h"&�|���p��ڡc��G��򮰋=r�Gg�%)�BC�:�+�ǣ�H�K�-�%q��/�W��2X5m�gF�ʥ,��*1�g�f���i]l�Y�;�'�mA���[Ӵ��,�k�3��ra�Y�ƕP���b?����Q^�l z�ni 3��8>��K�b̌5^$W����/X�K��ƞ�B�^EхG�������"�*.��.#Sl�{1���)�7��5Y�����7��NX�g�NF}_��Ž k/�̧�>���������g%D.���Q=�	:;��l\�*�d�]�X�i�gc�"�@��<߬������G��ŇzA�
��f��E�cm`BQ�Z/���/�놑Y8Ły �>��'� �쳻t�T���c���m1&����5�ٚ�nU���A,��6�D�PW��l�,r=�Wy�Q����M���9��� ᯁ��ueEVgE�mA���u�z9�I��a����'�w������wc��Xp����4n��dCc͞1�_���x��,z��1AH�Q�0��� �����5�����VގR�ǜeR���<_3!\=�.�(&]Y�|��u4�Ƹ���1�9��bG{3�S�pm؛o�JO���,�\���>�4��z�:�
`a��ӫ���mKS�}���xa *���b����= @h��\H��<~N�&� Ǻß������^B7r!�Z\]K���>�3c��d=��dv5�*���"x�|��cL���4sO��S��Gӵ�����D3v4p�W�|��D�I�yl�m����*����X5�51�ڰLP��s�M��fLj,�W*��MFǌ~�h��!�+O �LR��V.H�:��8� ���G�������1��%!���럢�6��0x�V�}=����4B�2�|�=�]A(X9(���RP/E�Kai鸁w��\F�2��pw��U'n� 5䜒2kh�8�X؞��M��T�^�Rn�Z���>�} ��8�!`x��6��,��I�S�X�ÉEz)=��V�T�pi� �%HLՕD���#21�ε��x��_��|�����!�Sў(@��$�+u�  ����-���m�ބEsʇgg��|���XW�bw�؎�	�1�S°!��b�۷]$�@�c.8����3>h�~�M��oI��=!�zx��uE4..r�X��+�༾��O<�È�f$�1C��A�+���'sy�?��}T1�'�4����Y�G9�&�de�����~�5���z��X���?�����g��=sb�k��@|4�S�p��.o�7�o��:̶���w�"��1v*)Fh�&$3����DG'_E��!��l@���!�H� ,	Ř��l/�z+ɣuv�A<�M}��Y�	�Ù�4܇ Dv�����ER���l54�޽��ͷ�Pc���8zT��}�J��%��fm�����=�]����D�ړ)t�H#�eZK�ȡeϘ{Q���[ Y}�!�k2a����(� G��`� �¹���@]D��B`c,`�����>�Q�+�Z�+�֎D'dQ��7C��u�5.4qBc�sb�ki���������6~� ����R����bU��+N+3�c����vc|��g�O>e�ͳ��?���_O1����DK�p~K�D�Q���K��,�Y9G#(Օ�� ��R���"�*�]0	e��_�(c)��4h��ƭ�kx����=���aqe���"��`b�:f���*�Jc��	�O��4il%���)����2W3�_���>1�y��G��x��:�#�)k�ঋɆ�Ū�f��0�ͼ��죎ړ}B8
i|��.����@�T��Y�*�¹)3�� 9�e����M9�2�VGێ�&��(��q>�p�����'7=m��Eb�~yqM]�G��O�|�u��ۯ��	&, ܟ�zG ��y-����r'䰡�w�u#ܰ1c�̊��o��_��v�#�,����h3^@�u��^�'�"���$��p�oȽjL{K�O��8�kP����Yν��k�&a�Lg�AE� F)"ł�$S�W9V)���?�c���$أh�7n�������أo�K��a����Ќ�E�������Y\c���F�$�� �.nr��&k�f\k�,	�0q���Vǹ��Ln����|��5Ǒ^N��s1�#��=���5w���vY��Pmu��lo!h��k�5�*��e
@-\0���| �L�5���w-��n���邅�ʲaı\ȩ�����
]����g��/�o?���=�����n�L�`�$�'�s�@U���H=��>�n����^?�o�����J?�q�F�F�m�SWf儎�BIu�~% ��Ɂ�[}?��W^{��cd�`Q���X�Ќ���w��·��u`�/�<���C=��J�������3���<��8�
�s�Aӡ�G�˳}V�nU�7uM�l�5X�|�އ�� ��G�޿�|ވ5P��-����β?�"�GL(��a_�9�o�6��kb�I�����_��ųN��my@Q�`�)����ߍ.g��"Xld���)AZ.�JU]T���#�h��Cg���@0�D`\���p ��ѵZL���D����4�	�O�����]z�B��t��]P��nwMTV#<X�W�|J\*n�p�R`m���)���>�1[ �sZ�����+q^]m�0l�w�%`��dQ��3�����܉�Ϝ����3��������H�!k��łg���������y�&W��7Nb��LR��5�?�����3u(�g����q���U���X������B19ػ��KO�>I��/�2%`߳kA= w��U�)�P��h�ִf.;vt����nz0#���j�!��Uj��v���1�CL�W	nT��}�!Q�i4К>C�����E�`D\_�s,��SA'����"�Ҧ/��[2��Y�f��#l����a�Q��7	��p���)���˼_y�j�{/�*'�S��l�x�p�����E����P�}#]��{иgx���Ku*�,�}HJU4��@�FN0x����<��J6��o�^kܟ� ?�/��� �����,�H�[Iz�I�Q����˝���O3>*2X��`��9I�0�nTX�AK���و�^瑷ڎB e���I�DMEA|�o�| y��;��"r�_m'��X7x�
C�V� gq���/��*�.a\���*&��� pi���f��3[���i�,@�Xb��0���#��|�~䮋���4�>��4����(���xZt��P5��#���M��y���/�w ��Z��|�����p��H���_#��%Ǿw=S���>����qV�Nf��+�o0�]\#�qn�U�9fTh�g�ݒx�kٮ�5E�Ty;�^ӱ.�1k��w-Y,3�	 ������9�{ (�-����k�q�'RUe�� +��WY`�v��zG�	�2��N����v����Q�BH���T�(�)�����*E�
˽�m��4>���r=�Y�G�w�%�$�����|�y�F���n�?�����1";�;��B|F<fC��_p^t��h�
U�Xuh�|����c���oix�?��5�:�§��n����E�x�7��]�� �Rf�GQ6�$�@Q��狟�=��>�Y)����W�Y���G2ϸ�\���׎�>{��, �U�*=��8�.�%l����]l�Y�ǫ�9�<�p�ԁ���NX>�a,v���	b�%����#�-�ÕA�`��LE�#a�_>�o��� pn�G�G�*��N^�sn���V���p���B78�������O�C�"k��U��`y�=����A��f	����؏�@����ߧ�o�p�����`:��Ff��}/ܸx7�!�Si��d�701T>�f�� k?w�]Ƒ}��r���Q� v<���L��y�s�=���T0�LA̜r����g��vʭ���S����ң�>M�7_���ۿ!Z�Yk^7�`���5�	�-6�V�U����/�G;�nv�^/Y���۠��)irE�iCPF�L�v��ޜ�&4v�I+�39�)&Mq�jcrD�#gn�DlJ�\��F@�Qu�3Y[R���_�\��}ޟ3�<FL�et�0R�e��?�`p#L��?|�\E�����!'�A���ڨD}����T�a��3�W�zH��֮���Jsb�B>t|�f�Y7@�����D�7%2F\oxڇH�8݇�
#i����� ���9�x�qP���P�6�z.ڈ���eD�$�h�kAK�"�L|`|����
&)��M7��=+�f�G�z��?,�p�M��U8I�x��9X3/_�J��" ,! 'x�*XN8#��s�O�<�H@���g�+1
�e��q�N�5��`��>P�(�p�m�5�#��\�0�ű�)T،ô�f���i&R^+�l���-E�R{�t*�*Z2o�A�.�NjS����Jc �AtPp�6�9�A�.���%����#ctU��P�(08�8���[hE��;w`}��`�aF����'b�c2\V6W��F���J_���������"'�����Ū��\����3���{1��$�9l���Z��.t��,�e�{��'׆���� D��-3�\���mR��|$��9w��-u�.�x��B(�!;�Iؘ����N/���{Eg�h$i}e����H0���ܣ��W���X#�HǐгPP d��`*��g�cY�U�#w2PL���+е�=�a�^�}F�l3cf�$�a`=�p�b"�{�6���q�*d����O�1�|�^���N�ݣW/_�/ ��c���O����B݈��<`|[;�H)F��(��ܢ]eP$U! �3%<��-�f`�`oØ��I=
J���H�y����ϧ���)�]�lZ��v�A�1Ǭ<F⮻@`[ֺ؋��Fj��:M׼f��a*"�����aP��?�Xc�߳��1�q�Sdp�k�.^�_�4�:c�ݻ"j.�JrU�����׊����b雜�F0-,�Y�QͻY�M���3!_�_�g/A����0�l�-ئ����Ç��\��g����5z�hd��>��
����1=ק�~xg�ĸ��cϝM����N�f �k�f��J�f���Ȭ�B���B,�n�S*���� ��d�4ʎ�v��=:Pi�u#f�⫌1��Y���Jl/��ؓ� �0Ҁ�b
@ĝ��i��@f"���b{�]��8�o�P3�~g�ޑ�*�/��4��z��(�Ԍ��,�����*ǣ���P��'b���S���$�ܸ�{֚}��ӡ�{���a�f�;�\�Nk��][��֡m,8ŹGM��[칺�2�U}��-cϟ��U��W"cl�%��[���.f���s��b1�Z���|���n�ܙJ�'G���dS�ռ[�����dFK
�NaK��Y��A�����ƙ�z*z�o�����Y�t:���s����p_|�E��7��[�3����+�!D��?���\_�yc��;�}X4k���Ά$^#��� m�hQV2�B�)��L�� ��{��p��ׂ�W�Kka��K$�X�"��c��B�. ΰ
�)�)i�� �}�;��1]��(�iok=�u� K�h\f��J�Nrk���H�~���?��cz�l��vY��c�ШYBA���/�:�g�4�J��V@X 1���C �خ^`D��ͳ8G� �轛y�v��s-��Į�j�}
=��nPvd��Ͼ2�����V�dG�{��u����w������y�����GC�	 ������M����TBn'��R�	Ș��D4#0C�h�D�Њ���p�G��j����qV3}��ơ�kw2z�G.�A}�J���<�bU��*����)�Y|u\��x��d��k�R�-���l��i�7=Ѧ�)�:B�"0t`g�7�_�.��gFD�$��r8�*�kA��&Fg*�����o��7�)���Xx�ћ����������>�A��#6BP��Z6sr�J�_W��!q[F]�0�P����A�d��rqɩ
+��l9B�/3��7HCvX)�1JU�~��F�F��9O�=�.�~uN�'�ݦ����80��ߣ>�s0fP��~�*� �<m�������h<=�����	��7��9==&�E�r +c���3��v%&�Zv���}��(�k�':J7��?�t�ߦm���N'�K��zK��f���m僡����hU��z8�-����i>�@�䀙��G+�	 UXB�h�}U���M��:�c�1���P�*�uFW��9�Nv�`�<���N��v��n�{��O=�7=��S�v&�*:�P��4�y`�]��Ϟ�k�?
���޳H\���%ZI��#^g̥�������=�i�N��n'elc8`� �HХ`2N�E�?X%C�g!��&)��QP��XG��rJ��d�h�)�&(@;��`-����f|��򗯹���(�xɅ��A��2�����&�qI�`�QU��A�/Q��V�{{�[������ݵ�O3}�u�)��� qUUf��{�="AJ��٢M

Y��ϟ�� #�ʓ%ܿ�HĂjG��Ҿ���{/�~��3��\FD'��Dw�t#�;�tvv�!H5����D�ܠ:iMg�$J��"���� �c�����D��$�8DҳAa����ɓ'�V*j9z��)��	�� �LQ0��c�9J;��w����� Y�ֹ�!*j�lб����HFȈB����ܣ\�6�U�K�(�����'��e-���|�=����0�Vݪ�����ę�6��9%p�"�Ϗ������g&���o�B訑s������2=-�st��.�����X\XП�Ęgڿ}.��QR���qB�O�F*s8��k���'],VM��]��dgl�ޒS�S��K�v)����~���홸�uU[s�iͶ���Xޕ7�\@�1�=�,G�>�>��3��O�i{���^���w���.����/����"�%ܔ;�H��Ҁ
g\��)�hGc���ǋ���:�z㱖f��5���Ṉ�Zb��q& ���(��z���}ИF_TAn���E<A҇�v�l��׼o�N{{�����h'?�3�DL�s��|h�{��:�%��M1,4{r��B��*��|���$mr���o�$�fF�������7ƈ�_���a%�$�%����E|���E�3Uni]��o�����;�w� v�IG=haR�ۊz�WZ!ať�+�Z?�zԀ�U"fp������O?�;�n��)v�u��BN��Mc�:Cə�ތ��u�2�-�ww�$�]�����YFqt�z9��sRN�����9��>"�
[�,ԦG����@&.F�P�r<$�p���� a7�齗�8R���� ���y+1lr�����[)���
V���7��eSdIP�Ϲ�C(�7����ox�bgwe/[�H�<6fj��~�N���m�9;i��0נM �������^y��y�˙\� L�8�ҙv�ŋ�x�m�hz��b&��X�6�ʩ�c�f�s,c�Ź��%j%0ԡY�����L�w�QM�֋E\�4d��/�xm��lT+D{62�i���w�,`��>9��u5�͉Ћ��W�5tsq��pf��c޷��������y��Z��bVo��lB.B����\�Й��K��bb��ϰ���.���E	��idI�d	�\���9�Y��ė:�8��Y �l Tui��<��y�*R0ԇK�3����0�[c>s��G#�8�g�d#�AA!����7����)sӖI��z=R38�0s��!���{}�j�3�h���T�r�:��g���]�iMp�+ɴ�V�6��䀔,~3]:�h|'����.�FxDW��H���\ �ˬ�tm�Fz�F�ႁ:�l-�h�BJ�� ����̃��������.�
)N�Y'ĝO�I;����8k�䆬��x��P��k��d
�%��B�(hg��+e�
R1k��.4�?�x馄k�pbѽ��W��A�ߵ����Zc����ǰ���O��)���:�E:�v�8�����=�I������q6� ��c6Y!s4.�Ś����2�	X��t롬IO�k��!�%��xv�z@�P�QrK�=����<���1���da��4�&�ҵD�`o�{11�|������8�X�nv��n�ة��9�����8��&��l?u�p�����x�"���=��B���(�����q|�1,O�1�� �q����b­K:@�eR�4K�M�D��`W��u�B�Y��{��	��5�~�t�Tb&Ej��b\W��J(�= �^�|�8�@�3���`�M��իW�Ν;V�Hf�|C(6���y�y"��LL"i����ۮ]d��֠�,�;��'�w��c6�(�������V�	$�`�v�S�U�8�������|[���.	 ����	�\"3ᣏ>RG=}b��R>E�\i*��6�P�)�����`�_L�@�(ȳ�v_r$u{g�E�b
^^׋�fm�_&PU,]6$��:�5���"�δ3AZ� ��ĺ]�w��|��㳩�}�V��me��KLN1�c��X�5�C��s#0��A c��Yu����G��s�7��~�m�Atn��k,�5��M{� ~�>���U��Km.ǒSEoN�9�T#&ِ����`|�d�<3�,Q����� g�֕g�R�jd-G��&9�Pb-.�#'"�R>b,�um�5ײ�ڄ�k��G���_��p����
�~��(r)+Z8b��M�`��>����p� ZHM�d�]�mbM&�,8k�Y��s:���HK�1�(�>��\�:)�͠�k�#ʻ�E��.�W�\%�:�70�hW86�������|��Y�Μ½Z���lb�#�>�*��Z�MS�52(�䒅Q~וA��c'��Z ��B��Z��ݑ���x2Aƒ���`4�4��+�p{K^�;�U�Z�d-Q�/���銅�&�Fd1b�}/�]a���`�$:�. �'��ЩAt|rd�2F[R���
�ot3���݁�s(2��\�zq��ʟߥ	�f���M	c�N�9�*g�Y������C}��F�'r��������gZKəHl讻���ڛk6Ӡ��G�j!�UA�d�rc)�Y)d�����x���zڰ�3� G�!aN
�<FyCaD�,l�X]�N�/ҟ�Y��o�n�\���t}��Ϻ�P����b� �[n����;��u��������lcngn����$�@4�FOz����8L6<~�0�>z�����������)Ѩ�1k������%��}��P��y�ѽ��Am�s?+K�|���������W1d��p�t�!�ټ�	�e+�VH;6Łt>����V�+Kg�F��A�;��]`����p�ޣ/��]�Bs����;������D�@�,F�֌�c�X�A �U[Z�U��N�����y��E�r$t��sȥ< fM���ϡv��yt]��*������<��6�	����iM5�-��1�V<j<Ek81�i�"��k��w>�r1�C�P���[��޽J0"��F�Mjj�`mTE��+��4(�Op�Rm���or��Q�h�?���X$�;gA	�*N�kŬ�O�h^��NJm�����v&�ȃ�6���s5i��`�ȅ*��:�uv�����]$�(�u����������$^UEDH�<ۀS�ky�9�g/����� u�VA��X� uv�2:���h��Du��m2L�X�6�U���y�N����?I��+2>��8uq6���/�=� z�����	ш���ۤ:o���,e��G��[;��[��z �sr�"���P�I����C>�򆰍�8��rR`⦞������KS�q�.��;��������e�	���� s���E�2��Y@ٯS�Iv@�N�!�@�d�,dC>�#ˤt��w�K��?�%<|�����QG�&h��$� O�o8�hE;�qp �>:YN!F�̱�������
�jj�*�tv�%���,�	��[q�=I`9V�J{�kM�'X��6�:����f�x�⟒#�F������m�������#�Xl#)�����*g�X�*�.�KW+�#�a�R�x�Hی	b��`�'	��hm�# �?X��������`�3��7��®A�����%7��U>n$���3�|�
A�7o��g��+q�+L$�xH�q�ݔt������;��E���E�	;�`F!�8���׼d���F�p�	T�5G&��]��b����^"�xp��S�>@Y�:�c]��+�fT��{�5P������;+�ĿQQ��Oѥ�ц�Eџm��d>���3�u+;�	./r����ox��/]��	b]�6��:kx�&$��&�HvP�� ⩷����1�Kg�<����X`��� �o`:gc������ڢ���AU�kƻ	�}o]b�x�¿����8�Ou��Nѧ�d��|�@���
�31F�3Q!�x�����F�.�{U�9״x�G��9
V4�ܾ�O��>{����:G��c;�؁��ǋ4&m�9|4@c�6v���l��=Q�=��A�<5�'�N	�O�L�ƚ%Ԉ'1Nl$����_�N����i�������6���"o������7���G��(�NN$*~5�I�<�s^1�q�Ίu�
s����_�/�hHp��f�2�t�\_�g��)���,+$�q�&���cX���Fg|�r�� �!��<�������V�Fns>���`���X�C�,���&����&�%o��d����s������͛ײ�-��@�ZZ7�n uf#�{g�;��Y��7�-��߂X<�R���F"��t{��u���5�<O`�MFs�C��v��͑����!� 泍l�2�@9��`�K �+�@�����9�|r3]�e�T��)]�ȼ윍�sMS�dE�Z�gGG-�(ϓ0�:��N���ש�3i�������i���E�E���cs RsL�iM�2��<�L�74λ�k&�-g���I���W�]e܀�4�ڨ�5x�嫒'eF� Zh/��Y���ux��<ܽ{��9G`�L�$xn��@P9r� ��|q� ���������*���s�ɒ��>�O����8K,�Z�F֝I���>R�q=��@z���� �Hp��e��M��tG2CX��R����\W�$�qd
5W߁y���˦�����a@�6�h���p��Ze5�WguN�O�cE=/�z��>�Z��Ac}�A��;>A���'
 2-8m�&��3�]]�g��z�i`em�3PG����H��߯e3c���>΀;�k��A�/0�֭�cM��'�9'����f&CP����X�8�-;��?a� �~�o�"���b�a�t�Ff���ފf���h����y��,�>|n߾�����[��/�Ћʥ�l�]�p�e7(��>���V�[\�>&�}jZ1M;V�7*����ϳ�/i]i����P�t����h	Ԣ�Uv}.�鴯��q�gs%Y;��Q�3�x�
ߥ����N��]x���uK��K`S��AA|���ȄQ�y�V�h����ܙ:\_*^��G�9#,������\
(o��#����n���O�e���Au|�̡���D5���C9b쥂���}n��v�Y�c0�� �y�$��e�9��{t\���N d�"/�5��Tr����{�\�vL�	�#�1�1 {��	�f����gN��U�m:��'2���<���捏µk�	��� Ȉ���F���=��}������R)A�g�_��)aŭ�zS9��>���7n~��>�����.�>(F0�����7 =���w��/>gэ� ���]�M��D���ƘmY�!'����'�m�3�ԓ2�G�!׺���˔��S�����<+ P���#�p�naS @�`���'��&�;��(�K��f��2Rl�f��b����d?��'�Ł�2\���g�2x�Ϻ#��|�N֘D`������ 8۱�3����%�Q�*�gq](F'�d�5�k��?|�^�B���fF_�ؖ�j���1b��'�Q`�e ��<�G(LR�b����� ���q0�&m19����>���4�e�[�P6J���s�b�1����TH����ddVN7r���3πښ�r+VY[׹�t]!2g�u.=�C_�"������` č1
��JqɬY��������͛7(�˂��訃]"��9��`Z� �3���YN����oI,�u�����-O`s��g��y�t�p��9�Y����X����z���ҡ��/yN��6�־s�m4��#�	!3ɰ?v�	��R�� _ffy�E����t��"���t�м�r�`&r"�?�i'b��p�p�<�_|����8cHl��l��p�50�oF�d��..�f��@W��ݰ�\;8���� \�z-|����߱ل����������	ݭE��:`���@W�kH�3��|ο�z������s��G�,��&K�W:�yIT��T;:�����8�
�����r�{��|\���$�}^K(�||Ӛ��EUqcqP��O�̞�hmUƚ���H��4��x_����{���zY�贃�t#j�?�Α}�]��c����`�y��h�z�E47I�z:`��	{{/�����@`�0���ݶk6~��ׯ(����+�3�dh~�������}��%�Y�R�06X������Y5c�����{��NҵbO>���d4�?~~�w�9 ��'7?_|�9�O��=�\�2 ć^��S���1�{����Q:_�>d�:��~�	�`�ȁ�C�
���7���&��&
ٖy��TCH��P�]C�S<�,�����+�`n�څ���Z��߅tmd�u  �3�TgUf7z~c f#�j���Q�ZSM�*����8V�={ㆴ��:u�b�i[�~�����JyWZ_�~��5��l��1?�&)X� �� �fQ�W'����m�K��t�|6G���*���� ��؎�Nڍ�<�Q'���g�������~��B��W��aod+g��
�n�Y�v4�����5�QJ4q�氧�P�jK�~`�!�C��|1�2m ���֔�*=߃7��k{)8Iy�#�&�:��i��c�@����!kW���P���/���Τ��#,�,�����m�{`}��� !}�B���'Pj��:Pa���ek�
ތu�G��g2�B�g� �6k@�a:�C8�z��G�u��4�kS���5wM���=�ש*�����g�e�:s�D�U�߹j$V��Bj�_�u!����B0Ut�;�yJ ��G����K���vUTq$i��삔��3�QT��r�;%:@�%�g4d��ւD8�p��B��ә=u#qT�XSa��s�-.�u
���8����nE_����Ϣ�C���P;f�'m�Xc Hir���d���B���p~�|�|�2i��Z�N/�Z�Z�%��O�%����3P{�OM�Dp���Ǉ���_R�p%��OJE�U|�`SS��V��ИkE��~��Z�.��ӄߍ�{µғ2�.O����|����ҝZ�g�md���XV��;(��FD���])8m�}���1F�.�$U�%���'�
�����s�s��zlIY,^�P�![�b�(�7o|���e2�XY4��
;���׿�5�����{��[֡\����h)(ч����D����v��}���?��G �%%t���{w�����<0���\:3bF�s��ܛ����Y�3x��L,� ���0��=��)V���-�5�xHP����`�d���[�֭�Y���Z*F��p
��d݋���3K�"��-�a}EvQ�x@g���רpM	�]�H�3{d�ưhYܟ�t�u�cM��Ȗ���=h�JM�ȃp�:�u��	�٨�g��:�Y���`]�w ���@FXm�����9_{&�[����ZfG+j�������FOvwY��z}dֵِlc�
�#���T\�����c���_#��G!�92��&G���F�P��P����0���:�3�MC�b�siS4�U�w.Z+W�� �d��B&C$�.!}�"�!�f�;/�������36��릶1�#�`>����_�[f	 xp�P\�榄�R�P��  �G�`�5x[HG �Ƶ�\Tf{�Jm���g�@�^�-*`G� �4��u�3?��o�%ǮO����E.����f`��2�Z�
�<��ݵ2��Ā%�å-�a�d�� �P8c��AgZ��Z�6��?�A��˗�LT�d�1e0bv:B���� P�ݪxC)��2G�frf4���x�*n��Xec+b�(s7>�s3� w�b�t�:�8D��˯~����BW;�sC��5��l0����n��ٮ랹� {�袹�9ld<�>=���4�,q���_��	?��f�yf4�� ?޻�����JA�%����k��A|�[�F�3 X�%�3Fc?�Cl��mͽ;�ϥ.��.��/�������:#Иdk����L R����^�~-|�� �t�a�r�"�1#�7���92bq���5�zK`���o�M�|W����W��`��"��Y��wJ�!�"�Mú�>H�
�~ L{������L@�W&����-�z��o�CK*���^��p��wt�\C�w��~={�<|���9	��ԭ�?����?�1���7n�O�{|�b2��O�Ѡ��7���)c&�GW@�H��+jM����[Z������sc��D���m�)`� �����99�bMl�qM��̷A=3X���1�M��(ʾ���y.#�kmb{�ˀ����[=��y}�ۧ�M�NO�=����k�ir���F�^�F����~!� #�S>?������������*6����vkMY�拏0G�.r��y�1I��IvS�kw0׵_� ]Љ.�=�� �7  U�<���s"���6��@�T���CE�-��7��b���:F}?�~�I4] F�Φ@sz�'�6vg��㣷�B݈���|��4�!�3ՙ]:��p��ɓ��=HW)>�ۿ�{����/��^��`$ϟ�0��S_�O�o��ܴ�{`��Y�A��ެ��=����mmAm�,c4c��qo6��Eݏ�F��b��k71	!�`
 W�t�u�;���w6����ly��I61(�۾�F��=�*���h��E`�H�D��9��x%�ћ5�	B�.���f'�	Y��t�ٕ�E�M�'���(k�C2{xp�nz:��A7P��E���9��[�(��"� c�������\�(ex=��D�*��L.q��剡��t3��IX��3���Es��Q{��������7�]�.��(a�E<U"��ϟrC�� f/m<TΎ��疔��;��jO�
i�:X֞R̪5ď�|���ԡ��`�;�fm�֤����#f��ͻ�Z]KS���`z���)Xł���ܢ�,*�Z�0t�[	 !;G��������|���Nu�B�d�3���O�����y$bD]uǪ*x�������=����oܨTi��ֳ]�;y�8�KO��,�h�wO!����z5g�z�x��~
�k�j���;N��i>7��`b�8�Y�tf�h�]��-��@���^E1����y��b�x= X����g������Ք�!B���@B�9��dX4�OS�����>%�i�I{�>V���v�xϰ
�)O��:}���Ӟ��s���� �ª!cn�	� �TH��p���;X����b,��<v������
79�!�)U�����ڬ��B���'��F�����FJ䤧"^c��9DeG�����0
h�]��Ae=�n0��ƺLP��iҵM��XG(<}$��ŋ��鳧���/�36ej2-De�<�؜mlv��� A9C��rkxc�e'�,P�����@ki1��-���L�}t�nܼ�qhGt�D��G�v�Us�虔�^{�?��7�� R�����~`���6�Z�]>~��y��+�+�4.��A0Ib�Ɇذ�b��8���{���+�q_�6�M��GN��qn��q�MsF���%t���@� �r�4۳�\Q�l��0 %Sl�l�z�f��0f;����z��)�nɮ�}E���<�>�M*�j�Yz������F��^��H��8��hAu�.~���ڂ��M��nƽ�x_8_[=w&'�>�pm�Rh� �E'�����`���uLl@�Nq+�����3A���%��1��&�C�;��(\P���s=u���W��U���Kͨ0E0Z/��>��6V� N�4B lxQ��"����>_|��x 6���X�����#x�ljMJ�a�/��ɺ8�5�r|�ү�A0/윭�{'��������FݼH��jZ~`޻џjU�N���t�P��>G��B�>�����;'���{�r=��z�u#扄z�S���r����_����x���b� ������W����J��H���l;��L9vk#M�:7���<�!f�ĺ7<�E��צY%1�5'Vk��{?�c��ݟ��!� &)��ֈ�l����,�~Gc�4/�0�85��`kNc!yd@��?,��>�3�;���`���=���F%QPC[ngd_���DLGw����Lg�l�Z�L�x����D�c�����u�F���T\Yޠ�j�d�^6�����6>���1�1�b>[�\�9>!P�&.s�&d�y�cxN�x��
䨸����y"sĽY�f�r 3 �	�؄��������Qg��}��N�@���������+MR��gM�$�}�1B�
:�Q��M��')�As�F)�)��E�g�S#u������e��%�+k�Ȏ��m�W�Y3:��hz��V&�!\K�M�W�s�8`�4"�(��sF���l���s���G7}��ژ�M��鬼I���mq^���8�$L(��?K��:v�Bf�m�1YӍ�;��W�����[E���{�'3�0���T�m�[Z���z����kk(�����^h�EH��EB�V�`Hy�HA[�B�кS.~@K8��aTLHA�{��)?tg`�&-\��!FR�kv�f\xp2��E��M1�⬳n��:k����cn4mȊ�	u48%�ʀ��s�р*&�i����Iq=B�0&1X!�kh�Hq��u��o=��e��^$M v^��]Z��ԕ�b<Ʈ�?7�	siX����l5N63'�([g(��*��
^�T��xt�
�A�|��)8�̦a�MD]I8��
?����t�%&/�;o-�U(�{:�`r��uvv��r����# �1�����������|C���Jե��s�;�
H��\�;�{�WU���T�mmų��;���?�T�8i9H��
��,��Mg��к��fIZ��G�ܧK:Ј�
j٘�����@Qe�.�M�*�o�Xy�TcLO�<�'�ΥG� �L+�������:fS�"Χ`�n!�:�7�l�A.OJ�~�T��'9���9��xw��{�~<�=iJ|]'����iu�{��RCy��n'|���`��80vp@0��w�ྦ��'f|�+����q�-6�����}�iz	���l"��F��.�����r̎e��G�F¢v%y�F��+}V�.�~�ن��A�T��v��X��������(�
�B�Clr@������B�#��
'�.��� �`*����!׭|�l%/X[*� Jnй7,P�Jt_Q����kvÞ�OR�~����Jq���	� ����fu;�v��:LbGJ�m���3 �����&��Xo���9:�$��&��Y�g6^{Tw���j��s�s�����΀��q�������]��hd���9V�Z���ܐ�¯����A bY ����N����$�L�Fw3VR_)�7�yGo��\���8y��
��i�HW���:���p�̱�)*�s��.R���X�1���Џ�u�Vx��XR�T�ⳎYaQ�A35�@@��rm����B���,[��w�'`k{���,`뱡�l�7]���*S�C���>�K1���k�@���I�Kp�6�8����qp��τ�����#�!������&��:�����O��mȢbk�:�G}�]���
}K�F�ӹ!6�QfE1fFz4G�wfv`�S����/���u~��;�3��������` .^�H�0��o��ŵ�&����r{���m&����%�>�	3��^�r1�� ��NBg{{`>$Ǣ��v���"\r	�� �>I���+ަρLM��4]A�E��� �26���/>:�vu����Ɓ��Z#XӍi�A���a��3g�s�.�&�y����I��Ѭ8|~��o�C��Z ^x��s�O��ZD㨙T��:��OO�L��Ð�3Ư&6��b`�LP����k�#Rpg5� ��`���Ʋ��F'nb�jx���l�xc�8`;޿�a��s�X#u0�g�"������qsu�3�E���`6al�霻���λ �hr�.��[W�5YJ�03�j���Mgn���%}�7���Ʈ��6�����B�h�|�܋�V\�3��>�\������H��F��6P��8h���Ҵ�r�Շ.7����d�|>��U�{)���&Mn"����'Lv$�׻v�m���C0��Ah�b� CT��R���6���퀉�O�=hZ�nL ��� ��{�)�;�*�[��/�d�*3C�baIz!X��[ި�2���yd�rn�?g@�w���B�I=!_J��o�p��}��y���N���cQс���%��Y$�˦�l^G{��^��J�+=D��N��`]���B�n<h\�`�$m�W��XP��NR��
��0}����w_���D˭��A�4&p܊.�J�&Tv�*Wv��QD�K0Vq4w*��0!�pe8)�޿s7�N�	 ��6-��Ժ�r!	�����L+��= Q�ʆ����x_S�ퟗefz�[;�N��40h��@���)ӾH�=�H4�N�
^76Z<�R����;�փ�Jt�3��p�|?^��h�J�!
�:]����[p �u|��'��w!����	zr-�^���������0�no�QKM=�������#�k.s̷�Li0�
�e�
��˿��8��X+��&w\ �� ����u;��4SP�k
c�!1��hq��j���?������?�	 ��mg�Ft��N�_=��I�X�2x�.~��=�Շ�<����Y�ã�<\�mT��C��IʋT��I�XM7?�8F :���_~�c8��Юq��.V��9ܹb��"i<N��>�<}�,��hݙS���������ǟ���y�p�R��6k���_�"��'�-���2u�z�5�͉ƣ�?���o��Yٞ�vܙ���R[�7!Z��JY��O+��Rd���>�m@j,�)��������YSO���~I6E]���K����n����=�{t�9j�s�PO��pŵ��	t�pOCe6�;|��w)�ԁ�b�3,�Xf-�k]WY�]����|��'��'7?�u�L;	�,�'`�z�,�l7�I�nxQ Ϸ@t�P�F�Zp�1n�`O|�x��9���q*l狣����s���dW4��k��=�8�b�n$(�p�Ө���k�`�t�(>}�B��H�D��
c;�W�#ڈq���~���{.WG��,��֖�����cI��!�B��bnq�& ��.�|.}HV�?�`̏��%�CT� �`��1�m��� x�c�Hj�{��
t1�v�����T ��~����#� 4c�,0�ͤ�c�UT4�5	�6�b���19��A��G��{���5�������5�jܱ���D'܇d�M�W8#8��v?+kLbh�]�|���t�(nWƠ��D9�Ĥ����u���0(����E}���!��{{ f�t�Ni퍆��
!8�!���hSN�!G���)�XfV��[���~0�r�Ã���Sub��)5�ڰ��PBn�#!egc��@ g�5u��y/�ϦSi�赂�{������\�H�}@�Lȴ��2y�&�tX��,g�M����{��fw�lD��c�����o�Z���ϧ�d���I Ґ�_���
0N��(tS�����o����	 �M|T�R��|��n%��@0�@P�v������8M�sd��2'8h�1@�x����wN��{F>��>���v޳���\��N���x��k����.���@=gljt��Hz����%ŉ �_���G���{��0��7������Xj��x�/(���ѿ�`�dpXεx���g0�B��5�2+�*|gd�϶��:��,PDV *�$��56^Kp�/}��ΚVxo+�5�[�c/嚷n�Hv��?|�؄�����X`����m��#N[�ٙ�MG(��J�5vafW�|��ܩD�4k(�XW�m]����'�AM�u�	\F��R���`��zԬ��ɲb���k �����{��;�
�b��wc���G��)k���UJ���,'���;t:q� �"��l-��%�wxÀ�~\o�Y�:w��Js��=�(�d9�Ao�S4�agk�t���� Y�i�xsUuW,y����Ԧ90�e�Q�:jkԧ8[1��`Ml��p5c�eUѲ��0��@�'A�O~=W����G��lY����AyC�������G�zessX��Ь����n��e�֭e��fg_�=�{/�( ����j�:1�"<��֝6y���!�/��2|��W)���l��
�"��$�G��{��{6�l�X[�re����M-{H�����p���p��-&����:ۼ�lq��c����(.�GZ�_`,mw�q*N.��t���M���{��U�d�������s.�1�?p�)�@�\l��F�Q�X�P1P� D6e|�)t�(�ى�O�t�X�P�QG�ؑ&�\:&M:ԧ���BnQ윜����k�MP��4��s)�ʨ�պ�-d���uz�&�d��:N���N˚���u�C�
����g�X�֛2��Ŏukgk�\��}������ŵ��W�Qf9rq���ic��:n��]��(�<��<��_��?�'�
K�s��^XS3w��CR�j �HR0��Bɘ��d�)�v�!����Fz|��lH�\NY��Ł������ޮ���n�kS�ԙPng��~�9Z
b����c^r=E�)ɫW�uܶ؟�kh���a	���>"�s��6�\7�T�@ UTޔdU�u������gtC([��Q���6a|.��Q8���;�^E;S"�Z��3䓩 ���u�9�:t���ކ��Ī7�'�R�Fg
ذN�=�=װ�}�;��dV��u���h"w�L�i"`}nP�v�8R�����?�0��@FG��Zk�Ng,���9�Z&e��>(�H��k���O<$����1c��U���	M�(�}u��N� ���f�Kx����u�f�"n® Vz%�K}�Y,NNLttm#�_p&�Ǽ���_aLc�%��6�@?��	�N��(e2c��1F� �(*fGSλ/���D� ���9I��,_�#�Xtaz���VV�O���y��	�:&�͠[�]m�K���s�Q�~8�Xb6XnR[�?������ѵt�Q0.[q���VF(��f/Hk���+�\aD�N��߿�����lu�" �wuk sqYs����|���ĵ�|t���&��[�
���[՜�����#��xag#P(Z�Vf�S�R�*%�;鬸r�
u/]��r����(0H�����ޟg�\�����@���bP߱�x��y���t^���0װ#�.�p���'˳6S���W��� �(Z6�Cm�Z�F��M6�������l+J��$��Ⱥ6~Wwasc��d�ʓ*6CN�%' ӫ����
�P��+���4���?J�"+��aˡ��k��hڵ�=�qC����+{;�Nx���qZ{m�p�r{]��qF3���P�����(O���� ��>�<\��1B���l v-�̈�Ks�U�"d@ǁ*�K�������ԙՌ�� Z�L�n?ܿ� �|�^ڧ�(v��I9�)���uH����!v������7, �C� L*��s�&/@"<S�%�����yݙ�}ǵ��q�i��2�
�U�D�I�ǋ��S}�.9I"�G%e/2fV�9�����>G`+��|����J��Ϣ��Ϝe���o�:�\����9΁���!wCkm�2��	�4��5��G��/^<%����[���tSL�OZ�x6<qfjT�����Y�l�1@�@.�m��0ȣún��Q��I�uѠ�X7N�8|�b�р��wpşf�I��k3��(y%��7�xf��v�u�O�ٽ�{���`���5K�*�?}W������ᒋ�c��h{��Gr���YOج�� ���|�.���L_�u��,}.�߷77�lo��&��'ҡ�H��Y7����hM��g�U�t���Ά�5{S�v�`{�\��pSIO4�h�<>�s��E�j�XdN����N��4'H��ؼ��W��5Z�r<��DY�̥x�/Y{�#ZW7�OLGG:$�˖�;�D�W�����b����}$�X�|�0L������&贸��iY��"�^�C�6[-������Aܴ&�;�� v�(~ut�9W��qC�������}c̴�1�  ���9�a�$�[��k6�^� tZA)��҅�FU`9~��U.0t�C��b��A�ǡ����@�ƀ���Z��n�Ka�:��fm�<�%;.M��wG�������=i�=���ݗ�,�hq~�^`��O '���ߡ�^�
g���0R��?��ۣ2�8�3�t�L]�`��cm4��#�n����,*Ce�}M�f�*O�=�rJk���P�����)�-A=�|btE:,6�vz��Q�_~��聒��2H@p}LJM#I
�α�� ����_}�E�������]?$���k`M�L5������pȭ`m31�n߾�g_� ���S����N�y=�HQ������w��Q \8Q $x����	�΋W�4��`Q����UA���,����@��B8��9�d�c�7��8�?�d�yJN��  �o �
*<��F�/u��L<�"l����w��ƪ�����|d�D���Oe��fޝ�q������Ь
 ��*��h�^��px-�(�)v��Nh�K\�@��suX�%4��	=�s!�����`�*P�|�.N�6q�h�VcZv\�h,:JF[�d��iZ�p�����ZTӉ�IoJ��`�pp�S�
[nT�clޅ��U�@���AS'�����<:p����ņq�J<�MC6����� ��*c|�ƍ���8�\��t)�H�x������Tlh"�.���P����S~+W!3Ҭ�}Mzs�@9>{c}	+���Mcv�fUU��ra���@�>�u����J�ncr]������X"�y18��Z1� ��yZ�pm���y�>�7�Q�*6�H6�b��lt�2�3�� l��Kק�!GP/��A�7��<Nځ��'�s ׶gD�3��#�ib��  �tF�ӕtǬi-5���g���X�f�J�-- `��cl:X줨�w���ȒM Ct��0'2�O��۷nq�����h�Н%/M����Ӝ X7���|v�"��bX4DB("�c�%�rm3����i�� ��\����?"p�>4�H�M
�i| 7��;{ݭ��P�9�=�i F��_��}���dP�7fd{Pi ���m!*q�ͭ�Xj��=}��txļ�es��Yϑ'3E�-}JcQq=�9Q�zR��YQ��Y��&Ȑ�QE> &�y0v���I@T���M�@�Ȼ�  N�~��W�a2Ay��.��&㳮s���:���ٜ�g���O���ݬ�����+�a�!�O&��`�lo�u~��r:�ފ���(c<��.c������0W! �`u�P�X�M�e�t(c���Z-�2g���2��~~6�3cF�c�Qc3u�]|OƴU���ի7���kj�B�O��h��ep�(����r=4ё�m�+�7g�3A�M�����HO�NO�.�L�x��cW���C���lL���Z�A{�Õ@�rʛ֢d< �i�A2�ςNW���S�p|tB֍jT]��	���#��~ş���9u�yB
 ),Y�KwU��~=����N�0�H�5�l���cAMݹLNP�8�
b�]e�B:z9��h���ui��YC��;3!Å���ڑ,���!7K��.���y��=�{��
r��@��rC(��~�c��Sz��P���3�����5�@��Q���0��5��6��;��d�+���|�b������f�B��QЂ~��� Ux0P N4bd��e���6��`��ރS�ٮ�S56b�؜�Y����d�to��b�A�w��g86����ʦ.�d��M��sԩ���A���H 1�����S1C���%������@�����u2���Fr����B������I�~ݛ��V��p���Zvv7򼸺}�h�C>l��v}> �V����������:3�ϝ�ϗ�Z1A0��0�Ь�G�λ���GN�
��4�,�����{a(z�Ȣ`�T��gf騔=�Iw�,� Yg@�m�!���%o:djvy���D[r�pHI��ի��[��O?�% ���;��*[Pҥ�]�� �X�r�r����߄��nZ紉L{ɼ���V]75w�`�{eB�5�#10*H�?��9�5G&���H?�������3�E,{���s�
m��'���Ç����b�0Ia�%f���R���T�P�O�{G�=!��/\�.|x���H��� ��%&����5����o�l����ȭ��j�� txOGa��K<�8B��:ne,�;�V\�a(����Y�u�ً#���j�(�~�z����w�UvCgs����� �k
Sb���o�I�e����\6��T	�7ĜR�'�J?1[y��s�(}�V]MU��Q>�)�o,�{�
h�V����`�5�n�*6�.^����99б�<J����Qq��1��xש�я��s�W�ܽ��T�aa���T mI���ݹݦ`\�����.�k�}�����rɂ{@�����X`�"�=���ꕴM �,O��Z��+�����S��L�(��M�w�z����~7ҟ�^��mm��h�?��B�M<�H�Y��XϾ�{�Ů5!|b��J�]O�k$��i�r�F$�PQG��i���c�L���_�Ĝ������b'CJ^��X�5��W��E���6�(B6fݰ��6P\|���+٭,�}����H�o�"�`� @�Pe4���q� p=�[�T�b�Ah��B>+��_�R˒3�V��[F���A7E�O����W#q�\f@�5����@��n�����y�&�[[F�`���ܙL��'��;��8S���� ���h+���������W�.Y������+�:>Q�~�٧�ڵ�|=�Y���x�T��V[�Oj-	�
.�JЏB�1�����ݴ�`���ӛd�u��"��J�ϑ a(����1���k�}˜�gs�, *4G>l>4W�ʀ�Yxݦ�n2#�L�5��,x��a�" <೜/t^�ѓ�m��� �ь<�B�؃6:�� /��2ˎ��r����d��#s��O�S5���s�|�h�q��X�S��
�m��diF�Q̣��H���ycvh#C�X|.}v�	�r`�5���P@�9h�u3��^����)�e����~��Ԡ���F|لi�V�jb°�w��=hj���+8��|�B����!�z�[�G�i@B�g���  ��IDATʍ�`0�����aMS3�a�4�\4�Gc͘���Wtd�4ţ�/ Y��#`�k�Q��\H�T8ؤ��gS�3u`��<F�������;�̂|�ry�5���|l��އ�a2�����#� h�"g�4���[k�t�4b����N�8tV��	4�ɚ�Ʊ u(ο��3���T�Y$X��ڀK�Pud��5��u,�Ge%�HA��\�C��k��k�'Ɲ��K&$�/�� ��{C���g8[�?Z����8c��N���.F勫���;�Z�2�_��'	�9
�ot���Һ�	8 x���N��ƵJ�Ƃ�w�ч�2�ZT���-_@�/m2� ���D�t��Ȅ��4#�*��j�uiI�@7ݐ���@����k��x&:5�(A�w��!%p�NQ=`c��ʺ��F�	��R0
�>��D��a�N3�xo$�x��y�x�C&�;�����7�g^���ur�����0�(��:x���i�7�T�;<�C�ݞ�ߓVB�`ڸ��������C���/(��)-P��u�@ 	X��0��*�fxg�1��8Fo�C��T�]R����QD+��C���v�"��{&�{:gi���,K��1@'����]KV�"X1�EW�8H`�y��������.֠��9�S�J�{�#>��фp���sr�쉰�F��ĺXs�Z�6
X�� �������(�щ�l&\�g\�-^�l�Yo�u�8���A�qB�H�I?��P���D�7hS=e�G
�Y�"�<�w��;�M4�<cH�N�J};����-�e �`]��>:�Y����Ȁ�Jr�������M��̳�s�2���g�q@x,���:��}0�@l�*��镹(H�Kc.�@4X����AW���;�d�(��Òd1��3ӪSƂ����D�)@jL+&N&x�C�"#��F��c���]3���.Cً�_][�7�2v^c�T����C��7u*�/Z�2��bc�u�ٟ�@��Dv�ں���c����F��ܹA<G�-�h��͙�O�%5-���X�1�#�R*	�C�:!��551E��^�v=ŉMc���dH1&�Kb��b-, ��bS1i3����j,���a��̑�hnl�>wDsܷ��h{%�2Ð�6Ē<�;��{�>�+v��i�L�#*�l�J�O��kD1J��:��@ �w����r����f�������5���3Ƙt!�
�ւw�Y����7��aLQk���g�7K0�_������J2��������g�}��C�Ύ�cM���л�b�T�aTb�8���k2��H/~F��ݎ@ �mn�0�y��<E�į=�TI�uG7�������#��2��A �!j��m��rc����=����X�l/;А����J^{M�7r��qb��z��-�dU��u�~ :��/
�/]&�l/���s=�s}�L3	�+�V|*���ӫׯ�?~O��k4��>ԖG׍<��z�O�*��ŵ�x�14!Vςm1'{�?���n޸n޼�}�q�t�jvU��%J:|�mkKa=f�"���	�$�3���(�S'�ga.q�[�!�LpD��T�7ر�O�+b�=�;�	\?t� Za�l�	�%wдV�LE�" ߵ�
��}��?7͌��ŋ����P��zz�b\a�h"be��׫��m��8�
Vo��j�:�}nl����ĵ���>��{S�(&�+<������2/W��Zm�/��^N��>:�[N���xN �>y����b�����9^?kʠ���S�YM	���w.}�������kt|�c��m5y���@Si�6��e�����G4��U����}�i��5�C+9�1�XA�{c�a�y�*o����欘h�m4�����"�����{w�k$�� x51֌[�:]���9�6�ȷ�����Z����Y��(��|bjgb��o���w�,�%����1c�`�]��cę����Un�8Kg�N�\�R\�B �-yL��\Go������"���b1=�y����Ga�	���
4v�T��
��?�"T�.�W����r�*�<��>9eg6�6R������Z;�YIH=)cwMTPJ,^R�
F�����ߍ5x[��v������t:�h��Ն��r|tx�`/_>g����ǟ�~s�R=Z���ӵ*�{9{J#?MN$�L�E&<���(4)��
_�����Tb����Z@<m��tƫ(`G��cA�� �1[e
`>hI � ��7␹)���f*W��%��~��.�*[��D6�1v�*�����aj.3�ow䵷�&�����R��}�U]��?�	��f�e�G�=e����<��ƻ�|��)H�6s:f�x��G���g6:�c]��V��U�F$H��>{��|?ܾ�3Y2�.u��Y�󏎣�CO0y]�v[��ܕt���ƙ�yO��n"��V`8#͋����E!�J#(rn~rS"��g82ő�&k���9��� �f�� �z��M�l�J%xkֻ<�6l?L�0�v`I#�X�oQ���T��
O�&��c��c�5:�>B����=S���*u�h_���G����-Tg�*�ޞ)(�u���w�@��Q��M�\���"1�>
'������8���ó�&o�����T�����RO%�x\�dm93s������������;�ZX��*r�8әf����Ӵs�QطNߟ���ׯ�)���!���� rgԠ�C������{�G1���\�V%�u�f.�Vz8���[+4}�����2Nհ�f�/�5���V*N.%X�9M�ؾ�}:��%L�|�mg7H����-�� u<Aw��cM�(^��0fn3��ξB�� 1cH�̗���8o�J��_����no�����x�i���K��^$ǞT��\rl�i*T<zH_��_�b^�}���X���U�k,�O?��
�)�wN7@�G��WםYÖЎA���~�	8D.�d��Ȕ��������.Y��"^b\SkL��rl�*��8��͟�'���ȭ�X���X�,��:��z��*6.�B��#�=kCu�+3�蘣��{�'�>�i�qvΟ�v��4��:�Pp65
?��y(FU����5��n[�G�y~TU�]�$Z</�h�umE��;
�I�++��O�U�&ߗ_}I= �l���!��BL3�,�������+�a�0F�x�,����������L�Kr�4��9<�ńEU+1���3���sè�Q�&�5CJ��l��P��4$7Ф�rMB�"Pks��(�V�%�&�j�j��-�"q>��`#��Iޤ����/�ʼ}�6�͡EI1�JL��td��]b}�VK����'8��\ZZ����K�x���p������P`M΍!��^�)����`����͂��tAȳlؑ���8����3�i��Q7�i3ӭi]��C�ޘ��֎"r&^r�{-h�����@���~w �T�s�)]�H�g0&&����F\�}�Ku��$~/��d*����[����и����TKf`ƚf���G�F6��&�>�M�iTd���J��]���n����9W�:�߽��Y��U��sJzE�� :@�#V�� h�r�����W8�;_l�؂O\�������J��9�Թ	7��#hA��y3�+P���?O���B�
M�c;��q;҂����:Ľ ���b.�J�У�:��8Z]։ɵ6�W�~�J~}��u�h\�3薋n����Z�.+�LQ/ȿ�� �R�:\D�|t]���T�7��V"UA�8��<�������(*�_��Dw������A݄�Jj���"q��[��-x�y7=�����]k	������@���P`p�3��0�Pr�U.l=�Ml�}��m�ޢ@��:���',*���
���;b�{���&�5�T(��1;[r)������^�M�!� ���� ��o�s�|�@�[>�I{���6���Z�r�rk�a��Ӈ�a��Tt���@�^ۨ3F&� �eu����~��|��rӜ�ł��5��,��ҙ�X��c:�3����?���U����
��)'���$*�z��.��W0�k��>z��Y`�4X��x]fp���ti�TF̠�	�5Ǳ���΄�x([����A�_�?��ԫ��%��k�k��k�ǘ�N�1}($���rד��.(Dd�����)U~��%啔�޺+F�v�s-�rV�9F�m���իEG�[�	�Y{�N.��+����f���N�H��b��֢)���6G.�!���8���\�@�
8�@��)bFk.5��D�<���q��E��������R�]8+m.��O?FN�uP��!�X]!sE1���J� ����2P�5F�A�;g@d�O�>���M�	 ���>ҳ�:����~�ڊ�&�z�F:8 �sU �(aG%a9t�m�������!�����b���In(:��m�?�]� \~�%�)�G����"=�8��n�mҍ��` �Ԋ��ݺ��?�W�E��@�Q��7f݌kA�G�����B��_�O�%�:Ӕ�&ڱ���c�
�W���{�h�-u9l��
g-�*8^��H�j�M�C���GKJ� 	g��(��,q�e0}��ETQEQ��D�^�BC��u���3t�r߹��2�@݆P L�����&R���AG�,НmK�:%�p���_��>{J]\�Fス��GjLXA��-t�\\Jk�1�t�!�-�mi!!�F,#�0�u��kM�۬ݖWl;1*}d�G�xs�|�m��[s������7R����.�׿�:\��f�>/O4�BPg������
/���xi������&mp�I����ƽ@�?��-�,�}.L���8��Q�^���tML�b������a�q=��@Â�w9�Gl��-
@4�ޔ#��xg� �[.��ш��O���P��t_��?�m�ȫx-�dqZ��	 f����P/^�����'����9������#���?�ه��w_���K{��?�5W红�ל�gw�HC
g7� �r�>W3����Gp�ĸό]�{�� �����lggKL�ޝz
�2�`��K16 Lc�1߄�Ã��O?�
wnߦ��~���gб�ؖ��Cx�cxM��a����k�VZ���FU`>rO󈵊?7�������t���}�fݳg�	��yHΛ5�ʆQ�qr��Vy<�܌u�ʸ��9+�u�b,`��
j �Z�̀;Q���눎?�f�x)K�֜N���Z�ni�i%p4�L��c{��Y�����ȷ����.}��ھ��X���Њށr�T�M#�ğp�����c�o׼��q��u�\ۮ�s2�.mw|�<T�}T���fq޺vg���������ȕb S0�	��s?-�쒇&jl=|�<}�)�;�m�u�ȌI9��+֘O�A�2�}h�&�1�Z��jTb��8z���頊1v9����k�s8\oU��g^ͼ��pi���t�d˾��5|6lV���8~�֧���Q����脃���1cnp�`�}���k�i��g�1�܋�\��Ÿ�T�'��on����9k*me]��o��]�r%���Y�P
���KϷ���]pfh��ktF���+��s�3�Y硝(��]��3�l������w�ȃ��%�6ϝ?��l�h�R���š�9�j�`�`�	�!���r�� &�Q�t���ȫI����XK��,�0�zͤ
�(�� �@aڊ���Ք��C����̨�_Q4�1
�Y
�d�5>t@Vp�X���Wژ����i�7�}M8������U��UwE�ϊ�����Dgō�;y�Y���l(�0�eok��8xU��b:�D��[��@�s��,���Yn4��ֲ d0�R4�.�٬'����8@����z��S_�C��i셽T���%اO����'&���ȓ���u)<;J(�Tͬ��#�=�3���N��g�]�QAF7�nt�W���h���
Te��a&׎�R;i�L��E4cM����4�qE���C|�$�GI�)�Mm�/HoO�b��0`�l?���&��:�Ē�������Z�x�x���^w<�V"�8���[��E+$sXu��biU���i�
��Z���C����?�Fǰ(G��q(Ǫ8:�*K��L&�ߧS����Z�ɰ|��%��_\�0%d �[s4������W��" c���4�	�A����
�ajv��^S""�ů� �Kj���$�c&��{�����u���������~�gn]3&5��� v���խ}Vdo
s06���rz�1$L`�=F�7��ڪ�c�I.d0�9���DA�"�hD��[��|2��>9>����[�j*t?�~��$��|��0�W�^��u�5dN����X���	52V��e��ǁ0؈�6B�Imh4�i����`�ap]�*���d��㪰|�(n�=��6w;c~�X����p�0���BwF��+2��~~#v�����lʜ�J���� ���dfg��n�=��%�y�]c�������O���&�]�F=�����7�n�-��11G\À�D#��0J�A�Z�8�_�x��K9����O䩙���>�<��+[CU��S˸Q���0)�@c�u�o]�l�|�u�ad@�)
�����ϥk;i�Y���YMca��@s*��Co9�;��ua*D�(f��}�#�l"!����F���UC5�Wp �cs��1���̎��m�1t+'c��.g/M����t�pV߲�A/�ncW8�&^Z��@ƺ}h��������?�<}~�{���I+�'��.�N���@���Ԋ�<H��]E�X&`ƃ��4�! $`"�����&h�p����~q?�}I��㣔7s� ���ݻOGxR��D�4��9�D ˆ�"�~6k4�1��ZSv"�`H�� ���7:����}payI�j�����`�2�� . �˗.�>P#7`�Trs���*,�:k�8�^b`aŚ�f0��N�V�J7�f��.pGgꈁ�(���^�ؕ�5p�� Y�]�s&}B�mF9��&��bE"��y����-v�r��{!� ��AӱR�ݍ�kb l#��<b�Jgf�X���Y���75�+��`cZ�6�q��ǽ|4ɝ�&����������Dg �u������	�zh<{���r����S�5_�p�҈u�.�a.|�NS��T���D�L��}�ѣ���b��sM���3]�s���i��{n]F��\ʵK,"���6�4H5Dkg�@���{f͙Y{]�i`���2M���C��m;
L���W�q��k6��,1�d\����X@���ʠи������B��c>�J�Oe�d���\u^o��Y:s�'��ZBW&�zbs����� �� p>���&Mc.�r:@6�N���6�^�ۜ�墅�Q�||���Q��v :���o6:6	�s+�J!z����iS���Da��C�H�m~/���atϋ�G�̤[�d��.
�l�S�V@��!�M���� m��P��I$�@����a��!�!X��AT���˩k�PĜC����Ո���a\+q(�P�r���N-A7g�z*�I��g��D��<kiKH4ٙ/��q�qF�\Ǧ��0�B׵M��W����r1a�=��w����<��^��5=ִ�\�(�Z]n����4�5�@0�D�l���S�r�C�6&���ۃÔ��Gd��S��%0��O��Y~�־��d+�;�慉��RV<D�<��D^2x}��/��������-F�𺃋����)	��Y X�����`{��XВʣXkv �A��+��2��^K��b�ݰ�� |����+1@���L�1m���F��F{֣(�)p�D6��~HM�W���k��u��̕k�=�{�8:���Q����k5x��b$e�hY5�n7�Y�3q��M�����|_�ʺ1XQ;ȑ�Ҟqg��6�
`����\.�0���m&�OSa�bW�:Z��h;�E�Dq�	�n&�(n������.���`��G5��j��;2>�^�i�(p+��/O�ƂH�E������yv�p���cw�a���͝�9G��rf�U�\�OT�E^[���qF�L�FӾY��ɖ
������{׋�
] ;X_x?�?�o�X'ƥ l{��皣��8 \�& {��z�>��o8��B�_ 0)z���\���^5�}��f��r�d�
p�)�!��5F�۱.]v�¹�6�,��L��P���/9�UE'��Fl(��>V��ggnm>N)v@\CDb�G6��u��`�����>��?β�F�hT�߻F��������駟�c��D�?~�, �%�&��,wg.  x\�D�f����j�d��C0#�˩��1�b(
��xΑw���l^�\�s�k���0��������k?��\���+xM|���`�OY87vvx~��ѓ���ΐ;��0�WJCj����~��{?�u!����ʕ�dD�������� 'H���-�O�]�gWg�`:3U)�m���wü�*c�XWІ�����,k����+tX��"������N3A�@�4kg�8v³�1���^�&�wxp�u��#�F���uƟh�{wu�Mq{k��\ ��M1F��!w�QH��8�� ��jЫqw�A�<��@�ٳ'l��mqfg���ۙH�1�av�SjsB�LK��W�H�}��L�G���9�s�:T̹�׫	5e�{��5�d�>�þ�{��ݗ�3��ކ���1���׮^���-��7'A���.Q�k���pz��t�{龿�{�9�u���V�*�$������<C����X�.>��\�F���>ا���J�ֵ;W�~�&� .�]�,f��g���NN@�v3��3�p߆^q��� �^�Fg�#޾%`@�޽����������9U�X.�'�U �Ș��n���`S�7�ujy����� [��1�ΛZ���V�3�љ���c��3pl-�C,NXc6P0�7o�XV�T��O�U��e�<�X{� ��\Y�C]�?q�o�l����W�$Ǒ%�!2�Dk�� ���>�|�����w�vw�!	�j�%R��~��G5A�����t��*E���ٱc��u�oՔ��q�u ��|v��5{Y�"!1]oN�߷́nc4��j�����c��!8�`�q�j[�v���n2ƨ��L�_tXs�`/��Z��rg��N�����@�Ů+O�_6n kUM�"L�{$)5G7�]>v9�A�:K�k6Xf^�]SY\��^���Z<�
0TG�~��p��sC���7��04JU�����,甦E,���['Q��J�ztR�l%�5���w�ݕM�G�qC	��ra��D�^�ʚ1��v�a��6�5�n]pk<J�a�͋�O����R�߈���A9:�1�x�^u��L�=z����6,��E�戛�Դ��c/�G&gR�G�����,p�����#�AW A�K&���X���J&K�qQ��(P�xu .�u�b�����\@��Zai�n�<+!���ԑ�z� �
j�H�&F�|*crG���]�!�Z�*-Ɓ��^�s�b#�~t)��;���f���S�ή� �����W�с���
���`
���<u Q1��|ExMb�B�1k�����D�)��$�~��-,���*��h��z��v wP�q_Z�Q�ܜr��\�E�4�* %Du�nֶ
��Ӧ��=s?����;''
�b@��Qy�q�J����Q��-��Y��N$���-VN�Ç�PXX7K���!F����6����]*����Y�a�[�(T�W�hG1������"}�z�k�Z'������j���J��@�}X���G�&�4�$K+��z���;}��z��@�Ya#?���}E|A����/�s���8�Ύ�crP�9Oo�`|E�+1v���B����\h[kb��et,3�S����|�q ��G�@��|0@��=�^U�9~ɟ������>]gQu��7o�Y���w�}�*@�����$�(�)��iԾ΅GU��c7�*C�Db�w��0���9boG�;lJ��']c�
1�/_���D�_~�Eq�I}$]:�!Z3t�����RW��T����W���bl�06�0�z����Y�����AB=GS�u���}���:�Sq=a��t�N��Um(L5���������K�/�Φq�U��n]_������YoP+��/��^��<
��b����t�� ݫ7̧��9(F�t��A/ob�����e{i���G	��d�=zL�γ�.љݙ�C�jw�Q8�6<4>����7���'�!]��V�����\yL�L������	��'b�XSB��]	{
�����Q���������Mw��&k�q���r?��R��ma����VE��gb4���v�m��Z�,Y�}XD��/���Y�<-��9�q��3�ëu�+kmf�*�;�	7�k�������<�f-&��@<}�٧髯�d�k�<�Hl��%WD��y�u�2"Xv(�p��/�Fr��e�g�S�!m�߼f���6@6�<v*@}��5:�Ƚ�`P�������4l�w5��@m|F�]hq�{u�L9f6��� �	�o�_��޾}n�Y��lP����q? 3�6/��&7��q����eF�@�;{���i�˓�<1N��@\�0刟_2u�ASc��� v=s�N��j�NԷY���\���_�:�mw�cE]�=���(�lJ��e0�'70�g�W���2מ��Ha���wyq����c�)`q��9|�9��$ٺ��\7��es쀃�����)�
:#����#�pٸ?�����z�m�.�T��~�$�������y	�đ�]*�q�F�$%���d��Y��4�Ju�4{<��� t��� �����S	�I��:�c4�?����;6�7�c]�uεo��zF]+ǵ#�{Ks�Nk&��Q����U��S��C�3W�}a�B��y��`R@4ї��'"g��i��4Y#Ǎ���g<�R�|��Чi?S*��競��z�Bsr����S��X�L4��_���Q�����b���.W��H����f�QxF����=¨�;s�4iv�:�bq�����N�dB�~���d��(pR�(��N\(u#��X,��4�'��n�.���i�����P����uFQ�3���%��O�!�$��m
��@j�Ti� J[���Ѝ\����wR�m`�L���0=%��z�.v�p�)��;$�'�ItyP@F;I�68¨���豓�����ݏ�`�/F�\p6а#�Kly�V0�����I�c��XWr��d��e6W\/l�yrlL�������y^>�u]�@Ɠ_k�膮��̩w|�*�f����i R�#�t���gm�Z������(�X:�j�H ����}8�k	� ���l堫b�z ���RM�#Z|߽��޿��kL������O�=�&v�|W���>O+�Yt�N�L<��;�Iv�ȲP�������#�IrIc�t���}pb=�Ϟ|�f��Vkw�.��[g����w`B� CRH�_�;����Me$֓5�����5����g���vI(l���"� ���Q�����~�p���2y X�o�-l��⡍�O�ߠ����,�YgA��_���H\aB��k$q�(��h�@���j�q��[�~6�l5�xl�$1.��ˁ��}ۄ�1���ø�� &�I3o�z�˸�YMx-tq�F���c�����5���}`�������Ho��E؃J�Q�U��(A����Ћ� �m���%�;��yf�늅�З��J$-HV�
�1_��-��{��ӓ�<3��Y�I�I9�P��Ι�8��b�1��8�Vlۧ� ���z��W ��5iJ>�E �x6���W�<��� q�/�|����B �Q��b?�����|���l��� @���w��k.�r*� ٲ�a1r�)N-���Ǒ��H��)�Wa���\8�, ���\��W�G�Is�4wX��3���vl�!���Ζ6���#��b?5<n��������S�-�s �׮�`����4�O�b.9C��E��f%��>[<��!\o������^�������S�92��
� ��w����'���)�� ���}�H�e��8F����(�4�sM�5׍�G�6�q8��@� ��t�!���;�;?��p.����9~�B�9���َE����C?J`ջ"��3���5~V��!v#6�Z�ۿ�k���/0%�h��y�;�=��;�����#}�g,���9�ٙ�G��߸��I�o���gX�)�.�2����lht��rJ��sJ ����~�G��֌�S ��0<�X;p,�c^Z-�p�2�,d>�#��%�kv��I��؏5v��K7��:�:�`1�IV���x��uL�뙌<�'^�j�<�X,�`BG�mE�l.�B����Pqޢ	4�֚�Q�L�W�-Ν�2�V�a�b1�kW�v��&���Vxb,�,%5��mx����X��`aD#�hй�P��^Ec�י_`�@�{������"Hx$���
cg] ��bz$�\���/�ZE4�˅��!� M����m��P��n������߃�
�K�a��K�j>�v��?+�
	�;n"�b�����'e�n}�$�F�@�V�F�yJ�ۜ��&yN�(ĩ�����ݟY��9E/�m+P�G!�z"��|3��'�0W܍��P���ز��Bd:4i�p��g+����:�2�/��i^<Oԣ)�ço�\�y�U;5�"���SU`��������)�C3�.�O�ұb�;֎A�P��Ma�G�O�u��#�z��၍�@��?� pǡ3z'*ޜ� �RS,^�!
i):x��8EM�u�Y�P�����xtisп�����{��@�|A��I����,����	���>���)Ic���n0���r?���0�Z��+8�Q�}:�9��A��Iʫۯx�oV�R����ǿ��ݴ�}�ً7M��� ��DB�a�CQ>��X����}Y� f���Ek�uH�NLbI�m/��T�]�U=�.Pb*���)P7�\�R��;5�	T�i|3�9Ж����5
��l��.<���;�T�P���VfBE�C�M�UӔ3��ޯ����qNf�2?}�"�k9:� &����.�^o�ں�]0��ꬷ�[��/ؤ����uL���E4��ׯS�d5�ƅ���Lr��������M�:��MY���_���8`1�%G�#1�R*�8$��X3EzYX����M�D ��;xHi[n��6 ��
�\ө3�����Qq����Wii	�`:������vXg}��_rO:�"�΀pq��/��\�I{R4� w�ӥf�����w��Mei����"\�:Ql	|�>��߹�	z@t������sq*8ոHiڈ�և���8�}jkқ���F���aC�B����E9���,`0�1xg�`�v����X��?J�����ك�V$FЌ�[�D��=�on�N7_]��l�S�޺��xнQ|��'k��*[g��,Xv��uh�(X�&gd���<��)�,N�y�� ��j�����1{!���LT���嬊�V�f�Ĭd^@W�i�͊�!�]]��A�]���yf��K�l9&��qЮ5�����읺	j����>��m���յ_�A���TovL���������d+��(]�Hn��FZ;���̢�f�Q�I as����w�����d���oq\:$�oĠw�>b�kt��v�J���(��8F5���J�SX{ ���m0&P	�iy�#��~�5���`C������~@���&\���s��@���\��F��ĳ��h_M^�u���k>@�>�� 3KҀm��C����> ��������b�8G�������z��t�x�B�~D{�,�Ѐ#�Xou�eMG��&�ٳ8b�p*@�o�Xc�q�
�fb���Dk7������#����p�����?����'�|̂j��,�tp�>MM������F�e��ۙ~���!����p�">�ݝ��`P_���
k��D&�m���=}*}���$�;Lr���Yo&3Ɓz�_�7l�|Q\�g؎�?Aβ9��m�Ċ� P�׮���������F���'����ೳ������5ĞC� ���_j����8��s����Yȕ����x��)�����:n�h9�i=c����������F�{"��r ȫ^�����?}��L@×|���E:iOR���� 1�9�z��(o ;G��XK�1��J�����?R��g�'�)@�wO�l���{tyt�_���J7���gH������r$�u�`�bM͓�Q�6ڇ8��ܺŽ��p�F�GCL2Ć�͸8�4:�:Eq:�M��z�:����qp��c��<��9X敱�3_���F)�fw�h*��6��'/]�x&����	@�jΙRe��_������p�Ls4[k�Q��W������Z�4�ͥ�X�jM;�W���C*��kE�oWI c���_y��JwwQ���d1K����¤7�.ǅ���f�0h=G$ ⥸(�5r�7�)7�n4j�H~8+l��������F�MfH�M��9�
�6X��p8��yK�'�#7V�� �u����U�䤃��ng$JEC��U�S���9��	�5R�5������QP�=A��y,M:3���q�h�ѱ���xj�tBoЏ��.�i��R�;�	62
noN2bWi12Ř���@�)ܯ�9��(�T<�� B�1�.�a��	Qnч[�)1>2/\N
R�) �x�.(x)['JM� ��Ȃ�z_�f<���uz|z���\�?�������:#"�"�d^�=I���@���Һ��6���9u^R��9;��
�0t��(��i��ۍ�K19��>XT��r���.��;�\�F�O<m5�y-J2Gv�xࡳm�)��G�·��Ĵ�}tox4�`�F��Q� ���� �n] ��XpС�{��$$��n��gY�%�3(�	�p�U'�m���@��)�p�n���[%�p�@�qs0�����8x�������?IȺ�⌮.># ��FH���@G/J���QTV�sv�),_��bךs�1B�buN���$�
6t�h"[���Q��u� C��B��7Gq��ky���<��a�q�f�`�\�����u;''(R�N�)�Z��ޞ��kѧ�z[j0Ղ���}�����h�o���Dn�_�{�?Ud������n�S�3�W���V��Z.�Q�Z�3���9f~�}Ñ1����H��Ɉ���L��d��`k�1FqсG���Ï8bf����g4�&�A۳�6SF�@�L����/	XJ���0�	_���θ�zXH�$^8��ڦ��H�2�:>�ՒJc%��И��y�2���x�S�v}�9C�9��,?z��Z�%wH�����N���JS
�C�#�bJ%\I���>2ƹF��`g��6�z��Ν+���^��,6	�T^�X��M��:��7к�zE�A�A�n�����Oә�W��BW`	t�4�YtJqN���e#� �tL����D���+��r����O�'�~L@�~���X��L'vj��/�;����Y}4B��_�[+	Lms86	��c���_�7#�9���xc:�u��L��ϿO?渍b�Y&��t�E�k�S��h���p�8
6��h8���B>w����`�:��t�(*�x����uދ��m(�a\�;w�2��Y4n� ��zX/`B��b�4��1.����?��u����/?I���W�-��\�OOS)J���g�v�����Q^38��&B��'X�ȝ�d��bm�k���[����n\8���oK�@��* �1��o��G�������t�$�RC�ުsNL �\���1�����Ȱ@g��'�;���H@y\#�r��:��L�8Q�Y�3h*�%��m��K�ދ�/�#ݿ�!o7���ȧ5�E�q�ʬ	gM�_=�ܤ����Kq�m�W��%h���D��F��ADc��U�i�s_��L  �7���_�q}���=��7t]�qض�c9�X�H}�q����������{�Gl�s1�Ț��]6�g]�Msm ��m
� C�YHVcc�E�{��L/hp��>���B�Z��0q^]9>����kځ{�"?'r�B�m@���f������ �9�5��S�N�b~��oh�~B�{2'�o1�yP�������|��uϯ��ِk	\�7d�][]��тΜ9t�����3�iLx��i��c�m����"���9�Bm��_�:n�_���7�Bn�'{/�qYY:M�rc3������w���_�����d�X<��̿�:Է6��>��
����f.ݴH��3	���6:G%@�D���O?���
8�qS� ���^ �a%�",B����|t��k�U�(XE��0)��s�Bs���0�$,2��P"'/,6te!���2D�n�L�{w�d@q����}�Z��f�y��X��o��5U<�Ӂ��MN�1�N��/5߰*fb���b̀�����uQ���k;&ƻ����Q����Z#�xu�އ����V�����д�@�Պ�`���i�h�v0:jP
'Q��,�*��������}0��O=^t�D57��7A���ݴ�;N�#�7�	�<�L�m9Y����W�,*������hWFњ�������kvGn���Ը��5��uT_��t��k)4o�=��<w��ұjRhS`}3��&�H,y(�LHG�z�Q$U$��x�Qks{М+b �~��t�4[�� 3$F���+�ښ	H��%��<��׎(�>4|�7t?8%��G�S�tb�j]�5�5��9M1��X�w��{ �3����=�t�
�4K��1:� �~��Y����Mw���A�:.Ƕ���s2��3�����d �Ф#>NsM[:Z4ӛw���,:)p��Np�?�Ҩh�:?�>����ļ{�:mrA�	�p��]_�?^/ �օ2��6ş`��܈���Mek��aWJ���\(`�Æ� �l���(�7�|�,|i�I"��u���<t�
�HH��r�ܵ�'�N���b�!kQT{����e]S�����^�� ����g(p�ڲYr,��߽����Ea������ qX,I֬�i��"�~�0�Y������� ���A@�qlr�O v ؘ��u7 7!�0��s�=�Q��V8���ȉŀ�P�u,N���6�E�d��Խ2z$�ۃ�g4��x�H�t>ĹS�:�e�$s*$Ώ�b�j��[0�Xh.�~� ,+ $�������X?�Q���Ya�K��c 7@�[���[���"-�(k�E�C�9�BĜ�e;��Eq���8�x�:�G�������0}%7B��Y�h<G.]���ϩ�IJ��t�|iOx�Q��+�#��MZ
1�z4�џ����!�k��s�j�߰Y��߾�Jsd�[�|I��)s^w�؉u�:��i5V`��8��i.J�O]�y���t��M*�#raivI�c��4CCo?�E��) �_!�h�`�gZ�u����7��z���4_?|�sr�^#k��.&�
/5j��+�K�X� �����Q
ݘ�{��>���d�;�ȉ��,����hV�D#z�l �52P�vJL+�Tr�Ɵ��|ê�z_�CΛf�iCc�b7`�{���{ͣو_o�bYķw�?�@:�X3�'g���'�?��(��3���g�`��Ch��WٹZSSaKIt{���9�y�)�'�[��̩�[�x�"��|/�6#c�C5&��]�]�"n�pC-�M���F���%6��t�� ����6w��p��-�\��ɂ�{d�@����hn�Ne����J��%KP�,�F6X5�2����X�O����>�E�c��WP�j��ћ�a[��o0G�/P'�~�*��k��-�E"����g�:C���u�o�W?�赅u5X�;�S2晇8dW�f�ή����]�w�]0��I�����у1�{��|=��:�ٯ�9���=	b���1��b�˲s82�����\�W�=����W�?���q�\��_}���gt�+��!�{+9�/����M,��P����jMэq����Q���L���k!��j��d;�2?>Ao��;���s�^���OX���D��J�95�y�p+a��:�*l��c�TЅ��q���+smm$�^h��3��ߓ����A=>!��x#}����"a��_IS�3J���Ɋw����ˇ:t::�(`BT�ꖴ�K��k�7����.�؛��x�4���Z�zM�
nwe��]��9޳��.S*t߶?w�:Q#@��aI+N,r�P��+xTRt�������<-��J��f���?��Y씲A�W�i(�-���J�Kw&�+쬵������e�2L��:��m#����pG��e� IŴ���׀ң�1��ݙ��M��La�(M��UqI׏A�(A�\P@�ᆭ\I��f�$,`�}��ǥ[���7���\�ޓ����\оGWo��A�x����-4v��m���v�1[��s��6�k h�u"c�����'�e�]M`�p�" ���/����Ɯ��??�p5�(�S ��8t�;��e���}41��}�$�Ȯ?XJ���M̽�(n�V�3��(��1��k�5r<6�}���2�[:EG����	Y8���I��,�wfK�<P���\�9G!�X�����d�E����0��Z�� &��z�w�5F>��s&(G,.�(Q���<�>�W�B��%���\�I�}K�"�0�'!$��t?���|6&O�����?�������2]rm`L��x�d*��qh��vLB�.,�`p�2x�0���E��j���+mL���zt�w@�Ga�kG=�|/6�q��ANf75Q����s2��-$�E�#����^�B��6�Ux���,HUxpY ��=���Mv�x^�Dy6���xlq������Èx -���oݝ��O�p��B�P��Nn\��1F�C�	����* �掺�o��~����d�1o��&  0V��y_��wy���s�����x�q/Y�:���̃�#�\�ދYLj��gw�;j	�OY��F
�B�p�n��C8h<�*�fj��k�� ����e������gU�`8�e�:�B��������i�[E��1����0�fz�Am�˃G�4��c �#�Ga�CL9X/�Ҩ/r * ֐�!��<��y�I�?���5S�(�
� �)�|����r��Z8��Qx��bTpr���g!σ�����/_�,b�O0E�~`m���ϋ�Z��jR��|�����5O�5��jı4j�����jZ�����7�r�`&�~� ����3
��c�{	��mo���t@ژ}W�1�n���i��*�����G0�,�G91A���TB��3�c�hy��v�t��9H`pqvE+�񼷠Ń�
�!��ͻ���"7�8�X4�K�_��y���7�� γ�^�O���>��b-���s'k�H�e���XF�8"L�g��9��{�1�Gё����k�6��Z/�1�4/s�TL\�"�9kt�y�$+x4O������_�W/ߐ)%��L��=��o4���!yrzL�9,@�?�(�Zh�Fk8�^aG�/H��l��-�<���cL�0p�<��:Uh,}��ߗt�"7҅�����$`w��ĨP�k:
��w���?N��O�Oҝ{w���_gc�B N�H�������۷{"�N�8�{F��ZzCZJKp�����L�zt$N�Cp�:9@[&-f�&�j����;V�i�:+��I۸N�Y�u�sAvҁ�>�B.����D�'���p��wv�k��/~�cdmk���bDU~�n��5��v�͵���k� D�o�G7=_ڴ��>o&5KFKtcS*�+��\s!r�0W�4#�^��`���g�`$Yhz|���tz��TD$�����.����*
���;������Aq���4r��j�Q*Z3�0mqH��=�4���MT����q	�l����>����T��(e�e�a	QX�b�
,"�[��-��B�jԭi3|LJ-ӝt�t, ��p���6�zʉ{�_h.2�}��bʋb�ә�2��$�(�C8�-o�S�ʚ��Ik�5�5�����*��o2@�&㊀�jD��s�Vb< ��҃0�����V`��+Z;���o�S-�Ò��� Q�)� �����@�G�>���H��5�u���q��b�>�(���<���8!��J8 ���5����I]�a�Kw�\�9��$�3��<�T�����T�y
'����ҡ7`J:o~e��ҳ�$�{�]<o~�,�f��`a@u�c@�j�8z}z��ψ�t(~����Wo�#9��:tL�oa119���i���JL��\�p��$�'��z]:PF��v.�zwt:�F�������.Qi�,2�`W�_������)�ʻ�����]<;�u��a�Hݑ;������"nA���ÇY�⁎]Ű�! ai���M�����,� s� ���s�~�믿��:��B!HЩ���TcMr�#8+�����F�:
&rg���#Z��N�:�<� ��* ��ctj�	b�s�Xk`�ܿ/݂��-��ܱ�h�����}�:8���������M�NO��<�Lo_�U�l�9�uEH[� ��&�ZJKG,�nJ�N�;�f���h�92��(���e^aWF���%!��(���!s�pX
=�8�E��D
M��V�P��i��9��t�4��b!km��-M��b����(@Ѐ����XdcMfC�(�}�
�I����K�V��zs�c�if�fE+c�þO���W9��gV [���I�;�
@}��)��*>���?���y�uu�XAUw��nY����8WO�Nlq-�-��r�ɖh��i5��vn$��`ݣ C��GeyMq���F,)<d4�5Ӣ�׶U�/��fF�����u+���;f2冀ҕ�Is��
�\�IOy����?r_�g���rd3��F� |�^����5b$4�~~�s����d�am!`<#@Kܣ�ͧ
�k?yԯנ*\Jf�����W��=� �[�h�T���p����6+���1?�#ȑW�R�����M��%�t�)0�-�/�&��MY��77�o3��nR-��ll[�-`���uN��ݚ�^�M�j��C=��q}�FX�y���T�۽�#�o'�d�����X��	�/�~vbor^�^�sv��$5�Y�6Va*�^�s��&�h*�:ř�)
l��{P>Ӑ�����1nB��ϟ��k�u���|���	 |8���+�*�|p/}����W�}'�V4/6)�t|�ǒaT�kO�=N�q>ָ�4P����	ão�K?~�cz��)G�	v�u��r�K�`t���34q!Vb�P��8�P��(�yOy=<�g��H�hE��zgM���瘢�'���֎����Xa�:����9�/�H8��e�^���i4�enz0�5MS~p�DNg'���;�b�aw�`0�JlU4��,@gN��W�Hd�<�,�6�`LE޶��x���Wr� ��J.c�!V��uA^��}3�~v�|�L$�)#%��7� |Jr�/t}PX ��W��&f�S*ū�3����z����N�X8��ƍ۷�ȾAj���Ư^� ��f������֟m�Y�s��/F9eIhx8q�C�f˄�����G��8�%��|Kd��Y��&��]ˁU2�#�~�+]� �X�?�1�� 7����>�d�������✯�	?b|!,�����l�oE�����I|[���4�k.��D�c-��W��M��"uA�.�9	Ҫ�D�J�FvP��5���R�[om���>y�W����'��T��dIK㍥�i{P�vipG���NIt5粧�e�kXe>�D#�Dg��
v8�������������.H�g�)�6)�o���H�2�u�؉�t��Ms�:-vc;�K�I����9���<�~�/4o�|�Z�E�+���V�	��Cpp7{.�5c�&�x�%ڸ��Kb����ݛt-�����H4���B�k�Zt�Yh�%\U\�3�&�ADa`�R�!�F��}�fi? ���S;��C��_@�T�����1�ߨ�w�'��94@,;- It�O$Y��d�E�:\���1�u-z��3.bo䱯�;v�х�����x�k1�H-(NM�9��J��Q�~�՗�Dq����?��i�()�9y�k�Fb�Nyq�2p���E^�H����~A��X�qO�cx?,&��m	�q}�@�	=
A褡3�ц|����v3}�b��;�S����.`���[�G5�y�X����w��#`��K���]��g�=e�tN���$Eke���%�_��u.�zu�(�������bB;)Ɔ,5�Ҕ��Z�M�ı� X�$&��[N�C���F�I�o2�\IbMFjˮ[�SJ�ZX�m""p?���Q��^O�c2�ñ��t6F�&�y�s��g�q��}Gq9�}9�8zD���xy�������{:) u��s��``S�)��#�ĢX����>�ʥ���aR\Y薑��򣘍�M
c�h�E��(���饿G�!u]y���}���I��O�W_}���(]��Oҋ��s�u?ݹ�a��O�D/�9'�JZZ�c����� �����._�~/�N�31
�`� �����A0�	@���KhXP�<;�K^�K��c�j�����)�����֚��,V��J�>X'���`���Q c��##����O?>ѨL~޷oϘ�	9�4�b�R�u����,�o��.}��z�-��~��8^&�Fދqf�(̝�dEG1�9�J��|6[ B�}�F9I"njO���k��;h_8�������b��Q�]�)lr������ni�����X�h4���T#�#/8$I�����޽�lzab������=x����Y�n��(<��h����`E~�TD_Ǽ�w	:�;��+X9h�<y�,�ɁM12�P�X`8�;8��Y�fr�1X3n� g[���H��j��s���;�"j�bi-��ü�{��ٲI����q��C���\Q�w`�%W0�zv���%�|���3�xh딼��~}��`1�5�<����ƕ��%�c�j}E����gS���3��67���ƻ���O�~���������y�y�o::Y�_��Q��	��uˇ����ٚA�{���K��oX��^��G'�b��w��u�d.�sH�;�v��s�� U�7���i:���*'20�ֱ2ҀK����.r����L�Z�2r�:��zZ��}m�9�5��$�F�YL����#�C&�k(*Q���5�+<l�D�%�
u�4Q�N�)5�r�Tξ�7l`n��s�e�i��H��C=�E�Ž/ͯ��}�(l��һC��^���sڰ��e:o�>�f��ӄx��Ou��Qim<��k��1o�e"��`�^�&��7Q4��js���8E��bIf� ��}*�X���Tu_�y���6��P�|v���:�{�ł��$cP?:ސ#g	��v�`�YX{3I��6G2X4��T����V��L8��6�Yx,6lPڃ��u���@�
�:aO��e��\`��0�D�0��G�3���!� �[&UfL �s�XU]��U�Li ԮO'VX�Τ����܅q�젥hW�oE����������&�Hck1�DhjF%��&	 ��|\��)���k@P�ߵ�-[�(��K@��8\I=����I�\�T��`e@��|$\�X��A���4vn�1�&e��VW�	�:���9	F��¹9�l�*�c�y!��D�Ѕ�`S�Kr���;[�ʉ�{�E��R��H���Q.��/�ȭ����tetl@�=�E0�:��RY��.S����I��_n�m�N4 �@��X��!��0y�s�e��b#jOm	�* �-w�6E�;�m�9N�_��Ĕ��`*�Q���F� x
[h��u*�i]���ߋ}��.�:�����/Ϟ�Z����Q���9u��O ���گ��2}��o��)�o�J!�щ&  $j`�A�z}tT:ı�b��s�3��YÚ���9t���W�ٮg�7�]�#�����3������gr����}��T�G�ͱv��f�c��0O���<`!�cMc���2]�(��.�b�aI��dw���Þ�g�Ӿ������������H��S$|�_ -@Y�Ut�����t���'7Q��3�u��N�l��B<h�vl�厞M���<�� �?g3��Cg
�T:u����>�_dr���	��j�Xl;}��xN�p�B[�]�\4C��� uޙ�n&m��ء�L�}%s�񾝦'r�i�^���`�c�Kv��c�d�p�i6cP\]M)-��ǃ�'0'i@���2h`� �����1=�6w�>KX%��� �8��6v%2LP
���B���*��UvYS�иN �p��ak�5��(t��<�,~|�{|�2Ƣ����\ �p=Ǿplj=m�a��C���BH6��F�kA��\ ��kC���Gl�zn��F�d�^��Q�bd�� x�~sl8;�E�/Ox�p� �P�k1�ڗtH��^�|���(�FI^a�: �b��C
��ݕ�?k�Sg�8�8T��
T|.�7(���٦<����~^�8|�h̬T֯�_���9b����3k���f��⎔��=\nјl��7;>Z���Qڶ;~�� ��4	�rȳ;I0�@=g#	�!tLԜ�׵2�3��iȲA|�wp3},������f� �C���KTg�T=>#����Y�_"�^�`� ��1`(����\�^�7��q�z�8�b�X��.��4,�s#�̄�������pk�p��b�Z��S�x���9�Xқa>��8:?�Ԩy�c��վ����x�����U*��Ǣv�RWj����GJg���/�P��f>CN؜=�Z=�=���7��MF9rj�}�ƐgX�q�|YW���xkWu���?h���E=Htb%�5�n�'=�9Z���b�`�z9�֎;�jKScX ;Q_k�w�
�N����5e(���Mc��Tj�QH�&*��Iv�L��#~?�z3����.����������t>\�W�o����ӻ�w����o_��ߠa�:sS.D��x؝���J�1(�Ҿ.y�"h��A �P��H�� \p��*�
6n����Â�"�ژ���Ō��ٹ�����({�VƁJ0�bƾ�y�YŖ����b)���c�LB)Ȧ�v)�	z^k�7����v.Ԥ/��k��P�yN��a�6+�`��l�L�є99� ;�{B$#|���@��h�M���T�p�%R��F���4Y�4-����RE/�����u�i ��e�G!^@��s�sa��1��ʚ��wG� ���<i 5�te��ή�% �Dl�ds�_<��@D��A��5�8��{�!��w����'��M����dE�y*�H�1J�.ܽ;wIO�8uB#x�ă��\<޽'+]��1�����PlPmJ�8�2��	.�g4Js�Òt��)K,��-���}^7+����v~[��H�ᆂCN/�Z"�\���z����P�!I ��W@�˖6�HR�a�Q A���Xj�����u)\%�-'����q{,����zM���$	��9�Н���}^vFR*:aZ�FZ4�=k?�$������u���,�ס�u_��	`� �s������}�/������������׿~â��1
^�U��e�A���4%�6����:�ft�rL$�?�Qn|�4����L_�)5V�_ԊpÀ�o�za�H�^�kt&c��-Z��.`�������`J�����@�i�k]@�Q"I�:�ZZYs�uq�tN�{1jg3 ���?�%}��������� ���;y����8V�o��5���"�o�A��z[����Jˮ�囹 O �G��+q���m�0Խ�4Wt�� ��Ѡƣ��r��Cx�Hj�d�����`(�<�`▭i�X�s�4Pp#�����9�s���=A��Qp���C���3cBg�@ A����@QZD}���pT<�- �Y+�	8~k��{AQAW����y�X�p[St��ؖ{{m�{��m4�ڻY/��Z�0�䄷/���hPLŽv��V�k^�:�#X��n_pD���<"7P��˳|N��|/���G�&
���%��e=+�j�b0�F(���� }������+��2Q�^�����=�s��@��ɑ
k�5Νi�hV��h�|��,��~�kV����TF��h���T�5ġc2
�o.M!0\����>ǩ6l��,���ݜBة��$!���pn��>5B��P��/�]���W2��>��O�y�|��-2H7�E�'�� 6��xf�;���;�ʘ�=zh���d�P[tg�5��H���>z��6x4,2�-�1�k���Wܫ�� �b:`��u�\bW��-�ҕzS����j�����S�����E��Ѫ�I ��Kj�O�!/��*v+ΐ�����	��?~<sm?��Ez�������y�7r��?A��:�W�f�G�@��5�]�wq��{ �O?��~���@�1>�e��0�a��{��g�Օ��{ժ���P`s�X���{�=�qʛ7���E�.�����||zBFϋ������m�d�G]b�Ҩ�\�Q��򢬃�������|6�߷!]�׆�E�&��~�j���n����st53�c��!�y���ޣY����mb�G5ûNM��MR�� w�/�|Li��E�^�A`ɤ6"Ǽ/I�����?�Sb��8�������_�ŰM��|P��A5�
�?}�t�J��Os�����@󷴟=�,��]�x��w�^o��kS��8�C��N�
���g��CE���Ѧv�Y<�Ľ=���9}9w��(O̥��;E^�J�%�\F�rq���X�\�����ǥ� �h������]�<T����5��R�V�f	:ڰ9��	n'��\�W��T��e'����!����1� YP��������{�}_0���8��t*H�P���F<�ڑNJZ���&j]Є��|e-.;K�3��j�%s'�`	O��Mf��c0j��[I��z�ǯbv9�ۃ�p�(��� n�`��Bvk�u��4k��
���Bh6�+�7XOɿ��8a��l�u�^���¡v���_Hܐ�í����;<�A+�T�_����t�Z��]�BLSY��)�eD�nl.Y��8�es�k�����:��G�u�s�� q���Ś��ƞI%��AIيl��-�<8XYP㤙d��ҚuW��w֌�@bU�7���fw����SӔ��Z����C)6�m�N�}Y�ơ���\Z\��P�8LoߝY�bm�n,l�lz+�t =���ߐ:����?.�E� �<N�L���>�����/ى@��,6��}�:'[3A=$: �&���EW�x�"�(���)��Ҫ��,���=���9+��l��a���="��į[�e��]�0ةs��(�pm8�B�ZzMw�^���]��Aߎ��C����=k��',�h���"�Ყ����������"r�Ǽ�}�����Yjb�Ա��67�'�	D��l��+�e2��br���)����^˘�(�[�/ �dӍ�mq����0ϙՠX�J�v�!�Lkp�tL#G�j��G�;'�m����(cǓc�������06�
8�0��ÆY�&�`��\آǈlq�C��skg��_�^j��e
�L�=?��*x(��Xй���)F#���y�ܭy�Vfz�1�4�`#��}�~^x�<���N#>�S�� ��6�s�ޕ���Y����:�kL�(^�M_i˯
�}���y��gZ�^YǑ��btȯ���x��F4��n]�+��we���f�q�9�a����6T#�@�d�����ߓ�L�J9>ʾ{�ܸ�e������S�|>�!
���V:�%Us�1�Y�Y���5�8�Z�n�+&9/�<˿�������f(v�����y�G>L�r>��Bgt�:�9���E����}a���s�`�E3l(@S�i�/�Wn��v{)V�k+��(�ڨ�����/�?�k=!@ȹ��3�`O�'�fϕ��^��k�]r򦎄���Lqr6j���0f�5�ɻ7��Z{�^<{E�{ @0��Ư�I 4+��%W� ��mz�?�ӵ?�z��MJ��x�&hI���{��_��9"��Ԕ3}`��x=����\��~���tã+["�m��us��Xs����d7�	4����0�dF~^� Ƚ����N0�O-� ��2| d,��Q�Ui,�3�k�#��3�E����c��G�~��9:�P�r��  uY4!s! �fDSu�ÿc�!ؑ��a�Y<��ZP���w���.u�����u����}� O�ڲ�O�����y�Γ�}^������gh?.Ȱ�ѭ��2�)T��c��Z&9W:���MY0.��3���: �\�ƜZ_�D��cZ���A�)i���3�E����cv��ݺ���d�Q��Q�r�E�t����@{���@�tL�`t;��~h��NB[���:*5��H�c �a�����Xܔ� )릱	���Vv�M�CT����r�9ީ���٥�2i�Z�z.R&��>���$`Օ9�@�Q�G�0MY@L�d���:(>��1�ܕ���v[�L�N"8ˢ�d!Uz�<M��9MW�v��%S��"6u�T���A�C�9�F���)��ч���8���Nt�Ŋ0��+M�+�e"ﳍW)_M��x\\#��c�&��u�r�M�p��=�+܊.ׯ�jM�D��;�;P�'M�����������k�	^s���^�V	�Py/��J��a#�ّX)����У�RG�
�t�?V���?��}_u\�m�V���z�h; f� ��I�p'��H<0��l/�@"0������s��ܾ���	���?���ƈN
8���Q�#%`!in|�.@v�N'5�A�Ҳ�&W#%[ϭ��1�_��kߍ��^P��.,;�Wa;I��׌�(��޾a'IV0�ʣI�'�8ɜ�i��+X��@@���L&h�@t���B�(��Ǐ$|#��TXL�4H�Yr��u�0o�]2��Q�1[���]�)�? ���K��TǪT̠��?�G�{��0���>v�M���s�m�y ]ߨ�q�����G�����(�z�Bg&·�^���sks) vi=�EE�"^�"?E�sb���svٔ�c�f,@
�{'R!L�T�f�+��Id*��kOP�¤`UU��(��M�����x���&���b�Z�,�{1���l�L"I�6&�2r�k�s���^�������]Nn<b"+o�Z�0ڭ��:�a0ޠz=�;bhn5�l�6U4t�W��Q�0r��Or�����9�H�d�Thl��%6�������"r��qk6�`5��ȣ�K�?f��6�>�U�H�cy��Q�quW���̬�U>&���ĉ�� ���b�s]�W����.���H���/�8܃�͉�w�k(���
p�13���G�4�S8B�VyG��20/�#4I��94�*���3�4�M��#�e�[o^��k+��
3A>PcT�O���z��%GIP���u%��+��OGy��]���ɾ��[���uHc�74ֶ�i ͒��ܠ�l�p�#�(�=_��%]���BkrU�2���b�#�+�r�bM�%[1�i&�ֲK�����YW���`GC�T�������-��o��������?���b�;N!�ɠ��u^�{;X�fح�1s������u,t�B���!D���m�;.�Ä�i��H$�gx���'2�K��� �U719�?)/��Ѡtx�5t�=���+cho7��t&��m��|�5���Pj� ����K�����^N�l��bVYȞ��N ��c����`�`���gk�¦����P��8�%�*��C�7�q���5b<��C�b!���(#�INx����1s�з�=�����k�5�rm�Kޗx.:����0�ЈEz���ּF���;�`9�R��_��@����Y�:.���0y~��&�Mm��)U���^~aOr�o��$^ڢ�<E�;ܲ#&�}���!�����EΛ�й���`�`q#��?��9^��W�g>z���2s�.�cZ[p��p����eQ��}'?�����0
H$3!4��?w||d��-`Ǌ�8+k_,
�Dƾ$(t6�q�1����ptX��D��[e@���������f�wv>Y��+�,ft�������{vk�#5?o@��+	C�;^oα{��+��\P����[S�֍�*��Tl�K�������s��ܬ@�_��x�t	�6���T� $�������qȁ�!@:t$�A�ɉ7G���՘�{��6WW>���zҘ�b>>��.s�x��n��H/�a�)��\n�
��^ރ�Z��@[`\�(Q�:*��c'41��Ti�����J�B7-�`�!8���%t
U8%�:�����E��)i�L �^ā��)Y\����V��>��GEē�s��0�k�I|������J�k
�#�m�E�.@M�#ֈ�nd>������#��y~�n|����ݻ���6e<�\��=�q :@��bvB��݉/kmVW;D�o�+p-a�ʟ"�=B�'�UA@�,o�b�Q�Ck�<�U�C��z�z�hW�w��x0�WL:%�s���\)���~���lk_^���h�_(H1�z'gA�� �Fo]��TCq�N�>$6�Sƿ�u��o�Ь(k%n�_]*��H�T�L�W���l���I��2F"bL���^�9����"���d'&�\]�B��4x�2z[��'�~ǸEg��H�������8�}�����/OK�D,�c[��8��8�/�q-z�} i�=zDP쳏?I�r�3�#����l9rD"�1��3+��9����v�|HWb�\��
��LV�%#	�&��13v��Ҹ
�D���`�ῧ��lKW�ٺ8�?ʷ��J�"��mx�hPNc�:�j|v	pX�E<�s��*ܥ�݈�Ϯ����,z��03��e�ށ�ea~q�����=y����_;_ޟ֌��s�'�b�EWt?��(fzKP��ۜ��2}6�K�{��u��j���Z��&�ljƚ�ҵ�M�v{S���ޥ���	�y
7���p�3c? �?z����!�e��`vC��XҦ���b��u�B�ңBl�LfI�j�	rj��X�nj׷�3��?�Ϯ2��6Q�I�"����H����fʷ��\4?%؆�v����6�[E�;�g� ��Z\'x�8_6HRWքr �=�s�@N��9A�#,?��3���^P�_R��ύu���yEh-��� �	Ιi�C����â��dI�Y��>h|#Ƙ�T�(�Q%���v����O?��zn}�[?z���$��ܘ��VӋ �\␇�8�RNWc^�x�8�~�<)��)��h���3��a�ˬ�U|��H,�u�^�E�w���9����e��^��?(6%����TW;��ֹN�|!/�f<�|ƾ7�96ԋ����.b���D�p%v��g6Y,t�[��ߋź"����_ �����u�E{�{��U_�&�Ts0�����'2x젎�H��O�L@G	{A%���0'ǅ�Lu廵���_�W��kg��4U�bԊ��p�p�P��q`���7)Pg���\�zFd��s9�
1��n���i;�R7�;�D��Z�<sڲ��� �9W��P�DM�v�k�d��>iԱ��;�O�4�X7l����ހd4%�y����2�uZI��G�Nié�L�-��F-ЎR�l* _�if7#���A`���T�������ng+,FPȩS����G$�ѕ/IX�]]l%�t&Y�@q�!lN8� �DW�G!nrS���J~2�7B	�հ;��$�R⌢{��Z;#����S)�$�q(�I�3@   `�ﴵ�!�O��u�A��`Ή���v���<��b���e����u��e���y_������b�V��u�� ��z�녎�l�L���q޴�'�펲!�pt�	|c�$�D�b8��k{IE�I�"�H�$�(v���~��Z�9ݫ������I�h�u�EA�ǿ�HE���]��Â9�
��x���#*"Il,2ٔkL��}�B�bݗ����¶���,�����J2�a]���-�u(6�=��)�1��wٻ+©គ���t8\�G����ޮgɉM�j���9���P��;
��b�I�/|$t��:�{�6)�(6�5d.``��.'��<��b����p ^R����6�T�qou����̂T^��x^ T���������C,��M﮽��h
\����fڍ�k/�pâZ1 ��6���~�~�Ͽ�3��̮@L<#��\��Pd�if\]�e�h���'��Ȫ��b�L�u�|�&���<��A���o߉	�9u�[�.lw�w��%C�n)Mcw���:9Aƚ�M�^k�~X�� ���_���H�w�����kŰ��B�כ6��K���n&A`j����{�]�&ݸ~� �G4�q��zN1�p�9׏��%*�$ZN6�Y���^�cG�Ѻm�cCjRt�ˈQ��{:� [)I�^.�j�hm.� 
$D�.��v%�����?��z(�����~��g������y��Yz���lU[`�L]]2��,��?bv<��e�Egl!�_�-���� ���vh��O�w^����W�����u�?]���^o��O�w�bd�@6���l��<��>'�� H'����*}��os��Izf�Z�_7��Ql�]a�;S�h��:���4�0��q.C	g ��0�`�Zl��}�QB?sl_�D(��}��E�z:>{�	9
y�J�j�@�pDB>̂���\��ȦF��ɉΤER/�PP���꽞f���<vl����s�F3:������/~C'�s��#68:����H\��T��.W���i� N]��Tj1�h�A�s1�\ ��R��9��vy���O�0C�q>�ف��V�7�>���&���#r��m����t���n?�!_�#���b^�t����|���X�p(���'�) u����+�|.ꂙi�'�yuD��q�?�� 	|�ݴ�_{�3�Mn;3q�j�#����`�.��8¶jJ��'h���񧟦O~󹜐��(��ON��׬u^�ϳ?�q,�1x-�Q<�����:c���'i��V9(/`3I�p?\Jg� %@Ty<@���&��+b������6��Buy�&�T,�3�s��SHW�-�?���w5�ΥQ�%�4��r/"��CTs ��u߾;��EHnX���|���]�C��H�;N��F��1�κe%]� k�Q��Ҿ��k�f*��bčt��+>�5;��,��YX �!��̧����4>�P����/r���˜�@:d=�\�}���D���qbW�۷n����h?� 4cA�B�K���־{�Y� �� ��U��n��'C"k�1��D�KNK��&�:�S�;'�&
!�w��^�x�i����8�"4�5p��pC�v��~\�hڐ	t�jg��Y�z"��S���5�����6��F�act�9"	�n�/�tx�c놥F�b�Gge�Ú�e�����hq�3y\�;�܎�yW-�b���P�u�|m⿹S�]R<�p�UB�ȴ=DX<�t؀�@}AÍ5��M�Z�|�,�4t��V�����R=�qx`�օ��@������T�0[�nH�}�`� 8���?(��5EߋI�3)��]�n6�!��p*v>@�Q�\;Y�P,X�VT~	��� �6秧�,�?��!gC��߆ H�����u�'����Iݴ.�wF���+�o lج�s�O k1���:�H��	�|_o��?PU7G�F C��� 4_�������:�+c\���fF
r��=�B�V�1��_F��y��]����P��D�H��Vڕt'�q�X�LI�Ѵ��hJ.�O�J�gʇ\`ѐ����\�D����#���Ǭ9'O8��S>�R_vY[��q�2'��)�Ҟ��`4�����c���F�;4}�0��];;M/7������k�`�{�6�ҕB�5>�J]�����`��M.L#�F+�� D������N�5^wa��1��D"�H6���q03F|Gks<��N|�x��u����B�*�Y�8k'`����kF�n�N�4.
����i��7�k����Iq����
�a/R_'lg����O�n0UlN1��F]$�<� υ���a����͛��w�U�x�4'�>x@�B�u��F�~��gڙ���	iҸ�na3�$%'b���J������٧��ɖ�����g}8fM��+�6xL��ѕ��]Rb[����o�=EwI?��}�]i�x�M�ooQdL?|��g)�P\C*O��/��*Dp����}vc�k�i.�ar �qҪ�ڄ�[.�a7�5r�	��4\Ʃ���JP��� �s��`cad$Q<k=�ƴi6eL����¢gX0[����g��[Jϖ�!:��Ͳ��T�i��EhՄb�&�6Hf� ��,y_u��r�$q�R��yu�i�l�CA?Z���2� �"�^?b/H'M{��C��TK�;��;�d����j(�8��o��\�� b�D�,�x�/��8ڎ\g'A&�f�!��~��#@?��#?\���f.���%Y1��9r���mt�oX,�p$_(����� �K�@OZ���Ic�P\ V@u�YGcErv���o�y@#��O�6w
-��9��rU�D�Ff
���~�=	�#<�+l�!�|F��L�%4.ܬ�`-@ˆyy��2�h˙�&��FM㵢����4�4'���XYk��X�?�>*ߡN��wCz��A(48 �A��a��^P\��^��vN�0HnN�ٚ΂�!�`�n[F�t�M4�8��za� }8��h��T�^ɪ��y��u��Z�)g9/zA��'������� ��׀�> �8�6�?=a��p�(;U�\U�tM���!���h�'✟�5�p��,<�}��4���{���ʽ/O��o�ϙ�dci{#b�"^hOE�c^d�In�;j8��C���4W���1�����t^(t���c���jnnx�����������
p��'��@��Mڮ��f-Կj���vr�=��1��E|>�]�ysf)��0|�6*an6�����,��Nn0��D6ݔ%���V5���?�pJ�O�������9j:����:�.�Gb��8+k7�����uE��y+�9����sMO70�u9�y}�z���% �)�D����dMS6#�]9+���(�KuD1W �F�c�ҍ�$I�E�������zfO�z�]�|��9W�N����4v�[� W~�{��z�$u���xb�s�m��a͵�H��R� 0�a��_�<Iggr�Ap�{��sl"Z���B���M�*�b��M�Y�2�Ǣ�lm��]���ښ6 �X��ś��d+��#m2�Y0^%
�D8�9�{��V�']w�I���0�̓�>�0h ��.xt¢�K*ۑ���!����L ��-EB��ٶt�*T�V:#H�p��|`^�����G���h}x̎�����uo��	��#����Y!�Pf�a����%��ҝ��͜�٢cki'��sY�^��C�B����������<�\%�;�Q6m��^�M]�QTXG$�aO?W$6F�$�'�4�.�4��$�Q%q�Ձ��zV�:�*NT��Uw�-B�N6��
�A]3�t�����l kJu,�)���ݟ� �$agK�`V�L�q\�W���~����?��dB0):VR�yMUW������/��"=��#S95�`��sH�n�����ٱGs���6��v"$m�3�/Ė_�(�/�Ӵ���9���+2f>�X��.��>�D�&YhY��gQ�	(����q�����B��W��	Z0�(�5hŽ�X�r���E�v��S��Fq:~�Y�E&���b<t�L�ɱ<��X�Kp��5<I\_���$��7\�D~��|��c	��
Ǧu�ErS�ƃ-�� �����:ݻ�L8�X�yK� ��;�o��������矧�7o��cѫ���Gߥ�{��?����ŔY�Y ��,��0����g�<(J��&��7��V:'�1��]׊$���5���A�Ύ�~WuW\��p/p�qv]'����;n��F����q�����=��8�Y��Z��h�̦8C�M�bv+&��?�Dp�4'��u������O.��4j�b��ͩ���0\�t#h�1�q{),Ł�s�������j>��up{�Ҫ��/eQȾ�%��P��r<m������i�nH�l���W������P �)<L]&s6�>�+���Ѩ̊�����}�1����4ʟ!:6� ��E#"t;�G�|(&�V�܉�0�7|�_#-���Y��8@��t�@�Lc�f��Cq��ںX�x`<儺:����s:4�R9�yN�k����蚅
G|	b����qu�5,���z�,�I�,Skģ��#�3� �:g���11v�<�B&
�Ʌb���P��U܆��@��s�C<]�L����5U��s�p�1X&`�So#�W�יOU���`:~m�e^wє��5>.�k8|��G�A`�ݸq�u���}�^�Iw*'ũ�b��{gWC�G�
����[�]B��r�3+V !�q�?�&�:L�K�
P�"�q�y��v9����(�}�=�Q3���9V�7��@b9�!̡����k.�j�1`�!��m��ArA�i2&7�=������u����\����q���?��n��<;�$ЯZ���Ctr\j��b�Bv����eˀN0u��U�RݬJ�e���c���y�(�a�v;����񩻈ƣ��4h7֐�8�B^�u�T15p%���(��1���Ѝ7�����[a�m���V��1%��Ì'�� ��n����=�K�i�J��ph��cP  o~?g�G;1����5N'����YiJENI���xv�.��)��}#��|��B>b�	�u)W�$��q{���%���o�)�8�؅ue��W��X�5��Ca��b����b)I� u�粈b<]��>�>0.��р_ i�ͫ�"
�{y��H �x�\����[%��Zt�*�<�yht>O�ue0-#p��U1O�m���gwk�=,wcAJ��8���ڴ�|2[�Q�P
H8S;@�l� "w�CT�5�?�������I��!'�ԥ�����Nu|���\U;*)�蝟9:D��R\�p�vF"��j���1��z��<��Fݝ� �����m;ϭ�I����{��]�n����40#��)�̅=��n�q!����+/����Z3���j�E%�D#ѽؖ�Mq��:��<6�=I�������eų�EY�8�K�F̥�sc����X{�&I��J����̬���9w>���?��/X����$�ntwuݙ����C�,��`�%���8���T�>}o`g���{�����Y��0���Ƞ��1A1���y��fH�>6i�f�V��ђÉV���L�aZ�����r`v�.�9%q/�މI_Dϰ�y�����J�v�\w�V.�Co&� �{i�Ĭp��Rj�I ��=��9�cAZyRy}V�^W�
o�8�m�)���Y��w �����C�G�^��9;���%�����S����b| ��x��n^�ef�2��cq���X��!��t�p��� ���(�ю,Nƿ�,�_����b(^p��i��4��@�vZ��`���Zհ�֫U�fZZ�k�����W_�����(,��J�LI�&uu�9���[���2�r���Y3M�2�^Hǟ�;��$�vrB���e����Y�˚8�d�r=����pj���O���nD��dBgp�h��é��{�1�#_Ocg�gZQR��dZ����lz�c*^�앸>(�!>K-�(��y3k�����SҐ��'O��[���wo��� �]�?���� (6��E͘g�vڻ�X4j�bvZZX��v<�ov�L������}Y/x^}f��o��!�x�a�-*��1�b�>@����zH���/�H�-�>'-} ���Ų��Nl �Q�3��g6�_��}W\,�XD�ɣj'��W��{������i��������H֧������C:N�8zNync��<ߣ�l2Uǡ��Ə�hy=�Yb'nF��	�=ѣ��*�2~��"���t���%iV,���$��o@��1F�}�?"k��	�=��컷��R���*�3���9QZ_��|���,EG|�f�U��+w�Kr�\ɧ�N��C�$�C)��@��x #,����m��ŏ?����<}����x)�Qp��,9T������cE���� r���>�j�Ne�2i�v�b���g�xu!}w�O�xi�a<wj�}��s���xk��"�$����Ŀ<o�s!�u��Osϟp'��(�������z9���g�۷��<r$�;�fs�=6X�D@����c,FgRFG�:b�Xr� ��O�����}(J���s��苀q7�~��)�=%�K�<x�1������ψp���Ǚ$�SvfCq} s!�cC؆.xm��:��nnhi�ׅH/�ɾA�� �)'�i̅l��K7��l
�q�nSk�U08C������EfWi��>y�D�(�'���������'����x]��u%ve�\�0����m�w��-��/�$����EM�\p\�(F�$�{(�-�L`,���>���R�_z��.�v��� ��l���)\N��G�5�Y�ub.$9�C �Y��=�>� 09�+�&�u#�g	�o���k��Y��Z�g�{<��٩	����0�BÑ����<
�T@_�)#������>�v��ܲ��z�];0ǰJ$w�\�3���#��*�s;����4��z,�9r�Ч�봎b���sjj�.r��Lj�CBXA(T��5#8���{�k���������xr�Q����Gۚo�q��r}������ؐJ��)X��7+W���� /�@_��q��PK"ئ˲@Oa�� $�A�%h�4�8PQ�'%o%aB��"H.0��q�q�����[B]�{i��Î��+f]�;��;& �� ���4�M�`�#���s/�����|~|p�)��(�TtPh��d_,���SW�-��cG�"�(v�z# ɱi..8�QHU�W�l}�����fЧq�r�,�푳�X̫��,�rpG�x��k,�HB�>,aY�Y����u�E(3i��_�h
���[>x3z$��Sy�=;v��0�l�q�j�>����c������J���@S����{���>%��am�D�ղ.�� �a��5���?pv��'Os$�h%���%��ᲊ���פ(� ���h	ڭف��(��GJ�G�(ɸ*�:��c��G;X7��Q��{��A+2�>y���/��r�����yS3�T�������֧22�m�5�ן��IZd_��.U�	��c]*�f�.L������f4��{�1��&i�����]�v��NW���8��hF�5�|��!���g� ��; ��{;&Ş	�1Fo�4A ������Z�����}��g�z�A�O�cz�ӏ,i3
��W��U�-�sXڣ#����Z�F���Σu't�#Ɇ�h�)~�x����-��?�VW��Ϩ��?�ۋ���=��� �-Er���B!��
�_ : !Q�"I�~�������s���[/�{��RK)�.ҹp��k�sc��&����u�`��`Cn!k�Y�;*BF�����H�V��O���J3��˞�,k|��M�ш�pDgD�mrMb#'j�� ע����!�:�}]��T��֨:�E�u�.�E*�k�X�Yck�^�!�c������eM�%��GX7[+[����t+xO&1c��Nb�GS�?��|�M#"Α��b����m��E���
{j��~�hy�6� R��ے�oy� ����ro;��
���n2p�Yk��d��-l(��ٌ�O=j^)F2������̩���;1��k��2
kɮK��Zr	�=������Vu��v�q�G���k�뀵Aq�te�����3G�^����{�I�y�σ�b�QIq�i��^�[�Ў�X�~<�ȿ�����Ę��B״em=z��쓅_�׬���#N�F=�ۛy���ȱ��c�3�M T��lD���&K��%�R����`$�8��2��d]_��)��Xk�¸9	[kW��K��ȟ�W�d{w��3���{nj����jW]��L������Ow�r�@	���`1f-45��!�k��^�9@�l��ԮQ�P��ݛ)t��A�C�5�qg�Ik��wH�wh:�K�]1��`��f�fu�Vc���`
Q�~(����cD���W�Yi���Z���KG<H��H�����>j����#eK Oi�MԤ�F�X�Ɉ�9�m�Ѹ�`��&8X&č�{��)'z��L���%�1R���Z�1��FS؃�y5�w��q͗�5ES)���^9uu {5~/p�X����/֭6����9E��g��¢ΓA~[��H���`O�^.�g[��L>�蚯��5H�M�_c�]�̹���+IMjnhS�Q��p��eNՅHoȡ�SӥE�F�z�6�e�k�������7oR��%���/��|u�{�B���YؠaD�ʈ�̠�B�E帉p�y�	����*�y1�F�b����d�:��5Ґr6Mol���.%�e�������>�[�s�)��VOQH'�}��T?���K־>���aH������t�K%ǨJ�)t��͓+�o���M�&�",�O��E�3���HkG6�{Bcb(_�>�Z]��@�b��P�����0ެn��NI�~�	j�V�k�}���N)8���?�.������\.�`��l ^u���a�O��d�� ��X�2�-�9V-Z=.��~�*}�ݷ�N#�y��Hb���H�M7��)"�y��=m�i5��!?�|�d�,�I$'����c�FU�Iqp���g�m�)�����y(l��A	?�d
��{9�H�n���%S�<cD*L:�^l�%9y��g�K�[@&�Q�R@ݥ��8�,"��A0s�N����uIɶ7B<e݆
�r����M=�g�6	��yֽ�E�"��-�y����L�fwl��v�;W���e�=
H���y��(@qrifX��P���_|�����ӕB��%I&h��k�*.�I���*AQ�?�\�Sh�D��b���Ύݒ�S;	ct�׼�g����,F���dv����
�?���:��94�M�����C�:�`�|��WKq��;�Jr�Z�1��� ޺�ݚ1�3�ܡw��$]��!fQ�i���*�3.g�M��LM�h�T��ˡ����9���s���F�gH=��!�n��刯%�w
�l��
�������W�Q��Q�8��l�RC�9}y�`�	�(Y8���Fb/�l���ټ�F��޾���s(@߼}M����{�#ǃě��U��3 {,70�3��[������\���R���1+��~�so�5����i"YV�r.�-��%]:o�}�=��/�&��|�Ŏ� �&q�	ll-l��u�s��rGu�h55���<�F
:7�#��r���X�\a�6k8aa��WU�����x�t�
a���w�b�)���r���<���zƨ4F���\���/�o�h��F���S�I�����/����r���ewQ������y���K�%���������i���1�N����8����T���>X7dc`]�2�&�6F���
��x��F�Q��X�}����F�0{�MB�l��>C\���\�h�w�n���}*M�g�x?`ɼZ�\��'���:.������w�/{�m)�g���=��e��7!����;;�ϑD�Eߦ�9�R��q�@��>�9��� ��O���*ֱ�m� xԓht�<���A���o�\�!q����}6r�@u���������rrM
Vp7�����c=�L���j���_���	�r1]�3�S�q���x�G��wl����Q�`Mc{>�T�+�Ix�?Y_����Jw��	�7��}�i�K6�({qOc���1�S�kt_��.s�Z��:J1�)�� <{;�fI��Z������,f��q[=���
=�ȇEV�}Q��Hu=FuZ>�s�	�b=wwv�?sW~��������9,�?�H����L-�-͟\�#蔼�ݔ���7�r��a�t�dE?���f�q�b;@�7���E���6��쉃�r���(�5��*��Ԯ�,>��)� ml�Ǉ�%���z��uC.��=p��&�(ן�Vdr��gD��PRu�i�Gpk�Bh߇�RV��I�������; 7�ts}��Fa:�۩{Ѝ%�	 �K��^]���a"��^9���7\65m���m,lj QR��A����1�sA�����M0/"�83�k)@|�]�-zz*Pȯ@E�م;i������)><Cе�F�<�����s�K>m���!<�*��^F'%u��֍�$��"�@U��� F��g�����n8Pi��J^�J-��#���� � ܛ�>{F� �A��C'�mm�rD�-!:�H.C�E�M:�5
�F���ap,�.��م[X�N~��%�8D�a_^� �B|Ϟ<#���hf�s��D�e֡=ٱ����q��.g����B7$z�����I~/͝^.�#�Cx2W��`��KP�P�2��<�H$��E!�7Kv׽�p�2��u�)�])m�|J%��(����$*�R�8x6��$�l���S�� elᬻ�$ Ԯ�恵���ׯ^���뗼/X?��/����#0{4�u��o�M�S5��
Gv�c�u�x%�B�=H�cL1�<x5�����g�� ��=�a�PZ�NX���W@����5�t����$KG� ��}�}a����jr���Ьϩv���Y�����ɂۙ;�߇��J��Ź9*6
X☯������GД=z�e���X?��A��Mݝ�����E�+wΟl��솆��Ҥj��t�W�� �?Mv)4x��~��Ba�L�K:r�	qnK��'Ԯ��,&��{���'<�o`;��u��ŏd�@{
�\8ʅ��,&�) � �H9���߇�܋j���O4���9����c~p�]o<�;�p)�N�\��t;���R�?0[�'C{��Xr��Ѕ�����_liы����YkRMC���A47�.���}c�sk�Tem��|����â�����-(�����Jg<բ#�b�t����Jѱ�s���9��h�7 ��ɬ����X�f���`�N5�(+\�A�����1��&�Z��1��rvc!�� ��Wa�Y�[��>ښ���lC\�S�zY�>�Z�|�b��PnY5�V�ջb��`�jm-)������!ľ{�����!�G�y>*��b6���N|��Q�M��e=#ƆV� ���p\P����=�^��o�����.� ���^�M.`��1Y�G���K�F�1+������������-�ŜW=3�g 	pf��"��8�\�M�>���a��W�| ޯ��P{��۲f0r,ƎD�O6��z�f��(�:�)n�A�s�h�H��*q�	4�;���DSck7���k�g�FV<���t�z�G�}%�p�I����UOe}X�D�k�uͧl���О�n�!UV����<�rewg�	Y4?MEH^�Э���i�>fh��H~2�8���?YPǹN��ө�ΨX8�ͱV�d#������Ѻ楒lCi�;H!��Y� ��;��u��T�N!�T4������{���q�����ؘ| ������K��+�[���]����Ql�T��|#�A��-q����GM�KR�.���Wz}����;���M-ڰ��40Bm�� 6�斀�^5�E��LP���@�	���' !|/
	|�|���r������X����bU�u�ŁH�p�<�6+~&~�����i��"�;O��C	z\�'!�H�ph���0�����u7E��I���#7g�]��R9fo��X��NI"��覰a� ��p����#.�T���i 7)���ļe��"���..42t؀D��.�y�|���ub�j�e#ƥ+�b�ST`\��p�'j�=�p+s믅v"1�;�[q�A�{�NY�1JP��� ��N��mz���EyO�L����[�=���C�����5�.���:b1d�r���f)Fµ*�51�k����o�A��h�#Sho/kG���8�2�|F��O�7�����_����v��~�ECp�8,�;���>�Ҍ��G_�V�;�$�>M�mS�4�Y�C���]o��J�}YS�����L�_Y�u�)��C�k�0`�^O�ڋ �8��#F� ���ϵ`NM�ሕO��(c�Ŧ�Z+�:�d��V���W}���rMZ�Q���r]_X�,� |�ĞL0^,-��--Zo�$C��3z�nǹfw�o8����= �r {�\��x+�>�����Nѕ��>��X�[S�<���$jY��Ђ?C;"�)��\7|�G�Z��_����ߦ_���t�x�F"��#F�9�è�,�%0

8�eү�����d�-��fMR���} `�5��e�.n)�+���u�Z&Z$�]�c,���F�@��T��H�j3�Fʶmp'���ԩ�����R��,��ֈb?Ɩ ބ�� M��S
�4���w��yq���J>����q��UW�`�W�K�� =Z�6KnP�(~9�z�&�;bw������`�1����ϑ	��OYW�}�����,�-e�ݯ'����	�$���N�N�����?q|���*6��y�w)����!���]8��(�w�c�\�s�V�bW���e������g��]v�}�ѢN����T4R��oa��.��is��X�֤�}tΌ\99�����OՐa��K������1� �0��J���O`��[gX���(K���Za�W�V\Gތ��)�L+>�W	���z��bd�p�S4�;<����Y)޹Ѻb�E>���s/!�� �3�8w�3�FO/�],u��!�. X����>7�.���zl�n�s@����Ӳ�ߐ��ݒW���O�^<�h�EU�f=��kf.�)��m����k������(���F}N�3Jlvlr`E� F�YE���9��Љ1�9���PL> LP#���uy��	�:���75����Z�fr�{�	��z\.����{[���p!^9�n'f�������8A���[�f!PM#�S3�:D�5{,pm�0�����P�:�¤����'BV�<�Ę3O�lW�~����3IJcX�9b����� ����w���U�{�`~b��.r�]�` �,�@A�W�Ϛ=�UP�@����`H t�q�����-1�W.4ک�"ăr#�r9�&6ߗ5Йaj�V�}���uR����.}d����OU]�S�#���xK�!Te�t���g4��d�X������d�`�j`P^�p��v�fyCE�����cn�@����^�����˰��\��;�"@r.�,P�$�ف��v��l+�_}Y:�e�� �`�\����iI,����~�{&W�[)��H��yR��u�s����֡ !6ԇX����9F � ��O$H�G����Ȯ��=�5#��~-vX�BL�u�N��6�x1�=v�&���l�!(���k_\̅�I�-DSg��5wP��d�_�#m��;y���b�h1��H�`7��A��l�%@��L5 -\�*-_��:X� ���ʟ��*L�ؾw����{�L_%8��]u����W2U<��ْ��o�A���>�Q���젃k�e��L89�(��;���cw��lI|Q�B�:p��*�їK��Yt�8Hv������\X/kw�W���
�`�ݻ%���em�@�K�G����{�s�^�0L|��xs͂#c_|���O���o������l�)v��+wI�2�ʃL��:��3�+`�&E�5Ǘt��6��� � r��e� �"��ňA8�M���O?����b��Ę֮���%Kҳݨ3��0��.l�R����V#d�46��n-t���P^W��c��:�u����
�
b
��.g��G�.����ǯ^�&��o�[���x"״� +����Z�ɀ.5ק �(�C#s�d�Swu쨄=ώ��4�� 5�X)yv�Gkk; ��>�f���ݾ��3���u�?���L���ZP��9��b�@!�IW]������~�����B�N�X��d��O�Nn�+��A���i�e�I4�eq����sI��,�W���E����t>E���Q�s�� g�����ߎ�FY�1�T
� �#O��.
�(���Cm�ˍ�z��K����Ѐ �z����C�9�8P��eN�����yCֲgg��P��_|��/�Ct�H�+�9�����`NP�d�5��1F��Վ��<��{�-}���eձH`�h�2�.�k�;�	5��^/��+�:���؆�ђ�A+.����oҳ�s�J�����V,�٥���v����O?�l���QI���z(��Ѧ��+��r/�ml��]��:z�X�P���b��4��f�zys-
��2�(����St̏�[^ �l����F첵�
F2c��.�r�z}�k���L�UT�e�;k�k���uu �!���
�����'���no�92�G6�e=�� œ9�i���'������`n����gϞS��c��{�t)�/�s@������:.g6��V�?�`���,�C�q����DG�Tݦ��_���H�� @�fG:�:(��t܃c{�N�ۇN摃�[���ke��@�5nD��Jz \ K��6Ӂ���#��b#W<`��q��%���_p��`w�hX��`��AG`����?h�[��l�
QTy�+#�x�W/_�o���ŋ���?�����q�Ps��E-���rӒگ���;:wM��Cv[���Q˞�vU�:4�qW�)�t�ş��<f�"n
��䚥��0���F<�XV ����h�)Y��c��4k�vj��T=�K�3�^Q+�ۿ�[zFi#q7@�^�-�{�����L%cьRͪ� ��C�����{�}�]�����������5urj�ʟ�j*�̡����g6�XU�k��'�)�,�}v���D(�ĺr���$��N��(����N!�9X��"O��F`�V�WK0��T���J@�D2,�}�M%���b�Qtc3��+�^��F'<�%�x-s�u��Q���V���r�ed����b����ը�P��v�"��:	��r!��i	�dd_��i4��)CX�Ͽ`g C�����x�|V�J&Ƶ�D�|�g�� �5�]I&�[�.^Ǯ#��q]�=`a�M�e���U�R(���^�����\&����d_J���$}�Aft[uM�K����,�;(q�?�`;PY��a�oQ�dd���FQV��+	�i��`��a�W^$�D�t��6M9̣�ܹqaL��kB�S_�M��f���Z#��;
 ���4*Fw���_�?���{�#J�1J����([����xq PI�y���FA�|g{S<~?:YCу���f-Mڑqd�M����P|�� �)�XC=�dt�*��6I���s��}|�Nw����x�P5�� a��7�V�k?�ss?�z��U�j<��]������˫�Y�"@�d��i�܋��Y���Tʫr�Lv
ӦO�.��n�r("���T�ߔ�z&8�(��]hGY v�6�o�HO�"P���R*No�c�&��7�w*��!�ufk�{˟���B� t (�u�w�k1H��D K�'��XӉݧ��=�pÊ�	"bp���7
�p���`qr�.���Ἵ�,�}1�$�ϑnr��j6����_������,�򋯊�-��٬4Hξ׈�N������~�6`B�����n�b�ra���3�T�lã(�!����H�FWV1����Db��ė+�zjX]�l} �Z�s��@�Y2���]�nZ� %���!�=��Fx,����P���c�z]�2�����硳`�,�A�)�%���S�u�S!�k�%�uj��I�1�vFV *���3�^�|H��z UV�O��S��6�����B�S�*-d7X���q�'�??E��NҜ�I� ��L�5��G^;�>��d�a��:�XψG�sn�B*h�8;lz�w�Ƣ���s�T���0�zPfip<�p({ �N�7�se�:�Tg5�B�9��fA��gW���Gw�nR��>�sTp��R �*n��M�q�l��3VD��f�,�[Qq�p���T>�Wf�4���ļ��+`��^��ao�ݞ���%�6L@R��9�M
픓Y ���_h�Ha�� ���5���.����� '7�X��껒���4��Q,��b_�U��ߧF���N���Q�OG���G1mZU�FzEc5���%�����*��o�����Y��� d��v�u<�䄋��	Fp�s%gm���� �*GC
���(N��~��8r<l�|c�����Wegt�}���LA�6:S��$��{�� ���ؔ�X���+���m�2�����M�h�l.
+{C�����T�X���a����{�\1}������;���2��F�ie?�@��xS�?��y4v��S*q_�'��S]�3G�t�����"j�BxHul1�3�)��@N�$�W��\���F:�>�U������*��z��Y#.{�c7qm����q�+��S�>'��A��4������`��k�� �~/���?��O	��lg���G�������(��a����%9����P��Py��eJ�NB���o:0���^�,l�ٹ�tKW�	�(��I��{tlW�BA@�2� |�<$7��Ly�C��	��f>)�v8��D�v@^��;:P�M�d�z
E|�c� ���o�Y�_3�x�TH>���Z
l\̲�,���.���ՒpZ�b5�]�2����c�J�0�0����:Р��}���#�Fch�4��.��z�(,�nx���@.���fˢ����o��@Y�y���z�:�%����,pC��۝lL��hΒ��(�<�JZ3C���[��1���ݰ��>����;��"�z�-^Hk7�t����љ�K��T���1���Bsu��a��}a}�*�;u!�F?RHpv'��B$Pv�)&�Ē�h1�"wE�t育���/)D���Hlp��z�f������H���Z0������/��h�s�f��<��ׯ��r�@ 0�k� �G�H��k<���G�İcl�]<�,fO�oz.:y`��b�'(�E�4Y����H�H�s�o��\�Ib���x�&���{�D�s��o�\�ug�'w,h!L;�@z{�>*Tu�� I~o���%�JuߤT�^�a��=�pm`G]��߯v˟�9�ݍ��~��zD�� �;Ʀ�{�5p�8w��~����b}�H�O�T@ݠ(ㅐh�ɞ�+�<0��l ��&��D�͓�:��$b��G-��MN��5�~<j�Fф��Yǯ�2��r��0)<{���i�4 ��{W�za<^�p��گ~����r}���!���DN1���srW���yO����xm٢��=t<Ua�< G7I+��*4�C8���8���X�<z}8�����'���M�ƆV���l]�P%C�F�Y��մA�>��V7XjI��{7@{'���Cfl��V�];�)
�8_|�����D?w\�<�x;���^�~����e7q�{�q�}���sQ�<�9z;��g��#G�)Թ5�C�����RB�	�{e�,��D��\(B��x��g��i�c_X[��*2o��	���n���^��� >��<�Q����S�"�0��G,��/�O��1�[�96���W�h���S�|��ds�����@�\��$,�5z9̓k��LN���;���P��p��)����p���Ȕ��Sh�[�6��2�c| �G4�-��t	�<����8�v�H����"���j%ax1]�Uܼ�4�M1|���?�nku����T�a��+���+� 0�"	l��Z�s|���h:kJ��h1� �1Lӕ~H����Ff2�9�^0vt�<*���=�ګWo
�{}������MIL���02 �lt��^�a��"��W����C����� ��:�X��ގ��o�p���Dż�)��I�.k �s�(ys�D6 Ǻ�j�����u���k�|֘A܈���\ ��� C@G0{
P�Ca6� �'��bHv�{���W$+��:���x�X��&��^�I���Y��A� ���l3�d	�ȃ�d��#��wl�9&�%T�v5!��e}��f
x��L5�@��3G4Ӌh8�j��hbL^+<g����Z�FX4�C;�/� ��ӴO!(P��tM�l��T�Րw�߲��P[�%����V�����q뫑��C�ByI*1֖�5`���q�:�5r�������,j�Fc>����~F�t�����^���B>���t�_�fD��$8�D����WGPpB<�L�\��Q�`�J�:�(o߾�zP���L[n�L��E�I���!ږ�Ua��Q�T
�#G���ԫ������em� ��F0E�"�n�n��R�����ۭ����z�]���5��-�t��XB���	)�Ϫ]|/��Ba�}��8��8Xn�$�����sr��8�j�;հ��v6θR7	#G�^���a_&���bq]_�Ȥ�By�!�Ġ�doڱ㱢>�4_0���ΠZ���z}�VRAt�������.�)���q��N'A�vk/U��6и����3u��g�<�^* O�����S���[���9]��
 ջ�6p��0����b.@&�G�� c�]���ltTrP�ס^ �W*ؘ����B�݆2�=[_I�<��`��]9�=p��BW?آ=܆��m%c=�.�r?�?޽{��'�m���s$�Ҋ�ƺpƠ=��k,LbxE���	�b�T��(�G���éR���|o�0��G so ��� `⠎�2�.[�^ɽ�C��פ���תP��B*B�+۞�.�C�g�|��џ�œ��!A檧�\�w`�,���LM$!(�� !A 3��V�F�N���X�����T�܇nIn��HT�����.�z�g�J�w�����#faE,m��FQ�.�>op(��7���KV�4�����T|_n��L�v9�>9�)�Z�L,��B:��{"���@��G�����=�x;%�I�k�y,��p
v��Z�j�W���l5�	����G��%Uͮ>ڃQ$�W&i�x�x�k��p�����\��b��M'�=�{�]џ��"�a�	�30q_줔�M&φ����'����,�w�[6]�� "^^j����N'���P;o`'�Z�W|V	���\Q�꘺C���4���io�|AW��g�C<s �QO�M' do��fJ/~�J�}���������~�&@[2������"�s��\��C�O�3�3w:Uw�`��(�?b�Q�q�cq��;��T�`/��滯�5<�h�˹��� u(/��"���Q׮=��Y����0�t~���5����cq�����õ�~�k{j���̻���q���� y�VK��M��Z�yS���%4�pͱ�a���tm���'���)
��`D�7���{N��#c���=��A��8��g[�������1.=�t�9P g�݈U��qڟ�ǟy�O�V����,g딯�<w C��)��Jj�2ͺ�\b��f 5R��M){LZ�>-���
���ӥaRָk�^=�|��`bXΠ�	��@x��l��:֟ǵ��]�o����"�%�^/�$�\��b�S-��8�aO0�=�!*�obN˦��]#��!�Ѐ��&#;�:� `�A���d������������x_'N���'哙���n4z� ��(��郻�6�-N�_�/hܾ�4Ί�rd�^J�_��� ��|��b�[Z�o셖��<wJ͏4K��?���5����3�|s��P��C�;����ڂUt�nv"��5wv�����֝6皴 ��!>f-R	���g�� 4i�E%������}�_���̈́y^��!���r�T�C{�eP*���a%�y*��'"���? 8O�<d��@H��Ӂ��������\i�JM1�KP7;��s�l�� �&fz����z�^�y���݀_������K��ْ�=}�+|=�5ɦ4�0z����Nb�r A!T�4��Ì����������Z6г��m�g��� ���,h����KR�eu=���߂	�\�ˮ4j����ϓ���!i����%;t� ������]	O$[��K��΀cϮ�0� �%�y.A��h:#���v�b�(r�d��@�L��g&��<��{���|��g7K7G�� |��c��0br�i�˃GN"i�o8"yy��l�Q�*:�$�aP����:.�~8�CQ�,��
�`1��L��A��t;yxX4�x����s�� ����A7oM���^��뫗?��|�5���pQ��;V�����ao�}'�#)S���¡^�:�f�8�ak�I�vh���ͦ���ʘ��+`W�_E���6���,=(������xj�G��n�`�������<�z��v�<�#oX�+?��a]/6�.=_��j���Db�z��V���psb��B�^�ՑcP҄�9э�b���Tv23�#S�3����I�2��m8X�#�!ˈpr�܎8�86�|^���>�,}�wߤ_�����g�",����g̊a40x�?������|j��.Ї����s�HdY�]W 4Z�;�q�wӛO<�e}>FU�&'΃5�J�Ŵ�'�l�&�>*�&q��}�5V�ӎF���lo���HǮ��\��7c{nDęU�✨H {;���>{�{�ku�k~�:|���y ����ߧ�U�v�I�+`� �ȴ���\��8�Pľ\�r�O�\#��z�^W��:�R�s.p��Ea+�Z0�l�4}�z)�,0�^ͤ�g6��n�%�:>x���Hx�~��cG��l��8�5S���5���|d�>����#����:��zw�``��̥�40��Vy���F8��>��!���sF,���]Rp������,+�g�x)6*pB�*|�F��Ǒ=��qnEm-b1�Ǽo+&��g�zJ�����`���fU�9��t�Э����|�R8;W l�����E�5v�u�	Q~�bĔK�f���@����v_��%&C/( ��O�^�_}�+M%�I����I5���Kh0ä��wj2I�cQuT�/Cp��^3 ��s�w��GVE���������9q�$�nvrAԒ�G�ʫ�����ȹ=��V�rs��k�&�ӟr&��t4� &�X�;��
���w�/�� �c6�K�{k��!v���'F<��E'�\��E�E���sܿ�z�͛w�R$�:�d͉���O��I��8��W<y�8}���)��o��:e�-jh�;��)��s͢�(�[����o2-��c�z��8��i�J��h<�f�B:��p�,߳#���b���	T�8DMe=G�v�$�ߺ�x�4��Ƹ���w)��#{�W��ߍq���]G_��F!5.r�Ç@PW�����Lށ�s�rL ��7 �6�6�̩H�I���?c=j�u����Y�c�yk�&��5�.t5���[����ԛ�w�����$�f���U�%(���E��m-'i��a
V
|�������(U���jC*����7�~����_~����K�ѣ��8& ��>kЏ�W�;�{W�-'>�?��*(�B�V�������f�$`��7��������?���M�KKee�8�5��
�o%P�r*��� u���%�E�	�$�(��1ir4-�({�(�������SW�Xn
)�I1�t�R�QwVN�״��j;c[fP��� �p<'\.�<����/�C<�:;2)����Ow�.�uu0�s���r:!M�{hM�Ͳ��r}}[(�aI���:�ד:�q�{������)X���y�)�pZ���Z�nƞ	���ݱ������{������x��$����|[�ׯ�YqA�ަĆh`E�Tl�M��p �PCCwW�xr��?K�=B�T�3K���Q�*nu�`-��޻��Gc������
a�f'�*:]�k�2~�3��E��� s�9(H\`T�%wV����S��u���X4uS␘�e�=bo�;OG�s��$��Ӏ\ߎ{�r=���{L�T\v������Pc�f�X��ؓG�x.YG�"�@��	��=��+��<��: ������q,���~|��tAL���cx/x�H��Q�	����Nb�e]N�9���ñ�JW�MP�Xk�.� b���t���(ߋ�?�g�KR0�g�K����#�#�ʛm�LJ���;i�>�'@-�+�1��J���'&[1u�v�ڶfǜd�\���q	qۈ�
�a��+�=��p���7[��I��u���P�r4���"�f��`�"��T���c�r��M4���芆�H0q�^i?�����3�9b������֋9��.b��[lP��89po�X�~����P���!���$�5�'�&UZq�%�>F��ܻ(��)�m�ծ�t�O��v�� �t��'%�!���W�s�+�g]/y����X��(��1���Q"O9�%��,/
����c1�КLeD�@ |���uG��F.�\O����ȷ�qY�fp�Y{�܆nX���#ؿx? �p�6f8�դ��NϞ?��ø�B���XY��[|�C�R+Ƴ��5C��>\O��p�Mϟ~��`K�9���ԎJ|���+\��ǚ����N5��A��ݿ��~cs�q�3��ŌM� �����&�_�-#Y͓
 �Μs9��F�hj1���)���̤1w�.�y� f�)P5�1%�*��sS�&!^c�FMߘkD����a���9�	���Sgs����jh��3�{B�=���xN���ma��ݬ�� 8�ׂ�8;v@+y^V�3�$��s��i$A�ܯ�e�.��)�t}G�-5�hZ�I}8�Vӆ�^4��p�,�]�Va�ȏ���*�z�l��DQ��S�\iO_�e4�b������B.�C��]n�x`�8���G|<ה:f"���7��<��c`��l���wv����b�Ԏc�n�nl/:P�dw5��W��W��d�:"�����|�����^�b0������ Ɋ�N1�BD7����8�X�)я͞R*��-N(����rC��7^����%��.貂�O���P)��r0- ՍCI��z@q	���Y�H�J���I���zI���J�����>��t�����ի�÷L�����o����U�!U/����-?)0�v_�v��֛�iPY��?���cvS8/y��K:���NA�<RG���a���6�}qX8L�ft��l<f;�w-? g��b��)��ɑTZ��|�=�Dnr��J��uQ(�>�[1�Z���`	�Eo�F��:�L�h��&�Id9/NԘ��Y���v�?x`}����VV�� s9�˞�mc�l�<KT�[�RPR%���k�
'j IFǘ��8�����d
](
 .���B�_)\>ewg�-Ib��N>��X教b��H��tL��F/���b�"�C���5Dw߽!+zVO�.��z,�	0�:TSaXO~��Xxx0٤FД�bW��|����ۖ�2P����eL�Z���%Зn~<8��n$wQ)�⤰·��.t��M�n�E����q�w�w�2��"����:U��l2�%EA9�p�ؙ
�+;��q��g/�-�L��@�~w���C
�i�4�%N�g<@�R���~�N]q@�2�hg�1;j��956��,�q��U���^:����_�Y��=���"�k\����m��/~z%G����<��B#ȡ%3ƨ4ϖ���u7\
sw�}w[R��:�+_sX0�q7υA׻�)�GԨ�����6�v~g�:s�^9�ۛ���`ʔ��U������{p(�Q�ihQ��O>x}p����e���@�1M)�'� M���h'�D����ܠ����h*ٺ�,G:\q�>X���%����*KE�� �z-g+�ۈ�y��ʲ�^1�֠#F�a������:��P�gl��bB��8�:bm�����-nm,~����?;oٖ|��������K�l�p@�K�N�G��X����K�ǜ�D8*��amH�E��'��Vs��z��k>�zrњ�L�s���$)�����W�0[A�2:��d��v+��4ِ�D�T3�y�$�c����#W���c�Ԙ��|��t�K3����"�_����:E��3���q���O�m���@DrӤ���V�{�׹����\4��3�����6�_��W�Y��x���` 9��Ŧ����\Q��YnA:S�ȡ��x�Qp�غqT�Á��Ԗ��3�h���,+��i��o~D^�jC3긜SYk��ƣ
m�RV��*g�e�,u)�{㬎�o���Ѭ<Y�����i_��0dN��Uь���g�[v��>�|1^[�qn½_�\Nd5�ش�!�k�ښh���`��Z=ZO��i3�1�O�?�#2�5�����b[�Rhw�Y���KM��#�gG븪>�TG/O���m�k#�*#�)��qL�6�����}O��ǌ�������˵�w��a�D������^�{�	WD���s>X;�Z��s�ڐ@���}5Zk����+'��]c�و�d�I�8���麳#��@M�V���U�, ��歜L!�t�yӔ�cEZ��ZW�7�!Y*�ZP� pT�U�����Ϗ>�cV�$n]�q�� ���Spt��f�]BAX�x#�T2����P�y���:
���cvo����[��5�1i� �����'ŕ��J�ݎE�uܬ�;�a��6��l��!�G���������?��A2�C��~�nQD�w�/��A�Dr�� S�x��-]�e��fI�*SQ�vsi�38q�83yB��⧗p�@�|$��@:*�5��30c,�`�H�y��+��֢�~��[
2���J/��X�M�qP���]u4���R�1̳����� �L�����{L����We�0�@�Ay�cX���z8�;kZq]F���KZ��&��[�Ǳt��6sT�wp!
>h�'S�	�ZL6�5 �H�Ǜ�V@�	k
+���a�c	���j��+h�'�U���fV.n���Q[����{�'0��`�k�џ��G�m�.I� �άB6�CMfS�o���+���5�1��~z��3S��ug{Iq+�C>e�>��%9�����ZQ�+8���A9����E����jI<GIE���3
�V$���o#��7麮�����U�`��q>�
]�Y�ع\7&ڸ���1v��	��C�c<��|H�x^�ڴnU�e�kE��Z|?�왋�=��`e�CG�Y]�^lQ�S>9�U�s�����Q�Gze�MJ����_�ҏσ�||�^w��%F
8�������k�UM�Y]'��ͅt0��5B���w�6�,:�����Q<�f��-šϙ:m�Ua]멬͈�5�V�"��gl�a��
��c���W��M��+�ZGS�	��{n E;�:�m*�H9��(��g[פ:~Ҍ �g���-�a�#�nDu��Ŏ�)xSQ�G>Q����ݧ�G8��33���6C�	1i�����>$�GͲ$P����ܻOqX����Q�`�Q��Rڅ`'$�}}��c��w<�c�h���B�,{����NM�2����<�J���k��Ƹ�#��?b�)�IȖ�s�?�$9X&)���*]�c��B3
�hL�3��Np��c+�ÿS5;2ƲУ�0�M��9+޷�,�O�Z�ف���Ec�T�2���+N� 0�U���x���Q�k9�,�*�p1��$��\^
ğ�������N�`Ƀ��soyR޸��z�̖�\��'����n>�����>�9��s=�h[������р$�;k4X��j�,���c��e=hAE\7 |�����./�����ܶ�RG^���ss�d�rNR]9W�a�)�,���@k߰r/���y���s�c��D��$��3u�]�d���U�B̡�vb.�}�� �_�&�]��H��nJNݼǂ��l�!�:U�N߅���l�������]��̯�樜�@�D~uͩ���@����IW�.
�/)����`y	4n���4ٔx����tl<�zK��!mƍs�v�@k?��.��<pc�M0S2Х��ߌ���_��G|\���0`�<�Tg���ϭɻʳ��b�?t��o�1����F ��0��Z�>cڧ�h��y���K��l$�Y
�(�ɺƍdC�P}���u֞B�cs\E}0_���b��Z�:�g���y�k T�u��a�S�����#��%y���,H\Y�F?���P�g�[���� E$
�YM�p��	�%6�!�Z�+�r�@g�(��q	� \�NAR�XJ��/���@󖀋�xW���L�ÝD����a�0i��Y�gO��9_�Y~]�o��&����q Ñ�w�����<_�>{G�<D5�[4��RI����m�Z斷��8����+�)��)Z/A����V��`��,*��1�$��J5�n0:y�t~v���_cѮ�0��g��T���0�v�>p��U��9G��kQ�~_�� `�=�aV�`�ˁ=T���\Ԁ��������x`o�@D0��8~v����	"��@�WgwH���x�8�:E���8:P;f�9r����]�qv��/�3�w�,d(�Guc��>���4�%�Hم=w\Q���n�$�蘃�=}t�q���;�Q`Ht�=���q~�J  V��э�"�y!�d��XمNĩ[5���N��I��FǨT�^�'�)yuu������g�IĦ��Lg�\q�rL��;a��>�z=b��V�4��L��.�;��Qa���=����<�A5�X��J,�V�����?d9���*n�x0W���7��k�A��A��b蠂S{z�����u�Ĥ7o��K�.p���f���rҙ���e�%�Z3�;ø��4U��f�,j�>D�?�]e�;�[��b�K���"���޲��/���kg�����{�/`�������v�Xm��j��tR��H��3e1W�a[���q1׼`�j�����fBS0(3Ƞ!��ۏ��t��K
��(������0ܬbL/�h���k�F!K�0΀���D2�f���LN|�|�)��ke�he*���v���#aF,0ظ�Rg�B���p�w7���"��"� �f���u5:��:x&�<�����l�`����aZeX{��
�IB㈱(�q.`_t����C)�����늋�����\p�&L^>�����O8������tyO������Ȏ�?x�⁳с9K�0]Sl	]�y
���Q��R�3=liY�ut���]mQ�W��5cu��D�N@����P~n��Ѻvj�Ʌ�����!p������P������K�qƅ5���wf��>[��H�]1�m\��'��|9��c�'����~���G�Y�V�� �4t�Ck������S�o��;�"�]W�PGj[�+�K�>�l��t�'=��D�/�,��\s9�P<1��=�������җ_��`�=�&(^�#u� {���9J^Y�A�J�T)K$���%��
�s����L�z�+�_�:��	FQ_����AQ�2��7���F߾y�}����ٸ�83�gL��1s�e� k.�{�*��|���=ؑke ��k'�48zR[�/5S<p߱�p�H����y����3���8�����bb%�wt�U�@����'����3�]��ePO����F�@h��d��&�ɖ�(�9���W�`�Ĝ(L�;7��}_F��@1
��i��� �����������Z`�������F*�97���ъɇ)S�َ;{���X�=ן�ǈ�h޴͜��~�2��}���m�O��>|�����{7��HN5����;lf��YI��M�EIl��#�cV�k!ϔ�H
wo���������`?�K�S9<˘͝��*k�.Y�
	���u���7��]=�_�����Q ?)�eѐb6���KM�%,9��I���[ۏ�(V�	��,.��Nϟ?c`�~ǃ�h�;�� n��k��@�9F�sp�s
�����[�%��v�L� � bX߉��Sw�]"Rl�����y�#��������!��FD*�Ş�'Rxd�<�PP�nF�pC�%A�Pu��AW�v��.=�#jp���y�Y�I�Vq�z3|�F��W�X���v��c��5��q^Sץ���{$Fd��c��=E;e1���	�}v��V��}/����}�.J���d���s���PsUg�{ ,��� FW�DUD碷ty���Lݝt�nn���ƉWg��)�%��}��֖ZS7���P��"�j�4�{.I�s�^�J�+wE��Ş��Ld ��nP�kq�)9g��IT:ͪq>�_��a�e��u�sj��Az'f	�C�����O�5���We_���i¹I
cL�,�.��u�4f���S:6<��s%Z�,j*�XH�,w�3+��@r�W����G�t���M�G��� ~�.[�RH�_��þ�(����q8�Ŏ��������,8!rz�k���ؼu\4K*�N ���/zj)��i�1��27��5��I�;="�;�>�O�욢;[��%��}��[������X����h��׽h�!�-p��|�;��Ӗ���̑�e�ȦT�R)bOϩ�'����>��ǫ^ָ5̴�֘Ye�Pp6%3.�.��������1�,�!@�Z����y��ۋ�Hv'Gŀܸ8"t}�~���tx*m'�Hj�͂�{�X"�r�R�v{C��]jDY%�͋ic�(�����ˈ���u��6�g4�y��*���ۖ�FQ�ς}3�/��b�_h,�r>וo
����:��h:�h?��~X_:�h��: �P�~c�E8�6tjr�kqҎZ���\�(��ڬZ�0�5З�M��#J��h�l���Y�H�K�a��!�{܉p��聙��u*�$��ڞ���XW����l����$�5�N�`5�Ʋ��G`u��k�)�g�����{�r��޼����Ģ
(� ��$v6�6|��/��u�:��w}����$����ɣ}K.�`�&%h�dę�����iE�5M`^o6�����M����$�î�GNΩ��Y\.S�p�C=?}K|����o���ZNQtF츨s,����	j.<��K�a�u�1�ԅ'/��,<\O�|),P0�f�˙F�m����oa�<5 ����ךMX2h�g?��s8�?Y� �#�g�:�]��<����Lf0�(������x�Qj0�E����ƿ�����e�������\�8hUMx��&އ�U���:���)]LŸ�-`�k�����.��������ڛ�8���T�M��Y��ȯg�V_��8_*c`Ca��]\n���E9sB3��c��޲2����=�Axk�@SѺKU��5� j��| �T���?���&���֬n�`yG>~�1���5��N����q�Gq"���s�ҕf'�C��h:��M��Z�.W�͘���Q���NU.\J�t�o��f`}`LK��;�͋���(���ى-	��UL�� �b�L��e�H����V�ǌ=
S����k�H���c5�� ������0��έ�;��!
�ʁ����q�FD�ַ�N��g�	>cP6����$��Ԉ��Yc��G���P�bHcq��}�9EN���b�AA��Ƒt�#
k�wr�|]�`ȩ0��f'�J�>�!�B�f���\�blcJ�<-Ϸ��L�m*�=6">Bvb���J�~�k��:s����<{��Bv)�R��>Ԓ�H�yO�T ��0b�����ج��|�M����,F~0��\}\��twB'��Ě��t��XN�a�Hy]�|��`z:�T;}�u��%�p ��R@�k�<E"�)n������F�;�޾��졺�ܣ���ZT0��RX?F����BbGp,��m{��2�������`�χ���X
@���zmC��n!q�=t�@��6�)��8���g��
H�{�x��!�Q ⻤�:x���S�g�A�!$��:s���V0F�8��@z:^1���g���猅���L�B�k���A<?�9s2g�(�W���R4�;�d��f�sQ;ĝ$Lr��=��s��Y��	ؙ)@d���8~�l��䂂��Di_�X�Z#51�x��&	u���CK���F�	��HfT�E����C�N�3��hlh-(��_���f���� ^t �yT���R3���m���c%�&U1�h8�%8�W7��9gՂ:��T ��m���<R��nʡ1rS�M��[�	
�\l�NZ����N<�U�0 �gJ���<�X6�b�QBVY���!3� ��O����۬4�)-o	��?~��5ͪW�m�]XЙ ��D��.�}�v�E���ϵ�D�ɣ�U#L����W�;
C<g�ҎE�XO��K~d[�}�8a��*�x�|ə>����rx�^�x)�l�CK�,͔���f6���HsE�7�
�s�z/Z���E�⪷|f��C.�	3�[ 3
�i��X��<��RRG"��),���K�Vq���O�(Ro-�`�"�����f��Նk���ƾ΅d ��iִ�؁V�NN3)p^+��"c� ��p��frZ3s��6?	���1^B�j�h�܀�H�X�(��gK�iI#�,!�#g�8���ƅa�(9���C0�����d��
�:��n�˟`��&=y�~9�n��'O��'���g�V�ߏ/^$��*����0���;�qߩ��1I���΢����1����Ú��c�$5�#���;���%�6q��i��b&b������8 �O�}�ޛ�3+O�}bK-�#]1cob��] q��<s1ބx(�`xݿMc������N���>~Z�לoJ'�%@�#Mrnx}���^�Z|��I��/YgP��Gn�� @��~�A�{e3km��|>�6���?Zi  ��IDAT���5�c5��m:��4�X�s�Z�;6� Ί�<Qql������:�s�:����z�Ǉ�+��R*�S�![|b�9J���N��^�L�t�hfޥA�u
�`\�Xo8gSRi���Ē�e�f��_Wr�l�I�i�yD*��9���W]���N�N~���9�u=9*���w7�5vbÕ�ē�s��'�#H� CS�� ���4��8<Ak�L�2\��ڄ�_],��9K��;C�}F� ��t!��ޣ����g�
��]�/X$�C��E�ٲP�K��AQ` �N�=f�~���֑�sA�;�`m��;��{�����)W�< ���e��N #Fq���܃��粱��m!9[�Gc&猝����������n��q�^n.�:��:p��N��ӽ�l�s��3I,�*d�D%F��ՕXk;�c����R+�5��M�������f��f������>p:Oe��j�ԕ�R����wG�����Y�+�^�������N��H,9뚒���VĦG�I9�B����ۻ[���(���=�7=z$�iJ)��{}����ⳑf�-P�5�xz��F�L�-��YI����N,�m
{�j�u(nO����aMV�s��}q-�ƕ�s�2ϵ[�ܩ�ā���[RO�9�ho�#4�/�����q��A�]��/�5��}���9�4��T��N��Fw0*{�/k�����uJ�`K��yЇ�5�K�h\�?j�i�}��
\Q@.�ےy�	��+:)[��ui���{iEQ���z��]��B2�<v��W�{`Bn]��ވbC���	������ô�^��ظn1�j��y��16mM@@
8�t�,A>�!0�ś�k�>�D"Kܽ(��C���}i� �ج�<��PF&���=�87��&��ъ`��9�G`4g�Aa���ڬ��K8��yp'~�* x�;>��5]�Ȓ54��}�.]�ܾ�T~�����˙�5��,�A�����J;ŏ� ��澾�(�r)��ts���1��9�bO���/���	@[gI��~0>�=�4���� *�/��Á����Y`�l�D���%�Z��\qq?C�d.������è���Kk&�	0����	�`4M��B�e��Z�2T�`a��*�o��[y	~�Q_�q<5��׋pS�U# ǁb��E��f)w���^ �&���?�j�Q
�6�(��r9�I׎��F�*�V� ��R쩡 P��t��6�� �&�)��W�cQ@?[�(���U�}7fS��v-:$��߁�P`#�]�<�`�>(�� ��Z_���i�g��6Ej0詝�Ri0aݨ�g�Fq��wP~4�3�Yl���9� ����n<�d^a�%O������5�.'w �ql� 7wB�yP�����
*5����ډ:������Ю;��E��{l�~~wiv<
���S������b���h(��ۓEѳ��"����8C!�#��B��O�e��F������W���Qn�z����^���s�`�EQ��4j�`��1�U` ����G<k�|\�3�ם�F.
e�Tcn�:;������-�IА}��	?/�-:;���g�\�x���=��)�WB�b
r1�&x��t��|�ӟ[\q�0v:?,͘�đ`�}W���M�V6�΢i�u��K!�ܑ��A�v<�'��9v��b}��.��m���ٯ��N��;����ר�V�~�߬HP"12`ӕ7�a��A������]�)�s�/��"0�ä7j�Ξ��R����Q���+��{�Hp�h�l�h�5�U��Ϳ���n�Sz��G�B���Ww`��� �!T��u�G�tp)}�ݻ�t�0r<�ԫ�� ĜG�"�+����2E<��\wJ@(�7	(����?��N�����,��`-�Z����w���>���4�Ud*#69[4��������޺�ǃ�^r���]�v�9��p��E�N+���3��B1m3�,�5����sv*�����f/�ݞ��6P���H��x]좯�j��mj�X6��L��8���F�%�'�ٌ���+�|�U �	����X7bwi\i��Wt"���W��x��)��z�G��� �&�-�j�nW 6\7�̇`���oe]�S��N�.V8��20E�  죝��`K z�['�?��e�����o.:N v޾y�.�Ѯ_EP0�쐵�ئ�V��T�ԕC��T�~x3�-f[�i���s1�8��$(��ʮ�gƘ�����3��¡�]�[��Z!~�)���tu�/w�����s$)��7v��f�ʢ���F�E74ܿ�T\���U�A��H,��f��A��z�V�
��!��	���H-��)Ix������D,��}�A�
L���У�mӽ�ˎG1ٰ��cd�@:]|�yO�ͺ/k\`�cLi
�@�9S�j8{7��+{�F�(f+(4W�e���nj�:?��i���ؿ�ѻ92�!x<���1`�}��K7��4[о4�y��O�q�\p��d"L���u�:�9Ҏ3�v��C� {h�kl؅��`qZ�AX_��DA|�*&n	v�{�0GWNkI�<���`an�l�m3ױ�٣R�͖8��Xy��o*�q�[���,��`�[�eD��Y9�4�p=��3�4���3r�9���!��Z����<ꂿ�uACC�ҡ4_�;�����OW�a=ѣrh~e.��&�4*�1��-D�#g�"��楞3�O#Eg7�'�+������Po͙:#P:{��P�3�Zӌ0!���rmW���쾛�~������*B��������X�6�H(tObd��a%��l����Ƴ���IB'-P���Y��fa�
�z�bl�	�?oo�%ו$�ݷDD�XI�;�6V������t�y�>I#MOMwU�H���5�-W�����L $��F��ˋ��당�9����d�+�N{��z){�޼=�Tܷ,�n˺�Ϥvb�X���ل�+#;���"��Ƈ��f�~�GS�i�闿<�~_�+�1�>���;����(�@&��1s�l"�i������tv��h3Yk��B.�X΃{��Z\`���w,������G�{��!����]��(�0~���\l��������Y���u�<og��暬�n�P�k&���[�8v��U #j+$�ܞ����A�{+$
A�+���(�z��,�a�W��ݻ����!m[�Rˤ!�\�Ɂ1�sF��E�b�/30 }z��;wy�. ��؇�"��n�[��ɘ;{���YN���>����MWΑ$�oђ�޲���GQ�S��k�=��F�z�G~A���՛E�
@�<i�U���m<P�M�T�e��HZ:,�����"=��FOC�mt:�GҺ&C�T�����b�[Y���nu��:L*�<�?G��;�I��)PR8Tg������T�}lZ�Շ;�
d���_�x5G��h��=�J4���$t���T�s_��4#�;�sC:�H,�-a�M�kㆣ��]Q<o���'��krP kc��.~-aE-B�[4˶6ntM,������[D�Q�>���ט���M]���*�D V7�;�l��&��� ��-\@��bJu�,��W,4��F���־Q	d?y�	*^#G�5W�q	����V�Y����tF�W`��5��1��d��a..��R%my!*	Pf_�X�0�6�N<PZ�R6i� ��	���|���5)�ܺv=I��}'���wM��@�V�z�D\�Qmd`808\�c�y{�@DU�j[�.�1��Ϩ��T��8nU�RM8�s�����9�6Z�Ne���M*��%`�6m��w�Ӷ-��B�n�ޗ_��l�:k�U6l��{�솾V$�屛J�ncG����F��!�g�\���"a�� ]ӄ�2��r<�����?R0@��O���>(���^����hq`�6����$�V�Ֆz��l\0��6P걞��6+M����
Gދb�h���g�c��߈J�'�n���V�nu�?Y%�Ga��ZB0p��D��hu�J΋�[��;E7�#Pq�ݧ:y�W�.
#1�x1-k�~�%����j�8���3 ҁ��<9�����Wc����%��d���Z�tj��<��G�)>��q-Yb���Ą�>65���5��d{yY��ތz�����c�U���X}��kz�n��o�\U��W�^�^�m(���V��Ob�������4.�[kq��X$LޢvmN���I�o����Zv9Y�\'��lz���ɞ�CŢl�ʑ	�O����9]�8���W����m�;��YNt �d�/�q���_�A�<<�ck�@��U�����3;���_*15� ������kR���6 �N*{�~.��EMq��$����H�;h���1�TFm���[���*Fh�jL�K��S�m ���MpÚ�$+�\GO`����0J��`g�*�O{(��om}m�ᄶ2z�V,����:f�p�����9m@�e�$�ā���|+����UÖV��p�N0��l��i���8aΥNOߦ��)��"Z��T����W�������yI�Y����'x�]��y,G&�䑄rd�j]���+�r��XA�K�Dr�,[�Vq<W�f)xn����s*�f��U�|��
��@d��5G��飇j��w�ĵ�6l����j�������z��������y���s?�(vc��G�5�� ����\�;�b��0bG�=J6��=pp�R%w|��e��鳲G."�ƽ����Ix�͙(�=?]_��Zb��:`;�x���qD��b#05�/�<�������ð7�^�g4�͌�XZ�՟z���	u���ln�̛����Ǚd)�k�~�Oy���k�F���S�噘C���c^����!$b��SE����
�x`ڦ����޻�O�I5屒�4k	�B�u�+В����h�]�6�X�$�?���-���(nN��fm��JTd���v��&�����ON����,��D۫k�P�~�K �v��I ��v��
U�2K�s˩?jm�sezR�m\W�H��Wo%��e��U�C`�0���S�b��wj�_YV!�`gL�Z�ni��]6�ݮ�5JdLqQ1O	j�������d���tl�n\ʃ!G�}�����R�� �H~�崈�<Q�]����� O�U8Hi���dq�AbEr�JC�{���gc��Z��KU/���wNX�E��9G��ۮ���v7�+%XC�,1Ї@�G'��x��ؑfc�U�;�n� �,�� Mu�)cR�w�f7�_���\�?���-	�Tj�����m��6�A����p�{�4V�/ކ 2Sx\�@�b ��~gSBd�݉����0��|&q#)��jK[7H,��#fw��Jf�XK�Tk�+����ۄ�� ̭��	������v�4���D3���9섯�dk55U4�>��>i�.{�g
1x��r~F���9p�\bNϞ=�=��c�'?Lw�O�}X��Q��x����SktE`v�d��Ȯ����37d�W�$vO���o%�nZ�f7&c��6����[{�l���v�0��S?;��˔s:(> b�
h��̱n0�<���Ek'�ec���ԭ20:B�-�YW^-��F|�}+�x���|�X�rh�0���!	]�:7+J�æ�+Z��Pv�]����n ;��|{�\��-�'�-�d�	���dp���ڣ3�9h\�������W��8�&�U6Q�I@��x+��%��[N�D��6���HXT����.PEz6A�T��u.f�� �Mb���i��4�4R]����iE��k�Eqm1�`-5nG���w��`�io��Y�*hL H&``�|�E��Ӓ4�|�M��,��d-���F�: @��P|?+`��L]�@6 �\)~�,xd xܮ�<�n��%���R9`X�ɜ��#�+(9�ELb�	l�۰��+�V�֞�X��cA�=�>�Lj;�b���L�{�5��P&�m�j�޶6|��9���
���@���t��X3.YAH��n,0�k�����)�@a��6�}ؙ�d����)^�W�k��=:82���|��i]�3Ar��m	&n�}{�)��T����$�q/�5�:��u|������ܜΤ��d�2�e3�{"��F���ئ����_���K�l�]�w|�l*�Иc�С�b�@xS��F<�YŰ�����d�"��^tr&7t��0w�%0�P$B�1- P�.�UBfXӄV��z�sa[�y1ltz�xquQ��̶��U��������ۈE*C�b��uϼ;��g��]��x����;5=��~�ټ��PLv�q���`�q8��T����7����C�Y��A�d����^�i��%'�7%�ŵ6�!<l�#���=�b�;������s�έ��k��ԖNV�N��{)��B�b���&���h��u{dj5�f��Y�=f����P���*dU���(�M��5o���@��)Y6G�q�(<d=�eP}m9����0��/�B���p�&����8n(գp'Ę��V��ťRܟ�: �BbZӁ�ZUq��Ѧ���#�tj���X�J|�8�{��8�֜��@ "M$I�����Bw!�ų]�OX���=`��W�5����h��f�=&��-1g´򱯆gmv�z���,����;Ciن�Ll��k���y6cj�=�6��FЮjȭWv��S[[��?��F}v���7��=�x�`�*o��C��� �!q/O�H�i�]������s1�>Z�Z�L��:�waLW6Iɩ��'j�r���VÞcRc�Nk,�+&�e,F`��W	Ъ�gb�l%31��Z��J�g<Fef��okaRO��k�5@/U�� �#&p]pR�f#� ���+&�R�ʭq�Վ������#'o��*m�����ʴ�&��ص����ׄ6���3m��������I^oc�R��Yf���C� �)��DЇ!�s}{��!���k��o�b-��x�XK��	���?��������������ɪ����@�q�+y��g7�к�֭�Z��{U�E߭`�ܢ��i�O,�In{�L��#�����6��O����gP����3��s����s>%Hv���V�<����A�1�T��ݸK�_Ӳ��m�--�Dn\p9D�mׂ�/y-����U�彭�h�>z���7M\�t�'���>��4aCB�]�t&�V�n�Ab�va_+eރV繶_i|oe�H�$1!��dK"F�������K�q�n6�sB"��-�МX������ceHr��ȆXk���Vx�`�&�ms�|�5���.c�W'��5��֢�b����@2��/��f�5�)v��,��իW��y�k!�5��l��)�$�q�~�k�M�R+�zm{��.�ʔ#)��j�Y�t����qi�UV�'�)XM
U���϶>|!�͹~�����# J��)�{��m��"�_��\�2���!g�h�b&{`3Z��F>�7�n閴�g��:
��M��{��F�gGPS"���5��q�I�)Zy�'�c/r�|GӉc|2M���p�\[&�J�^?���UFa~�m�O���<@��Yv�U�+V�ŵS�����e��~КW%4�&�P���b�4j��|�xѲ�������c��|-X����(�"�L�[��4�ܖԉ�V��\���8�w���m�`��6�P���]�Α�a�Ṝ�<{�^�6g�V�i�X~�6iƖ`��k(�\�α4#1�
1�Ǉ�NOW���¡�;Jo��ƥۄ\7�M�I��!�Cny�����6���'���d�K���Եd�/ T"&;�x��P&4�z�>�p0M2	֫�mZ���1=+/�r�q��X��"���փY7̜wQbm<��[پ����ݷ&`�g�"A����&�ݬVT�P�E[$���l�7>U/:1�u�f'��$a�.,t�i���' �şy���H}�~�H�c�U�M�*)6��}6�Փ�T��5��p��1�wM<j
pG��2V��0&�3����\+l1��5�l�,����DKQ[P�To5a(+ ;��gꀜP�
�I�p&Q�d�O&o;,бc��N�nA�4�8�+�٪���)�	:&[܀Sv���G�c� ���K��i\�1R�� |��
�vD`��s$��n9�� +۵�8�(o
�آ0(@�p����s=�5��S�:�ݭ�ナ�;K�����"	�Jt~��|=6ԉ%n�������p�ĳ]��
4׍���{8�: C0Gp����Ɠm�bt�N*P��{��0���,tXwN����\��g]1�|B����;�87�sP���F���N6T��dKT��R@��\^RD�Ńi�x5�A_��=c��M��!��,�$��7�+���3�*Jl�Z�f\���ĶC�uyqE(������𲼏c}4������	��y��H C�����6�#f`6�k{ҜC��[����J��z�|8��R�h	��`+�6����ʆ����-��P;ah���v$`dd���kvc�.�8:�cE�dُ>�4�q_{���.�\D{��iz�����)�ޝ����?/��ҋ�/x9���[�v�d��-��&�ʒM�Z�ǂ����D�&�KbMU2�1B	���gݭ"�_��d�Za@-)ց'Zdጚ҃���=�U��D`L�k���~q;��a�&(ؿ�t;���ֻm7`�t�m�`rrf�/�*��ɓ֯?�6ē݇��_���d�м��X��>���C ���_�C\w�g7=��M��b/0f�r%`�6}n4���#w�쩥& m��(�(N2�D'�I���ùe�ڋ5���K�ghAIwp�t�Ь��ȶ$0C�l*��s�L�s�׺F`?�G$J��^/�T�;�IY�ʔ@�F�����T�u����
�@��K`����`��~����؋g���kk�uF��r x�L�/ĥ��f<1��h?D��s$H<�޻��[�?��69�ԛ��8�o�,$Y�b{"�
η� i���A-��,�U����ND�`4����g�TL�4`����цeK-x��\ �8�U�Z	0��T1�9����Ź��Q�@�� �lU����i�l�p�B����|֜}d�hc����P�q���>H����eC��� B/��ܥ;6�]�Z�([�ޡnX��O(L@�g�y��F��e�ӌ�w,����T���Ԗe&ha;���@v���,^5~��u��k����@�H�����-��Ք�.���[�v4�
�k��qF��X�b�ӽ�y�'�����&�'�w���0����§�\0���O?I{�����yȸ�����`�����:�V��'ĖE��tؙja�uk������ꥀRn ��ɏ���K��[kT<���x���=���G��@��	�[k��=��"'��1@trQ C�홳�kd0}HM�fі�������D�C�se+)�2@/@�6|I%i�B[B<�>@aH�Y��q���k��S����z��#c1����s��e|�����ٖ?�����P��,�|�`�S�nnDk���S񥭐,�eGR��k�6X�k�+�_�2;l�rmS.�I7�P<mr1Ԇ�X��$֮�cB�.зv��+�'�%!~�ڤ[�`��ն=r@F4Mk�a�{��cSl�^�YT� ]���EC$�t��b:��걂�����u�JU�8ܰP��[Y�nU6G�{��߾'��ZE���挓S�e��p����������v��+�$[ �	�Sp�|��X�L����ڦD����x��bx�;q�Q�MĵV�zz�ėx�3M TZ{^�A�q��Z�9-�D��,[�H��`�TC�,6���_�ɘM)\��x�Y��+�l�̤`R�y�y U;5�1J�L''�)�dU;G���^��w�&1`���(O��� �;B?�	z�y^lI)��(�ʪs�������{��=Fc��p:ԛ3�-���&�<���T�����x���=2��ףּj����r[�9��_^fk	��县MÖ�Ϯ�$fݎ��*�H��T���/*'�Kk�������Q ���x^�h4���@V�saL���9�u�A�Vv�y�R��y'�+�ī�ج��E{$�t��]	�l��Fx&�T�T��4�3�n���DAk9E�F%��ˎ ��*�b�9O�Hu1�A�iv�u����m���_��{wY�A�����OuN����&f̏4��Y*J&l��d�.��;�f�9o��X��ڷ��&�)��<�3k[���Uؙ�e�z�ZE.�t�j-Y�k���\p'C7�6R�H�Ր	���m�FSW��a�Z^�$R�i��k5h��Q���1ߦ��4�n1F�m��X�|��r��L�) �s�����h`_gS*oN\��� �|���?�y�YL:/^�w�Z�}�z��3'�A/�����[��36�.yի	1���a�=/��'��(��4j�"gy;��[	X���
���S&� �8
��70x��?�������+:a2��?K����1�d�F�죴d������؉�F�U�c�����|�{Rq�+����k��!ڢÒp`��y���Ϟ�����
KrF�u{ЊO7j��l/�MXw�kPl��6�Iy�Q�6�V��m���t��j�Q�%�Ѹ�8���U!L��ޘ�\��fvQ�J���e�A��-�1�dM�m�y��l�����������>km�Q��vN�h��;�y	��F�A�L�����.�k:�Ib������m�g[��=���sb۝��(d{޴�\Z�����|l�!軉@#�;����a,���ޕZ�܆4m��_o�v����9�p2f�.@��z&;�������%gvQZFnC�� ��>m�=�)��>�l�����$ӯ#�������s������aOvk����W�� �%���ցpg?�|���CA�~M��;+���jZ.
_�Q�k�f�%Z��b�V��2~�V�v���W����32d�XV��7f��Ȳe�����4�a�|�.Z�z+F�O����k��n����l�b
o�6�V��2	��2]5�Ҭ*����,��\w��Z�4{���L�j�z�[��ߤ�_8?�T��Š�s��C��8���R��rmdГ�s �=�xֱ��'@� �Z�G�Ə��	 �W
���*���5�dGe��&ס-�O����=�{З�O|ݔ��+���������缇��	�0�m69�.�!�c��7 �N�%��`�o(�un�ò{�ౙi+5����}pQO���;*���7�,����rkd�7{b:R3'Cd��ex�K,U5��J�;;��ly���<N�8ѡ�N���&�iM$�iL��Ȯ���p���Z�v���% |�Fу�g�������V���>G82��C�S��>J;E�FAJ"#��;4A�'�j��x��G�������t���u^�pZ��7^բ� *W v.���0L4Ps[~94u\�h��.P�7$F7}ټ�<3����.S�a�^��)Xg��e壗;��9b3x� '�dݨ�Y����D����5zbC����B�KN�˱|�P�@�[�V�U��J��wM��DT�
}��	��ɢI��k���7lcA!ؼ���%������y<O:S��c�����R�A�u��g-5�"5���gJ�����d�N˹�a��/�!4��S�0N*�[o��E"�	�*9-۟!���^j�ƬVH����
�ͳ@W��CVU�@��p2�VS�p�zn�6�}���@낌�:'N��r���lTJ�X������Or�Cg�%������O[i��#	��&��c�8#�
<����N���v�%JQ�چ�6�G���6�4lv<&(�8c���%�x��L���J���h�6Q*@
�[E;/_�H�������;�/�d A`�OȪ�z?E[�5���*e��Զ��q�R�4����y�qV�ߘ
8�|�Ph��[[�k)�g�NɮM���/���Q}f�	�7[ѐ9�׀&��ḥ���������&�-fӰ�n#q�8��!��Oa���( �1f�\�Γ��b����<�M��;t��xU�>͓r�$�Ɋ8��v��y��q��������#�ϳ�9�����n�5�l7��1	�t{}Y��IS��}��g�@�'�Iv��:�{j�u����ѧ�Zb�T=!,)���E3h.����~��`�Y���`�z��k����_�X^�q�I@�Q��������ov
@�$z�rh��;���f���۠2�@#EGާ�P�x�V�#T�����
@�ɓ�V�q����jlL�&wJ�W�yϋ�m�c��CpI�6h���M���-;+D�+���[�3~6���Z�Vj�P�*���P�/���L���Ws������;��o��}ާH1�ţl���Rk��񚝣����4j!��Ֆ�l����G���x�ڇ,|쯴0<�Uq`ʅOq�.	 6�f�׶Cr��ȗ㬪x�Zhg�:?�u����u�R��S6{��~�B����,���]�1�1b��Ե�f��b�qX�Y���	�0d��%L��m�g�#[�D�(̜��g�a?�
�ӣ���	�]������ڦ�@P0 �Eoqw���l�|��q�dl�z<ƺ9ׯ�.�+Wk���V�oȌ���]/n�r�s��l��kj�&�"�@;6�S�\Ƴ�sD�18�?�ݥ�b&?����~����T�(Z��/�;�����]���,����d���sP��1���Ө3Ж��;�"cY���5����,z}R�#�t\4Z���:�����C��@��Yf�wĠ_�~Y�a u`_Zd�dz ��b�����)�x��LJ H���Ε�k���A�]o��5wZ��j�Cn�^�X+hA�N/������Ϲ���f16�c�q��4<iY��=Q�N� ��� i�YuXb@P :yL俾��,�����@�"�\O�~��n[���/{���-�y�D[N4&�H�h��\/h\�b
�Dx=���!-�i2����]Ee��^X��{�u��ý���T1�p�xȤ�m%��ŋ�G� Uَ��3���Q��f2�p��1v͂��@=Y���P��l�ƀ\�����]��ZFp}�Hp0���p/��p��p�Xk�*���ا��Eˬ�:g9<MGȼ�wڇ��n0�k��y� %p��x�Q�����1y�`�y�`�ʭ����r�}��bTvK��4�}��K4�k+��2�>U��v�:���%|��{�ӳ��޳}Do��< 1����z�@�{��h��Ǿ8�=g$켷�����`�h�^����FS5�I�|���*������]�x�O_s}���h�b���Y?4��dB���7�6ױ������7�)i
���;p��*�,M�j<B���eT�;�Kk��ٺ����\��X;�t9V�wV��u��zr��������6��9�|KK*g�^�� d�u�k2��d�,�%�S[�,hL�9����� Xr�i��u���bJ���%�g吀ߚI�l���1��>e���M��	_��픽��`b�Ю�����7o�w��A���O3��� &�P3����f�RH�N=4�S$:�[{��j���t�Fq��谧���ik�R�M�3�X����{�Hv�,�������z9-[S*�;YB9�Mkt�`&��P�WT��[1hW6]G�kV��go��I�l	��鱝�n��'e?wn<g>S�D"@ߊ���;�Z�5��{�g/�*��֕5���/�W���W{���`4���W�"c! @S��fS>�
Je�`y��.Z��y�jך��<K_�F�#��:]YQn�6�� ؘ�v�h�ز`��^�1�c����6�������1�@^;ځn*�o��x���d��CB(��]�No(��IXoe�E�Z)t�G�%7��ت�XE�Zz���u��]�ǩN��g	�t������Ė��[_�ja�{���jPc)� ֲ�@f��O��NX�����5509��se����b�D�)|�
��$5-�ߌ�H��n�יL����Yk>	/�GJ �����l��%��L/��$X���쬓��T�)�ƚ4���y�O�x��O2�q���I��2}�Oa�G��m�<����}��3� 8��^��P� F�#IF���G��Gd�d�nC�9O��9�=�-�g���&�b��&p�F"I��oZ�j]�$)̞�-|y�.�7��gz3+��X�!DgM�r�%
`!��z͸��i�S�ik0�Z�@����Z�I�td���KL᳽��V�U�|��&k�v�Ӂ���?���Ͽ(71����tp�o��Z� �f��Ʀ�Y����-�{�雌A�<�_,"�5��X��aӊ�6� �G}̽������w��-ż�����1��\7��/_���h3�Uw0�SkV,�l��&j)�k�3��Š-��D�K���+Ty��y0ug+q}��O{g�I2������c�q��3�(�R&�7+o`�N��36�-C�0s����Y`9^^�8�"�5�go'�����߷�~�ռ�]_���b6�j����ijj^�m� �̤2����^��&)�;�Fg�
!c^���6�*�B�x
�Dm�6� Jc��JH�Zz�b#` �o�Bh�ǒv������$�Vq�ƐfG2�ǤN=ŕ�Ʉ�w����jc�v�V�'G�
k�Ð9�1;>Z�S���޳g�q|x\��s"��>��*Z=���(G�ɰ���B�� �&{+��;%V̐�߽{�*���*u�m��ǿ�0}�vVe�?aY|�Q���l����y1�k��%������i�~'*h�z��x��9F�/{�@�5�����sQe�mt�Mj<20��[1X�f���~�s瘷��Ƽ2 gۣN	�nx�I!a�ٶ&^�+������c��G�%���	���I�^�1sma�k���[o6�a�� ��w*n�A�啍F�x]�5;��iDy�䱩���H#��mK�6��a��]`��&��@ �`�B�I4���GI3�#LF�'-��V;'����Ao)̋�]X�B}�BP�D0F�'���X�)���&U�*�SU�p����,��g�J�w�z��-`Q��ƂU�[��'���|am=�����C�A�۠�z�P�S�sڎi�@�)mԨ*O�
�L,�~����?���ݻ����G�q���� �
��6z�h9C�qx|(@k_���;����m�ʡQf퍸&гI���Z
N7����)Rm����%і;U��n %��[;V�d����(A�v*U��]^\�]H�������ro�|v`'I��ͭ��i�VE[Լ�siF�O��O���oi�.7������E�Ż��I�G��&�(ߌ�����?7[[ذ79�F�� ޤi �V����2oցq`��`hV��$����^3I ��H�"<1_Й�.1�I��v�s�Ǯ���޶��u���jq@K��V�H4��j�`�H&���:�w�?Վ����'wxv`E�$����̖5O��Xǲ�&�Tu�f�ȳ�Uo뙌&�Bbk��6�!��Vl���ܖ:����� I���k�xk-�����v99�x��9
����&����ek�~R|�c�a �ÿq�<џ'��9;S6��ۤ�i�����Z;�J�h �+)t��>H��b}��hݝ�yCF�ݻG*ƴA��Wj!Ļg�ro nS��
���{�kK�Uc]냅�{���Nk�W<�;0���Tog\z���^K���y��9Q��n,>@?��\�� �T�]ܓh�j�E�����g'��~��[};'I%fW�_i��}�bpe1}Ⱦ���ل�+�7�K�[6�O�F��mf���97��Â�Z�����0���Ĺ�l�֦S�V�,������gg�%�������_jF��so��xp6��O/�v�b��8m&���*權9�[ŷ�w�@���p_�8O��>�&�HmzGs�;9��߇�����nk�x��Z�d�o{�Y݈����_�*����O���o� H�~���ŋ���K�: :^������Ǐ�x.0sG�|vqAƙ쨱�&o�kC�^@�DfZ�6ky�v����Kh�oBi�����*���o��:H���_���":�.���W�э�g��O
����d�|�a���61�@�e�[ ;?C��;_�t�%���O�X�(Z�Aa�"����,���Z�*����Ъ b���rcA�h�&<iF��=��
�WժV6������tQ������7� f��SH �
�Wy�Z=9p��[s�+���&�����A#E�]�oۮ�̾pL�j�G�z�K��-�}�����y���1�ٰgc�hʀtD�W�mh��Z�yy���Y٨M1pی�,VNN.�h�{V��X:<:&2G���������f���\'��k�1ڂW�����UL��:#�I>n��}�����n�7�XF����������95t4�۵��osH���A��
<a<��쉸5l�}�dz�]@�hv&�퐣��G�����������^������n�y<7��r�d6�hF��$�H��=neI�H�.����"��z�����[�����ٳ�@�љ�if�x.�JǍFܣ�D}gc��k� ׅρ�c��LF���8������Q�v/�p�s<<��^V�Z���F�*������s�LZ:��8����Ϲ?6�;�g�w�*�����.��&�D�&#ւ��U�8��.Α�����y��Y�.,��M��wV��BU?�UN�X�6[+�W�U��S�o]mV`��]�o��|��' ���d�[<�&FT��>4�~�΃��-���#+���gO��8�iQ�?���9}����?|�`�$yHd����$m�����p#��t@֏t�H���\ﶦy}.\{�wȩY"]q]`}�|��r�Y��9�TT��Y4CPS�ˎ��G�f���}� ���dJ�����+��c����ҳH��	>+]/�����}@O�3�>��$nY����
�<�4�5u+�I3k���N�&�/�^1�	p��}i��O������^�6��/�d$5?Y��	߱��XYc���>��@7�u��]\�ɴ,����m E
ޜ�4�f�y�*���+�k�u���^@	1E�Y��3�iA�6��Y�	-g�ɞW�ӵ@�N�n� ��,�W�v~���L���m�`���&�L��5��<��D���-5#ޜ�
��iʋ�Pw�Ǐ>.{�3�&#��_��t�W�>�/]����h�l��I>Aڇ�������K�n|��7髯�f�4���Wob�"ۅ1~6�kش�d~[l�� �8sS�'��JTד����h* �M>4�a�˳�@�7�����?���G�h��0�>-��E�װ�s�Λ�	�?��ag�|jj<i�"@�qп݊������ܳW��m	���Ėڷ�C$����k縬��C����*�6��8 ����7���b���ӕL�F��'�۔���t�(��TF��qj� K�N�v���'�}���/�N��Օx�qyB?�X���V�[	>b��~�sq�����t:G��;�wy�K�;�p���Ll�n��v,�=��@���G|�,��žjR�H�G�sX
9�l��f�M�8���To����zC� �K�������R�iƞ�/*:�i���
���̙�5����OM^`ł�4M+-A����0���_��)�}��L�p`������+�žy-f�v\����H�]�?{�\Z��⵶(�f!�Mwp> ��_~���L��%�������)�f��v�s����ٍ1V��'Ĳ@$M6�L�]�L���Ea)s-j^l�6<���g��Ν4Z[��t�th�\��fӳ���i�ܧxi��Q1�֨�D �+���u{��Z�sގ~)*�#��0��)�Y����e��;���z���:��T+���{ɪ!��Go��WTUUm�#�!Z�+�/���3p�0�s��0�u*�o
F^t^��;
�T�!i�5ª\��|t6f���J�}����/���D"��zwj��Ê:0AC��ͥ����c�0:�h��d6� ���kn}�"��~Kg9�Xjg�7�h�Mo�@q:A"U��V}�΀)cCh����/Q��8:����M Г� h�2k/)���'�1`�!��N�rJ��1�w�n$�^Oke"�y���뵁#���b#�J>�zǸ'p�H�P�A�����(�#�,p�5ZLRȡ[��,r��-��B�-�����πQF���W/y�@y��@H�|���Ɛ�(�� ���C�~_��-�����~�aR�h�x������XpP�f��م�z~+�E�^��pXw(}�>z����h��}��û*k~w=�����Bh��=�W�a���q�j��&0@�)�+�/y_}�u��o~�`�k��2A;#�sE�	p�Ym�T3�v�l�@��T�� C|��
��qN��C�ߨ��u�2�j
`�����^����<	��b&�>jgQ�Wu�, %�s$��������#��CX��!$��*���k9�՗smj����:Y�^� ۩��V�܊!���#Ͽ��4 @���?�/^�~�ֻ@�)Z�f=xx�����*�d����k���}���ی�CL�C{�!��X.�ـ�v�}�J�S�ٲ�S"�b ���DYe�ߵ�`\?�[`*�Ý;k��۲���t��LsM�烄�e9?�0V
S
P齯��,}X�nNG��.�����@�е�!�٣"8�8i]��]H'���u�x���/.�=��v<pu6�3LǦ��q� ���1�"
YoK��c���K�&E�&uwdZ�\�\a��+�GqL�+�����@�I�,�ϑ<✻��)H��p.�n�ڄ�$��&���6?q|̺Wq�5�\��V���O>M���O�_����?�۟�˲����i�� �	�g6 ���=+�4�^_�� h�����租}����9�����>��,�����ϒ����#�G=;�$&�������b����q���1Ż�u��~����boT?r~vA�r�zj#���yL5 ��qŦ�`����i<ɀx
ٻ٘Ӳ]�E�Sh��'XIzL���ͯ��8�+�&T��oL*�~�zK^y�oqO&ӛ���⯺�k�����J�l�:�&0���Q�>.��m�)���b��l���N���w�MW�&D^acYP��0���x����ZE��gtxd���/H��)a�x� ��wP��+��Ѥ�r��Y�>�=/}��We=����Q0��~���6nϘ�]l���}��_�����Ů�+�vrT|���H[�S_�s5@c%�`��	��Y�֩����KxL�:�p����ly�4��`ls] 0���$o�o:�����!�v]<7 �� �C��w۞W��1-Y�,�NjoF��5	��uS|��S�Zq�`zN�
�d���aۼ�C��5���a<��������Z=u�1�>|ڈ�0����(�'�.�(
Ft�3GG��v�����ct��>��h��֑��mp�ߙ�)���3e[;A�� OV|�"�ǂ�.���a�۱e�|^��r/ �v�m5p@�ZA��f��Y�l�E\�p�6,�J��S�2#�kΒG��F�����H\�;$8҂���}c@��k��=h��_��"�1�~���~Uք�M�&-6F����E7M��Q�̀NY�
b�,"�FBp�1�Љ���7{�.��\8(�S�(?[�t� ���Y-Y�@���N�TO./�����~:!Q.$�����	��l ;~k#ygl���I��{Wv����1��xE$��9a�%]�}cNI�P����;Ք��+���^���+j,�O��)��u'P�������+M�F���!��µp����ç�:�Q`#�j~]p���W�x�ja¹���6B���'�S��&�e�X��%��p�oH:�n\�N��u��#G�O��)*�C@��,1]N���BaP���v�:3|��O�i�Xq!��7��c�/?OoJ�
���//�������44C�
@���'L��h��/��N��O��r�#Nǻ_KMP ��%��/m��h� '�4�  �o��+�G��5wĤ����-��_��6}��o��Q��L�[�Y$�H�\��j��:���s�����z������hO�=O>�܃�˝����'��
�� �6�Z �.:­�������&�G��� 0���X���W����K;� �O�h�Ob
�!��sj��DT{�V�w��Df�ƺ�����U�j���!h��daB� 	�`c��8��ɂ��q�����`:b��`��ۿ���W%�F���������lS0���OD�f��b�XCxu�/<AY��O�&�]SO�J��3��( ���	E\q�3/{ �	�(đ��2P30g4��u��z�@�`{U9W�]h7H�a#}�r�����O��'}������q�){����`a����D���U��}o��$��_X�5�C��50�_�ev��dyY�zWc/���}T
%���[k���y .F��:��ֲ����+�����HD�qL�m��%��l�p^���$��s��xk'�}�0}�����M�0^q���XMs�V�����<H2��������I	�8?�+�Y�d<)k��~`m@��= ���ѣO���S27�x~X�H�!��C9č`W"���36{zp��শ!�% i�6h�0�1�LKv��@�@a-��N�s1&������$:NL��X;�u�W$�'&����㘮��c�Ŝ��֊A`{��*�Z<	����g����G���t�����BO#��� eB潵456ɴ�d=f��I� {5�lR�Oy�� ���k&��%��O�V0���q���X c_�q�O~�x9l6�m�  ���'ưЯ��uV�4�	6��M���8��������%P�x�ӲN�.>�8����źj'�D���l2w k��3W�6��Zl)b�q�E�oc��ܸ��B��m� !��ݲ_r�Mj��8��E�~��Hs�N{��0։��7km9�θ봓�i��>�dQ��<L�Ҙ�Իn����׀	��'���|0qo�n�Eq������N��6�n�CP��ߝ ޚ��h��E�dc�䜈Aٲի�6�m�k�'����+	K��~�U��Z+�:#mE�ƍM �qP������oB���vCqB��ؗy61z�m���4��[M*�,�Ej�j��g�R���g��t��k ��acT͕M��������kG� c�L[��[�3�#΍���%˷7�5Q��&S2�uV�Kz�Z�M;E�PGH̍��j\s3�i��_�!�",��W_�Wk�����9���n�<�f�,N�'�"Q1Ob�'��+e����D�Rb��D�,�/�ם;�y�GuwYEc���n6�F�jS�C��ɩ�;^y�����K)��l��6�Hc�,��@.���͘j����ؼ�7�y�:���a���5��%���I�lz��[��&p��7Ԥ�ˍ����lĢ�����Ʊ��֗�,)\sٸ�} ��Q�@�L�d(oSU�j
�Z�n
�\��k"��I�B���Y��̟�X�u�j%7�|�����_��+���šql��bm�{��gl���$���f��>&TF3YІ�1�F�D��ϻ�}��p����矑��鏜*�>Sj�&,�瀀	L���
�8�J`þ��P�H{�HV���X7}/�r�#Ǐ�~���W���� o�r�+��S����>{�������~�[
�b����y{��Ф�<�3���ZU�=���1����3SŠY����/J��@����<��G�7*��jӄ3�6z��T���V6�B*�lK 7�k�
�>�\�T��󜂡� ��!|����:�6�vN�r����V+]�:ү�^�B�4	T���'�Nz�4���եck�A =�W����4���G @|�k?�8k0�H�}G:�l��,l���#�U��!A���w�1--`�`R@���p��4!�V�g�)��p*ڹF�"��|]��=eV��6����(b{um��	{F��u����P;�������.R�s`;(�;�a%ݻ�����s1b��4U;E[�O�JUB|��Ӟ(BY�KQ��X���$��ƴ�f�b�zY?��ygi��7�{���Y^�������b�X��V����67?�����F��*�E���W��u�I�z�.���E�{9��k����dP�/.L~��+�R�w�����W�	� �7Q_�:�˃H���K>[�e�#�V �����32���粽��%�����(V'�%w?&���Ç�Q�;HT4Z��� ����aJX:�=����V�����a�7���ɎI����2�L�/�L�[��;)v�����Ǻ>M4��\�`�lg�Q�Mw�=�L����}�z[��9�;-
���
�6B��Л�dj�oن1�}p֦�*&�e$cK�g%w"��D�u�,>Y T����MZ�Z�ќ�X���ٛ�~�3� ����h�ȎقE}cx�+��Si�*��žy��5�	bu$� ?����O��+;.!�{�8�~��p���O��Z���pǅ}C!�჏��r<Li�Ovk߅o�~��"�jsD{�Q8����lB�yb+��/�]`a���\�m�y��������qx 簈������ ò����MP!�+��6�tbЋ��-��H�z����ٶ���^=�ZZ�X��+h�D��۵�f�5�uk�?�/D���>����@�&��w�:�����M�}���Ip�J�Ɋ۲�V��^�+���Y@ݰeI��%�|��`���*O�1�ݵ�&Ӕ"K*C2tp�Z�Iڻ���,����b�Ύ�l��IR,�ZA�u�4!6�*��̏׮�:�oՉ���3����5�民f�,Nn O�?�y%��q�v��v%B�	����+K,�K��P�����\�6h�^���ܫ���H?�"�� yϋ���p6B�|����K(��'��^B�j��H��� �X}��:�띡�S�32�h��_r��D5W����������k���b^m(�8ʉq�VJ&�@���\�BN)�Y�a8h<�!���沘��*��z�����4G%`yp��� �@���;[������Jvm�0s�F�ʁ`�i����k���&�v������Z�8*��"���Ɉ�R}\�'���'.|��\�b�:��*q@�G��Q����1�=���3��]n�d�Γh-Q�}��&�(#;��9�c�V������D�]lJ�hlԺ���Bm�}�����V:&Uzt��������hs9>�0"I���:��~��'Lh�����(�#?:>d�r�*�����j)%�{����t���#E{`���3�Ƨ���"��P1Hp@/F5#&�t��;��A�����.��rQu���EGj3����I{B`�GF:��v{	�W¸��g�ɘCUA$��_�@��<6u���\Pn+AR8�7�/{�mb�`�d���0�1�\U/��a41Ѓ�6 ggm��{�l�CmL)U�����O�{PB��۰^��;��.���nֈU��[Е�4���4�I����<�8=�4�x�.�ӛW;�_f�8.�l�ĭ�p��V{��=�;U�gcda}�PI������v��}�
�K@�i0p���/�۱�����ފA���Ur�d�w1t��W����_�^���(���}2���q`������J�a��3]3�P`Á񃵉sg�M�t��MQ'�%��d�6gت�n0��+�cc��Τ�b��w��f����7��*����A�O'�ﲽ��VJN�l$�+�	�".�.�����M�߫-Mvo�{SL���u�"�~��	��k*�Hɓ�������1j��7���L_�@�����Ȕ�`� ^�NmC�MC�6)$%g��l��Y���,'20)�׶&��_;(����B{��Ï	��I �Cx�kkk���HZ�� �>k�f��n�vΌ%��ׇ=L_~�y��o����$=��ځ����i*����d�]��F16..����	�7ܣG���o��`��X��}��`�w&Dk�!�Қ�')�r��x���s[�]:Y����`�A��'�cN�|D�(�.X8a[D����^k�3�⁇��*>�(G˘b�Lvg2 f���/q&P�ؖ��a���}MS�hN1��/�&=��!�,�Q���d��?98�63��r�ř>z;�y���kV���I��h���?P����=��!��2�e��r_w��±)6���������:��w�� �g�'�65�m���� ءA�~e�lm9b[�>���XL{ܧ��ΥIi~�����&��`7��xp؆@-[r��۳#j]Q�m�}ź�sg��ˋ�}�❦�ac�5��~E����'G��ҷ_Z��I{hkۑ9$�X�> #��DVyc�c*2S#�d |ݸ�Ck�qF\3����kuo8ه�p?�{4�{?!�^�V�:@Ҧ]��nۓ|�z���|N��Ma����ۑ�Q�wo�b���4���]����G��ԯv�h�eS퀆��h����r�,-G��͕@s�`{�{���L�~v��x�VL�ܧYv~xl]צ��8^l1�34�=���i�����'Ο�X��e�"6`c��xL^�O�f|B�ĩm׾>z�����\�bV�D�l0Y<
�|��B��=�����l5��;�G��#�D�c��/>+�Eq���C�էT�1=w��� ?D�|�Ǝ��^Uxb#����6�* �3�J�Zkmr���&R�xٵFֱeb`��de}ओ�N/]Y�(�g�l�(E�$���ݮ]#f���OcB~����q�[�u��B��c3s��`�+�5P	C�.��ђ=C�$��O�&E�]�G����+�`�X=���=Վ���	4p*�&s"	��J�z�G�9��ko��uꪣΣ�_l�����p ��-�a����t�T�?��
$�`�"�s#<�`;c�^��*e:&�)���}O���irD������
���pp�b�x;�N��9��f:���q|���vu#P'S��
�r�&R�{	����� �<hܞZ~ ��`YHN�V���[P�_��x�A�BL�8~����?�L�}%ppa8 ;.�}��C	��	��(�%��\;��oEU��l}���ŅF�	f�T!����ߥ��_�H�؂e�i8��@0��5��k;b�`��\���D��O�Y�oؗ �*���n�ݴ�(&��9jc��H�)DZ��=��_�Bf�H]��rΤ����`�6�m+���k�������bۙ�7%��ӕ�ΰ/�[���U缼��M�Q�kj�v8�F��@�*���d�O-5���Μ4E�	� �J�!�\�5�Y�=L?�1k?�D>P��V�wu\�\Y$~}ɦ֘_�w`��`\'A�=���demL <�;N�ʷo%^y�*����_�8&y�����ި���ue��E���� �0}-���=��ZG�/P"S'/��N���������89�PF�gR�!|�q�H�)l{��g�+z^��a�Q$�&0�Xm�V,{�US�X�M�޽;餜���V�"��ij^�"-ڄ���ی��.<��UP���>���uwTa�dkc6�r_ǝ'з���؛�B�߫ K���`��s��ْa�t��m��@��k6v�d�O*p@�����qL_���m��Ѿ� F%�5�=Ȍ�����A)����
]<o�$�YZM��ho��ڱ�
��-[��#���Q���᯿��I �k*�������7�o��M2���`~��a�'�ѽ��O��ނ�Ů�m��J����=�SR"�=��j�-§�h�^��h�7�.�*�s0������vԐjlZ��Vܮ�'��ؘج/����m��ɟ�\�
0k|w/�%�W_�j	f����҄Ww<��jW�f~l��5�R-�6�|�\�F[�'G"��r}9f�l_�b�k�4 c\F�_^HX�� s��a�UE�������'؂=.��BN�&�_A<����&��w�#��~d�,
^����Z�>k���N/��>^+��,�W�Lqn�7*r��~65ҋk���`S���c"��K<��`��T#��ؚ�v�r��u�V{�Ap}㜭�7GL\�
����]}kq��c[�}����*�#�'��?�L�ǲ �@!֥Զ2[>�8+8U`ǘ��z���]g3����_R�<$+c�Y�)�F��q	�< '��@FKR,�Z^v��=2Κ�[.p����L��&�R���B���1\�f����p�cz#�+�!\�A��h��.�|	�n�������om�kRQ��,~�ۦ~9s��\�a[E��he�����Ćvϭ��"W[�]8��M�X2K�y-\�aF@2�?�|O� �^j��S�cy.�U�޺ooc/HXy^lg�f�>7��)��~����c^�_�\��{��C-0ݔ	��p�ġ����5�8C/#�k~�(Y��W?!�ow�a�hI-8�m���@� ��E�6>q��Ϊ��{ܻ7ϝNУq^v��6����z3c��&j�szt	��L�z;�}M	�l4��ѣ����i��Wk�����av���*�I	���N�N�L�6�PH�,u�	|�����D�P��"����9{{�QѠ�n��'tta_`�5����n�� <��H�G�h�����,b'��C`[�6F�M�]=�Bh��9ˀzQZ�����w�1%��|��R~x=������F�U��̵���[�i��Y �K���Se�YJ}��柸�km�q�{�e�&���̜6>�>� ��|@��C ���7ߔuwG� �d͓7g�1�5J�:����j�Nm+��ҏ?>IO�=%��������sVl5u��1��8_$��1�3�]�̜���"��:$���g;@#(�?�?��&�|��w�G#)�ċM5���mT��Q�Z�5N��'�1����ӟ������������a=R(�B�,6��C5L(|�{v �QuFe����ɌwӶn��̈́�V+�JU������
�g\;�-~HZF8��J-��&֡Wd#�XPL�	s_��lV+���^����kR�߃�}T��k�s��dU}�:�<�U����5q��Xq�3����=�����l�4��^�ml�ʪe$QY+�G0�ZO��,,�?l*Z\��Jq���������{��$΁z���u�.�ML�}C�� K"V �)��ld��5 `�s
�#���5�G@�L0yGf�����e0L�b��?L7�FR�ʒ�u�GG�| t�j�5�RQ�ӕ�q���.\.��b-�c[Ӳt��ג����ۭ����
QI �5/����8������������*Y1���?�'�Ims.</}��3�oV�HN������NQ�#�#9���.�s��dK��}�1����)����b�'��5alN��V�w؉A۶״�S��0C,��L �(����;R1�N��x��4�7oθ�|�	ַ�b�:G ���Ы�'��A7�+ː� �D<����hk�v���+_V�pP`��-�Z�PL��}�i� w�R
�u#`�s���O��q�W���$�D��R���ZX���>������n�>�90�<o1��6��V^|��f:����G�F�i�Dn=�u7K����me#X[���6�	^��+�G��9���2��/��<�p�`�2te �Y+�E���XbwO>yD�/ ��F�Ķ���߂a�k���j�)8KE�SF[	'��-W�	���wb�5�F�
gv��@�q���a�}��{�|'1�<�,��yz����{,��k�d~�/�Lݿ!Ց��i-��kn�:?km��{�8~ �V����@C��d��Т�*H61�֔��>9*ta�!
ԛ!�e��$�{mv��f�\��{	&��r������kD��Ƅ}�i됻���Rl(�� f�us�|g��N���4!�����[�W��b���N�� @��:M uP�B���~�Ԣܚ�Z�BۋԟC6#��R:?`�yKkq�+���y���"[�CZ��w4b�<�h �s517R�%�_Zm�P��7UCp6f���(��L��߮�r�����LҗR�Q��憍�{|#g��s�|�y�k��PD6�o}�^������A��:�]\\�U��141��n�����F3;e�/�x�Zc�O����~J-��]�+��S�ӱ*V�d�>��b���k�6�k���>c������}h)�֞��ЀR��ձ�>�7@�۲ʯqxW���삩p@s�L����3q�#��&΄3s�4��b ������}D�H@�Cr e��U��ij�*���ϘTe��� ���W��R@�� j4��<����{U�7~��}ko��I�j4�w�l��Qӭ]��Y7�~.��.i�f��}���%���g>s
ү)��o�h��EvP���`Lt�-��M�C�.PfԘ�$'�$�ղ����$ת�h� �� v��tru�u�yKc�6�pt�S�8�>}����ҫ��3��A�����U����[^;֨W-�0��b���</^� �
��g � ���a?A�=ֿ�l��5/�(��
R8!�.���ǟ��tz�6=�]������o��p�>b2Bav.r2b��w`F��4�g��0֠'u����Co�rѺ=���_��u��;��,����gG;6���Y�dc�M�0����v�h��CƠ�)IoIm<?��N~8&p�hI;�e�gk���N �[��	>��k����`3�GÑ���J&~�7P����JM_�j�8����_I�ˋ3�C����7����}zY�'�kA�G����0dkI���
��&@.�u0�;���3c�C�%�MÁj2R�1�ǥc��(��P ��3�����ϦQ����,�|$��祉� l�������U�i,��?��K�����~��L?�r&��ٿ�bw��\������WT�<7���'\NS����<���D�f�ψ	xoVX�7�k�����5���b~p��/���)�u�!�14 �	0Q�/�����}B&E�O4!��E��b����g���#cb�"�:���d�,��gU�3'����vBN[d����p�[]6LT����cm����_^p���p����dS���uq�|Ң�B\b�z���+&�a�}���7�
گVS'=�8ݿ�Oʖ��H@��űHL���ǒ�����b�wT�#�������r����Ih�;*v̂y�g*,u<Ꮒ�iZ��+�$�vx
3@2��/4�xc(S[h׹�8ۦ�%k����s�����W��L����~x</��f��
7���� m��/��>�?�N�ʞ>{�^�x��O#)����$���D�k%kg'���ֻ+�aop�A�#�Ft����p���o���Q� _�����G��s��~~�e�%ϸ϶�Mh�-�[.�wʕ��X-��ß5oG���'�1$6�~�U~;��r3�L����~�罅�N8v� !#�q��9Cf��l|��xA� l�i��1�bþR(x�m�b����7�86�|6�^�--(*�Nol�H����q<��%��Q~�����E?�I���D	�Q�4(�4��gz[�>��2(��iĀ�j�U'U9��w)�u��[AV�o3�gg����@������������ըGRq
�Ĳ�Ճ�p[�����Z�����YttD�Ս��s��x��/��[���s�&[^t���vVg�����W_)@�S8����Ƃ	x���:���.Orw����U^��j��R8����/+��Im�=u���|�ϴ�����Si^ӣrW'�,vY�WtB�jK�c�uM���b��2���4AI��g�1��k�*Cr
�uf ل��4n�ã�w:�#N� ���udr�K����#�7tM0.�`;���8T\�{��&�0K�A�,큃��tt"�d�@}�ݑt�?+�v��
�+���i��'�s^�ښ��:��b��^��Gb{��*g]�?{̿�%�Zi���Z3F���B�hq.�غVC�YP��Oٗ�*D���+�`�,����t�Z�J�H�`^�d�yIB��xΩN�R��b����#>}��jTP�AU�U��&�j�ފ���&�&�8ER��!��{xd����	4�����a�=�Na��4�����AG�
D6��U�>��z�������uU''
$?x�Q������A{$��?���#��&Izàf��>Xq�-�cb1h$�;�����,�*��y��	jomh	��X���1��-���^�&�? �h�ߪF/��*�g}�nR��J-��*��H����x�^p9uU3��ʄ��0��hM�3=;�,��ªru�f���M6l���� �� o�G��|6����6*jR�kgTp$�j��cM���<-���6�w�8���LBݗ���0��	L$�872���,������L(� b���J� ��t ��^�r��b��~ Q�sr�����|�E wS��ZK�"���aШ�@v����. ���r�:�a۰�&/���Im�h������92KТ��v-��QX���v�}�Lk�t�g��W|�C?c� ��e}�e�F׃�
p����DVe�6b�
ȳP�If��xׅ�i���d���cС�ks�'���6���CV��j:[mUu��ֲ0�g���x��Z;�{\ϩ�8��2��#�������q-?>y������qK��t6ء��v؉F��������6�m�Z���	���JI,���|K�Z���R?�I7@�em�4x�����כ����}�ncٯǵ�[�`��=$յ�E-��\�'��0gA,��26ml������md��	�����+�:YB%M�.&i��X��m�L�P�d"�M`x�V�s�TI��ْ���t�G�gy�; ����/��vWT�V� �&�9��WMj�=�sf��+	/�,\=�r+����<0|Q �s_���� �������zy4?�A(�A��y �3�LGL��Y|<ju��m�����w��$����G����M�\V�tL��<#_\%���^v�[�җ���m#���ٷ8�O[�Ve�֡�mRc�f�w�k\�m�y;�3u���j�`^'��&�\,O6
Zq�c���kΝ1z�鑖5������r߷��c���� K����x�laW�֦+�v��] �y�,��as�_h�S�����XQ��D���D�{h��,��`����꯮%�v�k��9��zC���
��]Y�äb7Z�#w@�m���e�%��bҰI��Mr�#�|���̔�=Z���_�����H�s���.�Mj\2A� �����|$2���f����n��=X�����P-*,s�w_^}�M��G�Ɔ�գ6��6��Y��VMw%����8�A���t��I��Ԓ�bH���?v;��GV��>���ZM��\�S��?�ރ͎c�̬��-�|F������0���YiV3���msM��c"�n�|�������{��"##N�8Tb2�K	��Χ��S1>�U�N�2q#��"��G:���#������wE1�+Ue
ҍz�eFb�6�_��:%���wy�LW
����UT-�n�^	���%7   ��wU4�wJ��a�e�����wBIU��=���Z
����jC�c��:�T��6Խ�-Z�a5-����$�)r]��[f����}S�Ղ�:��{P�H�����0J�p��β-�QK ��a򨊡�S}_��#��J�ZUq�>���f����;n�u����xR��b���[���(����J��S�t�iOqT-ơO�
�oq��O�/T������q���7<��� ���� �T����C�۶;8\ $
@�?��"�_���{�ǟ~bp
;��	�O�cTg�YI�N㭓�{��~����=۶s����R����u��B��ok���a�o;4��F#0��Zo?9F���?���}&�?2ZWc�Z,�[�߷\NI#нby��l�-C����?�V'v�N��c3���\���*��kW�v{��Ƌ���NŶX��&��5r0'��g@$A�M������R�F�9 �`aR
�W�
�q��%�P�����n�[#8<r��kA�{W�L��t����+�5�5��[SR@	���I��0�O>4�h�33)�T0���NO�ZsF�������kW�+��5%�S?/�<�����ԶZuiݭ�mR[���o2~o?���ç����o/��l.DE�֝�����u�vf��H}�t���DF;u��o���M��V9t�D���+�� <�6@,�%�1a
z?��h���ʭ#��xv~�N_��ˋs�f!� S�#��`�1X �{`�&��<���I8�m��ΗSB�Қ4򻋕tq��c�+�w=�a�`�;|�v+�n��'Ϡ(�D-8F���$1=��ھ�Dk�_����������a�EX��t����sj{I�5%���;b�yz�������ĭ�=.�i�����G�sY�>���g�����P7ٌ��s�c,�ЎRv2�_U�*�D���!���o�b�.Z��	12�-=���)�c����=�φ�X�/�B������SK�f��QE���Iz��U��E����S2� �<}�?�_���%�j�L�	`�l42Ml����Ѳh�ٲ�Ƴ ű�+[��o4mrU Z	������$Ī��V,�3^>QƢc���'��إV��b��WK1�<Cڟ}���ތi�pf���NߊCS�	���@n���߻S�/c)b���X��N)��xR7}���G_*8a��g�oڈ�����cń�Y��b����� �! ƹ|mp��ݼ����|���)q9�C)�����1�>aL�V Q�!�,*>F>�f-��d�y��%sr��="��t��Y�����������(al��ϐI6�욠 �y,�7�g:V+{1�)`e�)�f�-\x�N�y�M�����XTN���%d��2���h���dn��f&5��d�<Ι��?��(��Y��,�x��UǕ����D4b�*�P���^�@kMsl����gK��,��)�m߿s]M1�4{n�v�"��M-`������J��@ _j�J�QPYhh�L���F��^_p2���ή  �6	���_T�*�G�X1uk��HņvQ���3�tⴏ���>},�γ����L<�._'��PYL����h9�YT���f�J��I��eru�&PP`o<$C*�!NW���j�p~
���E�A�Z����C���f�팰��1:�*ک����Ŀ����?1������Uǜ�U�49heD�]�ֺ��W S�1��C9�˟I�*�x������a��СJz�d�����)=O'�������������^��g|���K��Z� R[{Ͻ^j�ۨb��)mӯ�sy]��#���lL$�{�ᭁ�@�~���&�%:�(�8 ��`����P0p`�;~�y�|A�=I[唴��n{y�?qO����o�������A�d�Vz��$�D\����>1��c�=݂�^��c���P�*j�;i��\�݅}G뢫�4�
m���_	��!�9����ꔬ���R�2纳l�9�^�rH�G~��� b��;�h죱������|��mAۃnƽ{w5=�r��n���61�5Fޮz��@�T��M� ۰v��[z���il�F�+P���3 �1;M��C�G�{ϐ�h���q-?��(����_�Ϗ~��ߋ������Ïާ���.�w�p�3�G�Z���[�~AB�sͩs�����N �?�[$C`�A�
ׄ�E8{����J���)aP�+K�g,��V(+j�q���岌�־V���^�{ҝb�:�-@��kŷ�;��hW�]T)�g�WwH+����o��9��4^�	Q�ZT��וuE1�v�~�$/���@�>��ip�f����A�5p�.��e|֒I�b� Nj���i�*�Go���>L�O>�"����/�}��,M���n4B|�)Sx� q� �ɺ�VZ ~��3�����7ļ�)f�-2��X�eI���_-��lgU8�y��_����+�VQ�"� ¤,^(�����ci?���n_~�3O$�=��nF��m0�ۆ���+[�cWFǙ΂b�� �r�{
,2�H�jzm/Ud\W	N(�;�l�}��'l�v���1����;Z��E/�-�8Kܮ�)||ㆀZwƮكN���X,��^��?���Ⓨś��_��>���?|?��g����!:�����̝���+N��YG)�(�=9�����r�`1N�6�v�+����?���b~[==;��şX���(䶍��8̇���i�lw��n
z�����{~~���"4F�������-�G,��Ж�ɏ�}�]�i:g O�t;�������3x,,�\|A�ةE�З��%)��H.˴����]nǢ�t[}�⁦���(T��~�[踴p����<T%��h�P�p
b�����0V�=�_Lm�wc����S��J��ܩ�����y<^4�GJ����լ��M.{���Ώ���E�#�E�k�����d�Ĳ�g<��~cݧ5�����Pr�8�;�u�l�J�c�^^�,ߏ��4e�P�V��t(Wv\�[r�Jr~l����-��MѱS���ֶ2�#��4��=��,��Ӝm��_Q�r��`�o��l���	�l̀]�������E�^q ��tđi-�S�W��l�t�VO0&b��h�ǧYm��M���!�j1RU�'A�������2
.y��g��c�����8��`p��/���~��[4���EN5��I�भ��*�l���d�$��5v�i����9J�T�����l$O���j�Ak���k:��C<��u�l����cz�ˁ���`�t�����㧡N�s2`�؀��J;4� �yL{�� G��ڏ���B��۽1�
�:HK���b$rq�s�f����싛��1���g���/g��>��pB�& :���UP�wv\Cc/��"6T��ra:-�/g�#ןæb��c���XM?[`M���t7n_9>I�����	��b�g���:�uα�S�,�ԙX�J�<�a{y�� Ϟ=#c��Ct�bnĘeh����$I@��RT}�C�4u���=��y�)?|����{�]`ߕ����w) �����?�`ڧ'ܳ?��S��ӗ_}M`�'Pd@�����N�~�
6tT�=��� �bd��M�Y��3Ю:��X.��`����89c��_cy�@'�o>� ;��,O������ݲJ٘6��=�0��,-8�5Ŕ�-��b>H�����Oώ�]�]�GQ�ׯ.Hg�}�Bdu��ڐ<-��M����#ű~ �B���l�74t}�o(�a!�>�UCj1�B����L��fy�<ғ�O�w|�����t9 n�����ʊ �:3=�Id�@���O9��ĺKbC�M�c[������o���wS}xy���rk�<��A�+F�;�>�E>չvdV_��j�������z��3�<W>�WbM�(إ_Wm�)=���a(ɱ���Gu��uxy�qp��7��,�4�\�-�:J�9��l�k���Qw�.�?&�1Q������>��B��zka}�Li���\a��2�qLw��B_��lЀ2���4�h��=g� (q/��uM���|�S6p����h��1Ɩ����z�znHN���*�:�2��	��j����R� �0\�b���u��j_�^�&Ũ��6̶|rH��'gj?�66<o����Q���[/"�{�������ut�3�=�� ����5���Y1��z�%ۜ�dD��1�Dh
��,���H��F�+%��,FIHk�8���p<���]�٤: Eօ��$L���8�,s�Q ���|���t����n{�g�x����b�]��%�g}͖�-�{I-'0�߲�p�~y�܌�Kw��6b�Ȳet_ �ހ]�b׎c���.���v��ZoO��	-���_	�f�q�rW�Uj�K	���Ǐ�  ���/�0���{=�.��E��X谱q���)��>���=9O���bQ��c���T�ʦ��Q|v.yem7�1LىiXur[R��)��V��������y���g��;�RL�Q^��>���A��/��vl���Z��.�?�՚�>'�zZ�����v!�{�O�`�2� _���p����T'EҎ�z���;��ڪ�4�3��1}�a�`1s�JB t�ؽZH�U�^O�%��bm�b��AV&��4ծ�pU��Қ�|sV>���c]��m��Se�7)� �'�)B6��o~Xp��׌�����Y��<�~�<Ο��ï�C����qr�>���0��8vl�Y�h�g�h!N��(�N�X��4mM?��i����င�q�-��6������������u�f}��eS�WV�I ;�3���\\�!.��D^X Ս�,%j��SRH{��p����`�D��gL2�2�>�~:<�p�M����ܻ��@>�Fχ=�M���F���j����꯿��� P��k:{TQ�|�ЛQU���gp48�`E�l�)k��PYGP*+	U�n��㑃.�{����V�^���t��H�]�w�J�gpK�;��U^P��M9�o��n�o��:��U�x��V�~�-(�@᳋�#�W�!٦Q�DԾuE_ O[����j���k�*�C�\�����QSߚD��;��}Л�y�&m[��D��~�����>}��7��~3�������9Xlt�Qf�@X��&KS�p�ٟ���O�`����$��o8:��}o~T�a{�{lH"��u�jC�F�����=&��n+�7��x����'�-$`,}���O>��3�%��?�������5���;��lR�sZk�:~��7�����R�
�����֎::�|b?�[RZ�N$,�Ȫ>���kC�`�a���<i,����`N[}XD�dC �g��B������E�=�ð�ܫ�}Z/F���o`
	lI9X;G㊓�@QO�
V�&ݺ}��y�m꒽|��z7�LM�T��Z[4�+�L<	��b�����m�M��zF�Z��I�\iǃ��j�L��9m��Q$��g�S��,�o���U�����s� �Z�:To�D�2�5bz7�4��Aw�X���)Gk�� ������RX ��� ��"��ՑFR_V�hN>�>��Y@u��>�@ܱ�+���~�&Xms���_%'1��f`q�oj��r� �<����4�B,%Hc�v�iLJZ��Xƚ���Q��)9ɯG@Lg��U��a�Q�,X`�~��6���V^+���<�y����7���v�
&Ŕ{���3�Cg_��vH&�!h:�����b_�Z�C���A����}Rk�aQ�.�=���#$��1��gҊ�f��� j�VJNr��֭��o���3#�#y/I�o���P�v�K��OŦ8=���*�<���y�?��ra{��'c�ǡ�ĕ�#���;���
��+���X�4�y�˔�S�$Yk�z���/v��M��^�E���Hpӻ5#�f5Z\,�H�F�Ū��c�6����	�7�m�U�b�c�jꂉ��>m������ԣ��D�]�'�|�Z���i$���8��ba�� ��˔������ϏuNv7Nk�Z�yK~~vG�Fc�/�\p�Ėj��H���ZS���Ȇ�lf��k�����_ӯ��DK+ٻ�j��D�b�E�.�^i_�)n {�-��9�U
qt�~�y:�o����'1^���.�j����/�ι��;�b�4�`!� ��6�suN*���Y9L�g�~�M�=�6����PD��~�?g��C�@���U���汷�dDL�+CXF�Q��i�� Pƶ4���㹾��cf|L�����P��v�h�2��϶��BK2��~��0��W[����B���S�����>���E2v����^�м���6>�/{:�֡v�d��
�-=Ɍ+�,F���a(b�)��h�,��h!ujM,���y�M#��ZA�Ā`2���}���u��cһr��e]_slW[�/4͢ 4���bg�>�����MiJjZ�X�*��f�GO��< ��Hm�3�U�@~��H5(	 �{k�����y�[�3��i�"���޸JV��|�Omȕ�v�\�Ц�MՋّ���`�v6m2MS�X`렭z��B�u�ld<XH$�h�7�PV��4s���L!�m籈*�j �*�ͬ�W��F��	6	-�b�q�n�� X�D�G�Ȫ����R�?��BL?��Q���-7��r�T�Q�`�ϏA��v��	�������ݶ�� tUմd��s%
�NI03���C��C���w_��}�=8�7އ�tG /X����v�����J_~)�y��)X�M�'[��l�H|����J�:�APH�I�Df��Ň�!����Y;�T�ga�ʶ�D���ŕ�B���֛,\�@	�P�Y<���(�;c:�k�8���f�闰��nI ���?��kz��'�a�����w&���CaT55t���\�O�>��4�/���<��C��G���+b��5���O8 �\;a����ϠD~�js�|�g~������o?L�L��yАU]`��X#�
�=J�~z������7����!�����5
��4�5�������u�NzIF�O=��&WC�bPtEv��U,��*X�t��&X��C�4cBb�,�w@i���+g��%RZa(&U pHnQ1���S��BÅ�� ß�	�̨֪@BL=	ԣ�	�_/�w�G�� ^nX���t��Y�vCz��yzz*M���d�-4�A���L�d9��h�]��lv��"�ov�G�Ƅt_���~S����j)Ը�E�9����#*(ـ�e�?����O�{�~��E:b>�&�����5��m�M
��#p�`��W���v:�Z�75�r �`��A�R��=G�2k0G_�@��fC[ػg>����R�н��w02	ne����-e�c�-�*�8��+�=��[�J�4�Vug4����3���HxeC�h�C�RMX��P����^���w�W��u`L?��Q (2����R�g`�(���%Mޯ��ԇ�z��B���ֽu}P�o��:91�\m�Yi��e��P��~��tf�:�:���[���ւ�I������Ʊ4��t�������G�'~�a��������( ^�">�dc�@S�QhF,5�0�#������Т5�o����ي=F��~��L����N� ߓ� p>P�����V�	8��k"��}_��(t!Ɇ��fK���`p�9�sݐ��Fn �ｷ��G�3�2$Bb _��(�}����fB��'U��k���F|���z��3�C�o�%�.���NOorMYS[��^L1�*��:���)  z����1�����t�K�p> pBA	��@P �mƭ�l)|����Fw���,2b��-�r ��O̘���i��1����T��g@/@�l0���
	�A6Ș��~�RFl���?	a
�15�n���,���OڊIf��C�9V��(bffz��oC��=����D�X��a�T}i
����3_^ؖc=��X�G"'�w����'�0�a��:Y9@��\\e������r��}5�cQ������ƅ�q���ݧ�m���|��3&��K�G[dm3X7+�ĹT������\������Q+�4�x��{��+>�e	�N嚘[_9�X�ҞK�̞m�3�"o���J� �Q�ۺ�6�X^,fT���X�����58��Y����S˲�?��I�~7���R)p��V�G�ixνp<�?v�y>���0�6�i�I(z�GN���P�'�f�A#Zu��1��f�"�;��B:`4�}��;?���}ڬ6�{�����oc��LҰ���1[Y��:G���u�����sYx6@���Z���j�|A�3�D�fi�Q�i�ܺ��Q�������X��Զ�a=��ѿ�K	iJ[���W�L?L�9�M�_Q�}{��42���X'8�Z�%��}/n���[j�A��S ��Af��Z��F��ф��X�L�
J7A����Ѓ���i��:�@�e�CyNu��f��<x1�����\S�=��(�&�v {�|J	�o|9�S  ��}(���<�vҜb��N���׽���js���\R�1���'gg��.ǹ0�N��-���=�ENv�߹�֝�����?d��������糆{���}"� ;�WS�|}��	���˫NaC�	D^�ݻoڼ�����Bb�{�s�g$�ǆ�������� �h+�۳��F0{� P�<���)_�/�k��U���&�����r��[0���N��曯��7݇�1$Lʊ�M���ܘj���_ӗ_~�>��s���������<�ӳc�������NJ���Xg��mH�����j)�nh�8ƃ��Rz��)Ɛ��A'j�`[Ͽ9�����Ǩ,��Uؼ߻���L�h�>�H*q�7���j�_'	�A	`e����B��������d�Ӆ.ҭ��(��@+v�b���x�6<%&�ɯ\M���ĸ�k
6p�v��ܠKsja��Zث�dNA���l�Ï��)&r��b��kᠼM��=H���Z�" �vz���z�����{�h꣠�g��u|���'�� ^�v��&^�9l���L@{�		��~|3���D��+��(T?�]M!J�Ob�4Ez�Qh���/�`���uW&��$bj�FX���z��2ѹ�d(ս]%k+�,;q���3�.����"���r&0����5*V�qi��65�����ϟ�r>�[_P��l�,�M�?8��l�`���[3x�^C�o�� �pZ袜��g v�&��C�r>Yp�>`G&�si�}'!n-�OX�Z�Ǚ~yq���|� 	�� ���i���.}?���S��`��}�q��_���.��Q:{����1�� <ؚh�㭶�/=q���ZTX�z�F��%IW�?��Lb���&T�=&��BL	�XВ3�x��x��`�/����� `g�Q�X��Z\+�6��*�O����$Q� 
���d��:a��1i���r�j$�NbrbL�b�ݗ����m$�J,���s|t�Q�+�b��F17�&ƃC�8O�׽����c\���'�'�|\Z�����˯�=�&;�p��'��7N1ɚ�ץx����v�s|}L�� ◟~���&j�l���a?x~�
��U�SmT"�)4��� ������{y=�LX|F����	ӫ�ؚC��`�k�������%������k�T����<����~���k�(��t�0Ҟ��[�-��f�K�$FS�f�Iyn{c�����1���t�GkJ����@B�S�苩t61���fJ�.g,� #��h��'�)3g�?GKkh�`/7f���j��|:�A܇kcN7ZhT���lՆ>,Eu4�-�Kp�3FL�u�Ea�`�|S���MLP����Q�s�G2 ��&a�<����h��e~]2S*�9ʀR���0(���{h��ա�8ca�j�t��?�i�/����H3{��^N�fࢊ� ^�4�+�u��!p_'ϘjE�o =3�Z��T�ySG��%.>�l����O,�q��x��)�� ���U;�����Ne����^�\����*�XcqSj"ݕ@Ɔ̜�z��jr�X壖��[����ֆ�V��4%�zaND5)���YI��S�9�,��9��΁���>�(����:O^�c�`"(�b�HO�= �c��,����P��A���B�nI��h��)<�<�2U�9���π���W����V�w���b��ݦ�����Ca�ov�����Ӹ�4��(��
۴���*ՓV-U8뺲��3�K�D�p��%j	Fd��C#OeV`'�f;�T�{ ��IW;��g�m}Z����w�Si�����b2)��<Jy���q`#�;RBU���_L����0�B?́T�Dv��@��:�vUm�V�ɷ����?{��c�.���;�Ï�4�`��j|�O�<�4-�#8D�7*� ��ǁ�X �V���a���0��I�X5������Ęc=�o���B�{#���q����Q�c�O�A{' 0$%�^~����O��P��#Q`�0�|6���x��Ӿ�����g�}����Kj��(���:sg��xk{��p�)�\h_b��5 H�CAj$�1UO:N�bU:�2��0v�'c�l��M�]#�!�� �&?a�ͥ'�틀��Kn8k��w��� �iS�WC�t��;;mXܽ{;={~�N���	94�Y�JZ����׺p��6N�8c�O����'_�F�_��������_=I(!"r}���;maN���@���HR࿡���DT4�����h��k�7ȋ5��iK�D2�:�zz?�+�^@ D,�[�D"���	��$�ۘ(2��J灷I�l06!a��$RQ��)�ih�`R��smW��>�����3� ���\�����8�Cۧz�
z0.Su"�̢�4��I9f�����,~w�p��#y�$�Ҋ�8�%d���p�%�ۑҢ5�ZU��k?-���Y��C��G�ťž1:}1��Z=�5_q��m!�h��@�-�`�cpp�qa
_�����K��<|�X$�H�� 	�h\{ @H���p��[|�.&�a������m�8g�$�w�;���0�j?hj(�g�j�A�Fպ��>�������yE�7g3��n������^����+f�$�˾��Q$�5����0ӛ(�Z�>�H*2�8H*Ѯ��1&փ���.�e�K�g�7�맍���~{��ek���M���`�����E���t>��ސa�{�6'g��������ׯ]X��/��`+d��Hq����
^�����Ze1*��21�1 Z%Ѫ��԰�U*f�������I Rqm� �hWj��w`�{0�����=����`Σ%�-�#
0_\�
�19�5��Pl0�`HT���\^S�F������ܷ:�.,����uS������T5��f�Bfi�2P!��\�]���nn�+��8+�񞇱9�\� H����O+������m*�������2�he�;�W�F��_o�>Fl��"��w�n6�%3���xpđY���S��.�	 ��*�{�(�#硭��`Xi��������b��s�\&�9ǎ��v�y_�+��M�9��h�vL�ml��K>NaG7��cH)FZ��1H �UC�x��*���2���9A`�kR��\�r�9�z�n�����_���N�#����ŗoCA:e��v���yܣP0m����v2�o%xڼH� ���h-
�b�E.���`j2\���.�l��&?L-��1K����aP��!��P��h"�/^㲚��쏇���n���I�>�f)�:8`.��z����'l�:5��1���<$H��kd�*�p��������oTfQ��� ���k�ly��� ��Pa����\�p�V)e��N�y{Jh��cZД�r�\.��{�^+"�1*r�k%��kL���b˪G�m�Y£�������Bad�8rv�9��)��54�iR���Fʹ��h�I��8zﰠ>'ocn`�A�QΦ���=�p#�%��di�fQ`#�W�c ���k�/�e��|i�L$�x���Z:6 �0��r`�J�����\1���>f�	�-�uTY?��Qz��t���sW9���g����_�����1��?�o��¦�fA"��������8�X��(H����doUq�8�b�}������OV����Tj��כ `�ܹ��!>L{�E�?��?�/%�I}���Ϟ=e�գǏ���&c�} ��d�~��t-�؁��ȿ��+~�ͷ������B�$a$(�?'���
_���OP[}3["���z���}�F0�=�}��3���1����� �E%�6��dhͶ5�c����������%�(�� l���X�[L�z�!:x��Yn	t"�q�F0��x�����H�ﾞA��hTeR�P��o������A;iw��8V�|�������o�g��AQ��`�h:��+��K���5H.Ѫ_�`�L������rFߺrkc[Ó>jo�m�L.$�Ѣ���{�,L�G�K����]Coa�u1b�e�>gh:��%��'��0�C�ـM�5�Ӗ��D�L͔��6����e�;+����`g�Pܣ��<n9T�e���D唶�H� �� ��:=˳�'��.k�Qp5��CP��̂+ȕ�o��G���M9yk�}*�= 1V����Jo�m#IAuy/���*�/����V�^ui���ޓm�k�)��m1�̿3��-��O&���P,\�ns�r�H1�nSR�6p�/h[��F���K��a^P�b��x����'_�>AM< � ���DM��3�X[�k?����{8�i<�B�=�&�,�~�� ����Xh?��,fi�2�j� + �+��i��J/�u����７��/�����d��I?��>�'~�E�i�E�oMpe�j#W�w�r���r��C��u�|d���}�_���,�e�5D|_cj�t�ߺ}���;I:_��!�S���Xrɒ��戽	�~�g��V@+|�3	�9vS�삅��_N�j�H�G��F�5�����׿������������	O�g���9��b]��Ф�`2E��:;�J��Ȣ�!{r����Ӝj��xRd���?R{�ys�1��??I�|�Yz���2���Ok�> K\ p��鴀�'���|��#�[h�a�'Zъ�gK-)h��lg���<��w���}8�:j��}��!{H�{)����Ia��N�舘�.Og٤������H��Q�
��A�R=��J��$����=�oH{@��9�eg���f�"�������i0�����A���\��*S������3������Zמ�����0�Y�%?�3�*֏b�K�vd��5F�uop�ţ��b�x-
�G'n-��.s�m���4�����!E���)nf��雫����?չE��fPς����f���{zfS��X��?R�t��hg����q}�I�~�o��e��m����o���(�GП]��%��Cٙؐma�!�������@N��j, �r4�ю�LO;��BF��*����W���{�#��Tc�Xt自��o�<�����/٨�XuYQ�q�C��dVl^��U�Ѵ�Ӗ���t��.$��>ZR,�iTD2�Dp�Ѡg?u҈�ׂ�|&h�cq��@c� WE�R�sB �?Ȟ�E_=�Q�W���U��d�t;J�޼N�O���np���NZ�|Ŝ�pzɥ�жt�����WL�_L4Z��@�������se��J�zG��$���X Za\�u}��MZP������%�SAiVIv|�q�+K#��-Z>�99�����������ÍwL�&8�1�yR=Ģ�Thɴ���rht���N�0x"����n��jz����S�Ql���Yeh�o�k����K��?XC$�2I� -�{E+�o0,0r��Ng���N��f
~��\�������������{��t��#����t�05���XM �Z��}2Y��nȾ��1陠�1Y0� ��D������<0X��_�SbgfN{�v{� �d	�.<�^��A�n����q2Yw�ϧ���`��	G�~�F�Ï?�����r*��_�X� 9&��H8��OL` �� ���l'�q���͎yp�O�g�o$��� ��1�[����0kN��E��;4C�i���R���{�;���k{�uֈ�Π-�5���`��~_��dK z�oT'њ��]��]� �����`��]Lg�K��S�|����-f���ƸJU{zN��L���+�:���c1�FUc�� ���+������[4�V�e�!����\{�S���ۣJ>k����������̢x�+W��Z�r�K�XE(�Ť"��^9P?�ȹ��_N��y�P���s�6�hz�`j��^�����,��D�p�� ��\��Q���T|S��z6���
螪��|�J��n��-2F�v����[1?O�r���:Ì�;��8l�eݜD��|^��ރ"�%ޙIE3{�M-v<�G�3c:]�;&J[�ȸ�JUZ��ʢ��zB�ȉ��`�~��6h�D=��@VZ�-e��]�����-�2	;!B��X�|�s����s�M��m��G�Ϟ���� `6��hJ�M����ĲS%h �/��?#��(�\c���>��zO�#�9U�AĀL, pL����:b�"r<��j�!�M^��	�����-]H��]
1rU�[�
��抭�2m���[��RV�Q☱؞�^Z�F��RĤ�^��"����IP�T y68[.��a��r	�Rd"e�4���l��B�Dv�*���`fRTv?k���$��}��ƞC1
~~}�f[����L|!��8�{	6���j�A��>V܀�P�(�k�^V�R��\ '�-Z�O��l<澄Z$m���}����=Oq�����-�x��L{m�Gd�-�3P�E� 1�H|��������f�Hk��31�\#fcK#.bh��N.��ޗ�ah��S�"���-�:]%4��l�&�Ԧh��n�ƌS��
{�DF��.9erIqo��R�8�ߏiw�{ ����*� ��a���"��p�@��t���⥽'���ľ��85A�9��A8�f�nͮ �o	�bG������~������p�
�F�A����8���?��E��O�8��y����	�\�ԏZ�
�SN�v{�A �a[أ!=�~&6ɶ�(͸�l��yS{jA�N-�c�kz[c3�t��W����H�{G����}�kC��k�9cՃ�=�Yl��:V'N9s"����sb"��}��[�w���Xj�ZTvpE��,@JU�SO0��wЊUh�I�or�Iv������ �}�z:`�O>/�R$m�"�Stm���)�V�KwL)��nr]� qsp':�z@)��k���J������������d��>F��� �A��;�XM;-��<�� ��v[t{T�Ut8}���`��A6��-b`s�n�rx�(����)a;�}J�~4���Ǒwٓ�$sO� �
:�ݠw�J���T4ԟ七��O����E����ӄ���s
zl*�
�7�?�\�:� �a5T��W�Oe��͓}P� ]t�X�nt_��4h�S$O�W��(&����tY99!ɬ�Q#� �8z����_��Q��E4M� ����gU������)	�������_� ��~��g���f���C���O8E�b �`v	
=.�㑝�߂9�V��,>UhaG���N��Æ��M���MgKU���y4}6��Q�B�[�S�1�d:r�}�`���Ĵ,L�"{b�޸���է���6��th�-����Q�d� =��X$�&������a��䊁���m�L��q�4��,RFO0Y�`v�=�P�7��5�/ՃH�#y�>�&�O����QEUb����_x�Q�IX�d x�`2�1��;�E%y1� X[�F�m� H����?��:$�,L���O���\^�N�ځ � �:׮��#P�Q��u���hbOq"�fcx��{���KS�s	�İۗq�L�{��j�	4>���%�޻]-*�|'�ló�b��/G��hM�s<�� Wq��d/hZS2��l'�����,�5$��v'A,V
�Y,-mb�������/h3��1� �����Ѣ=(�JMc�:�T�q��<��ρW_�ݕ��V`$���uML�:d����R�QU�&�L�s�N��q��bXD$��K��- ͝�K�C/�s"E��ni):P�>���&Ey����6�N�ɷ�f,�e�P֟0}��[������זV#��pz����1D��j��,��f��{�έ �^�0e2�:@0%ٮ�@���T}݉h��^K~J�}�E�{&mA����kW��MxN-bN����q�6���B�����b�+2�vL�##q��@���7kMJ�L}_ز�����c�t�����q�%�u� ��4ϊG˝��m	�\�ӭ��A׭w��@��籠�9 ��n�/{�NqS�:�K>O������S�ͤw�8��)F�ĵ�'mun�P���� 8c�7���%�10x[qr����2�3d(��.�3S�$�. _�K�D�ij�UirV��-2H'A��"W ��oc����\c 9j����#(4�O���<�)}��W����g1_�F�A��a(�,*��kl�{(I�m_���=�9 N�Ϩ���+���g�y�]th�Ƭ��}Zc�
|�'N��m��
�dWJj"��R�Fk��!7;�iFw�s"Q��#3��s�f��,t��|?&S~zi�V�Ft̇�D�轮�q��(~�� �ÿ���<??R���|+�xm��(���5N��9��o	����G��)�Υ�:P���
 m<I�2�`�E�}��20"'�G�*�]p+�����}o�e^��q>1�D;�m�]�M�2��{ᚤ�� �d�~E��5�b��=a��I.�ľԱv �m�U���F�5z��8ke��^E;�0$�>�b����]|t�x��A���������)����me�;&F?eY#}-��c#��8N�_k2��7�+�1Y!B8��
� ʍ����N�|�j��x��#��G�S�S;k�����ca�@ء�"�׺�PҾ��)qa�GD.���<�P�8����wy���m
��ݾV5�� d�9?}��kp`�W�?�����@��;�@_�ѕOc���FIǨ�@�e4a���>�08�=�:&�y�{K%�\S��V������+	�Fe���s��{|�{�֑�o��r�����r$Č��D:�Nǹ�
.��K�_S	�m�Č�fg��-�?ݯ��qwn��ѫ�}�=���´�&3A��߮pH�J׬)�U�HFzӿ5�lGf��[���u����%^�*�c�g�>��h��Umғ) AO8l�	޴/?�����W_�G?>b��v`3�i܂�ɠg�c��h��޴M.1C��*�/^�i��+Z6�_�>K?N����c&���RH����T�W��۹ڂq���v��Dk�DU�02QPe�1=��7��@ s�C��4� l��g��\S*��X�e��ڴ� q��_�)�C^�ᾰK"����ms�x��	�&L�RA��5v�H��zg�� (�4 ���'��4ņ`�H��� ��	-)iԨ��W~��{��*� ��Z�x�_�$M�E��|_9=����$���C<_�fL�ƕ�1��DԱ?�{vm\Y��e\�� �L2W��%�N)DPŀ8�D�ɞ>����m�����&:�	�T�Rn�ϛ"N�rpg���ֲ��0%6��إ5B䱊'g�K
�co�ຏ��h�Y�̢�`�^0i�pe�	���Pt�j�,L�����2����;��f���Э7�j�
��)��&ĳ`?��敵4��� ��s�?ΘB������̖-�#�3[�眒� s��-ߵLق�����c�Q���i��j����-
�O��t�3p����-�Dנ�^T�MC�/�+7��p��0�|��O�����Z��|�Ai ;` ����ݷ�	�|���t�&;n��s.�?�����駟�������y���L�z�M�	K`�������>����dͽ��;���A��=�����4��ؖ�N{�� ��6��)���5�m[j�V�� �c����g ~�U�y��&FE�	���2;)�(b�S.�Z
�Q�h]��Z������[(�EQ#B��r�}��I��b�Px�E:����ա�σ}�l�m(�^�o�ϖ=� 2� f�)������r��@�!kX�`�" ����74�bʜ�u��z��j�l��kG�~:�Q�Y,�ꞽ~���"�I�*�n�����v����p��ѱ�g��8W�7Վ�)���
�_ޙH����Y�5�/�D�z33	dnT�Ѱ�.���%��Gq�`�=� �&Z��v(v����&K/�M������uأ�Mk���ޣ����tc(��Nvӌ�@��b�����m�Z�5���3��ڃ��ǌ/�l8rsY�-y<�+�z��g�� LZ��b���W/��<�7��y� �����9���.C��:���l
����:o�}!WEl+Y�=������lW�1	�7��vBȡ�\���U�ǌg�7q�F���������c���HɆ�����󣞣� ��X�f�Ĕ��G�$:�r?�gn2�y��8s��&Tjڱb�Tl;ٷ�}�A1�z����o�C��D��й�/;dq)�,�I3�D"����ZԶ����4����1��z���3:�𡳟Uw������ڕq�T�����ڂ�O���8Mh�)Uy&x�!G܋d� -S�ު���cbK�R��}���[^��ߺ_��Rei�ܦ��b������98��&�l8]!z*�R\XJ�M��FJ77�X#���X�6�D�Z��ՠd�{�c�i,�f�����o��>��U����N�����4l:��� H/�0\xI�aj~i5l�b�׫�F1l3|���LI��!������R$F��l�l��U� )�%���x���_���M�	��w�5d`�]�D���%�ˡ��r����/,Jl0U��!�T��\]Z&*8�	���&{������vz�<���z�mG/َ� * ��~|�~z��Gd��8!����|8\>��O�w���^��4���q��`�:.���d-��ٚՆ�}�r^��>�k@��)j�p+Ɠ6��B��
P�V���D�Eb���)�t}��W%a�^I�EP��
���t������6)Ÿbl�6/��ɲ�{�.�Sr��'�gn������dg����
�a���ş��W�x�S#Ӭ Jo���ԉ�Ji�-p:[WfJ
+IAj���'! � ���@�=�IŖ	341���n�A��U���s�JD��C�������kW���O>����$�.x��/��D��ƀ��=���!t�����
D��-�]k��R�66�?���ߘe����Ӿ�o��������-��&���7���"��u"!��)���H��#T7[ǚT��s��x�:�d�@ ��@�2]#@ b�O�O;��m(N_�9�(]�Ƅ��گ0J� �s��t`l��k�q;�5 hʞ�M�+����Bgg��c	�􏟘�yPm.�MS�{U+hv���u���zM �<�V'�e�Y!��p�*�W�dp�����ҰY���[T�3�fQ��������p��[�O�M�%���J����!�������b��%&����]?���c�M`֚p�^�zŶaXK�A�4�٦�2�E�`�iZP�Ҥ9�2������ɧ�P����O���a����	�@0SLǚl
�#�Ap:��}�6���Y-�&��U���5�S�D+�b�*\˖�,���	�VU�C�V�)��b���"��e+ a礼2Z��.V���y����)�ӱ�|R]� Wk���m��Ω�
�lax԰��V���D՛��f���0��������[��9�(�g4N9�;�/~,q�`�BK, 1��ҥܰ%���׌[`�bC�=�*�%XZ-k��.XXQq�>A=�j0�Yd^�ueN��YS�z�4�U��z���o`�tu5R��//�\R$�~��[�n���O�� �p��� )�I�{��*:	عf�U�y�!c�[$;ǆ��Y�89	���P�4j�m�XS�e�����})�Ӳ �Ԇ��s3����L$Ii��.B$�9�����YP<
V��I�-�%�2�O�
�P�eC��PA<-��G�-�6d���+�ԁ���6y�S�j�2�=��h��C��im�Gbe�5�8rm�P����+��O���O�� d�.&�"���r�B,��t�S������GE4�d*ʡ]�J��ɷIp\�3z�M�&lt;�.2��G�����c� �![���o˟'M�})~�� 6�;.Ur(篁�������PcȟD;�S3
�!�b��4l�3<���]rX�����h38�#�V�"C)����`�?�%�ݛ����?u����R��^�EE��Fn���V�sA�R�P�~?R���4�����Q�vW"H,R�U�T8gѨ���]�i��sv�8��_�C=�k��0�N��S����(�Ov��ʼ"j��C��庄�	:U�VP��aÃ�D��"�'���܂��5��cLG�?1)��ȼ]Wd�X����G�ثJl�;�EDb{�*&`ݚ��&ǁ���cjU��s$� %�Tl��/$Fpd���(������IA�V ǥW��-r�@%���e��l%�|rE�*Ϟk����eH���2T�����,FOe�C�xC:�X�&<���Xe��fp��͌6@j	�𬊶��$Ũ�ʥJA��{8����x��mrJC��4
PD�
#и��b����/��:�k��b���Ӕ?I��>���D��'$H�њ��aO�҆��K��<p�h��$h'ة�`�:P�k�����V��<�9���6��3@A�����j{|]���_	>��}����u���<mM���e�P!�TTb��ɲ3�)ڡ���g�s�}��)�(�3Av+���\�s@�I'���͖u�}�|���U�w�2*;>���5���6\_��&3��}�H�𵱾 ��^U#��!@�ߡ������CR|��P������D��,��Drk�2�B�֔�����%@ �9LL�ZØ�O������gM~��h/y�1�_.L��.4�_� q�F5T $����}��[�v[�Q����0@���薍F�+!�`4����pF�Zsq)Wd�)��D8OIk�yp�:[���T϶������w��!~PX���K���3���x�(��jte�t��q�T��hK�3]�1*�B��Vl����yjZ�;�koH��CsI�bE`� ��ֈ��h�>���������:NӝRo"��s%���Z�q�f<�Z���PD5����{9�gaRXJdk�[�1�a:/pn1۩m���hQ��Ư�����<{�Ki]�ؾ�	*�dŮ�eN{\c]�kV+(D$#g��Ea�[L�Ox�� �9N�����E�x>c�|t՟�]2N. T�%j����$��^�
���ԜBB�]���>>��L�N���w�|�=��\7�<#&����XNMM(��@V�df���y v6bg!�6?%���eJ�5��%� ���~�ٙ�	:_�|߉ImL����=6�`OR[r��w�y�g�	mJ���eB�&@��aG:������:d��{�fd����d�h����g�����������c� �bM�|dK�&��4^��;��v����ǡ��{s�W�ΫZ �6�,D���/76��c��/����o\B�%?�4e�$��!���z�@w �߉�9�Z�G��ۘ�9�&=��ƀ�
f��n;D{yiͬx?o�*��E�($V]�� 0|��V<�&&����.���w�g-%�+2���f��
[iHY����H����4�������?��A.��\�3D���^��y��7� ����d�����o���<��(�U��4	�K%����P�:{�B������0�USh{Ǻ��*Ǵ5o�5'��9����9}f����R�nZ�o_�_�̗Z�u����5�Zܰ��\T*D��|(����p7[:'��&6��H�F��زgu�1���[�u���z��CR���ܓ�c�v]_ϪfN�,�$��3,��4c�5U�+�H��d�������x�/#�b�C��<����HDhC9�MI�[�8٠�8땦A���ִ}�ؠ¹5ݘVǢ��ac:�%Z�E�4 ���T�Vj;b�SI^'=��c�S|h������
J�	��`�y�h���4�|Ÿ�0�>N��z�ꖒ��4)*>-^��Q�y��0�B����[}ٍ�5�4cl�J�g�D��� >�p7sz�N�X<޴���O��`ԆRU�-w{3Ś����^t�EK�tz��8-T�8v��+Z����L?�����^v0]{�kL�����t(�DK*
�*�x�>@����O4�2��&K�׋��_^^yJ�`g�,φuY��(v<��5����PeU����x\\'�%*|&�Ҳ2J����d��+��BUwr/� A�V�e�]�B[^h�з��ȉH;�H�w[���9(��7�<��kkpSؐS�C|?�(�I-}l��ΆvQO=�a�0f?PYhDcM//7�y��6�{��E� 3w +Q����n�b��~���Orٔ�%k�H��8;WX^M���_�7�"��9��-�5|������@�V�ox�ZE�� �3���_�/�Ma��`���g�2��s=Z4�+��=�驉�ji-a� �zc�:/�Z��;��!qB��.Z$z(��MCG5��*�Z
|����(߹Lց�ɥ��m����]���#��Z��������;��?I@���+�C [
؂9AU.�Sρ�4.��� �T 8���;K���)�]���WɈ0#{x�6��'.��wLv ��V��p6nQ���v_�|[� ��f�:��LA\�'xfoM�L��f��a��:[����GMƛ�|N�4#7l,4�;��4��2��U`O}A��gz���K��>��?x{��@�����dv�3�ﾧ�=D�� �^	+�`fG�A;[0d���]��6�G8�z_gd�ܽ{{Z��le@�Ժ58,����,�G�S��J�/���T�:�<c��@܁��9K���.�c�S��Y�2�$3����0�`�o�d�~�����W}�z�d��?Ѕذ$S��d�<E X���v:	�g�#����I!�׷Z��ra��Db&���9	��<ز�#�*Lj��Ș���thCd�cdLE���V�[dɁ�����&�b�	�$��b`��i�b:cy��lBIr��^_k�	ځ5l�t 9lD�.�ܹ���֎Vµ�Ͼz��^[% �f��j��t&Ϙ	ź~'���_h�9���𹙅ޝ�A�	Γi����5}j������]�.Fڄ�.�V��,h�А.\�he;Ѳ3�Uoӗ>���(X7
��3c(�U���s2Ƌ�ec��/�Atdo�,(�T ���׼(�m\�kF1lg���ǌ�s&P��F1-����tux�� �q�y7�]�7j�^�Y���1��O�Vt�UĹ��?A����n?M5ƞ)�v�Ȼ��<;ek#�
�'�_� ��G ~��7��9׻{� �^�E�;v�1���'-�ץ9��j�E0}cx�t������ɓ��:D�%4��='�6d���t�w�j>�<4 ���7�[6|�&��Ky��%pi,��ܲ���~�矜8g*���;�O�W\ܡ�D��m7S ?*Y,�����8�@H��p;�'
<^OFq̾�H��]�6D�lg� �,��I��Ρ`�}����9���нd�׎1��̀V��:G�O����X��1ſ;�ͮ��Ұ*�%�2z:�
\�v��|gKV�@;�h�۷ϙ\5�"�FYI	��Eh�l��1	Y�"�AM5`ns�%FϢ�N��J�5�cB!%��;�Z�tˏ+u�$��h�Z;���S�����,�����cyq*���$�M�X���yP$Y}�����Is9 �`�ǿ�`��e�͉L�����z���4��f�>��pB�i����A�	8uP=O�'h@�FK*�8l�P?e�*C����`��G�i�wn�M�v� )�?�L:�ό�p[k���*O g$�����3z}E_�-�@;�+:2a�?efF���@�	�`�Z (C�����=P�S��#�����A�*��y:<�c�ֈŚ���:�\c�!>�+��s[?&�%��3\	�@���h���Y�[�����H�F�Z�}l� i	���!:
��)l�����C"�zz9�n�)�=8ֺ0ʓ"��d�u��:�.�h۸�A�r��TA��Ƭ��w�ә��d�l�C�
Z`!VI��m~�c�I����
���W�o�,����%�ĭ>�� H�M+k���x��ȁ]�r᳌2XW����!]$����/L��Z�=��"�,%�ۊM��>���Zm��1w�k��'�V�`!H��4����B��:����]L�9�|�2G��\����L ���#�����Z��g��r6'z����������N�S���
#�gg�K�!�Zx�$3ޓ�.*��}�7�fQ��P�ݸH�?c��[�$��w�����SP��~������k��F�V���@��sut�nk���A�`������^ʒ{��#j��E��ha(��cr���a�g��'S�b�	שU�������?��@h��ޣ�R����0@/Oa�	J`��2����L�s�65"�K�{j��_j�#�Bl�� �}@��Gu�]�/l8�s%�ci�������<ynL.���?�#�
��\}�a��f�Q�$��R>+-"�����^���v�3����{���w�=�.���}~g�+Z6m�p�v�}�G.��y"}H��dx}�b_u�BF�mCWJ,�c
ף�n��o��;w�6����ݷ쓳� CW����~���hork1��mF{:l�h��I���,��{hB�^��x�hoFQ�x��1�5J �m]�i�}j|������_��`���9j�
v�Xډ��u��f��% � 
�?Y�B��^�FM8�z/�J�gkO��M3ߜ�U�dq\|5�QbĎ*�dN9�}5[v1hL�*E{v�+K�Gw#)�#Yk˵� �IǦ���,m�`�� "��d��`.�DK�<��K��G��Lm��]���:���E��&�d�"
����?��=J��<!_���76�K��!���S�N�O���Á����9[?+|��ț���?���J�D�nafnf!3b&�x[������c
PF $�S��!{ڰ���H�5��8b
?����d-�Ƴ����γ��U��<��o���7�f�N}��)l�hR9$����Oz[��f:0yQ/�k<VG��B��1iaQ��,�W�M�����	�#$?8T;1;H�73hdoc蟘Ӫ�"%Ò�h��E����X�рo�:��,̑�54�3}<�rs�$1�%,[M4����7uW'O�d�#�`)�}��
�I>���w��^�0@�E�)�<4M�u����� ����hP�`[��% �ڂ�sY(z���K_[������
O$ iQ@;Y��&�8�!��瓻�6�&�ud1є��pP����,���7���x���8���|ܤYL�80�r��pS��Ѷ,��x�B$UbClhûY��o;vXGަ�=p9Htw�x^��"�!�7�	��Ɵ���r4wk��H0,��� �**Y??yw��wx����]� �)`����y��azkr��ca�P�A6�������i��<�/�N�j�� T^I��6�k��p.y2@��⾚�0���$\K<�x>|�T�����3Կa,������8VM�J1��)&7���u��9w6���@�簎�*�pX�}��j`�7�#t�����Ej��lan.��KL��e�:�:��i�?�
v<�6>�հ�`�A�����x Z@��(l��*��l�m��<n/{3.?���������~�>���� �ɮ�LA�)ڇ�O�MB�s]�M�ޡ�;����AyL0�QG[*��E�� ���'��|���`�hH>+�ԗJ��:���\^�"X�s���$�H���C_�1BV��C��-����T�xB�8�4cD< 7<�Wl�D��%H��^��dR��7���7������+��?����U��69x���{�f3:��b� �f�B�7ǩ]J�L���[���i�B0�?�^��@`�}�Eg��>�Vgg��oa���:��o��f�o��ۂR��"��n���yG-�ɾC�UC��G�[�?Ă� 3���	��3�n�u0Gb�Q�݌=�u����F��dJ8������w�~GPLN�t����c(�1�)����g��#::^1�{
�:�P�i3�#j��4)1Z�z1Lt0�z'�m9�dc�%ْؙ�����ĉLO�6�:%bFb<��Zivq�6ۑ��S|�Гwӿ^�joIc���:^�C��A���BzC[YQ�s�ٖ�&�ܒ�h�[ ��C�Z��hＸ*�?/v">��8�lEa�+��Cx��B�ڠ�. �m<�BI��R���\iD9�^�� �Bq���X�I��)Xah�s�������/�H?�,`�_�i��^ �%�L���d�]]nXP[.3�ʝ;��cяݢʈm��d�$�3��=���
�n_s�b����.�Ǳ&����v�(���֧�{��5�Cتb�5ǟ�(�v]�8�
q��Ps[�~��ق�i��ߑ?���{��Q`!�W����T�S碭Ӱ �����l�Y�! ���"�&Th�"/�]���j�Z�	��0�ƿ���h�+��F���f; ��~Lߛ		�2�a��G\��D����s!���
��۝O��޻�2.�w��l���Y1�΢�d���/��/>�A�b�/�_�8�Ml:�Ŀ�"ydK{4n�=�0�����!%S��Q!#��<��L�;퉦�D��bn�D�rP���U@�Qw�w�-�y����Z�?��ps�b�)R7���sQ�eem(��NʨZ�+�E�Ӟi�@,
c*G�@D��ۺ�a,�eTQIa��N��2E��ta� �E,KX��Qa-�]�@�GWI��ƇcJ�U��.P�p���}ݬ��C#�`������p,�n�����yd;���E�'��r�c��0l��K����sbb�ݻÊ,(ۜHd�	d����k�^m,�\�����;Ø(U�7��XÀOK;ן0�6�F���3�M���`%ς7��S'���
���9y��N�����|��y�1�R �3͒��oK��[���!�Ό��w� 6w�AI��.]-��Ĩt�(��ih1�
05�}�b����������!Q�d���`�����G�8%b{8l��۴VN�8��&��K�Y�s�t���@�����7�� <b\�|��Wm�3tn�{W�:�o��F������R<��'T{cQZ�ֺ�"Х����g��B���3�v�M7>H��B|: �D5%��l��fb�$�X�3�kw�䈠x��jon�t��/o},v����;[C���V�@4	�(	������(¯NN�#�`�,����:i�d�߻���7�^�o���Y-��7�5&�����ˤI����"��(�Y�;�#��oڒ����_H*.=���^Hg�F�i�܌@%�=�L��͔�"q����_�=K��^�4�`�q/'�H�L"�V�#�]6i�Ho�,Z1<��z�׊g´��#$^'|f�^�����cJTu��k,{���XmM���c����^���Ş��[��M�N$��D+N�!������,��c"	E\���V�m����uU�Tq��/8ysp��fl�9�D�soO�5@��)�G">���s2� �R  �L!��3��q7��bQb6@��RJs==��f�̦��������k �P���=�l��ϧ=��5��;d�^�y��)ϟ��}h#q�����2�BLљ͓JL��N�j��	۰�N���j�+�#���s����i6��V���6�`N�m!ϓ�X�W�;b�9��(%pȵ2>���}m	��j	�E�iU��S�CVO^�XuG�@�i;���s��<��͓�
4�u�h����f1���y�H���Y{t���dVM6�/�k�jY�m`=ĸo��!���w1�w@����i��&M����X���u����,����{�6;��H4"3�RPXzwRsGҝ{����=^��O"9j�6[�Pu�̈�f�砀n��7G*�Q�:Kf�������_��\(���p�|k��=9b�o��u=���,�!=�z<�O����K�~[c*����h�غ/��-��{\@�:ʤ����������l-Nx���`u����ALv0Cq%�\�#9�@�e@FW�s6_:��^~dMwkM�4��f�2/���m6������"��b�5 ��n�B�qrF6�%]:��#=��L�a��������n5�����dxh����c��9Dv�^zo�;M^�u��ͮ�������U�� �d��^�{?��9��D���s��b�Js��&�5;��A����z�x��"�Z��V�;��;3Vj5(ܤx�L'S.���u��B��In��.�G�ʻ:F|��c�MMʷ�U<����i��{e��z��p3�Lp�1���%Zx��+��R��19�b{P�Xbf+&���>�\h �Cr	�P�}���E)B�%k��>�w	��	�1�;�õ�sa���}�7�(�g�<��L�-IN��9����\�˅��b��yJ��bY��}XlLLdHEp��9��h��G;a��z��16ݧ�>�}�4|2�yq!�~X�ȭ��hi�їw�6�Pۨ�#��&'ʫ�&��(�v����dTk�����Z�B��-a��;�6$f��Z,�:�.��]yէ�%�����`	��-�齹�(�}�x���#7 �%}�XFM����%E�{DA�ĝ� @�<�2E�>��S�EwUg���y����,ܞ>�
��/����,Z��ǎ�\�p�d���>'�?����TV����Z�j�CDylA����˞���nwj�̻�X/Hܦ����;�b�)��	>b`��� �)�6�f�I�7X����=�^	�K��3�@`�31��~��'���Y�℥��Aa�� ��'}�KLB��bVx��}��m� �m�*�Y���p��>4#I���3��k���k�<�qX�B��d3Q��>= ����y�撯I�>�(&��+��X����1@���\(��%�ng�ȵN׮�$©Hj�V������]�b�H���Ѻ���mɠAB�oA,8XX�(^ގoik˙��WL���R�Q������U�=~�$u��Ux��uX�	�؋q2�L���L8(���$�'��O���l"��l�/�$dv��ļ7�.��v;R��l\���^
{��ek���\���#VQRv�=o������FW�PaO�r�} Q����c'E|�c��u]�N��ܔ
���7�S.���d\��������̺]�K�%O���.�5�f�;�a��<Vа��kh�0Jc�ƒJh�<)S�1Sw>�*�YO ��푵2�:�2@����E?�Х.:e��ac�3MGĻy�����nnߑ
�_�\���ݼ_�'����]�B ���c9 
f�2h4p�c�`�,�R8�50� �_�ی�;\/-�!v ����8	�Fg>���ߝ1��u��@�{��{���5����I��sy���H[P��i, �{ �bl�j�*:���zE,8��N���Ӹ33�(P
��Ks{`���r�^��!G�У�=�q*g�g����Y 2�M�Fssc�8�h��ЂD��5�H;�������Z����Lsl^�g�2���	�j�T �
�����ҷ�lb|��ȯ	�<��������|�nM4���{x�0��W�����M����?�g�>�)� |�r�=�{���mޝ*��_�p@��|������D��L�$Zۼ���B& � �v�K��<o����{1����P�����W���F�(m�`���X�PU���n��b�hdy��c�C/f�F�U�l�������72��1�<�.饈@|�ev�:p�f��1��iP��8w��-uQe�rK=�tc�
l2�S�W���h`u���8扞s�֢����jb���8jM��(�J��51�G��+��a���h9����S�:�Z�5��Ý��c��_���_s��֣C; m��t���g�nΜ�_[ ���Ǡ5X�Xv|�H�^��À�=��3��.[g'�\�����'�=�"�����~M뎳�7s��N��6�f?x��j��}u�qh#<'��"	�w*c�j��.�oTO��;}��9��3d[z�ܺ��,�}����C<��Ӥ��B����AI�
$d��LhBY���n�����jI`c�m�,�|�I��`v������Q ���ǜ-�,����r>4�н3�&tۡ����fw���%��8*[:�!�G�$w~�VT��wH��fȸ������J�i��_�Z�7+��Z�x��]�Ѯi.�hX����|����N���J��n8'�d9m���d��i�f���L+�?�Q�Nws���P*z�p�Ձ#"C��1����Q�{�����:�	�$~�bﳫ�,��.�|�}���o8r�ϧ�I��Ї��휀�b���/��|���uBſ�����漣$Jg�\M56�E�0X\��s0F�:`申Î 1�����*r�}n� �L����L�NZ$���b��P���;c�����v.n�p��&g����P>�d���ZQ��m��@��o$+�w����^J F��j<&��{<����x���kQ j��]���ڟ�����4F���1�e}��ݧ�n�ݷ�<��_��{H<S�f����G��LSH��A�P\�=�X&F��`�dx6pK����P���!�yG'�y�ko.o(NA}�HU߫�Gq�.U�8O|XV A@��.���ɍ���K`)f��C�� }Q(�XL�c�ׁ��'&��󖅺��@��n#@l>�K�q�V���E۫��!v���5����z�&N���d�
�ΞhZH���<�]�dr������}U?��fj�c�L=�L��
���� ??Od=�(��E�@�8 ts���9�Y� �A��܄�W��͉��D�ou=���yf�e���2���9�x�CG@����Pr�z��,���f
�@Z]��h��?�l��݄����/_s?Asב��A�&��F]h~�Hm���l���,����`�I
��ӧO��:��(��\��;[� 5��{c����a��)�d�z-�Y9��G�廣XZ�@��[N��L*�&��:���Ľx)c���6<���5/ � �w�rsY?���t0�.����N:jv�@���o(�7BE3�n��s�0��|b�ܹG��3����G6��iZ��.���9�w����]p��N�|Z-�`PSL�E�����x�Z���`�W,����=w��1������;�6��B�1����/�/�K�I8�vtջ�g�g��͞׈�Ҹ��9�h�,UO  ��IDAT6�Oc��Smд�� v�����hf @��P�\�ĚL8�2���)�	��G����;kr���`K_H%�>c���؈�����:N��=oǰ�s�ͱ-��1ǀ�-����U��z�=��/˝n����bp�a7�������/"�ћ�T\s��u��y�>+�{5@��:vL�P��ۄ5�Y�
v��l���P����֚�b<����55�������A�`����K��HId�y��5��L��8��ld��X�;(b���#P�h�6S�Q�F�3�a~�>ёOL�j�SBm��]8p���l5��x�[Va�l��C6�{V=���4i`���Ѯ�do?�������O�Ԛ�r�K��=G���c�<=����q
�tBZJ.�b�H v�n��X�{n��v��W��G��QB�2X0���q�B�tk2̳n͢���mOt���	s"����r^@�!"�d�*�C�ng�^	�14.�]�dZ
�J�38*gE�w�iw��t ��'Y!�.��Ob"���X=p�B����t ����y��$�>�`A$+ɀ*�� )AB��I#:w@�����@��(��A�r�bT�w��6�C�fƓ�Sg�{ ���v.�(�_G�:11��פeԺē��\��S5����X�Mxq7���`�a�G`PKǫy��g��՚�3��>1L�4�-���ﴟ\XN�ow�r�0{����`9�խh�Q
����=(�JVU�p�
��5^�`�+"�
�#퍂�f�����|./�sq5����OË������ի�}c�E�/�i�L������ML��=h� �@G%���X_�1]�0*n-j����T[o���2�Z���h�wMwt�ڔxt�%����x0���5�^@g6�*pM�2kT(��2�Q��6�12u�� O� 3W�pxk{O`���:����&�������X
)��+e�������C�Ƿ�s����3h�s���*�˶��x0�Sx?{Ym�Y����& <��b$/~��s�G'טv����*���ҹ-����:�'r��P����0�ӥB����:��x��q�3��ф"��3V������� �5��oI{��{u�Q�L1MЪ~�5�;hؠ_X�n�8�������+��~(6� ����c��<��_��2��Ȯ:��E�W���z8;\Wg֎����cVۻ��d�Hb7-X�����CȔZ�a��ŷ������`����-I�wْ��N���[\��\�\�1�����c�X\w��'�|DZn@�����پW)����b�k��q@9Y�yֹ��3T]�q4�L�vz2/��GGv}�i��|�c�9�a��|�5�}_�������� >b��������\��$vo�.���\o$*�)��h�-:��P\}��j�a��b~�c�b�Ew������S�қ�IB�d�ͽ��=��b"�}�X��9��P`�iO�|2�!s%�=Y�0�5,�$0��KCo^�N��=Q{��7	9׈���< 4ƺ��<�0Ec#��lԵ��t���#��;곏�����張�fٌ�?o]�y�}�0��'����NU6v�_�,~�I�ltVv�Jcs����Ar��|��`V05K��軝�̥�+ƨl�ACr�}�<X����Ƃ�T��g�KB�fO��D���p.�Y
���o����=7!�[� ��ӟ1��oׯ��H�\|-6F��sxX�BCk�׿�U��~��o�?t�����1��틺.�7Є#����A#;�$�bU���
zh{6X��a�	l�;����:"i�������x��'�Mk�v�RU7v�����]��4{�x,�����2|6�U�r#�В���o�6P�:S
M�d�<����h��'�U��3{�^�`���.�,��'3Z��..�)��
�qu��F8�Yzw�����v��ʙ��d,&l'�
�ǜ�}!\+��>(P�!�(��-e���a/^�/���q��� �tȵ�W�h�Sa.Paе[�ɪ�#��\�eK�"C����sV{�[m�KtxGd�qҘ?��{����AZ�+�3��e��j�_JP�&�r��&h���N��'��q�8x��LCn���e�m�&戭sO��aS�a�+�!�o=V�dT!V4B�|�c�h��� 4J]E�+�+	An0z".���F�x�_j�Ǯ���(��ę&,��&C��\�����;��0���a�����Goo/l�Ǯ��ݖ�q�"���@�ؙ�=nNE�7�7�����\�:5~�+�e��$9��.mAf�äk�#�z���v��Q�&��Ӱ^���/�=�r��L1��*���H8���sv3��gdH����?�R�5?�4�M����f�k�� M�F��ցol��q����4�$ʖ�B���w�C��'��y���������tʿ�|��ϖ�za�
G�h�Ajtk����`�`#B6C�I�ER�}�.GY@�W�F}O���޽R�6s��9�t���>��{o�)�(ǆ�>�s(/� ��O������#�s^_߆��0G.�2XQ����I��k�tx���1��*�.�4U&S{�T�n�S��>^���dos�*�QT��@�Bk(Q(ဗ��()�֮s�C��퉓��2���hZ /�110y�H��CY�^^��{3'�Hb��	6F^�zM�`c�P.���6ٺ�zO�m-t]���]+���@f�?��o����I�871��gڇ�"~N6^������#VWW�}(�i���i�4 Ard�x�������j�d[#?U�� S;Ĥ	���-�#ݷ��f}C�fw+
e�q(�k�}*Nne6q�ݯ���J�ϛ��z-f\�������M�i$bd� �3�U�	����+В����Ϟ�T���3�[��M0�1���Z)\,�6�ε���8#�h����yo"~�noy����+�� b��[�-��[��tX�¬����~���CZ���8��2��7��`NSX�,��e�0���m�@�}��\�����ʄ��ό&n�&�m*P3�[ ��({8'؞��#�ƈ��\x�c�C���,�-��Z�b0� �z��@��aM��r�/(~;`�%�h��9�:������%���l6@ߛ7�s(6��L\��Q9g��M3������}o#CEs�q�K�ڻ;c��֭}��g�F4�Cf���ӹ�0-�_�@f�F{��K�s0t b~>�e�}��1��Y��\ƀ(ٵKX��|�_�|��b��)y�1S���Z?ZAΆ70�4 B��ee�9�飽��A�K����b�վp;r�.U��i�|ѻ��9�%cqM6 ���K^74��/W��7�MZ0GE�8]�[1
\�w��/|4-b��a;�0�� A�~�Wӈ��lhb�VvmΕ�#������ݠ �/
S: 2�b��O�ٮ��.�ۚdb=�`E����w߱�J �$"�xƽ{:��g0��������_�,���?#��yKF�;�g���c�E��� �|�y(M�>4��o���څ��=5R�Aݨ��;5+� p����qϣ`��Z���'ӔK�ۿ�� �Z1"I��sӑ�w8���W,|!L&k��L� �;cu����N&-bٻ��{�*{�Ӽoox1���P �3�7}Ԩj����;�º,A��.b��s�F��i�>�M֤���? o�+ݫ���n�u��h&a"��~��fw洊n��1uĄ<�� �?�[492�u�M����~8�p�)����s�O�3��70s؊uv�Qx���m�õɚe�D�\ֆ�:��̝1�ޕ�He�{����K���"N�}�����a�b(�"�k -�uؘ�џ�,���De�)W����F�q�t�g��i�9��fcFc	Y��bGJ�O��^�Pʽk��jm�
7���⢚�w/�����0��7���7LN�(=���C��"�t15�+<� �v$7\�ws���0��*6�k����� 
:;�P잛-����x������@ʂ��օ4a��֥�`�E/(|��f�yP��~���xGdtAF׸g�\JI}1,,�ס�۬�\�$0-�J�8�e�g�Ŏ1q.uGJ1��@oqmK�u0��:Q��&N@��(��7��F]3n�ܛ}�>r,
v���c�ؖb5�+�։:]Wցch���~�����k v�'�����!X������{ԑ����6~%����vM�Fbj1}_t�#��)Y!9Y+J�n�[$"wKF�Io� �9$4������ #*`�`o^�}m̅��Ӓӻ����߄�/�	���Y����C�Ս8p���
���/E��܆���� @-�-	\r�H���v/
%���^��H ��"*����8���;I�%��/��[:c����6�OS����K
R"�)�������PC�ܵ�z�f���6
p��@@$�hZW�q��,U�6�Xcn���fm��0]Ѱ�|�l�"���D���|`�ܢ0����g�U��'��`ZQ$b��4�vI`z��׼��`�qͻӚ
��TXJ��s�d�����}_��OG�b=��ڬ�%�_t��׿����o�)�k��eP���%�sb�w%�O��8�
�G�3Z�ɢ�b>�(�Dӎ|����V�l�FV}������A��~�s�N@WW������A<����×�sFM~�,| Ӟ�F]C�٥��'_�����e�F�Z�^kX�Yt40��$�`M�>��.&y8�d��q���X�"���{��x׵�Id�XMq����I�\ژ�����p:>Uv�K�<3�"q���F�1)tW�|��{���Kx��c�������s��K�YZC�ӓ�{�������_���|�5:�o�0!?�}�����Ds�gd>5J��)l�3��U=q�ƃ5B�`s�_�v��'�X#��DV��3���Y��rv�����cglp������`�
����W��ꆧ��[��W���,��.O�;��Iy�Tb�톦Hi׻�����1K\��u�8E����\f�������%���Ӵ��x�{�X��A�V�����6�l��삹1�����D>��Ωd�e��;imtK��׊�\��S>������:s�{�X6>������+Z����ʉ4���i��z���g!�=��S*S���� .��F-�9.�n�,��g_|~�/�O��|����zxI�2��k9�?W�������lZL����(z�Fz�S���@�T��d�Zl��b:߼�c��v���Ӈ�<to ��PU͈ϛy>�Aq3ǻK��}�d�&��%L20�1h\�������BzF�s����k9Z�F�@WB�p:"�望���H�F��6��P� ⧘dr<t?���dgc�9F�cƟ ��僺ӯCg?|�	����q��O
`	��7;�Ɛo �������S��K�t ��he.�8�����Hۃ5�;rd�G#e��[�-u� <�c'��g��={��c� @���p� ���{u�<�R���A��{H��v�8M��z]њ�rk�d�r�zP�eõY��R�$Y.���7���:s�4�2Z�s3�|�G�p
fcYC>������ouː+�@C����8�E�᝴���P�V^dwc	��u�+Y�ApV7�.A7����y��ds��̼�8��IX9[c�Á�6�;�1�n����,��7��ϳ>�;�DԞ��B�������"�:��Z����9�ݻL�B�H�DhW��[,�W� !���켃�4ݡ*Z���8h!�g�GW�d�jB��sd��V3�7�$X��ї��X����❥\�-IM�Ц���ӓ���&�\�#�%U
� ���Mb5`0��>[��qTh��:}e��#C-������j9Z�N<q�c?.�5*�2 N����o���~��|���v��g���t!�|��KpP�����k1�(�:���IE���S�0vK2-��E�O�A��nN�ބ���7�Tpq9�P)�j��c�"O�Z�zo]+n�kJ�cQ��N����_�k�&�F���}]�`T\����p��&�ʧ9�֡���u�N��Y��,.���d"�����>�E�zX���v��.��?:�d{ͣ��ս)�{l5����TS$%؄N��'_��f�ϓ�:��
�) ���@�|T7�x߃s��P�AkY�2b�H�P����b,��Hbp�����*�w��K�����; �w�'`Qf��\��c�H�;�\cu�)kՀ2����7*(���(����D �*$��� [F�K�|��,�Ͽ���m���s���5;o`����/ÿ�뿆������Ś���z������� �Ci� h�M��Y�&���!���1�*x��$S R���A�.��pܫa�V�1ANٚ?��H�E��Keŝ�)am��B,��r����#��}��^rJ%nr���	������ �e���븆5���+!��8'��r�4QY�⒃W���/��S���O�h���	��>�Nd�n�:��x� C{����Eы������;��a���xQ∁4~6�M/䒏-�����֕�#����o��ቂk,�	�"�Ћ��%h <������<&����K���U4��ѧ��ݖk:?`F�%�qW,���
]e����&�9]�9Im�)�t�K�i��&�32+��@"��T��j%d��u�\J���V��p\n�/g�-�����O����"�r���|T#��d��8s��͚�O���I4�������Z�{�L�M9a���&��ymd???F��uݗ�C�S!�b�>%k֍�����a�<=�H}��
�jX�=�I��ί~�s��G��| f���D�;k$r�qr�F��{c,�����e�5��쑅����L<ϙCP���Lhq��u�B.�����%�ˋո�#��g�̚��nX��6b�������僽�f=�K`K�qo�g�E�@,�c�>fϭ����8V���2}
�����{�� ����ƏlV�?8��|�zxŘ���	��J-*��-;���@@�;d��n
��4��F8��εZ������{�^ȍ�����R��8b+���;3^�jmr��e6��f��G�G�V��5?�I�g�DN�fN����1Egk_r�d*y���W-� 4�O� 7ペ@1I�����~_�ޜ.��і��r�����;������`�Ip�<~x&ґ�s<lS��,Qo.��_���'ߨ�!�^�󌬯%Z�O'�
⁺l�r���$:�>���_	��(By~���D�u�bt���y�����++� �,�I��z�3��;u�12A�,����}=��q�뷟�?!u��(�Z�:�H0vuq���$(���Y	1��/���	T-��iJt�`���+��~��gd�(����Ư6fo*���X�Y|ԫ�Y�RJv��\M��\\*J���2SQǳ�>1p�7tl@���ӎI_�W����I�g�Gɀ
���4��A��s��@O}���q@ǿ<����������@�9XqY��Č��!ڌ�P�hX��"�/NB��4Z�O��t��{�u��ې�I��Ͼ�=�?�{�[��������f ���p2M�`݋y��n���
ȳ���}����'*��,�9\U�4�p`lG���r1e^�\�&�֩��P'�3��8[�wMX7Z�爛t�VK��(��C7֗d.�-`(�|K�{�׳wڮB�V
��su��飏�E��J.����+8� X2��g��������=q�2�H��ܵ��Z��(8��@v]��:v��@��5����K�`���'�皬H�l}�PD�$ńB.d���5X�kZ�G� a�q�&�+�\k��ل�c��e��s�u[�#�(�o�����E��7�ԡ����ة$5~�& �{�]���o·�~���?����_���=���|8�������-;�8O ���s�'���lY�&�xgI�f.�_����L��FH:%��Xк�o��J��đ"c�ţ�Ə�M#&x3V�(�8?���jX2[�m<L ^W�
�cϘ�4�������J��8L�/�P��LO����F>��9/ H��q!PT�g��r@!�mZz�Y_H`)�:�#�[��p8����᷿�_��c����?���o�?��?���?q�ץ�\�Q|���L��ԛ�o���Q4}�_����0�%���ND}s�#����O���:��72_�&�9*V(4�$d
�^�1f`���Ix:�r`�@t{@��ب�FW	 �[
�J3k�}�y��6x�+�O�M���~8P�U���).�3J]ܙ�VD��Ri���byTC���1��p�6!�\%Q�=b�bM ��'�R��dTAr.�6[4Rw���P�l~ރr�`�����A�w{6c��e�9��M6J�2�y4Yq�AL�(���ϱ����.t+����Rk�&�������Y��YtC���F��������暍d�$�jY�K�&�2��o~���~~�˟ٵΌ����=���;칻�Ş�;дo�IN��<0�����e{��d6�.~��~D^��F��c�<�@۩����X4$��N����ᐌX7����`����މ�p�3�G�;i��[����;�U�{�F�}�� �m�os�ڐ���|�7��Z+��qb���(���Ĥȹ��0E�>;:�&c��cu�*y\R�!6�^����Ad˶<��Vr�}�&F���$t~y~i�OȌE�,Ú��n�/��
oY���d2n���[��ZuM�z�z��G���y�#��Q�U�75M��D��~�=��^��mp|�����c��*Yβ tz�G����	GH���P��=�)�{�ٿ�10��t���&f<�h�=�	���X+
��;-HJ:w멳��c�Kp;�es� �.%@��5'H�x��.*!���n3��%�Q�?��.4�&��4�=�=]N�\����r���Pɽ�QJ�u_,�V�E�r�uxS\.'��,�0K� w!
�i��F�m-��͉��#���2�,tY[C{��ސ���}zo��:����^.�9
�sN��z��;�L:!.���Yq$�l���ב��!��6쬫�+��t.�C���ߙ��*XS�hT�c�����a/�����,�[:8'��&��A�P"��@��{�:��[����h�b=QjE�ނ��
��O�DR2�<}�;k�`���fE�=T�A7=?�E�և���և�U��v�~ �(U������/��s�>ʚ�u�ʚ)���$��{��s��o\#�<v]���Xb���.8R�!�mtαG��&鈡x�acE�'��ntsL�ѯݑPt��FQ�*(�^C�K�FD'g�r5�u�Ņ��8���v������ahGN������4��N����}SN��)��wFgv��a�î�z���P�/��Bn�M>ݷ��2�0ʻ�@���y��HAm��>X�3Mː!�9���ׯ�"�C��f�uM׶�w�~C�s3��ӗ�_��__~����o��X_�@�G�����"�Q�	D�`�3}��N��X� �p����o��R|<�{1�BF��]��G��X0`��=}ܹ+��%��
,���K*�	�&c�������5 �3�blJ���vI��+i�q�K�\�`�2�PF����/�� �3�H�؂��CmKڱ��p����|_S�����7/~.<����~x�;�[�����|���xͻw%9K��ňm[`?w+���z>6�V�Qu��"?��P/α���x}�`��S�1���/���x���c�5�!��G�̥o4'!�{����؄K�q]�g±�tn����R��& ��.=_�=�&G�.cK�6O )NDͳ�I�k�E��s�P�l����H���� ���l�P�U9(sa-��
�ix�=�Ϝ��q~�$ ����ܖZm��$v��̓�c�\]��&����ށ�^#�~��]a�9���Ǝ������J
��S��sU0�d̓O>�t>�ؙ���b�]ư_���t2�(cV;k4zCQ�	�:˭!���,�-�A�����<�������]=�ۇ״���{5g���:�+kdj�a��kn��@���	!A1�s]�Iqbʪ��$ 6N�1���%/��e��X�&{8W�s�r�O걮n��-6�2&�?�5lq��3�~��$�����+���݂���
����S�xۘ����	�E�LY����4L�<!K΋��9c)X�xP��`�j୹��0 cYV�gc���+q�8��G 	�p��%9�����wA�7]ӄ`���(�Ha�%M�97cO� ��s���'4d���F9��U�<���>����u�y����P�����9�ڏ�d�e�"�g�P@��I� &�1�7?���A�ȅ	
K�Ja�Y���P|�l���@����\�f����:-P����9�qe�u?eS��3�ƃ��$��j� ��K��֑�[���P/A"�&D�.�\�.�n���Y�}�	ǩ\����N	Ue��piL:lm��5W�MO��SX��k��n�V]�3����̃]IJ��Sb�C:����&~���B�jO.�����:�_�����,������k�#�^Iˬ�C�����e�x�����>*K������R
�C	���mڙ���4�@@Dg�V&�D�h�d��"Ȩ������a=�'��9��}�k�����ի0�A@m�S���[e{��<N LD�G� ��a�ͺ�^�vl��a�FC_�J��ȗKc�d�~��A�8�C"��!@w�� ��� ��T����1����˸f"}g�w�{�h����G/���� ����v
�xѨ�@�ӱ3�Z[лj�Eu+�)K}˾0Qw<|�{� #ԝ۠�"֥��$�U�A�n�,�(�§����>Q�f�p�EP8:+��|��JQĄ�s���<��(��N1.�ռ/��,:]6[��|N�@wN��M������;
�|Y�dՋ��$g�B7�7`���?�S���7G�P�߾{��N/x;��|�葀E��dl���B��ݐ�\�]�p��xn1�j�}��9�Uq���U�Ħ=�r����u��	�,��22�ē����?�w
'g�Kέ��sɳ�X ����-;� 5A��tQY�Ǐ�����:P�5�! 6tm��=b�A�b["��}����6�i�5�Ֆb������Z<߆g_<?���i��m�(`| r0S b����߽��
��`@�]��r�2Jm�5��:���׫����s+um|/�3R�K^��>4�%�h]�a�0�
�_l�a��RZUX��Bn�1{�|m0 ���L0��q,��W%����Fyw1}�RkBU�x�EP�{ѷ����g�4��X=�qg{";�!Y���au<����9[�y�g��ay�b�-tb4}��k>�P��W:��t��HQ�=����k��[)0��`������=OG��X����G�c vpvPkU\gq�&c���Uw��1=�1Db[9�� ��Av����K@l�4��Ź�������?�i��Ϟ��C�҃�XcmM�����a'���w�t<B�|�zWng� �7���\��1��T2��7�H`�X��g�D�7�=)�~�i���8.f�ݮ_�����Zl6;6l��?�'g��y!������(�d�!w��0:�j�<F�`IV�G�p��X�,D�]���s��$�@�`�=��~>9��A���F߃���tˣ�+u!j;�dd��q�^u��P�=o>yͧ�uK���ьE��I�X����| p ���Q��}T��Q֫+����i�ɳ/³���%xY0����~/��w&�AVQa��C���nޣ�Ֆ��Hr����S���7y/�
���И��#Ɲ��q��2~Λ�+�p�o��f����g�|���ݖ;����u������o�|�����о/�u��������"���bs�s�3�b�q�@%�z��:����t�Z�bt�A�(k�uۅg`���6�7wz��$�U?$BUæZ�2{Z�E�t�i��}�/M_ �R���#:�H��;RD���Ƃ���Ҋ������E�`@��V�������zߣұ���:1�r�H���I�LQM<�+�DIܵubэ�ߙ�Ksa��k�Jz�q��:�������D�-S7)-����S^���0���7��M�qʮ��a�b�~�7����V������%)�9}�v|�GY����|(U�d�=��֞�R�b.
�t��,=g1��1:��C��Ѥ}#�|��>}���ඒ]o�6��(��ξs}��.�$��޻����qߗ{�����[8��k�DŚ��X�E�"'�݉�
���d^{�/�x���A3�r�Y�-���J�T~7gs5N$�

j9�O�$����uЋyg��k��H#ޛ8���5������{��\qp��
n�B���^����H	~� ��`_`\ �_s�2Ӭ��d�Vv�Z<KR#���^,$X����H
�&$�{�פ�Qi�#AQA-�`�ȱ�Ľ�j����\�~�+s�LA�q��}�uy?>��2���R����2-����(-�`��~��� ^gcL!.��d������'|��di��b�:h(��x��?�9���9��5��WU����
����~JKg���_����� �M^S[�`���k�K̒�=O?�#�ӧ����Ɵ��9�����Z�s�l�
�����!(i�9�@�^/b�����Oe<��"����_�<� ��|8:�<�i+O{�J�<��ze���4��F�	��������Ma��x{N6:�ߍ�.B��{��`��R:�' Z�|kZ9���oë��|1'�?��k���Q(4���/��ڃ�7F��jb`�����hEk��^�7m�1��[ ��	�pK\Ro_�Z�����+�"M�[v<ńt�An%��-�Wp��R�Ŵ�Iu�/\��ȵ+ <#/�> �����Ί
���m�mC�s%�S�S��Js^x��or�ΰ(@���T;��zU-�W�F�����`M�cd��W�9chg.,�|8z�OV�G_:3:������Z8��^�0�Gkb:�Nl�Xbg��蔃t��5�F$k�����,�"��΀\�@`g_��Հ���=8 �������r��Qc�<U�F�L��|*�zC�G���n.��¯�K���D�)
m:!�-�Jb#���7���|a��������g�����C�Cg;.쌚R �M��!���8Ce��{Pr�qj������>��bz����R�+�rz$�"����5��hLc_���Z2�F�����Ql�{�g�#�/��}g�avNb2c�c�AZ`$s��`� 5��5��>��H<o�� �d`m`�L�K��$	e2���~^8ێ0JKRu�b苖����2y`e2A#�h� �3לף.�т��b�
���.� �~����"ښo6�y~l�d�=�ы���`��|�=-�0A�uE��<D�c�i���.�Y��=h���+lG�3�8O)���.�C߽�����@�Y@��s�|�6��vφ���p�7�E\�$�;1$NU����,b
 ��0d����h���w\]<�IS�ЋF�nw2�q�����'X���p�d]�Ū�0�����/lN���%�8�x�J ���/��%tWo�ܑ���f��k���N���tE�q��O:��BL����6�)��՜p��9�@�N�(��Q�"l��YOB#�Bx1��Ȳ6Or����n��{GAL�:��!@�:�����ʼ30�h��ıHq�(���)���8����u-����5���B'�-�ۯ&��u��v��h�^�?�N����-�H�Ӂ`h��)�s:�U��!�I��w7Z���g�uJ*��l�a`ڽ��b\�s��B�Yj��(�*���T���w@mX���H�{N��V�Rǂ�~7��^�E��C{O�
��u�aΔ{l �._W�_���	f�ђ<�Iʟ��\��p�EDYA�ٵۊ2N���:�{�`s�!%���cIZ$((>��)�� w�HA\�5�B���W�{X�xI:q����=�8k� �>�G����ax�n�I���_�U;H��Ί��싹Y�-LX�P>�~L����fnZ�MC|�W����d�N0G..��n>	u��X���/A�=yI�c��Q�;P�A��Λ~��?ب������缶o��{�
���qh��4��6L��y�$v:�lq=��-��?��\���ů����٩����~�o���_CS��ß��g���7$���9y���P��u�X�J��}�
��ϟG��3?&K0�5��k��=Ę��Dl�F���[�Y�g��-��mu�N�ZIb�q��?U\��;1b]Q��\ ���E���YwM!ptp3�z~�>�/������#�S-�տI��6S26��N2��'#gX�F�[-���L��0#E��w�4����B�q�Fl0�~��o�W_}E��?��+j3A<�'>i3�b>�3�3M�ۙ����5a�X��5��:��f� �B9C��s)ݏ���]n4ϴ�:	���[(�#]�s�u�6t9(gs�]�x���|��B^����k�k�/0�}?h�v,򤩣�ʭ��9C�α��T<��5�n?���l�����e�E�a� ���\��h�9�qb��r�Jܳ;s]B�cb�ޅ�n>��6�9�P�6]e� �Li�Nl{��V/�.;s�H��?j!������y���Ff:]��U���>5�,,Q� �[氍L�ӂ�jg��%bOf�kSC#��i<�D�Ў�ϫ���LX��X����F/��/ȧ�{�e��Qd���)kg�s�����l�$#�F�O�����1�� tv,����{$����	�O�Hn�c�����]4=�3�M2���.�<�� @�����n����F�dhYPj$��������w�"[Mc7>�+�o�[+
�#s����߻�k�R��4�"��r��=�����6�Pl,�Uq`��ծ�i�!�Gv��I@8�<�uC�+���<�����d��@��f
�i���+�x3����}d���i�H������?Tg�N�:Gm�q�z&{�R�MZ%d�n�u�N~��p,�P;�߻�|p�/9�y����;Se����4��a�Š�N)�w����!p�}x��t�pӔ����e�Ǐ��=�Ia�C�(�"=�� ��/�V;[���43�9��N肜͇��!��Z2���Y��#�	��N	L��Co���	*�`��&l�I~ƭ�J��$6j�(�.M�r]�����a-Հ_�0���F?���Ű m�m�Ã_o��������ǣ؁�М@QL�IG�5DN*�#��n�$�e��m���Ɋ���c_fy��a�v�=�s�<1��B����� H�Gӱɡl���u�*��8��*�瀓�·������D�+��T;�~�ܹ�6��b]�Ч)#3�#��pbc���h���U��J�y����l�J3�}M�sq_������$�-�& �kئ�N{I�2�����@s�L@�\B.l?��s6� 3G��Q��j�t��Bu-X�ZЫ`����l + )�d��]9�Q�}�y�8O�>&��ɧO�  �_�a�3��՛7,�^�z)k�9Q'���(n�K�umS�~4�_�@sr��{�g�g��#�5�H$�tW��|����.��<��y��k��T_t ��3:Fu,����B��boU����H�B�����D�w8,��i`}u������x�X���I�\ϒ��w}}��|{rk�:�V
<c�:�������&������M0�@e��oGV�����"z��!�� �]��`sh���~18�ݐ���έY��������4w�`�C�N �dg���B�Ȋ_͒���~�)ެH�^��ƺ��P����@���OCrǱد�3l��y�r8�	�@�Fb�45a�N�3ptVL�m7w�ژGK9���9���^�\�T�^ ��H�����
��9�hd�Ϳ9{����� 18�0?)�h����.��z~��Y��8[���P;�c{S���>ƣi~&s�+���g��f^��Zϟy���J�Nhn�_��؀xK#

�*.���SG�C�
�rtaΉޚe��ww����:xk�;o���^eM�ɞ.��q�c�:΁��}�7��>}��X�/��uiz4��ԛ`� ��|���@�2����o(���Ŵ�}��ޅ's.���'�=Y�n�>l��&�ɶi`y& ���9h������\�z.��U����*h�b}����^�������,����F���^��a�qKw��dG^\�q��u)��/�H4;l8m��*&4,�*��;��T��u�ԏv̄l>�'x�
�м�ڄ;��?��*����ĺ�r~8�бT��Ը�[���l����KDy���h]�PxNj�	�1D���MT��'�>�H�>p�s�X��Em�\���QB��Ϭg�����>G3�� ��jm䠭��{:�r��`ų����8��zkXD�J&�py%� �]}��'��{xEM-gG�ъ�rӒ5�-4t79r�'˨�	���g�'|�R��m�CY72��8a�B�!GknSuw.�:���K��b�1��Υ�u�3>�,��B����g���\�����|�I�s��x�������?x_�Z��\ߜ����y�Ó�eM��IͰ�N�n�~'�6Ż�3ggK�;��[���6/���
�Q�F�tp�ٻݑ��� �V�s[�@��nۅ�/�Xr�Rዅ����B�bJ�&c�L��`V�eY0Fu��ͻtC�� s�8ӽh�nXu��;=�G[��a{���f�!����|P����(�ɴJ�b�	|]��;ɺ���T��O�^���S�N�����Ó��$?%�yQ��Q��~���6xc�7Ϟ[:v�<-����o�@��?s>
^t��Ě˔8/�3�g��U��;���U�x1��r��\	+�#ppR�z;S����`<2p���˗,�.!s�^��cTW0�8��]T-G���i�c��;��]�W��yh���_�����
e/��cE�&_�Rh�����3:!�=q� 2v>	��禋1�7�/�k�
L��on���G��4J��\l�z�����^���x�q4U��"�Zp�'@�m���:<݌*�[��qY[��߄�������w�>��\����$��R�ضl��P^�����v`��E�u'cN�ƶ�.�}k+6@�{��!�S�5��\�cMJ�
���	�=�>������b���.��?�s����ozMƜù���,vSR���{�9�c��(`���z~�"�&��_(f��4��+����-g��d]K0� �Хd�����{WD�sq��z9�=�ᇯ�X�^g	0TaU��1ԑ�'*O���{\��Bi�0��z�"@��e�������>t��� �6��:{��3��@�qiNTkk^u�-v�%<c�:��L$�l4����#_�}�� ���fһ9^�����D!o0���5��+�Nv�ŝ5�=�:�X����8�m�dq�@�r�jl���"���"� o��?�k�QM��(F�{���x��Exm�97p��L�q��B~�Әk� S#��\O�+���@XA�h QWد}��<�s[s1�qW�֦p��N�=]$�3����b�E���i�[���Ns8���n���2<��W�غֈ٨4i�ѝ 4P�县�����g,k����˿��m���;�xȡ���;G�_�� �k�0'�h�.g�)To5	���,#�ao9��}8�A�ՙj��GY _^��O@� <o��ywa��<�l����	��T�+���*qv�7@���9e��#�~]�g\�x}e��p�g�r�H�r���"���$��Mk�tf�p:��, Zi�p��Ǻ��~�I����v��&c[�0`�'<g��n5�P/�r9f��~ϥ0�����,A�O�/ڵ�p�����P�
>��#�4��8���#��Ȟ@J�H}�v[��q}��}�t�����g?	O�\L=مO�B�2#�^��zw�ߺ�&��c(5|0NMGRw��������v����烎����ֹ��|˛���&5��=����s�'FG��cfmC6���أ�?~>=�^>��p��Q^<��k��e]O�u��R���r�wG�U$����&(�?���fos.���W}A��5i�K���cמ��v2��h��PLK�/�E��9+�m����uF�㗻c�����ް�JjeW���F'�Fl�Ü��q�����Y������C�C(쳞�E��"�#i���ՁK�\<жs#Q6�w�J�F)��9Ճޓu)��^)�,�L<iפ��o���bYm9���WP��v���[D)�s�������G#�{�X}x�-]�����{>,�= �0s(���h������uO�O]d�,�yn�ӃyȽ�>[�cո�k��C�"Xv�6#��V��Ѫ�a?ں{G�{*�#�
�47����>�Y�ߞu,I������q�{O�5�-`� ���$
��0�����	�?�d1A1i2ud#��ڑ��.�y�*�|�Zv�����ةx��J�#/�mo��A��u��@��?J�?��~iG\w)4����b�����]�~�Y�U�9+�I�-c�[�k�멋��������0��yH&^���� ����v�,���*�퀶�&����}��?��Q���]$Mc؛���F2���=���F2�R�� ��o���kk��W�^��u �k��6��`�,.sV��w��2�����2�	� :kH�P���ݳ붓�2��4_Z����K8��i�y��B���Ҿ$�uk��׆�{����:E��>�t*z��)M� ;����5����k�4W�@h �L�0��Q+�=�`����u�c�	��d�l�e}���.T\�r4��u�����]�~;N����� �2��3{
c�R��o`�v}(��Q"����ޡb��@Ü�c&He�f(2  �1VG�q^`XHq�`>I�v�J����7���f�`0Q[� \ۊ����{l����Ut��\��u9����86��5J^��W|}?��`�����JΩ�j�&����޼߹o�}iś���ؗF���u���i���\Ků���ݱ�h�Zo��r��>_'�0R�2%]��-�5C�M�'?�����R󽢃��]jk{&����̱�P4����4p�v<(V�(�5�?cL�&���>~rű��G	����\/Z���
��[��lȶ,�I����1���W���^ �e�^~�y��-k�_�ǀ;��;���3>b�������G7�{����=T"  ���\8���` -^o����ƪ^U����ϒ�������h���e����`�h���C;�{�0I�{tTn�{?��O�� P��z1[,��bb$���^�'��ފ���)1�(L���{�XܙϚ-�{��M��:� ܻ7?z]�9�9�:�E��<�f�VL�䮊�;8�&N)80���Ļ�~�X
��f���������O7Vhb���G���~�c���d���jc���qa.u���	m��	��oH@ ҙ�2-Aa<;���>�[�q4�\�V+!}��E��c����@�ms`����C�e��m�68
ڛ6:��g�e�gP"�DWk��n
{�� =uw	l2�� ������q/��è.+.E���p�\ob���.ʱ�\�j��9<&�lB��Sck� �0��V�bR��� C���S��ϩ�v�T\!�u]n����;���{h���?�j�������;^����-���ď�����>v�}l���Ծe,@���
�"vg�&�&�z$��Q����L�X����Z|���tNJVg�r��n�ȽŦR_�񢴭Э�>��ռ���o("
%#����D������Z����y1B�O����~��i��`�F��hs`��+�%A��K�#? Fm��O)27��&D�_�xA]�D��J�� ] ]�,�c�}"яͿ�R7�j8^�����:�(�'+���j�a՜�Sq#Һ
��X�a������%� 쉁e͘���W�����Xta��	<;�������^z>�9�{	��Q�y�)q ���<Z\�ѝ�!���K5��7��N��L��ّ�P��wQWt���ݷ�o�7�A�?�w�/k�+��8�������ܩ0�mv��]h9�Xۏǅ{�;7�崃4����81֕����셓ѹ���g�_�n�[ud�+��k�8����r�T��."z|��������wEG�g�sr��=��0�t�(�4�<��d��&�����ps��(�{�X�Z��� J��[ܡ�����Nk��P�ȸ��J�*�}t� ���w꺺��}��:���q��{�u���5�Ԑ���1�:hP;�lűL�.��b��B���	��aڙ��!�ɽ�<_�9���;������=Ły���caIn���>�g��/���\�c�xL�@`W*��GyB0-�_M6� ��e�μu�[ۧ`��3羸�8��&؎��F��x���s�V4�M�87:�����厣p�V;4g��xk��Iw�S�ᵐ�ţ��a�G����K2�,�6�tP�4�u�cS���&�>���lL�^���t����t�N ԟ>���ln�\[SI�K�Ü���i��L����w������y�N9��|D�߁�x�l�^�~x���>����r���x�&����Ǹ6�����jK�zcqB�b�.t�2�2�<C!I`i^�bRN�� ����	����!�o,kT��3 ��9�y�Iδz���轀6ޜ���ͩʯdc���k�n/�s�j4J��?:�ά��\C?`�����,|J������;ۛ����52�h
�� 4�d.v�?�G��	���}.���%�	&����P���g*�G���Gl����$Ph���/�Jv����bx�J�?���#�����\�:����A#�TcZ��2�$fSo�Dk�ޗ��vuչF���6 mf����x�*wY:_˅!��끪�DT��l����_μ��Ŕ�?�f`�X��~#��b�Y���������Lɒj��Ζp+K���`6�j:�U��RX�.
�Z���d��DZ,�(t�\kn���l )���d�i2�i/�`��	�y'�#D4���C3�>fpJ�lG�N�l�`�����2���P�������s��[?[_����?���&1=�/ �nZ�N}�5�����$�Y�H 1?O��T�!Bꄮ,��R\�����pP']tP�IN9H�D�d'_õ�� ���ʣu�^��ǯUo9�ޝt�\��5�b��G3�5D�a�H�蹐 �|	v�\<c����;�<�?�޾}޼~�d�;�{�E���c�f��A���~Fק�����,�)V?��5౳����?�uP�JB�	6��X�
���.������"�E�H.�-�������̯s@��Cg�&\���9vXS��~qy��sw�;ex�ظ��{�}�>���ޏ��=��P瓕:���7�t��uz���;9ǁ�u~~ɦ�Ȏ�F��}u���r�\� ?�����5wI]��R����N��7�s]��%b !�0�KV��1�b󌱮�sͅb=�wƉ���}��N��w����3>J�➤�g����>b6A$�� ����l_7�{� �OG5~�[%��bc���ı�ܙ[�ǻ�� �$j��8�����Lne5�;?�f�����	�X�*r(�K�}9绾��\�ǣĺ����nN���Y��y}	�rW+��hdz��l #��쀩s��+�5ξ��)WRS���bq�M.�;�����<��VZ:���]i��Tr-�{�X��7��-��A��qu�wc�V���h���gC(�Y
M_��qi���E�������\�4+;h�;E�c�������$�x-�x��*kl;(���u9�(`$�;F�v�J%�O�� ��4���?)ꛆ���-�� ���)������~v�s��Kʟ]�Z ���ظr|ɸ9���?~>��,t��/4} �=q_k���k�e� %0*�~��uxg�9_G�#�;�,~t�y�@K1Y���p�	�{s����Cyt���
9+�3qRSe/󃲋��zk�(���Iu��ڔ�>r̞g�m�7ZT�h��s^������d�K����g���y~��@��dc�U��jЧr�i�ig���>w6�5�%�S�H�X6vL6i��Œĸ�!���52X�/�l�i��O����--.
N36����֖�! ���m�S'��ߡ_oJ�x` �8��S0��?pa�?<K&�U-�u��kN�t���w:;�����P�|?W��OZ�� �s�)=nt���_����Y��PͿ�GS���5=�:�|{��6�M�$���Y�����͵�&A���^��جyc�i��h�D=�T���W��Md@8���m�b{â�N�6Lк{G�$=��s9?_�$2��g^���t)Y���wq��;]W	� hk����is�<��i�$��_���)��R.ͬ��
O�_Y� ���
'�� t�\��y��F"c`	؈������&���ʁ4Z������釂/�S��~p��<[��%[�#���u�=8v�C����}����ߋ�y��9�j���q��{x�Dm�?qA(�ܨ�����΀�Q�[����
��w8K���Ţ�G����{�Pe>%YMO��ju�;�x�M'Ɋ���]�`Z�;��{צ��?�0�����T��_o 0���9�ʡ�	����9^.�P(T���8�S������,Л���k��T��n� ��o�8�� ����VC� ;>�u�=)H^�dw\�?�sz
L.�>b�Cu)����bң�$�~8x.H�R,���ƗȲd>��{�.�����{���Y|�瑓R_-��.H���G>�'vAu�QDf�A��FnS�\w�]�q�	d.\�Jx6̸絣�EJ�fYl}�>�XQ������-j�BG��G�w�йa���k��ߒ�J��LǨ�P �ȏ�e��5%�Eb�h�$��z݅�Zk<��_C����~���k]�'+�;����/��x8zKb-Z�>0�45�'5��ŁKc�t�b�N�g��PXd�#e0ԁqt�b4@M&R߇cF���y���uO�F4���'��|�:��[���޳Q'�h���&�7�������m��̆���5t@'�a��d�w�z�X*{C�A+���\@ό��\�ܺ�ԟ�|n��҉�h����=���N��47���+���(+kl�h�|?̝@�3-ܪ��w��* �g�7[|������5�v@��I\n�Ǫ����DM2��{x���" ���6;�z�%	��$�Wh�,	���C��?�K3Ł4*�Fs��kh9Pah�C��ɴ��.�͑�"{�P����LBB���]m���VV/�ɚ�]2a���������b]��fϑHX�?y�0<y��L'��b?��?�^o�r,� ��d�� O�8������K<��%&@��D��(��$I���5���+~��>J��}�X�@L��c-�"��Fg�%5�t�Ú{��Đd�ދ]��^ҁS�����g����4�Gi���؁�ǁ�cS���H�3 �w�E ;Kol8*5����+>��g�ΦZ�dʍ�/�NC��1@��aG1b�U.42Ȟ�ba�q���9�o.&;2��4�O����������Ȳ���#�?�!������u]2����~��4����ɴ���F&�T�<>|�l�\H��3b��J5�),2ƌ�~
��3�9���BP��4��jz�Qέ��N�`��:���h�X���@<C�L��"
�Lp��	��u�h`��I\���yz��z2�T�ZXFӭ����m���dK��삂Y {�9��e������`Wt2�\�A��-��-�iaH��)f���$�!�C�A�%��)�u�������4�|��n�����w�ը|�s)�XvS�PLw��5�^���fo\[�Y��l*�â��4��=��@��l�L +�gV��JY�jnx'��9�������!�p
ܔ��M�<Jo������O.�w�|a{Fi;W�1L��ȱfΏ[ڀr`�O_;e���\�����`��ء�ߑ��~k�R���jG���%�Xc��s�������w�>B�y���%e����=mwpvQ!"��u|�L�]�˝[s�����;���u��BA�K;'4�N������ZֿG9�����������.y�c����cƗK�%�`�2��
TkԤ��������#pj�R�{�K�t�0�3a��aBY��$�.�{��]}-���V��I;l"#��)Ea������,`#Ug�����m<����h��ݹcw|v�����3�s��Zz��o�`D���C��o��"����IgLŗ���{���w�AI�����~�>�4	t�J����D�������'�^##�8� &b�D�*�s� p�R��\�}�ME�ߣ@7m�wņ� @��5Qf��!�[�fBW1�r۫���Fx��m� �w�����%N�"��m�t �c�D��3f�3�r��K�n�5;Tv���+�TA��A�pSĵ��.L�n�#H�FL1y�kMgl~1�z&��Av�o��]���ƾ����r's7��A��:���{ҵ��i���&10&��c�(�i|��1~��֩v����{��ُ�JDrE/�� 	�����ܦ��=��Vr�P��F�TR�m��e�@'�� �\B��5&ss�/�Ve8��1;�Ӕ����� �ǖ� ����s��ưd�k�B ]u_�{��Z��
4��v>�[�ɀ{�26$&�^Os����u#�]��O�R7�@�7�x�}�i��9��Y��z��1,�4��)�{��9�L\ƒ�_����΋���l��`�����\�4���fG�R��q�(��7Se�x��=����J�5�5w=[��׳9�~��',�YC�q���ݧvԎw��⬓��2�e�&������{*�z�by=����Qk3��s0�%Jz��k}�м�}y	vx�������tR���������r�&.�s�@K��՜׈o�\�Ŏ��W�#����������L�ؒ��B�K^���V�����%��-٫[�$o�v�����w�ȑ4Z�����������������ػ�G�� 	�.2#"� R��/l��I �������c�::(a���}��+ž�u��7�Nj���ߞ�p���>��qu�������*��gf���h���gW� ���8$�!4;�AZ�D,UU�;ĕCh���O?��~x��� X1Ar��Ies��%�>�f+��l/��{��œ�����<6�B�J3Bs�bj)^c��(��܉�u$���|��AܛO'Q�����d��{͑�F�r�8t5��Ǖ`G�#�ⓛ.���=}��I�m�ވϲ$�w���i��� � OG�b��3N	d��BC���p���S?/�0�F�nDJ��"s|�O6ӁYEO�oMl\e����O��Ğ=�F�ۈ��0B���NN�<T`�J#��`(͡��g�go��e(�ڲ:�#a�����O����� �rG��@����#��_��h��ׯ�W��@��A��e،�Lf|���)�!�|E繧�5N8ʦ���3���b�D�m���cp`��r��$P��
���'�?cfH���l����W���Z��[�����,Kư�߱�K�/�@�؛�����f�u���������V����� �k�����6�խ\0���2wP6e�jy�g���v���q}׹����/`h���� ��>Of�:f��1-�m�ݹ�{|� �tR 26�p����t����Ļ�	8��t�`��u�@�0�r�s<��qh�.v	����"\�/ñDFT��@M����#h������K~� �ur���f���m����t���8��R���ٙă�>Ƴ%o$�"�f��t�ܑ��'D������#��#A�.u�h�\XW�|��_�PsDLP�2:�-,)���k�!|;�ѣ���
ֵǲDV6�h7�p��*]!ezf��S<9����)ud�Χa"xU��{/&
���:�v�%8j��̼��9�e�N�h�{ b��(9����?�_'s��һ�~X������K��d{�;��`�� �皃i���������;st^1GU��s S�]3|-�Lx������p�s�L�|�s�ws��y;73�zeW{�g^Ƕ���t�k��k���2�2M�~������/����Zޕ���@��d�I)@Z�-�Da������L����Y���b�+����CPg��9��vW�	�-��D�82�S"�nWh����+ ��1D_�sȹ�����؃H��%��1�[��Y:�\%έ�l^>��B�3�T�m��-P.<m-�ԙ��%�l��<آR5���C���q&��d*����ص]^r�!��;I���� A횆꾋[* �]��b���+�숅rH�7C�����׏���ϩ|@�w���������J�L_(�ke����e�'�Ki�;ߜ�:�Y��(iA¬601;a��1l�5V�]A���W�9���$�T�.Q�4OLJ�|?Wt���f��sݜ� iQ��"8��`���3����ɜ��^9#ǻ�.���9�����a{�����kA�B��錺l���������o�?���.?hU��t�`R���8�#]�wX�p�ٖJ���~�j9���&�|��8[���1glL��k^�˺>� (��X!ї[�"b���5:4�=�J�zƒ޾\~���g��L����b�vL����do�Y?<tJ��2�%����1���G$�l�x��8�9x��N�R�|���G���{CNhx`eE��ʩ���[M��u�Lz=3gů�Y�&��@��P��0���q�'Ӹ"0�\'%��`1�im�����7o��hI3�`f\P&�%̗���Ƕ���}�wpmw�K%i��9���cl4Rl�5��I����P�$@bK��#��95�ZG|�I5����I=c�xg%�ڏ����fS�w`}����e�+T����z�u3yzOjBE���C�.w���G	
��KQ�k���wȔ�V���z��7�#�L�<Y��6��TJw����¯�ʚ�q���.ȼ�e�r�N�ر���!4 ���2�IN�E��E��ϴCe�Bv��HwΙB��C��r.��A�
+�ZZi��d�|�۳���ʨ�����*φ�vQJձ�l�"����憦����_~q�d��T�IsN�IS	��l�<0k�j���S7���u����nn����-�e�0S�lMdB�8�k�2s��T�l~�N�V{�[pj�>�M���}�T�X���!o��[Ӗ�Y8P8΅�Y�]AV� �G��5�޳�Ӄ?{�B�n��*��O�	� ��v�oN���х��Av#>�θp� �|�`zsf�R���mK���w�堶�HY��t=^-@����|'+�����bs݂	+U�`�7�[�u^z��J��A��D��c����G�9�w�39>�H)W�bdp'-����[JV�!�M����0���+2���ѹе�n~�UVK[�4I�`^%*���Y��.������Wj����s���=�GR��`��a��Q��vZ�͔�b^-�=��n��%��te����a��%@��~Ƅ�zV����@���:6�g�7훭�yL]�ϗ9�;v��v^��M�@6ٜOc\��O�u~x�ځ/I����y�l���hRʏ.���bZ��4�1QfE :#�`Ş�.�l���>mO���u{�_�ܹ������l"�+	�41c�N����B{������y�r����bEh��k
�^�����ʓ�$����$��Ŏ)����{{N{��!����qgэctOS�
ּ��l�J�oｮ)j��{�����R�!��B_�#��:��QƜWm~�\׎\������S:B?�����#���z	���9E�$�v&X�li@q�pi�p�xv��:�v``9���co޾Y��[gY{@�yb�[d�����]k���7�sYL*w�������:�`����[�?�k���]�����>�YZ3�gף���ݿ��<pݭ֑l_����O=�/G2\���'���Q��,R�(�|V������D��,����G�<'�>�:�II �]���|¡7�Dff�q�ˮ_�~�%UV�jI����>'G�!xt2�.�+���&��o2Q�_~��}�H^���� @6攃ؙr3*,Hv�toy�V���h�������c��vlY��E�t���9�y�>֬4��0�{�YY�sP����ſ���7!�e�U���U���>Q��*���{4\�5``ȋ��d5���#�g&��Pf�:F9�=۟߼~뀜�t��Ԡ�Ʋ�b�(
��@>�����bc�*Y\���i�y蠍^���~/���[�2m��i��bw���6�X��X� KX\�m̗{1�'c��ӧϞ�t��tfI��(>������[* Z��sG��6��S�����Cف�HeJ�4��A�9:f��N�]�f��(�}A��p
ڥ��{z~�G���ѿ�J��tr}	(���A@�!���`�}uR�>d8�u1�?�{�H뼃v�g(#Ł�fȮQ�7E{����e}��эY�d/���-a�OF�{(�����{T��Bg7/b���2(��ސP&19���;����	��� C睭fv#8�p�V�	��
� ��g:e�!���uO}�곬���߾�!��LP�]>�_~�Ło��l"il�edf�(���ɐ���b���]!�hس�Ők��Å�SSs�|	g�����4i��N�io?�[�k7"�C߯�3-�^�c�رC�L�s�����ư�͑4@��7��6)���mٙ������^h�2��6��n}��rK�YXǬ/h�l���3֙�J�^�pJ�ir�Np,��3��9�F\�ÝGd�}��sX��b�T	�r-��k�Ʊ-D��Uu<��C��cCFG����r�B����Kc���o���v@lp�hqPT|��7Z����x<F��4�18�(o�&�{7��̒�v��ٗ6��!�14�րh�a��S�vmm�;W#�	ͬKu��`�� ���z9=�O�rsR-����Y
xJבn}N�����������\����i�*�M��D7��B�\��O��5h�}_[��>�q)i5��X)� ��6�`�W�jԝ<��X�S�<?��lL��������駟~@���4'���3tE`Q�L�/���i�k�G:��DHk�d���-���ɀ}���;jH�V�lKn��F��뵴�a�PX���	e4S��@U�a��x�V��F���_�&{�V�&{��脬Ya��<�X2�y�����ӆ���nu�Kd�R�㱏�$]9}����8Yǯ�s���@�/T� ���u f����pK�i�sk#�%Q�S�%�:��v�~r��íK+g4s~A�lL��3��յ�ϐ��,��	���������}o������7�W|e�t5)@ǘch%ypJ�^��|�!ރM�
&�϶l��=��$��[��o�v`�-� �=��3������W���d����Ҳº^l+(;x�옰����W��$�k�u���B{-6��ȓ�f��Qwh�	�� `g�Oh��2���
�z
�"�G�uO�X%E�&���c~�u|�:o����G�J�V��*�{�:R����oA�u����ӯ�w�&�IZ��| �wtM�e@�L�3E���|�����!M$,��D�<_��_������Y����:�٘��3Ӥ.�cH] 7�����]�鑀^��E��2��Y��&��v�zu����m�[w��	�� u�uvc`�>�c�H�!�����?$k�sw�H�3�f��M��	|�5^>����;��l�b�e���8�J�������[�jw��E7ё��w6O'&{�ǁI {�����C�1�'��4� w`��N�g�-]V�
g��:�9�1��S�d��	��{���U�����N���ǭk�v��͹��K�vY��`���o�.��$�D��K�y�w��[�%�F�P(���C��v�*Q7�T�W[�՞Y����B�j�1�y� �p�;u��/��'��hYh��! �]��&�=[H��,�m�$v^���3-��53����.v�G�ޯ�x�t1�lȇ�K!R�p���w��f��?���FBP��96dG��m�W@ZI�r'�R;�w�f��c�Q?���1΅X�S���h �32�������+A�D�M�L)d\2�l���@ں�k H̛�����eƤT��O�s�"�-K�~f۶�i�e]��LE��U r��Z�тNW���W�A^^{c<4���Q����:*l��7�r�L� ��7}t�j$S��'�(�_�#G�4b�x�![˪��i�a|�u�9���z��1h�C�@b\6ǥ�f���S�KҠ��v,��S�vp�˘f����1-�s[�<L��)Z}�
s�"c�;\�fM�e���KN4���32NE�e_L�K�]_׆���*����N$� e�(�?���g��.o]��y�-N :]�{��d4|W�rgݿ��3�CЗ�,H���_�޽w^@� �д����S����Bbx$�5��O]��Fz�n$>�k���>�`9�JM]}<�-W�U��g�oLN��~s��#i����]-����U�����s��u�`������kx��!����S��j������愒��{3�݉=��{���4�S��
�T�C$ԛI�Iԡ�!&Ke����i�I�Z�|5���G�~�Lq����a^>��9�҆�`0/ ��Se�(#82��;��J��Y����`X�Ap}@���Й	�ղ��&{�ܞ�Am����_Wp��l�5#��5�b�nO��S4�PZ��3�.S-!��U��a7!��W�X������ν���}eh���4�1���8\���g��-t��r�q0�9vb�Ka>�g� R��?s��yF칶���jr�A%� 6Ҍ���1�k.�,	�_d�}�rqVz�{��ne#�f[�h�4��N�fg��l����	�;�W�	�\�JN��l��M��l+a�O��S�k����ģ��	B�7��M{�X�uq�����ϟY&�屉@���z̉ Q�@�%)b�iϼ�s��:���O���I��gTp�Rs���V]���u��T7��Aܣr��%D�ud����& N���V�b�9xg@C�6�h�1���Z>�>k��i���{\�]�s��gd�ݏ}�<������cS�`���=�/9��+��L�x�����ؙr�ԜG������ƿn� �Ҁ�$i��� x3!���f�&F�󊑯��*2Yӊ4�]]c��p�l�Y1���I�+������u����l��R�O~4�B �ENo����j�#���C��������>�S�Q];��qϢ��pʊ.�zI7�v�����E�������#Z�� h8x{�D`��Ƥ��rk]���wl�p��������tp��O[�b.��o=��RP���� �\pE =��C��l��-"d�Q����j����):9=HB��Lc���A�xF�z�z?3�R�����VV�`F�Yef6&ǳ�*��Z�R�G��ɗ��=�N�lE׶�n\/�ܪ��}Kg��l?��l+ ��F�B��,���S_�gj\T��߮ܛoNðCu*��;7b�K�i�gj���B�<Ĩ��X�s6��y���ϟ�^�L�P�ydvAL8!�l ����dK��-���g֙��W�C<�e2���R��D�1���J�P�!=D�鎙��݆��m���
�ެ�ZΚ5ͬ� �g��o�8aL����Z�ä0|ڮ�g��^k�5Мİ!t��(���:�sޖ3/�pY>��)�g���}���R��Ȟpko4v6��Ό��ݮ�M<7��.�����e:	�����
x|������b7�1��r��І�ۀU���� f ��9P��h�F;�6��u��m��9_&ph�Cu���+u�� �;���gO�Ի+��2�F�<��1 ��`)��9�}2'tu��\n0]��S�(�����o@��<	!˙�v�u�
~E��5+]"@�d��u� z�k�/�]g�K��6ÂJ�g�MGd���	�iV2h���c7#�T ۹�z3��q�W�㾏ϯʏ�o��(r�d�7�ڝ"��yc����_�)�:%2;��-����WB`��G4�(3�i�h�r"K��1�� *�X����m)�fӅ1�o�J/��XN�Sc���̈́RHP.��}3ub���]�N�I|�0P�'h��ٝF��\ D��j����!Z?{Y��i�Ba�%�^�agy�5i6[A%�Z�:�$��4����������X��,_������GgkƁ�%�T |��㱐)�����n��4����1�]o����p ���geS ���gW��B�V��v!y�%��Hc�㇏�~�ٓ�
yx����4`:��3��k�9����߹�~]�s�Jk|�k ε��c�.��1�>��oUv۲2d�TS�G�#툴�fJWhmv4��6�~xoL���8t�b\�����	��hs�$6N�#���;2c��s��Qa������<~� tUO��Zb��Q~h��%�O�3�	��GVS<�|��}f��6o�vs!yk�� /�d���[��{�Y��޿����J��P+V!J�+��?Y���[w&�` �}y�Һ溌���%�!p��
�ܸJv_����Ț)��H�DT�6��=�i��G7�� v��R�*�S��I�
3)9�<��m0l�M$�&��ω��ҔLh�Q'��tfս���>0���W���)��^������{�X(�;�ћ�9;�&�����x�k��[Ƚ��POe�'LՑL������.Ou�u�]4uFRM��z���x�H�;DM�m��6��<���7��[��*'��qOO=�R��(��<�rHd��N�����$m���S�1(�j3-�.�s�Rg��rs�ӿZk���֞b�l�}xi��2|�m����N葉�S��n��7T��| �{5ÊR�>6`|f�d���|K"Yɝ9*Ͱ�{wg� �p��3M��E99B�,�j�Y�F�,���M��������b��D�#�P��BD��j�b�a�q�c�%�Z7 J�̤�?z&�2/����t�YN�5��	�!�Q��pA���B]-�N� b� ��Q�"�R�s@m�!�8R������k�v-Xv�$�59d��T�Wm��f��Cw��d�mv�i�	̚Mo�8�ɻ�y7ƚ4p�#3lb&����� �o���%�ټ�%,�����eu��QznS�=�~zg�J�V�V����]�&�A�����XJ�;=��)�
X ����N��8~�gI$Nm?��:p�����]e`̡Ã�~%�^�۠[
�}�l ��h0��5�v�
AΔ���̦Z� !%�Jn�� �9*X�}����h����}H@� �������r:d�wCW���j�k��с�X�14���q��11�K��Hi��f��tA�Lߎ�#�"�Oa���&9�am}�������k�z|x���=��d��*K��[q�Ԝ/��������t� +C0?S�C� �~����iFM�xv�&�:-a��: ���L1��%)x���&d�˄���^P>' E�h�'R]����ʾ�!�qG��f�>����� ������;k��l;����V�/�*5���M���l�2�{�����.�}�׻w?��}Fc+���q�a�]
p��)�oO�Bf�L��|����k��g�e�f}h��+@;`���Y��O�ا3Iy�O Ԇǁ%f�g�~ 8����"_{����oY	��/wn������v��|���/�]���¸`���~����ե���qH����^����9�{}�6��kK���
ڟ���c>�7���%��%;������lx��p��}��z�ch��;D�?FR����k�	�g^���j�>�&ȉ��!�&�~��;D̤D�۪qD��np0�ʩ��H���l��k�쇚XGZ�77d�؋�8�h��^��UŅ ��k�"yc/B���g׶2���~����<�d�6��_�1���\*|dY���r�����ʜ\���o{>I�=�j��K��S�ߨ��q9��T������p:]�=l�K�u� ���g�]�s���`��5�Wf��9u����6΍8� ���t�<ަ�/�K^Y�/6�0�ӂYS�yE��f�l�=76�9���	>�H�s�W�t����\�V�0�@���.D&����;r0�A��@��� �L�ό����u��l�D�D�E����_�8�����<����'*�@WsA�����y���i�
�%N�Õ�d�ȩ���ʾ?��V�{J1ߞ:ZPg�q��\�����R���ܴ N����|J�������=����V���Kl��~ ��8|Fa]��M��i}Y{�m�y��Q��+�4���ڎ�Y��17�W�4V\�F!�t��i�y��䮎�69@gt,p�w ہ�����z�% ^$.��-�TC����	b��f�$���3�s�}#4����,��E��Qi�W���YL,�r&Kվp1`�V<��"Ü�H����ߚk�����:��:�,�9�3J9�}��t�Ye��6�'+[3'��@ 2��M��\���q�MT�|=K B#�TG�����E������j���X^��y@���H�߄@��'��Ȭ1�����λh�|K!�a�#�����Y�b.���茂#Z���_~~t1S���
[�UЭ������T�� ��(1����8Z�t�O+������e��Z���	*d�O�>��#/�<Yl�zl�,=�E^r�[k-�����;�E ��'S�7�mXQ�#6��:t��f����������yIm�W�Y���h+�ui�j6g�^� L�!���K=�.�7{j0���Ӊ�}pF�`cd�>�)���:�Z~��p�R�=x:�i��`J�� �%2��|�U���&�!�c ��Zve�D�9Um�'�[Gf��M	���)�L�]1�*KH	Ai�M�v�j�%�j��fC�e^-~cw�u��j;����	d��fI���!�	�J��G^����}H��k_�N�۷o��꥝�����=C�Ou��v��Lf��<��>���Kن��˽���a����%���"�1.}�>��Ϟ��A�a��	��w�L�b������:%���6��p����1��Oׂ����so�󮺉���;�^+d��Rj}��}��[�������}e�K�9\����8'�:Z��Q����kpKFMϦ����͚��-�{�k��yX���M@"�G�;smُ�G�jo�o�&�-�(ٴ9he^ѭ� y�]#`o���Y7�l�e:F0�d�&�N ��T� �����E� �J���{�Jn������]N��Rz�.�1�������ʺ_ k�v�n�(��>z��mU;Vl+��g���_u7�f'��)�#٠�[Y�:����$s8+�ɹ�돪 DJh��ݓ#���Ua��6.l��o������7�ٿ	�hc�6|)�#�:	r�|�2����F�	t��5Ԙ�E1jhg��=�$ɩ���j9FFLIt !6h'�`� ن"���<C�|�׻{��EY�9�,��6�W{�ɷQR[�N�V0@-N�9�p�V�� &D މ�G�.ݩx�{��̢2�ڰ�P<Z�仪ϡ���r�ܛ~��F�D���FmP�>��u�j'�:8��g�5)��s�YŘ�VyQ����G�b��Km��:-��G�,�^fP�5k˷�����-K������ymƣ5d��_�p�R@�_|b5��+���fW%�?(��@��bY�xBK�zv[pa�3�&}8�:����v��/!���^Srf�2I96xh� ����n��̖���q�l��(�ٳS�ֳ��ȝ�5�l�	��=$u01�m�z��ď���I'�<	��.D��R
��L�N0FX/�]ʑM4`g&�Ǿ��nv�@ku� $��\��֡o[��m(���p��5���zͧ2��8�F+G�?'���lIF{Ld?+ �q�N6�͵��twK0�1#�;ҽ��~�>�|��>�Ł5��+{j7k+h�|ON;6��2���lf`s�p�*]_QfQQ�O��9mt��Y��@�a��6���A+Q���_'��X�#��g�;�7�訌�f�J\k���b�+k%�� ���;���-��>JB�T ����ۙ��&�,� �r�K��M]��������9��>����<}��sX,Vdxk (�����ް�:���|��s�9Bll�9[���z0�'ѾJ���X[*I_mO��w]�j�(|o��:(u��h��^W*�R�:�/V�{��I�]Wx4�����D:�)�g+젽a-~-xq@Ӄ{D�ׯ_�i�|-�w� �tJ��˲�����q�l��EP�@�6 m�'ʔ�+�d�h-U=�	Ϻ��@ߝʚZ���c>A%}u�P�EQ�UYe��뚹	f����I��G�/Q���/�G�=���ɼ��ZFX�lm�?�_�5����8��z���3X���M�X�[u�Pv)HB-{�"��煂�*��8F=��8� T����7�S0���Y������y���cgW�����##�+E����Tpy���~�vĜ�!���텉\���>���Yh�~�����
�gF�5��d�?�c��B�]Xw�m�c���Pee�����P�Y�pt���D��x>.��i�Q#=H�s��f��b���w�9��cؕ=�J=A�I#��Ig$4d��fϚ��E�}� �=�eF�	DF�}����!��)�
�*!æ;ct|d���0���p:���{���m��;#�΁�̔����l�ɮ�@`�;�"7p�D��,���=:zvhX" �0�|w��+�)�m0۹�J�Ǿi�D��j�-c?v�d�;*Aɠ>E]m�V��$CY�M�3�����&^v�~� �w�}��v�,��Ŧ������K��#o��1����uDLO',+���`�M���B�2�w}�4�.Y�w���=��j�&�GQY�Y8JjBV�>q�7�'��{_f����̞�צ�U��T'��Q� &�P5�gj�(S��Ú����U���.O��!B�DPp�j���G���C��n��|����ֵV�i�{�q�0��;G	`��I]ED��'��%��J3����+6�sU�O���t�R��{���8Z��Q��=��IH �V'G�ӂ%[P������LFv���sR� ���8�k�m��������1,��;f8p�e���X6F����Pr�&֥r��p�Z�程��$������ޮ�~@#��%7��D��9έ,�6���!�+�N��c�\u�����S��S+z}��H�S���&̔�Ch/�v#�OQ��(1��Ҫ���v�m$��Z,�ڝWA�&�'v�yjÀC��"H�� �?T0�篲|9�O�d�sH�f��B²*�r9�Y'+�p�|d��4����Y*�/��8H=�=��&�gr�z����y(��6x�Ԇ�S��z�:��v���k�ao��X�nŝ�KA�?����T��w��zk3j�-�aY�#�� ��`?�1���ʾ �@d�u��о����Yd����q�i?�����k<R�7���Y��a�ֶ9 �k�L�DeX)���:h��7V{uH��a՗H|���IH�#�|aكl�XW>��ZmNg�t��tҫ�!�iD��仍�BD>T�J���s RE��o*�͕�h��\�vi��a"H�*�P�~���=q��6E��������T�����]��Oy�����ʀ�~uքJ��s��m���]��n�y��e�Jp���.��ކ�K ���@�����!إ�����RUЉv�W@V���j��/�²:&�ܼ�V��A�=g1[8�8�,n<�B�j�Aer%O�^,R '
2� �Q��ʞ���	�b|n�ZZj�(KS9�a�g��F�v@<�Am������z	,e�=�{1��(��ND�� ���9M}���^�eq��1��}�%�Ԋ�(�#�6�4�\�K�[��',>�x�����#�������`k����F*C~�u����sg�l0��u�ҿ�f�� �`<汀mb�G���N˸{��q���q�u��0)�HaL��xv�*��)���.��L(��^X����B�ky�浯c�`f�.c����=�(0� �me�%�ITQb�������� �)m� �z�
�v	�C��� �|�"p����u���=�c�=��y!�m3�F�G*���e�Q�pN0jW{�&��Sc��J9�Lឱr})� U�[�A�H�Ӑ�&�ģM�Tn��Ago+1f������`6Ok�ꉭ�9�V��|�1r���!={���la�KL���ڂ��,��=�x(_GS7u�����{���jbs���k�@|J���K�#�!M�&����-ߖ�����g,8z��?�GS�)d��;>�
��h��1��}X�g]��?�R-U���Y;�{�6yY0&,7
p�$uV��ﭕ��O����\T�[�sL�FkAz�6���(;�
�L��=I( ٹ5H����p�U�Z����m*��c�?�`���~�ݘZ�[��E��Z�sl�-�ǣ`r���l�4X�R��P������B�@������ȫ��n"�@e~��4u.�&���!�:X�8(�4�_z�얏M�w��,���jn�:ffO��a���C=�ap�H��!�NKN����rge�DfZ�@�f0��<���'�|w� ΐ��J	���ɿ�~r���6�+�Z���}k���#���S`�3��v5x�g
[��1���i�'RƇ&+mN�n�9�)2H���~B/w�Rf�	���A��|p�g�@�T���jt�V�fm+�aSP�+�&�)�s�9ґ-�G�So�ZN���N�}tb��6�͘�\�k�K`x	@F)2ʉ)��m�,�'�Lvp�Qʠ��/�N���-+�3�.+�Sy�J�Ū*c��*��3-�Sd��xa ��5�Is����r��a�A�3�[0��� Ƶ�*kU��)�Kd���sPaF�эcd^S�
�g�.es��L��1Y栗�];˫Ús�s�))��x���mu�
(�X���*�(�Sr��ك!Y.y	�1��g+lcY`����� 0L�Gv�Gv�Z��#|�EHm�*^A�`u]Ow?�����S��A��i��y�I�� g�9rϚx5(I)ʬ��6��.���,@�B����ub]�|�j��k�]�s15Rh;�����=O�)�]'sB�i���LM��h'o`���S��J���7�~���KZ,1c��u"rN�u*�m����ǡ�5VM#�<��
߻�}v�n�H�V�99��j�7n�sыHG�����zB	���k��-�)Y��1:���;�N�9l�����Դ���$"/�b㷮:��*՞Ȑ�Z>*��8�S���i�X$+T�f���,�;r�ڗ�6�w�n��r�=|�n�<{�1Y���������7�%�)^?Dr�M&��ϐy���M7���n�zj��Im�����x<R����g׎b�7{�V�����(��s���^���̷�6Ⱥ��1�>`��gCҍ����~������Ɉ�6�Ɂ(�O��fQ�'c�:�M�'�!xn���IH��[�b�H�_��܂�p��a���g�W�8\�Qgu�MuN���e즔���h�14�j���.����X�S���$��xY{rM\]� vt+	"�tX,C�l�:{�#Sk��zr9\G�=��򬶗tG��mOf2*����4�u�tV�*7���<����⥗cɑUf��
��R���AL�i.U5?��-sz�� *��;}�1�:HE'���������+�VJ�mt�8S<�����V�w���l[P��<�3E�Tk�*���Ɣ�%t�G��(��0�k��=��CxO*=��پ���ˌ��8�
ڂG-���ۮAn���]�GEN�z|V��<'��#G`GF[YO9vب�Q���4zn�ٝ�¬���fX��/�c��_�c��т������k�0���}��Y������[��8�u�M��l�&�B����tKT���;Wa�y�b��2�z���##��=��3J�©O>	�:*cA½�h`�TƋ�
�\����Q{�h�.6��?�� ��~�Y�)7��uQ��_��Z`,��������V.�wǍ�C��βg<>� ?X�`��C$�l�9ӎ��^�=2�� ^���⳾������	G��!'ğ����u����|$1F�3̤���0D2%N�C������C�st�*��A�C��*��Ο3b�zfe+���:��%��Ȥ����e�%�|��|���z�]�=HV�x������e�s�2����>�@�iG�X���%��:�u@����� P��dS��k{N�����kff���ڔ~8����.�w�__�ˁ�%N������<��G-��g6�w
}w���v�*�-�/{�y}C+u@'%�Kt:�fќ��vN{^7dm/�n���?w�r��3�s�A�˼��D;Ɖ�9Z�h.ҼNə����#�m��l�ѩyA3��_8��q�z�6����sP6Xc{h�X�D0�"PX%�a픚tk}�<�z�%��s���]��K���j����M�_O��� �]��r�����;gC�>S���6eNHV���|� *�>���E�b��g�Fu���2�h���7o�O?����}he_��@̓�#��Wq�icfe�Y�L��}w�ՙ�M!�#W����Z���?Z�U_�͙�<u����`��j��'V:�������W���{���?zY�t~t`�s��2 X�:c`�;g��,��P�u{{�"%��)#�ҩ;�.�kz��%�߼~���@�&��Ur��C�ߩ�4��	��Ѭ󧕈~�v�;_�b�@���2C����a�س���Ä�s�� �U��OS�UU�"ն�n
�T��Y���_���dM|T�6uɔ�K��y��t�2��H�B�S��?�\����k�!tꊘ����q�]9rJՆ���^�d��\s}1�� v�8�um'�ą�!|�r��*���󰽃�V�W��2�� v�9�H�G��"�\��ˢb�����Oc8y��0��� qU-_�����K �A!�w��େ�|���?yg.[3��j��[��ǟd(�:gt,_U��fxt�����&�S�zIkvm�T(f�6��v]>,����_~�-��˯N)6A:���N;8tw��s_�\��f��@�2`G5�)U�J<����{_���x����N�|���c�)p��r����k��}O�Px�5G��z�~WT�Ķ��{h��\�����`���� cW7�n�R릝�{��閟�	pb��P�ϸP:�g9f��	ƺT�� BR^;��mZ�֬8���� b��U�a�LN �I�6:��m���zfum��	\
�[�3 'f�3'� 5���8�ܔb�촒�?�E�,�A���d���ϥ��KG�N�<t�2� @�{L�!D��v͵�>gts�n�����J�T�����2�P�Ctɢ�˖`�X@ P�j��*:�a���_�~ʉ������U��Z���[3܍�[2��o��?����V���u��3��]��4���ܭ���Q��K��Ym��+c�2�p_̹��JP�Z�睆���;g��P���I�Oe��l�lr���A���*�vt�<�	O���\[7���#n�1@1�#ǿ)�,U+*J;�J��YXb�%9 ړJ�Y���%�l���c�{�{F;P�u N��j6�Q�\I-���������>�<S�dN�['�|�Џ*���^�� �b�F��3E0S�Q:!m����5s00�[���[$M��"��,���<X�t��!6eT~�s-��k�~��a�K�&&D'�U�\F-�(�&�l��?�����?-��WO:+`��C��ʅ�}�}^�5�-v1�*�#�:sd��g�,�~��
*���$��ŗ�����Q(��_�n�me�{C��Hn��֨:�E�����O)��aε�B���9�4~�a�)^�z�B����_���e�X�7��� �p�ϱ�XVJkA��P����U� �ѥ���a���r�FC�_q��y�:4�sUV����!�$�?y������W�\��Sz��_i��à3j��N��r�o�7`������P�<u�� ����g��r)c�a��7o�:�h�uh�q]JF ɧJhY���"n�޼M_�~�Jc�؜��#X�S�eڬ��f�*Q��%&l� +j�}� �\:HX�էe>~����K+�rAr�5���p��E[4�y>��yc��h���f�tU6ưl��؟3�Dh�U����s*�;]�k�o�G�_���H̵s=Eq�?�[-��6��&�����_�����g!�RcL�R��i����E�:}e0]���Ǩ��V�:��x廤]5,Y��ƹ8��"�t0)���|=�I�_���e�({�����EЈ�z�*����eِ���k/eTW�K@�P�9Q ���s��8+` �o ��:F���?��G����_Y��!=��3�wh �:��i��V�6�n�X[T���6�$��Ale:R�ͱO�HY��1�ϨNN��=�`I\s�u����[c�~��:�y~����1�(|�~7m��&(� ���R�r��֟*�@ɐ�s{�!g
�!���*�w]��2և����/���w#r}�F��V��T�L���J�'�:���NVX��\��84�{8���m�r,cv4�=�v���pm��"�G[v�LA���*	1�9���k�Qk=ՠn7D�"&m��fӅ���G�N-��M�]]#nw���cn�:і��FO�ᓖ�mx�aC+bԅ\T��m}���,p{����9��(�5)����)�����Q��#�]��
D����_0Ϣ�/�I�%����'��I�]q��il�Qv���ERCG�E��$���5����y��3N�������:&��`�P��`���Ǆ�/����s��wm����g���A��Ȉ�pas����������(��-�ui��=�2�`��
K�3>��xgkq�hMNf��Ao�I�H���v`�̫k_�������ҞHM�`��9ҥ0���ZĆ��ɹ��ɽ:�uB�W
�a�~���Tv�%Sv}�E'�iRk���g�,%��Ӕ�%��N*%:�80g�Փ�(p�-�z���Ľ��[6'2���>�Wn�
&( ��sW��ѝ'��˩�`J��[�u��Z����b�����.���+�_�dџV��q�6B�c#Aӫ4���6��.�x}h�%;^���Fĺgw�I��b���GtR,����U�|�p���o&�n�- iH�k�#]�'�7"���9�����oL�����r�o�~��{��Mz��?���'Ɣ��������_���s��O����G/e)�G
Ar���L�x?�I �Aa>P(��`���깤j�'�7�	�6�yT�/�����
}QO�QR�5�&$��t�]әs��(�E��2�7G����,���	쩁L[+��w+;b�30�?:c��>~�`g�;օϯ�潑r&��bQJ�Ld��j�{ŀ{UW��ۇts�l��Q#���B(�V����?�CG�`��J�fƚ6.6/?c���|�����)d�G��	LkذĞg�]i<�R�u�1����s���c>���6�+c�ͅ{\�o��٥?��H���K�GLO7��$qj�.��W�7�����7WD�_���J����"O ;�BF5~�v3Y��8�*�ެCw�tI�ok_�0��~W��TAE7�����tP\.ē�w/��l�od���ea�l�`n6dwرF�Ʃr&,���'ˣc��N�t�ٟ����F�����ӑ��e�����E�r/�k�M�ڳ��L~��jk���#����������ٝiC���2EJ!Ȓ� ����zW���Z���@�Y��n�����Xh7���#G��?1VZPG��S�,�V/�{�;��>ss�A���+ՠ(5�M��ބuL&{�b��	��N;���J�vA7�N��#�R9�����Y���Ύ�l�d���[IGP�f�S��OW�e\�Z��ĭv��|^�-����^\Ƶ=�8���r�&SgO�L�΃6�i�S�9m4�=Bqd|�&�: uT~c�"ۏM�]PJeF���`;s�|�w�)���ڱ�[P�]*��a)�j3|�3'Lu��o����%�@�!�Թ�e��s�I��l�zl��=����,@'n�? ��ײ,+��A���|���:Y��B�k� �uP�9��3J�s�f�f�W�����)E]�$�-��o��Mj@(} �e�wh	�%9���޻ �'%��	s���л}�@$��κ�#$;V�i�o*�{�D�+�����c�-�i��.��\�p]�w�3��vm@;�o�q��Y#3��z{`�K�o�QOK��˽&ԑs��C����]����];�v���p�ňFL���kg�f��5�i�:�v?j��	��6�Sxn��.�z�YFSe�g��8�5�ϰ+�2��̀l[;{f�_�~�~���?�!���?_c�Hrf�����ћ��k��S��!��{�reۣN�"  T[.w��18�\Ipm�i����8�3���ׄf u*���-��g��%e��Ё�K)r�d9O��߶/�u��s�{�bؓ���yR	/���8=�����=��B;�6jy�3��y���m��ĕS�W��Y�����u\���* c+Z`lbˮu�L�]����L�￧��������[�����h���c���غ%�̏:z�$̙^���f2�+%����V1&=I��u������Z�絉�����&_z�����|��ǵ�X�`k�l1�L��Ć	�|��+N)f���s���a�������vC����0�����LH���;cfٹ�����8��o�������-�}�C�x���ym@�A8
|^^��&4&��u����O�>�_~�9���_��z�.p9�wg���^��,;�v���pI�>�O�w����W���d+��z�ę�	�be������u��K
��y����w�r�e�ԇ���c�m�9]���q���c5g=�)�=�MIT�d
�Z�0��=�C���
�zʅ�g4�;6��
d�ï�����+�@ߖ\o�ی:m�)�2�9n^��0��D`��1�@��/���&�o"g�UNsR�	7X}&�{��9L�:8%nܝ�B�5�̅�|A6ldlCE��h�\�����װ��oz��YV?K�9�$4�\E��]Àc� +�V�;:أ���P�@j�g�l��{w�>&�����z͛C�I�(ނU���_�RN�p��!��o����R}o�U�����!�іn�5��䬔T�������6�B���@�۽ȃ0�Si���R��"��e*�������p��$�7Gdm�����0R�b̖!(���B�p({�&�G��T��;����d�g�7l�(��}+�^7� V�6-JÖ��"�@� �G�aCk�\���87�"�z��04�3Ka�	2df�qo�FNo���t��hl��G��>;�ͪքA��,� 	�\�z]�0�g��9Sj���۞3��ؚb?��"����F��AP4"���D箂�8g
1p�:-h�8xr,��I{�����6�S��ʰ�YW`hn�/�]�6�f��`(K�d��fծb�y
�2�Z�̆��� �?O3ʏ[ +g�L�ڵ,�;=Įm?2F������1�>�C�g�$�Xֻ���K�_���	�P��hM�)Pj��ɝ[� ����2ߥ�!�/�$]�զHB��(i�6:H5�d )���C�O=��v�
D�i?z�}u��^]A�`O��^ǉa=\�|��T���=ð���K�C_℗�^=�L����	byvT�� ��Z��9���S{j��s�3�^���yz�β�(�F���{h�Y�-�����QOq���<�UF55�1�# �ŧ܍��w+PY��3YY Bˤ�QE��ߛ�]W�Kw������7�r���"��Y4�,q��JpKM��央#9bQ���b��T�W�k�1IwJ��ֽ�!&��J$�p�:܋X��[P^��%�
���1������ >Y����d��we������=��?~I���[z����q��XplL�o��=D�ŚDI'X���ۛ�.���!l�Vk����n��=��e��'n�Ֆa��__�UTCQc��U������:u�Y�ԣ���ce�3[�O�0+q}ѽ�I:�{m����PK�y�d����Ԧ�G��p`��K���б�9khc�^���l�K4�3z��;����'�67��u�<�{�ϻ�H�߿O�?�i�`����2�|��g`�(��Q*�͍Tc���ҫO�>�xq�u��s�o��I�8{ge�;��7g+�5N�Zv�{R�jY��?�}u;G�ܯ:�ڟRyލ-��9�I�{^�_?����y��^�����sT&N���
`�\7�7�_�׾zs	+&�W]��v��u�q��sr#�uh;8���F0�`d�+�,�,!�4I��:��,���&�۷oc���O�`��8[�����m�i���-�ڙ�$baBO�>i����)�I�߼QEW�I`0(���0�1�Ё@-�U�>������訰�u58Y�5��|�Ȓm5-�b��o�?���ő��>@�x���o=��\������� n�q�~Y�P\cL��w,r(���X Q"HiK_�g���]�&��#&}c�M�Z��]�[vMKI]}~s�6�REŠ�t^���Z��Ht"V�0ͱ�Bmo�Y��J�a��C `��J���X�������-�[&t��;���X�5�z��t/_��L������wȦ�9UGw�1��p.$|܅ \��64v��C�z��@fe�R�K9l-pg���`��m��������X���x�A8��T�r�g�������y�qR�i�Z�2��2��ǅ��)��E=m-&�6#�$�����s� DN����/��:4�5��@��|�8
��=$ſ��F�s��vv����#�tI��nb]/�����F�7��2�1T����!�xy���@�u��g�t-sX	@�:�& !�]J�]�Ar ĞqF@B��q�d�b�%�@����*4&\��昳p�x��|`κpB�Y~?�pK�r��=�I[�U�u=���a���g@��������^>~�삐 ۲�S�YJ�o����2�*t��`�F�� q����=�OѦ��.�Y�:\|0@x�hQ�Z6Q��|��ASЂ3�;��9v���F�k5��ײ�j&���A�w��{9țW�X��/ӻw?xp�r��t��n��+�b��e^�%���%�5���b-S��^6k]6j*ʬ�'l `�|��b����,6~X�lԳ;���&�]�L�t�b����O��HXy�/�Of�L���R_���n����N�(Pu�B,����u��ۡ���L��w��\'vِY2}�Ҝ����wdߓ��2��ǰ�Z
���)�T�U�z��e�Į�=�T-�X����s�s�O�B2��b]�l 2F��[����]�պ��EAk�	�0�7�@����f�8��#�$&H�Z��T٦�`[G���S�aZ��N��7�i��V�����l?�(�
ΟЕʙ~���:��Z��6"�r���JC�>�'�L���X$��[P��g�g��Bq�����XŒ��Xkf�O�G�W��2���8�����g+���v��fi�z>s0��W�^����,�v�ث�Wx�浳����h�hϖ�����OĎ�\�)|rݚcY��o���<k{�ɻ��/2��;���TNк���ZH6����r�~�������G�׻��,!�C����4r|f�H8؜���~�)���~��s)�?�۷ڹ�þ\���'�7�h��d�����쬏�ƕ+3�G��z��zsf��	hund�f�VŊ×L�h�L������SA���|�,����kO��|�����rI賥9�~9�YE�� �����A���#�mzzs̈́��\#{ɇ(�1�[3��b��kGE�r,ƶ_b�>\�ƇQϤ�ca�j�K���Y�L�|�2�\0+ą�̟�AKt�@ k��=�
���{8�nBl�� �in�P�ho�	m�Ա�S��K~�~}����9��2�I9�s81N��[�d}�y�ʗ-r1��T[�T�+qʹu�\�fa�i�|���5`��۵C�֕�u�=� �6Ҿ���JsK��L��k��k�('����[ٸ�����uP�֎�^@Cq@�7�L�d��V<MS̓��wym`�Eȥ��mQ�J��Ƞ��,�s��������A�.����������;t)��{K蔃]tfI�9�F3U�	���Nا���[��~�cm�<7�䢅�>ZV��Os�[�����<r�d�$�s��F��{�'v�4���������c�/�ƾD��1�S���k��7����&؋�PR r�lnp�ch;�:U `��Ϳy^-�ֵ֖׼Ǽ1]�+~�h�YwmC�q��7��qq�n<(�	��dZ�U
0f>�Zn�{[J���W��#,�Sip�~����N�cS�>��r.��uK�-���~�V��s�/�R�d���P�i���DdYn��w����}>��S�{�\]�K^I��-�
B3�X;,C�b6�о>'ck�u��M�δ���[�	���V���>V��,H��� �G��8�����_x[���.V9�<H<�ͼg';����O?�K��_<Ӭ`�efLcS����1���.�g�m�'�BQ
8W�>)�����i�6|O���	%@��,��{��\8�3ڔg0�ls3�W�:�ӥ[��_0}b,��Ġ� c셸�#���sPծ�a$v�6�mǼ2=�s,�Z�C��,%�j��&��$ݚZ�;x�*�v����gg�j-��H�s�\������&�Z�J�әg9�5a��k���-2���&>���Kڭk�Bj:�g�fM��I��ew����l ��D`P�;��>���R���k�2|yi�T�^B��u��Lh	���������ڻ-��?�Y{Ҁ�ؾ�g�8��!�8i�,3���SE�Җ��^Ǎ��뮸�q�g�Nl�ے�v�/c@�OSg�$9��S�|+�bs�@7�?���3���o�gL��&M�j��Z/ o�_��|As�.1x��;����r^vN��:��Zg�	]-A�~�<�_�^3�oţL|f?�;�!Y@{����k�^�`G�)��dk'n�D�Ly�J�Ӊ�;g�X����{�{�5Li���xy�\������Q�9��e��,ؼ��i�>�@��KM�vc�,�x۸�����Ý-d�w�j��U��R��E��B�_i�	g�����sL,�qØ�87`眣�R���^�Atm�\��_�[u�k�k������§�^G�����䱥�4A�Ͻw�Mȍ�Zg{��M
��V�(nH旻;�0�©�y��A8�R��ւ�9��.�Gzn���Νg�دkⷆU]F��5C�MX���޻J�Q���|`�4:�P�b�����JI�D{{�]hQtB�9����J�H[��8Z�I��I�4�u�������/��挅����֚#�7�[Ə��]
�j*�h�t����S�R��u���e�o�q�y�k3ϝ������@�xv�3����jι]"Z-��u�S���0����ɹie^�%-0�~4
�q� �DC��-�@e�~�2�°�������2�����12F��	5'���<���8�.*P��j��f*��'E-�v�W^=oJQ/g��֚�`�����`Z�5�>Vז�U�s���T�uލE����Ywy��WS-hl?�������986G�V�Z��+�Oޕ¾`�' ��3����Nk�J� ���˛�,8�ce�W�L�~�*��z$͘	N�@xO��w�ݥ4�J8ȕy����P��{1U�D��c[�9t�l�`�U�Y���w��r�����Jt�Y$�[֘���B�ˀ�V�l.��Y�����.q��<�<����X���|T����s8�6��\;Fڬ��-�	��~r;�ܝ"�@r���1���t�2;j�S7����bK��< K���y�vì:�������	l�){)�����F�f���WF y��ac����*�  }�{�&�Hȯ�����[��)Qk�8|�y%&��0:IW=�� ܱ��8'�7��nˎ̐���g�sZ�͞��J���8�\�3�2u�j:\5s�]�*[i�x�t�d ��E���i"��q��-����|y:lDMg���T�Z�B먋2�o���y)V�V> �2���Hp�E��,I�i��3ٔb��.�Qy5-qf�(�h*�ޟ�Dm�띙q�Xڍ��xnɌ�$���}�	�C�yӊw?��¿R��6��M���I;��M�[	s�cwk-�;���{��3P���Wn(�qGu�3ƨ[kޕ��h�@���Jj1և���@^ӛ7G��8��7�q]ӽ��.�l�+���
�.���B�=מ��y����C�z��E�����^��}�"�~8F�D?ڔ?����j,�G/�B�4|��w`Yi�Ab^�KD��v0�f��#2*{Gw�i�n����l�֭�۪
\����sJ)F�Z�{��Y�#W?��(9���={���?V`�n(����B��h)����Ε����Q�,��A�6Z�\��_p�D�/,��9�e�Е�j��-�����-N�e4��?9��˵��T�du��t$:	䉎6�<%�6:��:��B�w%m��
�
hk�	��W����H��3$���d�4Osz1�suX�|�
��+]��cU�����^J�g�#^+�z��I�/�`ch�A�v���瀝oO� �
�ԡ�Tx��� v87WH����\��Z����)���U%�:A�-r�.{v�b��7�G��z_����V[١l3M)�I�G�MgՍ�?�Ti߼���>�+X�g��R��}MP+z�n��u�-�M�2<Y����ѳ�1�]���B���s�<~j�k7;9L��n~����<α�8�sHYQ�?f+���=J D��-(��r�����۲qTZ'P~��r�][�����w�vXyqG�Fq, }��}�����ɫ^��XJhK9���1�家2�sDf�e�=~0窲���@:�&��0cA��䧖T�;��)�?䨎j��<��3� �$����~Y��$���d������[�~N����fN�T�	n��CΠkrDW8u�Z;}���VJ?��y��ڂ,O�)�oP��I���_�������G�`䙀�(I2��Vv��8�5C汁��E�sX9��?}��p�$�:�EW��µ�U*�>����@��H���smK4_��,P;�d�ZrJ�#�b
�Zl����Go���j�C���
�
ݪsU|�R��R��.k0"�ta/d?OO;��m�.\�P�����(1IԲ���L��%�k�|x@I��W{�t�t�	O+l7q9�D �1_�'�K� U�5k�q�j��~� ��}����J�f�g�o�Cxµ�/�]�,�2f� ��������@���w_���$1X�6����;]/��8+���J������g�,m�d�C;g�M&Ʃ�Y�G�'�]�iρ�y��t�=cs�[�� �/�D^��VHY�icͽ�=,З*p�bn��������d�0��;��f\����-�8ο��U�*?vVgR�����4��/5��c:�R�x|��u�@��Θ��{��*���@��25I��W�X�jY�|s��*��4N6L��Ջ��n�k7���c��ssϘa�7c?J�՘�?Y���e���v2#��;h��~�}��ު�e�8k�T,�����3f�m���}���Q.~��#|�_~�u��ށ/��D%`���Tm�w���~�iW�kU��P�4w�U��[Y�r��!����RĪ�����+S��oJ��>�R.n[?�7T>O���YS�Ա`��w��mS�lH׉�:uf��?�(%nlr�Χ3�=_;�hUf���3̪4��1׎Ce!C�._@Y�ʴ,�堐��M� �DYp���D��fl9��z�k`�0 �wpJ���՘�Ɠ_iο��ƱEw�Ŧ��M���f��}p��N�ۖgǡ1&��7 i�U��}n�D���v��6ԙ	��%�4��y��]��As��i�5�.Hv�lt�̋mP�L�\LD-�0J�;{�=&fu2�<r`�L��T R�i�NX}�9:��j����c|�2�9U�#j�5��q���� ��Zn^������p>ZDY̕�(�k����qT��f��K�� �عl���8�ܬ���3����i�E�5�N���W;�Ql;��+�3�׏�W�9H/n_�<@y���}����y�f�	/z&퀒��{u5Ih������>Z|w�V�{��ӵ�ٺ���p*�&���eK���%)'�����Vp�K��`�2�h���D �%41�R�y8k�Tq1BĜ��4oJ�6��/:�Xv0������:+��c����r��=��?����y��g�E ����Ϙ���|����(`g���9Z�c�{`�.�^G�_�  ��a�P���:��"����Ĵ=PJ�%�xy��ǲ�V� ڿ�q+��M=��]2:����PA���4���޺4и�nB��
軞G�v���}�� (����� s n�F�@�/��5���!���$�7��9/��S���4'��nA�6x��~+�4��\$��i��H1qWn��DW�>�a�:&�B�lZpd�{�0S�@Ä��졿z�T9��_l���y��Y/����k���& ��ЀkG��Ao�S����JD�����g�5�vbg`̰�+`�����1:^�w�m����?�#Xl���y�1�̹g�0z��$ˉ�ǧ�>�7��w��Ϩ�]�=��-a/��RM�;ˏkp>�∮�1��>�=����?{BJ:@�L���&��Џs�z��ӛ�Y��M&�(��=�9#�T{�Ws$��+r��2���a mD��� �8َ{�5�}]��S�ne+N�&���#�da�ߺ�^.-��<�z�	#K�����Wg�[|i������(�V�R�p����¦�����j�|4_�:Z���v�k#�_W?{cc�������'N��@[��Ν~Y$�K{����-�ӓ���-������ N8��Q�=�Y\%�fw2��p�vt���])ڷR��ɋ�F��,�4�	�"8Y;��)K[�0&���M$6���)צ��E��(؝�JW0eX��x|]�/��s'.���S�A+`�����Χ&I[Jc���2ƍS��a�:���pP����F'��(�<u�!]�(�������;��ָ<��[�rs�ߘ���V��p��O��7����,�N#���f�%��T����;^�8;>_e�m~w����:��e;
;'e�ή���PK�v�f)��z:����b���6l$6��B L�-��ctd���C?g8C��xB���6)Ռ��2�~����![�5%#מ�5���k��MӜ�T� [ ��6gN��u��� �({�y�*�Bs�6��:[�t{��7O� ;�Y�>ГM� y����������� �]�}q�����% �۴��N�4ޘ��@������U�m�#�u�� ��=��K��(��m�s:�V�����4�vd/dޟ��Y�t�u�M�gw m��)�?	׍��8��{���&�\�9�S��ٯe��g�Ҙ;ۗobf��i=�kso�d����xEYF��)��A\%�r����\�W㥘�����6];Wq�����&��V����s��g���� �Cs�x�hYh��_�ސ]��kl	c��X�&����v��DV4ZPFQ��(+KX�r��hZh�ڀ�EJ�n����ǵ0�jv�`z)��~%�!Q���
5J��|ӡ�Ka�1j��9�麴����ڼ֖���դE��mY`|�l]���XV��"�Ώ�0�"j�y�#��:�1����&Y�e?�}y��[�>M��8�]���;�{z���u0�^�|��؍�$v��u
�2F����ϣ��J<�v���O)�9v�v�>�k� !��j�<W��	@�f�w_hK^���o)��.���-���s"9�l���������ψMv�p'&JP�](���J�<����;�.Y�Ļ���N�NFٌ"�S �掘ff�F�ꄖVqjn�ES������;&��=�A�l���o=)���m�|WoS�ꅗ�8���,(Y�@���X|�j���Fn2���El�[�.UV.�A�"H���e>h��Fb��铃�_���O�ӧϟ�Ml��*φҹ��������{�&G��L����YU�U˞Y�R�����c灏|!w���; ��-��T���Df5�V����n����W\�H#=�i�p���x/|oO��vrEb�u��@�A��"�� �%�f����#�A��s��a����5��!'����\I؄A���^�Xٴ�]�v8���UN��yO�"���V
a��
��/�x곢D��"C&4��҄fe�d�$�geS�$^�xC��$��Ч*�ϽĦ"�����W�Y]/s�6�ҏb��y#U��)5ó0�$��=�g��Y޼h�ZMp��h��IQ������	)���_;�r���l)����o}�n ڿ7�L�B�}M���
���>���s���"(F�P�״,��e�jped1k��/b5k��"���&��{b����7	�����Xz�^y���8_�4�`lTb����n��2v�DqW+Z�Ã��̲��I�,e�gOӬ9)D��pf�[<�z�3h�:�ߢn���)RAD�lе�yW��	C:�א�UW� @�=��!�Q��c(�c��0kY����G�`X�v�+��8�Ŷ.iR�6��lu^=��J����IqdoOA?Q}�L}�p*(zLx���&jZ7�
��y�ѽ)l�����a����Y<�&݂�7՜V�
��H8;5T�wv�<z"Pi�º���@B�7y����(e�;\��s'u�g�aז:	7:s�%V4�m
U���������v����	�����9�^z6
��(�|�2?Y@�e���М�
��㙯#�TF������-+,b�>�w��=|`/3��t6�g$��*��w������}W�2�I+߱煞6o���4��ؤ9�hlM�������A���5����ӣ�+�8cQ�O@�3�moYn�������]e\ψ�k
?���c�X�/JE�
Sr%��~y���p����?T�j�( �E�Vc�� ��He�	���\���_�A�!K pJ�j}ϓT �E���K�g)�Z.4G)j�5�3X<c$i��q1d�E�"g�.��6��.����ߥ��M��߸�9y��?�%g��Q�+ޘ�g���%9~�X��T�L,d TcC3�Mρ��*��9�����	F3��p-9T���x��">/ንe0IM!!Ǵħ̭���p d�{��|�e@������D@��48>�L�D9�>}��_��TM���j�y>2O*J;�A<i�m��\-�iG�L���ːl������!����h|OO����&M�\G�8����������s��d]����K�̋.<y�1)2��ᰆ/ыpm4�᜸�=;O6d��^O�@l5֍������u ���������4[���SJ�H�D�H��Ad�2�S{/b7�y�T�Fm�׏6>i�o�·�! ���w(x%�s�c1�~�p]�����A� s9�u���T3�4c7[�[5'qM{~�r���M�C���FF}u�Z`Ѹ cU%S@��� Y�i��ƺ��\$������Pd�~~�d�"33�\�=tɧ�2�_�\��Yv[\��ϯ}�M�	V2�L�C?�z�1@����2��?H��m��������tg��ǹ��v?��k���u���B�>o�
�C�Ȣ�᰹�k{��d�����XޘA}9�,�bQ��CH�[5���bR�
R���O�a��8T��"ڱ�E�3�PÁ��]k3��V�p�4Ϊt �2gv[�0�T�SG�
���O���y\�ݖն���:\��wô��BH��>�I-?T��Q����T9���=�+.l��C�mT� �z����������y��>%gT|(.H�J�'C��Bj%�7R�+ &�^�h�F?2����B�L-��k�k%?G�P@`t����Cg$�u��(�d�%�Bl�5.aj۹�UINi��#�UbUU8ɯ%`�ҘHK&G���y����V�E¾X٘��xM~XL��X�ҔR���B��Q`�AI�_��>�͌߷
�?ا��EN�<��ז�:�� �Q�5���M|��P#ߖ<*^S�w߆1̬@�Ya�,rH�R"�aWƷh��gK�z4t���#�L����(���G����΃Z�A&�Vu��
�8K~_�&�x<bl�����X�~��+HЬ7x�� C�T�׶�Xȳ\�&%�{0g� ���SDq���L��l��-�^x�I��$�s��<��.�q�g&͋��Q�+J���p`E�*=�z�����r]J�l�GB���9���ե�q����l9/�T ^���* �RA��s��Q�X�y�
n�uC�Y����6���/���Kh.�8OOi��Y*c��*t�^���ma�F���bL���:�sG|��c
~g<�����Q�p�2>�>S�{`�ix���e0Z���I������=s�[3�HT��dLI
���>|��<m<I���W��E���;D(����tz sw�QZ�+�^J�J��O�t����a`��ʗ�S̒�k�s�G�j�'�x$_h�`���*��4�<��2+�a� ��k���]�7N8��8yV�;#^߶t6v�.���g�_��A��7�d�DH�Z!@�plW�3��x᳏b<�Mbd )�u+<��1D9薊�T���F$L�fX �C�9�:�_,�!§3;���<r���u�1����0Dx�9ĵ��X-5��*�����ҍ�\9����Q�5,>��9�����b����j�I���P��t��<�S}|�fQK� q�*.Ϛ�_��_����K�mz���"1Ψ�qfk�b��Ѹ�^r����Vxy��"}l��߷���	�a��C���y��X��=��ԝ��xk�	�![LSSl��� O/C���2n@)��x�D�*�a��G,Kƨ�k��LꝗX�s�(C%E�;RT0�k[qʲ��W�S:@�<sYn��>p�F����!����4oU�������ȕ��(!,X8 �y]*y.���Bݢ�<o/�ک�B9�p������CɁ;�jV�%��$�v���S�ٱ�/�	ˢ�}JFGB�r�*3Mѵ�_�=�������4/ysM���HQ��Q��D/�H����)\�}�'��ؓF��yM%����@9w��cY)i>��j](Y���3g�4�&�k�F-���$�Lz�d��\$gH�������B���������7��Lcyo�vZN�|_��^�7Y!��}2�q��{g�M�j7�3z�F��8�Z�j��}��c,��:yrTΗ�`g	���uU�v7<3�1_v�ZR���@p�� s�q4�r^�Z!�y���]�D �f0�V?�/'	��e�R�vJp��Yʏ��5����p��a��OR~�/��x���݁���֖sJ\���J��PiN�'�
�d��#݃�D���P�C2f�hu�Bn���}z��
�tT�bE����N���b�51*D9;����� ;2��*�sBq��l��}VOâ��}���Ea�y���*B�
L�W�!���4�V�HG*�&}���F�iV/ ��C�e�%���tz�<�t�Z:�3$�,�(�Y�j�-ˬ�������Xi�Y �����h�~���Ij����|�����.a> _�����0��A���pkֻB=Dj�VV�4�4��]�;[�7@����R�_���ᓽ��:8�kF��S�FCh�e��ٳ�˼�d�Ť��ub�K��H�.޾�X]�{�I5���U�
N�qV��z߽K���{z���L�F��6�ޕ?k�S�44� d=�b����z� 5����?���AC
!�
�Sy���˯�ˋ�̋��N�>�A��B��M��{J�Oԟ8��Z�W]�w(LԦ�oH2xc����ݢ���i�U�&y��EA�� �G��l����8jB����2�sH��(��������s���S|�$ܮ���l!�zv��#��\�"�5�"N����=�U��9쭗[m��֊��SI5�W�Z�w^���f ��t۴H(�Y�YD��ed�/���:����}����T/W�lDZUH�.���&K����1�X!)��Z��,Q�|�=B����R���(a	d��=|r�9���r�׬��c[)��<�P�ܯ��?�f��~XIܥ��؄��s ����[)�߃���Hm�Z V�Ӳ4�}p�ފ�;+{�I�4(X7W�pY���f�V΃0�G��X�,����jT13%��c����Ĵ؛�;�%��1b�k�HЫ(Q'^g]�W!Y\{>6h��� Y 0�� F���X��aJ[�G+�m�I[�+FV�gf� ^L2"P.CU��=
p�8;T��(PR_!(�P�Z���E����y��n����/G(��X����*`��Ja:���o�o��iV�%74"�=�r$�t�0(��I�wa= �� �>_T�������>dQpfI��n�yS}27y䘁�\49��`�l��:/���*�7�,�{�K�	����JVr]��[ �5��/����:ڤ��Zӽ'�.�LR��Ӟ9�}�"l�X>����F�������"!��B9����)J�,|p��.�VLcUe��UJ�J�:a�f��ːS"�iY<3mIz�%�e:��8v/�N}��а�3?)R�7D�YYC�����:E9���%9����9�\�� ��ʨHp��(�"l&ʶ[�K�#��Q8���|�y��X�d�����K�3
O��&�N�L���(</n���UT0�ġ��s<~��8�I@��^6��^��i��U�+*���L?X�N[i�?����gɌ���	8W��E�a��e	jQ����P]Ph���7̒�u�]�@ z�n7��W`��M�Y��x%K?��ږ�����������g��y��0�Ng���>�t��0&<L�lH�t���^��|/�E �*�3=��� xgΏ�T:��9��*�R�)2��1�WU�5��4�L�[Ձl���|qÿx��|�=D���!�3�z��\���9���-�"����j4�?pp={୆�q.PV���N �{�-���������k�ޒ0�M� �Xo��qy�<y��nd��ʪYe�e����(^���y���PU���|�2o&{�?9��W�=ݍ��x��ٲ�҂@`�#�}�P !�9�*dD�u�M6H���ޓ�r����n���������ځ�:ZM �����w�`���Xr�ˑ�!��2ku/��ݽ5�O��!�7>$��ǯn4���s�8��}8~��d����������1*>(s���r�}p�)�W�� �p�:){F�+~�o�?�i/dxτ���3���.�Pc":[�*�c�H����'�p��9v��˯v��͵��ZrG��>�ə#��GU�N"����p
���C>i��P�BR2(�����O�r�1q���$��i��hoT����?h0z���a��������ow�3��hi7V:�!m��f�1�v��)�|ъgvM�׉��~`&(�+V�_� ������ 	{댬��ҫ��G��EϤ��o�y���Ye���V��!ڣ7��9D��b�6�9�M<�����х
��_�z�/���yJ��I��#ywjP�T�H���v����2��;%��P�O(��g"yY��~��e:&E�\p��W��<��u�;U\)\�rJ(�6o��g�t����t� ���d󖒖�����D��s���aة:��,uNr���&'��(���9s>2�9���_�X���T����K-G�b� ���#���9��@t�%�E�� ��g�/�����E���^\�PK�}(�B����T	��"�b��%:ߑu���B��J�^��� �b+���oY��_4 D 2iT�y��6��:N�� ��%{��k	�
�mTC�"��E�p;¾s������@t/���zBɚ�A<	&��G�؛�o������!EL��t�T~Dya �E��Y�UrI���qQ�YB��S��vx�r� ��5��I���$�H󚥣X9�g������b@�)��u������f��<�Q����:��{R��i;��~	����d�Y���<m�6nE���"=�ШȩA���pR��tٳ��o�
���|9���C�-�o}IE�%��Uo�9�p����¹k 9�忍�^��� �e�r�k�R,\�+ɰ?|Ho�����A÷��������&��X�"#����bKOg_U�ַ���R�?劣�ӆɿ�Nۈ����|�ߜuA�F;�	.��r���j]-����q���A���+h���*���#�h�vX���n�$08��"؂)�k�y�j#`ݡ� ���}��w���[�u߬��3d�j ��֢O ��,H���#l)!�⥿�b��o�}`.��
%��)9��A��B#�Bt ��[��9���ػ�ڒ���|���/��(sv �@W஼��:
��pE�J��a.�E붍kж�]�hٟ�&P>� F��P
���r������}����9�=K�6B�4ǉ�>�^ ;&��Z�z���܏r�(��=���Vn�D��U�o �l	!�Պԡ��X~�Ԏ^ы�Jt���s'��O��vGˤ�sD����<ۥ��Vü��Ҁ�U����0�5X@E\Y�P��8���P�B��9�����7Ue�-�ԏ�i�y���Qx�I+ҵ��i�����^n��z��Ob(��E�|8!��O�Y�\*ʙ����)
�$����3W貱$�V�2�z4��H-�Ƴ�.}En�v�%���5�}i�
.���!F���1-66�'dD��ů��/)�L_[���X�t���
�󥭆�D� �J&�A���EN��x#������9q��>(�,1+$gʡ3��>���z�J�9aOHrgxY5��$�n�+^o����0��#��F;�>|�Eʇ�L�ӣTZS�h��AH	#db�2Ģ�G~�^H�ʲ��@�]����س;2�WOЯ+�ֽ1�aE ��kv/����t�% N,i��:2L���@q(&������tR�U�R�7<�8C9��yJ*�y�*ΜY�i��A<�O�sS@��.���tJ�;Ue#��Bќ{%WM��z� �����̋�Ka/�� �OaTP�N 4�g�� �u���<�*ψ���r�Κs���I��#��0I�zyhr�J��f{^��4zء��s�2���y� TD�R�;n�;.7��l����(��/��(9ߒ�����Ž� 'X�H� c�r��v��W�����Ⴭ%�WRc�)}�DT��6��7 �=��0O��h��sf���9[Z�TD��@j)S~y���� �(3�r%��㕺=/�������	i�� � d���k�1��W�����-��ߤWtZ3L��A-ف[���I :��*4��Q~ⲹU���﯍�n\a�%��K��Wn����֧�����M�&�}�� I�`��r�5iV����� /�%y��͠;�Uh��1�M^]��aq᚛Ƭ礊+�0C��e@[�W*?��򓳗�4!1��E�ݰ(�.L�
�ʇm�#[�B��
6"��
��/k=�A��g�2��
S0ׂ��[���N�G��Ú�ɕ���LT�E ��M(�+�2�[}�s�0�^��5�����bc�W� zK (I�<�>���O\n�����O���׬�{��G�_��yNF�M0���Y��WU#-H�?E����'�>�Z�kPF@��C�▩�喠C�x>==�r2 PlZ�%�=����[Z�*E�֚�B{P	A�H$�P'��f]*��Ґ��!�#��<w�9���6�"�{~&���3���tW4/cԐ��VI�M�8�}��߬ը��8�vp�=91������3X���JDאRQ�+�'�T�AsSTST%�K���#W�E��6�����VJ^"�Օj=v�P|�D�4�� �^+�֋��3W�U���B$��X��U�+}iۢ��My��B�Kk~�(���C���3�|+ǎ�R�j������h�U����A��K�����|T���,Nw�����z9�I+X��"�o�G
���_��0i#j�����s��fI�I�9{����݃�~~���f/;��`�RB.a:&��������1}೹&فc�;�|F�<7�y�֞������-��K��x ����S��<Y�F��Ɋ�4�>�Cz|Z�=h9{�U�kU�Z@��7o /�cOO��t�T�Zd�X�9�{V`�~�{,w|6�x�� �?V�G��Ā�p��9 ELX�H�3\hL<I��:3�R�����M:�_���A��ϧ#{�1`�`��<�|��e�q<#�T�v�	!WU���C
<��.D��TI�~^�mA��������(�֫yk�ݠ�V�s$�2�	�|�&_s��t�y��Le	��ꍗu���Fr�~��|��gB�Z4�S�$>�����ާg���ܐ^EMr�5f�W�y"�x�}�s����K��ޜ�<����T}����������#�4��ǇW,_0}/U�y6�ϟOܯA=��
'�5�lw��Y
c_������;F�|i�s5yrw^�1�D�H3��#
�"�yL ��L.�h{��i��;�g�uC��}v�<n}�>%��L�-�I��'$�l(�S�D,/�ƛ��`d�O~����6�\M�%뽸�J(��ȁ��qHZY��V�ͳ�bT�:kV�x��.�Q�0N�R��`�ݘt<!�=(�8�na�_�������!;e̸ v�^E�y���`����熾_�]W���M�ݵr��>wo��������w��k=���z���(�?N�7&U.�՗�?̼i?�b��\W牁�.���@c/VŇ��(a�e@"1TX�cu`��,���� �^p���ӧcz��sGJ�&[cT�Ż�-5�h�-k����ĵ�k�!.�gK�<��C���)�#��k]`�:��]���-��{�B�[~�����U�?�yT��������������  ��IDAT�\����E�|�mz��K�J����1頡�)a�kC��baH9�"�K��]Ҥ��q��A��`��xM���IϢy9�U6e�=hM����H�X��-�Ҁ�E�堿�1r����Vn�I-����<�5K��T �z~7��K��<�-�w׮�87�L__�	yb�z{O
���b|����,f� ���ڬ�i$��s�z;L^+*�� �@��JW����95qg],�0��}�d�Y����ʠT�E�v�<`Qi%E55t���4����u6~��=(���ޚ�{���z��}������k���H��TSi�ρ}����b��V�w���/=��l���lݫ�y3��Nî�Q��ݣ��>�,�x1����;K
>r�v��������蠑h!UL[Y=B�$��-�/G2�Y�q͕���$N�o��;�(��d�ӧ�b$Xf���`����C�"�_�<P��� ��
�{��e�`��J��� �D0�{लB����-y_5�;Ag��F8�,)�޲�Ai�l�w,fl���OZm�@�Ys�`�Mg�2E���A��z��L_�=�C�;<�����,�R�2���^��8�W2��$�\lY�iP��ũ8�ee�&>#��{T\�Kz|���6�Zg^PP�D�=��AW�v�=�3Bf��0H<�U�x�#`�Eе�{�*mi�2�{���:�7u��.5L��ͼ�w	:��Z�0(X�`�&FC�&,BY���]��U�pI28ϒ\�K'0Y ������pE,���xR�h��#"��n��,��s��S-AY���3@s�R���� �>[�z�!P^�(Չ��֥��6?^jF ul~�⹷�u�A���BR/H��F|�׷�q��OxG���3���P�2�����u��|���:bx�Zu�A��J���!@�K(��P��Y�$	�(�ق�Mc���0\�n�&a�	}��+�9[hֆCJ�Q��溏��+	;�C����|���K���T�����hA��Q(R�N4ק��?���r��q�+(.ܼt� ��j�54�0OJSɁ��%8�@E+J 9x�x�I��_uP'�Yr�,��] 4e��@�Y�|}���"3D��r�S�5�駟y�dy�P�}P��zE%��G#)�*��Z��	,wK��V�I�T�S�+�-!9���9/���y:]��϶.U�0�`ت��-C��е�BΜ��CI4��(ʎ)�5Y�UY�E�Y�5=�Ҷ���� ^��J֩�y�
(���X�^1O�M���X��Ukm΋��0�1y��φPۏ�Z5(N����,e������ga���U���	�F�"���!���SQ5@��*V͓u�5�Q����r+T�����&�A���wo/J�o����,�+��A!��S.�3~�MI+e�p-�9�����_#�*�����"=r� Lx�n�dѺf�*������&z�)I%�;��Q��ٟ���*9m��bjϗ¡v�jDC�yq�� �:������uR���q��*��C\hEGx��z720�@�z�K���独A^�b0��*�IRM.1�@��y4~���������)���+�3o^?rX"�/���U�����3ī���&�~�
f�h��fRh#w4��Уf�i(�������
�������Ct����ވy�F=���f 5T�)�׎����p�����y�P��O�)$ %���}�}����?=~b�;s��%���O8b��R���N��R���Q� �F��I�u_x/����L��㯿���}��:(�5Y0��k��0{~1N';I1 T�mu��
�i+��]���k��+���	��e�԰B�r�2��ʂ���Q���σFT]7�(�m�7��5���̍P�M̾@��$i�
��e�mr ����#i�c"U����䦉	�������k�^��	`L��CPڋX�$ߤ��lH��KP�eL�E�u��J��'�tS��T'���''�Z)aB�k��#H����jv�Y=��KD%_�d��۹�S��}C�wY_��6G��{��'[�'=�FE��X�`��=����]˪��@�k��5Jݾ�SnhH�J�I�V���G
и.�ۃU_�Z���$�%5�ϔ��	Y��P-$��=$�z�"�`���⠎��e�~��4��e�x�e�6�؇�&P& �<uD�����D>��Ş�;D�	^8	
xh�~֒�dȲ�����U��ќs����C_�[P��ėSk��J��<��v�>���e�ˎ.�5�,cQ(�{�r������ ���ȉ����Ăې>C ޤ�sJ0��e�������fwE���̔�BY��c�� w����Uq^(�8Z^9�Rn�_�&p�^�fL�4��9o���s�4S�"^(��Mi/�
��@����L���3���/ԃz��ܱ���y`�|e�Q�^~P�HZ;�0�=H׍��3۪W���Z���&a���
{�A�-οSRB����sz��W�9���)mHVl��j�����@K����l����� #G��*e�������9�/�ɇˋ,�dI��f^	0����Q�?��hij��(�� *�5��ᱳ��k����a�"_fN�M�uzy��~���U�K!?N��+R=��2X[9	g��MUV��J໨y&�W˘��afRɧX�q>��.�\L�����s�����hj�r���%�'	���뗽T�:(�c�x�뜭�ŌU�}�y��8K̀\5�
�:CW}駟~a���w�L4퉇G�I�[00��P$aNH�z�ٙ���Y�Y.G��b���˼c�V�EZ@�QO��?	�Z���Ș���A�������k��2v��嬠� 6b �2)?����= ���%%%�r����H0C�N2�fƌ��Ղ;a.z]��9��-�&��g-w��RB���t��_�Ͽ��~{�>����C���(�c�H�?=�B�$���JU��F���j�%��6�����_{B���v?�Wt3�ݖ�T���k7/��(�Z%Ф�)��OR�1���w.�f�a��|���8&LT7R���Ꞻ�#�悠IPf�v	P�~-:@�@��Ɏ��ֆP���Ie$��IM%���h�����ӟ��g�QH���x�s(K��0��>sF�s:NG��0�Q��>�u9��rq�+�O�$}�����%3�1܃���x#zL�T"�Y�w��`�)������P��DOì����>o��I]��z�,���m\�f��[�`��5�7�ւa��B\cz�� $�����W�P�k����Ow�lp�|��ݛ��{�������"d"F��B8>����\�M�6�~�m �nN��B���3c�)��Fgj��R���&܎��bi�Q�p[��R��(�}2HաY]2��J��a�D��J"�� T٭�19{
�tuW�.��âT��R�Qu�O�-f�@��:L�=���.Q�7�/X�,PR���O�����=16W0d�Op���ۃ�fЪl��$=��n�.X��Z���,9OG`��w�	eP�x�"s��âژ���|�a�.�;ˬJM��g�;����Ǐ�`/'u�ƲBa��@E�9�*�4��jc��W�ˬߣ�s��#��W�[#��M�;&	2E��Փ�[U�w� ����9La�g��f^��5��%ѤV�1r��6DÙ����,�
����ŲF��]Q� ���X��0	ͅ����2��`��3W�\��H�@�5����!����U[(�L0GN2
�����Փ�F�am�z��cfŅ�������%�����?q.=��Ӑ�0���k ງ+�����%�S�P���z/������f Y���Z�1a_X)�hq��JzM&d�Մ
@lW����4�<���:��[l��JSl�ü�w.�q~�ɳ$�0,2� ɞ3��2�4��G*V�A�M��<L�$��?GZ%-) %�N��[P=wa:u�C,�r�d����x�Q�E�����sb7��)��o�4�V��i�Ξ�,oi���CIPN�[�������=F>�b_�%����ۿ���*�x����2�>7�f��ULޖ(�%�iFl��Ϭw�W���e]ɰ����˹�^]^�o%�O�F��c���);/7��g�IU9Y{8Zо8���ʩUs�M�<��%G�~����������ӇO��<��������
Z��a����"��	���S��b��hN��2�C�~�� ZC�ׯ�G���V�]��9z���p��
����f�;4#��Z�d�$�-9�JeQkS5Z����æ$�'q[��%�B�X��C����]+L�xW���N�{�����x��`N�>ؤB��'���H���!����^:���WZά<y�<��������s����>ɛ����J$����� �?HJypv��M�]Ik�L��G�1-��$P�=pho0��=wV�=��L��6�Xу:Ѣ���G�^Z��>w��ej/i�>熹�]������\����/��=�,�3��E�A�V�XO��Rў�C�D��t��+b��*��e��<�>y� �� (>Sg�`��r�sk��5�u�*��<�TO	�qJ,���ˢ	fsz�
`=�E��~�<�+u��}�y�/�]~��y�1㰵w����w\�@s�7h'(Mk��i�?��;�?����5X���>>f�wV�LRl1���t%�ab�N^;$xǮ�Yݑ�ɔӆ_er��b�7ev��V���˔���7�!!�1��V~�����l�\��Z<�%Ɗ,	L�г��*ct�^ۡ�{(�V9E�5��M�%R��m��Јu��Ġ.��PA�+�7���~��3{t�?zvf�c6�}0]K|͌C��#��@��Y:ƞЯ��ϰ}�t��zC��`�cE��$����aP^���\���!�i{��|��3+:��cG,�ѳ���tRF���IYsuUWY.���&��8�1}������a��t�կ 4�L�H�1�u�27��k�_Sҷ���[���׷����;=����}�н�ʋ���*�W���zNәO%�kv��< �*���s�K!/D�����K�ex��<uf3j�\d9X���Umμ�E`Gh�r���M�5���C}���t��nȈ�TY�9����jIo�衧�ԹO�kypIb@[Vt��{���D�5�wѽr���m{�-q���=�~7����ң�wQYs��8ZG�l�������>W�+�R;H�E~`T�̌�{3>T�yGM��_�f����n�N2�R.��ϧtb#��~V������p$!Z!<ҧ�e/�X_�p�t�����eU�Y��/l
}ܼ&a:KM.[o�}
��y,1^�=�@{�KQ�w
L~��d�������u3TETӲS�tW�h�L޼y�����X�\6����`����@µZ^�B}���zr�^0��kR_�Zݳ�le3�$�i��U���
A �t�n�~�K�Ÿ�o:^N4]�3yK�������j7�/y�>{�ND�{`G���i�3Z���6������ ����5������P�;�[P�,,��^������T
�-XO`�^�S�e�E(] ]/d���;z�?t� ��̳&��HB)�ٓ*���v<�U�� !V�{�9i��A+�<h�%�FB��N��
W��O�a��mZ�Wa�w���F޴�Y�k��x�}�!�]!���K�t���^b�R(��2qI�a���Yʕr)��}��A9R�G�QQƫ�]��s���ʕҵ��}�`�&H�pE�
�-��˘��[B0������,!oDKD[���1�^/V��r���nU���I�T������rU��aAE�1l�-5���f���?��p�*HՏL���ͷ��˚[P��� @`^�I��(
e<#8@tB
����	ҩ�y�X7!w�W�6�u�<����/<\e�|��$f���1����yV�e�
C�>�(.{�p�H��bΡHx�(�t�r�����ζ�^<����i�u�n�]���ߙϯ��Ĩ�:�'�n=�P�<X�t��0*N�zQ�߽{��<�z�j�d�y` �o6��9 G���d�����G�k�[gN����	�O�a$c�pX2*sP�Te�L	���_-Z��as�� �]?������0���{�N4V�ۧ{Zܛ��[��q}���W
 �D��N���z%}x�|>'���k͠�e�	��|�S����� _,���
}�� ���ৢ�I�a�t�_���~~��Ο/��ߏdD]�����8���<MI�����!V�Ȗ~�3~�4����_����-���Ͼ�݅t�;�=F�����T�A��E��oE' �� LP�H*�F���*���ݠ�d����B�g_i`^�W4,*�"��+�_��q��:h25�M�%"�A!ʑ�@��W� ��٭�X*9�eH6L��d�Hq�ؑ���Xy���>�����+�zO���ư�����kǙ�lZ�Cz%`n�o���|�m���h����D�kg)�!JE��:��D�GV�
9Y8��N�ƒY��u�5��x�g�xw��cF�T��1k����4:T'X���2N$������i�]����Cs/�਄#��[%m��=�Y��-V��p��Yn�ڦ���_y}E�Wƶ	��Mұz����b~��^�c���Q��i� �i�Q�DT�2`��j2iy�/�ר��p^ZH��V�+j� O�#{MrV��g��Ȗ��y����sQ�(�&�z�aEA��	N�o|�>��� L8��E(�~��O_�%�%�He5Q*	 �pN��;�x�u���4���ݎ#ܶ*��ږ�	��*ݒ0��<'Q<%q1���8T���v$7�z>�R,
��ᡳ�K��J�Ҟ!p�ǀ4癁����r��g�����G�|
�(J�hѩd4��^���I�n�ԍ���aL/���� c����V����!#��Mx�������kz����.��t��,x[�?�j�{a L�C����EQoz�[~3��@C^��֨��H��^�̓�r}��R`���|�O2�L�m���HBV�Ʉ��	����k ������o�[ �J��[����!��\dFV;C.?���>�D�;yjW�=$��y�\��;����d�]2c����V��(��h�3-���+���B%� ;'6(�.��'
aT@��2�d���2lE� {o!zeNQ~s�?�R�wm��\Q�pD���vn�/e�d�j������Y2�*��3:�ߋ;{P����/��?{N�w�qm�c�R��z������}��A��uX�QƐ�5���ƥ8��j"�>UĪ�H�+Y��B�9������V�Mq�y01�\F����	3<�.�-�<��+�_ڲE�$WNE��ӲO��޾�]l��������E!�i����MI��6-(�6���6�у;��{{��3�k߹Ǔ�	B?�O�k��,�D����U���� ����ż���|E��8�
`�͘�䓠�X��e"�M�P%=�S��]->`�F �|㚜M�qP
!"&l�X�V�
Jtu,�,��4�v��g�J������-���@�]�牠C��7�����~�@�6r�@��IF�����Q�PqmQ`��j9��Q���64���,��r"�!�A@W`��|N�S�Ĳ�Ҵ��&�ZQ>/�^����ϑ���d ;rq�? hs�?s����c�Yd�kl�Qt)����z�����WZ��
��?��9��C��}<dee�\���V�3H�p|~NH�\�BMa"*}y�Ϗ�TF�;J
��p�.r��kJ��1�@�ʬQ_�N���G�S��*c�@��#�>[�j��d,�x�����>�a�{g�-@� v�5\�3�R�ڶu����]�[�t������(�Dq��4ě���z4�YX�B�����82�e*Rp>�ϟ���9��(��;%��a`� ��4x \�#�1Dͽ:�k�C�����_g�|����`���/���QǼ)5�ɟb�v��'7�6�vpN�;��{}�=j�d�/iͷ��a)�0&!Y85��8`��_��!x	
����T�:�ݐ��)����!�л�^��.E�r��᭚t؊�TD�8 ��oN��U╶X�";E�G���9�:��#9 '���|���E�m�S.�Ec�?䆲�����h���4;�C�.Ǻ��}�n��T�
�zk�ץ���Z=�%�������U���G��RG��s�k���k����0_��LR�.�WÏ��Zy������.����9�3ob
k�8lD�mr�����bJԽZ���87ﱋ�&
�K�,n��6�!��AI��k(�)�������7�e���������IF���N�`�wu#�RG�5&�M��0����&^wَ��>F�E/#T�������^Z#���-�蚠ۿf����`��ω�ؓA���(�Z�8�5%�H5�^�)Ik�N[T6S;{`mI3%��/K�T������ªP=	� �P��0�<��(I@�~$S����@�s#lm�gjh(�s7Zl��'��yMr�sy��о�G����}�{����{g��0"�jQ��RN~�em���Latg�h�G~�|�WF�'Շ�i���I�������* ���{���*	��Xnyy�C:3�^���J�U!�s;�ϭ
��{�/�9�
M�B�x��Sp���������|~R���2��Y�,�Y6��mz��Ssu���U����Ց�bo���<�(�N�PmI�x�aU�P6��>;	�Z��*R��Q��[L^�ճ+�g��UT��QEc���\ٕo�&Țp��(�2|$L�,^��h�xDr���K�n�q�sr�L�F7�Gý�Lm��@��{]��ʴ��
%�L��r�������Qs��9g���Cb����s]'I$�C��U�2�'FL�n�xX�qe͋�Y7�zU=���}g������w	=�:?^�G��p��!�����֢"q߭ql�m��3d������w���[���>��ye=��R�����l<H��k{������O����	��$�L�6�v��:�Y˼S�¤���q�O�A����`c ���;�效�V&1,@_���t:�T������$J�'�����LV�9A��n'���8�4вKy��Ys��М��?���mYs��g]�ӠG>S�{�z�-�|�ou�P/�.�.�Ƕᱣwb��Z��-�]�o|^! ��m�A�)E������T�U>�� ��6-Wβ�A\�X�X�)i6�[=�ժ�0�*Z�G�x:N�.�)�/eu�W��؁%J��bK$
�b�٠a�Y�ᰒ��q���k��L�H�&��Q-
�[��`X���[mعgC�Y-� ��f�9 ��^� ��Ϯ2��)%���-Z n0]�����\'r[>���C)DM��A���\,�}��oE�����H�I��w6�Q-��s�XyT$�.��B��9\%�B=K��(�H@5,xH�����WB��C#���"k#�z)i1E;���M (�/������n�/���T5���5I�=s_냺X��Q���Eϭi��ee�!)��E{֪mW:�`��?��5҆��^M�� Qk��l%�월2�&��X�������+S�k��z�*��"�=hlOO�����א�_�O y���P��;9��0�A���JXZ�\�h���X_�)G�珟8� �9=$�+I+{͚Wj��JjN�����V]�V��s%��}=��E���,��
�T��z�= �l����]�U�5an�
C$ם��{=>P)b	�b�6�=��K��^Y޺��~Y�������k�qԉ�'B��z�
�LZ���Z߾}�>_~F�8�0�)x�X~�Z��ś"�9��!�Tے/�3��`�AI	c�㱙�r�)�@5�R^ ���`�]��ŎN��� ��\%��rW=H5�(��m�k^e���=P'~Fm����r��$9x�Bы��}P���[2PqY�ǧ����xE_��!�Ζ�����������FO-	�B��C��$�,
�����_��n#Du���e69���*_��cg�����{Lf�gȏ
�2�Cc��u8b�8���bǺ�M��ؑ+��6v�Y�z�ɍ�~���ך]�%���@��޺�*�������e���οX̩_-�_K�,3�J2$��Ɉ�T�vAo�����MKr��SD�@X�[;��>S��X�`V�f���C���I��M8�꺋ċ9o1�%��{�u�@�`n��j��˯�۶���_3&���s�#�wUq&gM���2� ������lM���䬓�X1.Jt�t�P�W�d��D:#���C{�ܙ�o��G/��&X@{_X����d�鳽�<+�a�/���5QQ�Ͱ������K4�oRe��"�G��
�4o�46WRΘ���m���Ca���jc�)؋��\,?�rM��Ft҃�{B��Kт����G�G�	�=�|є��&�ȸ�}�'��������ݺv�œ0��������LTh��=�Oa�Ֆ�f:��!�f�k�*��j^ ���ݥsC�-�gU汳le �O���� � �pep�T�-�P'���]�[U�C�;�3���)Wzm/��5���$��3X�;2[�l �0�����v��º�kR��)�E,�Xj:��^��0TR�R����j/�u�[��xc�~u�YgR����*���O�a;J���`@wr�W:I�?��[%^M"�FO���ˏP���K���<�b<q�`��Ey;�`.>(.k�	�{�� +Q�y�>��Z,B�Fȋϛ*@��03M��kS���w�n�^�^
�gH��~��n�K��SB8QO�[J~ߟ���+���s�����%{�rX��&�:�F*:¹�׊z�b�'�\�`��\���9���r���8x������o���)���,(^y��'���(W�h\��+b���$�����Ya�t�ޓ���
��{�fO��㙠�8�5��a� ,�������Ɣ�w^��X���0U����:���t^����3�HնA~g��R=/���̼�£�NiRAЅ���3��	�
�u��ݫ�	Os�`Kz>��,�����"�d�C�!�<�ȹZT,��4S�X�-�`[�+��h-O�i�j���oύ�:�S�B#��Us�����"��d�x@�O��.���f����p�*;5Ɂ����P�Q2n�AЙ�;�3���l&k��~Ugh%{k�L�f�٫p0S)����1{Rb�l+ڴb�<�	�B5��M�k"j��`
	!�G%��II}Uxyȡu#Go�hA?b�(�1˿�H�V�PK(u�u964vHL؛T@L�s��a�Z���jJy����z�p��swsw*mb]�����v�2��q$A�>�Ȫ��Z� Za�M�!pB.�KuYS�a;�]��6;���<�i(uOm}���E�C�����$$7O�s:���r�X��*c��0`	-�jA��7��פ��'�%>��'����5��Q�)��,���TK�	��	J�tÅ�-!�-�*$��q���bc��S-�$�)H1WCo��p0�	d,�5�mC8�>��#_�����EY�u�<,ڛ�l�
���j�
!�la�N�M�CEYSⓠ�9	�ι?jU�R����o�Sɀ	 I�.�`��=��9{^��]��3�&I��Mi
a�I��i���%�XH\�dX3�Y4i���k���P����S��s�����nJ��/�<�|q��
:�@zo�Q�dY�?zol��fK����*�������g[}%� ��d�>Bp�H!aYua��yr�ęJ�Հ�l RMF��u�� } Z0Dok� �L��n^�s,U}��ȉ����V����յh��[��D5�U�Ķ-��'��k-~�'j��Zũ�_T
,wM8��+(�r����)�;#I�L�-`�+糝Y7�S�C�<Q�$O�ɽ���(�"���)��J??�ޒY�%��[��y�꥘��r�؉�Y'���^��ܢ�3���.ɖ�����\\
؍�������Lu'�:�/������޺���ne�x������]�{�����!o]�
�A�02t`�p�(�'�ܡЫ��D��\T`��?<$��2BǕ�rDo��n���G&��k͌�v��3��g�2�P�a���t%;�U�$�\;�N}����\��2�	&�K�'���y׻UltL�/��4����l8�3�Q\�^7�k� C��<V�Q@�c �1BV�!���g��.�y�'���8��,T;�=����ؑ��z\�O�z�EP�����y��
Ԫ2�P�>6�&'/"@,�����^/�;�R����O�(\��\L9l�4yoT�HGz��n�5S[\8S�E���c!OFr�!h��B����I+�ƛg����m���$V�����NV,�];g��܆���&[��a��#\)i����蕶 ���G<�,X[��ލ�L�A����7�����sA�=�u���B��g��³�+%��y��x����} ���C��=&UĞ��gF�x���֒�o�y�G��ѸеPU#�	��@m! X�>υC�Ț�� $�g��2���++y������v����u��-Z���&?�����[����T��n��ā
�H��@��I�~{s�l���5Kk���sn�=q�� @$ .
��'B�/,��ḀۖΌTaH��ɐ��0��,J�!ߓ�K!%"��!3��*�E��\������{-\�����e�X`d��]���3�[l	��7\FIv~DEyk�=���^�Ê�\�����k�S��c��t�x���gB3����#'�d�Y�_�rQ��ƹ�Q4�Zz��Xkd��͌2�q�\����5�9�n�!��\iK=aS��g�1>2���xjcO#�k�p5�YB����\#�Z��[�;G���xNy"��[uK�����q���r3'���=�3��3?P��ׯ_�9H-ʰT�ý�pB��(W#yB�ƪ��J�\:&KڎS>xQ��d�������,����DfRqf��ă�Y�a9�e�2�j �����V0"�������[4��n[<0��w�-�����d��x��]�1&��d����>%�=u�Ozd���N�ʫ��}��f�|v��rwm1t�ܙ�Pgy��A5��F�0?=�*�;T����j���y���2���1-T���Ƶ�	WubM����b�=��LW��\uE��꠯/i����꽦��������Dd�P�?�E[�J� ��q��s�n��
�,.aJ�	�|�I�F+�]c2��G<yt�f�Ɛ�^�R^se�6)r��||ԤY��.�l�lC�7����s�`�e`��Xu�;XQ�˙,��:R�Ԟ�]����E�89�WRT��n�ph�PkO�y{/�͜65h��� ����u�g�� hg�[����A����$�|�����p�@Y�UF�-Q�1��G̭�ɳ�Fxq���Ͽ�@� �3�Ж�*X�e� ��k�8�x���xj�d�{�(��G���>���r���cϑ���i=I�+И�a�v�oh�}XC4�.�ͽ��rq===�@���X�p���݅ϗ�
)_k�hk�������8,�{<Gzhry�s�B���R)�WSTy���C:�T9�J�'�:C� �� l��zq%{Q%ᬉj�'T�Z��9�����}=�&�Y�2B�N�*�����I����)nР�l�A�+
�~�|R�u���VS�Eơ_�u�L49���^u��k�C������&�{[�N��؞���8��ߵm��]�!*����7��ŒBC�c�B֩
�򝬴�e�)!wJq���RJQ�0�$wŠI�cyi�dcOγ���°:��h�;�+��@9Mʠ2�lT�]�±n/����P�ׯ�+�dʮ���=�):[-����2 wk��o�~�F�W#��@���{F��V�Vf�ܚ{�5�Cs�_(*�y���Ƣ�\�rT�r��b򬨴�����b�1k�?2
��Pv�k^<<uV�ʳα�~3X��2��K_�@�����_9����d���V�5 DAF��9e/�\v\$��4�[���*^�Y)a[��~��z_[ɚ��4a ѵ9����%9�^�3M+ڟ���WP�d�s�s.�y��&G5�NN�.��`Q���:��h��M��&�x��KA?���c �?�+U�~V��Ĺ�e�/k��6�26h�j�[�;���IF|� 91�eR&���;h(�ΐy�,�
WՅK��|�2�<k�s0Eq�Ւ���FhB�L�$ä�^P��R{��F�M-����Xx�N�L�|�Ӣ,���}��c�C�BԌXuX��f�Nj��7�nf|���]��_�����:���doڸo��ɾ��0p� ��9���8�pGWx�	��\��!j�k�	Nwl~|�p���������ρu��@s7g�j�V7MGN�h��,C�_��.�)�ډ��5}�������հVq�Ih�\J��� Ed`@��L �w
�b$PF�Z�n�l�m}�
����#)8ʲCX]��Ǥ�u��tU���"0�B�Z	S	AJ����%��� ��R<t��Z��J��W�^KE�g)�{:=�Z�'9ؕ�a�����A����Ըt/+;��a��G�.��C0�,nH��Ԥဳ������C��
�&���7����n	�[ݸ��޻ժ��l�#-+��)Y�Ȓ���s��B��P0���h���V
�:ͺ7��ϻa�nvC�|;�,���
đ��k"@8Ͼ�Ei��R)^��*����ʦ}B�) ��n���e^�:���^"`��*�N��n�,��-�/U�zJz��M������o�
�(I�O�9��M@v���E��0�x㍳.~�
���{��v�Y�[[~謀�+J��l�������E������~Ho޼I�>N���K�駟ҏ?����i���	WҺ�*�od|m��J�)Yr�l?q�aAha19U&���|9�H��+�hAc���	�ע�'�����B )�����l�/���$-�����n4N�u�k-�Z7_{�٣���޽px�߳E}�b���9:TP��C��������`
7���?�l $�x�K7�AyH/�@,ᯨ�v$'�>�S��v�����κ-�ѵ���ĉ�G��[���q�V�J�6B���>޹���e��S�ⷷx0�	�aZP�����n�u��ӖVIC>߯����6�h��`Y��|,\!#��;?<eC�%��4(a��p!����j��e���L�c'Ogv��ˬq��)��8��X��&?���S0�6iQ<��)K}��.��J,�!�Y3o0�Bm�w-�<cnxq�w�ͅ
�2�Œ��b÷^����vg*ر~.��]��1��<��bm~\k"P;�掄�����z�ioA�mQ�A]7(��l'��Q�����-\��ke�E������۾�>���9�ӥÖ*fp�7�%�\p!
S�oB2Vj[̻-)�}�@��0�mza�%'�O�%�!`�PG���+%J s��>�������~a� �nL<`���ͭ�d���Mgd-���,=K�����	����k���bR P���ϖ��G�;��ڪ@�4�̺E{횃��a�]��ә,|S�0� �G�+X��lLIo���eJ�d�q]C�'��bU夜+�m�\J�Y�������V+i}������ح�����d�/�)�	ed��y�籺e��Jo��[xƖ2��ӓ�c� �׌�6�1vχ���3����A�O4=��$��%��t<s��竧ל��@F�&�\G�Ň���~���x-?y*k�
���84Le;����e�u=�������)��/a~����������L���_O
5&gQ�6����m���:��n�ɷ�9�~�}|� Қ�l?g�ɻ��[HHn����cz;m����?���I�����k��em����-���+�N���o�a9��MUn��"���vqy����=O$�!4�?���v��"���Χ����T}����_�:xȻ�o���n�Wk�)*^B��^Sm_빇3!��~@��:�k~]��2^���m��?�AJ,Ck�]�5=���?�����?.������������7�Ԇ3C��t��聾��T�C�N�̚yv޽�μ"��̿'���͍�cz���
d�3ˬ��-�<��~&���Q��9���p$��O3y���o�|5i?�~�L�vz�7���ƚ�N���/T��!H:��Z$�,L�.�d('�,��-�%��s ��Ae���W2�I�br#��!�L�$1V����1�61�\����D��Zi����&ՀH!���BAwA��kr�(����q �`A=h�5|���俧�2�ч{m	�����y9���W['XF��R�-lM��]��[��I��a(.��Ւ8~F������/KU ����	�!���G��b.�a�_�^"òD-��.��Ґ��I��ɖ�t��)�m�ǭ���3���}y̆��A�xm_s-x�����ʾ���*��U��F���6^��'NZѲI"xu�0�uv��:rR~�]ly���J�
��=�@�;߼?	z��,��ǎT*���+li��~�+$<���
�v�k��T5_��G��E���	S&g�~���`�[��lF��ĭ5������������\�r� �-U���-��~*���W���MOߧ�QrK�[7�e �(}��s�>����|����J�,>����*V��9%(bU���"h	U����o&^6��\T�d9L�t뼰'��@�^�����Y�i<Ъ��C]�֞t��x�V�������pmlrm'�v���J�ɴ�,�9Te�}����n�=P�/M���sLn���>�����o����!	����G�>������UJ&Ϡ�+�m�jU�w%������,,�e�Z��7cPBj�&G��Ȼ����� h�(X(�#qB��9���΍�/wG��g+ZP��<��=��Ҿ�۠�E�I���J��?a�3�ց@�7�߰��~�A�ojp���*�ˍ=�'��K�<Vo�L���W4�'1����_aCv��z��؉G�L���˵}����-a:�8��{.m������;x�+9/�3����5���MsN�^�ղ҆g���v���� ��L.8����nơ�i����rX\0����APDs�K�`��L��>�Ut����@�H���A:-]�5qf{��M�a?�` ��'��W����h�	@�Q-��.�	����a)�1��aP�P��W6�^PkJ�vd���,/W�q�}��2Q ʹ�qh�B��D����iN��)Emu���Ⱦ Y�s�"5
��I�R�	ױ�j?����0���Z�{$c��?�:T�,6[-*�ߴ��^���#'Z'����8]Ζ�;|0�����k�뒽��V�'�WX�YQ�k��#�Y(:z!}��yiszr~Y���>�ݙ9�d��mMr�=��}���op���M�P�S��~ ��b"R�'Q0 �RZ<�ȚOB��r❷H�Eʵ�hiq9��yY�6�a�}�rH�A ��\c�6w����kk�G��S\x�jy]:e^ps�]�������>���:�չ�/�ԝ���=@���%�5:������>�Ӿ�a�"��>ll.�5M6j޷�V�s�iX+�8�(g	��;�.k�< �b������r ���@�;mk>����E��ְ�3J��:�E����q�0ؘ3��1�����#ې�`l4���;}�n#��s��ϣ��'i�{떼���9�^���;��>�Hm^
y�H!W�gZ���=���G�������֍�v���H8��s`RXÐ�ˁó��0���
��#@�^n��(��hP�}s�~�����2QF�7�B>(Y�ƿSi��~0�v^H/�iq>��~���}���-P������!�Z��)l�QI��%�1�9�U��U���o9<������Z �1��ޚ���z·w�*��7�#��a�\
E�z*:U�(]J�=h6�e�H�k�v�g�� ꦗ-�C���.��o=����T29�q��g��ș<�D���r�,�n�=s-��Ξ�7R�9iJ�W/�5��y���$�_#UX�6+�q�nᒛ��gE^T�%�v�w��X�g��u��@�rOĚW!^[��9��UXx�e=������n����!�-N�C�.���?�%��܀Mv��ٓ�[��2�tZ.�I��Yؽ�.��@�;�����S���9���I� ��ׅ�����C����z0�77�%�cJ����� elY�B:N4���!]mUo�,ON��}�ۃ7�����a��^X�wT����%���s���R糲�õ��[�Z��0�� �h������/� ���[�\@��l�C�v��{X8�r�x��_m_��7��9ߞ/���?����;f�g��1A�OpT�f�/���!�h~||�\pE�'V$(4�r!��#��${�\�e�Z��f>����LcȢf���٪}P�p�9�p�c>O��e<.�f�V���`�8縫�w l�z���;��y�ʻ=�Q�U�@�&W�rX�b��w�#���![���d�k���R�q����]J���S�ͽ[ѿ��5?V�>(앖�"ͽ�#%�����r^���4�s��?/
�8����	��3�נ%�!���SʗFN�P�(Bܵ������~�ш�?N��Wd���p���p_�id�7�3�?_^r�F�lx��/�~=�z2^���	y>�8��I�����^�qT=���� �z�� �_~��׈� ����+��֋\�-]�=�-9�9?���{kj2��:T����B#��ik_�iJ���c3u��/g�e�=><�+�26���zC�j�-�@6� )�lzJ��w��k���xl�8���~*���_	ޔ9�`������y
�Ԯ���t�.�xؠ����Lt&��=�O��(�):`�M����������a�`�1m�'�u��$$gwL���d�*`v�pV�|,q�EK0�%Z�p����=�K�A�5~�W�}!k���X��܊�;|d2 މ������zL��~�o������V��`,���B���}�h���/sAk^t�\��F���b|6��=c�X�ᚵٓ7O�,�<���9ZD�S��<<����,��gM�F��O���R=S���SVz��8
�Wr��3��%n[����{=<Q|,�dON��f� ��0wZm=v�;�|���aX�a�S*����I�!lQ�X*9Z���Ғ��N��`�Y]��Z�*�W-��w<@�p�p�>Z�p��J-g��% yHJ�<%�{���}�ۨ�oU{��b�8)�����g�d=�L�����5~����n���s����z�����3�-p�ZMwp��h�a��*���=��)=y2���NR��H���ByMi��7�bic�'έF�_�VڋV��gw�D��#qlV}�:=E!�@%vU���C���y
h���oj���@��e�_�L�?"_wPn�"��,�����H�"�K�,��]��>�Z1 /�G��?|���ǧϟt}IQ��=t��'�ܻ[l�.�*��j9��A���5�J3��3�*���e5�p��o���E��2GP��p�G��j�Z�����P��Ҩ�Cs~��s��Վ9��WS��u�]�AA�ǚg��hN7�:�W�C>u�%�!�SF��e/��\)B?@�q�|Lr?ً����#��y��L�wm��X��Th��%�4W����Y���9�p�{*��&g��H-��Р)���I�j t��vq�[eI
N�����5�PD����y�}��ɔC�kY���VF��d�(��z��9��:,��1ܹ;�C�}�E@+�������Q�!�lM����V�`�	ءP,��>�]xZD�#�j"S��*fQۥ�/��J����E	�3�L�}k C�U�s����w��xF<\���Qd�̆�-�3v��ɍ7��Y�P�P�Y���/�A�
��B���|knM�T���x�#yu8�Uf�L�4>Ǭ8����զ�IyP &��8������w��qB�Ϗ�Z����G���;`���Ƽ����d�]Q] r��Һ<����8�p^V���$(����B�>���4ݢ��C�a���P��Z7e�uS>��'A��ַ�vk���aN�~��.#�n��on��{�¦�WUnT9�Z낢3��7������s�r����2>t={�l��}c� ��d�����c+SU��G��U�wQh�C�%�SpB��v�)�
_��M"�rm1��q��۾�R(�E�����aYc����������`��B_��eE����f���_<�)(�E�a�[��; ��M���;�P.��ak�֩�;��^����q��"��f*�*3�V�l�o� �!��$�Ô FR��;VȊ9��WL:M��L�	�j�y���
a�iM���j�/4#m�V����m^��y�P���D����!�]�'��~{���4�MJ����>W���m2|?a\[�w��{�~"�jkB�c���sx�R�6,	������CRˈ���W34c�P�����
�ӹ�����PƷ�`z=`<�PA�M���	�	�g�	`��>|U9$+?Y�%���$^,Y�T��_���_"��J���}����Ih�>���N8R�R�t�^����� K_� ���$�5{5�`�«���!�:��	��ժ�����%55V×��?�m� �;uK_�J����l&��h��,B� �`8���P%�����I 7������ȹc4����R������s�.J��8�(l�Ȭ�i�c��?��wf��2|s�%-	����=vH�p�� !�^AFS睿���q�_��H�<�c�3a䖪�N�m<��
�pbd�i��?���a]%/��+��S�-����.ia*c�� ��uDF����)�?��'�:�Xe=&��� ���5�ZR�n'�O�%���c���ͱ��I�b�(<����&ߕ�a��Ȏ �`�
�U�J)X^�k�M�'e�i�R1��.ar_�y٦�[4"�[���Ɵ�T��P6��F�9#����}K "�������ɾ�3檬펝w������4:���a,��P�>WIЫQ�Ǭl��d��c�"M�H�^�(~e��G���7��!�ԃ����#@�띂��t�t�=/��?��\��Pz����BJ��Cs�J�L L��8��Rl����'�8v�`�����Iy,�^�BJ��ңI��|=tΕ׹� �c�0�&,	B�+���ᴄ�����	
$�91��*n\@�;n�0[ܱ#�s����neM�;��Ov�$Լ�ui橌�l�f��m�&y!
:)�ґ'8ԭUB��5����R|������Lɦ5��XY��͟�3�6B.#^���Q�O�P��q�Ҟ�����ZV3c� ��� ]1��\x��V0�s��9q�Sg��0+�KǨ9`�1b�ԁ1���CʡX�N���Xv��b4�u���(󘛑�TS�k���&q2H�Zq����
z�6ֿ�L�>�(饬4���Z��4��0L�K~�����lp�_��kK'���s�����b����1,[Y���U�ǽ6:�s��&_�{��C�*���F��y�Uè�����!�x�ؙ��q�~�ϖz��]�qK�8u���\h�d�՘��O��1�g�[Ms59w�Ye�6��cꞢ��΁G1�>��r<r���}�t���(��$7���Ց�C����
ܸ������ /刍~�o���\\>�~<��mԣ��\���;do����G��	0f:a�0���l�YG�;uvɒs~��zv�'�l|�>鯺^4���ޗn4w�N���6,����������J��p�H�ȝȀ�84ޣ�P���A�筄�ɘ�����-h?l;��e�eZ#[�i>��p�8����]ʜ�czٯ1RM�3����c_y:x';֤慎~��ќ���c�����#��o9�\*�����q��tU��#�,�צ�����l6�M$�ȼ�` �z�*g�h±�Q����Ӣ��0C/�5�����6�j���<��W�M���?t�2b]/I:2��}�\m�d��������k����8�<�]��<t��  �'Mi�zԽYY��M�*BY.���ؘ˘���� riVe���.��}�o�ʆd-؏�+�*�� ��}(�6�mbr0�$����`����ջ���!���F^͑u�S��l�˳�V���Q�����x`e����\�lLݞ�(?��顏�㋣G��5NZ#�W�W$��4%FBgD���8���mhna�=W���eG�p2Ꭳ���8�2�tH��Q���vJ��b���u�kH��*ٸ�m�+e��Gx���7�*�?�=ɷ5�p�J�`%�e�O3+�b�����T��_Agb�U��K�V��2O��Y��d	���l���Ǚ�9�{c
��:msݕ ?j�=�R%^���/��I��۷��uڭ�4�G����� T� ���$�"��~ϕ�*��A�>ݢ�we��Ty?�b#�vZRB�~�s��Fcxe|�q\\Am0x~�dY7��gN���(�!���v�u(��w��'�k:�k0F~�ȩ����"
w�[vb�qE�ܱxE<2���éǹcې$��A�8t�k$C��7u$�9B�n���g��ǿZv�=�z2HZ+��/>\v��r�/2���Y},X���v���^���:B���9�xQ�g�iV-��"�U�gu!q/r�Y^�]<���+��E���|�2b-p���~f�	u,T���T��I�w��NĹT�O��$���f2 �9�.�#"gl���8�HF�F���N��^.�j����ҡ�@ȕ4�#�r۸��>,E<&~uˁe;/����s��1�$����(-�����>j���/1#w���8v�P������Ca���(�#Y7��Л6��҇د������U�S�N'\!�:�S�	~��^��9OM�� ���*��c�	<ձÞ�>�]o�+M��>��a@�k�ɶ1���T;�7(Z����ҼY�'��~3ݰ���=��&	s�,����PZ�w܀�@�خrU8ﲣ���`2t���u���C��D���3�w����T&�>�V�ɝ�b���_k~����u=a3�F�1
d@3�^�{5��/1e%���y���!�����Պ;u.�9�'���۝Vj�R�X�xR8j�r�d<�HC� Ɋ|��v����+�g=��<��r]Y�tr��o���8cY���Zf!nN��xb���<��>gfД?���q(`%
UC�e�A��nv�lk�#��|�Ƿ��5�H��K�'"G��E}u4Q�H�?����.��2,� x�Ա��`��
�\EF`�F)c�k9z��(f�f�)U���b�D7D����5�X4';vT]���rWB*ɫ��K��a�jzU�y�6�w��v@^�<��>�*=P�P�����.���c��GN��=���������:~���������V����������4��_6����Jv���3q�5ى�̱sU���a�4�bUcj�1ȅ��s�k�؁#�����_��:���^q�\��hD�~s��Z%�c�`�8�	m���4<1Ϊ�:�$e����Yڼ@֢���挟hDT��[�:;�7ar�����<���:,��vw=fVL���y���ȷs�Ӥ�������� �Y��dB�����W��y�>��E������zJ5\��PGT�Br�/h��ݟc+��p�����[���*N�!��2��b��+��@�uu�Ԗt����ͫ6Q浑�J��8�I�uX^'��:t��>;?����f�p���h
�/���1�}�!���0�V���`Aq��(���jI�Ti~����bt-D%!e���"�2Ɯ�&(yA�y��Q�S�˜,�V	�Q7"|���r���^0����g��������V��f�g��f�R��	Tl��j-
���)j��A�-#!Q��Px��	�C�A����c,G������f��#!�>3�1N�D�ŷ�Da^��PZٛ;h�N�r�#�%f�C�`�{���`����"xU^}���l��ӄW�V���$��Ϯ�{�|��(��8��t��ϊ9�l��&��%Ae+)]��:oΑP����?��?Z�c�/��9|^����*;���\����LV`��\m�lY��1r�c_�Xm��O���u5�nl��!cw����%8K��X?����H~$��C0^�D��+śk��O����Oʔ^+&�0'|[����<$��a In
��mٖ�IsX�Z�9���˪�Ͳ`�i�>���dީ��+��=l7X�\��׮���V�g}���>����-�-�R��]�F�s~דD����x��؂��@8����N����1�����_��r�B�����S5�j8�$��S�j����/dg"t����cg�G�##�mr��^����t�.WF��v�6j���;;�Z�~������
#���^b��ٕ��\�ϼ��/�Q����_%���}maC���/(/��v���<}�5�|oc�|k�z3}�I����4�#{4�߇�P����I�������+��3�p8��Zw>���}�z��1B����i%;v^����:�[��w�М;5���f�>N���$e8��u�;��;�\���_�Y뵹�� y�JI9s'ǎ���A��X=�Y������\1bW�������k��n �2���aݟ	������)��=RO�i:p#�� �6+ʭ��L]���&���#(�r��*o��?��3���laY�Ws��x�,[���3�Z���|+��.]�H)�O޲�r�M\]���̺�~���,�2h��ĸ��;"�q<,>�FS&�}E���ӷ� ��V.:Ͼ���r�\��
J�=�ifE��;����-�r�"u�.��0�{���p�Y��M?���ؼݒ��T9e%rݦ|�R.���B7��|���*��-E��20�.���.x���ȹq��Z����=g�6eNx��'+qw�Бχ�yq���W^���N�Ͱ!��M��nHwC�IF�Z/�W�!tY���9r	����z9n�Cp�N�HB.�6���au��4vؖ�"�C6�E7>z�H ?Oa2��N���(1^#�C�����)Y�i2�(c��y���r ��Z�c��(�Ǎ�Si}�c�ַ<��|�9|u�o�G��yT͞J���sD=����ן�Q���q0�-8s�O����t�mW[RV݌X���F6�wee��d�֥ {*x1�'ˌ��QW�Uy�s�
���ziN��ʦJY`���W����f�Þ�xC�]8��qZ+�e���yӷ�-v��r����<�虣1v�Ek�<"���U���n�7a����0�Vd��sԍ��>�@l�?·[��>�ؖ����%�I��<�sE��\[G��ݹ#��:_��cX�q�p�>�vpQ��XG�C�ُ��׊u�oX.ƥ�7�:4���Νі�0���8x�P�V.�T�u��)�}];���	�Ϭ|�A$;�s�"W��s�����6���=X`��Y��{�j2���&3�L�WDu�Z�|d��a���bE�UA��2MZ|�����8ʩG����H�t�@8�Q�5�O�B� ���P��9�D��R�甹�ci2nUXN�mv��h
vB�chE�J��� d��m
2��^ۆ��g�}6se��I��s(g���X%����1������
��q�S�uU� .�ɪ���{.M�����z?����hv.��f ������o���$��7/�:��O����B=�S޿fv���3M_1X�nez��WN��3��#-;͠�t<��]�0eN�dˆ��#��#.��L9���z�v��[�ۿ�-�����x�P$�0ػ���H=I}b�%:o�6��h����]��У�2������؇�?� ��cs���٢�pC�tG��w_��I�E�.(�c��Q��oVk
�V&��P�DA�*�pld[����m������[�>xY�8=OV�T~����cV�1�毿~Xd�h΀'�����uz�N�"s>��o��*�1�즅�&OH�9f�Z�xMu���0F���+����X���d�ŷ�~_Ct��ޫ�6�y�H��T�69D��K�fί�Ga�L�̉�I�۸��-"B��������䃩��#�2c,#�:�,��`d�a��}rA�V�Äȳ�~�>�J�-�($?�Q�
8v���hł�8]��4��ￏd��_��ҏ�~��].H?�f<����84rK�T�F��/������k_u�7C�ĕ���B�fg��]<�2�;�c{�>��`�������]>��4"���*�vW}���|e,��,�h�a�r,�~���Ƙ����^�h�_���'��cKq�����a��]�VNK���c(�[�$�5�C!��}���1�ά�!�#}^<j�����o#Ax������sз�OoAN�Zo;����	1�Jr����a���?2o��*�/p	�|�Ȑ��6��'@~?��}'#��E�/9�Vs�_�i�v7���5r�8�Ʃ��O�h��|���uz���?���㯑���N�?>���}7�[�����i8����e5?8/^�{�[	6�.��d�Kn�Q|�CЉm_	�vPԡ�@wQ�m�#C�f�-�=rқ����܇q6����`Y��푝�W%�K��90�Zp4�#�ߒ=8���q���!?x���ef!��w�pW���ȩà:���|@
�YDG=`{�]����ľ�l~�Iyt��`�%*BM��Gϳ�1�#%��uo�V��e�~ܬ�W0�F����٪�0��ƈ�9��� �J�.yz�	
+�e�h�vQ-Pх	:[E��F�ڞDVn���J$;B|Gy>)R�Z�c��j��%�����?�M����!|Gd��瞭���n}"(�k��Uɑ;���P�EX�ҍ��M���K�1rC"AÉ$��';��3�,�mu�3�㈊�B�\)�WNv�}���b��yG2^�0C�硆q��'U�H�.��u��c?V�~��v/;*�0��j�+�����v8���g�Ź�bV$*G�#/r�}?!	QǞ�A���2�?UN�`�S̀t��	ר�~��ysTc����?��
�G���D��B~�2�����}К�vK./��pv�i��bߍq����w��s���ٕ����޿�G8��~z8v��Qn]�l�pļ��{��58?�k��Ph�n�~�J'8�cl�U���fΜR��)��1�Z�}�C���3���A��@�_#�k�-:�0�Bj��7n�}�*;^)�Ym�?�Z�+�����^�9w d��`��gt���ٙn��:m�Umu:��|X;X�f�;�Ǽi��`�5ukc�Aw�|������o?�$��cq{��GK�'��o�?��o�h߇��6����gc��a�! ���hv��E��4_�gN�W��]q����U��S���S:�9��������$�r[ ���&����U$�l�,�%�Co���[�ˇ����
>�4�	'V-��hj`����:�ʬ��6G.��s΃�/�:M�����VNp�D��m�|��@t@ᷪ��\$�_�c`<k}q������L���l��\�'E��_iyIĉ�m��᎝;����#�q�O�-�`Ѕ� �{dbw���k8t����w�4�^��?��-�H�����w$�=K���^����%�#"�P���WH_�!n�j&O��N�E���z�1��sYrddK�Y��YH�A!��'z4��|RХ��lNDBɎ����gBwڼ��<J_���p�y��Tp*�r��H-DkuҸ�Ar"w%d�-a�>�8Ɯ�~��!�S��f����K_���z�e��0�ЗAx���#�>d�{G��!���ߞ4�iUd�Y�� �3����Bt<�SB�&"M�R�%:��1 WƚC��V�&���k>��R�����1v)Lk<)(6�zXߧҊg�ߵ͓��$U�I0}~7�%G��9�����!�mUT�a��?����'�a�}{|S�;m
���7���
y�����$|?0'���U��������gCVN���=�+�u�m1�~2���s�lUV}̰]�,��	֍���f�ùs�T�d�#�����m�W�'H�j1~��`OB�9v�NrQ̻����Ξ�XhFz�Q�!�-�n�Vb��9�J w2t5o5}����~S�,�o��;���JG#`�۷�@:lE�Y����$5q�*�����?l�ږ6d��ۇQ{>�?��*)����n�w�l�y+H9�g��Qyc��@'ʑH��;�y1�*����i�ӳ���۝9�F2�������$�qr���o���le��]W
A�j�g�9����ƱS��D/�������N�d^�Xw�]� ���Mq�6E��y#0.b��h���}b��ҏ��|7�:-�}����]�<��sV`ލ���Y~�������#!=nD{}��[�l�S^�����b��g&�����fG��A�S7J��)_����'��`���1���*����˾z���۸il�F�ݒюC)���M8[��y[��> ��WV8��'�S��k���2`z`<�Vx��=C>дf�,��j�gDV�����0�M�Fw��4�[�8�͊f��#���������zYG�F[d�8�hU�#鴈Lѣ4���J6����)դ{zd<�l��e1�;l�(s�S���uc���C��p�.w�u��?�����Կ(��q��g���Xp��t�:����֯R9hn3����ق��I���HD�6X�_���5	'���j]Ǖ���~z�����Z�Üy��\/�3�+w?EڦyƜ1`N������>.���������������/:</U�
�Z�ϙx��Ȁ��}��G%����{;�����l�5~aC�!�cR{͠�\x��1)��	8���a��1ӽ�U�y[��Yq�_����d�P�q���̹��8�n&�Q��g��)�糡�Y{��Z���������D�i��� ���D�8Ƶω��+Oy�+�f�m��3L'+�4^��g�*s��ˎ%v�p��c���0AU�̨����HY�7�sS0�������>[�|��'�6��̫�����ԇ#�8��#fr%�#�Y8DJ#*��?���i	�����=��.�n�J�D[�p�����8�'U̈n�~4Ԋ����NQQp���u�Ч�ސ1����O�X�o��v��o��ߝ���'~4���M�y�S�r�i���R1ȉl���5�K������L#ְ@��bR��Jd�l��ʷ��6{��<��7	ǸA��U�^�ϑ8�0�N_�g��j�ĝ�ϣ�"�Ӯ��)�\O���N7��0�x^��ǎ��yφ���Yٶ|;�mAt�U�����U���D4�����^��CsC�6��#�VN�Fx8ɡ{#gG%8��ނ>�W��q�X�팋^^���s,��spU���<�V^DJ���D"I0�������騳5UL���lҧ�����Ї���pП�>�����c��}�f�8l����[ъ:�j���m��yn�&� C�u�QG�i����| ��c����IX��2[@y�2^��tۨ�c�Q6����(=��<��hu�/�'�G������RyxDCd`c.����ߣ�6�z��a1O����[�/��p�q;4�h�@��F�#w�����ǻ��IӷY�nWߝ����6K_��fl-{����ﺈ��2����͝���w�D	�uA�;�;�:��uV�/�H�?�F#k���;����8H��Kj�s�lS!>mtX�m �ǜ�d2��N�S�Wrx��掳R���Ă�
^j8��))a�����_=������Ag�.���R�A��8�����i���*�)�(���K������������à�V�@��c���L�)� s��OD[�]|p����2P~�>�оV:HA�E@�F}�`�9k?1����͊�G��=w��1V#�D\y�rq�m�P ��� T���hj��'D�S������O�����h�s��Y�G�4�\���9vd��t(3\�~ѱsu�U���̹��  �x��<���1���/��cl�9L�软 �3{�S�O�V��&Ҙ���+�my���v�����r>����S�8�"�W�Λ�6TE^)ѹ�Ǭ��w�|;M���\-*���B�'ƾF���
�?��K������3\�d��L�4X5�B����V�q4�7Q���x�lg�-�&�q�O�7�2V��wQ^�R��#�=9��6oW�'���;w�gHb��@;�TS��f�m~�$�oc[·Q�WK��w��<F�]�t��SDLX-���n�-K�q������M��~�G�;&�pd�*^x����y��M�QcK@=l|��R I�'��Utu�v\wcz�S���X؈�J�;`d�����a�k��	}���\��S��ˑ�;�!U�ۂ��8�:Ou��|�q�ؒ��E�o�8��ݙ�t�Y�+���p�b�d�i�KZta�T�;�({F$&�����V���y�3|�4�K<��F!t�-��G/#�o��������~ʣ-��t9R�;���	:�ِ���8���r;^%����a3�X�7۾�ӓ��Q�F��o�	�'gc����L���Qh�"+�o\w����s����}�!C�J1�����o㳷��:c3[rD�(�y�~U#�_���N�쎏z��,���޿yE�;�����D���#�o���~��y��x���G�N<��Q�-m!Gmk��y0A1�Ҩ,;dbo⒳n��t��r�w3����uTOq��\�r��7�یˌS�0�p�HU�8%|�nºØ�]>ު�~k�s��������nI*�˗�8kO���|�m��� q+V]}��`��:nJ)�����S�f��.�(������x+5�/�,��e���٩Rq�	)\˺�R)f���֬���.+^��R�����K��O�q6M��if�7�c�v��ҵ�F����k{� PV@�b��~T��;o���e����+�F�
);]i��J��o�x��`�����s��c���Z�F�(�;�+��W�a��ӣ�Z��"+"��-N�������U���`�ߟ(,�"8���9i�:C�C�μ0�mkC�$�<F�'4�K\)�E7d�d�u�d叟��bEX@OR���f�0ݔw4��c;�a���s1��Y-��7#Ti�a;p{��aF��7q.'4�U�x�UƱ<F��aޢ����:����֚n;r�^(O����;Iٱ�����i�*a�?�c�ɭ�%�+JW�>,���)Y�)Fh��#�FS��� ���7�;z﷛�R�1��g([�f���|�w0.{�	8�Ǽ�CS�.v����84|C�%�f.͝i��i�k�prMLC�o������B�����G>��O����1�99Ԙn� eGI���kI&V�X�����"���ڱ�2�w�3����ڠ�g����$���~��� ����(�'�N��Q����JrJ6Z�n������7� E�O���F�j��E|ض��s��ж;1N{}<����q�'m�\���W��0FTrQ��t ����D�����N�̆�}ȩP�$�sf>�N<��x�]���c����Ϛǎh(��ɣQ��4x��e=k��#C�3�&{$������p�������4w�*Ɠ�IzC�mŀ�Pث����+��g�Y���g��lݚfZ���yŨE�y��N<���a���m:��S�n�9�@jf�$ϼ58�J�i~�#w����1�� �a�u]���5pV��pHT���éS�'�قطw�w�{{y��e�Yѱ�16g����V�A^��L��߿��0�@t�����?��+��D�22ZQo1(e}�p�#T�a����E
Gs�g�  �֐A4��r:��~g��;�/b[���_�q= �B�TܺP�W+$�Aa����9>��'�v��8���5d�\|v�z!�g/ce��Q���Q/���G��4�����(����ޭ2��ϖ+&d
=�χD�ـj�zb��v!�S.�α�3�#҂�^QިJ\��v���6M�ui<2�od��rFC�Hn��?ʟ��4�	O���������'vG�ѭ�'H	J/�rLS�V�x�$�c��;m�r�_�*S5Oݑ�pg�n ��S4 �e��.�S���)�	)��}LA�Dzj��'�Q%�k�Y�3���IՎ�ǪeU��O�(i�L9-�g?��]5cܢ��^_��98�,:Uy�	�"�18�zG�!�J|(U�o��}(C#_�_]��KC�5?��f�(7X���%:@��\-h
7�.Y��@B�FrP�"��d���1�z'Z�1M|�����Z�-J,f�g�ܟ�h�QnnH�RBߜ���+��	o���Cs"!�<Hr����8���e$�z�L����:(x�;���d#h/l�+���߷펜bòX������H�K0z%ڟ�P��R�����Q]2�A���'��q�?��T}�C�?8��s�8�,4��8���Qó.�^���q	Vg��a84ѻb����S{�qA�PU�����!m�q��2��q��m��F$6a��xu��=;#/l �e�Ћ��]q�},j7hDO�%�o8��F0p��]��,�&
`&���z;�@DT�����y*<';��t��������d��������?&�׍ܺ��d��p���O�yΑQ;�~s�؎���bם����H��6�;7�+�.8	�ा��4�n�!n���gyh>,>Y�Iv���>��d���B!+D�B��L�K��p��t����X��]�&�����+���3�R�?T�w܊!X�k�FK����A���5d]g�P��L�%N
(��J
��k�<
����-�d�n�D�>m,�����&�����B�c���`�dS!3�񛘃Á�0a��7�p��1�Z���h�h��BW�sǡt��6z/���1��T��QQ�o9m�A���;����WϚP���ot관��|a���iҔ����R�#*`k�ʎ���q�m�|j��qZ�)B��w�ɽ��tG��vuRRS�,:�&jq'>V�,_����;�ގ%�"��m��w3�jq��!���;x��c��Ѩ��X����ls�ҝ
������l �7���!/��VE�l
$�6�@u�o�c����t��B��8)�%��S�4�yȻ�p
��xG��`�qS����9`	����eWl�VY.͢x�q�W�b�I^؂mʽ��m�x�:oG;�tD|C��1�u쬨UC�#���9@�퟉�;�Xb�շ!i���$��c��x�ybF0"K��s��>/�;1�8RTh��k�u�J2��C��ö�)3�z��@�m,)�h}�uX�/��.;�L�|?,�+�N�eVm���Y���i?���BV��Z�SK���I����*>I�ɉ��׊m��q���\g�Ӝ����ͷ�BΡ2�<�
�8�Q?;���z����m]^^Z$�z\�MH7�g]mfx�O��G���|OΫ �=��qR���z��`����c��g,sU�Ψ5��Q�G<�H^�?�Y�9�h��L:M�c���0l�a����5,��y�(F��k���Ȁ�Fp;������TTf	4�݄��35�tj�X�[a���/vز��Q����v��g�N.C'��bL�ᮎ���������Ǜ����PD���ƾ���_����Z�������\r1�H�͐[�K�E)5�ez������<� �lU�������GTZ�f�ᒃ?����(��a�K,�>�[�j���OSw�<���G$PT���6��M,�1$6��л@{C�w�t�d<I�'�q�Z��?۽T�w\U�����U�A�A<����r�ت,5V�T�_��q�Gp���v��c����Cѫ�V}<��
��U�����d7��1�_}��V'_�+�r�1䫼Ҁ���N�z~�%��)p�4>���,8o��i<�m��J��>7�i>&��R�o���`�F-�-���pR�#'�¬N �y��c���&����������Y��т�Yr��������8`B�R���-�X�b�a�a��6�]S� p�dse(���6� ��
�T��o
D�5	���o�b�(���Z1?�C�E��.a/Z������J�	��)ѐ*v�Ve}�폴�7q81�7M��1������OIҳ�x����q��M'N[���'N�g�_����o8����k�w��%�j!|{���JS��@�r�,�dt`2�u�B�;}̈��<#��gU���B�o��N�<����=W~Ǫ���k"�.^�����S*-b����]��tn,�P[!�8�?c�{��ϑ�����V{���=׆L��c�۝o�q:�}��c���1�B�*��^�F�0P�9��Qu�P�Xtػ������^���>��&[5M��V^u�x�Zla��,|��=�T����ƴ��rƌ�Q�D�W���xn&]��8��A\Ξwa�E����~��v����Ȍ7����贿&ə�d>S��Ӈd�)�\�@��滹�d�@��Kj��EQ<ލ��zg5\�M�9�y���|˷�p&���<^,+"�V|Ro��? ̈́>9ʌ��0f�2�����LJDo���+v���ܝi	�|=Ҧ�l���+Ǖ���i�����:.���l�pz��߮St]~�����c��)#ڵ��� t��J8���66�_�N;+�iEc@C��� ��O����|#\R�e��"LV�[ۓ�$a�s�fi�-�:;��pA�Ӏ֣#�-d�| |�&��]���}�l��0X-�^����h/�.��Tx���2�xf7��fz ����3{[�nV@��w�GY��AV��<���ڲ�U�6�6�1^���rB+�ǧ�9�CN�y�4����~��p�7*OJV�l5���\�<�d���ɖqX���p^f�-䡇���a���:��x%��xv�l�����h}���zӨ� x�w�A��Z'��Ǜ�9\���'̼���qPfĀt�Ǐ��;G�@	��ɸZ~�[i;1}�5F"D��i �V��d����^��`pY)߾_Mqs��ဓ��ٚ���$�)�����M���!��ևǸ��4c���+����#oNO/��[TDWw���c8lz�㹇`�䓞��]9M���{Ύ���c'��%%l�sR���#�;�}�R��0ŏ��QmΧW�_0�hl��|�:����if��|k�i��$�9��x�t=��+��(;E�wd݂�6��y�?�3)�f'\��u�C��4F�s�\i+�T�H��l@���B�}a5D�5^X��z�Dl��I1[�	�K��EM�e:J�Hci�&G�N�舽����3��;�-#���l֩�0[uRi&�6.DM��r�B���u�ڲ�0R�7������8��zňܤ�nN�RZs���j#�$�vO>����t�f9
e���M.������S�5H�zB�&�Gl[�:q�Lg,S˂��r>x��U�`��E:-�ݣO�g)�"���;�w<�n82�٢Lm3L��T�٦X5z��m��\O�[�Y�/]V��)�k���"����:���M�!N3A�����Ǝ]�'�#�T�`U�����|Y�@��Ġ�dO��f�����`��і�WP��!0(n��eg��<��~� � �s9V�<�%Bh@��`����0v�To$�D�������
Z#t� ֖*W�qA���	Ȍ�槫&n�8w�/�3���a�f I�F(k���Å11(���ŉ�O�f�9�:�O��*j��uQ��	�x�h3��a7e�	�u}Ü�J6��&<�~3]���T	-�����2�3��D�ٮ�X��03L�<Lx�uS�a��,M���N���ad��6x������`?h_�?.48(�=4���!L+V
�˕r��5]H�&�YS����ry������[2P.��i��\4Ňߋ
�J��_��반��kj������������!_�*o�����m6���I�y����Q��Dt�O�ִJ,)��Z)� �MI�ePǅ}��`\-�H� �s��/\��;Ю}�6�������Z�;�R9p�?f>@*.���gK8
�n��e�>�'����HƧa|z�{�͈��Q�����A�?�d���c8����ԗJҫ����KԿZ�Â�s�cs���K9��hKe�:����Fsp�$��U�;my豓�r�;7ލ���rt�mU��@��%��&�`s.��!O�%q�� ߚ��l;�K�������3���"�oX,�s�*��-�W.t4{�i�����Ӿ̝���I�T6�W�*3�On<���g��-�m����r�~�s퐺�b������d5�鳃�d��a����w�1N5>倔�͵~��_7:Ѯ?�L���??��I���P�]p�w2�����[��.Ӑ�����Z���p��
�{��0	�ˤUd�YQ���`�W�γ�`��S'=�-�=nvB�'q�g��'�O�13 0��DU\�&���S�KE��I��cޤ/u�y8���Z�ro��q��\���u&���;6�ق.���B�C��	����gZOI�h�%\���C]�O�h(^x���p�)JL��^�])��m�Gj�q�޹}��.�˩�{��+G�T(зv���]�nž텡�'��8/��Ό2�^�]�S�*���v��䂾����a	�e%.ֵ ���b��+f0Q��D�K>u��,_`�m�e�)�0��jX�mQv��W���6�RkYm�!�xn0����.��X/S��z���2�`�G
�C~�s��Y�Y3�����B�BR^��q�śim�*�?������{?p�>'��ø7O'�YT@-�4������h���P���~]���Wp�Uqs�녭�uz�F�l�s���7�sGM-��9ͫ�.�m㧘Ё�>y{[E���h���1э��6�gΣ��q�=�����-�~�h�I����S[d�;c	������=:��V
�5U��a�9���"��h�J�Ƒ���q�h�ջ��G�s��$��,�z]��]βS�j�m�#�p�P:6�މ�s��n��M�������S���l�^i>}���z�@C���"�RK����������ad��{�1#!��s�R$[i�*&ݨ���\���(�G��mW Lo�����֓�"��Vq�ک]����4|ʢI�+d�g�CI��L�t�ș׋��<b+]e$M~�r8tF����u�ձ���m���J};��:m��}qg��~_�׽V0,W�F'���&��Z��D3Zj��jGJ)�O9��ś��J/�FSϑs���	�%'B��
��)Q�`�pm7�nT8Ӭ$t=��nO����`�PJB��s�`+�)ӱ#�E��k�	�D�訦$2���b�d�[��׿�=vִ4�<���AHW�}�^�c��m�܂�I�^�����եϿ�-嶦�Ϡ�F	8�S_�J������q%�,��:|7C��������)��]����m���)aũ���[�v�F[�r&\����͙O�T�۠/�n��R}��'1�'HƸS1����C�Tjە}��/9�Le��������EY�4.��v5�uO�4�"� �<a����'h+U/�ĎG�<l�{b�_�=H���Y�Fؼ�6��qU���u�<�9�`48�c�q<��_���K4n��f���Om�����X%q�k$��2�l,�! �.p��=__(é3�t�r�s|������o�V(�(1�Σ������o�۳��� s��Ay��n�x��ۊ�?Q��|�;NZ#]�e&;�fG���m}5���.wp��a��z�#���yz1z^��4*���Ƽ��;z����~��v����o���;�a��<�`�ا��.j	��ao2�`�co��c4䣺Xl�uu�݋�K�J�I�^h ���
�,5m�jק��ƛ�SY�.w{�8x#>⎬2��S�������~�5M� >Yt�9Z�y7wJ�м}-���>�1p�#�z�_�EF�У|��[y���Su�79��_U�h�WUI3
W��b��p[�L�����Ď}��'���F��J�9�R��J�����s�Q��8AJ��n*Ѿ�����ɋy��I7�ܰm�:۱���j���I��47#>�������ǙS2>v�Mx,�%qN[���a^����3�>C����y-B����\f#�Y$N�zV��Id�������N.��j>Vo���L��܏���I�V�ϕNv��m�����!��k!�u�U)++*�ə�TI�é�bo��V6�b�P^qލJ#U�89�:]#Z�<
9AȑA|�K-dd����-(eX@�%|��#W2t#�{�F���+��\),��8;u�
��X&���O3\�R��uW���i���J��e��y�M~���{�N���E7�ظ���N_�EZ�)@��D�ՈQ�Z؊n���j-�.Q�gu�/��73���klb����ɒJ�-\^T���Pu7pPJ�	��)�`�-pC��c<��Fs���P�h��7�Z�-�L��	 �M�&�j<_���|�� ��<v4}�tg�KNyng�!�fky]�� lI�Ns↶�4#�D0�>�m�������U�|��}�#���vܖ�1���`
��	x����X��Vjz�O�Z��G�w����/�9�񾀡�?�*��5���杌��LS0L��:DΧ��=���1��C�M�1�{Ϧ�h1�� �4-��T�j�@?� 	�@����x_|���t�M;�P�=�ql߶SU�P>�z��q�T/=�O��~�p�ߗD�O��0��Xscv`^Ք������U�/�������H�
,��X6BքUu��?C�f�A��>9B�ӯ�c��EYث(�9���Ō3�O�db��ʩӦ����M}Xt$��V/^z�SE6��*�HOut�c��y��~r(�����zv*����a�Q
�ByQǫ}CF�p���O�
1UM[�r']Tϋ�������Жﯴ��Ai��\�8�����D�:�Y�6L����i�k�*J8�M�?��B���4�EWWG���=�QML�#>$�TeɎ?y���T�;�$0]�� ��q�1�cǢ,!W�ρɱ�J�m5��d���t��ǀ��Ǔҟ��e����f��V'bA?�jݿ��Ln�'Ŷ9\C��KUBM���ʫr����'�M;���w��[�zBΦ�Y,j��D,=�o��h.�# ��lp=�C�hǍq/�X�2G��h�D}	ėK��j��R���!7�-�����K:����fڎW��k�����I������q~R��m���,Gd{���3t�~��b��{I���nD:�8�)�7��#V�7#�ZX7a���E�����z�gt���Փu��<� ��)u���2���b�ʦ�n����%W�֧�g2�(�-h$gDo���=+�����I�0h��o;�]����o��ա�����v���a;58��G#��J��0~���6(�=2�ongT;b�n�Qv��M���t� ���5�1���|��7��7m�~���sKl�=�o�O�~ޜ��&����	�"�?##�YB�[�3z?<��q�H�^��VE8�ju������w����[�������`�&=+8�d�p��k[�p�w�T��C�#�ƻ����*��P��٠�,&	1�Z]��_{G�'��p��dh�I�ވ�k����y5ς�oǺ�����W
�&Wja؅�f����r��7���*3�Z<�1i�W>����w��΂SF�c�G�����t%Bv%�i�+G������.F<����׊AB�hf��4��ɟq�\:(�c�����vb	A��h�Nא�,5�7�n+�
���nn� $%u�����ʅ�F5��Ew���Y.T^���5�����<�g����/�x����.��T�|5�J�"��^՗Uvݐ���,�>-�״� gY�1�k�Kx!\W���6+Z��թ�t��}��i�s�o
\56a�D���k?�D��i=pZ�;���Ay�q�0q�JDP�Q��t�#��i=ٗ�nx)�<��N�,x`��ڕ�'�n&}'WФv*��ÊU�iޓ,�*O�v�A/�:�[�4��N3|P����x�eŎZ��:�|���h���Γ���Rk�{�	�Y���y��F�q���'����/��㉷3n�߇8�4�"���F�s?wՁ���R��5�����X�=���x�kƏJtd�X�$�n�3f3�J���CU�4�}ȩp� �})���Bǖu�^!���� ̭��YL�*�&"S���	n<=�y& ��"�9���ޅZ&g��t�N��S�-����q��`s��]�� ��.���줝�6:��9�h��o�?$�eD�z�.)2��;?�Sl?�S���M���=���.��q��'u�t���z��l %�w�{��e���
��+LԱ�ѣt=��_#Գ(я�R�;�lS"iL��-�fr�	�7�F�����"ٲ�-�X�K�K��O�ԙ�DB��O+T�b��|�7�o����iQ�^�	�ˆ�}��*P|ǊZ�v�	�0�[T̃!gm���.�&�/��H@���LNx�l�п1.}��z�����F:i��r���^�1��^���<�_�>�W/�;_�_H��`��Ld��S��|��"+�SFLu��p�Ċ�r�P�z�%)��h5�;+�N8$U��G��ۍ������<.��t�R��������EֿM�<�:�[' �gZ��~�	]���ݯ,���,�l��@f��j�>�R}ֶ8�1��%�s�cGɉ��l��NG� �[��6�J6�^}�^ϫs�<�����?�,���\��q���?t��:CHG�i4p�{k"�k�b�S����ӭ��W��HݔW�9��Bմ�=9����V���`�+�R�~�O�]����J�D��V[+���,��4- K�طۋ��1���:/�)�se�5}��o�O=��U�U�2s��1�}�88k�
x����ƽ�9�Ꮨ�P�'�y̼�q�d�@��*������- ]&�8�qf�_�K��-�Nn��]r$�IT�y*�(kx��O3F���~M�Z�-;���G�ݝ����Msg�8���3l�5Գ`f�β�d3^�h����2Ե�8��2��5�oRGuk=9�tJ�!�W��s��Jc�T!�Qnz4��_��q	��Q�R1-1_p�]��KC����8�f���W�t��tg��e(eA�vH.ݛF������r�0Gt����p�F��L��?7�������^�~E���?�x�F� ��q2E�/9V��������B�y��ȗ�rPQ&"�NJ��� ,�h|~��˞���i��# 8�1��5�x&2U�Qh�J�/�pYN"����t/	c�E��
����V0W��[��������k�ަѱ	�V8���,���$�͏#3��^Av�6�Uɠ7�?՜E�2s_��|Vx>Ӷ���'*�kL��<�̮�DT}JL劧�l�v�^3��d�}�����6N�H�=:�����$P��e.�	���L��aȚ�K�3�{֓wn׾���L	�m�g��[�9�1�y�����)Tƚ��5.�H��Akܞ&Ǐ���߉w����Z!h�����^�}{+��a�8[�D�}�͜�����
Zֹ�0�I�9pCMz^\�Z�P�ȉ�4C6O�g�_2�T)D1��X�Q�����Dk��A�_
zBK��c.�O��3�/<���c%:w�2ms,�n�0�g��$����U��>���)�u3��Ŗydk�nQ��|W"W�)>ʹI%K��j��l��}_+��}-�P�?ԁ%�z���a��?���0�{��;Ȃ�h�hT��ܒ���_/���qğ�z<�c�Vk�g��zZxV�ڪ_3���i�]��Pw�ǵX�.�3�#�\I�5�vK�D4�����ڵ��$ؽ*��I`�4/���I4��U��0��� ��!���Fg{mĽT�B�!�ȧ�%<q���v�H?��(rR�XD
��MN?$�fe*z�{��C��^�=��.�e��;�,���1��Ws�n���~>c�V�E[Zl>��4����'
�T�Ѐ��zl����u�<��K�Mj���@�Y)�lȧ�@���j�F�P��yZ���Q�r���@4�j�:o��9���X�v��Vl��������,w���\�W���u�9�R&���o4�yE`���1�ꠋ²l����OG�A0�*j�sW����]�DI�ȸ���F�X�S�b_hj|q��P��9/�_G��ɋ� z�颴̎6���,Ŕ�����fge�,pG�yn��N+Q��ʓ��ʘr�����n�j�����<�쬹a}L �G�qv�4���F<��
�31"�x�d���� ���WeJ�<+緳��������*m����ۈ��>z4l����ₜ���ʟm&n5��3F[dq^�g�/���ȥ�^�j�?���zjSG+��<0݅��>*�50[Q���A$�_�ߗ}2uGg}��rK:�T�q�k�q"�8�5%#Y1��Bۮ����Ԭ;N+�Y��񞌖'}�|�ۂ��LV�y��Ԁ���՟�����I��P����.f��x��|K��9gN��Ӆ$��M�q��l�(�����z�1�v@��"����D��ye���ķ�}�T��r�P6-�Gǚۓ�8X��jT�a�(�; _(�#�0�l]�,ƕK��./�G3�/8Μ�j���9�����O���������?�z�	�c��	{�k�p�"���������U�9��;U��Ӈ'C�T"�q�N��ΎF��,�؋���\Mv ���(.�˶�'�΂��80���OW���P3Jh���{#�gǎ�?��W�+�XQ�Z�T#a޴�^W�d�4�	U�%�Y9Q�+1�6�fu��6Z�7�)���GE�0İ_xr�U�?�"���L�B�	j���ҝ����Gz?U����mb�ڜ<�������$lk秧U��u{���E�k}36_��BN��1^{�#�|(D�U�5-Ĺ�8�Qyx���KpP�-���3Ա���+Nm�g�y�යvD���i�;#����_k�%���'���sౙO����S(C��h��%�fp]��ϛq���o���w�S.d��|�������#�߻�k
�'=ݠ=W$���g^�J�Fm�G��R�>#��v��z5�\��f�=�yf�.����8��a>O�O��ʂ�y[3C���?��+ ��M�߾���'RmZ�_�����p���][��1��˺�k]k��Z�-F�:!Aئ+�u^t�V���)�ŀ�&.;¨W8��'�;6�7�wo��c����T!� "o�_zZ�ū�N�ׅ�ΚDS��N��XmpT�XyY�mu����{�#��h��	��j����d��L�Xyr����K��ճ$wV2�Ɔm����M��`�y첳��O� s�Qk�6������N�v�g��H�ʩ�L����ۤ���*�ŕ6����	J�؉3��%�p�&���>1�n��LĲ�*��d��'DP��&9�z?{�&5Qc�n]��1����RU��J[qbΟ6�F,
���P5�6�5��V��X�"�����U��4�0���*^��*U/&��.xҙ�;Y��ʍ�{D�ض0�yzL�sSo�~�KI������)�Wۚ~}�1�h�mݫ�!?H�~�+����/Ŕ�d��)3���J+a%�D�Y��<.ܮƕ�;��������R��2���_3P��~z7+s���מC�뽼y6O��#D����ϲ���^��m�\��*�y�*|$4��7��6�o߿�?�l�x�X_��%��A��Z^[=t��W�V2mE3:BC� WQ��Q�4�eϒ�W]��v+��2�^�e���s�r���u��{|�s��~��r�t}�-~����K��e>μ:Dq�e�T�:����F���=(��s'-���C�J[�Ra����N͟1x��Qyb+E�;9*�b�|a���I�튂M�N�2'��n>Q��䮬k:kf���U2�t�i� �ٟ\�B�_��lx�гI�f��]�L�)eG+�^��-�O%G��n��u�e��#`��!y��D�-��E��j|���O���ǲ\��7qh���z~2��j�O;�����WBO�p��o� �����u�w��A&��\���8�����
d�*�aly@+�e�4�$ت3��%����DSY��><��^]~��J�M��\��n�'j��x.��o���,���b4FV�E�Q30&�e��LuR��VJZZ1O�c�DH����Ͱ���\�~%^+��`��;�)�K����77�j��f�@iS�i\t�� ���GsJ�u�eh���XN\��4�2YiOͯ����fE'>�@��rLt�*b'��k\���W���)�	�F��lv�Gb~�ڕ&I��>as���t7��S���	��cٱs I&�S�Ü,H���Q�)3���̜ezgDc��4Ǟh����yRDoP��y٦^���:;�>�0˜� ��|�g^���Gt��`��l�/�_��O�?+�u�Ʀ�(�w/�
�~��S>gh	�q0M>�JTٺ"��x���:]��,2���k��g{I�ϪY}��x�Rf��ˉ��̩�3�7��R�@�ʖv,�������:js5C�U�#ҡV��C�V�=;�a`s}�SB ���}ΰ��7�'r�uLX0�3�޼(^;a��;H@k8��Z���f�y�Ժ����j6R�'tT��ŭ�]���#�X"�m��Q��{��C.룣����X��j\����@G7U9EV�PV�IZF�I�N[�>�O��<��i���+>�\p�ƀ�M�6���>�h��z�V?{D�R	.\(��u�Xa�}�xp���ٸ�k�o?������b?�V<[� `��8����2�0����I,g?1� ����5���Ah����h��Bf��B_��
�'�Ϊ+´]\
��[ʥ��ʀY5���V�~a	�����0�O_I ��k�%:%�h������Fh����n������gD6�#��~�LZ��V.��a���{dbΈ_��
H�t��}��h��hզ��P$m�+:� �p�Ԯx��6Y�[ͳ��T~g�;vW�z�=�������5�ev���_���j��<ߎU���G��Wq��F��I��ߥ�d�=+�/� V����~F�{��^*��%��K����"a���)��vP��k�����	�s3Qt<N*�Z8�hs�Ӥ��W���_Y�����l?G1́Q.��#!�O�OS#z�Lk��^��{`�V_���9?Z�_Rx�E�Q�Ԝ:�{�8)�7d=_ʁ����Vj:������wȝ��.����8�vܔY��xa�f`���uQL����-J�o�s$������y�}��2Ohج����1��c��ld0�c91d�`�s�qߴTu?af䆺����&��w��'f鉝�n-�g���LG�0V�b�� ���m�h:�&<ꡝ���ё����nmQ%f���}w�b{��ʓ}Y+���^�Wl0Y�bX��ʾ��cz��G6ʼ�T*�5?3��܉�^���aO��	~X�Ɯ��$C2��O��i��k	B����F��B�f"��l�r��f?����`�X��a�>��`�U �h�1��Bn�n)y��ft��*�l��?f�̳�����.�o�����iRە�Pw03��vCP��Q�;���f�%�hTԊӡP�s' �9��8>�Ӕ�5���D����������[y�о�К�H1�����}E{�>��+�Ju|�OKI���)�bJ]���о��{i+�����	G����]�oGkN��F�3ɜ^f�~�5�Rn<��JN��
���\U���ҩ����1�>��uk�	�O�y�(�?iIV���D����0x{��yT�i�B[=Nާd�/��PY�����wMv�+�Ԩ:��k��`�1���|�/�Lo��D��iΝmMĖM]Iσ���$�4?�������y�#m�}>�����[��e��i�S :]ƽ-�n|�t�+-�u��g�6���S��y����DF�{��/s�Aί����J��.��:�r�-��/o�Y�b0���ÿ�=q�)����g�p��?��U����x�Ѕ{?5��PM/?��~y�\�h3�������(�i�~Y�eo#<C��q�R'K	+�U�9�oo��۷G9�ͽ�'Ͻ�i�k���Ҧ��,,.�਩~�*C�V�F����Ia��n���5�ʨ�s�Jp�Į#���-��/'��î>�`��6���</)�Ʈ�d1��S��`��'�@6�Q����	/~�*9K����7$oj����#�0U���
� �c���N�F!SOzټ�ub��~���V@�g���&BS�
����>x��Q����+rg�l�5w$��kV��5�,�ø���F���γ*�X&M��LoUsC��ىL������G�I%8�-��+�g���np8f�d��~!�v�$z�o�b��:�SU�
���]��
�`��9��_�:�_������e�d=�o��>o��#�+K���'�ӦFM3�KH������$�6.�rō>����mge�!M�f��mE�3�bzx��Zea��%�\c0vce����iq�G�W�j秳B�jǷoy�ܑ�k(|q��LȈ<S�6t����4��'G��N��,�;�a�U���B��i2��K�n���o�d�ugJ\���x?,H�V��O�)E������>ù�w|�y��iXH�1� �Rs�ͰhH7���An3E7[t�>D:�0D��K�/�����I6���2(���ċruz���2
���{�k[~�r��J�5�I�l�Tjoy��S�h��c��p�_��2]�x4ٵ��w]�����{$�Rv(z2���v�|�Q�1b�Ȯ�U��n-� ST?�k�B��2ں����o��o�����<��(��6�_��9�z]��m�^�;�lD@h��h`��� �U�t�v��=�?F��kzi��O4�.�
���P���x�So9Clr΃�c�P�����a�.8���}��/�>��o�������)�7�K �`�M wZaJ��:Z�U�V%}_�O�,��L�>���XV�O�zg|vڇJc��f"[j6��	�a�>���6M���� S����<	��4�B�C�NR"�7&f>I&o�]���4;ucP=��g4Yj;���<I8�����Z�g�^��(�g���?�9�	=5 �M͹ ��oe��OrZ���Q���E���f�w _�2L�S����F_�[�������@ӯ��ڗ�nZTN��@�椛�e�HT�U�la���8oM������ٰ��Q4�]z�t?_�
�Y�U�3��r*A��s�|>�܂�qqx�!|y&fޗڰ{��l�g�n����'���^�I��4��
�.J�4���0��˪������>����[�y�A%��:E�K�C����N@��Dz$��%�����>7���:��A�pk��E�s0��O�W�>��uL@z&�A����q/�E���xaq;��u�������*�Xb�c|�)E�6e��=���ܸ��9m,��!�# �f��Тg|V�:���"�+~(:�^���é�ۿ��Ώo?J�������ߎr+_+�P^�}} Q�ᦽȺ�'_i��*���M�Fv
EK�i%�.f�Ea�lH�^u�4�=��>8v6����%'����.^�Lo4��'�� ׌O0W<����'oAR9c�����[W8�����$�V�9=Rg�?�6�;ϑ�dL����_��Ws�нiuOﭮ�����y�X%�	��J�<�1���`��������d��'�4��{��	��\$%az��Q̹�<�<��vqq�X�;$�.:��b����4��X�����3s��7�l&�Mq@�cPT&nW�^�M6�͇����OuJV�KV��T=Ye�&�#
�����spt,�.�Y|V1��ӦD�OFЀΟM��gĔ�i/Q��G����@m*�=���t��%�@߳Z[�8��w�^��|���|Ux>�5��1=oZ��F]���؏�:��<��s�Uw�-���P@g\$�3;0W���ރ0���!�Y5�CUlO�����@|��PTǀSG���(�)H���r��(+���.�^�f������zʀ�\���7�?5,�Ḋm���Y��-�>o~6n�-�ȱk��������f�.E6#�@�u{|��j������s̏�����jyAm��=�������>�} +;⬩�:�a�}{Ν?���j�q(�2	�>��~[6�RԘ	m5G�<�-bcg���x+�k%������VRߢH�������V�(Fp����W_��S��GN�8���`Uф�����׶����'��ܱ����<�;=�Y���<�/s����Yi�Wࠨ6]��J��Ĥͨf��4�X����_���<Xx^*X</�i&�
�,F�a�/+�K��,Btg�*h���d鵟�i��1:�:9\�ފ�1�A�����溱"ӌ�v��K��|b:�{��YgB��To{����Q�%eZ�y��=j����	�Ĳ��Q�pM��J��3��WJ�J���tG��,����5�w��g���ה�ӰY��(=tu��I�r��W��<Y�j3_��&�m��ʴ���3����Yn���bo�q�y��W�/��_� ��c�b�3����6%!�d����n�яD��}�8�>aK���'�H�x\��x��qZ�Fޓ��NW��u�=�X��,:�U����T�?H%ɼ����i��l%y��oͯ����庎k��J��
�ώ	��-(����ɨpl��RD`���L���~�SHF�Y�Ny�,ZԠ�0C�4�O5����[������A�`��y�"�y�ې����x�IWi�'G�;q�e�S~� �?G�:�&�����'h������r��I��ÌU ��ĺ6��3�}zA��2��H<1����G�u,�����+�R�_cR��6Qx���"�[�~�
�'c{����>�J|6��c���S�
)Eƺ!�EO(�G�k;`&�ؑ68����Pp��p�u��8�)X�	߅� G@�b2�c�Q��!r\�P[�n��T���헌9���!�βfB���X��nl�?�JI��uѵ�"0k��*[�@�Qw�L'���R���{GU��˛�Wc��w���'�|��bJA���g�_�ْ������s���b�����6F=_FD�w��1_-.w��$�}���'b=4j����Y�C|�
~>ٳ�N��X3N�_�����7�����[��J-\[<���uS9x|�I�(��9�sqUJ�/��7��#D}�vH-�L���l�m:ތ�s-���bs>��T�\4������|2w���s��g����̣/T�<��u$�:~�7�JV��n���Z�ڻ�?���1;A�`��9�i+�{���u�<,�q�89wB=�^&�e�8w���^��8�:������7�8�>�ة���ΝR%फ़��4IN ��Sl+�#Er��0��Lv�O=Sc���YO�8��u�Ó���}qa|e,^:v6}���������M1$�O9��a���AF�7sN!zs)��p���!T�SJ�Gs�N��V^P�)��A�OR��+P�v�=+7�����R�Q��[Z���8
�h1:��\��W����:0�;9u����������1-~��@�m�q�K��+�U��ۭ�X����a.�� &�U��~�g�!
��N������a�|R�_�r�B���er��F�֝q��e�`����K�C�+��+��FG�|{��y��闔�c����Rݮ�C|���������Z|
�t�Xy
s�3�m��Ј��9u���� .�C��3$��D�o��A�'A�\�P��0��l4�%��ך"�\�o�_u����;�J����ߋ�#�.�s��e�z�հ�b�M�Y�+ı��q��رd�
>�ܒq���|��2�uֱ��
��S�0���J5BڮBd�F�Di�"nZ�#ɜ��T�>�{�Y�<����OL�d\�#F����SVD}]x�L�C���Fs���f����V�xby�g���?N������>9�$�Q\�?E�g�N�X��$�^Y$qۈ�Gij!��m�%��l�3?'�R����	�ŹS�>��dq0ɀ�B.�g[�!Õ/�8m����kPj�n,���U�z��w�~n��8v�j���@^����ui�z���9IIu��Q���j�ǭ~a��>��mv��Ɉ5�)8m�3޽����mN��GD��f��:���OH�&_�VӱLl(Eal��X� H��N�[[�ʙpA���:�&' �!)m7�i������d2��̈#PL�. ����O�C���e7A�q4I�3��\�d��&�����~}�J{B>�s8u��,�36%�p��V�a�y2�4�WSnK1<c���e`�]`h\RMP��9��Q���6�m�+�����ּ�U�Y1n��_V0�.K(*��bf�/:7[»���/����P�"궎�s�]8u�g_`:_�X8�FWk�+h���b�G:5��c��5ۺ���
t�p�߳2��1�S�ƛ��<����}ȅ �KN��K�0����/�;�	2���_��_<U�S����W�/���f���_�2ϩ��f��Rˊ�<c���\4��o�v���eߟ��|E�I�s#7�O�m��g��w�h��� 1�r��9ư׫�0��)Q�ql��sb"�>�//ɡQ��m��j��)[u9�1ۅ�:��l�s���Ⴌ��LlO�Hj\�V���&1�9�Ӕ�3�i|���i�������؂�5�?1P�9'E��Bq#�����q]��y�@���X7���9�p��6<T��P���"��%��@�L33�	ǩ��������g�]#�u,APvf������ܝ~�J;$l����vVuϨ�iGH��j���̨�Q/�I���/��ԙ�w$F[���?黕T�:@L�ū�:�*�@�Zf���*!�V����Xo汖��a�V~��j�5�ɱآ� 'Ŋ_8|nR2\��}WX䲽�U�_����Ԡ�/#��-W���=�F0���Z�}����t�D��8�/e��!TX�Ƥ`�?Z�B6x	fW�gm���_-]���"Q�Ϧ�!�'�ߪ�;iNN�r)��Ԁ6��/�~Ѧy�`���/���[���b���i��)��?�CK?���]Y9e9�S��Y!�z�<��}��.�L�/��ܸ�p��>X �f� zԏy��'a5��gnzԨG��B�N>4������$ϋW���S�ӒX7U�D��:)v��C{sR��Eȃ�q����4?�&Z���	�_�Ki�b���H�F������څU=��B�q&hi���Zn�0�Rc��E_�F��yu�XY/�x m6��f�В����BA.��U����W�]\��:7'�#wUO��mMi��;����ē����߄�j!/sԺr�EU������s�C�Y��%��q�B_������	'��)I�q�,��&���?Z�<)����9W��'�./f�]ukݙ ,��?�i�Q�V�d���w���6�7�/�ql-vЅ-�Jda��cv��L��fjʫ�a�]?���tꃯ
R�xWo�ؑ�W���Ф��c�=���k�;}���R�
U8��3e}b��ʯ�����v���j��,��]�q_^+ �a�K��yx2�v�ԿY��:X��ʿ�:�&�iA�| ;m�3��9�c-�RKe���e�GU�3����ԩ!��;�o�(Ǘ[�r��5��� g|!/�~���S�>�L�������CeM�yt%W԰$N�t�	-���s���_^������Ē�� ��%^�B�?u���[W�q����U��{Y3ֲ :N�Q��"��I��$��T�P����\Y2v���Wi���7��#}Q���� �� s��L�V��]��i�1���T�Uɵ�m������N?���(�U����K׀K���h�o�Z�Kfu��gL����̊�ϗ}���w@a)���ب(��e�2�C@���-^���\��'��y�6�*��?ϴ��W����,n.ǘ�^K�c���IB��V�9��~U�ԋO�oj�(�x�g�\X��k����p�����~����K+�
_�/]7�ωD!JZ��3�.��_7�[���J��2���9���7�V�o�8�֘*��iӋ���y���_���I�'(�7�W�Ξk����:�KԿ���)C�#�T�nyo�D�c�Voj��8�,�`��,
L�4f�l�A�Kv��'���P��m�ʾ�s̭��ȋ�����=��~�w�)NI4�S�Z]t��%cN�������.&�)��	�2p���76��B0����(�;$$.}j�����.߭�J�{��2�Ɓ��	���8��k�տҌ��l�7��� Y�X��ؿ�i�Jc��A���5���g��Cע�|sf�c;ڑ!G_�ol*D�1��b�.K�P���c�����;���||��D�$�׮�����q��^��f��3��O.}UyG�g�kݪx<�$Q�ՐѮ�7y�mh)�P�鋁��ۑ؁(KA���<4�����G��Eg/v*,|�aC�3y�gϮxs��L�2^J#yq��W߸�/�ۯ�ov��jV�����d����x}���'~���a��$����k�h��
��Lw�k��><ߥc�#99��9������7�'��׮.���]|����7*�:�\�n.7�Z;��T�i�����>}��eV��u?��i���M����N[�sGY��s�8�f�!dp˟�1+�,��1�� KmB?ӐZ��x�WǮp�A-`q���|kp�����_��+
��'#���k�+!���u=<�B*�8�੢2_�oK�5]_-��ķ��s����>��S��Mہ��0ns �)��Z��������*�*�U���tѶl�$�����y�y~�N�#��H;\�g��
�3${a��%�ݬ/W�#���r�EW����hȡ�g�<����f��c_���	�DS���A�?q�~{~��s��FLs啣�S�X�����X�>� C��Օ��M�ZOK?�Q9�u�^6�,Z!ZOp�e�ȓ� �,{��RXK[���齖�\i��H�,�j����+P�&I��ö(뼼���V�S���o>�0��qb��MaRfc���;*�qF�-�T<�6D.�&�y��9u�1�,2ͼ�e�����̣�tӵ`���0}KG-���G���L(��C@^==�x0м]����v�V$�@���U��>��{a�M�R�A��LK�����hh��~�me1�?6��(��K����5둺���ԙ_�/-�
U�K���]Trq�w:�����|Rs�%��C��Vk;|�����<f��Mc�����x�t�r��6O���_���	���$J�kV�߸*(Y�@����̯_qz�8���FMrf���5���I�b[�v�j�����SnWZf2�r��K�8`j�ِ�V▏��0�=tM�3�XX��n����(~m��y�_����I�3�^?��nN�0�o����!>^�}|��� ����<4���uI�qI�/n�	�GD�mk5�f�@�L['�;m���g�kc�N���dsv�yn创�F�דc�d؈��ŦQ3TLۭ8��Z��>n�ԜrAͦp���$�o>_�����<�}�����!;Ž��|�p�[zzz<�|���F��n	]�z��5-�WEB�G�q}���1�ƣ{�pD6�b�g�=���x�ze��~n�>�5=l&'A�L"��Mߺ�ӧ)���5���a�~m(^6�'���x��yS�k�� q.�F�F6: ��g�-��`��c�S���m�	w�0�\�4+ �ϔ�-X���7��Q��e(�Y>U*��QX�|�D��J.�km�ɵO}L}���ʊO�NRTl�hl^1ێ�b�^�/�I,s��o����$!w�:|��J��4��g��`�| m�P���ƓzN�w�/��hgs��sE��(���'��|��a���,�d��\M�+R:������Qg�i�$K?��uq��<����+���:��II�������v]�k���&Uޟ��8�\��I�L�&[\���e>�s���[�~���R�ҕ������M�q���:ﱷ�/�3��2����Fe�/'B1N�˓j���g�I�A],��F�[:>=�mLX��
���xv�~�m�O�V/.�on4�#�	�I���Z��o^���Y<c����CB�0q� >	�����x�xȠ߀KR���>nq#㤿r	��1���?A���#�q9�`��fL�,c۩0�ɘ�fi2^^ ��}�s���"��ч���.�eZ�߲x�mY*�jz���Ձ��,Q��(k$ �m�ߜ~:&����Z{�%�D�4"�۩X8z��3c�c"�֓���b���!VL���b�8ςVɑ����]��W�"�M�aP��i���ץ����ϸ_@�]	����gr���bB���w��	���L6�w�{�,Gxy�ȩ-���,Yt&�	��A�$gdr E����j�/_Y�=�ڌ�y��o��|!�]�2)��
�\��ŖH"Z���s� J���`zk��P"ݘm굡��qn��~���ږ�d������d��>9/\���;�k��&�����x��\	�9jW8�ue�t����T�G�P�	� �;�lhk�d����:ک����pe\���=Zg?�#vH���w�S���dTgY��R9���{�[��8a�A>M����Ky���ݜ���R?8�|�R{X���������L�q��\7�o�.db��sn>|�i��wS#��+$;�IN��e<���i��T_�(�+
i&��K<��%����va���Fr�թ�ӿp���STV~���Mʿ�U�`�S��F������!��w���L��������<_5�ԫB�w�7a<�O���O������{�����V�Y<P���ɋ!�8��)b�kѹB�i�ڴ���rw���8�� ���f��߼������3&�W�m4U�:];q��x���1���˛����.�z����7��h-9-PB-�����}����`� ${��s�ǈή���y�,��4).��(���0���*f���@q���'��W�8޶�'3���+IJ��>�9�� ]u��D<&�s��-�o���wUݩC�8`&ڌR��>v��-�<5�H;2��o�݄3���ᙑ2��o��T.�k�qU�j~z��c����ۦ��k#�?GEA��2�=s<Y��W4w�7��m�3ec'�G���Lц���p���s������{�J��1���R%�����4̇a�{�p��h�K��֫K�Fs{q�e��c>�kY���x�I��̀�Gf @�^�� ���������v,�JƯ���k)�	�԰�J�~��c*�L��ʘ=DTy�uGrFfc��g@Kݡ�����$a�T�˫��5�+��e�
�����8���2~�Ə��%t>�6䦙�#�$�_j[ψ1>S��J��;�����q����� ��w�!g�W�|��R�-c~��� ��2��=*k��19�k��$�ǰ��722yrr�]������gv�s��q�����̷�,�����/f��wze�U�U�'/��dK���x>deC�^_ͣ�/������c�͓:��T���~r��ܪ.s��I�^n��l[�lA�ߟ?7��n~�ú���-L��f�T\w��C�"T�H�$�DBN{�&ʼ7l+��q�U=e�q�)>�-L'X����A��__19r�`U�@T�=�<ocy}!E\\�`�'�����MH.��8� ���7&� ���*�L�1��A)�ޮ�]Y���6#E������0���K=��8f��W��~����%��pZ�u��:��{���il�Q[3|t>
�7��)1λq�h���(�^yttw��=<���UUY�V��w���:�>ʆ�hFR� �a4(�ꨯ��W#O���o��58}14���Z��i�r~��/�	@��#�,��3Q�� d���rl�����y$��t:�ȇ�lw*���?��	<���8u�̷��N�$�kk�Բ�tt�������r=�&�Ί��Ѭ�X2��}�|r0���1
����i�|[�$>��5����	O��UVz4:�=�3V	�����u����L0����u��'��re:䈿��#�*��ܓ�s���)�&��Jw��LfN6�(������c;���\{/ՉjF�d��$��z.�/5��l��eC��ߨ:z��׮E�;�ŧ��Zb�u6�v�0f�-��q{����l��R��h	x�iZ�1����To~��Z`�e'���.N��~f�;�Լ����r����~�[�y{S[�o�F����?qݯ��2¦n�����vk�pb�]�!{�0��%��V+�P�G�1@i�ϝZ�J\pq�<A�����`�Ei�r޼|�2�"MAG.��=���p?o��5�廠K�����yiP�?x�"�@�"I�Y��>���69V�&I_��=A�����L�h�`!V=3�M�3�$�l1t��$Մ��A�:�I�<s�7Ί��p�e5����Ic���-���c�në+�)}�u���O��d���YΚoҼ[�2}�������f�?��������ڕ3O���ί�����`v0�g���w��Y�p�a�>��a~����IN	ǫ<�("n�Ƨ�)U�M׭��+��tl��8"UK�_¦h�-F�oyЈW�a2u�Q;����uoMs�.F�������4�E%�	�U�􊯂:g mi�ӣ'%��u���[%	�m���w9�N����ː�L/@��ƺN����V2,C7�ت0:uf(�X9��Цւ惤�������:[���rС�݅#|>�t ��ܗ��C�����!2wPmuC����x�H�h�;A�>#B��b�`��c}Fn���Yv��p�eS%�<�̨Á�C���z���x#�¦8�씭�+�l_��R�4D�v��$�N��������knUiK+���d���2/�� �P��pֽ܆�ε��p�WԦ�A��i��&9� ���}.F���ۢ_ȝ����R4����x��}զ�$�}��V�[�s� 7���f�.���hc��}���9�-�!2+�8Ζ�c� j�u�(��ߡ�.:+�q�x��G���y��]��C�LJ�O®?���r��@x��r�u�ў��G?t�~hӤ���;���Aۏ7���i�!��~6r�͘H��J��ɩ)�7�%�h:�^n��no���`��y��w��֙j�Ua,#�Y�p��ZJ�u�ZXrRhk_{u<���8ܷĄ��k��N�}FL��qф�4h	(2Zk���*]���z9�8�r�nT��j����vuFܲ�s��L�s�E��#����x�f�J�I���vڥ��G��}��8�nw�>�:�D�~�آ�g%L�O9a'��w|�b&�r{����)���Ȋy�r���;�Ȍ�a���´b��������jU�q��ѹ3:���V8�JYcS(m����#�<�vh��7�4%���ws�ũA���?��Ӌ����m�"2e�]��n[��S ~�
Z1 ���x.���P��yA�(<�^�EL5rc�[�O�LU�2͛�O���6���6���n]�������q_�D���y<�MZ�����1@�xwl^�x1�0���sn�15���ӝ6 ���]��ع�������x|��b��=�����N�Vn�E�F�D�!d<� �#� ࠦ��Z"QTW%:���N+��RA�s��)/��&ߖ:6<��q�픾S�o��8Fpn���~b*|��G���Y��:;�e]K�A�2��`��8�2�虞̾�&��ɶ�z��Z�W�ū��g�m��	ǰ���6Π9'.򗇆��4j>�d�W������揱�yR���w}D�e_ ���eUf 7�Z�l�&�ٱFr0�W�.����g�h��@�%��:��m⧟��Eʈlg�wD/y��5ϫ��_��p��i���Œq"��?z����c|�'Ե�k��������:�@��W�(���vy�X0v|V˔�+9eSmW�.[��C��'m�/r��Y՛�����Bw���PeV�k��8������������t�� ݱ��D?�Ͻ=�a�r�8�M��a9�ɳڹ������J ��2��^?m�,r�!D�f�Ț�����ޏ�}�e�mH[@�����br�jZ��fF���2�h>�fFi6C.8� C$BZs���#�(.�Ə���9���lWW��� xQ���,@�u�H.�Cg�bF'Ϣ��ə���݉x\4^ƕ�?�9=F�+���}���C������χ$ؼ>��E���`���"�

3�|���́XV��-�H".�6�H.�N؄�{����9���گK���י��_ԯ��)�u�K8E����A+$C�xs4zp-�
��?�����-I��v_]L���J�y0t�{��~[ݾɇV�����uY�����jK>�iw� $�6�I)��B����ns�e�xқg=�(�5� Ӌ�Auf]<[�|j���L.[�1��Ƣ?�8�������7z{{����B/�s�|�����3F���;�p:��V�[�Vu3>�>$��>wQY粀��_�tu��C�)e�~꺨3�7L�2�V�s9(t=����F�k7����ђ^U��>��۲شt����� 2l�H����7��E��EJ�2�Oϣo���W�P�T�]�Y���_��\���݉o��1r��Pdb�M_���`��rgcs���9�>�N�I//�\q��ߐ��sc��b��<��P����遗ˋ�_�~_�̱�fxm�W��g�2�1�oa���LX���,ؾE1��r�)�+ǎ��[�#�v�1�}]Q�v7���m������_�����̖x���X�<BmT�u�Z��p]��ឨ�84�hU�ʣ~`��)�El��ݎ�q�_�x~�
�O�)��_%!F�C������)��&�v#��=�8n�%�Q8,�B�(1ʟ`�'Q�_�Y���k��&��	�v���N�Y���.��eRްJ��0>�����t9ir.+B[KQG���-�T?�`��k���W��ftz�5z�\`kg�ǎ�YVy������x��C�4����*N�iEW��>���!��� ��^� L�:A7\�L�Xr	Y������X�j��	Ի��H�����չ8�í��r���
 ��u�ogE�����͛��֜-�+��5�/[��s9~��H�� i��mZpu�����3��U䊫h\9p Z��y��l��5|!��5�s�D��*/5��$מ��e9^iG���P�p^�hgc��dOPwҤ$���x��A��n�t��<�$���
]�����z8�����p��q�;��7z{w'��?���/��t%'jF�`aN�7�E�B�;0ޜ`b�EQ!9т����<�����<�m�&W���}V<�ǋ�?|�ǈp�1F͖;���hq$x�>�Dϼ����F�Wkn��{�Q	�w�X�u�x2V�,sbL�ɺ�{ߚ����b��J-9���Pi�=Pk��t���1:5��k�gf3\�rhou�^���rӮ�scAv9RGk�ʌ�g[}����ph�hC�2��\=��oS�~����s�Q�k-".���?�c���cEM؎�5� ���m�f7;����V�E���8d`�o�!�mj�6��P�`<�M�Go��TD��roӼf�4&OX�L�"?k�^	�	�U
±�1^�a��w;ңp!-H;4������;�;�������α�( ��=ӿ���pRD�9ۊP��u߷{�c�d�@G+�j�M�\ҶS�D��+%����P�G��k�������]>:�GQ[ٓ_��4�A�S�SO���\r��^3��q��c�<9�cw� �8}�z@��O��ȣ�GְБ�q��9��6�V���C'��x2VP���'ѵ#V��N�lPN�`5WJ������<�������U&.������^nlGR"�ϺP <R����ӿ��֌�����x���a���vj���]���o���4"	@��gl�XL�o��]����������B��ᑘ:O��U���O �� L�Ǽ��<^$���՞:Fx��i'9t�áx�u�c��#����?{("9h��}�v�3;*�T*�;j�����>>>�ξ��r��W�SC������d��ߖ��.i�τ�ڼEY�N�	�\g�Q�M���Ͻ��uYP��ksi(��E%yb�\C\�^[�|L5�_Eiζk�Vƚ.�̵$�l���-�o�64�e�I�&��|�I������'��?��"QT�dr8���	�,���������^��K�]� ���'蓓;Ry�F�������h����t��ĖTu�� �WݢA�Y������#��*���(������1�!9N��:������D��<�T��,G��W����;(��1>�7�|�(R�cTs��6��/H��"��D,�Ӧ�W[A�٩�6��|	�_a�]�7�_��T�Ȓ`��N�J�m��pK��u���A{ӝK��Y1�����礆�h�'�����=<��+)�+�d��m�#�z2�}�A����4L�4'�QH������2{�����n0<�0	T���kN66>P�w��2]x�׫�Q���Ƿ�Fԝ�ń�o�
hg�݄�&?�[�s!1L�̔'K�I�fO`I�J�=�_�n f�Wr�ֺ�5��U�^�����y�6�DI�LK��J�LS��V� �Q��z���Yǝ��o��E`*����jo|(�įk�\�B�MW�����3]��7�p5U%Tޒ�:HO4�U}��: >��h���/Lz�3g�vz�P��/a��PS^�$z�!��+�xf!#
`P�t�$��*������o^yx
"@��$�~���%
��N%B/��0��^;jt
-�2��'� �[k�ߜ�?���ܚ�c=��'����0��ӟ6:[t�N������?����]"vt�V�0_�@����<�;�l�E�F��%���(�n3�k��8��[�M��\�&�5w檣@O��}ʠ�D/�ʠ�-9C3�PzVg˵`�8C_$	��b��ӹ��lD^d������"#�!] 8N�y�Z0O1�F]%Y�s'�M8,��9���y�E��2��t6��f����_d��<�g5r2���K�ʛ��1`��*�������uKy�њ���]L�;v���ƌ�'e�{�h#s`�H"����<�k����:q�S|�
�U����/\�&�*�&틅�@r^�j��+����2����43�Xn�%f�9��v�=yp���\���޸'*�HoQKmN�>%�=r˭w�h��w�7�4G
�nVs��I�NO������cQM�C���"��~8�+m�Z@!LV
��W����'���}�����T�)R1m��!Yi�H}@�n;���T ���#A�Fx'�L��M�qq��ibg띇Ʊ�����\��Z�{!����L@�'}��=�IY.�W:7����t_�Gk>�G�,Ծ�Rx�;��V:2d��������2����]��Pڟ�>�M)��ܛ��2i#s�H��M1� ("�2���VAM~����`D��)N�j.�d/�� ���&��'}�6�����'���ؑrt;�r��"87��R��վtW��v�;��2ŞAg�K.�o3VcB���᧌�� F@7^����;\��$0X��8|�ç~2�6E"' �'��Մ!�
���k�zN�ޛ����վ��$WW����lT��ǈ�`�^D���z��%��>zL'�\\���?s��OQ_�����v5S\�.ԟer2��ZJ�E�20��K �'x��ϔn/_r�0�������_r�~�k$��+{��f�}yl��.0��H�����7��蘏Y��Pw<s�}��\��S������
�\�"�-�M��E}&T������kX/�R�����'��Kj�<�1�W�t�ͽ���X-z���lk�_�DӐ�����>�L&v�ݶ~x탐ȳ_�����X���Oe���xF�쬳���ݩ�B3�s�O��lu9l�^�a���A��|}�ET(*
8�yK���W�Rڂw�����[��x*���ة��3>k����Ϋ'
�2�հi��[�K�)~��@p�a�Ʉ���m��'����_�If�-1͇��I�wl���wFN��kSy�E./8QV�|t� ��\�t���9UD�l�o��9̦Y�y��Р�}?����I�d6m�̺6EĹ��������2�&�~b�=�{��M�;]��\8r������w.w�\��М:���$eФћ0���<&��F%<����<�ޞ��fbٲ݋e{�m;�ʌ�SǎJ[7W@�Q�>u�ܱ�P^2e��?0A ~�D�Z���i41k.vͨkǎ��3	�Z0Nv���p�$�ײ՟�_R���c-{�K+L:��oi���d{���
��G;��Z.��F���ߍ�+!0tL�fc�rF�FV�0���!���~����<�rj���k~H�u	�K+��OV���N��/12��-|��
'����4�v�2v)�l�W|Uo_�������S���7�'5���Wx��
��	)�˿�+(<�����C��C���o�w�ޜO��.-%N@&�d|}��]�����J8��Eu�v:��Ю�t���D���SaN����k�1�
�HZ7� � ��b�~*�wi�b�G���Ig� ������(+�����NV��G�۰�c���Ӱ�x��9v>��=����5��DG<�t���Y�8S���^nT�uA7��	�A��4d|��-׵*���Su�'U�Ι(�Δ$���F�Բįlu�1�V�t�aΞY@qd�����;�!7��\���yӋ-� �x�_��y,;OqR���g��w�o�V;�}kTh��F�b��ٽ�1�Pv�b�M��泌���Z�ؙ��|s\��:gP�H��uҺ<��9�����F|-e.����f�9�X,<i3��i�>�e�͹ӆղ�v��`�9�m�� Ձ�h�,�gt(O�mn�~����)e&'g�vs��7����O�����&Ip�]�)�g�jf�o��gv�z׉M���!$Q��k��J/���+6�tF����IvRt�S������m���+ږY��,���(g]_x���n�I��W.�%�7��V�@�*ئ�]L<T��I������(����0�G�~{�1�U  ��IDAT�����Hbc� ��$&��<|Xh6U�I� ps���E�f�"O����b{ت�'�u�_���'0�V!�"��H�l���gH��Ǳ�}l��/�U�uAW�F/v#�Yy`�'��]���,�Z��ۈ`�*6:wּ�}Kc3cΎ��j%��Tj�98۱\�B8�������C�:" ?�j{����8 #������l�I�\���\EA�͹��Ò~-����t�� !��8�#kz���&l �����)�,�_�$����(0� �j�I&z��a`9ݏv��k����$��[+�8�U�A���fy� w�a�kr�g�j�'�&*�?&QVr8��!����#Nπ贈=SB�D��o����zb�S�a�Y4�f��e���sD��GSV�����'���8W���?4
ΐ5"G�ӏ5U�JN
�gh׽����p0��i۶�L�a}�F�:c�(m��'v�L�~����fG�")n�=�ґ�ulΜ�8ݨ�'�7�#�g�gul�j&.-ˉ:�vg������ő��.b�țd�;2\�%�msr��H�<�s��E���l��Ru�<]\I�{+3N���}~�y��E4���d��<c��|��-�t��H�,��bA�x�'���󖬌��%�����w�M�����&��s!����n��2�4g��f���K8��+ʀ�-&�n�����Ji��to���	�/���-�P�BK�W�ʰ���29q�W���ؚ�����O�-:=v�����^:��\NT��}3b��$�\�_Db��(x�E��r�1Lrh��s97:=����y����s�v�9���3��1J4�/s{Ƿl���*X��e�%�s�-�ĳ~n��]����"q��1uJr@��š�m��[�p˧D�!�6�)b����� �MŮL�҆��J���&�`!��c\N��9%
��?6�M�!D�˸���e4Q�.���<*���Ý���䅖;� ��t�	�W�hhېݞ{ǟ�X �P~�8��zY�����.�$`�>`݊����[GM�hI4y���MoǂY01�n�Թ��������C=��=^߾�E����+B�B������D��Յɥ�dv�}�1ۈNڜ��Q_E��Gic8����y�h�@����̱���8�O�{�L�]C훁�̀�f�����-vaB	Gǡ/f���1hm��O�2��Uf��'Z�Is�1˄<�:���^w�$�O���!+����ӟ���ኛ^�m�bTP��''�[�I�uϺWy��N�Һ��AW���D/�(�.�%q���  ��w�t2B��'ƜL%|����%�pq ������~�GL�Lf��~��T}�ӆ�zF:�RDbWJMh��Q&��'�m���Oi�F�o8���V�K{�ղ����^�y[i7��W�?�R��]��x����fFz�&w���ѭ]���5	*�򾙱☴yq��r8��fPsh(�,w��:o�y�^��c������b�f�>��0�]�& �o☗��&��2����	
QP&�I�+�x��a���S=Q�z�±���[�&�����s���֡�b3��Y��R.�uu����c���(����2��g@��2`\�
��G��_�4&�׺��$z��gs6��������\�;�:�B�G�|����us��o9RHFE�)��#��M�,�1r�.��ߟ�v'��y$>�B����/s��☌OJY}�u'��"{r�G,6��aD���4�09�b���:NB3�C�~�8��p�_��c/t]]Z��������5'�Q���g��vr�it��"�0��n4�iԝ�-��e��gM�*"�	gC^�k�;����L*ߦmn3Ƣ�\�F*��i���'dY�ơ%^r�=�F~�4v��s[��MϘ�������"�y|Ùw2-Fy���-V9~H���A�a����B{D��i�ȡ��,�ݛ�������m���O�yH�������y>����#�Z��rQ���-�l�<��ޚ��Σ����[]I�]�ĶaN��Y�`��.��h��gt��N�����s؆���@W=�Ȫ�<*"�_��ʤ+^o��Oƹ	�l���=X�����x��ݫ���ͱ� �f �pv�����ߞ
������ǿ����H��}�M�:k>��`�	ppq���!��m4�Vc`ƴ$D�����+�r�{��Q���� �����YL��k�\�D�(���0��}�!p�N8;��VpMں�f^�2Z�Ǉ��X��_���{�!��������}i�r�؀v.!��yU/���_)�h.�(y�n��x&����p|�x�5��G�����v3�J�9�p��8Na��1��aNr<��r�١���v6f_}~��l(�zy.lN��s��_j��=�c87*��Bh���#��W�vjP�I�e�Y_��c��Y�.ی�|.-��f��س��#�\֟p�ߊ��#?��<����|A�#�������'v?,Id����+������Jt�暁<�6MF�� @4��_P�դ�0|��ى^��q�o}��ˑ��>��z��ׯܑ�յ�;5R��4>'<gv�r�����O�B�oۛ �~i�͝g��ʢ��q��5,���x���-�^�$Fy�:h&^��"�E6����t��%243Ũ"]�g=��8m�C9�銾:�g���F�r�����&��߅���9��Uߋ�n��؍��D���>�v�>�����(t�oݶrZ2r�������
OǢ���	?B��\N�7�ZDզ�������}{W���L����c3�Ctޜ��a� M����B`J:�1��?]'�[󶟽��+��2F��0Y���&����t��u��l���g�_�;vp#�&͝�kZ��E��u��c�o��b��N��i"6ܾ*(�����u�'&$p(��?������gu|��	;���|�};;Ӑ��a�*]�L�*�|�Q�=��4B� �̖�J�SNv�QSg�є�}*���� �\��/T�S����9=�i��Zo"ڑ�Հr�8��.+3����*�E!2/��I'l��G��w�=ex���}��Hr��1�����h��(�Nw���n�v��	_x�&��kp�Jz{�G붙cg׎l��ƒ�`�*�gqoL�ڡpv�����~<1�z��/���_��������E������3{W�tlZ^B�N��Jg�0�������+�6U��)|��!��G�bbʘfBk�rZ�V�6D����+�c���:1Қn�+k��7d�`(�V'��BergY1r!�M�K���{ χ;i��Ȣ�����V����oM@n��Y;q���s+���F�P���xa���S)�9�H#_�A�VE�_��2Op���኷'PD^�Xu<�}9?�<*_'^߈?�祱�t9�z6�$�N�����8ue��\��Ϯ��>�vs�=���m��w�|9��F�m��V��l|>�ן���_Rd��(i�W�N<8�V��;��m�&�>ʥ�+��
�Vm��{ߺ*��vN�ѱ�M��D����~w���-��|�C���8�B֙��2��3���h��}ާF��N��1��L�z�y����ӫ�"�<�pw#F(�Fl�٩�M�8�6�Lt����x"5z�.���)�A��w���۶��������廴Fho'����￉�/�t7l�����g8�fۆ���>UNt�i=�\�$K��`���tʑ�<���vM�jc\�������<ֈϘ��G�o�o]�)4�A��2[	���ש��xI>3�cƒ��>�̑�����즎��P����y��#�y
���K�˧���D������a�ٻ�U�iU�]^O���h����i��7�?�w���[�-��f�f��	�,����dd��Qdg%�/�a���/�s,;�8��FY�rs�|���㗖����%���Ö�ܛަ)�Gn���[T�v�o�Xi��Հ(X�l��n�ˆ5�D��"���g�Cy,���Ӡ/+� ��ݣ�p�s��RD+�����]�ƚ��<>ù.�p2HlC�nk�����ȗ�>�#��l�ЃF'FN<����L�g���g�?�K��m�<^l+�c����<3�H��1���CĎG������ޟr�.�!$1,��P�o|+{�S�gF��n�i_#@��j 'ɨ,��w��]i
��< j�<J�ɲb)^���~t��D�H�ϭ�f�K7a��������'mo�o��p���D]�7p�x�g�3`�����$�T� .��r��I��֭ �M]��*#_��+��V ��*Dv0�.��M䃱E���G��U'���B0�!v����e�D�o�3B�
z"���N�a��I ���C�#s��]��1�Q��9�?�5����	J���'�0�d[���� b�g���H �����q�=�F��Y\Ǿ��Fr�_D'I�hgj(Q�e�;�kW���?���:����QL�·�n�7�gF�;cG�ǜM�:�z�WFyӀM���JØ۸�2����:����C�ROƒ ^����O��/�#�	�����c��Z���G5��
���a���r%'�z]�"yr�;�,�w� �Au�tE�$���R��s>�o=a�N7��=��7s����m���ဦB��7��ꐈ��uj"yA����%绍*��D[�r���N��u �3��>���g?d,o©"m(;v2=��#�g��Vu���e�mȚ�ð@#���|�+�f=(�&��m"=4��� ��TI��y{b���"9�deP"�7��$Q��}[��/H;�#R��k�1��=�Ձ��#9�]fc���l��1��Ă�q*�&z��{1��s�����9l|Ý�C͕U�DfSlND\�w	�a�5�s�Kˠ2�S;(���e�8^>?h��[ːI�0�y��9*��1}�c�x�/��1�r{ ��y�ہ���G�U�L"���z�3�?<�n�Eg��v}���y��8v�q�v�C-��,����6,�_�J�Y���&D����a�'N��������;���}���mzf]6$��U��_�d�Zc�o�M��Cw�^[���h��aq�c^t���u!~W3R�s;��V�E�-�P(�E�ρ��8ڮMh]5-q���{c�ꐔ+˰�+��\,�0�+]�x������2>ja��,E-+����HB�c��~rU翾���׷��Mo��{O�����!9�I�so�c8[["JLS���c_����z^��������g�~nE#�{(���رU�ׅA�}ix���O�#{є"��n�v t�	����ލ�w����HԘPf`���p����GQ�/I���9s�T{'��3]�NI$�V6�Osƌ�ֿ������lX[�l8[�Є����Oit3���H��$ۖ��##�ln|�_7sZyK�y7y.����wy�����C�@a��"ؐh�5�7na��p'¨�Z�'6큗bTx @�� 5�t�����d�<	@K�5͏�]`XS��T�t1�,Q�	o�1y<Tk7c7���}Sy�Ǽ��sO�>:����q��%�ż�ו4k�����0u(
�vJ5���.ؔZ9]<��%�����a����(#ո��yA�`�JZ��,Q�O%}۟<՝��oNc�s	�	 ^H�h��ɑ4�6)ajs�Q��.��d�j;�����H$��췼E"Vř�1�4���$����x;f�K�se+< ���.Σ��Se���Z��͙9�h`rp-^��!j'�)�i
$'
v������s<���뿞?�쉼IO3D�AsƎ	��0����ItےsG�}Xd��r�&�^�v��r2�D�6i�L�Mf�D�|�	]
;0�����������o�+P���襮���W�V��"�f��@a+�GTC�`厝��Ts���tC%�tǡ
�1�:��;v.�&�ի�X���i1��%�����ݖ���y��3.9vn�9�nvj��^�w�u�l�|�ӷa(���n��>e�DW�C����;Z6� ���Μ�����fBw�L�jQ9��P�`���5AM(�iHé��ܱ�r~�/�3�:v���]\�kN�����h�u3ǹ�N8S{_Ttl$����\/8����;��u���~�R6���ylH������v���ET̢G�ͱ�$�}�m꺥�g�5�̥e�N~IGwj(�ܩ�̺��F���-n��4�����(����
MU�H��fJ�:{�����.�WY��ƉUo><��˗a��y!�W;YF����o�-���U}����ǻ�|����y��I��v����O\EC<1Lw�G`:�o�X#��ey���Y^M���.~�����H��B�a@��YY2��#��	����wz�iΝ'?��>��$�Lv�v�!e���9yo������ٗ~�DO^%
�2��I�4� "� �~v`Wp8�1pb`��E��8yj�U�����;��Ý	8"�/�%�WG99R���'Z�PȘ�������!ڷ�-��]"KX%GG����/ƃ�����V�/�=�{��Ⲉj���:��K��B����A�v���k�˖�Nҹ��� �e��"�K�j�Ow��r1��I�<Q�8�:y�Z�.p(�\�N��͙K�<-���[_A�&�mç����3@�i@I���Se���X�7�a}u���n�Z��B=�T||X�uP��;,�^���Aq��UOs^�_�#�[ �n��3)��<h'�,�#?ǜyh(]�Dn������|�l&#���W��a�W�}W�Sq��G��/aϘ�UK.�{��OP�}�p�ɶE^�4�#	"��]���E��S%�d�-� arw�l{w�|JT����fMI�򧾰,Ǭ��آ+�B�Ki���aǠ�i�!���ԸZ�ϿsD#@!w=�`������9���/Ϲ���ܭ��$G�t�D�z��c�[����$j���MpQ_,��$�"�M�`��I�d�r۵�!���(�����H�9�����.%�/Q E���Cl�AD��/�'�)O��������,Y#/��d^��=�}R��m����#mU�����|�~�m�ZF8��䤬��� W�>"�-�g%�����Z�Z[?��Z���x��rzB�+��q u+<�S�ta�-=" �\1?���aE��3�-ۿSw�������_�2�;���������+�_^� }�y�v��Q��o}{s�-���*U��)j#h��9�UoA�ΎX��BOck������ٱ�X�l����0�X)��\[
�*�;HX���P�=
��R��M`��{�����n/��s{�m:�֐w�=�w�艄qp,<�DD�|z�Xi�w?Xr/�4�zʰ������_��#'��V,���i���ـL��"f�
vŜ�l�ˇ���7Jϭ.fɄ��,IP��?��򡉕�3��SC�{ԍG <n��[A��(�͢&�$��J�m�=�P��˼�@���^=�4[��Y��x˫;c��?�'sb����J�cU��"�z��D�D��}�P�v��Պa�NP�r��
�Q�b�>��1 ��v�;V�V\T�É��L@�Qbj�F���������m����L����p<m�H=����6�r�̘���a�daS�!?�@��I©��m��X����ۛ�4q�!nS�N���P1���l�*��3�y���a�n��b�UȲb-2B���F]�~_1��-r�8� �%� � H�T,`hE���5N)K�9o�o�y���)�Q1�\�Db��v��:թ.�Y�BO�Ϻ���s�8Ģ�$��.�VY���|������Q���-��|b�4�eBi��
9��m� $+O�!����h,���{�z�	�@��O :�a�9��a8��g��@+��'9���18����䀌4�k4ӡ�>[�7�U6z`u���������C����� ȓ^�9߻<�6��٤%�dtBޜlh���ݶ�������j�yrL�!"xA{6�KrXu��P��mo�.�|��C<=��ov2[#$%��)�|3`�182�����"НH�����L���"*�X�#�_��FS$Ɋ>S�<KE��5�\���+�VDo�vIӘ�n}��^$Rj1&�4��C,�c�JY)�_�a�V��ѩ�7f�Pzb>����u�>li�muG�V��s;��DO���.xp���ݰ%h�'��w�c���{O�Y���vD>�!bg4P@�"+�230��j���b�"���s.�.9D���Ζ��0�3V�.<1l{|���t씶�������d�Y[g��雵�_�9�O��B�V��i$�OH,�;���>����k���B����Gͦ$D"�U����gl\r�seY��ɴ�s��4���k}��$�0��A_��ǉä�<�������_�6���ӗW������}IO�G��rZ�3"vo&�/6��f�T�-�}����);t��n:�թs���̍��EG��z�Q�}���[�#&T�eD�LY6�$���8������~��������	��c����T�?7z?T�=��D����?���_7h6�2����׳�7|Yq��;}�����IAٳ�:�w5B��+��<y����S�~{��Q�2�H�(�ٙ�9N=k���
������Gl'Rg���x��M�;��q�$L�N�I�G/�}�&�ԲL��Ͻ�� �x���?tu�WE��]s��R5o��;8A@Chmyp�N�B�q��+����\8�	���b�`'&��ѕ�#�O<����0u��@bq$4E(�E�N�vܽ}�W$M�<@_Wj-��������u�QI��>���4��ǧ���#������ȫ��wc2VH�Q����+[j���d��wgG�0�n��:�X�JJej7�N�/�>���ց>�Ӆ �$���fڞ��苜�� H[ ��n�'�+}��ŌU=.��9c���?����W��W��9���к=y3P^��t9:���孮6��]'���R�Ι![h�<�S�q��EY!�$�� ����[��>e9/η��I�v�3�n��S@�K"�¦��7>M�Á��h�{7*��o��s�CM{�h���;v�����[?��L}���N�a���NߐU�'�������O�����ǮG����Gl/4cwm �UNl�w��z�������|���ӟ=�SϿ=��~z����?�Aڷ_}>��}�^��5w�A��o=�oѤ�jH���^�:��+k�
/zp�l��fQ}��Ƨ���(�`4o���}�T���/-
mWc:��R�g�����j6�p�}J�r���m��-$������ `�IΦ���vӭݢ��i�S�yH����@p�#�&��3nFL�iΗx��۪H�1�d�-��$Ps�����IK*3m9����5�ݼ�����#h��T�"�M�u����}Ȟq��g,�[r�~H!�Åz�*�΄�xvl�h��V¥�
p�u\4:�a�73�҇�<`9�S:7�W� �;��	����d�_�^���4:^ǖN��l8�Bp�a|=�6��i�#i[=1>wH{��0��]�-K.[$W�!�6�.D�A��M�$�Z[o�Y�!pAD#�\���!:�J�I�_�o��if7�1 �;r���3N� ��B�'�޻3��'�4|"�'�HY=P��CO'c-��v~�V-YxqYcNʇn�Ʈ����f�/ij���YH@K� �l�c�w��CM�)�n�z� �Z�2���]�?�HO�|��}*!����M�a=���/�K�'���� �щ�ɲo���CG�1������Ɠ�?�S���ww�������-�X��t��Ձ��&�CV�>�@����~�L?�Bǣ�c�;��� ��i{�����F���a�*M�����30�b�����aY:lq�H�Ӌ�81p���>��x�{W�kp����М=�Aޚ8�J�{�A�Oߝi�ɇ1��e��$0��C�Y����S8��x�y�Q��!�~��aa�ø���)�-B��3$4Xg^=��#�ZQ������;v-�ٯ_�s��<�H4��B��"���2�씇 '�@�����_C�^�͔�9w�����)5��ѩ�!�6���В���y9 �}'.���(p8w��p�|��Qv@2 �P���l�����L�S��[CC�F�
����Pl �̙������)N���^��_N�oin���!0W��sS3��f<�c��x����ҿϲF��F9_�R�	�`$b�K�n.��f�Η���E�-U#i։l�H�Ɏ�h=iCe���	���t{�I7�7ѷ�<�d{�I��CJ�vܐZC��xD2d���4Κ��n�C��#�������k�ey��)��9��[~}<���Nǧ�i?d\n�O���	�wY��:Lp�+frLГ��Ug�]/d#���^x�lЕQ/2C�9�WsFgX��,��X�G�?��!���	��+�/����[�fs4��nF��G�r[��Ŝe�w�P�3�(+��\��b�\7���Mr	�ݒf?�z6�D�y�NC�9���V�w�	���y^d�B5�}�Xg��jdf�ȃC9�
 �:�2�´�g|FA%\�Y�Uy�Q��x�Ѧ�����#���.��ڞ劶��ӡ���W���-:�,�y��|�4��szi�H_��� �p���m��#���]Ϙ���Ł&1G3�ù��	n���L�rv��o���ى-~���1�^=�/��~8���|r.��:��FӼ��S�޲��<�"�	�j�v�"�k��Q��#��N�d8xc��o�v�De"���e�w ����n۷I���q����"x�|W����ϲ?�+1�mm�o���^�<T[�{��&4�-�����a��&�Z�M�%�M2W�S4��	����ٷf��מ`�� ��?�՟:u��*������Z=�����_��¤�&x���x�?oo?�y�:�;1�|��#"�xy��N��i7�ؕ�9�؇D�0�noo�lrʶ�u!��G����=�S���	�Lx�������˧�R��I��<`bK�P�UvwH��D$c*��!�Z�6�s���-���l�K��� _d#��H�Γ/�%r��F�G
 ��N��p���Q^yS�q�Zd���3���N��E#�"]`��Ԟ�_$���(K%� "�"���6�~� �4b&A��oŲ-��YsT�z�V������߽ms�Ԅ� 1ô�.�z�.�mOG���qکBٲRI%��Q�l���%��Z�N;�{�c`_|���� �s(A��8��{D�VD`z$ϑ�w(����P��fr�l>F"f(�M��ǪK8o�h`SB֟f�ٻ�ضY���w	�XɃ�V��K�lj-����Z~�IZE�4�c��u��;��Z����,{� +�D3o W��ӶLu����P��l��	ԋ�0��u�ۛs���STb���MMlP+fuO�||x�&�3d+Y���\�\O�ڝ<p����(��x8`%9V�#��4R�ͶK�c˱(tv�9�m[}^i�M����O���)#O���)Oo�	���f=*S�S��mo��"R)�!h�b%8/D`rt�XtV�㐅�(H=�g�%c�>Ң����g����\B>W����<���"\Z �xM��?�M�I��mz����4	��>VX+���'7:�/�;�L ��Q��zU�g�f8�@��Ω� ��j�,��H[L^�V^�u	OKԧ>�D���xM�A/��)�;E�/���c��In�
��s�"j50���ly6쐐��ם]�<�t�8)��VO��Z�+O�qW�m������ҡr}��`/�__|��ꬄ�3��qZ�*A]��z�ŧ9r�}�r������Y7�0A{�5�V�њ�����L�K�B�!)~�񸩽���c3�uK㢲G�eN�c���Z�e�@y �/J�c�v&���}���l~�p� �>>��a����,��1���ޞ#0p��U�u�V�]N��ѵ}��-|?�M��?�{�|ym��p����b��t�#��4�d�~�|���=._V?3?y��%��d8��{ǻӲG�H^�714�6������O�gu@��4b�;x:!�Z�NQ���q�d��b��Sǎm|؉{\EK�1�x΅'�^ӂ'8~�jfP�{���@�O�S ��v٢�P��6 ��c6<�n��$�c}�RH���j���p�1�:+�V��U���T��b�vO�*/Z��,:�TB,	�,=}6�	RGO��KZ��q@њ�79�f�RH�v%�"Z�o(7|`�\2�M���6�j7�
��Ը#���	���zd�cp$��ٕ�G��tOm�v�;�;�A�[5�
$WM$�N���t��vS������~s��v;<����!7�����s����<_;"�Lj��!J�&����B����ItP�d$���Q�i<����3�B�A�����D�NX��&O�z���<��ڇ�@7W���x�!��(�mK��H��0\U����x4 '���ј����c,���(E��]fC�\9�|���iL��)&c��ڶ4���	��OJ�0�y
Dt�k�A6d�f�46�g��SS���:N�'x9�q��1a jK�x�'�s�o����������{r��|�^8v�I��]��HT��;M*�g{�&��.�����U�;�KL���N���o�����/���6������O۶j�������Aq��1pCN�c�h�ݰpr�;�8, ���U��iL�xf}�%���|m}m�r^1}f��b�(��xnN��ų���m�<�kq�?�~�Յ���c�}x�3Zl��s��n���J�� y$0)�<h"�W����:��'%]5��� ��5,>NC$u6�|ld�q�htq케z��
�8�&d�gxMP�%<^�k��	ry�>A�HX�ơancm�.a�]�qw�%g�*����GY=1��n�z�=��k=�^��(s����s���TrzL%��x�&A�Z�mP�ƯU��h�$Q�:�m���4˷�N�H ���y`&9ষ�pz�rg}���0��vH�з�XT��#az2�A�X���r�?�M�?gz	�6�T�v���W�A{��C.��<��4�� �〃Tm�Z�}>`s4Y�D]�R��ί�P9w{���������E����eI���\�.�[��>�����e�Q%�$����ro�}ƀ"��\)���՞^�XV��v��	|~ү����<ׯ�	�I<\��C�`��ϧ��ٷ8unw!�$�mw��}|<��̡�v�4�#�p2@_�����
�l1�U��a�5�ݒ �	�J!b�n!����(�V���o?�zR R�J��������%�.i̱d�~	X���P!���8�
!�y���å��/�ʷ�����?�Ӕ�q�:�a���t�'Z���D~ � ��ߝ��OMZV�`�����o���*s�Vӛ2&�����[Dꬔ
UP]�����;H�-mxԼ6�!8��{?b�3�i#ql!)$�b��7�����&)�7~�Y'[,�!��,��`<����a��)�0`J=�z��L�w?���~be�-�qC��ŕO�Z�T�M/��av�����m�[w�pVz�U�׳���!(e�z��I�V	;_��^t�h�EN8� 'C*6jgDx}	��0�^�1���@���ɘa>�t�/3�ܢ.���id���g�: �Eed���ڌ�U���؎e�SO�|׼���,����_���i����Gh>y�C�v
9��Kd�A��w�e��A�)��9g�6@�}�����_.{~첩��eܻ�Щ�W�~}��E��9�{��O���dq�z^���娳�ri_>��I�w;xa�����9��z-ܗ�lYɚf�č�h���(��V�Me̓��#�Xr v(�S���1�@c�S�ɀ�5��-�眫����;�j9��Z �b��`p�Fs�_��'C4�E�c.sv4���T�N�y��.�: �1�_%�.�^�.�F�����>.��9H�(R��A+�y����@����|�I��e�����'�^ʣ��7lP�L�����v�|A�"�U��o��B��c+�����oU����ǖ��͒�W-��\"`�+�сI�uٸ��=0���d4���q��O[�ۙc��	<�	�Y�\)�a�M���سW���M��~ ��
�Q�ݴ��G�:���]�t��s��y����=�/7�0�����գ���sk��0�z"��<-i�*��l�T�� �5	2t������{���`�?�cI���#z�"z|�I�I?�����8.$�l�!�]ǖC5����1�;��اi����<{ѩ&�(8�"���<�]�vڇ.
��o��Sv��n��{��FjlC�L���G'~zFm�ۚED"�"|��~Oے�/���8��9 �jxzԋ��7����-Q��b;�pL&Ť�K�=�遪���n�58"d�L��lt��ʡ)y^x��'���(=�;�ai�xՉq� gDw�l�I�_��a�vB���l���i�wx�s���<,|6��#,W�� �	(��I�Hc\[r��|��F������b����0�������\`�h��:.�ޛ�4{^�Y���ʖ;���WN)�~)]�o=��;���caԠ��_�v�%��q��QvEp��\O������'-������W�r���&(�3(�GNr[m��z��s^�)�~���4"L���n��	���J��M#5<ʕT{���ď�>�u��W�[K>*�R�6�O(�"�� Js�J���F8����(�I�ֿd.7�Sz�[�����Q�Yߜ4��^�?8��a�L������n:��֯������?��������?e<"�գt{�ee�]������n0��y8�"j�.6ч������_v>t��S����q�'�}�:l�Vpl����~���>�n:��4]�� �El��.3�a �SG���V\���YJJB>���y��A�� �x(ۋu���1^���H=���<��	P�D��]e�䶹\��Cw�a���ɱ<���Qlp����Q�S�������8�).�\��A���o����,�n^F^�~�<#�N��8��c�<����.��驄��N�b��I��`��؉
||@W�ŧ��'��Ϧwʻa#�ЏB���	|jr�����<1��-����ގ��i*��!����[���:z8֋ʎ�'�E>�)���f�����T7:��hɮ�ovDx������;���N'����m�m�"����2=Ld���Z�L�<�m�J@�B���ǽ��?�]�-n��Dy��fE�EW�Y�}��dꕲ�pzS����Ճ�����x���������h���VzJ��$7�q��,�t}�L8w�������9t�u�Օ3T��F�!�);Īܚn=Qp�4��E�{��)	�nrz�n2�&*�"�zߤ��l�X� BFsO��I�$�Ni"DۨhO���Ɯ���v!�&�q��x(`��v߮qpjӉ (ܛ��je�ñ0<c��e��3�՚��f�\�0c	�Ap�߮��O��ډEip�U�y�
��>�����@"�-9�|\\�[�%&N(C�0朖֍G�Z���01M�z�@��9��Y�o���H~��3d�Aԏ8mG��?�-�P��#�i����cK"��I�4ϟG�mV��Ͷ��9v(�Uu�h{�}�>�X�,W�#��h�(%�8�*\�����`��Op^�[���lugߺ#�*N��7�ަ�1ep0����v��'plj�7��eFᡙi���0���O�#g�������ݣ �
6N�:R�f�-�n�5R�-V�AsD9�|h�S���heD?�8�?ˇx�+2�|����/��~\ݥ�����<�L��>!w��)k�jW�R_���E_]�H�.�P���(�����-�e����L��"+�i�7E�N�A�;%���77<�%��g����1'���|'��0\ݠXѨHB����O�y���������y6?����l^X�}�[hM�#��vרI���m���?�L��ׂ�6�C�|p�x�7	tV�o�_����Л��)xo���&��\Ou|��"P�a�h��L�\����tO�6m;�'��b��Z] }7��"$�W`���҄�7��9�>�V�o1Z, w�Z�i�?��~������1�v�A�^�L�U�����~m0z�fr�HvD��6H<��2i���>~t/�����}=*�egB�1�N�ҎFٶ���")���.��M�FI��$��0��Iw�g�]u�\���WvK.e)^���+��������SSuX���T#����F8� �>���R�X�\DO��{eL���G��'�ߌ�����x��8r�� �%�"���0Rez�"���n+\�����i��^�X#xi^�j�|��s��	:"�Ϭ�٦��h�%zKf%���f����{���X�䤭�dz=2�w눜���qe}�9��E�dyu�{葐�$9*���u_ �$E�.��W܉ђcGku�3�#�<~<��Fo�.7��Dp�4�*.C`�~���p�]V�ě�x���a9m89^<ẗ́S�~hG�H��H��Gm���dn�(G��;Ğ4���},���;&�z��!�����s?���V�]<�����S�%e?D0p�Ap��"¡���D7�H�6p�JL��<�H�&��J�|d'���Uo��8�4z@Yu>|�:(�+y -��x&f� �a�Cc�8U�o�J���W�ۅ0H�wgF��8c��uGނP�2}��l[�L�ܰ�>���-E#�xı��)U�cx�3��W�b�{1�V���5��/V@�x"h	Y�0���������Hm���2'ɍ��v�&������.=��'H1T-���S�N����(K��~r�S�mOyNǛ�'6��v�U��l���oj�L���y��f�y��Y�^�6�J�g\��hO��鐑C�ٖ@�`i$W����9�~$dL:�ٻc���s�o�C�M�@���/�
��H��	��gs��f� ߰�F �)�(���j�N?f�)r��;"(I�suV.l��u�C���%��b�·���:?B�-�]�>����8�]��C�u��F,-V����ω��9�r�`�� 4ǫ�����mF�$�{ba{�:��dyU����臘����wQp�ֵD���N����й3;v�T�"�,����8g�aҖT>A`�;G���S�+�p�b���:�����u٢Bޱ4d�єb�G��1�	[ODu
dv���������@zJ��}�`ޟ��"���|�
��G���8���Y"��/��TJ��8���?N��|1Ŏs
[(Z�VW�[ݴ�95dO,��P���X���-{e�^ѹ�ʧ�I�:�rk��|+S��0$�V������T'ƣ9)��G��>0.���H^K��_�g>�gv��Yv����#ŏ��� F�
,�0MqZ���T���.ek�ӣ�skǶ�b E@��-lGX18�@�8��a�G���+�:��{ԨA�HR0�v�f� ���yԁ��Y�:��Q�m��mま����܁��;�������)uD}�rG>,T��Ϸg9]�#���5�4l.��u�3����B�k�q�����ng�[���8Oʵ�*��
��Cv,L��E�jZ���Yצ��v�E���`�+�5�G�p�xEA_��q��\��Z��]0K3�m���, �c��m�|��p	��k���/ ����p݅��:H��3���5�B�*A�,<� �W�� #�`�Ĳ�
3Ǎ���1�f.����o�ӑ+X�{���9��~�ΜֱP㚥�h��%�?)�hV[4�@;�ݝ��q��~�C �p�&Ŕ< ����
%�-G�A�xT�A5K��G�B?tw�{	E)XX�$3q�B��'"j���0 ��A�R�@L5KaP��S���X�f��*�9Q_z��e�X���E�:P]�;�iV�s����ٓ�-��:�v�b�/b���D����}��t-������,�=�֏�מ�]Е��SV��|����9��)�a�*#�0
%I�D�cg�U��*��P�fKϯs3��
�'���V�YI�;EL�,A_�
���NJJZ�#�М:����O�#�8�o�ڱ�FMq�յ�O<Pآ��|ԣ��'��e�f���Új�S��s��'E1�4zw]u��k�w��0y�#\�C-.������>������^���ql� r��Ae�}�>ߊq���QW�,�F��q���+>�j�[��P���{W�}:^���=���>v�q)����l�.��:��q�1���r��՝�?��r�˥F�D�t���|�����(��7�U���=���#/#�YB %2J�a��J0���&���P]3���*��Q�.K�`�Ѩ{?���/�v�+��h����+�_�|ͼsT!t(��`�g�%=���#�׆8�����h�Vӧ+͋n�T���)��?Y����,K���J?Q^��1継$�NC��
B�_�/c�@�L�,���U�s׀�l߬��Y����c��Cq%�c�2�E�=��]	,j�$kl�l�A���Z�8���`4��M���b�dB[�6�R�:�X*�s��t�MؗBs��]����߫��R��Q�������MK:�h��:�E�.-`�ޏi��mS���)��hn�/��?���r�uk��H�+Ɛ�_,j/L?ѫ�ٙ{���1����z ��EDzqk�<vJĵc�Κ�OQPL{��4����r7�ި#��x�S#	�N�˙�ts>R�0td��wWa�s��	>aHna�pі|g��,�bN=���F�1U��-��Z9̿JA�W��!h�~�zyd�D����)�p��O�u(~P���6o�H������U���cIt/��++	��B&���c�U�i�.�:�T�s6=��D�����1�I���2c��'�;������|3��A���a�Xh|�#
�_	W!ЊvO����Ϗ�\����s=�բ��\�.�Z�GR��=,�x�"�[bAUUٲy��mB��fi��n���n��[H0IXc��oی�ۮ�Q(��;�ܒ�5�l܀�66Vi���`#~��]̀�R`�dI��U	>��k��%!��Y2~!`�J��{�H���q�
3�O
�o�sE_�i�ə*�Up?��*�1+��c���/{�������+�F ��I��>���~߬yZ�o�mJ�o߾uEw�1dE�#�EV�	��Hs���cε�cOݕ�oKN�#W�xE�1�q<q�H�D���8���^Z�����v�
滖��l�`�i���� r]jR,�	Zf����d֔�}�k���q,+#�3�`X,��L�P00����|�����=q<�,^���(����g5������8\z���5J�����&�1s_b���x)Ih�mj_F�Hz��ɕ4NeEsr�zz���\`�PqC��
��ͽ9d� \=ZQ���!Ú�����(v@d�|��,]��C��*���w`�m�J�J4�l���)CW�:�q�b���%���Zmoz`t���m�N�}3��f<R�]�V�+c9�KF�m�b)��W�yк��<G�@���"�ֶ�S:�^�:lS)��}�������}{γ?�t�q}�=�����JW�@�`j�l��
���<�?�{3qv�����j����Gҗz��A�PG��v���]ՃxU����n�Ab�3]{�v��W{�S��N��A��~O�#�Xn0 �D>�|t�:��0Fo��jT&}_ms=N�xw�����Zg9�� (�oMe�k�TY���n!�Q��HÎ�:����k!�:>9�MʇEd��@2�]:N9@��gl��(�r�^y�y���C�v�`�k0\N��(B���A{�,��*1�v�EW`�2nŗq.��0��^ɗ��Z�
M�$�0�����e�T��&�}	�:��x�}Y'�Y����L���o�>�L��b��aM��l3���]���
�#�3���� IĬn������ظ7G�?%U��tH�x�^7`��)��7
ݯ���
Џ��ų5+r�%��O���Bt�_����<D�?7ڠ�Hf5\G+���y[�6�M����)t����_�`B({(Ew�	hѶ���c��zb��;LU�bg��y��k[(^-J�+%�x�)��}��2�#�8��\��"���E�Q� ��<�U��ADFgkge��.R��"�U�i��-��&?��h�]B���|/�ᣗ���]���.��g�"��A���z!�Q9�����<�>ҵ���(a��k5��́!�a��Imq���2�+�2��`0�rht�>�������h�>�}L_�A,ZG��]�?a�����~s@���Ou�ЎU0��+s��n�[��ޮr����lwP��c����qŎY�>s����F����7t�b��X�iT���l�DB��3�Mo5��:|_̎أ��D�c�0�Xdѣx��C\�a+3�V��>&��j�l�5����E.���+�o�gn�5꓌����R��$|Br�����7c�4�+G���Y�v�cg���M�"aЉ�;-g
�����i���q�!���n赮5գ�)){�k��|�Tuz���{1H�R"���!ט!$l1/�$��"7c�����j#1�P'�r��0�o�ɚ�8��K041U�JrB�;��W�f�Ӯީ~\a4� �F�N���;@���빡:��&��m�,jR�%�Є����0���O��FS��1<�'ed:C;�������;��L=�Ȍ��ɯ�r�~W �cLD����`de�ر2�H���5%u�k�O�]��OJ�{��鐹E�y�:�%���2E�)�?�7{���S��90�Żձ��߼�x��ʪ�, ;�¿�B&��� �Y���|�J52,�{C��U��$���]�4/x�����o���o/�rPِ�e�p�O,М�n*ϗ�4��Q��%�,ͼ�j_�������UX�:��i���b:�����T�R��sT�X@�PzX����o�a����G����U]17��W�]&�݊;�g���u�M�S���?�����~�V.����,��.}���+.�|��w=�^��O�T�!��W�۞��+�Љ��sI�nQz����� �r�B��Hf���B��AEjR���Fʊ���P��x�r��Y�1��N�R�|�+�:� U�	��V|ˊ�Yq��9z53pqK�I��V���]��D���BX3�J�yr�_�ԃ�e�������TrȎ9�Ǽ�C�ޏ��zD�B��]o��[��0����n<��
�m��j�Ӈ�_�B�+�k'�iVX3/��X�w��6��w�(2+w@#.�����:�F4�e�\	���u�Ssb��	�U	�\ş?M�l�E,�*��~�?'S���{?g�}� �����r{��G�ʝҬy����������xe��Q%a&9��~��U��Da�g�t	�V#s(C�$�
vM.8�v3�l��B��`��TE��� ���V�fg�A.h�i�յf'�jt�!ש�X��BuҼ�z�U�n�*%��!�'�"�؎�I$Aw\��%{�V��K�|�=˙�g�k�-E����Lpվ�M����^W:�fu��]U'��m ��i'�3��f=��+B�1M�.��Ij��L+�b�8Vo~ŮUM�r�`h��a&7s)�,�Vէɒ
�Jr(����P�2��[씉V?��~�Λ9f��B ��!BC2��*�@ɚ����w�1�Ԅ�����!.�v+�w嗈4�g���X2j�/��[W�v'�W�����|~��°Y,h4�-)�;�ߊ9#����ϡ�捌��>J���G7J /��+�s�_'̠��=�z�Θ��ɗiJ��]V��IPm�/곥ώ��T��EX��QZ<�\��N�H+N�:7t��&t�G T��;ÛF�4�L�_r늝v��f>E�;Zﾩ{X��h=^}]!,�,�2��o������~�a^Jqg������Ja�e�������4�����9�_" �M��9�L%��J�s���O����e�],2� {��_���%��'_���Ţ2��mc� ��m����WC)��v�u��d&B�;�jg�3|��\�>�?�AQ��y��S3O8r�(��{�G��L`��b��t�W�4r��o���d�w��(Nb�뤑�'r�CV�LSt�T�Z��ˏ��u�X��]�д.x��u3�Rυ����][>��_�Z-�(�V���� �nP�5���+��U��뙰O���H�VO�4��Av��)�
���^���g$K�������+A'�S/}���^�:�^�Y�|ًP�M1˛�woܠ��*g����/j�Ӄ%\�t�D�4�JF异']S�;�[S���#��(V��r�ƻ�%����+f��?�8-�pb��iN�����C��
�ݙ�Z6\���C�V0&0D�����������϶{�r�S3��羉0����T@�0<_���ǯ������s^�FL|x���o�{�h�甩���3�Gi�CE?3.�(ŪS�Q�_�x��Bê~���i[�.�j),������.LV�5�cz( �m����*ꬫ���𥚒������r�S$���ST���O~��Z�\��17f�����W��ԫ=\�CI�eD�Ðm/�B�>��+shѮ���N�Rs}���tV�A����(/&�;Oܛ��H����M�����G64�͢�5����_�0.b���ds�fW��/�����xb'�^�_�@*G*	z~�.
� �T�����3b;I��(O��x|�z���K{f0�k��"�]��o��_M�"�9�T���H�xF+���j�����Ղ34��Î.��
��^�#�EyD]*�ܰ����qei�s��2��1��|�
f�'h�X�-���*P<몬NK���R��u�܄p4
��q����,��������e����<�Wd���~����#n��bNL�1~f9.w�9�>
�w%zv�h���qw��˕���Q�zC�&-[~n��R���������2��o��<��Ls,ɜ\��(�xwq�.��:�'խ�(jӻĂ��i<��V�R��a��Ǝ�°�)ٯ:�[T�Ɨ���ϞO�򉵢Fj�u$j��Jj�f)ycm���|�,���ub�RN�1�꫷���︄�Csf�Cm^ ��Sz�\�$^b����k@f� ��!�Y#��D�;�Rz�v��t��S�?�uy��g�NR�Y\~/݌[��o�A��r�C�Y'��aמ�. M�dQ!�>B�ٹ��ǳn�X��/�α�6Ъ�<���p��i�&��-+��Y'���� 5��*�T`�ڠvs��d�t��zZ�& ���L����Y�
)�y�@�-X6u������{� ,�5;ET��rT��Uf�����Lf���R6A�J/
0=vWOz8�ƛ�j���ԭ��lI����۱������!Ⱥ{���=�d��s�J�	3)�c�+8@�{�'~��	������x<��<]H�a,�)��J�8�En|�l�T���>�R]��|+�ʐ_}���[𼎒$�����f�^�EWht�|�]L�o��i;f��_g�ȵ�2�oL��}�� )1&<�CKfrZ��n��)�9a\�~~W��-\%��g��� i̧bt��3N�u�Oʢ��nx;9�",�)��<�C)��9������K�����}�b�J
_/d�2����O�r�cL��>�������͚{�����o>n���͂��j:�v>&������W�9V�ne�����8�N0+aѰ�)�GWI���}����M�*~�dY��I����.�|�?���vx?�:N�ʎ��}�ͳ��(�ݣ��qY�d�1XE�5��j��#�۴�cU��,��%o�\�	}��B���}��3)��,V�X�g�䣏]����?�X%Vt��>J<C���A2��u��vc��9"!7��_�7f�r`����G{;:���M�������~���'�Шj�P��������T_IIuy0���e}s����-��>������e_�UH<��b��n����A��m�����걁�18�r���B5��6�r�X� �up�a���f�^�5X�ny���ͫ�Y����]r�g�<E���i�$��O�sZ��P�7o�pH��Jg��w�-WM9��Y:/�0 1�������Z��PA���f�����Lպj�J}�ۖ�0@��=S3�R�׆IX��r��b{g^0���I������Au�6w/0��l��?싊��y�az͜*m�:M�
��!��m>V��U�Lj�LU�8�p/Z�3�����	�O:�bQ��O��� �q�E�P�9\��xdz&�iy��*�ݧ�	.�҂��:�`%�?|��j�ґ��e��`3�o�'|Gb� �6�����5���/���� =-�ݴ-��x�:�o;O�zA����c���|�]���X��L�A����������X��򇏞��ǳ����6��(Z�� ��eZb�b�yX����y[��8�=�$���#L�+9�/ԍ;r��r��(6�)s_������ʽhu�+$�v-�1ZQ�g���6��>�{s6��B�n>yz��/u�y�c�����K���o���8��eNh�Zy�s�F�Y�o��	�Lf��J�)7�^HA�t�<��	�c�����U��/�$|i��T�F��c�?Þ;L��5�l��v�#I�����w�XiU�ֹSJ��|"
�k�>�w�Y�$������Y�Zzֲ��À�cZ��:���-1�v?��w��Ў���� ����Er��� ->�d]�f�WlU�_�~��k���\5�m��[�$҄4��P$���W�NE�M$f���Ex�� ���{t_9�|V͗���{teP?�u��p��y.��^�hI�| ����*<�i�%�V��%-�$�P=�W�����CWȍ	���Ӽ�t,�h�=��ȸ�i�:��1��nƱF�Dj j�/�s��e㶕�����[6�[�?QV+��r:ؑ|-��c�C��.��d�Y����%wwk=c���\c��T��x^���}�q����#j҃B��7�;v�t2>bqTश��H[�6��lJ�k�Y�-�Qg #�T����)@I��4?`=�O�����	g� @�l8=O˴��� Q���Cr�P��/������]�%�iB7��`w,��q�U{0��
���ʜ�f�Q���Y�{��6Z$P���AYإĜ��2�@�S $�&��ck�E#�aT�%0�֕;~�Ύ�!Lt ���ص}ϴ'�c,�QY?(@�#ş� �@��\�>6�v�Pq���o��$��D�N2ʳ ��v����է�x��T�u�|Y����K������ғ�9�iN1F��Z�z,�Ў�r6������A;��P�m���~yJ	h�k5
п�������}�!��
Uz�� k�G� /�\$��9yȫ���+1�x���]�:���>#~;�M%�s�gQ[��,�-��.���q!�϶�� H���Ͼ�ls���_-����L�=2f_=Ɨxa4/V�}	��8:X��<wڛ���`��?��b����>����-r.��ߟ�⫅�m���G_�w�ΣE�kml���]�yo;��jf�Q��nq��p�m^ �9h�[�l�0�C�^!���ڿJ�u�<����=;�o|���IWC~�܎鿕��̧��1�:�������ł[�sO��c=�Gmsh��@9�=�c��PI�	�[Z�����X/ޓeǂN��˟B߸D�e�3���ؙl�:��k��`�ǱW��1�{?"\�;C?���D��%hL-�v���
 Ojp��9Vބ25�@���/�ZI��2�6�9�`e�1�]�*�g��sl_[�p���j8<�����L�*E�n┇�U��G�3__4�~پ�r�۟v�g��˓�_��xk�hm����$�l����XWT��2ͳ/O/~w�9�HS�`��  ��C�Lg����:�����>���i��	���;X��.�Q�'�i��Rw�6E�@�:n��FK�(dO�����O<4��ܥS`h���r݊	����jZ����b��J�)δ�#�% �V�j����EptJ�HM:k7wl�t}'�	���:���?�������As���/&�nJ�;�ШqE�!���BvL1��	�8�U_��ɴ��.9�ܜ.�v̅�X��֓=*7���7�h��|�S�]�T�T�Q�Ȓ���lLa&��iIژ���-�5�Q���I�tB��̆L�}���i�۠$mwX�T3R6���4´-My�q��T�Q�<&�}Ǡ�:�!��P8��N&�1.[�<Ż5�i�ig�Q@�C_L����ۏ�� 4ЏF���ę�����uC_��^�(h�v�5��!
> 	D�91��m\�����Wa}Z�j�y/�NîN�����<{�̡��N��s�7�k����^���%T-��r���H�b�+�n��{�Q/�ߓ��>�O_}�t"�>А?�����[����B�GyS���ó�\���b�KkuG� ��n
��K���p�8���o�K}5��%h:y�e	��?5���9߼?�<P�4����cO��������W���0��\�Q���^�"�����t�>1�ɓ��u�N��r�#���M��Z�]�$0Jډ^��S��N�G�0E�SH�,�:M�EU��P~�ɻ�>�����'Koy�%�j�l�_h2��FQ��!���5Q��ܢ�c���	,C �TW�[�+���fz�]b�Q�h�MFn{�;dH�"��c�����\W4�Z��?�V{DL��K2�z�pӗ�U�e�b�f�}�k���##�$����Q:Wv
FT�q��wQ#�c�*�F�z+̨���gQ�v�������}l�6��*���}��W�~|�["c5߱�������x�Y�<��}��$o��>�z�J�1>�m[�N������ܣ\�����,��9�ЪnQ��ו0�'��ku}�4v��ā�jD�����~i�0�-d�U8Y�к����8)z���ڵF_��ع(>�L0,@�ǅ�@7?y�NU9�45�Z����Q��:�4"V��� �M�z|��&�4^�W�㮑���Ķ���w�U��s�s�z7�f���U��2����ۤͶ|��΂'�����e��4�0U���SV�lf�V��;������\�A]�y�c~/�-*`~Y�af����y�,��PT�05�Lk׶���鳷��sz�1����6�x���b`����2CB��2�P�D@��({h$�؂fPG�(O6(Q�k�bg	42P
�DW�HH�~ v�9m��;�1B
�7�\J�#��������A�}��/� ���.ut�2��kE,��ԍ�X������Z���')vl|7;�:����#��Rs�sN����f�hԚ����u�:�1ޯ���;X��[�>mGtWR���Q�ZU�c�Z\9ˊ_�P�;.�y�y����z �de�$�@u���T�@O������U�7e� c���ᅣ�rƕ2������ߓ�zSy���1��f��6-�ʏf��8h��!����x�������H����<��@3&��o�)Q���L~��\��Q;������I��9&�� c�o</�[IL�л%h։0�$��:����C��KY�|���`��S�m�L�B,�k;L.���~���bx$��q���� �D�����AP_�p�jA���2���ܟ^璺����-Nm��=��穦�Ò�^7���OD���/���B)��f�����Kԡ�4>�u�iT��cs�M�Xm�3�����⽪���[!��%6����Ɏ=��0�H��3\r�x�� ތ���B��-�̧PeΕ�f0x�X�U	�H�XuLK�g>m#?x���V�w��|�];_����ۻM߰`��v�#��s����b#0xx,�����b���oN<?_?��+��oRi��X�x/b�w���c��cQ�YJ��Q�����YAT</�~�J��ȼ������Pƿ�.XB'Q���i�^��q=B���[�2'�f`��9OK��!ԙ�ﻙ��*-�i�ޭr��I)�C��Yi8�U�m���BJ mF�ӄ�S팷[��kv^$!O,�g�THh��֜���<r��! a�4D�t\���5���p� �cH�� LУ��j'��d7M�a ��T8=���\c����Q���\��x����
�VR� �RXUx:��yGX�D٨#��V1h?,w���1�aJ��,g�z��m#03���q캶��P���h���u;b悵]�ypf|�)��܍��=4w	� �{����`�9e�c��D�ܗD������ȶ���x@��W�B
3��0����Y�lڼ���G�$xծ�B�]I�}���f@��c(?)�I�Ǩ8��\�J�+���Y�[Dw�j+�n��u� T�􅰁�<H���?�(wٞ�z)\�ɯ�, ��/�ײ�S�d8&p)o�^�]��L��H�M���kG�ڑ�GC0MqS.�N>��}���>kq%C_2bk���T� ㌯v���o� v��$��ɞ؀��!$4����
�Y��F��0��2��
f�/�I�E�g<��' O�`�����*�9PhnA�g+�?B-���r�c���kR
m�{lI�c�������a��.: �p@�H
(�G�����p�y���Q?_Vz{�Wn%�	#
�U�\�f9k���	�,�g��k�����9�y�ˋe��@F�zs�פ؉sEQ�%�F>�,(E�:����$ￂuU!�����;]���� b��ʂjJq�6��*����y��c�m�y����I�P騦����Ly�0���ߛR��w�GL�z"_Թ汦2�RH��_�������q~ d�S����y���Ɩ�A���U5q� J�~(�#Ҽ��f�1�<��l�8�o�����C�M���<L%x��j葮��uf=T���|���˩¤u\�3�P�4���	R�HD?m��Z�Zj�h�y���F���젨���#�La@Q[�X�S)<�iX��+��f�,��!�υG>�B�"�/�[�q&p#��+�
ES���2p%�	1s0��-�Z�F��w]����R�l�'E	T~ޞY�o#��+�u!a,vY�W��_�0�Z!0��#�\ �,�IAX3�Dd��8�S2]O�&�����l>��#�]6]|�H�e^?�I���R=�IT%"����#��J�u�5ϥDWC��u����D��.��٢_��df|���|W��B�����>7k�7Ӝ͕T�wI���]@��G�J��v?�}�o���`��x��ҳBx��c Bl?üÁ@y��@e��I��g|��[���g藾S��NS����BqKW�������N������񆳲����ic..��z/��`.E�aeӣh��oe����<��S���������R��I���a`�r'-�0ߍ��&W��j8���l�,؟K]���[$YT�)���ԕ���;����ԣ�Z��N~=�����2,�/bȅq2� ���C���ʟ|C�k��
�	ug��s�<:5�~�3�m��R��LG,Z�����<>�7GcLR���dz&�yr}Wo8J���u��NϹ/
0a+Vv���{no�9mYD�tnY�V��7�~i�\촂$a�z^�[6k�G�K�����t�����.���?z��/���}���LX�І�9>oN)�~,5�}u%M���һG�jk�[;��䳟��~�;P�R�w$��C7ΆIVL�ʋ�t�^ �_0Ej�Aи��r7�����=ʛ�����=󕢳L�K@Ew�\LM��4�_��M�4!�k��¯lX�|����#@	y�X|R��颖�H�g�]���xh����+wв�SC��5�.Z�ewpSL�]��3�� (���U�#Ou���f�7*v�yFL4�Kt�?�g"
9ڭ�J��1+Y.�-~����Ѕ�Z���A��ͽ��Ǣ�u�R�09�iA�<��M����7�2 <N�(�򸡽�PoP��#��פ��|�P]���A�1^��CM��2%�����駂�fY�xĔ ����a~;�]� ��:ӱ�P-z��a%��e�o���]�禖0�-)Sr��V�X�cy�-�Xp�Y��Ymiޏ���m�)��-���Z���mP��tK��S��EP�Z�\� H̵ͯ���;^�6oEw�>>>���&��Z�n�`	>w���#x0�!�%�3�;���p^���`,�\��x�T@;�5�V"i4!��tCڧ*������(���h������ܸXz���TCǵ�1X�$�9(�e�����?�~��W%m�<�w�7�M����'�a~��rs>���'p���yo5,E&~+��7�<�r
�c��.�NA�.��}}L7����,ϝ��/+�~�ʧ�)j8��5=�Q9�`����#o�u�^�}`�D�bT� o~���Lm�x�D��:��Λ<��uʴ�E%�ܪ>慎��SO{����F�My�u�R��!��U~f����ךm�{߳�9\�<W�цM6m��&�9@���Xި�#/�6��²�D?m�g�������l�����e��ś��>�2�`I�񗆙�wEN�|�^�@b�v�����kU�O9o���ؚ)��sY��;����f�Ԡ�w_������;Ќ#)6�:V�xW��{�ں{c��a���^ȉ����_L��q9�F�e]w�cǅ�2�.D*���N��%� ��Oe��Ҽ��ӿ�1P��u͟jE¯׭�K5�B�]��X�Q�ա��ק|}V�������"#��6�h	�����|�}�_�_@�+>��"��1g�jrJO��X
O��ϋͩ��g���
���N�g�F:bΤ]���:_0/��ˢ~OQWH�w�-z�����뤠��@��L�hP�8n6�`�+�n�+E������g'�wH9uլ4Ժᨗ�E���b��B��"���<:Z���ImX�/���bi��粗��� '�*�ۇ{zV��~�c���y�1,��ݜX0�a&e���ʫ%��T��םhJ�e�\�	�:���X�g�=�7)�[�غ}|s�{��_���sD�F�?�(�{c�Z��� �Ǝ�4B+��;R� ���7�^I:'��I�#g�LX� �q!1(�t����!�tu��7AGX4�#��ۓi_��b�%�x�����o��"9"�CX)��s�7�r�=ܣ&�?Bz��Z�O5o˦���ވ�-ʬ+�G,���D�n��1��Or1�!?c�^��9������*��v|��8Z��XZ[W�z��N�"�6�f�R"?�3M
ɲ!)��)b��a����*����F,�������X�U�"��C�����\= �����ūn�m���L�:��5x%����q��y�[M�[߷�^4�7��9�����U�{�㘮��8R,���V�|��C�.��X���eN�P��-\���Q�o�.�kQ���9K��iJ��XN�J zl���GV�h�Z������=�|�ջF6�}n0�V��B�[����cz���ƥc{�xW�џ�~k�SqF��y���6�����&k<���9��|���u�$	('��;"V���,�!��f�B0f��%�s}�&�|(������]O"0XŴ�vdu�ͰK��u�WyO�='��L���P`�����/�}]��땫j��3j�Ė��V��� ��v�ڂ��-� �"�&�1�J��1Ǆ�E�Kk�8�Y�V��X���;<�x,��i���_����
������A��*$��yL��8`6�b��#���1P�>u�m�|��L?��x�`�q��U�Ж�oQ�Dp���wm7#�J��X+k�>7L��Re^V��HA4�F)"_.�y�g�Hm;R�@|��=AI��EM�¯�?Z�Ȟw�B��}ꭶ�>h��%ʚۂ�%������=�����iկe�J�v�]r]Ʋj�4/��XtՉX��Ɋ��?�h���U]�RJY��}]�ߤXv������gs x2:o��i9�%�(Fi4-��p������S1'�D�������qY&ڟM���YS�@�
�@7��d���B�[�HY`�6w��Nw~v�G�a5 ��@KMn��a�"�h��Gc*��չ��le�2�x��/�h�c�+$�N�1�=�bP(p�B`��1/.&�U5쎀T��4��]��a���ͮ�����
�sƄ�b+�Z�s�����\YAk�	X�7��v~��f��T�9/û5�`1�NJ���V� �\���:V��湬�9�L"9m���:��q����l)n�Ul���ś��!~�I��D�gsK7�B�Վx�HV3�c�Qlp���5��H�_˸K�2��G���?�zse���T�~[��5ؘ��ֈ�ߑ~�* ��͚�	�7�:q-m,��b��t�|��{���U��u�tc�cx{���-�Jb̤�i�����Ay�����g��.���57gѱ�),��b꧵ل�R�j���x�*g�@B�ݮ(�Q�"���1;�����)��_*$�4�<�j�s��Do��q�i��>�.�P��1��
%"� oE�v��-�5	�3�P���	
�Iy�ghc�1�`	Dy�c��I��-�u�_���Gم�F�k�>1ɿH��g�=��xm)s#�#|�V�&' e�Dv�x};=���b�ReL��>g��]I��,�eֶ���pI0�?LEw����S���|e%Ϛ�v��C;2[�ځ���i������)�X�T��wJ~���<H�X�V�DIs������ �6��#��-����b��/����'�Ѻ8"�dO@����R�E��~���"	}~J��)�ttѠd��r|[^S�Q����N%�B(��l븡ʒ�V�:^�b�Ws��X���<�_[*o�����a++�N�����&��q�"�K{����������4�?��@fI�+Ǥ?��JI��B���
?V��v����X��l�\�Ц<�7������3T����H3=*4�l�9���I�ۀsj�G#�Ge��TT��k���'J�_�0�yh�8?��qV��]Ps]�G���W�y�mS��$����4�ݬnұ�-ɰl)��a��&мxke}����V�e�)���B���J��͗	���k��]�����Z멖nP���h�./Hu&�js�9>ҊΉj�2���򰚜��sLrd�d����D=#�0����P�t��Jr��k����Lky�M�Ld��X����{X^>����[���,b��~+�����3m�E�R�bǯf��xl�ڝ)��q�cӏ�o�X�����(�c��QY�~���6�;Xs���*a�YJ�ܽ��f��W��<�����Q�+��SI�s(:���Kc�P�#������.�d�E㜻�_���B��_��ӕ�5|ڣ���:?��Q̕��:#R����9nj���ύ%�d�a�X�@�ϛ�(P�b�b�S�N�Z/60����l0t1z�:T;~�p:lK3��_8��F�[�`�8���[��8�"��Q��6PQ�������� ����������6qʴM�JXY�0Y�钊Jr!Ӊ���cU����vgvK�B���\	�-ϻ��7�y�8����#C���~�:�(M]o���>(v����7�εq�C���q����e�	.xv̢޹�Wx��_�D���`�J���h!����[1=�������D���yngտ�r������lǲX����wq�ei���V;��ό��t6����!3G~mbN �#-�A��
��OAB(��U>(wPo���3�r�Ě��F�2��W�3>C�9�C�>ɠ5}�%� Z!�E�B��*�]� �[?n~������K�@�~v`A�J�ݏW�f���h��&w�L��w
���k�9�
�WbE�G}C9��)�R��@����h)��YD��o�O��A�#��J�!D�;�S�!,ʸ�'�TU��(�gޙ7����>TK��U0���m/�{��oE�C�,��2�»��� Z4B�N^x�e4R���ט��m���?k	V�]�
=4��\Qz�TF�"�P�>�1��"�}�uڹ�E�Iw�)O��|�;:���66('Z�>@�I`�^�k�����ߕ��ð�4߁Ib3����WjqE�â�n���Z�/���t%����?�}|�M��op|��ߖ�~���'��=ſc������� �2��� x�k����PL =V�*@��ٱ&{�'��F��G�`e�:�-����jzw���+o�N*��G�f,u�c�E�\�+���U�����l��ª�����[��`���\D�&Ԕ>{8O��2Y!iY��|����7LȖ�}�� Og������!�s,�*=�f�(ם�c_G�1Fl�úV�mxVLle�H4�*��j>6J��{�����nsq�1�@!*�ј�S��;ȡ��B���6��~��A�3����/aK��R�p�XN�?�J?�Kn���Z��P��c��}Q6�����kTI@_ 5���- ����_�3>UBib�b�ߥ�ee x�N��-`�[�D���Z�Ŝ;�[�����&��

��,���O�f��}s�[�@�WoWC�v||��'U�� M��i~IR��]��wE�"��I%��Ք$^�e�Ӽ��ϥ���L��5�l�칗�&��l���#���-� ,D�K�hR�(��g�.�/ʋF������������?��q��QG�BD�#���v����i�|�8��y�ORZ$|��d�p�\~Y�E\M�2��w~�"zn�!��,���s��KG��W��l���L�>���^����D�J��DY>+���V�o͕q��W�٪��s�T�7N׬d��>w�z��n>��߯�M�c>o�6�P��gYM4��ː=�@ͳ� �͍�\" �6��T>�U||=���hCUl���� ey�"��LI���}�k�;Xw��[(�՝�Η���=~���;��)kl�~ʶ�Zo!�(N�<��|���k�9��U�+v�y����V^Sa����������qY�C{�7v���nF�J(�D����$�sÕ�F��Q.����'�v��~��?�T	vD7e���;�؃�\K<��4HuxOd������($����ڝ5��^�=�/��X��MOK�4`ScV��i���ktHZnE���v���P숤�azD���� ���3v�E\��)�_�Y���'P`f�c�c�K,�L�s_e�@t�o��c�,H���Z"���*�6�ڝ�N��μ�Pf�ZCA˼C��?�z��p�8�r R�s��ǂ�wN�φ`����u=��tR�5i�1��K,%���	:����h�+������c���pQ#j��.�*�N�[[��;�O�������(wj �=����?#�C�*�}�A��
'���xp��������~�Ji��zAZ??�3=$<]s�nʲB�'���m¸�ݨ,�
�'�<T+d���q��Rg�I ݾ���1%>��qɾ�]2晿���X@��;��;��'�`Jt�MR�]�,����f��Z�:�>;��͚��+���ʖ�r��ϡ��>�9�	��ۊ��l�'�[[�X����j,%0�Lˑ_���Uz��&�rא��ҡ���rҶÂ�KM�Z��I��1k�X�ͤL�=�j�.&eB�˒����mj��'C�22��d�[c�Y|^�{�t\@�=|L|ȧ�QفF�)��9�fj/�c���{t�y�6\��<,Д�T���IQ���-��U���V^���vI��7�n^��y�]u\-�fS�����Xw��1]۞}T���ؔHM)�>?�}3L��ӂ��������V��OHkٖ6��~��̣��y�]�tj���5VtL�����V�K}�1�E��*i�,t=�k�N/�E�\�`�2�避��9*@*6���a��ߞdB��C#J�(Z[!p ��:��a��$ֈ,�L�"�L/s���1Gjt�ԁ׏��N�/4� Ԯ\t�%!�Dt�"+	�LM�;X��HKJ���J¹�z�W�Ff=5/��-��t<W����Q|���$65]��ڗJxM�5<���U6�	�1������Do-�����v͐��O�e��,du�Ț,�z�[�Y��	Ë҅���,T������\�u=G���������4?���P6�u��a ��e�Hi�}w�(��9�n6��W��0�zqZ�	�i�T�8��Tǻ�E�Bg�M�ÀT����V������2�c����Ы�]<��֝~��w�����.A�;ߢ����Q)��P���o���4����Bg�**�N
I;���<���<u*��3?��f`q� �3�m�߉�<���G,�R��v�V������w|���\\j�`�l�G�:<���_���-Q��/��;p����g����#@��D7�9��}�P�;�YȎ��G�+���,����}u*�Y*�vw�:���i�"�m�CZ�ۏ�?�C�e{��:��qZ��7������M|�8S0`� ݨUyؔ�:G��1f����:T���u�K��;��(Ȼ(�NNe,`㽊M��JH��p*�r��-�S#��_��ݔ����¹�bq�ñ�Q�ܝ�+v.�Kխu$0Z+ G{��"b%_?m�b�=�w�`\����7�w�����Z;�լ%�#����{�n1e�މ������n�s�S�A�2��ͺ����{�&�=Pw� �$�97���:&���)v����R�y�Z�Ez��(qPI�)�B�B��"l��ڒ��6�M���v�p�b� vA74�;�;#��E���y_���������h��̻@y�`2W��Z��Bt迾�Ba�N����,�28J���5�C���[馕X��ߡ����uA�8��o��	���9�m2w��G�z�w^q��ުD���zɶ ��a��|��|V���p4�1 aZ�a��.l�ܦTb\�zp�a�Ҟߖ�M*�*�cP�( �-�mG���n����BIb�m����T��S7w�i����J�q��Qw���o��>Ԝ�����,��YC��H�"����%�׳m�~t��$ÑX����]�ߖ^������A�M�O�����g�̞~>aJ�f��@��
}������ru~�Nh�^��;�9��.O�n.�<�o�N�nVpm����e���x����ѭ[A��g_��b��E�d�O�V�Yz���M������g�:n!Z��4�Ŕ������D����K᳦��8���������e���~�b�ZݝGs?�����x������ca�g<�rN:��+MH�\Y��w���Y,���}�~��˪G��\��l�,1�F3P����'P�5U�H������u�/)��x����yQ�n��nau<��?]1��nѡ���c+�F��s�Fhu-��8�u{u���wR������}�����~p���b�S�_kJ�p���j�5��kG���/Y���ar3�eZ��o��G��Ҵ�
�qN�K3T�ӰF����tX`�P�KS�����oxW����cYn�Ԍ�ש'���ʰف��wZp�<��;xZ��x׎9'�Č��r�6���-vNw.~�\"� <#anY��'d{�ae������o��OcV� =����T+S��FX�M���03{A_R(k&��$�tiܯ�l��O�2�gТ��p�\	K��>I�y�;	����H�c)��99�[i���C�������P��lV"Uo�L"c�����n�4����8��	g�ĵ%A�[����9i���⬼�4~&�Q�:RzVi��T�O-s}���@eT�5�K?G:�^v�.�Es2,vj
�{v�A��nQl���/��Ԃ�vg������wH���ͯ��Yk(L��~��f=*����-���-<?l�-wa�N�p�(
����]��M?Γd?Ȓ�\�0M�Ǻ��2�S��Nx��z�L(�|��?64|��/7�p��~�5+�'>�mXt�b����|mw�\�y	�!"��Nb�+����&�f�
��c>�5�/��ܨ�jК��E�*>ٲ8)6x���Sh�a@��O�������oJQ����=��ZE�K�Ut(xT_j�[��ҍ�������_���&W��PJ���[/��p]}1F2W,����Ҝ�Iz��2���������3��W¥Q66�������g�����r�W��hs��ŎE�kV78�P�1w(�G�E4�#5�D;���~g�n�5:kXfNe�\�������~1a�pDS��ͮ�Tiة���ߛ����������zC���o:����."�ꦚF��ԏ��h���ؤ���V�G���q�eے�)C�/Ej┿�����h.�ց9��Nӟ�Bl8��j݆���f�����A�dm���3�Fy!G�?������;`G�L��֢}�9�\��J�EqM	�S=s����VdZ�5>��i��˼�芸NU�����D��]_=b�S����M�Ǔp��|�*3����iz�+�dZ\�Ҡ�3(c��:t���6Ga��B ��B�.ǻ�h�")~��QZhP�c�ឃ@/aI�^W��ؓ��0B=��gmx����M��f �}ӷ*����Z�cR�>+e����FM�K�D��Z�����O(��M(�	iiѳ�2E^ɱXp�����^����֠gf}a���\V���n��mi�YjD?m;HX��h0Zp�2���Z�_k���ȭ,��n��=��֝<�n�<�rQ�j7G~��U?�L��3�>܋�e��#�M��BĞ��^nR?��[���ϭ(�UI�e,��	�PԠ�ch�ݹ�z��,�:��˕��y��.�N�.o$�aZW��@n�=����:;��Jʆ��a:'��w��>���Sxf��Y�,��nJ�8���?�h(�<%N]�C1����VdD5i��R�{[����9�����Z��:v#�j����
~�ʎvt�}y�OAU�ڢ��"��o�����%�L��%�wn|"����ń�o�6�l��|/�_��UI|r��}|�+������W�*��~8$^�$�Q���*��	P���΋�%ƒs}��k��+�b�G�F��,+���Tj�4�xJД��]�3�hSY�!�P�w�"M�ed��};�4c��GB�f�;N�񲩩�S�Eom�֧ۢ]<_K(l6��٬m:7w�������A�ϔ�=���&�S��I��6��i�1w���(��O:�0m�FD�1�T��"��Jp���͑���\��]�ڎf]��6��������!��fJ4�U�j�f%wE3�����T����R�HkT<����Oh�!{�~�Kw�[�P�<Cp>r�d<Z�<��D�4ZݰQ�t<�9��"�uo.g��y��L��"o�3�>�珗�}b��gw�@hd�±��PyR�[z�;H���T�4^g��9fq��x+ӄpK�̪���w}=JT��Z��|�@��zq�%���f���؆X�����nV�D�U����>O�VӀ��/"	�m�5� ]�)�;����ʔ4��suF-լ�r�r]cA����	.(D�@j,�k0d�ߦ�X�S v	9��6 �}�q��w�Q��zo��%�93���?J�p�NS�E�r�E.X��Y�������}(��X�?ٟ	���L@��{TiZs͜�[.�t��Yb���;[�X3���B�U?�|�[�t�>���¶ɼ@6j��`��QZ�eu�}�`��Zf�Q&z�d�������kߚ#�f��w�?z~}ǭ`�^ev���X�Q35.�3�s>��0���x��P�/��q�Qĕ.kzh���ƊݹZ�����)92�D���޲r���-���!,\�cu��	��v�jvw�1wV��IJ���p���jδ��mٻ����|�Xg<����r�#VMO+��۽���ڻ�d	%�0���]Q�t|c�R�w޷����zt�xb�+�����ex�E�B���kz>�K19��!=�3}dԡ�S�ݫ�.1�{(s�����Ł�����ԫ>��(/��vkz �`���2e��L<��t��,r�����(?��i3T/�s��X�U�x��=��`�?�o��<%�h�����' ���P��5U�(��Fa�i���X��b�3���8�U����V��?48^v��]�eȧI� D�:u���9��*=��C|ޟ|�G�������Ax;6�1֍��������o����|�������?���hVAu�{�a�i��vO(5}�%^��:t{�V;�|�Hc���X��T5쩿U�49����hlt.��p9I��K[�v�j���Y���"�G/��m�ׄ�^e6Z�BY��i���;R)E�ꢟ�2Oa�++#8� �r�K0�8J l!xV�f�u��'�:w0^�
B�����N���v�[L-�bċ�ݿ#/ΗS/c�d\uςP֋N o��o;�<^L���Q���j������פ��K2u�Z�D����A��2�O�M��)�҇���v���0iw0d��j�q�6�P��>W�!'1!zrL��.��g����^�]<�V��6�ΰr��kռ���ݱ>�ˋ3?GzJH�)�q�ͥU���r%�ֹn��ҭ������B5%��)��o���;� ��6�,s�[��zhe�w�y<����GF�K3i�0��
��������g/�;���E�@?�F�ĸ�`\���:�Od�1(h��;W&���ۈ��0EZ�1_�3�t�Vk�>,���C�Ww�����RA̿�^�g�"�jl�Cȗ��2�z�Rxl0\��h�<��)�*�����G_���� 6{����!��e�'��Vt�?M1'M�u�N�;6�j�?��վ�¾�Λ��L�i0��d}Ω,h*<��O���v�ur�jEG�bA]�fʤ|��I��lO��]���Vh(�Z��ǘIY��|�wl�����j/y]e�߬��8��h��:�&��|}(�gl�i>�N��|�h C�� �U�Wu	�[)�J�g����e(��*�Cl�i����E�E�&C���ԫ��`��{ �y���Zq��;�<Aq�Eq?�o~ʂ���ȿ���h�$BP��,�����!���ƛ�GM﫼���#�}>ۺ�[?�m|���-)�?U�@�^ݒ�8�#&����^�Qy8�#R>s]��:~�`P긅j�#��9p¾zb�f�ڜ6�Rѱ\m�d*�~U�U�Ս��b����o��ì����b��ۿ�L��7�b��I~����'~�x�cǙU��ƎC �X��qm�C̹p��vo?�Ԥh�j���Q�r*\���5n+-6%�h
�.vDow�QG����7_S��S{�H0�L���i��0{�+ۙ
�7.rk.| Q����[�����B�o���Ӂe�?�����|J��B���@��ʂ�?���?�)C2�^K�*̀c(J?
/N5���:��賈od�1��Z9M8 �4
�B��yDT�/>nlE����x�h�D�	f�����R�8�]�!�]a"1O�g0|nZ���v�:�V���p����h�4m���]����|��[LJ�ˬ;��esA�#@XA��;�
�ڕC�t,s�6������Kn��>>���p����G/��Ǿ�Bb��{E�~�F���SFU谦�C�󇸞�!�������:�F��Z���b�Z���̪��u��g�^u�~}.LŻ��g_�H\^ j���gy#�`�tՊ�� �;��M�=v�^��X�R_���B��駫d}Z��P�"\Z�L%Y�0��@�����}�"����taP9v��w��,*��e}}�I�s���9 ��|�c ��b�uZ��k3�����I�P���K�Vu�Z��L�[		/�;���ߘzS}s�>o|x��6�"b������Z" ��'9�˴P󤶼�\�s]Q���\��
��]�)"U�p�0nfG���a���83����N�����|��P��5m����R ���-嫛�͈z��5��_�r���,`�	�ϝKRf��j��I�ݱ����[k��~n��ѿ�xWkf��u��ǛE����{�����ccL�Q��&�;��ѵ�ZdW�t!BہS��u����[�j����1���:Ɏw%�+�iί���?��;�r��%"*��dxa�ܴVL���<����մk����.j�]�ج5�����YYx��[��	�̘�;,\���FR�ʨ<�� 3�Ҳ$ ^/�{f�?!lv�״ktD8Y۝":I�H���v�e��@���CXg� �:��*q=�w����6��g������,��JZ��35�`mgL<���P�"�>�נ�>z"�Y��_���~������.<)��4��0Ё@�t4��;��;d�5��������P�w�J6��|8ߝ�a�pҹEǦ��BC2k�#խGx�)�hʛ'h�0�zk�o�u��2��s�a!?�9tQ�g��J��w�D�Н���G/�j<��h]�;���O	.J���q�_^��K��Ǆ�j�q�w%U��R��q�%{��<�`a^���}>U�-������P��NkwO���*S��;�+PH�5�L�l@�x����+�ґ���2�ESΧ�9�%���nނ����I��+Z"!s%���0��p��Z,j'�T�qߜ}0�`!�����l�|�k��E�x$�;��Ez�s�F�ҥ�)��mZ��zD�������0Su�Nb!@t���>���oN���6�6Mt�^�J�?[���k���9��u���x��p��R �c�RO�K�í|�_^�@ ����;����G�<7�Ҫ��d���@.E�E�xS�獿��W��_I���MIs����p'���CZ_�ou��~q2�a|ޤ�:ICq�i��� C�H�]�6��H'=TQ�xx��q�n�`�U|%={҃ H*���YVR殆q��B����XS�Vh��G�W�M�c���n���W�?��G� Q�@�����g��}n��JW�x{�Azm���ho�F3�f�{��Zf�X,zk�k8*�J�W� G�F�`.��g%�K�5-
�����'���o�B ���Ð�S"QO��݀{𓬝q��$��͎�_�Yvܯ.{ ����V��3}^���c>	4��5�ηk}gY�~:�92ݧ�yH���>I�z}��a���rcASJ�pv�LI0m>(G�:�q���?J�F2�l`�� ��}]�΢fp�9����j�ʞ4E��-�|�\.t��߿˿���U�������E	���&л��*Pgw�g}�Y�����;�,}��(9,R�Þ�g�mWÏ��z>E���sٵ���0~�"��q�jq���uE��f>�?�ԯ����W�'��3h	����\�B�"�"�Бj�}��U����
�F�C#����*�	M��&�]~�)ث��,�VӽE��y\ F�Y�ckAd�wR> y�KX��9�Ei��C��?��_�7^�t�h(dMd�9/���\ �Wba��i�q�z�A��~��qyT�ԯ�<x�_��&VP�12��"Z\����/I
�23[N�[��g!Y	R,���?��F�.���!��K�HU�cC���Z�ҁ�q��X"�2Ȑ�ۗM1��x�*�/��52`�km�1$��+Cej4����̿�!i%��$.��yb�n�㏈L�,�r�|�^`)R�'���jW�O\��~��E7�`����>Dǹ����X����������e�;����J��#M�7z��`�^���1�E�Ƒ���ݕ:�ѸZ�ӝ��iY�Q}�\�w$�*,�9_�g�O*u����$A��
EXS�H8��?��<T��b'3�L��ņ¿�"Ǧ	G�\*���N��q���"��$C���?�����t��uW�O��S��h�Q_ �a���A?�{;��y"D+���Wj~"�P\�� X,���Sߑ�&+y�����ѿgB�� �1Z�*���&.(���ڊ�/$�����EɰL�ϊ��u�	$l�pg[߭J����u���H5f��Ҝ/��+R��Si�Ou����Q}��#����G1[��P5��U�D7%..���,1^�Ϭ�Щ�_��}���]��w=�iº�i<��ሯ)cJ��S}W���w���oͷ;",=�?���ބ?�?�~@Vi�yZ$1y(7�A<�3��_������S����L���uz���]�]#|����[)6���e�]Gn�7��B��W�}�ȴ'I�+�����1�\��%a�t<��h���O��1�y'�E�=�`�5YG���'�d�b4����:t�A���"�!�^
�e��:[U�L��yY��yp����s�˄?f������ձ��ڶ��5}�:��6T7`h�]�����a�1a��{��~"�����-���'��EY<�/��:S�g��'��m�z�WW�u�q搐�	�[�t�*����н���I�>��1Z�d�7��a�#��U�R�[�3��������낻���T.�/�t��m~w�iڽ�M�S�F7�dܫ+4hK�^�[��믿�߳v�>}n�>ls��C����q���w=�m2,j�׀$b�G�����8�,9i�h����};G��;6��%8�� �����W�:|������\
.�u�������~��g����(C��Nآ>ᢐc��2�&�/�L@�W���?���;�db�]��KA3��v)Ky�ύW�3Vg����	�Z}���0��X�ߙdhV�W�i��G�����{�&�""Hz��5�'����@U��[��܉�BF5�+�O%b��F%�~=�H�<���\|�WhW���ȳ�:�NM����lG����?̂��1��L�x�l����@Ӆ-�;���=W��u�5$Q�uzf]�f��b�膣14����G����Eϱ_�2�	X.��cR�'`1��ˣ"4$T,�����;<R�|@��m��1���o��?����o.1	�h����c�K���G�����lQYV�&��;���l+Xu^�v ����B�.j��}��|��f�5�W����#<�L��,G�\�Y;��5�r)GŘ{�hm �AeM��q�?8��5�ى��3���"@����S�a"u�
�x��p�}���Z��Z�J&EW\GՉ2��п'B�Lh.)@#��4�����5H>���VGn�액�G���"�5�{�C�y3��q���|����-;�/��J:�����%6��j�u^���%8���Ju�:H�W��N;ϫ1(إ�|�)Zn��Ǻyt��u�xE�%�c�~�M-3�H�z_���q�<�M�fW��X��g<F௾���:m�AJYW=..�6X$O��=K�*m��'�h
������e|Z��	����Z	����Sfo��o{��}kG��7y�r�R�?m�����W}*�ik��l���aD0��*�@tC���d�1���r�h��_��
���ơ�M�J�`+�O0v�(�e��9�dx�����5g�/s��ϻ�_mH���~KWd��8�(~�K#���Wc{w~� !Z{G6�	:Q�L֞�4A���'?u����b�Ίk�C�AQ����%��L/A���΅�!a���~g>���7&��J��x���R _�NX-��7+�8zv0����!B����ƨڳ��|~�Z�{��Ĵz�{@����u?Y�z���5�5�Ξ1C��q�v�~B�����'\�R�S"�)���:�vY���������;��:��3��hG�a��/�^-��hO���yt笠�#w!��=,y�,x��d���]�Y�_wɮ���g��D4�&��K>?����;@����]����|�|�ٞ����@VD��Ʃ���ra:<��.�O��B�#��U!�OC�jt���fa�%@:�m�P@�Eˉ3�Z�f�P���n����b��y�h��o����	)2�`�;d��R.V��V8�����*+���t~�����G�ʿ �c�Rǫ-&��f��d",4�ɾ���q�c��?���E��(:�����"�C��Ub�o�A���}\3C~�4��[kK���y��ͥ���?�F��f]��e��ށ!!X���漂�/
>j�Y�g�_�7�'M���0����iX�1�IB���f�ԧr�o影҄c�ث=�����!�j�3���H��@;
;��T.c���9��>'���}��X�1_!�����&�D-�z�-�� ���	�:6V��ˮ�ky�ul�UഓSƹc�*b=E�O�s�z���,*��y`I�|�Q�l����l���X�S�z���fF���T��?z��F�G�^LXU��0�U~��9���7�U�Dڮ�g40O�X��3X��9�{Y�s�����a��w�ߖ'�����?*Y�L��X�UH�i�G㫕=�<�W�R�_���O�-hm��O�]��A�ir�m��w3k=��;� `:*��b���8��3)��;eL(����_0��7��m-�m�.>�.x+gC;x�L~%��Z�8.�����\��Bys��y�]z��`�Fz�n�\�У���J��H�Y8&��p�r>b�`n�j��O28J/pB�Zx^�y3/�Y9��r^֨X;g�+��Z�9h
ͫ��2O.g�����O	 5T�_Z`κ~�.��F�U@��;C
3�V��u�f}Ѩ.ff�@���E׺[�[-]6=��@��n�;"���W��Քڏ�}���~zP� s�)�H
N�5r��رEғc��R�%���Ԡ��u7��4\�浻���αo��6i�ٳ�C&��ݵ{?�՟l"��@�.��0����p�_��3��@N[x����`Xs��yPa�
t�<����Y&6���m7�{� ��*��cѱ|��tE�喎s���}���jZW?+$�:��V�FR�픡�H���ǲn5)�P�c�_���+�93��!M�,i�7Q�}��G
-��*&'�����#����HSQ�C�VGyy�<�+৭_MرB.2�0-�'oR���Ul2 ,�|�~,.N;L�<N4�)�cP'��D��ŽO�9Ir�D�P������D������̪������ݙ>v��L[��q�C��tV7�����M����~$-U�ČZK���A��	Jى�X� ���/��y_}W�2��]4��,��Z6`�p��|�1��|�+\ϓW�
�f}B���fe��2��
�$΄���v����Γ��U$l�|z4��,�[�8�z~z?�b��r��u��8pH ;y�%��b�X���k��*� �S�:+nX
(p]��-:Ӣ�O[�����%�R���K$^�Wl�K�>v�=E.x )p�iz[g*.,��j!��)�SR8��ͫe��fb�I��o�o��\?zR2"]����*l��b4��{=alF���R�_�_�먄C���܌che�b ���P�� Sa�xc!po̛��ʠ�IlJ�VqŻ"�����X��_����zk����S��S5��rF��S�;fty�&}���|�̠�i���@>\�q����[R�F�����ʎXb@��vNd-t�ߣ��Ɏ��X�̧����NG{f�/�-�u��~&��3P�Vi��!�.�����5�H�L!��9(U�kN�eI�8�s�6Ҟ�П׾���xI:�ܕ�����Pۺ�?6��CM�Z�@˟I��'��� ��8S#��V&�=�;%��-m��cޤ�t9ry�Y���ҷ���;�ƭ(,#��5AՏkx(�-߯�M�P�[=�g}6��*��� vd�ν<�k*�X=�\���B7ӂ�6�tHC��뾐w
˔�ys*�.���ޅ��-)��'�&rَ��O6�Hu?e\q�e�쾆f�����+r�5I�>���T�S�͖����σ����n\8��cb�D�lDJ�� �4HD.0ň�ۡcL��X���G�n�+�B�v��0�k�:Q����`<w�_��pdm��ԫ��E�.WT|��`=��p�DGiLY�����J���-W��!z��@�(Xa�O�|��,�e�=a�ڄ�O	�v�d�4=�����&~��&����u~��w��M(\�y7xMQ%�h/�W�7�X�|�t��Q`@I���X�6�z�*��M��Ӹ֕��0�u;�ږ����b�c�/}_b�|�|��ǚo�i��$���|����o���A->dw�
�D���I��Q>gR&�).���o9jv��3���s��v$���q��*IS�GM��
�ڢ4Sd�.�8PV�36���)9�o�6u�e�r�����'�AҎp�J��1��=`���5�J
�Wo�Xy��"�Z��b��vֺ���*k��Wӗ``�|���;N����an|w#�e�#̵�!#�(��F����>�o�s�����9Pn=�c�E�԰�ū����eU�-��z.%���/y�"�������y����ⵥ[oTk����fC��P!�$K9�,�!9�q�>��ȶ[�Zd��D0�Z���,XH�hrkG�[��7�����#X�0���c.��G��T��+t�.�=�O:-���/���y�?S���+G;�ZW3��y�Z=˵��+��۲��9���4Go�K�x�	�o�B;{}T,�����8��	n!��-���)�r��@���f�﫦��Z��~,�͞�g%��"@���`r)�h��n�*�	wU��~�����hs-�w�p��(!���^��9�fF~]��`�8�j������CR�Q3���e�ϥ���pR��hwL�Ҵ��]��nSJP�]�F���쓭��oM��T�۞�����'�cB3��]��pɑ r�Լv~ZfV�0�-_r�<|}N�C]���d�=��đ�hg,�����A��Uc,w^R�7���ή��gV���WtT(g��� �{:_CԄ$��|,�#&�.$�o�#��<�P1֛Z��<�
������R��v6�I���O�(&�`��3�J���Ӻg��t���۠3��Б!�`�ؔ� F8�6�%�=�\nR)l��t���o������cl<��<)	?��/NZ�m·Km�D�n�Wx�0A��G[�;5k��̷�'�"/+ƌOD	C�Α��l�:��:�Ŋn�[�A6�rP��;�G�{��Ȗ�MώAN'��`�Ǐ�O�a���j�ڀ	���]�zׄ��k��R0D%WČ���v]V�-J�~���6�m���C~�?�ն��{\�y�=�������0fT͋ҁZ��{�2eak=���<z��ͮ�FZ����P��+�ܒ$��^--tZ�ӆۼ%��Q(w������L�WOecT\}R4�E@\�!���O�ڜ����:덒ɣ *��<����s}��n���ܸ�[���(�U�y�ֳ����#M�$�@�7�,�k���>�n;k-� ��#�uUNoN����&3�e�
�|wY��('��CϪgeKN�A��� �ީ����YI��FƓ�(e �`��#(hG8��a4�Z�:��܁o3�nJZOWܱ�[3���:O֝��lq �eNg�L�GfЩV?�ʫJ�R�`e݌0�I^���2y�D�h��J��=lӆ$m��
)�_	�%?ՏQ1;<*�J��q�\H���j��������0�K�#�֨d��}���V0.��|��1~�N[IB��d��?�23��=��(��-u-��m��EJ�ZD�)��ս���<�T��1zx{
��*�+��ǫ����Y�dk�9�s ���	�X^�rG���	0̨[j㽞y�.�g���f�b'?G��.�o����9�w����ew�&�C{6�#�D^�M(Ə�Mvtsj1D�"o�V|ҭ��'}{���7����Q���x�6�VڞS����nY��R�9�R�HLlIDaPS�Z{�W/\�ko�����n7>�����	�z���*L�=����K\���k�]g�^��i��;�(��1�8f���ǝ�ŵ��*�Z�{�l�Lr�U
�:6O�)�x���g��
�Q��9�0�Vp����)�e��ʌ�yg�.����N�@W�|��9��"R��~��"%�N�c�<�q.&%��'_��s���ˡ�O�Ժ4�~��D��IJ�?`b��;��Id�4�����*�ߡ1ŋ�)�}sd����
��%ON=����<r���}3�Dh�n�GzK�؍u>�G$J�c��(HLN�*�̪\x����J�5��4r4,�D�G(*����'L	�J�؞8�VӤ{��*�o�0̣��ZmM��J`)D���V����X>ͻ�:)����7�򑹝t���>�.y��Fj��ʧ������\� C��8{+1Ϥ���	|Տ]�)"k`�9e�y����ʝ��Wf�VBw��X�b��e�����zap4<�bQ"K���9�����M��Jì��*�X9��o7ius��T��V����Ɇ��8�rg�#��/��\�Ö�ɟ�&V�c�;U�~zt&���p�7'�kk_�va�M��&L��8��$��Y�$A�a2q�n ��Ǆ�0�㢋&J���(��D�B4���� ����k\%����t��s�/�&ĩ��_�L5P`=YQ�z`�f����aT}�D��+�q	�zojzv��1�����S�� ���9u�b�������<3{~k$bE��u�3�WU(����v�j�t
"��bl%��A z��סW�j�oc���#���T�:qhr	
P��=xd����(0�;���钁� =��N 9,�()�e����Cݏe�(�U�����RXo�) ���dW�����l"�}h������l�͸=G���(֕�4��0V���mА=�N�5uN�����6�	*/��ۓs�L#�s��dG2.��b��K�V�G��2I¶�<�q܉�K:�M:M�|������$�_��ƽw�='���z~���Y0���`Sf���P��#�;��Y�ޕ�=�a�8Q{��s�aN%�û������ZG�va���Ë�����%5#d-Y����"?q�)���&Tɓ������ѫ�$�]��Π���5X~��#9�&V��A�3_�Γɉ���p3S����~ek���UCݳ�.)3�\4'a!�+3�^��b����!���YǬLj���z��KVV��E�TR�`�@�@�M�8��J?�fH�S��B̗t�[ӵ�;�����a\u�(z����+̕�_[��8ե��ʓ�ª*�))e��I^}%���.�0�O0>�!=- �»I$\9��p��2
8�V3�8ik�:J_��\�e�,D�0��1������N�I�ᝢ������������>Z1�X=��(��~=郰�i�j�����'��I�m��Y�چ�A@��U}#�jw%7ܹ���F�@S�o�T�G��%�ا&�e�C�Doq%��3f
<�E$Y���u�����$�m�� ��w
׵;�9�o��삳*�ӇK�g��%	C�_
E�a쫵��� ϒaУV�s�$������������~y"V�����) Н*ǳ۬�QG��?���s�aKÊ�)�d��REQ8�?�1/��Ә���q$+��Ԩ�C�>��,��`
)*w`���R�̃�s����A� ���j�����C�Os��+��&�mƀѷbY�O|F��	m�il���'��M,�~N�_@�����~��\�:�,��|>���s&��TF�#�_�ר�9㊸��y�:����$=�#1�$��x%ڔ����[A�
�ўT|w_x��� ��x��{߹l�e�KIo��[A���I��u����/Ȧ��b�}�4P2%��r���z���ؽz���^9����`�J1+�!6M��r��i�?�����۰=W��~�y�fO���U_	/ӵ�m�.zo��u�����������R� "Z��\|4��I��n4�5x�f�q�|���L�s���T���[#nŉ���5X����E���?
��t:G�ϟ���Yr��٫����0-�`���8�)���S-u)��<A��N�<���i{\p^���i�̡'�v'���$�cl�ʛq������Hx�|ԩ�P��9�����:�C�4TQ�E#Y
Q0�a�ʘneN��Ɏ��j�a��������wew��}\��Ik@u7�E;킡�~y��AMJmV���@��e yY&){��* �A�Nr�`g�IF�SnA�7G�04�����X���@���z~�A�%�)�_�2l����UJF�1'?g�=P�bd�S�=Ԧ�}��/��f��m���~���x�F�mV����+Ǘ?"@rG�����K�6弎�8��wד��&�2�<OR��
W�7`�lʝ�~|9�����N��E��Wj5\o�۟e�l���n���>v�URU!�l�NYt0l̖�a-�}`�R��P�(gTѣ;L� [�c�j�0�N�m���g���(R�$͊���|��\1D���q�X��»z�^LF��]�3G�`���i+���D��됝??=q��ġ�3�yxX Rn�ã�`:�3e�:WSpMb�#�s�Kqhە�5��A{!?����~�R��ELkw�gc�����kf����yY1�����0�C�Y曘�Ӝ*e�����Ͱ�Jj�3A}�pB)7J�(T�Z*�!�F

-I�Yp�g��e�Eq��F*y9�&�a��ٙټ����o��3��׌t�\Y/B�QF�����
B�ek��~���ͦ�%;	_U��۩��Ov^���N��7�\���*���q@;�W�hn�`�4 %��*(}tC(`������L�jVы��`������N񁸖Y��^g�6Χ�w�L��� pN$E)w�%�����W�$q�"��%g��w�
�u��|���`�)�Τ�x��7}�򅎔͉�P.�cH'�XS��xG��h�h`5R��ϕ�FK�c!�%��W���mJ]/���|����8�oP�4���6:�y�,yzL���:�zeeӸ��;�v�H��!+�l��(F��f@O�d�R��d������Z���c�:��Mk�@ �9�A����J6_�E$�Q�� *u�f�Zع����Bi6A�ȱ��䴦��Z��9��I
�b��Qk��9�|n|�(i�)ޞ˱�ICyD���6yh�]}�$�C+��, ��2y��oP��HB:�B��`��N��QK ��,V2=D�RE�*
�� ��S���48����ɛLc).�9��Ԓf�(��:�)��L�q8��J����(���49p
�6��5�TS�IB�3h�Z��X*)v������H[���ǯ�x�5���E��l�_�զ��LQ^>��n�ߒR2}E�;�W�G��3<>��|:Ӯk���i��B94���+ʱ�y���.4em�aS.���a�6�?TJʎ�m0�u�2ڿ�k�WY̬D����V}=a�޿L2�j癣�y��0*�!���G�c�1a�~������V�%a��
�˺~�xD��i��!�'�����Q�a���e(qw�pV��h���7��Rg"^O<$o�<2���f��4f�d�u���������2��]��X��wh��L�x�)����W2v��c�,�����Qc�Si��O��`�_�z�Z"=0	�������K�طO7�a��MR$�@�
̝<1�F��#x�ȉu�p�π�c������ѽ��ET��m0A�c�S�� *����$��M��Е;^��J7*�k;u��U*���ݷ��[s�T �k�@0m��G����o�Լ�z�Jݯo�p��
ܶ���#/�I��������]D�/Zf����à�]1g��o.3Ɩ9#{.d�1}+�D��#!>��DW�C�GIÈo. kEh�N�@T�Y�Ѱp>,VG�~`�)��J��t.,&�)d"�Ґ�����j
p��X� [A��		[�pb�q35��W��n�?h�0��ć��*���Ҏ�<�쮥���Ì�{�A���o�B {?����D��zl��pB@��I0�:{?T��1
�}��M�����8��AX^�>xK�765���-��R��,V���^g���C7v4���A~��z/*^o��ʇR6!^gcƄX}�h�Ϝ�(~��Ù�}9��r�l�$�p�~�ܠM�̗���Y�T�|EOV� p���� �U0�`~�V�AC��Y�6�s�r�c����\K��}&^�j	�l�DJ�+)�rЌY�G�>��z�j�D>�r��_i�{x��7ZQ����A�������{Z]���NM��Ul-4p��!ȉ��$�n;�F^ l�@$	�J���߫����S1�D�]����x�)w�M*dwM�XHt�c����F����8{���ML3���^Wx1#_���Cu�RR8<����׺U������3P!;��P�q��g!��@"��Uő��u6���v�6�f��-쭽�I������6����N#���4dM�����D��FR�$r��AǳR9�GC(3���7T+kr;8���D�9���?Q��.:�D��l��F��#�-�U�1�� ��\�]�!aP����df�d]�Bičk6ia�{ǓU����F��c�j4�&�����o��QO�]�p����9�a��GIn��,���t��H �kX�%=�k�g��[_�·A7�:k�g�Z�$���3�ޚz+�>P�K+wK��__/h�;QR6)?;�=��2�Q=Z^<*&�oGv�)reԋ�@5J��^��_E1$Ήs�e#�Ne73�̼z�3=C��Uh :�x�F�"��G�蘹[�c�3�_����V�z��W&�����#���c?�vF�����l��_�d��!ohd+�av�$ �/zS,����O���a�3'Gո]�G�5��!_E�E�{eڒ]�~x���_�x�I��Lvr0����a5��_��|O����ȁ&dP��=�\:+��(V����:P�C�oZ�B�	C��@�Q�;�^T��/�r�P*������[�b=�����h�BuJĎ�]�؋�v�g�E	�S��V[lg!*t���	U�\v��+������P���B�%W��}iZScc)Z�T]͋��WD�f�v�b���le"�<sra�w��a�#==C�&&�QA��S��\�X�d�N��!E3����)�(�T�1d厼��B�n*v�/�nj��ҦY��� ύ\�Y�(J,��qZU(w�[���A�V���ϼ�ur~�y�T/}�5��:�����z�z-��`����HY&�lA��0xs��[�J~f���=����/wP�|Q�j���O����/,�*������g��Sa'%�s��B������r-{�x>�6��w�҂(��fg'��<\�m��B�.��,J���C2ءQ�z����b���*�t�*_ǼY4S�*��Fj5�� �NIn����U�W�F�Z�M�ܹ�$N�g2pƌc�1ìB��m����qKR��=��!+���虍9�qt�I�*�{�HW02�<�6��y$G�T��#���Q�N����jh���.7�^��Rzߕ�������S����FL�	؀D��A8A�	9�Φk#9;c7�o2�>@
0M�r��50*p���"��	> ���?��ܔ��i�w�V�4�[
���21E|�a��?ĴJ�8:7�����$�/K�����_���KJ	yn19t�Xl
��d6��)/*_;��)u������S�� ��'�?s�\�r���R���?���#���^E���G� \)4���t3������KwY�q�F�f[�f�1���2q(��<�_�R�.2�����7��Y��G�y��4���[S!���:���ؚ��&��>j�y6)��.�s��+�����/�#��59��D=������DP��jm�j�GS�:=�7a���}�b�v���)���bǎn����K��S���g+��%�w�w� �!
}^��(��=�lNv�h\�x3����8��c6E�`��Hs��B��ꜙd�ٕ�1*�[��C���hX���kހɎ����Jky#![�\���mP+�B�}��i�QR>����ǎX�jpz����m���e}��է�Z/g'�gxx|G�;�_�j���Q��FJ�]w;��82��G%B�ϸek��D��s��f�O�0�Ý�Tv����&�L�r�Z]�S��Q�m"PL�?� Z���"�� �O�`��H�T��$S�ď���g��������"0�UC5_�o=�E�q�>&^�&c�R0�>i
�m�h��1'p��n ����Za����,J�	'2edW��Ol�+�7Px�B�AArL�8��3�2�������t���w}ͬԙ5�#f�5(e`�N|6�����fcw�_2����_�b��;V��}(,w��Q�i�8Y���j��s����YφcX������ �z�(k:�y���ʆ���K�X_6����Iٌ�]�(��Cxt��uV febVf�"m��P�ߙ��Z3@-��u��\�N������a��'V����ڨ5ꩼ�m~�=g5�[��8�G|Ɯ����r��J:��S��u�Ƭ��hl��u���o�w���=Ƙ֗��N#�D�GUdqJ����GZ��3��V�L���tk�r���#:QmR�V�G��	��.Dh�E�ȍ���2��r1ڤ�>c��('g��p��'˘z�Ma���)}�i�ЁZ�o�xl�V8��7X�i5�D)��;I��A�D˓�r��_R�p�a�Q�&+��.(x�׊�3{2�GRD���%�;�So����i�_<7�*�ʃ�t��iHӸ���S8ޝ��r��?���B3���Nf��Y���o-����bc���]UP(����;�Z�=���Q���^��#�g�hDY�Z���};y���z����%'%B��x�ya��I	j=7��NQ�g.ypm���T��w_n���KF�q��?U��7
}�ڥA%����_izӗ�Α
f��p����mhobFmN�TN9�����46g�&k��4��I0�,ŗ��5�%LT�\�Y�7�ϴ���ȸ����S��9?<�ٔ--�I�� ��������n2��c](O��x��f�!7����ɎA�JqȚ�(�X��
��L�=��ҞVLa��&
��k�Ʀ��&L��[�T|�ʑZB�.����&�fj�V�7�P��n9A�g�1�H�s�P���H�5� �WY�#�C[gI�@�p��~��P{o�DH%����7�ҋ��o� Y�w���c�����)�F��hu��K�8��9��Cs�r~!�����|o���<�u����~�f_��L��u��?s�s���c�Jw9ּ`�z�O���):J+e��C(��9�z�"ΛL9
W6������$;�Ȳ���wR�Y�$>i0f�yT����;�Ja�����_q�2��i3�:��RH���gc��b�vY�E�:?�>+�Ώg���$Rz\+o^Iy�gԀ�h��ߞ��4�i�(������	C�����~��O<��|����w��}Y��� cP�8�}�.���bYv�+O�MN5�خЦ�=�=��w��p�Q�n��/��y�V�=S1�V���^�(L����4�Nښ���~
��~�X���V�@�I]d���ڤB�ZHY�9�Iꯚ��NaN��N�
F�d���~�O�;��hM�h�Jvw�ձ,>�C��*����V2g>o�;;:쳀�l�{�O�.J=�r�Ȕ��H8�$>sr��|���<.�d����ʥ�zc���4�����)���y�����Ȼ��W\�%t�7�1�O:�ce�Di���!۽P~9;��F����aѹ��C�SW���j��*�=��zҽ�_9f-@�.�\>��73v�_*P�(%?�tz$����Y��*��:l���>��i�O��D�H�ն��;4�v�߄��@֭���������XK"�$�^���3��g����Naݢ��˳��͂_���aM��0��r��[���@Xs��1HF?��]�(3JDM\�I��@7���y#�{�/NNjYC���W�����T�#X�C�s�:p&��'�s�N���Ԝ.�ܜ�P�����C1(���/���۱����_񭓏!3&Yd|	򐭋q�c�(~v�(�㽴�70q����|�#X�hS?�)�2Y�5��AɻV+MKXͽ�i󭤊ץ};��ڹ-`>o��O���_�i�2��2b����_����9|YzZ��\Opy�n�5�#��Q�b�)?t��\����*�[z��Ʈ'<��f��C�D1)�#�Elw ��	��K�_�5���Ϸ���+��`�p��B׫ҚԈ�:*u����2�K��L6���F���โ���3�\�L�v�;7��h�Y8AqOClґ�I�XM� ��O��/�R�ق4����OE�M��<_I��ѵ�I!D�F��r�������OGX��Nbn�l�ZQs�����L�IzN#���(�,�^�@i(��)*j�����i��t
J�ڇ�����'I"}���x��aX��C��<ɡ����i�9m�"y	G�95�A�`!��4� ;���ZO�7�@f$,u��/�7m޽k�TP�tW�Uu���)��/�f\��=��w:���WHi�G���J��Z���>x-�2�C��Tt�l1Î�����L��<Y�2��+e�F��5׫��c�d�C�eJ�{��I,Xr�iU(A�7��^���N����~rg9�&ٍ�R�������ٳ���O�Q�(e$%N�ś���C�0���)jiұ�<D�&����V�}U��/Ԥ�&��Q�'0�9j���;�2V-pE� ���yx�����e�'�.W���+]����L���Y��y��*�ǁe���4��^�(u>�V�@-���	�?��{����m�׊�a�ά$�
�*����7��:��@MI�j��@緦�4=�R�e�Ԑԗ�5��%�$ʣ��d���܈�1q��y(���U e��@Bp>����%�8�ҫ@H͢l�Sa63����Y ���/��.ы>��#�y/fG|��P�<6=o4P�-�&c����E4��bd��֏���7�?�i1�w������f��7�� &݃�9wg�kJ�^འ@���X��ݖK!���dD���
F�9��p:�ju�|f�f��@�>�w���D۲���eX�l<�J?9�����U�R��!1DB�&[�&�Ȣ.��+@LX^P��B����l.��������I��*m�w�/q���y��	��OW�ۻ/O�L�_�Z���W�|}2��Z�P���i�8Z���R�a�Υe%M~�C��dᒭvf�,����l�]�C��+��uo!#�9[���]�{�'P�~:����8|��;�@,�;[��FT��Y�)w���\R��ǵӾpu��:Ի����ʝ�L<
�;G 
���N��hKO����i���8������gx/�x�,qZ�~�O�?�y|��9����8%���|O���6&L�+Ee�Mzz����o�bO�|V��;+�jm�`�CE�|�@�iߢO��{i�Z�~�s����w�Cb!��h&��<�Ja,�K���]3�Scx���'6_VaY@�e�eg���Y���U2Zݵ��2�r�Y-M�ݒ9<�QPqbVM�|��
;�V�(w�����-�E|DN�3���	�R'�}����)�5th�,���lz~vzJe�zD�Rl�c[(}���x��T�+M��y�[���d��mG��ą��p`��f΁9w��?���z�%˪���j�{E�P�J����PZ��;n{��"�P_��Xt�#�[����m�rJ+r�\�]�r��s)�BcG���*?��>��<�#NHX!_���3)(��V�s��Q��a؟/ʇُ�3\s�3[ܞ��(v8_$����H"> �k�$��Ό��n!�t^�~��\����hu�����[Tڃ9+���'WMj�!��Β�V��i�,�5vf�Lv�e%e\��E�	{)oF�ݧ>v*�bu\ض�n��_V�i�{<=�y���O���W���,�|&0�l�y���|� _�,�/ȟiQ��S�$��D��(8�0P�J�7����/��<��*�:T�f|�&�Q@�kuCߨs�a���bob��Y�+����0fvC�*K�Gފ��栆ɎX���<Ob����W'�&k]��e,/���Tx�F4����������,vNd�C��;�Xz �v"�R�Bd�Rƣd�?��H�J
��J�v��� ��e炗�'�8Gd@�t~��W8]Ϧȡ�5ic��^eQ�~�>�)���Y��k��r�)t�{��1G�)v���
;�m������nc Rr;��`J /;�R��jE�VB5�G�F�V��8/svvk2�2؂a�XE^�(8�����n|`v�D��c�u~qO���2���,��^�W<��k1U1��>=R�P�k2��ׯWӗS������f��~�������E�$�~��	2���C/���KͿ�K"^'�M0�����ӕhcMS������Q�(�`�@;BOF�ǳ�o.��u�f���u�v�X	�1MV������2���r�������Ta�#e�Pⵒ^ߐtx�A����ޜ�o�F`����l>�1�"Z�Ҷ�i����dK�Q��$�{�I����3��C�oOn|T��ͮ8��T��b���P���a�v������L�S���g������'�����lJ6��9x^&_~fX@�	�����/_�|���uٳMT.��K��檾�o�E.��% j�;	k��B�����p�@�+@��,��O�y�7U|l%��G��G�(<SqɁVy�y=	AT�w�T>z��=yR!����ׄ���<��:mn�5�G����J����O�Q,���#P].�lF��mA�gY s͑%��,N�����U�R)>����-���]Y�\�(��b�kK(�lْ�\�]�$&R�p1�{	��f�Arcb��!@
���h��U6����|��������>��;unhǄ�JG��0�g}Vm��Z�&����ܒp��#��@���)�㙢�L�	�?�|^p��O�_�fb����Ȳn ]CJ�Մ��ꑻ�^<�ʟ=@��XG�;�:b�B�W���)(u\y�йmEa�^��__�6�Z�p'V���b<�b���J���߈��)�k,
�����X���COוLU�ڹ��!���XM ��}�m�m��כ3io�H#��B��T�3�č �.v��Z��Fc�f�o��a�P�	�<_�1?m��O��̾�8;�u��Ǥ��HR�X���bp<���r?c��1�˖��X<�,`�����$Q9E�C����-�%ܹXW�&[2M}ʕ2�+hΞN��t;���Y��������<�V7��S�� �<I�!4@W4�#2a��#'���g��������;'2��2�D6���!�$,}��������:Ӧ֭������&`Ah��ݻ0�婵[�= n��?W�*�r}��l�)cUoC��e�SU�N���t�=�CW�m} �D�U�aQ�Nf����2[2��3�G���ulU���yB�+��
V�	�H����W;B4e���Տ��@�!7�V�x�.�?���Y���щ�(���r��.��ά�,���X�H(�xԄ�#���'�Ba��Àj�w�<�v}��~$�g�t͟3���$�,�,��2�x�G�E�|&e���9��s� ���������|�f�>7�B =�a�M�s��+�Lͮ�әL��Qò&q�8��+�ky�
%��D�X��'���>9�H�+��1��5D�E"�v\2�S�T�z�K�ag��w��8ߛ�j��Ԯ|y�vRw����ז\1�.��C�Eu��n�h�
 }��b�)΋ޮ� k3��nc���6�K&`�~���l_;�Q��%��wS���[��f�z�ӿ�l'��p�$.֦�*�.vE::�EmJgтkk�n
�L���r`oW���h�aw�T1q;>�f�=�2�Z��c��&�<����B�SL8���V�w�6�-���s#~_�^���)��_P��/蜟,=g�AJf��2(�ș�EMf���2�7q&�
�&H�t�K�7ypfޙ��J�M��=�S�A͵z��F��ͅ�"���0y}Ԣ��&�qj��G�c_a��A['�L^j"���k���%g�͔q��-#��S�}EcJ��b���c�0ﾔmV�+��C����)�޷9��l���;q�3�K�g����>?��_����7�\��d��~\��L��PC�R'fP7�s(`0-�n�=iC��م2m�+h��15C}E��)�ْ���=�j�N�!��چ��o����}2)i�%�a��X`�4����]���p�_�P�m+��ţ[&?�ꗠ�"�mh��4�Izke��`B��%��E��T ����q�aȳ�p�~YY�gu�n�nhx?�4�E�ֳ��D��*�� V�$�0�jƦ�5���S17B[Qvse�]�8�-۽�[�>!�Bw�"O��CmDa������;2�ώ��͉,L��҄���Bq;O�ʊ$V?#�c��R�(��ݱ�Y�G� ŏ<C #ӱ+;Α�yfK��/׏�xd[�_����O��rgz�<G9�4ƈE��`
=����4i؈���;Ԅ%Vy;���g���n-3��$�((���F%��KdE�A�)��HM��� �89�ѧ�Fqp�Q\lrui���וj\��>VO%[���m7Yzw�ω��oMS���7��(2�>^�uS|c'o���oG���u	s��7�1ҿn�<_�o�����K��%@�\�I�~��ZZ�]Ϻ��צTg#��'W�p���U̩��5hK�YC�����^�ŰV_,����Sws�z��~�tn���b
���.�QZ�pni���8�a��k�����FG�F��i��u+�iw\rk�Gqc������~�JQ4GN�`���}ߑ���-g�y]��l�sZ�8��N,r4m4]�b0�bu<J�0v�G�/�\^�(��P��1�!v�oJ���|̦r>���4X`��`���*�m����;j���`�a`XE�J��z]iT�S97��3��8q���ѐDfF�CkѼ�>���wr�/d�e_Kٗ1E���f&e�j;h>|��N�n�fz�\^�r�;k��#\a�_�~�������_�������X��R��w�$g1��uR�'uq���0%7g�	]=�a�B������R�-\���Ƹ����ӆF@�LI�Ȝ�B�b����G��	:�鰘>_�@����EB[�c�*I|�ى����)��xs�`y92�wy���0l�����D�)�h�k���m��Z_ޥRT������g,Df`@��Hֻ>�Y5��r���v�'�.���zGF���\�t�������̔��_��-;-	H�k#Hh�,:�芋ٔ(�X�]�H��1���$��3#���x�)+�Tq��ɠ��?���	���&��F�-葓�����!�r'4Z�-X��Ҟ�5�R�D�,ܧ�(��^�^��<{[o[�V\p�b�9,G	oJ�$ι��<z+~7E�Hr������i�%"���6ܴVPy��{	��s��GX�]�*㭸���K�ص{�o�=��0j:s �<��J,K#��:�=�/��V1���V��Z�-�K�r�XY�K-yB�nC���_��_�#$P*0�⋯(�`Z_+�9��L�p����wT�u��㨂xuq�-X�}�V�i  ��IDAT{!�7���m_/q{t[�e�d�WR�<>>����� u�HW��Æ�_f���^_�?b��("���r�C�sa���O�L����Bd9CA#�������[�YM/�����k�1k(#d�p��Y�+xk�]�m}��G�ܯ��e��*���6��6��tI`(SG=�ی�+���p�0�Yt�f��N�ű@�A�m.f�p���
_�����_����|���y�����ϟ|z�r�a�O�H�u'�@n��ڻQ�BxreD��Ť��&�+s�p�!���ݞ���f����Ca��]� Ԁ�@��I��3D�Eh��_֢�>��v��+�,OD�AE�B߀��I(w�7�+/NX}~`����k���o�P��`�<=]Z���-0V�V)%B���7��Zɯ�@ȧu.DEZ���
`��գ���ݭ13��X����t׷�T9;�Kb���l)���Bn�����Ol1��^���U�3	�PS����3�pte�'�� ��~��b����L��U��982ٝ�O+8q��Q"���צ�^��r��*�� `��t򳿈� ��`��4�o�;u�U�$k�_1;��3�`�:U]�6%&�{Z+[QX�+�+���V��R�_��~�)�W�����YB�;�!�I�/�̔�kOl(wLF�Hf]��w��Γ�K֛
�z��A+;�s6���I�O�,)x�?��Nr�FURޝ1���ew.�0N0�;B�st��\�f˝a��(ސb�p�K��y�g�&V�>���Қ,i������Q�c���<�� d������eG��a��U����3&7�����6�c�H�*���3�����ŝ�r��Zy0^���o�Eb �<]�������3|�����/�����C���>/`�yy~���=-uyd�Ԃ��(T:��;fPw#=���a7SM�Y^����D^f�`�N�Hȿ+J�6�ץ�*8
�-�!�<���P�����	��M̤W�(q���EBD�uVh���,%���[�֡����q'<x/�^D���8|A�,ׇ�����esF~���l:A�ԙ�e��w���{�PV����ۛ�%�MA��me~��|7�z�|WG� �]��N �����`�c?[��">2_Ȁ'Gd�;]�Pb���R?��Y��1�����A�`�`Rw����������1/��4b�F�Mq_��S��� ���Z�͔�ϖ�{���Q�7�Ϭ�-�M�Ѭ��hs��屵㋽ŕz�-*��a�ό��!Ň�wBWUϨ1�s�'��D?��M�R�S��E���4w�P�o�~3�|������Ȇ�Uc�V��Ո�A����ozL�Fdo�e���Ƥ�R�/�/N\.9R���=AA��Y&M�U&�19T��ʾ��Oa�p�(�=Z2k9�h�/חL,aq�L>�4�Q�9�T���w�K�c�j1�%�3{�z	���[W�	��@��V������ͽj���:aC�>�
��J�\�jj�n+-��n�c}��[!���n�CA;P:!�p�r>���������7�/\�.������r�<gb�2N�?9�Ff��`x��:�tOڃ���'�q�F��ő��F�3�j�5�)?����#�)'^O{�����8�3��5!cT;�U �L<�jq;?&��u��ȁ�iHIŌ0}ES��m�_�|w�</v/SxV ��׾2�@ل�e��S[��[�q�YC�k����њy�I��i�*�+�Qc�� �C�W@}q4�R٦�{��>��Y�|t���
ډ:W��dN��o��Bk��f:đ���.�/�fQ����S�r.{����f��V�2��+u�j�<H���gd?���C�r��3��<O;`�MED1�}s�Eg�M���ZX�B������ |��=�G�œ���6�~�T`� ��g�?�L�r��䞀/N~|܏%�7�~���~�'�����>����=�
��u��צ{�R�h[�,�g����r����^»n����$�ꚤ���<�}�
�ޓߛÒ^2��J����IQ���](�teG+!0\�ב9�tp���͓Z5:d#�@5�r4kt��/�� �+Aq������ۧA(4���ř�~g�M�¬���Y���[���0�(aԭ��s���}V�u���ޘWJ��F?���$M-�+^T����h��Y�d,�Mܭ�V����Ji��V�.]v醔'�}z~�����<�_�~���	Ο�	��G��AA�:�	8������U2y�q$�9B�d��;���oԐ��1�V9ۊ�M+3ǵ}�pp�w	�N�L�$)8�Ѿ�<����T�A1�����3���dµߝ����r���E�Kڅ]�"<�
@��2��-���Q1��2��=�-�������	`8Q������0�%�zו;ků�?BC�h�:8��h���(u�У��4��>�Fpɗ�7)|Fq<��L�O��Xyƀ]�&J�\Ď�#?csi\�T>�D
���E��9��c�XxHm����,T5ʗ�Q��Y,�A\��� 	���[�k��0pZj�M����x��rG-s���۷��K�{��C�j[^9�oLu�1��Y�h6�q�TV�*.�E��mǖvLՔN7L������wK�����M=���x_����.1��	A]���T����W�o�\�"՛�5=١ Х�kZܕ��z��X�t�Aڞ��2CH�F	9<�^�r�T	wX`�A���Of�3\ ��@�(�'�śJ݉�X�&�r�}�L3)v�|e�Ȍ���4�$��Q������w�Y�	��Oǉ�ჩ�ך��t
SV�����l�$�P��؉k1bO��m�r;gK{zx @��/�p�˵��/d��8"�??�)y�<�.���	��(��Z�d�Q��r�����R���&j�0h�V>��D�J���BG��r�[%ՎG�N��tV4]%<�."��(�D���6T��kPaC�m�/�a��dk�mŀ�wGM(����3��5�7�&�����^���B���8�^D���	n�N���2��q�x4m�U�/:�����0g�X����Z��_a��v�x_�~��bx�I�ގ�Ζ�a�)�BhMI�\9���lG��^ā���OK�O�t���~�O���ebV}Ɋ��+�]�D��Q>���&j�I&*�p����:��h,Ek��N�5h���#+/�;7��^�^ӷ�4%�D�c�����!��w�TzQom֖����:��Ij2D{���/��F��5J��I@��][KH�s�
�M����ؚ��WȔ�"�>����X!G�y�G�4'��Q��*�*u+c���:$(9���ˉ,����F��j�LG��$N���8�7?���Q���m�`S Q�k����]Y���^���pN�0������'R��Ěg��ĂB �;����>x�g%�t��&4ږ�K��˓J���������h'@� :��'�c�i"7Ȥ� @?��oiuR��Vm�x���} ��.?�A�>�3�љi{�'��)h���ĜP�Љ���q���]��b��E�)5&���44l8f���(A�m����N�C��Màu1���)�f�� [܋ʆn�����S�W�4y��)n��P�_MqN��s�S�T�vo"���!t����)�tJ�f����+��	�LJw�"�>�G^cVDSfV���R�H�S'���4ȕ��L��������=\��E-o��U���7Ngx ��|?_�t�Pyl�sa���eL���	�֌
�꾋}��Vjq��=�h�J	" wB�G��j�ڒ��PF��6Zk}�-�~�i���d ��oz�ϝ����X}v�z:��מ1�ש3=�z����U	X}	����@K���>�<���ڶ�d�$=VҦ���c�X��jYF[�Z(=�n%�G~������w������V��	m�5_|2�#�p����ѱ��Y��K�K�z����_���}���� -�����$(�6:$&�߻���L~�hmaE-�n 5QmM�
*�b���6�a���u�������
\���U�/mVE�"�:�DN^����@������'�i(:��=4����8����2&9B Q�浬8��{�L��6�� ��R~$P��$ QT%�+���'t�[I��l��g:�����F$���餳����O����vR�/t\������������_~%�kf`y�s��֎�`Z�1;w��W���y��<ɱ��"S2�Ωx�;MP*�@}��͌�g�U����-��j�@����bg�#���t�w�@�6��./��Obw6�+�F�R$7;sA$�~@"���'�be|H�r_.xB�D�� (t���-� hh�͂������Ή�vI		�x��YA�B���S���}d����'�����ˡ�x��F����;c��t�`�1E�ʭ���T}Í�{�b�����D
���(LC[��W��~d��6op�f"��h�2T�F��G�x�CuNZ�,'u*Hf�3����o��YBS(#oB��V|�;�4�ݙ�d���ɟ�9�y~��X����G��)B Gښ��B���];���IB�R�+�?��b2:��\'��!�K�zǯ;X*&�Wd%1(���7_����4���@%�T�H�%?�;I�c��$E��4��X�Ի]�^���]B�E*~�㘑&D�
��J���G�t�Gk�����'i��q
%4%oɉۺ����m�m�u���t���u����}��W���i�P�U�����y�k�,P�-�
�W�~�wk|0��"�J��~z�
�U�^?j����c�Hx�K*���N��k��U9��[K��I�;��%�$�&m
�3e��A�ќ�4�?���E<rF�%H�1�}��d���`�ؙ���U�'[*/|7�y~x ��6�>	?����;o����@��Nf!M�)϶��D+���p߈m 說E�F1h�~��S��7�B���Y�2rg�|����|��=g),���A�E��.'�:ׁL2 ��� ߿��?�ax\2>(�8�4��<��4�i|X0�yμ�I��t"K���r(��)!�hCm�|ו�k����cѴ�nj	x�,k0@G3��V%*��é�z_�7l�R����P�f�"���1!X���bջ;+�����Lj���@6�kB޾��Dn��*�EmwD~U6�Bp���:}�:��(�^����R5Y�7B����⪲K-���|g��WuI�o���e�wH;�J�U��K�G[l<{�"9Ga@E�\Qg(��k��V~�vd�f����3_=�*wd>��������lgЁ�s��y�S��$9�`Dם֜���Wl�0��L�aNv+3��yX��'�$�&����r��#o,�u*+(�Q,���Х����YGk��!����gܕ+h\1�U!E�`��^-��!���1�A;�s�6�ڗ�)Œ��N�;�K(���r[Ȁej�m78�]��������N���]��X���z�����齥Q���9m��;���E���K�elS�J�b�wkk�8���mx�t8�Խ�N�h%�+�NMO�\bަ���J������oa�D���t����SoP:v~�����q���"��"wم�mD�3o�L��-C>ɒg	nuP�4�H�o6̈́U&��J��H9+zL1u(�W�j��<�p3|Xx�LSB�o=e4�䷖7�{ڝo�j؆�P˫�-�'¶b�O�j�\L�?E���Gb�tB��T�����!勅	��k#�gb	ΧG�˟�?>� �����H��t�.��X���<}\�9�ސO�}xX&����^��Um�-.^7��޳6k��&$'���H�@�J����mey8�B�% ��\}�vY�٫USQ� v�!�7I(`L�q���!]|~���k2u<��3�R�����r��h�J�Ա��~�H�]��|�� ���;�ZRNU,nɵ��gP!�r�.�O ��N`G%� �_M$oL����T�uOoi����0�z�����\���Q�}1�|��H��J����2�&]n�a	�&���Q��t�\�f���G�L�"ML��^�'ѵl!��Q��
���_-|�N�]�|��z��5�l ɭ��UKD�Cf���ӄ�ڂ$bsh�z����a/%/�]��I�'�N�� �lW^�5�v��T\`��t؁j�g�Y�=���f�FSVg��4����/��u*�
�"�@�3��zU.(�A���jM�k����[�����S�|qL�W813���V�xV[�ώSo����-��[�T|/�:�VZy��P�/��Ld���2}����k��ەc�mtmp�� y~���ɕ�>9�Ք1A���?�ב������ѝ�[�G+"r��+�(��u�/t�%G�L'��tk�E�_���x&��6��B�YD�#4V���Q\��(g1s)U��
�����%'���|��9yeZّ�f�UOF^T���ҭ�y���`^�A�����Y�BRh��}����������?�����O�P�9ۈ�R�q�|p�z��^�����R������C��v4��vS!�(tzX�t"˒y���l2ϖ&�C���ٝ[F�oaC�	��u.[��G�z�cm)�.R�~�6��Y6�� c�/̅T- �$��3��f���2�f�6��v�0a"饪#0|��A�@;	J,,uٝ�*|q?����:�j��`�x�5���O��;�(�T�^���n����/N�@ �ȿ<!�GJ�e��Q�n�9YR.�><���,�&_�鲽u )]���H+���~e��q�c Z���wg�_8;}f�ͳ��05%9
ܶ1	�֣Fh�.y���92���l���2�{xx��i�}���g�<?Y8t���1��r������?~Wu�-���[����r���u,�P���#eɎ~����<�Rj��n�	�t��m`ĸ�$����
V���e_Q)�M%����]�/9 ś	�?��nq6y����h^�s�ƷWv�o��i��z7ο�Z��a��S�KSP|��\�;)�E���[�Pb̄�W���c(&b������S��6+�oY;R{3����N#~s����A=��d[A�5���W����Z���Tcl��=r��6�A�%8��{cfl������h�G�e<=�ܝ�sg�!��֡��P����s?��\�U�V�/�ޑM0ޤ�=�J(�+[<�yc	V,]���p�i)S�P2��Y�=�r�DCFO-�)�:&�׆�n�տ��zc�2.k�aN��h���2D�<^���v��L�Gu� a�6N�U�]<�%��|��9�����G���3��O����������qy�~�e����_~�o����/W�<�l�I}ށ�#Ynb��8;��:Qk ��<�.<��r �UR$W�p�t�"Q�ur �J��N�cS`T}UQ���+a4����Yl�R1M�|�b�5�Cx+< HJ�9F����cXY�� �e,�y|�{k���g�:�|�BO��x�h堭
�T�����,��ɺ�	Z�l���*V	�P��Wam�2��T����e���Zy렛3)1�qpco�����<��
��v�{���8X�X����W|��3M7��X�kTb������{~�L8�]�/=�ٯ���&��h�H�'<���ӗ���sm5)l.W)xn>s���<_�����gxX�>������O ?�	������W�����_~�#Zt��'x�f�tlh�?�|t�L��4���Z?�='��9�w�<i��*�'W)Z 9�
�v��yA\S�+� �H��#�@4��ϻ@pl����=�{ޤp��$��^]��n�)��~���Ň��v���}#s��}�T��� I���,P>-v�1�㬌Gx�A|�9,u�]���5�̋T���mX���F���`�������:2�=YSe\{���i,��H��&���R{y�?^*�6�*�ΰ��(B۞7~�(wf�ܙf������I4���L��?��)�أ�9!�id�U��MN�r���4��",��$�ˤHZʺ.B8E<�.K�<���U�7.�AI���^RGW�M(�����Q��0*n��gi�!���V\Y7��f�/�;��+8���Dp�Є��*IX�|f0����a8��L�����O�������	�_��4������0]zE�I�8��)�!����90&�wP��¶� F��3�HbՅ�s7��� $����
�mj�q�Z�l
�*�U�s��4q�_GF�}^��|?� ��B�E�1� G���Vf�D�y
�y�b��!����,�H�v�o^�C>r��Ҷ[�xΤ<�����B����9�,����g����(��Ѯ�|Q���OJ�Y,�yܩ��5P�����au:r�|�z�#[L�>J�KX�wU�$a���n�#��d1%q��o��)rԨY�9�ŐY����WS.����(X�*��k�[�=??/��L��4�����
���( �7�Q.�:(�O��zr�?B�w�mJ&�(9B�i��Tѵ& �s %�;��%�R�ڛp���c}൙������d�?�xm�uԪ������[��t�Ҫ���>��$VC��V�VcW�R�R�;]��a��+e�~�z@��?�݆E�{�SWE����j˹��b�M�R[�]�`�Ǭ�cǧ�l�u�`��kh2����b�\80t���@ɻ��IR�oѵ��C�(�˝�\����PXt˃32l6�l�G�x��BIV��N �@ �NR9IQ�7�(&��i�4�ěR.3xA�ۢU�,�/�h9�lW+�� ���E��jĺ��VOZƩl^�h��-��^u��t�N䌐
��D?Z��S$��ٓ�zgRԀ
����9/������LWd-��gi�u�����Xm0QT�݂�n�*d�Q�4��U�G[J�h7�k
�B�>��?n���� �l���O�\���u`3ES�h�SdU�y�#AD��h
�Q!Q�+'
#�//xR���9��D�3.��Ě�B#��ШWʘ�_�
�P�|W:fۯA��h˳�c���n�y���L�"����&��\��8�����GC�� �P�Z\�)�vj��N�*]Og���&���d>�1��+;�%�D�����.`{��E}�Xo�WK����e�.����G�|7�Y!0��N\96ͷ�� uC2�y~����<ydP�}�\��p��A��jO��E�(sΏ�p�ײE�4�*��J�F�w:�M��6�u��inn�H�\6e���ɽ&\~�II���������{�R��B��YI����j�`T�F�Y穢A"䭰��u��:�P�B{��V���A�z��e�ˎ9�*k�h����Ȩ`���+�x�)];�.�9�����!j����/�|���a�u�
����y��6��0ɹ��o���>
��s�-���y�x'.$�+�T��uÇ-jf9
��Z�ț$'�O?�쉲�Z�Y�	�BH�&ɿj�,2�I,�r�i��$��@0o�Q�t��(��F�p�A7%����,u��t��5�r_bZoU�%ߐv����t����T1�^*L��\c�8.���� �����~�~��W������wR�\��e��7����#ESR�bQ��S�h��R��uh`{��X��>��On�j��apEJޖ��F�흦e�8R�%���E �x#K�I�i@`'?G�S�8��I�?V�r6�g���b&r ���#n��gE����]n�I��5���U\x܇� ��Ki��/[��h��5WT&�e��O|�?EA�u���Ǒ�&!��?r���v���R}>�Ga�3����Y$�׉��	.�Y��ק���S�Ȥ`�W�#�UE� p����c{�R��e)���6a��{� �-U�f) ���m���z��Y�ߒR��b���5�;]h��9���s�9�鎾ǘ�vU��:��4#�<���WP*�~|��<�:���䞮_�^	���Ύ��Z�.��f�
�8�VM~��}d.nq���
��Fic�qw�˅]�e��V�X�F6"�î�6��۴�z�}��=B�S
�zܬ	ؠ���*�&�V�9���H�ݎ嵲���Us���jU���W�yD�U$��/�Z�O��Z��X�:����ƊB�#�%�w�a���S<���c��ێ��j�
��������f=�G��b��k�lGAQw��:ką��7Dr��X����i_�ڰ���0>�
��E���^�8Z�n"�*M?�R�zH^q���'�塘;��ّa�N]Wӫaiz�]�yk<�~��=v)�˺�t3$A�t �1fE�B#(z��zx8��A~�b!�&����C�)��W�-��|�����cɃ3��˂Kr�v�w�1-�s8�k<D��=�@7d��
渶�ʀ��sO�`�̭_2��;o���q�ʾ���1Kս��ݞ�I�(�k�(�Z���A��d6��x��39�|^&�/��
��_�r��f��c�2��L���tY&J6]�fjȋ�3)X1R]���(��Mk=-*�n5�U�%u����#���>DO!JWtH�g�ׇ4�����q��5(W�tW8���W&(�ge,e�K|�A,s,��ğE��yȖ##�o��w�� ��'��E}`|��<��C�v����DuǨ�[�����E�x�i�)�m��S%�* �:�+��W"�#ڑ-%�I�?M�Ia
+Vc��&1�L�]�,�D�'sh6�@;����Ov���"�!L7���c���R�آ��6�����J��Ą;W�Ƥ���/`��
�l�	�7����F*���ŚJ���p0�����` �e��I�*l@�8�_��/T��E�6�<T�8�)�9�;�D9�yB嬼v�\��������?
8J���z���U��i�gU�y~�i��T6�~˾�ӑ��3 u^V¨X�^f
�]�+�^�-U��5��s�S��V��6쭿�~���J��ͩ���NAh���K�.q�b}�x�����ao���)�@[��س�^iI�(P�����is-�C �o�7�:%K��%�ﰫ���7�a'ieJ�{��q��]��Q[�J��p�]zS�0&�#�lZ�h�����<�{�怼n���޹a�ԸV�X$�@����$����	�e�b�5ϲ�gS��6���єTY�Lsx���6N���a_��lH�����0��1Fخ]�N�=�rC�}�';����ǔ
�Q��U&_i66��z];�*}{<M�7W2_�ͩ�L�}E;5@���?�:�~%P��o̲&�$�$����Ã��y�#ᓞ ��6�0��C�ٹ�*B�qs�3���ʝL��fq�'j4<e�r�6��1mO٬�ij�[,�9�Y���qe�٬�-^?"���HZ��C%�s=�P�#��^1E=�=�x �H�/;|�:�4\q6 �<]���~��L��G���W�?���r��w"�N>�w~��"���.����	���tY�Ήb���5��S+/�~��rB&�����R'��RU�_l��7�Ͼ�2Htr`���~���,6HJ��w
�
���tHO�"�,�(1Y�C��Rvޝf�@�%���Y�xb��������8.�<w���Ll� L�|/;���+̬��� G�x�u�2q����d>��B,�c���;�Ĺxba��D�_��������e�V�{O���ЦW�ޗ��6�7���(�G~+��yA�ë��4�4=�5��0�%��g�
`(�0Aq�K���7��dA�'z?%��u!�Ϡ�a�Vu��R�<??-���BS/�����C�֧��Y1H���=�z5̯���p(���N~��Y�}+����bEk�٦�s��.���J}��I摙�6��5���5�2m4����*^S(_� �P�(�U�q�����v9�+��Ə��cR��|V$�aJW�>m$x�|��7XBK���`�ݕV�VYn�<�oyw_6�:�]7V}�P1���R�2eMB�Ҭ�ڭ�yd�6D@�ѹ�16P�D=7�a���i|M=�t�q���-!6��t\Is(��S�6u鑯����3���&�a�;��â�٧�l�φa�L5�	� U��řQ�L��5��&�ce:��(|�`��erN��I�$���(� ���m�7_��E�4�����k��oL4��l��.���S��3G��Tt���2!�/O��_~��"`>����o�����/��N�ԁt�O?L��3�EH�c�W1yZ���-`�J���/Hk�:иh�����:j��,i^Z��v��Rr]w���I�s"m� ;���>?}���=����D>q�s��%<>�I�s�'V��k9Z����#vz�ˎe�C 4��h����~��-'�j,�@��d��S~mz�İfX�3�� �X9Gn����,gp/׉4�(VO���ʝ�����������������$�>��I��&�	-2�_�6)֝�*fT���@?�`u��=�ΊP:}*�n?T�i`�y6f�;�J?FQ��8e/gb�:��"���?��ϟ���Wx����� ]`�����E;�X:�ybL�.��c�s��	;oQ��G���/��֥n��0�;�9�q�}��W�S�L�ޅr��ҏ�̼�b�*�`��n	�pf|�AEU�NT�*v4��l��>'�^||C�d��25��z/ɼXS���<o�-g
��ˎ�p4g�z<6�GK�*�Q��KlQ��=;�|�CU���PdfU��t!��:��߾�I��>>��Gjz��E��k���`��☙=ͱ%�b����i�HU'��_�V>�|�2Hu�짢��-�V�#K��0dÙ�N]�z��]>N����}��S��d)����~w��� �t~$�G�����I�b��8Cs���T�������%�6�b_F��C�<�|�/�����i��������)1[�_��A�� ��rm
B�R}(�C���[W~5N�zY!��6qK^��D�O0�S����^�z�F����Y0tLJ��tg��C�R!G*Yy���Yy�<�'[�2'+r�޲��Z'?�G���}�0]O���m��n]G�	0���%�#P�0�ܪJ�J�S�Gsf]Q�l������⑺�e���t]%;�5^�Y,�l��9x���Rrh��>Y;R�o\^��v�K�w�!,W���9 ����.0u|QR���T��bg���bm�Ϩ3cV��&P��#Cx?�nUX�wW��NQ�������~��v�2]�Q�2 �f������'��Ŵ)�M�F�w���̕�+F&�J=��[�/�:�[�`�ӻ~��ͫ�Ih�TW�b�z>m��&X=�$w-y�"숔W"��q��*x-Be����@�O����z$ˢ�"}γ�2�iW\��;�0)ƞI�3�ʠ��$�R'�kG�X��v��Sp�4OA`,Q�[HtB�i6��|\43���Gd��g���oI�❵dR��g�M�$Gr,A(i�WDdV�TO�����������vweF�ef�.q< ����ǕY+�!v�J=�(�ZK�P9��$����p��{.XW�շS�r�W�|m\.V���Z/Ԑ~�š�2�ă���K�!B���bUI�Mvw��fU{M=������RȠ�WBO(M*��"ޏ;���<�t��i�̍԰�i(wĮ.j����{��e�Ɏ�m򋘄�t c���J	/<�����d��F�ۊ�w`�b��'������?�_�':�����ʞ��"�/�|�k���p���0�ǠD}	[�GWƼ�5[��$��oQ�x_�`n�;�{x�EC۠53ʢ
����+�H�P���)�S�.=�bQ���o-�wwt���gV��(wv;S��2�̈́RV�����������*}����kږ��עm��j��tk~Z ?tW��I38��g��m���1��:�4�bǀ�F��Ė��u�91�(P\�H�?n
�-��^�;�?�\ib�\;�/g?����(�W}��S�d���`D㠎p��n$��)��K�'�q
`8P��A+g˫y/���I81�lG���MY��Vt iO�_��噎��d�1��t�����`.6�Ŏk���m��(���ˏm���-�_���?jYn���+ͳ�"��6D�F-v�����Z|�ɱ \ֱwIq�J9���ts���/�AG��լ
NО�cH�� TY�|<$~���2X�>�ΎH�&X���<��w2WӍ�g�t@
�8���\���pS�D�N-�Y�3Y@W�3�c+��Ⱥ���AE`�<!���4�[�?�l�$��p[�"����[;~E!��M5���܂j:��� ���&Y��vě�<&�Мc��oN.�fI�����9{�B�!TfSF��)���������jV�!`�3�-4�1A�se�.a���� �X�>��������B���Y6V�ߟ���OtÙ1�V��rօ�:��	�[��4=?[�����}
C���1���	w��R.�˓�5{��D6u%�N��i:�~$�Y5�"�ǳpH*�YuUҋ�3���?ܪ���n���������V,sؚGc�3kG����݁�6����|R`�;�QݮY9fw� 0���fb#��d��A���"A ���Έ~_y�t��(��(*p��9�c�v�&��i���;�9e��p�ǧ���(�Z���ϡ�[L䇻1\�Y�iˊ׈m�_���7I"�K��b�;f>��j����J��T"�r�bg��v�3�b�iT([��W�/�q\�������$�8����������ݔ�GQ����J[Y)��Zb�@�Sf(x5��*�V%�ӗ��J0��_\�D�Y�e�����-M�g��X7��N��)��q���`�H���f�f9{�T�(߮��`�C��+*F�T%��N���n/�M�����I�
���>a�"-��K����4��,��eC�f�5�N�>��>��s�|�}d�ű¦iW�S�
�U��(hXYc�Ŏ*�����ga����zZ���t�q��r����7�+u�s���qm�S@$�ЄV�.��pn��c?��2&�a�Ւ#5J@3��uI��Ӡ/e�P�^t����يU٣.�s��T�8���Ms�Ze�-���i
�1U�VW C�\�y�WX>����7�����!W��Q�lg~���3幺 ".�bV���~�e�4�|���NLx��>B�CP�A\snh�Q����$D���[0ϑ!��}x}�I�^	�d#�6rI�HkJSO�Դ.�R�N���`~Ǣ���I�2Y*=U�H�^#���p��>|��'R7;��]������EP���E8aw!I��tno����R�n~DI��(;	�l��ڴ&Քym�sD�Z�r���1��'�@����c������A2H���?B&�8]�1��q�y*4If,%<̞�t��9@�ϟ����'k��-J�C���{�O�\z�����~�S�l��Y�d���n��6v�@j�m��.[�b�����3h���Y��3hVUe�f��R7�Q�)�� ɬ�yzz�=zwwO���I���BC%��r����ӓ���%Nϝd�sh���㿵�N�_���V�����5�l��,�`N�{£�<��*.�q��� S�����S�`��S�?������ʜD��
bՙbg�������e+�������*vv����I����FQ
m��s3�~o-vF}=cE�,.X�Y�t�X�������5�>o�~�Q���)"�rs�A���x������h4��Z�X,����yy=-����B�q�#���g����7!���_���ԩ-�l�n��(:l��b�W�^S[����璮�ႃ"�\|fV۾���bY�*qӹ@�c-مF�!\m��lɆ��8��Xג+�f��C�A�MF;����bRq�v�OCKک�	��4.����C�4G��׎�s�r����j��������RHT|�� �z�+���>����˿�M,��D/O/����tdz� LE5�N�EEOV�i��'���$9�t��٫=`�W "����������$�|���2^m[�].*ܪ�c�0�B�i�Ժ@xT�5s�b7���~a�A�ѹ�!�g�4�/i�s� 4�<�EM �����$��@�փ��?�LP�`)�P�p2���Ŵ����="BV����#�����D*f	�Y�0I�i�I
�����<7�h6�km�X�~~��ez_^^����yF/:��D?��}u����U��8��JA�S3j�v5�[x�M��[����R@��!T5m�W~���o���wu�)��Խu����X�a� �5�C������-��~] pH�Ν[�@���\ޤ�6k��۫�N̏gkU�X����A�vNlR� �������a,N|��Xa�\�F��QW\����R�g]���&J�;J��-��bIB��dC����jt�����N��o���pG�(��Z4원�xԍ߽������~���N�W�f4µ��'�u��֌v���gm��ꮂ�M���m�����Wp�a;F�^TX�`,f�~�
�����-��*gT�V�p�Q�R)����Pe��&��"��Z���|�����a't��ڍ�K�V�ӣ�NP���N�x?�'��;�����a����D��`YT�@jo§ᤚ�z��-����3�.xF窈��
O���h^UCö���zyOyKh�������+{�{�#M�>�P�t����5X�М�N���8cT�i,�6{z�9gگ�ua�v��U��U� ��5ۍ4��Zk��&Sp�L5y�VW�(Fe_)�/��"�:��Nv�Va?Ԙ_
��F/��(JlV�L���G�w�a8�� ӻ��E5���� �o���t���b�Pj��jj�߀(�>��z�v�]$���T�ٖ����[J�7,<S�S<m햝/0IH�%����Z��Q���'Up������W�':<�җ�������1wǥ]�����݁\��n0*@Xbؾ+Xܗ�`�"pՕ1l-F�ȋ�A0T't��[�����o�@���M�i�v�ώi'ѩ��9[�Lv�����O�>�_~���X{6���GlF���a6�	����&�2@h���[.�5�|KP�Ȭ#��4	�5~F�@����t
nX�¦�\ p�)%�a�'V����*�r�'���Jj�Y���Z��R����8��'��V{9��兞�����͓��W�(W_���k�;�%�Vi�f��gx��7�s����3�F�q��K!�]B�=����r�zm��=�HktV�L;��N��ݣ��֙g�<�T��B�cG�Ji����;��:�@D��uIN�&;I�n�Ê��/��<������tw{G���\�/OO�Ŋ �>���+���Λ��&՗,/���K�J��R&��I�,��t1C��T*(8�n-� 2�EU^Y92���ڞVRM�����f5׃����cټi�$��ҹgP�*�_kW2�H�b��ݫ_z�ta\�۵~|w�*��+	��U*�9�$��ٛ'�D���%2|����ޕ8{�'(�w)Ó5�n�C�7�5a������q���z�+KG�|��~ϟ����;���/���E
@`e�=mB�W�ŎMt���ig��^�=����IP�"����U���XG:,2�o��[�ZlQ�]Ye�)�b�X��>\Ï� �] ��ݢ�W�{�]7d�[e�5}>3����5�*wPY^7�K�7ˏ�j��y�J\U�~�<"?�m�tէR]�g�2e�{{�"|�
��!؋<�CX�nQ\q��f�{���]��1v�l�!���9����j�w2K��J?s�n�(���g�-���!	����qL�jkb�U����6w�Df��Ē�Y>�Z��HI�rw���g0�yW�j7�ii��d�(Ř -�4?LP%�v��������G9�a��=����.��S��
�F�kD�ߤMd���o|�Sқ=�3��.����
ogKp,4Yd�MjM��0�qPSc���������;�����5�^2��Y��0e��e愢�u?���k۬BqZյ���2O��f�$���;_yv�C�=�ӛ�.���o�;������Gd�R�ۢF�3��L����E��^b~����L������hr4��Ir )��c�ni�C�կ�o�:?����r�R��s�^ZR&a_l��b�3�K����z��w�s��B{}�m�y����ѲԞ��|m���a%e�C%w�ͩ�i�n��d��I,�{0�av�t�m4F�ם�����8bI�Jrn�o�ѽf�|}%�8���v[�F=x�B��s|�������u�^)MY��s���&e׹�k�_�C��[~�Q�f�]�űZ���}�&㢋�5���y�t|;v��큵Y������}�}"�{��.�{q��i\�o�jG�$�^�jv��+P�����q�n��v�in����낞�N"U7 �FE����T�������Zא�>T�X-���p]�|��ز�>F��"rҌXb�(��<f잊�^M��gҘ>��x1ct�/�j�/g�]�F��tK���bM����öh������N93�t���I��S�GE�2I��.UUI\�؂��I��r��?$�������O7��{,�a'u?�8:e���S�Rc��

�vc���C�"u����*���3��E[.��j�Y`k	���e���F�t�O.c���2+��3���$�N ��p<��$��eG��|�����s;M|B:���~�{�^fz�X
�Z� �Z*�/��Op:q杣yq2��&�f.J�;��3�ZJ�n�@�RN�%w�O��|����������^�d9 �끂��<��:\��1u��̰p�)v6OI�b"$8��Y�
7'c�cG�M�t���P񁵠�4{~:4�ͤ��X�h��H�:C!ڐ��^�����0�XE��J�A�F,�X�s��URf+�~��d�ݮ������i����r'���ї��R��ךޜ����^!b�*͉Ξ����G)w�������8"(�K+A	C���0��$us��s�}9��[�L|B�Seq�T�by4Ƞ����$�b��g�P}y~��F˞���y�f��^�W,ԣ|MJ)}^������3;��K(PB��@p%̥��w��{	��qu\@T^�ѩ4�P��}��y���z�ڶ�in�-ek��7N�6n�c���Y8�qq��?�|�☦��_a�V��V�0ֹ�5����eq�Z����KP;��O�!�T>=9M�8$6���J�3���J#�X����5�+�5�G�Y�ͦ���p��U� Lk���0�g~�:�-�������a+��Ѳ�U��;|@�� ��V_�1�]5?/)qj�����R�w�kAm\������N�� �:��~���r����J���.��j�g�A-�W���a0[���<hv?uӞ��ŭ��f��#��D�E��
�}fQ@�}xC�W����Q��P
4Dipq�3ܡ�x��zV���ƿ�S��6c[�}	,EֆM+�xn�������h|R�5#���>��r�	�b���	��M�d�!5���-㎳��EȧJ7e�hn����B�/#=?�<>/��Y���H�59��-6�A�4��~��C�{Ӹb]��� ��L��z�g^m��Q�6��G����|�ž@��s���R�^әk�8����w���iV?jҠx����n`�-�o��_{���c����V��P�?��BM�����q�i�Z��B&�<�
@�;"0����:#x��!ը��kf����IQ�ؙ�d-7h@/NA����}�B����>~���XA�P@��ʚ4����m�`��nH'�N@㮭��,�5O��m?�$�&��ۃ[6?�~Ai�������n!�x~��j�����3�~ϵ�y_�Kd�؀@0��oיuNݝ��${�jV�+.* )�C�$�N�k�P���3�`p������_^!��N<|� �w8&�벇�$��d�c��L<k7���8ߡ���Բ�|UJ�^q#ms��b'[x� �,l%��V8�\��s?0z��;�&J5	Z��x_J,�8�.~�@]
�~���'�2ɺ�g�h�F�ڶ���r���8y�E�Y
��Q�Il�6��Ȃk�nl��n��7b���rG2zJ��b
��y�� �d��	�B��;t��})�IK~ŵ%L�M�K�	�O�1��J>�E�/��U��aZ��յC�ل�0�k�>�7�E����2�_r���J��:9-&���i�|℞l��Y>�R���;(@g�mcQ���R.����/}�i�c�ǆ-��o�^>��s��������L�R��R�a��Dz���qEaK��b1h��X��n�xsB-�טd�:��b0+F f{ڶ�v�����)��Vs���V���BО�`Y2��.�AG��u{�Ϡ��c�rUάAHJ��.A%�Wo"���㯈��o�]V�X&��@�%�M,x�"�;ca�n�ӧ�{��vwK7w�ts{��,�=>}g���i,�⋯B��c��<����b+g��o3W8�*J�ڏE����m.Έ��|=��@�;jq��!��Y�c��������p+J���IKA�L��$5�>���ygU\�*���ڭF�0�&ĕL��ؾPj���;��gW�(�*Px��8L��e}�Վ���.Z&l�@]�xx�Q�0`�.�+"��F����S�?��Ϗ����X(�]�ߑ��OW�����2}{Z���@�ʝn��z���Հpe ��l�����eEW�x���d�������� ��wX�ןS�r;7�%�w��A�������+5��L�U�ˆ�Ú�����;�#ʁ�q:��!�p��ߡ�a04%[��eO�O��c������y}Y~�����x���&�q�
A͋/�o ���v��&d0�ht#y�=�b�&�����j�7�'#З�p���}s���n���E(���[�Yzeػ,�l�i*�b���ڹs`X{��V΍� �HQ��A��e���4��.�S|����_��\�%�  ʡ�Y�����~R�ǩo�T� ALG9�Ű&S �D��&���c����W	A�W�6L xb0���N��8� re!7M�;��ZHg|�Q�@��X1���o�<��RŜ�	|�����X������c�l�0�҅Wo�����ۻ�������䙧n@��y��r��9�t��IXi��w�s����~�?����gJ�쇖�������N���8+�5oD�vҬ{��f�5��9{�D	ǥ��PMi]R��3��$W� �y6�U���%�*(�Fġȹ����gg��<߇3hA^'��ʫծI(�J`�8'Ǐk��n���OZD��+���L�B�Sʳ��!,x���a!ć�Nǣ�xX���mבI�,�X����@�����f\�K,Fw��&5�]v�*3��-��!�Ap�3�U=��������^�u�U"��Ŋd�+�ߩە* ,��(tNTJ����4�it3#��J)Ið>q��%��R�p������6I/�R�ld���wk���ڐ�9�;N��IӀ�TJI9��!bHA�:{v�U(���[���Tc���$!g��gq��`���C�0�_�|ĹV�>�Np��YݵR�6h����]2f[�����U}�%v��/wݾ�>�(�<�G�8c��#�	i~puoՒ���js���+Ԡ5�,C�|%��
t����(�rKvC���(4C��T~z�{5���/��akh�.^�?�`�A5�����!O��
#�P�+b��+��&8�SJ�W�E0�Z��-�P�J��SV�ԧY�a�/�7��ڽ~��\��K'o�٠����e�.�q�"��	q!�A��-���Ç;��ݙ�N#f]��eVQW�cp�b�Ӛ�c�8T*��<)�+�LADy�_���hֹ5��JTÊ�4]#���G��c�b����h(��y��}���9-x<���qG�{��@(���׷�7�?�$��S�)<2}����,d��/.��P�?3>��W��]C�26�����|�������k��+5��XGWEM�:\�Ȗ;jQxp~�A�K�m��ǲ		Ʊ�}7>�� �d�F��,h��\,S�4��&LO�G�A���e�,��|_\����� {M}��~tKZ��������
�*̢�~�ʮ�'���8U�"Jx��r���d`b|�<;�IN4&:.B�?����7��y=����l����*�V�>6���(�k1��T�kf�@U�g7=k�ц�S�U�Yo�^��J!u���s�^OX8����Ye;��i�O�b^�no^&�Nm'r��jd��.w���(szM�+[����i�WcS�'���1��[O/N��a���1��	�4����G4x��gƟl�<�h���� ݄�j���i^^����L��/t|=��X��+[��kvA[O���+j?�YCMI$ +�K�����m�W`������-�3��Y51k<]�A ��{�O~s*[#�!�x;7��[��S>@��ݝ��j�X�G�GR�W6ǡ�S��������GN�$^��͐T�j���Vܘ2�i,T &1?��px�����Ța�b�&	%�y=S/,ڬ;kݗ��Ok8Xm��yc��[t\I�ζg�+%�@I��$�z�+w�Nn�%�UǢ���Z6�^w������g�&yNu��L����,��/ܔ/�?gA�s�C&�)f%')�9�(��w�w���AB���Eٳ7k��'#&���5:+es�,�\c����֬�!�-f���2f�o�TZs$�o�Zʔ9Ď�L=�H֫5��bD��� Z<�ð;�ϙ�2h��(8���i󰀇����ڮdn�2U�:�E08�q�-~Gʊg�&��R�+�����]9[���K��=��5.��_�?�B[��+�uZ[E��-�hQ�+�G������ڜ��6�{�	�iJ}�&���#6�,c·�1J�V��e��Fs�N�Jt���^�P�Trw�b��j���6�Zg�v���0I����>Uq)'d�����>I-�˸���6�Y�ʘ��ϊ��6���m��zq������Zk�댔,���B��RՒ`�i gv���K��z���g�������?���8����������W�l�:���#J�O���Ҽn����N\�QE_R�^ט6�F'�	�/B,���7K��u��+(��4���Iέ�]-?~�_>}�su�R���L�w�!��yTNyߘ��R����}v8*�oq˜~P@����k^��'N}�{ʀ4XjAp�&V �3RؚI�<�@RN�d]� �%+-#�z?*��3�t<����������'z}9J�Uy>̂�Q�˯Q��Z[��j�������?��w��*�=�H�6t=�:¯i��w �'��XÙ9�쩛�����پ���[c�QNH���gz[�[�ڸ���9p�kR�g�}SzH�!�@�z�,"�UM|�L`)��A�s����)�	x;*e�ۚW���vHɢ��GL����񕓤7��̄�>��sw/��Ӷ�Qݴ�[3S2-�-�z/t}�W�[�O��֙e?��|XÄ�����4��ϟ�,���R�E_���O�E5 ��h�R�yOkg��Њ��e���z��k?��Du�HQ�B*^a���0{������k=����w#O��|{�{�x�pq"tfV� ��)/���[����x�����Ý*uH�Sō*J���+��ٞ� �i�|3.�]7ʰ�1m�mA�c|5�:�5�ߏfjT\Ј1�:�l�B)��b�re�i�T�_����)�+~[�xv�d󄬢U��}�l�Þ��J��D�O/�����g0��f97�*�����Xj�zn�y���i�P�[/Ӛs1�� �e��Q��}�c����-�Ͻ����T��^�5�
���r��Uw6�9���e۫=�+�B�v��>���ME���:���t�����l��� �4p��0i�%��ĸ[d��Q^_��\>�
Kz�)d�x�������|�$��$T
���\f�� �t�N�����Gu
D�j^��p����&�+�_��m,[�0���N4x_�Jm��s��A�k4�?������f�PYg4��j�O�DwLXc�J��h �a�3��z�V��������<h�����]�_�0�$xb5�F���g�Bq�s������U���e��`�UөeiwH,�KM?#�����5�I*��@�
�� �2�,����?~|�_>~��$+��i,�`��,(�.�n6j�x:mseh�Zt�`���t�P����ͫӅv�e+��)A�)c{L�4��+��¹�����'���P����-�b���i�Z�(XE���sx?=/ �c������dYaZ�c�0V��2O�APN��P��W�#�.o�n���� �t����B]?�"��?jy��"n�
���B)ٴ�r�L,��b�ύu�`�3J�lp�����L��+�d�ChKO�g��pn��q�58{�L+h<(��A��1��N��'�@�J({*x��v�E�G����fߚgF�Y��Q��ݽ�d�e����nE��aease}�[���l���N��^�۸�	�#(�3��R��:�JJ�!�2%RB��KR��j�-%ӦJ.h]�>�>Ř�8���(�N7��NC�g
�>���wf�H���=ʹ��ބ�sg�ғ�P,��c
�R� S��Z��էO3�-���%��F l�,KȔ�	�ޔ�́��6cM�p��/aʞo��D2�{ m(��&��r�r�mh	u_��|���[|��Yi���b�#޲�^;�U�H�\><�@ɯ�ӂe^���E�:%���S�kC���[�vO���|l�]�O���r�s���չY`c�e�X4��î=����<�9���������k�:g'��w���T��*�.����) 3j���(��~bu�r�����䌾�����4,~i��D^��u�q�|8�b���i��W(��+���C��^'M�NO�w�U�ny.{��:Y�z�>
�׏oX�f%7ZBv�}Kf����W~���[k��h�*�5V0�i�E��ܱ:���_R�Չ��EA�a�ƛ���J��W�������g:�%ȸ�[�=L7r�r��E�W�F�[�
��6^�6�fRB�O����²��Ԩ�H=P��qܣ�n*�<f#e돢&����s\���lb	\�ZV�[ƉR�[k(�~��r"�U�.�m<�d�=(��ɷ���-�4�{ �+���]?�t�{�����w�^K`4��;?��a�t\�]��,����������^���ue����rTt��#��I�`���wb�љ�g�X
l���/�=�IN�K)?�\�=	�|�Z���ge���w[ A����)%�S�nQ�E��)�*U��~�`��q���W�ZK6���l�7�4� �����l�s'���;%��e"�{{��J8o,��vD�`���l�c5���vJ�Z���,LY�;���o��zޣ�%O�[J��t@��l#�?M���s�NC�d�S%��W��f(n�n���V�9��s��'V���֟��A��E��L���5��͒!l�.	p��N�|&X��]�a��va�#���s�1�1-���*�*|�t�ݮ׼�����A,M]t �"��?K��{��E��D�&� �O)���bR�2RCB���I<����m~`��WTe���T�;�X��k����{�#�*�"<��	�8�'�A�&�,1A�.AYQ�e��^u�v�I�fKU+�.��j:
M5z�<[@]�j�rg�,�l���FǴ�s/�ҼSR�eoA�p��ƐS�=S��Ck���֣5.G�۟�o�rE��:(��-k�W�v���W�l��BO_����zy}���W:,ߍ��nfvO����&�ۢ�N�2�~��=�Q��1��_:ٱ6T ZJ&ӹ��/M��ߒR'�i(k8Ȗ����Y�Q6������T�u�8I'��wA��-, �g���^�f�<��L�5Z����j���iݛ���xL�1+�YI�W��mTh�k ffQ����?� ����#}����u��o7�dK��K���{�K�]���3W����t�Z�и������w(�⊁�΍��\�~��t���.������˷�w�M�K�U��*ĺ�ߌ���)%�+;?��ϲ �2�^��8]U�Nq��̶g4JVM�$����iٿGmg,���}�i�0I�n��2eR��:�A��\����%��)>�[qA;J�R�TS�$�E���ݩ�l����ф�I㮝		��6���:ck�{~��Y@]S�ʷS�rᷟT|�R���?�5�/�v5B���@���{��M������u�.	�J����S'5�l�a�8~�qA0�6ş�~w�?ԋ]�6�
x�'�M:-뼍�%�H2�4R�e�����N��\�
Y�:,$;�g��N�+��{��?���/�Q���ug-zz�um	|ϒ�#8�{���
\��;�#ͅr����7�WY4U{�0��n��!���*r�V��4�=y�T�i��F���Z̿A2S�����ӂ%���R��"�1,��i�0X�T_g���[�8��WuNQ�C7u����qa��QO� wn�>_K�Z97�e������3z"xKd���������Nu���[Q����e�eӾ��pM���j�Sܯb=s��E����o��w�S�e�kJǅ�޲vOLbY[#�4���%?�L�S���x��G|S���������x̶�Hm^�)����B5��qV�������=��=�gV����~�Xy(����M��B��F ���5j�4�����1`�e\6	G9۷j�9� ��U��5��?ij�R����W6af?��#}y|����������z	*9���a�+C
���6�d~�b�tc���և���Zi	m����;pz!����t}��s�Xo����a�m����Q��u4����r��󚢴_����zN񌚪�
�i�`�_�Gݘ���d���3��N[��ZnT4+w|�gS�P���YlY_�X�p��b�*[��-��65�$[�Hp���tL{�s���K�XI�㔾�t�VJ~G��SW�@���S��8�Ʉ��^椸�8�9��w�z�~:�'�"(��|zL��-���T�ʖd+��Bߑ�^jl�����Ͽ�ǯ���H��Z���P�V�p�䇇���F�"Y\��};@)d1 T��a��9N�z�{A�N{k��W���?o���A�.�_[�u�}�����C�.z2��ە �>[=�b��H���L�c�ǖ9/�#==?����,�����-�+ѕ��ӐxY��W�?d�r�؄o-����1�"���� �iC͓� O��D#(QP����:��g���+����-�]c�G�p;��c�Tm�|.��w���KF���,��0h�+���'Y�-��1���Yi'�ñP�a��eq�dJdA���Z��5���ll_1��#G���!Wo��?`��Қ�KT���W���F��I�!���?�EF��t�<>ӿ��F��N��q���������hUi^g/d)V��Em̚��Ĭ����ۚ_6���٠i���D;:�h��]�_;77w����+$j���#q9%�X�\R�P��W�n��,�E��q5��ϡE=W�w��o��$��Uצ�kv���mj�3��L�#D��u �z8- �S%���A\�fX�����Y�K����?�n���Ԑ�fKj�FU�Q����>T�1d��*.|	ݯ�n�Vg�΢����g�����JzxjWV0t-l ˹��{y�zA�J3f���ʺ�t�����[E�82��Cn�n�P��	]N��<H���C��ف�v�~���Y	�<���S�KܺA��R~_�<��O9h�I�����P'd���@a����W����r�3䟓p(�g6����
���0��1AdK�\Y�Q�ыbǭ>-�t�`?د��G
v�7hY|/�|^3�j�/i~\�t�z�ҵ0����6o�Xw�Ɏ]%6�Z�p��[�F�t��U32�]��ڗ����)Y�J�+���n�u�?-��F��xSe��6¼M�����e
��I>��z�3f����q�>�a�Y�IN�\p�����<�b���U�ɡ��4@� ����?�����v��2����ҹ�θu�j���^I^�r?@�TJ&9f�qmM�Ow���5hg�<�V�&����m�Z��&�\u�|�\�D��Qݢ�r�,�'Ku>�5Y� '̒�E,o&�
��4�
��X��8����͖�����u2dnw`�b�tCVk^O�
T뗾u���59'̇'��;�?�[??ͽ�5���k�|�7W�T��񿁾I��Eh1=ԍ���b��J֒�/_��2(}~y������.w���8�x��7��Uz���Uڵ�YJ^�q���߱�=��X������|���O�����Lq�� *�0)`�I���1aoY�\׿�5F�}d6�`��ER{@�5��9�&�M[�	t�҆��DX�O"͜���0���z�<���Yt�D/��b���ʯ�����L�.Q�]K�,��m��U?��YV��oAQ��1&N��1�o�~\"�[h�$='Z���9��K4�αf�-�@7���.XZ��Lӭ��u+���W�$R����j��v�����t�\b��Yə�.��+�
��s�_�z�����rf����T
�E���!є���H�ӝp�:�ܙ����T�3̢�6YM���D�?s�Wu��Z�l�;0�sD�����9�l�ŋ\�,v�S�u���B.�q�gs�؊����n�=�|&Y�X$k\W)�[d*�y%I�[�s@EM�zo)_���o&�$��(uMkф{[s�~Ŗ:|Xuwk
����V2�d7��j�Y;��z�3X@�j�^�{��U��W/�e��)��bO�����]-M�7@�9��kŕ�=��oc�~Zǈ�仩Zܱ�}%�N�w�uE0%xlu���I;��WE�4ľ�=Ѿ�\��r?�\b3g�u��l��n@=���w�Ҵ���6+��l��Zۺ������m���㒸[5���\��=�nY}�d���bi�r�)���v�"��T1��T��ܵ&Ph��Òx!x4��Js��U�Tt����5�K���/��4Y��ZVR���3�!XK���`�-��z�����G�+�_��؉�F�,�{: C�=�Pw��N�<j^Yl�|���?�V���T�1!�u�d�*i�'�#��fKBY�����Q����'�YZ���u�= ox�F)�����ڣn�i���oU"�� �����P�t���q�n��W�����	~M�u-W��p홢�cJ|�_���v�*nu��]_��p#>�:`�1u���r[̯@�����|k�w���[�Ӏ* z����Ғ�rZ9pZC&�T,�k�%0�G�|�WZ��|�N� \W�d¾q����u�h���6��|�P���1Zw��3���}�ږ&��(�𐖸�R���>E7Kssz��v�/�~�mkZ��h3���:��*�֙��%r����ks����>��|�k?�&��T:���f	�up�;`������|��SK�i��1��KpA��ò�w;�2�'�A����-e�~L�8y~b�rEF 6��R�U��{"�y]�& ��z�G�%o	y�0p���Yf���	�5V��PڣNO�D(��������A@������hV�L�ZJ5GS0w=�Lm�Y�L��W@e�ܾ7���f�U���oH�;�m��Z�Fb����J�:�w���Ϝ����f�QpB\D���f�tJ��Ξ ������(b�8gId�����j7\�->ts�A9��:~��ڌ�k�'cϓ�.+h�u������gI�2&z��^��]L/�D[�;���z�b�! ���X�3�l��Xv�;����Jo�Ӵ�6���<�)`O��#�D�;3շEOһ���={:IjdF]�r��>ި�kJ<fcb�ƻ�ך�4EI� .��$1:ˁ�,�9߄Kdj����h�!̺�y�<�6�����S�0x�
�\�b�(��ǢmPV{�������FlkE{S��JfM��}�(�ۆ`M]x��J^�5��z��v�
����Ãy�������]�͝�X��7
֖��>��Q������<=�e��#v���h�2��2�SQAY��Kz�AfJ6??&:(�����Tg��՘��K'�-�X��w���@v����a���7�Eմs�<�����`�� u�HN��ؙ}��١�i�l���4 ��d�R� iP�Tۓ(|���`�fѵ�?Ư� x�)����<����ul7R���4a0�6��2�h�1��D������ǁ��p��/��EҜ8 YY�~��t����v}����\�pۍ��s���5�NU���Du��ńr�i�4�uMН�����J�������c�u��S
��Z�z� �m�a��&�f�t�Op����	s��඀=��#�k��\!�o�0��*��joV[��Ҧ9/n���C1�[2:�@�� �� �e��j���{�P�P~�`����9���P�5k��ߌ�K��%�fk��G��|nkJ]�����!N�"��^2�I5��$����?��z���ds0�+I�5�'f�<ն�I��ZѩOB[� ���;�p�R%��˜����`���g��\^=+��t�>!(�"3��)]��k@��Ӻ�?��N���Oݚ��ȥd����oc$0�jL�p���"�F{���	i��*� ,��<�?f�%�~���"��F���JL���.X7�vO~�Z��m�S�VG������=d�3b�$��un�n�';��(��VqC���1�u��FT9HUW���b��\�7ܷ�)3e%�6=��R��X���I2{>K��_9��gɆ5)�a7���z,`���Ii.���r��^���Ɯn
Y_�
<��f��C�c�9}w�u��犲ؗ�p����FںT��S��F׷����b�WC��W�]�~j0I����(Y?@+kSOi;�'���D�)�����c������g�%d?M��I-q�����_$��F 4����!0)d���q�����ִ=�L�f�s;'u�-DDĔ᫏-� =�1O:"%�����o�)M�~�P�Vj01h�Ve.5syf0z�N����B�<>�]o ?˵	v��JX���=�S��'�;������闿���F3�"`�e�>}�H�;U�0#����Íh�Xݗ��o+=���no~Y�==����>�b�D��m�y*��=!@P��XM3k���j�d�������Z�wbYc��h]���P� .5����Ib��io{?S�B�R$ϭj�然4k����=,�+'�?3�}�I��J�O�^, ���	nR���)��M�9���&@�{�Oļ�c'�%)u7�J> U� u�R��߿З�_�<�R�$�kt��h ��J��g{��XtX���~pT����,&��M�kL2U��Z�d%Hffymb}s��js��0�����`���9�Y ��[��$��UAq���JnqzR���l�s�iAY�}r ��J�t�!4kO���L�@	�޸�_��H3͕�m�4��[ ¨0�AMI��4Hy�U����qM�bL,tq��6/Ճ���0����`�H�M�����g���"E-��W��#m��Kh6W3b\P�S��N����aQ �_��&Y�A����A�__U1:R�2`��OX�+��紥!q�b���в��,�|�Re���9��I[�5u�ǒ�u!�!����-&�������j\b��}\-���Z�����K�w���V���~w�SoQ����`�v�>�e�ym^���]̙k*��I�XQaP��a_��<�a\�5����gP�Fn�k�l����Sݭ�d�mc��M�^��Y���S���ꮶ�n/-S�;���nV�ȡ<������0����%p��7'��#��7On:��:s��K�
��pa���
{l�A�b��Y[6�^�9Իjĵ���Dקo0�69�&�|s^H.]K}%�m��]t׺�Rbj��� ߖ��0��=bT&�Y|��s����$^�{[A�����t�����M	0f~F�p�ڈM�`l��&����)(b�j��ܯ{H�3�@���\�?�,a'2����K^O���ʬڵ5�@&�(�1Pzzqx��K����c<[R��_�+~��剶b¶�P���ꚴ|��A����үEV�O&�YT���Y�BF�P�Е��Z�&I'y��@��o�L����txz�����ϋ��|x�4�����J����7}�4Ӟ�<� ǽ�o���H���n����@��������Ł9�k/6�1���J�7 "�������Y&o/.PUn�E������^ʍA��rJ�t�of�śZ3�!�2�+6���\;ŎR5;ֽsƼ�
/��]DMG����UӸgPdW}�Q�[ݾ�S��R�P@C���;D|O=&FU�>N�A�̍��T6�H��#I����4���LL���<�-X���o3]+�rPG�b8���i��N�>�z�kM�-��`�W���b�-'vE]�J̈́��c��t�5��#����H%�y�u,����$'�	��8*IМ�mn5�x):��u���L��������jbl� ^�Qj�`4�� ���}>@ ���P@Ω���A@�u+2%�����`mߩ+�[�[�j���hV�`{
�Z�m�0Ӯ ��5={�<�9�%+
�԰�^ �����|99�qݫ+j�H� (��P�`��j�"y�������Y%U\
N��"�@ŵuP	`N{Aْ`0�<�פd�:N-5�������9��^_!�7:.������$��s3�N�1c>x�M�@�o�R)�o���J�(�0z1,�	.�A7�['����4�� n�{��~[}�Z� �J|�,X�2����A��V
�ޏ-� �7�N0N&��]Qh{=+�����5�B��V��f��x<H|�y>�*�ؚ�bpI��P,�sK�8�6��=&ݏ���1�ʖ�aM{�4O�ȄW����Z�%��dƳ�Xŏ��2�ʯ�s��|�����Q
�Rg!e���]��0��Y��4ChV�N�t�c7�W��[w'
y��d�LUz$!'�;���͓�<SP�����	H�}]�Ք1��8	�&랃��F�+2�#l�,7Y#� �ِ7�Γ+=$��8����)^�T�Rֱ۠ǃ�!5p�jz�
��V�j8x0xn��8�ǃ��TҞ�d	���+a�Vq��t�[r6��
A�-��Ǜ*�{��e�Ej���T�
8�Y=$[�����BG�Mr��ꂿ�Ƽ�2�Z��y��O����|}V�j�Y�qu�y�8��90^i�W����*�U����}#D�_)���q��o-_u�C��5��bӄ���-5�>|������s��d�zz~��>֓��D�������I����=?=�[����?|�_~�'���_��v�,�����|6-�D�)�=?r[����\�h�,E=��N��S:��X�z�;P���64�����9��\��"�����T>�SߓnhV"���T�Y	!F�<(5@�p�. p~�K��R��\(g�	�[�T{Yo>�i,�\�7� �Wf'�J�J���z���IKl��*n�ɳ �'S���j1v�74�o�ߪG�h_+�=���8$���q�Z.��u�D�Lѥ`[�*O��tfq�SӚ����9�Q!�d	\k�)�A.a�_,���	�����;��`��<�J�ֹ��}�J�\�S�*���*k��r��Z�{��3ڤ4��%���������Ua=d��a!e���7���-�J�ZQ���*-���i�&s�s�lױq�5kGV[�[��=L��N ��M��YȟQS_�ɕ_P��궲Z˒ ))���(^�l9��������yn��Σ)��R�R�g"6�� ٬Fc<V�2MGz~|T�Q������Y�M1Ќ��d?y\+��GW�4%�d�)6��z��XǹΚ�V�>�p���NM�6�������Aͯ-Xn�"-V�@l:���:w���2�>�Z�p<3���
�~,�4z��H����ť�/�����|���u�o��W�y�X�΍b�G�{W�jw��H��0���[`b�V�2�a�Xm�Cs�.���`]�aG�7��Wk�A��+���r1��;F���� ��~�S���q���#���~��3=����p������R�]۸�c��o}��G�R�;��N�Ǥ�e�uE	^A�|N6��Է�',�3����T*�iXj���1P�����HrS�5����:�E3��9�IH��=��7Z[�|`��r �g^��T�4���e\Կ��5�e�/�C<3���A�D�֯� c'W��n�n�$��u`��_����?t2��הl�����l����U�F�Vn!���R<s�4/�X�d�n���:�{�+���Ԉ��A��a}(�Fc~����]F��p}��>��S���
:Bg��n]J�e7l@�\K:���$'$b��D��/��U8��������L/��:�鷿��no�Ç�bB�.���Lr���t�r��^� ���]�0�7�䟤l0 �!��0��%iO5K�}�+�t���0 ��I�*v��Й��`%�0{�d�
v,;Wŉ;��*E5����c������<�j7�YȤ'�:7� �P>e��k���B� isG ���ޏȞC��)��K����3x������CG	2q&���N�`+Nޡ��4������
�1��������V��`�e�k__F:�[� ���҉��	s1	SQ�c��X�#Q�+��o4L��`��A:)(��V�`�� mG����8�zMh�X[��Iq��g�˖yv@�ՊJN��~�D������J�I��h�͜2[������SR,����ƩU1�aVF,�fU��;�����c���Z��9K��h+ -K)3\�j�F��*��`�D���'���B.��t^�[�� �E�e��ڭ�jm�2��h�1�4`�*���ֺ�c?ٱ1�k�~�<?���l�d���Rol&ϊe���t�'�w���f/R�2~�>?|�$��dVc,8i��w7�����˳�^�����q6�2�c5ܠ�4Ͼֲ(v�!��X���r��Db]i+��2\a9(��~�$+�ӟ*m	�߳dU�<	�y���J�O���b�)��W��V]�\��8�*�^u/��h�Cϓ�ݜA���m)�yN�dڶjz���q��>��wR> �&w��G����)ͳ�`��J| ����d!4�R�@v�Q��cm�˴�BMc+e��5���������I�%�"�8�Hd�2\6�;�Gb���r^�[��юun��4g��M��i��)�Yu�aX�E����٬V�hl=օ��Ҷoi����Jۚ��C>܉�����3��j��Ҝ�i�\y0�}����.p�nF"c@�H��5D�-|�K�N2�'r��Hvc�1V<��N�1)�Ɋ��W���c��=]S_ڱ��w�t��*<ϰ��q��-&�Y �!��`c]$n�&D�����[��ӹdZ_CI;[��GA>���JA+���Q9�.����~���=�6�
Ch��n��u�w�0��'� �
�R�fs.�n������㸔B�;\Ռ�Z:`1���D}Z��\��b���ǧ��
|?��;���U�qae��c]���ˋ+u�d҂'b��L�p����#N��Z�Լ�̺R�|ϲ��7�	�3�r<���:cA��{r�@~��~g��v5Q�X�t�;M{5���z� RC�6<V|f�Y�о�����`Zܕ�j3�N.^o^i{����B�J��t�UQ�\}.�[� ���\��0�dAU,<&����q/J�ǮZ��'e1���#�<�H׍���d]���1b�le��@�j=ff�U����.$5��L�/ǅǟ�=��VJI}���i�G��*m�{��/��F�g���m�"(s�).��,�R��+��5Eu5sփ(~N�H�072YCg�~���oe����kZڱ+'3K.���@�Q�r-K�v{Ā2 o�Q�Ns�W��{��hϞQA�ö́��~�W05��V-6
�2b���J�ͪ$Ŋ�A�*[�ۓ3��Lz�l'Gi� 0��ka"��D�m�b�8 J�� �`_D�y���nbY��D��S�|����0,'�n�T��%=(�6P,�Z�X�W������_&:F�p�].V:mn[�^��X�TK
�����	Hs��kE��M�£bE�����vi0����%vY�nO�D�E�]��?������!��-+`��=m�K|_�=o-��Ĺ��Aws�M��JfЉ�4S�['�#����X�t�
�H�P�P7s+��~���3V��v� )\?Uh�֦5�w��}�*3n�}[b���g$�JrX&�Xv#�1�
?��
[�:�/h�c2�ZM�<Ne�U��pB�i�̞�~-.�8�bgƮ5�����oX�5�����`�����_L�T��%����	dUM/X����C�����f:\ϼ���|'���d䘞\	�jZ�N�s���yΉ60_v��Qǅ\��f�����&H;��%j�C�le%*ښľ� 9w�C\�����n,c�@�p����#Ƒ���|�UY�X�-��(+7x���m?��0�8ia³�gQ�U�xA4����S�jzp!�A�/n6��4N�?�C.�Cߴ�[���}F�5���1^m��b_?��N�H!�7)��
Ϸ�\�2:ѩ��..����������XV�'Zm9�;��v<�JE,�
It��L��]��k9�ī�G��������xpk��}A�c�f�kwZ�#�3�J �@c��f����&v��i���:�.�����U��X���Ї�;����Ϯr�5��(v9E� "y���B������q>0�`�A!��+V��t��P�L����^ŧӽ�:;m�Wu�)C��2����ϙM0��5R��N�/N���+�&����.�����K�,�r�QA��~}[�bQU2����I�!���q��=�Ԟ�	����%#[���Pe��� C6�g%ˑM�����Ё�
�]݉�N���)nDy9Z�̝(G�':^�X�!� ��}���*䟴su�SO&`t`�i�1ͼ������Qk��	�Y�M�p0�9iTC|���~��A�y:���qRa�Ý<_�+\���:����+!���Xধ���������5�s�%H��`�+�N�VO�z�u&
֝��:����U��Mglps_]6IIQ� q��S��Z^k�P��xΣ�+@w�.p�7�U�15��Lv
�2�~�D�o�mg���y�O���V6�?%aQ�Ϟ����51 �n�߈p&�Pc�q�N'S�)�0���ʼ�^]j�G��#������ߔ] /����ƥr���
IIÀ���̚�"�͖ ��;5�K�X�r�����`n؏��⺙�(��na�@�C�K{ß��i��`9d�,h��i
\�� �g�:��=�b��gk�qd�} �B02��[���p����J�8r��P�����%�e���Hذ�>׾��?��V��M�|�!��,�Z׾ē�����9p�樥��4���,?,|y�\��O�D�5c�WGo)��B����2uE,*˰%�ĸ����BCd�q�q�w������\�`�3R[���Mwh��3�29g�\p�3f���B��hQw�$]���u(ݧ���^�z#f���F�t���+jϊ<�7�@eD�s���[�ڨ�����2����v���h�8tV�l�EV�uIeҺ�z��e\��2�ޜ#d�ɞ��|+^�:��u��4�=Y�t���gzC�M@�<�氏��A7Q);�,Vd�b=�B΃�������3^�C�$_:�"�+hER�e�%�?���������wXi��������M�\*D����t,B�O�S���T�����?����gQ���.if�!��(@_P����Q�f��FF�	�ݺ��ҷ����r������̭��ܝX� ͯ77{F�u.m8��mB���(m�zN��N� �J�)#����w�"�P[\�s�z���c�e�L\+�������d�*����<?g6�]��zV!,][6>�����pc��A�U�px=�a8*0�*�n�4�	$K��*�����J�^��WUh��+�M7�f?�z߉�J�{K={���L	��P;|���N�J��JX!��*j%�s.'�ƌe��TLr/�#~��^�{X���4Mz]Ɣ�����R�<Vn�f���.v�J�	*�'��=��w7��X9�A��j�&�Q���*���jMqG$ի�\�����r�ĉ�'z=l;�5���v��S0,:˾�<s�½YG�[��f��gy���E�"���)ux��j�����pK�w��E\f9�D$���u�:����@�8@�xU6���i�/���>��l��>�sc.aVE��ʶK{wq��4I{����y�ƈ��S�D	b�A��B���f�/ً���t�t
'��(��{FO�&β�8��8�Jz�(unHZ&:,ߋ5����^صP\��A���
��c�1+����)Pw!dZ�Z7q��P�c(�}d�Z�z�B�+�%��M�.��E��@����/�ha������צUv���e��uA�L5U���GQ��Q�/b}$���\�{�wS���P����Y���k�5HE)����MB �݉����.Kd�?d�>,&A��D�;)�2.kF6_O�r��u����(��F0]P۴���H?w|l�2���*��)����@��i��m���H���]:����Ao�����%G���F�!(g�vWE��ٟ�o���U1#_{�$d\n�x&ء�������blg|�(	�r�b�����hm�!N�Y��8���|�C��8*���͵�GW����c��Ԥ�3H)�G�*U�Wl���5���0��f��i�<�:��H\~�GY	 ��.J�����-��@ю2 ^cV���(�
gl�����Lw���V]�K]냻�������5��i?5{X���9-��-�A�{:PbA�5���5k-c
�d4u��!�XV�A��}��PjM��uѸ��3͚Q����0����5�&/�l�U�Q�q��P��u=iTr��_��<���4�]]�՚�������su�N���{�.��7�/�=A4�/�1�|zz�WIѺz�|Z^od~y�B���������uw����ӇE�(������v�*i��A���h�60�s�C�z�d�8���8S�[,��K2P�v�b�{��{U����D0��	�����}0��N�I���~��,r�bL�L����-[썒������z��b���z��:�f*���i'�_� D�V�ɫ6kʶ�)p`��	1����8��f#�d���r����ߋ����3���Gq��d/���V�#� �u9��ƒ޸�;U�b�ȉ, ��n.J���k3�����vz�)�pO��Tr'���;�c?=}��)�.��'\��A�jk�?��˯����0@�9�2SW�2c�'�Pa�����]X8���ӓ(���B�'�6�k��I����?��_>�e��13�<��ݨ>?ɖz�Ta���#˧��̓(�>-��/����������;��_�<.�.c�<�)E`Y9A):Ij�Ċ���w��v�K=Z�9�у��%��+_��2R�g���Gv�e˦W�|�u���O��>}|Pf_T�ȱ��Ĥ���^�����n�yu0�:�Ӹ�2�� "�VH���`��kJ�����X�H�x��F�'QF����0�=L��e�=��'���	s������8ŉ�՜�F���,N�#�׉=[ �ݠ�7N�� ;h]�~���d�c����o�K�ʫ�����u�"H�����pS��tXrvj}ʀ�ܓ�lJ)n�������B'+I�r:+�ʅ@�;@s k�U�-S7���lo4����j���m�v���'8�U) �9	|5UO5뿕��򒻀�0~����x0inI|���)xN1�6��� ��K�q����b�c��*x��ִ|���Z�w�X.:,�q���XW�}报ʋtXc�pat�=����U�,�a���h��_�V��ϋq�j<[�K�Pte�ck��}P>�Iי�#b���[��0��$8�7z���F2@�(�ҁS�D
�ǽ���Ø�&�^m_`��X˭�1*�e9\V�t6"Cn`�u�)�(�4#,�jq�5�ީ��;C&RR������9�/���ە�����6�B���Z�-�\���p��3�R?�严�/��v�1o��VۇI	����͚�����8���T)[k��������bX��0���a�.y��aЬ��=�a�$����(�Gu�ͪ�����Z)�/�&�B�T��	a�E�|1�!-��M(ֵ| ��,���?��<�	=
�"�;ut@�
̳f%��4F`ww��[G{0��›�t��[�. [�i��t��Xz8^��&�+е/h�>���OãW���}��Q:��$"($&���ϫ?ic^�"ԟ�V����w����im�pdKQ��R2����k`f(��@�U^�̤Y �es�Q!�}^^��*f�a
Z���L]F�h��5Z�K�v��Um1���~�f�c/l7ˬՂŪ{�D���M�U����@i�d#��L!��"fx�bb8!B|���J��Z�W�r!��l��5����=8Jت*!�C����R�Ѩ}�lK#�ҲZ"��\����ry]��,j��+F��9�P-.3�� �9�yk1�,�轁�R�+�jF�����ֻ�4F�׷@�  �iv;ĩyUKV��vfY��� ���ט"�,��O&X��7��믿�[��N�}D�BV�Lc(��]'���FQ�=?zy�����ce���5f�EO��>���1U虭�ĥE��D�0L�Q������Z=<���̖5�p���=|y!zyej �����0������;��s#J5n���Y\+M��G
lX`�K����a-���fig��K��"������iy�(md �
�/�b��V��?�a�iy�3�4���+�c�*���7��%�Z!�x��"Fl��`�+vX���x���l��]7���$b�͕�h`�\ ��=]��~Wf��j�{ �-��Je
p�.�������;U��(§��g�"U�+��ݽ�`~��œcQyݙ�i���=~3��,,nƳ�ű/��Qh�*w����1�S������*���� p��k��_�6���[���c�kg��Lf�9��FᎵ��Dl�UP����l./�nNW��.���� [M������t�����|~1Vݏ�SnoGQ�3}��_��������;E�7B��-�0Mf�k
�Yh�,����	.��;����ڡ��,�̬R:���5��=�_0d�|�����f{v�Z�:���J*Ʉ��p��F�>Q�^5X5ܤ�6�ݍ�{��E���3c�9�T�[г~_��Xy��M��s��*����Ԍ �2���+��ØC���O�wK��,�J�tm���DB}(�|L��qf�+giwA��bV���zTwg���֔&�+�;�/W���2�r����x�%= X�ŁG4�C`v�Q�_�v6��,�!Lb>c���H��X���	�,е���g�XHfmDھj˺^M�8\WQ�|�,�C�C�L�ę��WQ��~_�֏gW"�@�
`��+���`1��&�ҁ]ٹ|Sy�2T��_�S�>�b�;��"��4���C��ƽP�ﴍQ�J�K�\�j���l��x�D���S�p�Q�;�b�DWV%�;�@;N�l2�B�Њ���k��:].�w��o|Y���'ԍ[vmó��O��`�~�Ƅ���Y4�L�D/�Y�R,4JuH�X	Q�y-�ۼ�xi�7�@btm,������h6m�J���i֠A%��A���Ajٚ@��X�,�h����J�e�јo�v{r�#'@���q����a��jy]솑�ܵ��xq����R6�f��K�`�)+�������9��=�_�R�t��6b��	�2����!��DG6�R�ా��i�i���f�@�� {'Jin��T����_��И2����ӗϿ���V��}���$�-�d� �ʟW��T��hL�9��+�Vw��˯�.���f��]�^^����eᑅ����n>|�WU�wCaN.&� U,�ĥy}���{%��eY,��WrF�����%�+{��eHvw�@
������p���bwW��$2c��`׾��%K��&��y��LØ}~ũ3x���;�-8޸d��1Rb�gp�E(iß��q��d<��k}� �˨1K�вrE��i(��X��LK@É�2���r;�g���� S���t�����@��P���>&�u�M_��Lc�5����M�X�e|�Zr�D� �D /p�eo������nk0���8���s	|m�I}�4�5k�褴I��.�e�Z���b��Xyh7���N�*Z�$�F���1�4h7���Gk��l�	UI��w��C��uǌ6e�@2���Ul��`[�j�AndDk��y�{ry�ݑ�yz}��` ������,��4W�>'�`��{ٝ߷��9^��S��}�=�v�����Wv��iܪ��	l�]�ը�Ԧ�T�B;�?;�߹U}��w��b�2�_�w2Ծx��~Iys?ɺi���6y��䥮ز�}霙E�Bi��`gH�;nR�ᘳev�L�alK"L�;ϵ�/-K���W-��m,Z�O�2su*/It�<J��3�<��;�~��Ґ�k�E �)�#��pZ������n��@y.�cr�m�G��4�J{O�3���p���"ki�GNީ�Ҁ,)Z�řt<�u�L#���J���3�}��pێ� �`)`%�o��	.+��u�h��"��B�G�,X��:�x�<��D�;(��?������q�)�X��v���=�A$�uAg�i�������@�X\/�J�<4'��܊zDc�f x�'%ͧ�s��3�5�������I��r��j?+K�̚{�S�Dh�����`v.G�h���LkI�(D+�3G	�����"6���L��#���,^�Ӡ�q��,�Fi8`�q]�kƖ�����V?�ɞTw�x>l�<�;	���>��K�_�.��*�H9]�7U�V�3�V��`���cw�A��W�8�� ^A��%5�����;�#o��;�ү����g�請V��il�Y�E� ] r�x�TR�F�FS��5��3M�����؜�����=�ˌ�@�|��r�f6ƹ���i�r�?<n�v���{�%Fr�8��vFcg��䜭:�H����b�Y�@�k�NRfb3EW(og�iƨ�5��֖6�����P߻��
�>K��(�r(Z�:su�l.�z-�H�H+���W3oʍ�"?t�_Xs���g����F�(�QE(< ��/F�Fif'
�gv�i6�H]���^����+_o��V��0j8�s�O1�6����?�I�P��n�΋i��l]/��j�y���0�(p'G���Y/��<Ⱥy}}Ioo/"��� A ��J����<�gV�~�P��P�g��KaY�z���F;2IX"`1�,����|���%��ͣj��L�{$ɭ�Bp�����rj�]�mVi�}����!�L�23S�d����,59yƈ�΋k��XOFd���Nc��!�EQ��<g7f-u�h^"J�R-����/����X\��"�aJ%��솬�&���I�>��;d8�b!A���('Z�`�h�����yGp�G.����Ah���o�]���-�M������"@s�����:��|=���x�Ձ��$��˲�5�4W*�&3���\R^N��D5�� O5�����H���0�܊�	vG�[^�	��w8��;lP-`6�����;���A�Vw���fvP�۪)�w=WJ�|<(�9e�~�[�"<qa>on���nעó+(e�omxW��:���=KSٶ���\m��w����>��	Y�v�Lɛn��XN�]�9Xc� ��3L��f�\��8c��;�	`'u���5�Xm�Vj���y�fz��(/�/�O���w��s��'��׬����Z��kr��X2�I2�m��eAr!�]��?�8�S�L�<��sP�<K�.��1+)���o��iI�:�<dlv�s��t,� &{�� Z���2���~�L�:(�~��"�;ȵS�l쬪q�/$�f{����I���Ljыs�d��4��GC�큥�|��d:�Vp�{Y�k�\�������XS�a�����h�0�X�1;T��]=�Bx��>؄�x����1����%v�'p){�)|�
���ğ8�G������K+���/b����ZL:��M�{8z����4���l�C?x`@�3�=e�y�����<�` p��ۭ>W=���鬡�\����7�Аmz�8� ����|�����f�c<D�=;��;�_ <��E��^��4ڸz�cJ�;�H�@��;���VT�]ߦ�on�a9{�ȵ~�/|L]��f�v&��m�{P��/�Db��Vmn�-&#{�I�,�i�L�d��n#5�R�1Y�o�����d�v���AE���iТlCD�}�������lt���5��?���߽]{�>+�����2�f4u��W����̲��{(�G0UNe���\<�].}c(��1T�H�
z��0�����qxg�����ƵN,�����m-%֮�k,���M��W�\�RIջ��3���97�[���/Y�z"���t ��k���-������p*��f���iR�&i�S+����6ݫ+KS��Q�\լ�"^�K��?�ڟ��NO0ߺ��̘���=�*�eA��s~xz$����L`�m�FP�����oi��j
�nt�;�3���@�_��(`-�*�+�L����q�ӿ�M��A�d<i ���v4���yVe���KꜤ/ݳ|������m��{+kKq��d$qrp`�}����ZKdΠU�(#o3���:�6{����H�j:���������@��([�c�i:���*���00�<OO4��}!c��p�M�d;=���^0�7<?Ҽ9u�}���J�j��%��U;���m�t��NY'�7^ գ�����/	�c?=���U���I�f%�����6/�k��ks��3^�PPA�_�:o����s�����{I�hp]��D��2r�4��j��3��I������9��r��̹Y�?��)'رmI�g ;���p�f���u��㥛?ruxD�{da�͋l�{@!׈f�T�>�������m�p4WG��B~���йY{��s$�� ���eK��Q��  ��ߥGʪ;��y�uv�ƝD��{��Zf�5������WK�C�U����؍(��9�`��fS�q��\��)Ϸ���gߛg3��<~��{�~��<����$k%oݙd����3N�D�����]��AO޵D���{ɰ2�=x����Ec����Y77%�/拁L��$�W���aR��z5�O��'sr�-��8��(�L�:��� {�4��a���ހO�&X�Ț}��8��;f ??~J����OP	����������H���rK�q��.j�� ��g�� �<���p�G�f76g/�&��]C3����m��I �q^C���8�E���3��މN�U�Ѵ�ټ�ｕ {f�����^�\�#+�Es��۰+�Z�+���^���Ҟ�����5����; 'q��zҩ���q�
w��q~2p��|r��@y喖ܰL��;4v@���-�+R��e
��ol����� [�ʩ���"eEje�k�_��^�������ru�ٲ����+ط(]�5^�8Zcڠ�?����!�&�Qw��|���{G�_	�\����z�㻷8W�6�g�l$6"�<p��!�
�6(-�K���3�؅N�;$�,
��쳛��eھ��Lw�]_é.n��J��Q�����zc;�3�w�={�+�F�|��1wke@�Ra�خ�����B`�r���)J#�\ί���nAΆ��n޽�@��KuA|�m���S�8Յ�E��x%5i��
��7/ ��&-�<��2�	OiB�T�J�`���`��[:߾~K�o[:Σ�N;Ir�9e6�!�^�����6W?[3�ls��ٷr��Q4�jvG)�}.��G31�E�^�<���n(��<0HPr���<�O�UjH_��1�� <P�NhY
E�ޖ�@/:��D�����SF��� ��V�:��]���@�º��]���́#�}۰$8q�O$MF�5�<�����3JʦW6�t\�� ���~7]��@�2d�xY����`A$
Q0�p���fw��d�gx"��:]���x��@3�n:��o/��o�p?�N�<gQO��IѺH&�a\E��]����*+S	�p��8���o6N��8{kR�5+;��=��:�tܔ�Q��n+��ߢ��@x�@/��(�0h��U��5�9�&Gܡp����9��ǁ�t�ۨ|"0j�o��;����\�L�!Q<����Ֆ`���[���|�W����~�:8Rȯ�,�2VYT[Z��:���k�1�P���hs�~�.���YtM�\?�U�f�J�{뚮NY;>�u�Υ�o߹��1]�vN���_Q|��~�Y6�2�e�kqm!�Y:�V������}�{g-;�WV2JuAu^���
Bun��<� �����:�#�9�TI�ǘ���۲����}����Z�k������3v�D�)@8�Cpe˦��'04X�N^�[����@;�M��.%�Ν�p��C��<f��xon�̧c�&r��w9b�4	p���#���+�'������9K�L���˅��dw6X_�R"����]ٳ�M��܆�E��d��!�\�Y��o1�|Y�RCKv1[�yN������CWi <����Z)����� ѽ2/����#x�����w����8��o���`N�O�!�a~�?~e�h.yg^,F���پ��t5�e�T�`�:��~�캇7�5��Z�$&j�ݤ��la�$�g�
4�!���u&
���q �T�$^I����^�^G��)d �^�`���!G��36K	�$V��(\:~�e8�7)օ�B���*Uuײ�l� f���V��f� k��fD�u��L.ܖ��Ϯ�?s9{��J���c_��
jd#~��)�%����E�4��N�$����[t(�	���x��7@l�?���$�N���3�̈	H7C�H�̲l��/���X79f����|;���������ւki�w+*!9Y���h��jqn�Q�ȼ��5�V� �
��(�Ӯ(�$���/������s�3ըH���3r��4�;�~��)�Q�A൨��9���̕S��Qگ�qz����4�4�Am�2v�|�c��e#��8(tm n�4u�f(���ǜ��{l�|�(�4u�A'^2EwŔurΜ,�bZ�2ze ��%�gi�ك"F���	��3	_w_�?��w�b�nѷ"���ty��L?����I�{m�~�;SJ3�Z ���t�'S"�v��ػt�!��A�yT�qD4��t>58�,�8��!��L� ���WT��*���:����3�n�Kݧ6o����F�b�~�9��v�4`:�͑)�e*��!�Ә��@㏐v��.�|�����-�z`�l 9���'8��c{��-�'��+^��g'#��O���,���צ�l(��M��Ǘ/�X}�b~(Z�GTs����i�<O��@�j<{�fk�N����n�Af������gI�k�:��[~��R��3u<��r��s�!؂��1Jas��Qӎ�Hޛ�� �`g����V�/���\����Lr�p�X�%U����>��*��_�5vP�{fg�1�"j���\�n�#�+��/����h�֘�Hpt�I>E ��V�ԁ]��	2Y������q<�كG��>��Ë�S��X�&9�H
9�g6=�9h�]'��a�cz�l�;u��y�}s	άb`ծ�<��]Q�z��c�e�eϾ� Tʱn.������1�D]++ǎx٦���:�%2�b�=��N� �U�_�οKJrڦm��g}����Z4�Z������fN�{!�x�h��N��V�� �2+��g�����˨�i��n}Y鹲�TmPh�(�$�'��; D����}t22n=KO%=r umj԰���1�z[��gWXf���XR��`]ɉ�� � �? ��A�o�'�FGe�`��<?�>W�⑾F�.���]�F�+6�1����Y��U�����'w�gJ�Lg+��Zð7����������Vj4��Z��Ԝ(���	��M�A��jcY)Ÿ�N��ܱ�,Ya�>��0�xF���0�cg ��d�r˥xg9�-K�48?P�2}��f��3��:��+�h�w�tR[���g|R�SP�7Wr��R��r*7.��K�L0˖ ��U����5	�}��>�K�X��e	��g�_�Olevέ���	c��[Q9��_���Z��+nԜ:u�9J�����!�蠭�f��N���_��j?�_^��n��u��_�;�ޕ��<��8�㓛����.4�E�t�jjnE�`�.'a�,��5��+)��"� �c��x9r�;��.L��kyr?�AWoF�?vN�h��ָ�Qo"ԥ=F���/�;�;��N���u������"���9Up�A;3���T�d��^�V���$�(B��T���l�� �*�Y�KMO�K�֎Ua�_��'��I�P.����ٺ��'�9ρu�c���=:���р�ZQ���`�OPΖB?���(W�Қa�<�4Y��؎̚�Gv�ƹO2e�)sm�t,�<vkQ�K�p\T fN��LM��q#*F�Fљ��!(�ZuL)F�* ��9Șr>O����ی,q�.��-�#��Cd�	/�G��t����ۍ�t^����Qu�95��o�b�i�h�|4�W�s�����E��#=�m� ��E��3��\ok:�@�w���� �e����^��]:�
9���t�����%�~ۈ��_ ��*�6��e2;�)a��:-�r�]Y#�S��wJn���)ԸU����d�:���ָX��f�����^���Jշ���ճ���ʲ�<�ey*9��hǖD�� �߃��h=�Կ���,�<�,���Qm
q#�I:n�LG���daIh��b�G�
�h���{����̡5��X��f����\'�P6�t�e����~W�,���w�E��e�fk���^f_���xg����ƚk���j��'�ˁb��.>%�� ��z�#��`���ɢ��k��8�bnѧ�d8�7�Q�Gɜ)�q��61dg�@�O:˙��ld��͔��p�u&�ʜ��y`(FEZ�0��wf.�J�[�~��r6`�H��ygm�j*�P5�D�	�w�J�58Xٛu�b��K��by"��m�*�>�q}�W����Ϯ>�]?�!��%Ǜ�� @��	��/�/,-����`s��h���u,�C�?�	EЕ\r��"A��v�]CG�x��&`�`�ĉ�"xr��6>X,���tB��Q�@?XI�]l����2{�,�e��	@�^����qdV/�9�b����_��{zz~H��-2]��g%U�l`�^�����c���:���� t� G��4��8�7h���s�<)����jY��]��]ѐ�}Ge/ +�}�ܢ�/�U
f�}m	���cs2�g[﮳*wl1�_�u�BI�� CS�����Y���`]+q�a��hע���m�)%���	]_Q3O��bHF���C~�y��F'>o�?��>������y��"�8ˮv�1uV�� �\:���g`��-ӭ*��ݭ��qN�=G�n|�\O_�+�g�ߢ��go)�,�Q�}g�߻~�ى��/kG�"��!X�D��L_.���Dd�}��������3|pqo�����?���[z~RV��z?	����v0�]��e��s;Q�Z{��=�+���ݛ��O�l»�6�I�"���/ L�h7~J�f����'� �r�{����aBm{^��w�x���b}=H�E:|��Z����U^�3�8�[Cm�Hq F<''��$�"锪�r�a�i:wg�������p�ې�qN�,�(�H�Q��"sJoFW!,�ǳ��h��v��,�3��o��fc8�(p�8/�Ț����+�k��r щ.Y��%Up"A�ǌ��a�	�����L�?�"�b/:2�ph���;5����g��ֆ+k����ǹC��k�yy�Ce�-p$D��4U�I��|�+�Wɜ־;�-s��~�hZ�g9�#���2�p�ǧ;K��L��zˈ0�atz���n{`�׺\��f�u���H`���"����o�-��͛�*�� G�dR��	8�n���f$�����Dd�NI���-�Ti�a�A�,֞����lM���m�/���5(�ٱ N�SF�8���`�
}���}z��%P
 dRev9��;L��pʌ<�V�4R}]� �N	�冬izB�D{e�S��0��>-}�ù[*���m��te�����#DR#t��Ͷ��a�Q\��w�n.�ޜ��9�u��4�ul[�)��0Ù�q�V�����R�E�G
��34=�ϑ�gf�y2���T� �q� �	�;������%ˆ4��F&�S��|�AP���O�32�uIf�c�w&�:#Ϊ��ى��ÅwAΘ�������2���*Pg�?R���c�J����w9)��82:���w����bEr{����:�?�D����@�@��\��b�p�uc9���%p	�Z�V�}%Gf3B���D����h9��:�~���#(p�)��ٖ��j�$u$3H\�8����|���Y
d��6c�UB�����H�P���}C>�p���=�z6Z����-������E��Z�S��Pe�n-#8b�����xo�A��x	ࡻ�+���%J�ٕ�e0��eDb��(=ZO��C�E�����&6o�뗯������3S�<Q=�ӧO������������єN��T�N��7���Z��_H�m3�t�n��(����ˡ/�i��o����~K���1]������x��i��2��f��� ��+blם�c���A���5��Y����3� #�	͛l��b0��C��ԍ5���w%͚��� w��]Zl��}�,�Ű��C0�\�Tm��:�K�H�
�%�aɬ���-	��j'}��$ٴ]�;���}rL����zMu�]���Z��D��N��g��t��+���m�L �؜;�z�XfY�.�/|�����X�Q%�f���W���?|��&֔�@�q�I�캖v#m��	�V�0��s�7J�*fS�b�w��]c݂2W>�"�x�B�?w�����,��׋��3�]t^;�"Dm��9�*q0�Idȓ� ����������E��X��l|��$���рW���t�'�z��$φa�M�FT�P 7�f9�?��
H+���-��lSd�L �R��Ԛ�D!�Z����fĒ�x?�67^k���p���8���.�?����bgF��7gȘ���݈v������r�����d�D[���Ԙ��<=/�ܽy-v&�G��me�B���-�0�j�w��;��Y��@�1�#d��$� ������+QI �Z�z1����ֆ�|4�����׺��Pn�|�n����fߢ� w�8L�ȷRT�?��\A$&1�T�R魝	�dY�])��3�D��_(md���PmsM�6ܩI�ͫ4)���&��Z�3��"9tB&YeF'��l�Y1Sa�
y��,���] �����c=X����o4^�1�/ ~��� �y��5��|��$p��x�a�r�+ʸ��u�}�ߙ��F�1<0WB�x���"묃����������6ۯ�Ɓ�i*1&x�t0��DʩCu���.Q��b��<kK��Bз�8/HF��G�kj�;���vU2��rsk��>[g�F�K�i�>��,�mdi�gX�1fـ2����ųv���#�I�уw�d�K�N\�3���&y	d����L����X�����wE�yP��Qm���{��[N�a������et��ַ�J�H�og�]���^1�܃LX��?�5�_w�+ �H�Kk.l��8�J\��]v��i�(��H��#��eXƟ!goE�%hQ.bvk�\���K�W:���.�b�zl >^��=*��7_������H9�������֚:d�{���L�?��g�J�j���Ug����{W�Ц�ҩY�^1ɈCVv��]n��ˎ�� j�Y�y��IV)M
~�|���_9}4�W�9~}`�x7&eJ����%�Y�eV'���]s�Yb��[y0Jw�U�R�޲��	*�l������4�?�������J F(����u��[�2�J�3��������&�����F��8�XξZ���D��cd���*)�@�+d"Mv�a%��bA��� �^_�pz�<�q��x#���2vF��Mt��� �j��:*#SU؇��o߾���Q �F# ��5�8��N"HN� _���We䞱lϷx��gN�g@� �y�#3��M�wG[�@;v�2�� *�i��:ZP��GIk�����x2������>W�;�7䃜lʻ��t��9�ܷ,���џܮ�E.�����#?�y��vYɐ�W���j��1��}$K�����]�z�R��,H0��cC�y;�f|~t��0�]��R�� �|�7�w�v1�����'-���0v���u�G����p��8����Ŵ���m���������-�zJ�/�2ΧID&�{ ���RO����������L��CzC����T�{�D�1���/�?��[���Lәq�R�9��A��ϓ����""��+�D5Sf@�%|]����,�.w�ڦ(g�[G��J�n�T�#)�X�Dx9scdќ�Gζj����������T~N{_Rֈ@�yb���y�������"���(�-�j�&��}���r�;��͎����l�A{�<VB�`D(�5����Y������g��_�S�ǋ�<���;d�S�Sͯd�)�Gs�sf�� =���"��h��>��h��z2�����S�����M�Q~���/�)���Qk�[*�rpAw��_qy�đ��I6��)���="�=�3T��9���FY�}��D�2bH?�:�~vs���GJ���G�&�cxݳ�j?]É%hh�
���m�rE��\�����#\�l����J5��"r��"N�Yj�-pG䉋�����c��;k��;�Z�:��op��u�N�Q`Ϣ���L,�Gv���kYP;����7���gV�w��o����7��YK��ܐ[6���q7�{�sq�k3��%�)@B�ELc�0�:ˮ�@�ȹF��_�.!�0�)ozoz`_������u�t,��� 9���V`'��􊲤LL�ѳ���˦y��R:?a��;v�,B��κ�R�k��d�]="H�r������j3�������׍�6��N��J�W��!�3�9g:��Y܁^jr��9�03uh�tg�9������L��.�͹l���b��c
�b>�c�3���A9�w�iK�� ��l'/�,�z!(6�ٖD����2���><��R^�̣��\$�l��7���/���Ƿ���W�&�]�f(��sy��q������k�����?k���4VS�G��FĽTp��-2Gw w�e�.L�8�Ͻqs�-����)��?�3��������R[�����%�/t���#� ��N��C�'e1(S������.U:��W���`�,���s�s��I�>��x<;k�>��N����1�� 	:��?�D�@���d�!��_Ƴs��\�j��������0 ۪����t�o��A��lt�S�I��������t�G���J��Fa��z���N(��*A<b\�h�޲2�/n6��?���}t �ʾ¹ ��F���D@���^JY|#U���<��Ӹ}��̬?DּPv����(�{z��>���sQ��g�T�<��Wl��R{�L���q�vM�8���k�����~m�����ܸbMN Λ�/� ����і}^\S�A��ߵ����\5��翟?��s�YE�ʱXZ�	{F�Ƽ�>?�����!-�������_��|:o�3w�ސ�'�^p��2���t�]�^޳!�M�逰����R����+ߗ�֞3���"f;�I�f�o���J؋ѝ���heV��-Nx�?�#��`�r��O�Kq����f�vI"�q����5%z���s{�� �5�v1WM�O%G��d H��f$@ћ����}5�7=%st�v˞�L'�j�ŕ�#k.[)�V+d���&a^�_i�ޱG�-v�)YcD���gҲO���ύ��_۱��S�~�����'*c���x= H��5)}����2)�|��3l�i����_�1��ʒm�I���e)@�r
W�F��/�i�zev�	�3��ஓ���I�6ȁ29�ӵ�~Cf��]Z�;���?1����erz�������L�9㤞��d��F^$:Lٌ�-��;�x�2���eƽg=���yMY�d�!5�f&��Ӧ���p�X]>縷�=�X�7w�59m@%�O��n�`>x���㤔x���C��I�!��G�pg�� ��#�9��NӘ�&�i�)�7.��+��L�[�-o:s�<��ůcyKh `��k���+���=5���x����=����'H	�i�� =���t<�K��M]v�����uY���W��Y����<:�Ϣ��?�řM�m��`���fw5]\ߵi��*xX���%���}�|֐��2�ڦ�^pՓ���k�\Ov�l�<m�*8��M���|�^����r>o�0������7U��D�$Y�V�
�|o�y�$��=_C RJ񰓃j�̵t9�K���̲n.��lN\��f�_@	���v�jtY\p=C�Ӗ0�1��\�]p�{%ѿ�VJt�k/��,CxŲ �����vL�^�*Y�lĳ���~ϞM7��ƈ�Y��Z����V��x��/F'A�c!@g�<	����0���鳮�'�$���p����E/�G��+r�<ON���Lc��F;�!i/*���u��
������5�k
:�a�/j�l�2Q���-L/\?�b��_�A+�Uf��]�����~�,(	Ee�T�}`F�"-;e� `zbY�5�'k��f�*f��4h2ՒM��O^�t=��>�;9�c���Y3�N��ԛ�2�~�NR�G܈�}#�3��,�Rv�٪�c�\M�\�lC��?�	�"^B��=�sge<�s�܃M�l�,���^ٲ��
"����f�:�W����*-�i�k�Rr�D�J�/o�bЕ���&f3�}xB� h�z�Щ2%dKPm���;�����9�?�Υn��.�`�?���'?���^7����NV�jpF#�l�5"�LL��x-������+�����TӉ2��^�����-�e:�br��Ӄ\Ȁ��ĩ� _^|I�Я2x�B�������|�B������[]���%��P�.B ��5��|��ӓVx��u<�13 (�,�%�#��p�=K~�i��Ͽ��g��J*��&G6I�ݘ6��Y�����U��a�#��g�X6�=��<�`DhI-��^�4�0����m_�H��i s�=��;������Y3�g�?��b-��/�M��k�{kL��<=?N���vq� p��h��W��ݳ2�@֢O�~(�Q�"-�7Gs}c<��{�W���%�~"'ϐ�=FF 8�є�Q� �*�x�O�w`w�����������{���4�J �
o������.'u"�nU�^��A�^%G�{o^���)�?�)�D�}�M��Ȭ���s#�T�5+K��擨���ON~dD0��\l]%_4�O2�#=̓� 6�膣v�+^�q�������5m@b9����24W���sz���������'�������༆D�tKI���nο]\�i����:O.�ޮ����2tLη�8����g_��A�6&b�S�ѷi�ޑ�1�k�
8�T��a���,���/�,e�s�'��v|}߸����~?���)�0��k徯����#IYS̫���ͺ~��>)v����z~,�����k5�Q5kf�Nk���y�+�r������g��`U�/~"KA�N� O����H)�2��<�5i��esov_��?���[s9se�3n���h ��E�z��v��~��G��,X�U��r�?���'�#᤾�l�BV9�Z[˞�̇�GJu�n]������n��;M��+̆쒵�����G��aE�7�F.���o�s@���%��˼u����L����Z��wt39F�+E{r��L�᧕�0B�Ѹ���=�ck˳��(�w�*V�ˇh��~���U֜q�tɜfeX��?3��,�k{e����#�T�#��e���}�H����n$Q���ˍ����)�A�s"�>q��-��܁w��㼌�6��i��;K��vL�U�A��D���뼪�9ߠ+O�y����Z,�nN%k���x#�V~���5�R���:�G������K��[�1��[���	�>����)>C-����2�4��f�'�R���WO�V�<L�>��I�8}���?��s�T<ϛ��X�2$�������inm�^��_��&���,r�F�D�α��4����$g�)yh�&2�>��4���jBW�����S9�Ztb��yOb)1�7'w��0h\�|�ڥ���j����"Zw��Lc[i���h�b�Y��Ѫ���v��͜1�Nug�=����=��G!�2:�9�ކ�Z�,>�@m��!���E�h���T���.��q[`B 1�i��ɅBq���L�sD��x�R��InH%S<�����,��u���cY��3�؀�Hɱ��h��by����R��Vz�7	Jj0w�����Q�;�.)"ռ����h-�zH�?}��z�L�����,#���-9�g/�%y��֡)�u`0 �V��������s.|�A"Δ�k性��KQ<:8,���R"R˻�$א�3�����W T{��L��`L��,kI����z)V��E��b���ډ;/�#z1��� �k_~��C=R���õD���T8�f�{�<-:��\��:�ln7�3:��1���y�E�"�*��{D���4N�,X��� "��������~�:{�=[��3���Rn���{�o�7�R3�d��Y��p�2l�f�=�WD���Sjfը72�s];�����Xk��X�C��<(R\�و"��IX��ղ:7�kv���`�!�~�>e�vv�혷.�`/s�:F�_�x"߷�q�R?�V���30>7�ί�%���n�5c�?Bn+������n��{s���ydF��Q͹Z���]�k�T�*�=yV^����N:��U�7�A�=���-�C���R	9ټy�ό���N�Ϫ\~2����3{�vl�ٻS=�~�A������.E�1�{4���MD�d�`(,�ap��������O������N�,�8x��^V�=�L�jp�����`�e�	'#M&�	l���� �|O�w�����Ё��鉁��vu�4�<�q���R�/�F/ś/|U�.ʗа����-��Y6.�΢�f��㣌��5�dv��W�:\���y���F9�X"��Q+r����J����}SY5�juA�]�u��e6r�;c� Gf 7�&��Og����΂*A&!otzLa3��P{�x��X��a�����#J{It6�_����`�ya?���	f���v=V�?�M ��]Sm���(�{6������
��ܶ��l||��B�c�f��̞m�u�����w�/��a�I��s[�d�*W���XZ�Jq�\��g6^釷sW��q}�N�f1���Ai@��KS�#�_�|a��=:5=>��I��H(�$�<���h�w��g*F�C�䜫4bm�`�={��l����Mپ]�ϛ'nm�����-�R��y���H��=���D9S����^�q=�ec&�O�&�Nqs;��U�3v*gD5����s+JԵ�<E����\��H8o���ζ-/R�X�ˏ>�Ղ��f��A��=j��s�OEǨG'0��R�j�K�&��$�jqQu��|�j�9���]o.]��cV��ύ��6��@�ز2��N�g`�cM-��J��Ǉ�����uv p�t�c�u������e���9*u�H"\[ۥ�>�?�<�j��_X�c8b�Q���D��1Z�"�����T�i���X�O�@�;�5 S����H�) ߏ�0����'�1y�:1]�3J%>Y�������Â�I����8�z���f�h^��(KM�1�eO�j�d9[��}L}��=�R�e�A0�:>"���Y%�r��~`��=˽���6��o���������>/��ѲKy/���\���=���k7ٸ&�=�"�:��5 �d�.C�T{��DǪ�\&��}�k6[��F;6Fn��`�@�CR�
����y��/�RD����;�cg��>�M��v�c\��2T�pʮ��۾���׭�̊9�W�`�.���x���y�<���� �?2:\�'�{��=���-?�D����V�+ɯb�L�uU�,�a\��t��^��:�;��Å̮�n�b��R�7뇪�s:�3���ʇֵr���.��������+���{I��-��]���|��4�_�]�;K�$fYb>ekU���?��ޮ�u��#ttʔ�,A�'K=�j�Z�lx.�������M��$�F>:�����Gg!0���?�F΋}@��'�^An&Y.����<L�������`����
k-�Fsw��m��-�cdO��}p� �5G`�>��#�2�#�S ?v����z����fĀ;uqώ��&���9�o��b��}��dd�lO���A�=�}c��5Yc�<���_�J�t=���o�n�R<3��@f���k�;��'���q3"fd^)Ki�.��`�9�l_k�{CJ��`�R����/d���;�#/�]Zw�b<{ʂ߉8\r��Q�{2J<�)�D]3�r���R7���ópr��[Z`�8�Dc�$������@����5���ir��S<���@�읐+ef���z�q��5�֢��n�b��ď6�^q;�����;R$��C���
���]2*���To �h՗�۴���\o[hK9
��ŉ^}���a�_j���m>�������~o���a^sD���O�@��d�߫��N-�!9�m����iG�צ��mfCs?��o��Ӯ���`���>��-GR��]�!Yn^u�.W�>3H�'�x�T� K���Y4�')�=��* ���p�ϓ߫ ,��♐՘22�Ƞp��F�ݴFF:��s֜��qD�HX=�,�?O?ݤ�{���߸�>^|ףn%y�=%*�I�C���'ŏ��zN�&�����v*�����R�A\���*[��p0R='���=�;�@���'3P����5���F6<X��>ڱb��R�����zE� 0M{��C��k+�� D����S:B��̼Q.A3b�Q9���\ÀPg�����͖�����s O�hN�y�]��A����blL����,���ж,;�S�lΫ�!����܇���������S�Ƃ2���W{�����W-+;f�� o���k	�����c��������'�&�c6 ̌1d� ���fk�B=��F�-]`��� m����V�n2�+�Y��ި�vn��XҞ�������t��:�Yύ,�d��`g���Ǝ;�9���|��֏g�9�1����A#Vu��3��wsJ�Vֻ@��<N�Dd�ʜ �\>��̂��[&��w�r8���Jgr�	.��jnĔtZG,�����"(�hҖq]�Ν�����U���rϚǿ�ք?#�����4 p�VK�:�^���w�j���-Mכ���/���m�W� �<�e�c�w�4w�30�����.@�����������4��K:��h��c�{�(c�	k-�!�Ʈ��xW�d��Ǔ>A�frP���Zāq��+ceL)��SȬ+Cc_����lV6�<��Y�n���O']��H�@��П�w�a���^�=���?J��Kv�C���y�}�n�~��3��e�2�j�zF��喓��Uc�<#�X�O���3��ŋ�㮶�V��u�ѳuHt H�,�b��&�>G�g6+��<����:���5P��>K
Ё�<3� ���e/��s�){�7�m%��,��k�J�ʛ�1stŭ�W���@���q�V�feR��H�68�Z���"�/�r�q�o� �a(/���'fG[&;�����1h�,�u-�3�J�*d1�dD�y���yG���b�*.d��[�����Ȱ#fgkty�mѽ��c7V޸F���z>������E�a˹|?�56|;5hd��ӵun+��W��i�1&����z}k1��_g Տ<�˃�����!���Ft�ɱ�ۨ��h��8_��A�΂	��ϓP��l�;�-�<� ���-i5->'�tc���ܺG-�z1䶤�\���"_�{���X[b�f�Ӧ(�ou$YP�K���}���(&���1ImBύ���`Jyj:xfL���ť�;��[b�ڿ�5#.,����fG�Qw��VD�S�V�gG̥���l ���j%���DC� Ř"�[�N�[,�,F'��_��zB�I��.�\��!�_n�=[R�E!�}w��Ⱥ�����«H��S�9�~Q"�ýtP�F@W�;������ٳE��Y�/2, �����n`h��ks���[�ΊF���vKb�Fv�(�j�O���;�	�'@E@0E��Ti��td�mMb[����o��J9Fz#�UW��v�c0F���ߏ�{�Q0i����4&����5�ׯl�y�,D�N2n6 v� E�a��)�N�X��}Ntv�a�h;Q�e{1�-s��9�ee-F�ٽ�"H��:V����0R�5�;[���s��t�v����A4Ȳ�a�|ϝ��Rt�BT��%J�6V�~�:�5��;"�*CE�:` zF n����!�?�Ѩ�n�Mt�5b�ƹw�3۬��P<��	p��b�t#;
ƴ��%��*;��G]}W�1�L������հ׏�_�'g�2�����j�\	2����X�Y`!H&�:����]&Xa-ͥҫ�`D+�J��s ,[s �\�"�-h�:A���,�h��ܡ�����9�c�Y��2=��ʖe�]����ED���q��]b�i�_/�|N�5s���j�Lް��k>;7c.���P�>nH�Uo�Q6���Dۦ���# �)O���;8@�:wvZ��_�3��[��g�ە����٘��1�'϶�����ud��;Ag�_l>���w{g+�}�I�?��LF����o2�OΟ��C��*���VO�d��Wt���=�ن�<(���S;r���2��K�;M�:_����r13��U ҚՅ�@6�@p ��=����PI%d%� ���}�u�$gّ4�
�����S%��s���8;ל����`��7{#��Jb�%#���&���=�,��7|6�1PeG��c��~�Nu %�~�X�g���v؁R�.�9�$0�rЪl��`�	� �x02�� }t��x,�K�� ���3w��x�~�6]+��%׵�/[� k�,�>2K`*���@'�f�QYtQ*�5���)S��RT5�1>}�\X��[R�����&��^	��0+ʂ��cVv�xl�ݓ{�h%f]��5�ϩ)��h;[]�Z��r��i�P�T<{�T��̎Q��y��Q�5^�&��y����sr�^K�ԡn�\5���(j��dVV�ϡ�d�����6;�����L�X����k�9�d�!�x��c,�жj	8�ሌF;�^H�g��op�ܯ��Z/�i1M�is��Gs�Y���AC��v��	X<�9�c�s�����H4�_�Ϸ��������F��R�ܔ��V����#�9�ƒ�R�s�ǍKNN/�3���gjߍ?}�޴�~u3��WZ���ZT'�sv�zl�.�������O��]� ���MG �xv�%�㗸�4���s(�����=�Ų�t[]��J���"�{�<��Ɖ�DD\���̑pGA���,��?�D�f�eIV�0��N��Ϻ7�#w+e����H���Kzy�K��뙊Kd��܃x2~"/�b7$k.1Z-��	���%����
��ܣ$8���3\k���ձ'�쌴�[kf������)){h������s�����I�Y�@*d�,�׳~��ܔ2�M����Y�C��es.�<v��|�VD9�#����y{��U�ݯ,X�T�yܿ.ҷo��kJJr��[W�az
:�ID�Ɩc'5WӬF[s�-��a��Z��4�.�z�a�����!��?)9�G+�դ�y��[iہƹ�غ�S� Y�+��*������8�;�&M-0��R���f�7�0otp���]��g�n��,e�O�޺~U>yb�7�o��s�& ｋ�V!'�Ϭr�V�Қ[5��3l����x�=~J�?�/�KÍ��Fy}��5w?��D�\��J�|�^�D	˸�n4gׅ퍝]���;����4Tno�i��\��LͰ��Vֵ����l�9��!}�������ÿu_��m����Ȳ_��;�S�n9>r '�~�grq5�C_�V}�*]��w���v�2��ɒ�pp�\4����O����陃x�lt�A�J���$��b��_?y_7wm��|.��t=4�e	4�u��5:[���0�V��Y���{/�O7��s�X��� �
(~�uՑ��et[l��{ټ*��{�/�(��ǽ����u|BP�$��=�#�i���ނAGf����%_�L^�}�C�Y�-3ȟ8ێ���l��sz��`vs/�i���%;��#h�2 ��Ԕ�:���[r���:�٘�A�*sG�;����3�<�����_Ӿ�lRq���:V�M/��h���@M�3�"�Уq��x���co7�~{k���9§n��]�On�hrW���Qz����a.��ZA��DT�h&�r��ٕ����E�
�Ϯf�g��Q��2jY~ev��l���#m �����_[�?�Wg�y�0?s�١`[(r6�����"���P.�y ���0��:K�^��F�e8�����?:'�\�;�2���	e9�g�>?"�����Om��'�	oE��(k`t�r" �`��ូ���|�76e;����~�K�P�(oo��^C�}�W%tB���+5�����s�"JW�y��ŧ�������d_���x^�c!��_�Z�@�	3�N^�����<�bi���9�Ħ�{��$��X%s��w���Ka�\�{�e�e��"����`��z��"����X�uH@K�t��bF	����^����qEPgpczAy�rnvd���e>$`MW�8���(�:��0ػ��x��ȓTQ��6�"2P�72;n����E�퓲�N̐IEmCݐ��O��|��  �r��@޻���ҏE���܎Q.���:c�d�aYB��4�id��W+�+x!Y��+d�`�?~Nϟ�y�V�����I�kǮ�gJ�:u(�ge[Ǔ)�}��-�vv��d���,�y�5��r�����m�  ��IDAT�C���S�v��uGe?��WH����]9iJ=�O���n���QRb9_�t�M��Ø�rٔ��c�yg�<O�Ϋ��d�w��a�U	c7��Q�0��6W����]��td�M�����<�*�heC���;3��!a�4�_��,��c촾m%��v�ѵ�Z���>��Eq��$M�Q��x�	��[y�}�e��K݆9�<`�%����+e����u(B
��N:�ꂵf�C�����q3�5�|�D ���*&����L�לo^o�9]�ָ�}��ō�0�/�W�r�-J���t#��v���Zf2u��ʗ:uL�N�� �CɽE�ѱ~�o���X^~%~+��\�Ѷ�4('_���;��Ћ^��&��Z�q��K��A�d���-�
�4���,!3r�#�����O��f�=߂:�Q<i�^���Ż3���Z����5�^bw�SϠ]?"�W���	��q�����#Y�4���Mu6��t��t��Q������.V&�t��e+���/��L{*��ejd}v���2_<����F����#푖A"����fe�'[/�����;�����n�,%�ԫ��Zޥ�{���4=��7r5��2P�����é<*�ί��6���J���5 eh�f�^7G1<;nl��߻���Ն�oa7�<V�# F(kPV��Z��k9d��U7�=[�VF�*#~f�O���'VM��E��J�_�q��4SiWݲv��.B��.� v��t7�|�&��ϟ��nPK@y5	�ez�V�aS�9�����s���/��VW�^��y-su�R�r�IP�޷�z2~ ���q
N�1�d��n�5'{��7*���L�{�9��z�h,n�]�r�t���|�3��6�J��DMVR��+g��Q��򼊫^�tr��D�5	��2��nJ�Z]��w�P��N{���)��\�Tب�B��#�S��V�ۂX��O��Wm [u��@s!ta0�|Aq�����K{�tÁ "2//�;��ݤ��@+��a9f�f�2��0E d���q�.Mc8�sg�:����ag�;*��rM�<�#:#�	�Z��f�-'�Nea���f|���@{���;������v9E�Rf�~?Yf����vUh�2{��:����T��w�:�@ݳe�f{�Tߓe
9Ϝ�[�4�y��b�:k�Gi�$'��*�¼F��AA�Q2�)�Nh�P+K��R��t����������i�WO�-���Q��m?=�m� F�z�	ܢ-���4���ǃ�Wq(\��	𛟟;fy�g�Xioh<�W�Œ�՜�z��1,�6��	�FT<�#�Ц��@�����d�����R��U����z��Ȕe�(Km�G�����>.�|t�J��ڒ�rU��e�F��I٩��i�t�?�@"��ۚ�b�,�>�s�S��v�h�Ek��D��k;�go�ήlNZ�j�e+᧣�R7�:,=XZy�ˣ�H�:��+�5��J`|��bNi3&��e���a��)��9�^�5W^64���s���}�c���
���f?BNeR��J������8�L���������rD��ә}�������b2�M�;'j6��m� @$Qo�St�7@@�6�	��u:��1�D�2� '��ѨrD���6]x �GU	ծ����1r5��ΕG�*�����:`�F?�+��:�l��	{�dY*P�g�~t/�O˲><>�F����(�k�qGЉA7�u��8Y�l��i+�&BzZϊccs�-�ߩQ�',�K�7ud��G�)�!K��l�XhC��t��r,C��N�-� �h�'���5�����+"%��S'�|Mi�s*v���f����b��CY���q����ms���&8Fׂ@߹Y7�v5:�_]8�u�jׄ��]LR�3�h|7ʚ�Aa�,�:2B���g�a�]_��!=���m��f�:vM�@eZ�u���=��=4F��m���0IB����ٶ���(guB�gΘUdvQ���kHA�B�^ϓ�>~N4�ǡ$�SO�r��}:�6�l�>8���/�收�z�1�u�V!�d��J	x�������V��m��*O�yٳ=v8����D� �s#��ŵ�t]�p�{(�Pk�?&�X��u_@rQ��V3v����맱�q����Z2�Xxe���,+evM�0�bB���gv
�y'�Eȼ��\	؁�?�Y��v���)���r����V���26�;qq��S�ZM��ۋ8��Z������_�ɀ<�z2���Ш)'�,x�N//���,2���Ⱥa �i�b$�j���7����:��H�?�J�S�dD3���@9�w��;� �GI�x���.�g���!A��D' �R�a���2�������� u@ �q�vQW4����M69� ���G�z˜q������������I��/'�b͟�\6�a�ɐx�l�9�1^�.f��u��k��ղ1�3Р-�ѪjZ����.�f�����n�>������ATv�vs���^�A/�M�[0��r�\�t��FB-��F4Ҟ��J�gi��m>��dj���hٝU�ҔL�����8F�>3�\^9 d ���}��R�lM�|��\��}n��U��D�y���Rs~4�
�csR±˖4W]t�й,y�o���j�_Ƕ�x�=���3�p�<����~u3Yn�Q[�&�'cs+�z�Z]���$�_������s5\�O�{������t���X�_[��,d��{m��N�%�q<����lS�c-����l�w�|,CN����XԽ�;Zc����y9��ax��~�u:9׾�8Ds�l���D}4��٩��{}�����x�H�`�~�rfi���Ǆ�`V��a��B��cn�GG$��$���M���F��q�۸'/�?J���Sd��Dp�P_��I� ��w�<YWKrmN��Y���x�-N���s�XX�1�g�\��� ��1F��b��N�+���ŧ,�AY�����9��z�L:5�P�D��1��m;�	@���B2�v̎J�/�3婻����ٖ�Y ű #8���S�ީӁ�7w��v�D�A�b�p��� 2�C��E���X'�w��'���3�٧�x�25����Q�
2rPr���7~���,����������I�����7�\�.��չo�ͦn�n���f�2�j�����:΍�EPj�H����_}��A@�$�\:n���ܢ�Kg�V.�y`*7|8.�o�w~�����6/������Ĺq��_�_h�)]���"'���I-��2_޷�[����g	�b,?��a�&e�3kQtt��L�rP�>�_���q�5{���׬���ɳlbx��&�6t��Y;_'!�ݿ�F=����n '�t��p�3�#��κ6
5-��N�Zs��_Gʻ�3V�{7#b������n,�؜�Q���Msn�4�F���sC��=Rn�80�V;-Õ����"�eD�7��K+0�qBE����ך�����R�۸�g[O^��Q^��)�Ϯ����#�1�RAL\��&%���#?��'*R �K�i�^ޖ��� [e6�>O���d��ǒ�IUtf%b�~e
�#����F�d~��_�S�,�A��Č*]�8����0���'�� JU�;E^�������C�Y�*A�8��4�*_<��פ��C/�dN�m!"E !$��C�]O���^[k�i^p�u�)̖��v���<�,�|eu_N����GH�ѕ�ϳi0�tod��Ky#Q��J����b~a��N�6B��F����6*S�[��u� ����~-c��5'��N�{�U��#��D�ޱ��3g�[VH+�9(���A؅2��~�e�0�����$/��w�R��[��B���-]qP��'�lx}U��n����Cj�������)��f�n����������.�R�=��T�|wPY��<�Ov�z��Y�:r���-����s�\��}��:�d��c�~r���Қg+�ҙC��%Ͳ,L�w=�v�g!��^�#Ȟ[2��<����6&Y�����?�izL����m����XV� �=r�(�NM��gY��Tdｬ���Q7����r�Y,�7-�su�������}f���]$s0��� �ă�Ҥ��˅ԭvE_f��l��lz�Z��˿E[`D��𺭒<� ���`%�n���L��9��tBx<�U�2v:�~V�\�l���Ï��#d�v����TЯ��>l��ٻ+.��>�,(�v��K�lk�%F�@�~�'�kXbA��\vl� �ᕲtMTƱ��,`6��D%��������9��@��~΍9Kgk��z�K�9��*�ߣ��nVK+}S��{�j7{�3�2��/����ܸ֟K������53��L���!�Z��m��+�ll��8�<����#��גw�i���#$A�b��ܿl�>�G�1��1��2�]�:2����1SN�j7n09V���9�4](���>�o_����cڼ�b7�C>Nii������r�_�M��ZI����&C�r��w��d�BÇ�=����,!��9����>_���Zt��bdJ+�6�G�{#i�����o;"T���'��Aq0���ڒ���! �m���T�JJ MYF���8vFfy��.�@�#�Q�a�+g���̵9�s�J#������6���R�s�r��{��A��rQ�m�oOy0�;2,���JۥxR���5	�"�Gs�zh��:,JUЌm7�q������!��L" .̤B:93��c�����B���{�������Z3$U�my-o�������ipe��,ƶ��a����Iĳ��N;��;9�.]S��F�I�(�E�
H��o�ρ\S�4��H���}}M_�~K��&�ms�s�/낒�A�uHC6���bL�����>���B+���STO2"x6R%2���Z��9짛y�)
:����Ď_0�[�3N�]5=Ӂ��G#ҫ�H�U�����ڔ�v�L�C͟k������yD��]3>l��(�aސ0;J�,����dYB~�v<���Ʈ�2���ۦHW�摕�q���v�NPu�]��4N�3���>�R�O���SĶ�p:�9__C��1���w�jd��P������w@�tv�3�"̌�>���=��WL6030w�x)g���\z||�L| q�@��*Ii�pz'�涓��\۲�q��>�%_m��w� sJ�u�Om�2rě:��S�T���ٓ]����@Bs'�B�a����Y!�<r���?�oJ�吏椩t��0=�	X\�fM��88��׶لq��.b���3�_Jaw�`&�eΫ�=3Fȹ���90����!��*�U�$�@/���C��9��L�V�S�z}�g�شrGv 9a�P�����#�~+�����c 
_�������1v��W�X:�x���yٟ|��r\��ʢ邳�����	�S�;t�ZZ�� �VGϮ�2P�Q�ʎ�f:��A��)8���T���:�l�ORb0�3��Y(��z*��]�0�xNi�[����e>���gI`�|��-"ӈ�4���7A�U�ԑ�U�R�����WZ��T��R���`�͕��X�E����ܵ5�b�Y~%<����+C�L�V)��f�����m����مz�N�0��$�k<���o�E�����>M��<&O�\�?O��1}}�L�I�*�p0�5��z��uR}��~ߍµh����ڿM@�ngwA�J;��l��d����V0ʯ�5H[�b[3~
��A�/�� 亡΄����YJu���\8UP�=z�?���E�k,V��4�[9����I�7��Q�3�%(��l(���oɑ� =�o9(���탎�X����<n���){K_ݟ+��ڃ���c�c7y��:i#�L?���G6��%�JX,���1�@elcR�LSR����v����
BY*�u�ǔ�T�ט�4������#��Z��ZZZ0�0���>��c�Z�-�-�$�1m9��O(޾?�~;d�`�/l��ظ��Ɂ��'#`>2r8/	��p��	
 ���}z���9@���۷���@���q����C!8"Vwӫ�����kz{}�d�͞��CO��������o0#=��N|Kc @�}Q�	N�x�R����oDE�!*[��"i��wZ�����:O�H��a_�#�U8j�ad�n��K� Bp�E���vL�e���۟h�y�����c�� �`�����g� ���惁Zl)��)d8ݭ�A� #�f�F �n�)�	@��N���@��t��d|#���r�u������y?�����a�Ӡ����q��Q1��� en�4(0�'X�ǱF�CL{$�ejH��謶��cRǬ�@X:�uX;���-k�$�FF���JVn����[��EQ"A����׶�x]��D��+u�E��O�3�4j����v�*o�3���hnr�v��g<��0۰�A2�K�jf�2�����6��Dr��/�K�̖�E�TR�N�PW�xe�e��s?�˕+S�ี�K�읺�k;�L"켃���BN#�zы�UA��O,	j�3��]���[�}��T�%ӥ���cc�Xs�2?vk;�kG/��I���g_���F ޺��J���}��n�w܁Z����Q��r\1�1����|��Iw~��:��o��0�l]+E�ȩ���9%k���#`�ݸ�R5�Yq����IcD�9�ȿϡ\3z횖K2A�$��Þv��U��ɎB���cz���Β��]J�b�qO�o<0�U<z
�'dw��p�ew5Pe��.�!�5.\ȸD�G�~f���p��<G�M����7�m�#ϒ���M������Y\���ǣl��f�^�e݋4Y������ӧɎ(�5 ��ގ�Hg�x�� KQ��w����9�$_��4����g�����Q���q;��-=?�2x�a[�����p�c�7��e�/{�e�*�&�`o`|єj����i�L�eR�[P�����ALf�AM�J?X������>�=n��NN��Ȉ���U��M&����?���V@�����i�g|v�������t��k� ��C �e���0S��m��;+�9�_��k�ʦ��m)K\��}��� Z�_���mB�g�̹^��y��a���{6����;����9ed����]���H�R�i�7����� �З//�__�N����Ͽ��ӂ����u����\h N���yI�!Rb`����W&�&k�A����T�Cd��|��cp��jD;�Y(";H��9�]������H�6�d
���,�H���1��ޕ��W3K!�H�y�k8��"@&���hIyP⃜��\G�-��}:#ɜ���YW�����4�����*8�g(qJu�4�����7Q�I�� ��f0"��{W��kgD�{�������{z�ܝdfF��,B<H���]��z:iT�n8^�����wZŠ�	J��T�T�~���h�!�.$z���Xӳy��NnonEC��thV3�4
<��)Ah�mo����!���4$DyL#?ߙ�MA�V���i;)Qj?h��HV�7^!)�`�� V۫�L�y��WMo������7EG:;{9��O㴲�� �..̰s.�W�5 ��T��uk�}@�����/?�����d���:W`����M����?e}~F��V�8O�yU�^^�����|�+z]�&?��o�8\�&ɳ=�jV�i�ӷ����W~�6�
u�#��@��a.M\�J�D嚆�>�a�$3i~�2����ẻi�6(�ř��Y~7ޣa�bV�_ƨl�y��w��E&�$?����`�!����S�p��(U�w4 Nc������w��?��,`zX4M�7D~�Y���;*�|ٸ�3Hf�?C�����x����B������u�����ϯ��Ͽ� 7�a��`%��������Ô�8B���  U�]��-�`'��.��0�:@RN0���D�Ux_=L�W�u�s̉�Y���ڸ��e~��G�^a���sG��S�K�m�$��D������R�֚�9�ᅜe�^	���o's5>�,��4�c-�{S������f�6/�ZT�&a*�#�EԈ��0�����u �xf��0e�M��6��\q�CD��0�Gk��\ZX�a��>�r�H���C�֑s�z4$�T�S�*R���r���3]��VM�X�lgcT5�c�8�N��}�R��H\���C�;F� xu"�@��`���5��K��;��RZ)��)���:n-}����d��0����C���A&����ތ�;��R�q2����H�73��?����bO����rA�PO��&��E,���<��q�M��K읝q�8�/�-Uĺd34�1iR�I�N�k��xN�ͧ�ʊ��g��3y~>���+��ng�r#����w�@�:&���4��j�����9��l�4y���S0Z-����烃
�����C��j�,�F�:�.��Jiʖ�PG��`�4��%�d>43�x�7��~2��S��?����A�6je0�q��nT܆߳x
U�ۖFVu�(­{�Aq�9��,
H"��i�3~z'�������Q���y̾�����vO�*���,�xvM��C#+����ZP���T� �X{��n$�3R��v�Χ�iP'$R�@�G�o��J�����F���+y�z�(��?�Vq�}����6�3���6J���
i~;bԩ�r��ݥ�0����R��)�I��I͑�������G�W�n�8��6�x�����d��Sf��g�F����S���\�s�(�kG��7P9��pZ�tκ��Ɗ�"��}l�9�����J��o(K���lfp��w��(��p�Q��u ��t&�|���B��]r�3 ��H*�T�|��=�\z��n������aKG�0)��(-��k�SUb"v!��,�/�@���{�E�7���3�n(����N@Л���vn�9��&��W�b��&rX#��i�)�+Î���"T:>�����q��Nu�AO�B��/���S�t�X�;�%Y�%���tҴ�R6UØ��[y`���+��lm#I�2������@���3A���i��l�b��[z9�B�����}�����N��Jrc��a&�G&?�G���Y�;��΀:��("AW���829���#<�Tn��r��N��o�{{M=Tn��9�iĐ�A�����jК�R�4�[:��`=AA�A����n��!�ى���E�hpD_�; ��nit�jK�au�Y{�h��D���ƺT�d�7�o�Z�r�/�o$�-���t��0B�����Tzg��V����ȨK��H �}���~M�W��Z�&��;X�v;Q��|���%  �5=�����͛rܰ�B��6/��2���lE��J{� Oӥ4�z��B�qk�F���>�s�%�e�j��3bF�ld=�
���É����^"f������:Rn��=�Txnl2��1��u�ϙaG��:) F�΍̨��{�G'�N,I3�9%t\Y��������ؤQ����KJ#r�H?�g���N��a2-�.��\7&w\��G
%��y'��
pZu�z�~]�������5\;v�����V���SNi���hiǴ!���efi���ûeB�[:V����9#�����n�7Ua�O7r�DH2�2ߵb�Ԍm1��N'U���Rs�E�N��q�'B'���N#v���?2�y��)c�Gǜ2�(�I����W�]�����goZ��ǹ�P���g�H�é�����Fó����Q=�ך��J#39mDy{&�K�>axй��D�s��3�W �6vY��ԛ�T k+�=�
3P��,#5�#��Y���J#��_qEGˎ��0,���y�s*�^�<;�X�VtBI��O���j0�?�8P1�FcL<�ݣ�1+�%j���L�_�-�_(�H���w��~"F���@�ZK�]X�@��0��gث��B�M��s����Цr&��Q#G����x@$KC��R�n,��U��F�Ku4��`�n8�!a�C1H��T��MS�5
JtH�2��|�G��V��hx����k�V.�#ʍ���++7(�������"��a�96ؘi�C������,jn��Ԧ�v�T�fb�	�粕C��+Lf�,P�I�vhq��z�"�H�� }��;YF����6�ht0����Am?�t��B�C��+�Z�|������џ��vۅz��fUߍ;��ϋp����3�F <nvo2laIL�y��Zh����zya�������KS6o��1d�m�HZ{[ F�6��1,��$	D�H֠D���T�^=�u�.�9�T�V��k��ng(���"�&���;�-lv�̍,kc�m���%���������a��L{��L�N��Q�>��m�Z�T��0LP���,��N��)��A�ZՄ�e��ܵP��*	�*��D����;�z�U����ϙ���).�y�`d@3�cuLEv?x� �a$��������㊊5+���3z,l~�h Y���du�^s�1����ܰÒ�g��k���%Du@p�nnut=��5�p2����H��\d�vC����1�7O�#�4(�Yp�����m��t�Az��r�p�k����aˌRY�Qg�3^���ձ��a�'v�$R��Ak�֑���c�^^�l�y��Q���6���n�䯌xAfߟG���:�>�T����3��|��"E^*x�ޘ�¨,��F_�ɶӴ7�\�W��G:0�Ѱ3i�9R���onVj�q���F"O��^�J؎ϥ)6���	�6����%y37{5�L�y� ���\h�6�W�׷G�����{�r�5M�F�=��
�������I��K��j��r��?�����9qB^�'�@D�ෞ`ZSAu[-�]S��r�dF|�a���܊V��?s���M�, �Z	����q���a�T��UF��f ��Ȏ����pE����D���2���_s_/�� �U�Sexq7�� s�Q�����~px[��R	���w/�����z�����	c6�!KI��0R�&��Ip��#�R�_8m$��l��T�0D������81�˴uf�V۪�ģw��}��� ֧��9�	�O8�ؚ,�?N���+������u�"���e�T\t-#>�����q�(1�*�(+�TZK�垝�תR��YD�*�b�ȑ]��ޜ(f�ή\)֞,�%�CO�w�r�T��C��#��=tuL��^��5Ӟ ����g	�- �?;��ψxėFLk�6�\�a �X�)cBO޷ܤ*o�P�V�d���Q>M�'�4}��f}����'�����!�%��{���������{��Î�,	�r`��n4%������zb4�WM�U9�Z��#�3�]`g�ޱg��v������8��ϓU&5��}��)�:0]��tXN�aI#CNc�qqYʔ2F�\hz���p��(����x�����3���(�3K�R���h�1���/��u7�x��rmj�FҾ���Y�F��e�ISP)�k����� �qǿC��{�&5��\ǌ0�vn-+�����ew(�F���aGyZ��^Ѽ��g�hč��x7���M�|n�� Mi�	��	2����,���1��� ����#4�	���·(�d6z�-�-]Y{�\}V?p��<a=����d�UF�l� �7�J ��z,~F<\�%�;1�U����!��8U��EHm,Yv���g���
��p�E9fe�Wf}�~���y��.)�b4*�4��^J%�4Հѕ1�f�r	UpX�or�g��R��}S�&��Ema�}�P!S= L?��"ie�d4y����W
� p�UIvC]J��x��
�Ai�G<5������]��//O�,`=�8 R ���3X��4��	�׾����;�K=����PZ�C��~��[���ɖ��z%������������E�;�:�=R�0��^�l.ΰNϫU� p����o&}y}�9xs{C����4�4Z�!�ҁ�	�Ƽ�����������vJ�,�+���\SP���r�T����^�`#�u���h�F��H�lӯ�bf�_��c׫7	{�<% D����-҇2�������(��Vƴ��K�Jb��̌))��0��^�6"�D3'��(4z��:�ڤ{6��yO�Bȝ���>�<����܏/�h/泧&���������,e�t)�.�/��Qa�=m�`_z�g�)�<��c�}�q��vK ��x4�Z: �~^;�w�k��%S��P,F�n���V���l�qE;�7��0;�5��-��"���D�d��F�o�h�rQo�z�T��`R�i�B�3�����fݥ��vU̠�k�ܞ%��}���no���Ӊ��b�R��?�#��j[^��R,��37�;T���3j�S{�f? �1�����x�DI9����RKܫ��\�G�U}d��x� @����\�Ȯ�ؗ���Vƛf��ط�%v�6�.�&����W�!N��1���峥y����u���O�,�k��\��F�&�i�ߩ��D��*NP����E��ܝ�<�AGb���̦�ȌE0,s�Z$���q�E�P�1C
O�.搛xu͙<�5����"�;���.�j�hT�sB�Q*X*0d4��Nu�a*�wo�l���yo���n%`���h2X��N��:*u��7����eb%�y�������Y5�!��z8�ň�]��T,ޓ���4y S�u�B /#�&�I����V%-G���.�4q�)�j�P�B����At�hբ���N��F��]�p���N>VS�Ǐ�j��2*�GX����{�7i�9��$7ϓ�0�`8�6�ӼW��.h��$�vO����p9�հ���s�m���X��B�x�dH���sv�b�1���Ϊ�n,�$?��'�N���iّ����:��3�S�&�e�w7���ݩК$�BWW"?e*�:��1��k*�|j*��)�$�^�N�x�G�6��Ѵg��Z��%-F�cHaV(iqDu5�G%�S�T=�J�T��k�0n,�ISS�_L^��o���gp�g�41u�Wf�_<�gj�q&���xV�@Ω@b�sϒ2)%x=���O�ܻ��.b�����f�Ѥ7���H�܀��6�~%��r�fD��#��l�9&Q6�9tϐ���Wr��N��A\k�q�<��/�57(�茣�lT]�)S{mBD�_�a���t)��@�,����
4��ҧ�"���a�
ț���v~]�AG�O3���=��M�����F�ƚ��ߨ�����Or�ȕ��V�y��e�
Py^���׮�ØA����r�GL�(@��	c!�!_�Z*ٵ)iY�	F�p����q�*�� �J�Q#dG����|�ˍ��i<��P6i�^Y�Л�ς��U� \�3 pe7)?�F����&aй��e�"e��!�ᓙ棆�PLI��u�j�z9��A����� $)�&���2Dh}�<ӈEέ���o�����[dKj���d)�
�a�j��y�.�ٗ��<&[�bUi4��7]��wc3����4���o0Α�^��D� <�M�t��Z����JY�ݼ�| Y>3�:]&��q�&r���y?�Q�F���D�TG�CNj����b�kM����.U@4�~4~W8�*����c�:EAOҺ`Z�Rʫ�9�KI
ǘT�ʉ�"�2��5U���v�ɚ����d�X�
f!�o�oĽ��f�c��<�ϝ�TV�1�yVH���8&�=bGR���ӂ�~����O�C�3��W�� �5KO��0Y%q�P�*j�N��_����=Gmt����Sn�c��@"F��:�X:�)��z��q����9��<��ZqE�׽�.BԔ
��?�����k78±j*���o��5�(�����x0�����E��Nv|ol��裺2j*4�h5O|�(�̤�̝;o��i�A�y��q F���5��e0�<D�2چ�]{���X�'�8K��:��ڽ*UZ� � ;d�����g�UԸ�T�l��Ɍ;nTT� 	��ޢ���Yt���Z>��~g��k"t�5F�#�6���P��\�B�VT���J�~W�|�G_�=����r������b�:�̐4�π}X�e��!	�����t���7p��sf��~w��S,�u�4��k�̿b���G�#R2B���3���JQ���:_����6猴A���/�xeE����n���5�^��Q�������|�i�A�(����d�>�il�����rq��� >f�8����0� ��ԩ��@�'(�����O��m{1��p4nP��"]�J�`��}GnK��޻��E4�ix��0�ވ�^�`��q��Y���F\:�Q�3��L�hu����S1y�7~����*�<��Asn��?�Av���{�;�J���r�+�.�C�N�z7�\��cQХ�a�"�����DZ:�4��Î����T�N��Ʌye�`�a)�\-{��@^��J(��ð���5��|�T,(�S�^��i���6�h*�4�����蟇2?*���GC�;����88pE���t<U Ը2�Բ���5�ZM��A�N;Q�˷	o�b)�O�0S�����ѯڷ4x!����������{���+`���-$]x�s0���7��F���6�Z��рȈ����q�o/o�Y�G�,i��M��>暦�u��?ۦI�,�=`��BE( ;*�(%��c}�ex�1��f&�5SR�K��P�jYꉃ��j��$V)aC�ү����!�����j�JZ�3�Pk9g�������u��s�>g���o�B�e�^���d�:�{�t^������� ԕ�%�'7��@O^�J��]2��#8��"�'à&NJ+�Gx	��������8����DӘ �Ġ��N2���%L��>ρ��GY�	��XB�B����o���S��@�V�kf��y�ggWJ~;�"�H���&0v����sk��$fsy������ S��J���z��u�譻;��GZ�3S�0Ϙޅ�e7��7ry��6�Y	@T����*��<?'��ju1��\�s?a�D* @��u�8V�0F�����$O�n4���� �p���9�x\s	�V�ݪ�|�֩A?��|��sܟ �AN�hG��f@:�P�U�����=��U� Ɲ|ݶ�PEd@m�
�K԰�o�������!��#��}��_�}�]�E��Q$��R��{�o��)xPZ䝫�y�ejcұU���v\T��8�3���"8"�!���w��FK��Ǣ���E���Ԕ�%iyX�&�sN7��4۩­=�@?�Ӆ�pT:�#<�ΝBŰ�i�1�c.�3P����N���F��W���ΰ�*1��_NJ���%S�p�(I�������Nvg���d5�\^�;�**b³L5rfȿ�KM�ޛ���xg�k�osKަ �w/�m�=����W�'�ږ"]�7����r��\���0@�<Q�gg���rF�Q�1��{z|$.D�1i�$q������Ϗ�p@��m�nw�)c��(���a8a(Hid�J8������g��D4f�l�;F�
���c�U|�I��ψE���~/Z�d����������:;����*#n�;q4C��g�T ��θl��"�o�gs��kZ��"��f�#��9��>���λ��}'M����'Jq \!DaB�R�"�"���D�}A�C��q�i4�Or�9��9Ɖ����@�bb�>�5�H�����z�8��Nw8ᴃAF���KJO�>/�Y�P����qh����NnAU$�s�u29n��pF�F�X63�y�t4X�m��_�
߯s6�d���"&�͇�C�U�.^*z)^���qU��/�K���Pt��ݣ��5�jե�֡��s��R���y�vEW����L9�+�����Rrcܩ~)ө�Q�A��f
�{�1�l��ռ1���&ZA��׀������dl���x�dM���';~�-�W�S>w�1��tΨ����[����&�rƘ��IgQ4H�nA�B��� ,�Y�D�L.��y�q���2���9�-੓�a�b��i?}
f_��Ff@I�{���7�6���}�v�X5[�6s@08���ͷo!��@�Q��@���_�_�P��(ªFg�
L�j�`\��K7�0�w
����fy����_R��ZJ��%O�� XI�_�=D���F2�튂���Q��E�0�����ۗ���qF2ͻ6���Z��8_�"\U�ɇ�G�޴���|ϻ��F��E�f\@$z�i��v�)b��<>�m�Gg/os��/�C���Wڙt�Ԧ�#($<��}���^�VAy�6j)#�(�1l}�Z�f/|Ǝ!睁��-:��&[W�*YDH���^�q�ݵU�@�'10�HD�����<f�`��.ț_����A���ެ4�"uH y��s���hxVFv{�H� ��X{��"�py�Թ�������B���$��6��مyx�{]�H��p{���9{W)ED߈��vo�~��k�(ctԸ3�N�n��G��#���9pBRe���J<F�v����mR<�2�K6�&
��R�4	������a����K� ��n0 ��캏�6�F���@C��s%�\��z+f�#]$�8�Y*f�X�ďps��k��%���"'�3�j�^�>��w���s
-�UPz��\�������8�ދ)5n Q��Z����ؼC�v�,Ǯ��s>�j�WmJ�p��:�}�{���ߩhbS���bYj4��'�	���Ѫ┪��!����ZN�����7��r[W�Z<����2����+QE���h��U�d��7�j� +@7 |���V�~�J��xp���#�=]|���:*����-#W1��h�5��#�����O1���*���3X4!�N"�D���Z#�:-6�T&�0Y�Bd�;Y+������'��0^VTedˎ'' FC ��;�
jL�z=��~�6�~�h��{y~y`E�g+o����c�u�9��d,�j������0����� �v�>��hC��Yn_mհc�`+�}�����eM�~����V�x*�&9�q��Gr���<�Ȇ���<��Kbxa<�"�OS��%yV.Ԁ����T�wp���8(Z�!
^d�d��"�qÚ�A�3CHOC�������K��T��*��M�ڂKu�:������0�Ή��X����_�=�^Κ��~���|��O|��Q�(���]T3�A$E�����k�LǖJ��r��^m��%����&i;��5��Le�a�Z��T�%z���8bC���|�]��0��O�1a8�g2�a&-=���s����T�yr~���*D����G�ܬ��YX�]]���]E�0�����3���f]�J��;���������T~��V��\��BN1��o��в�,R���CgA�YK���Y*d�N��Gc�יn��[�]{0�}����?��3����������΁�L��J�3��@}2�R�9��=UJ��w:wPp3���XR�6��ɪ�.#{���f��}<�&A`)��>�S�_gM�,Mfk��u�q��c���B%��68����C3�UO�^�K� /����C^��c@�L$���T;�͌
-��z�v����~��混w��8|��&I-ʱC(��Vì��V=u���޻��z�ӼV�ga3~��7��-XTT�S����go$�CU���
<9�񍠲7~ %kv�^��^�����*��O4 reP6�=����!�����.��WCN�K��3K������_g ��������� �^�sb�u%�T�M��g���y�_^ �7�)I����@f�הo���FW�0��/,�	����3	��o�h�!�@&H ���]MCC���X?$D�)O����qn�#ˀ�y�Q��$I� �:4����QֵW�T��5J>t�:��x4� V<���ջ�1�^o�n�����EV�����\��$�E��a��C�s��xnx�0gp�q���f�� ���a9v��s_r�?���6�V� _�3���Y���\\ѳ�)�'��X�����>���=�Qf\W9P�C�^�)����?��ވPqh���F�>���^��<��n�
xI�,�/l{��2���X�i�ZԽ\^�JFAfZ��ِ]6�]���Q���T��_��ISA'����&�����{��Q`���:�Ij��OoC�%��i�rC)��caR�+�K���,�=u&��!��H�1p�,Z�ci���d�_�ዮ�T�cS`�p�:U�M)E�4�8�p��3�l����ؑ��i*F}��dǎ�{���zN}ӝ��w�~7�9���J����Z�ASfld�jv��9�"�����hkMq�t&N���j�H��J�r^�j����%#�^��"Y��p{ʌ7��vP�~v���8�U�E�v�&Ajzz��c���P=�4�T7���X1,���"��9q8��4�����~���&Cװ�ҙ*�4�_�~;7v�al��p�J�@'L���*`><�0e{%�a��׿��i� �}p��1���0[\c#�3@dЋ����J8-����"L-uG��v{���~�9��yo����'Sfs�PґWp��|�~��`�Ǽpg
�M'qG7��:G'yی�&��	x9���7����alѹ��:�Z4����
�h3=�wT��KvG��b/^:>���*����BoL3�\G�`6��e��
3 %Y`.�vZx�5������hz��X&V��s���;+MD�MT=CuOrm��n���Q��:I�F|�Vl�/�˱[�TJu^~�ۜ�"
cF��5n+߿��Ji��+��
�t�����6�����M�g���4���H����r���y?eq�������{���탴�=��3|8����2Ɂ�m���~Q�&� <�Yٰy~��mV`��`7�o�?h�6#>��S���V8���B�K/��yOH�\趃�]Ŧ�Vy�/b�`Z­ܱYhTqB�|or0ڇ0���蹻bއ�v��i�@_�ә��q%a��C�������CO����Q���Ш4E��=S��Ke�(H�E
UZ~���d��L�D�x~*=�n+�?�=��J�#�������de�18�1o���T�G9y*���7C��iO >�+�2ҵW��~~���IyFz�!�y������tS�V5D�h�kF���Z���OD��i���a�����QgV��9������s�z�(R��+zcג��>�-�z4�Ĉ���r�swfQ���&���^rD��s�B`b9pEH��*��{��쪌�Ya���}��
A��j�_�^$"��S��h��FD+�qsX�
<������� ε��6�Mޕ���a��)YR|rtoo,��~F4�F�h�
�
zN7Q�����gp���F9����Hۯ��#U#�|�|�=��y�4��	l����FǍ�v���<D0x�ގ<���H���mve��{������Vޚꥡ�jI4�pH�\�H�R��l^�\�Ӄ}���O��!iry��#T���ɾW7�v�؅K3C����JE^(œ�a�:׫S�#�>����T$N��tS�[87�4Y�W�x#<ֺ��l 6���'K!���d�2��E݌�u�nd}e�����N��I��;�ni�%
gN���Ï���"ee4�Ȣs�o��Y��ˡ����؞1���7��<s��
XF�e�ؙ_W�XHEX��\[H���ї�88�s	F�it>����v)R��m�E\t';J	��a�������	l1V��W��4���|:q��,V�Y_㩼N�c�}����Ʊ(6%?ǾHǢU s|½x�4�4�!5���b���꒒e�OV6���L1�Ϙ򂱿D���%��A8����n��VS��������ij0�\^\�s�F���*�#1#��bB�_ʓ�}1��l��?����XU�h�9#�S)Ɛ�ث4b�S�ə�������J�+���2���&[�0��e���!p�|��SD��� ��ڠx��fDپ(�����������F��5���YQ��xÿa[��|����9ez��au:5i3��v��fV�Vwu��ѹ��}���ŷ8�6�w֌�;?h�A;�;u8���id��X�Q_0tX�Mg�C��w���-FS+-Z���^��u�Ȥ}T�������q�
�Jp"�@���ՠN>��Q��q�t��+��|(�0,Ŏg��Y�Q��6j8�g݊�\�U�S�r���بz�GG>���BR|�BEr��N�l��8��������F3���6����)��P S�O�AXgMq�ҰV��JɃ�0���O׷=>�&s<���^8"%9����׸V8�7����$s�q�#��$_��� G�{%�2sI�(/�7ʼ�+���b�Xr$٬�7�~#O�e~��Ӭ��7\�R�~����Ln{Z�� *ŌUρ'w��uꍿ�8����r�E�n��w}�2��[�W�e
�〦��l�)U#�I|��h,�⨽<Hbj��?\�/V)�]Ӽo�R���=��+�pLEiRi����L�P�="Qv�<��4-^�ʗ�V��!�I�0{{R�>��|���
2�PwV]�d�*\�2 �fB�b�p`>�r�3S���u~6�s���憞��0�b)�NۥR��� �������/����?���;�����ә��׿|���/�����<q{*�P���;���dY]	�w�F�l"��=��}l��^S��]G;�SiԒ95tzm��Jj���k�7�U$�W��9�i�,ق��_�j�*�����v� �c��^��;�\+XB"A��-�>[��I
�F�(�⟍�,dHDSh�L�+�9���	��V��\�oh6R'nv���~�A���0H>Xj?��0E��Eן�A*�"��<�[�6^%�����W,v]QHJzE��z�ў��Z�u0eb�3�?�g+?����V�3��Z��H���v����b��QE�!�����)k35�@��m����� ,%�.�����fu��(�
1|q�|h(�x�D��4ܟ�����f��`��w����v:L�yj�+��q���S �����z���YT��ǔ�
Շ�wn��fܰ�U�7�T ߉+�N��=�2�f^�����+h6��������j<l�d�_F���o�7P�*�Z�x;t�C�=9�1�Ɠ�1�r�yl�d�l��F:�^}]p��qm�n̷������ظ8ζH$�a�[��"�$�L���Em�R�ʳ�QX�sq�G��������4U�Xz�������"/��tz�b���F���[�)�CP��LKz�R��'���΃}�qژ#j����8uƩs/x���P<������(� ���ω�Q�8g޴*�r��y1��?�J�2����y~�"+�����Q#�;�E�-�N��_A��q���հ$iT��Z���f�E8��?���0��!
J��yTqB�^�2�웽E��	�T�*�؏ܮ�����;+5m��ӓt�Z�|�H֍����{�>�S����ʟ��QbTh�Qek8)7Jb;��9Z�6:�x�˫Kb`�4M�Fڳ���'��a�Ua�Č����~x�=�9����<�5zz��� 93Ҵ�Ϲ/!b�|�Y����J�}�$�����w����iz��}�FJՐ����(�sЮo��x��ww�h;��bD_��5����^l3�s2'q��Y~��<�3��p�}�c��|P���[#5�9<"RJ�f*�N�r��]e����{��TE.�wxլձJ&E2n�brNW��G�WHA���Ce��R���0W��ph�*v��s8&4y��¼ov~R{�q}`�Y�j��5��P��G,�����}��ʫ/ru~3��M	NG����_�8���g�ϊ�У���:y*B�1p��#8������&ħ��lBI��6�� J_� 4����T)8'#76�E�Q�D�6�uc*�N���~�����y�}F.�-j��񓃕�.��<�n�����5�7��̂ܳk��@Ӭ�T���z��CX;7^��LFf�Q�&,'�B ��o߿��dyF��<'tb- گ�< Gyڌf�R���۸�vV|AE	��-/�y�
�� �؞�	�\���w����X�Rˑ�����6���+a�Í��Ͽ�ݝ���4��o?���ͻ���wǀm',�gu2��(X�''��5Y���OgJ8s�A����������5F�#X�7����Z�� �K���x7JHQ��c��βg�/������K(�Ϟ(�͙#����mT��
wb�x2cS3�sQH�j7�	��0V���pB��������յ(%��H�P� cxv��b�Ju��qߪfW����2K�o��\��0ؓ�  Blc�a�Eu��e{�GH�V}ɻ�^��>����z������p ݤ';�@�J�%�N��O9b\S��Cq� l`��5u��iC�׆�bd��H
ft�H�S&0Ѳ�%��g7N�o}���5_����o8z#��biJ��y�����h���ZX����ɜ�a�GjD�p�5^mU���b�I'"v��Y��~-뷪�j���K�S�� �'�l�_�A(nĲO�o��mS=�G[�l]nT@̠{9�3ܰ�D�ì8uf���V|�Rɀ#�Hc�ъ4��'"�>�>Z�����"��c���?����Ӫ"�.���s�]��g��<�>�te�m�dYkF�m�<���]��34*���!Հ���'Kg͌��鐂����C�Wa�ߛs��D�������G��P�I�>ӝU_�QY�%�,�4����q��[�!ve�љA���Γ��+��h���,4r#�+��]j��5�X�iu�ior�}b܊΁Y;f,�AS�ðD<5�����j�3�gr��}��8�ި�y��P��n}oѲ�p��,�����/wv���c�Tx\���ƃ�"Hr88����'����2�S,#d-���ʲo�,�8Z修��%��~�򂔴��F��H���2��6�2�>�O3>}�|y��'�_P�ݢ�`�A
8l�A����ΩL�'J4�<=����Tt�z�SF���9	����L�b3/��t�x*�D�L�g�֑�:���=��}��[���_a��#��P�܀İF1@��U�}��Q�,li,���_�i�D�}�2j��Gh�?�:ՑL�)�&�,%�э7�W*㶧��\Hnܱ�ڳR���u�9���2z��%`B�	��1�Kj�A���;%wa Ytc��.nU��&�u���/�J3��F���~r��=���ޢCFnn
��hMlx�h�dü�\ 4�?�[D�8i)��lz���dy�vޤ��ay�4�b�>�1�I0坕O�Ҝ�fٍFh�
�\��J�2�aʺ���7n�4K����`�^�0�ƨb �"�r3��:EI��
�^Y�$A��%6vx,�yq�T}��]�,O�ƓG�������^���ٗ]n]�keG��C��2-��	���(�_�����8چ��S�4t�(��У�����o�Y�U{P*tZ�.��� �%O���]�򒮔G(�,�4��� �4������,����!�y�����O���ZJV�zá85ۅ،�(rc�hB�7>���<�C��PBKH<^C��J*�ޓ}=� ��bE-�S��(����8y��S�?e?�<�hE_��i�珢l�iZ�>����5�[�|LCB��,�n�BI)᪀�%!���S� �������&BO��li��Ԡ��u&'W��DNo?�!�H�Y+Gװ������12uAd������sD�iǰ���"v2���E�鳨�����7�l$��G���S$�?��E��#�q��<h���ΣQu܈ag����Is��^����{~}��x�L�S��^Ƙk]�Tv����#��XWU��d�)�4��{��rkl0�{i��7����l2w��V�-X(��d�><)ѥ�x{�%����(w!e�<2�'���� �v:@sÌ�g�|���~���8n���yݪ��]��t?� ^�5�v@|��z����0 �O�˾P����`�T�8�">��ܛ��1���:2�3�w)��+ <R`���^|�@�MZ,�+�d���{��iS��cv�j�R5�@'JV�Fy�D���.��*�e9;��2���J��T1���iJR'WW�YQ=�ח�y�~1~��Zg�g���x������{�Tq^1UQ(h���<>�6�_�]�t	�~��F%ղ��|���st�"��Ҏ�4�<�/�Q�)+��@����f�W����0u���~e*��C����Aj��i�'�4;9N��߫���N�OLۯ����ᠯ�(���݌c����ӂ%"�1+�yor����8���N M����,��0n�f���8j�}����!(����
�-T��s��D��C��;�ؑ8 ��E���F�{�s�h�1k��
���`�%����3�D<>hd��Ŋ�UM���J�ڞ����QfX���������DZ�?���<<<��	���� F���S��)R�� ��vV,D��7fD�5�ơ:Z�`����q#�:b�u��Xu��$�.�b��؊ը.�M���/����E�J�|����ůT_��k\�O��u���뮋gv�뺉�?)�Z�]�u�7�ߩnJy%��D��g��Iիzj����4��y�aGK�ж��3�m��=�����7/���y��ơ�,Lw���&�N�x����6��)©���]����.c���I�R�;��!�KVq ;wPQ�}4��'eFI9,���S~��4!�K?ׁ�jq�R6����ڴ�&W�<İ�Oa��=[H��|�b�*)%lN�8�������Dԣ	C�|���
�^n74����D�H6���D�ı�Zϭ>������8��`Z�\����w�*������y���yAh0����r7�(Vu굼9��R�j����o%�|^�_��1
�{�T�p3J]�[�¯ ��â�P�;q0����g:+�-�h��(Hm�(���Oeg���W)�SR�_�5/�C�Cg�������`c;:ߐE����AmW2�V+)���/'&~$�d�Sj��}�Qw������F��U�y�F�KT�W�P��B����� p�L���0x���o�6�	][ʛF4���q�V��S$��6�aC]�=ˊ� cê�6)L���Ǧ�aTM��e^�H?ZT� H:y�c����Q�|q^h=�D0��3�
OV��r��zf�x^����J��]�S1�`���D&R�QQ|I��ҵZv��sI���:·��`h�.����0ZN�pxdQI�-a�*�_(#Ič��G��q9%�}�"�ݠ�{�9sZ~;W?NE�uU ��D�����Bj�R���r�zB�%��y+�Svý?���O���8g�,9�Q%��O|�Ͷ�G�c���ag����z�ɉ{ò����xxω�r���h����َH��-[���Gu�x��Gh��X�<5���'Sd�E�F�]qH���E ,�z�u���i: �V�AVCVrL�Q�JX,4�랼�t,5u����Cc����-���C�Q�g�4>��=_(a�
B(�����U.�o�{���w�"�UaB�
d�[���<c�Q��<����=��a�ĳ�������*��\71PJn�1La U�=I�
u�uGa��׹P��T��=(�fe��.�>�|�(�މ��vZT�u�h^�?�z�^�ۣ�G���W�Γ��}ì{r���I�/jt�Z�g�^
ͅ��X�J��������[�	��Q"z�g�AfGc���R�;����i�^8��V#�7cY��-B�FǞs5��.����)ˏ�<ˢ����/�Ӕ- �Z�c}�*���3���k���G��,�\����F#���h9�W%s\H���{�)��8��@ ����Sz/gL�m���
�2D�'���{���v�c�o2jo��?����hO�����b��S�:��ɦͶ�'�$pC��Ӯ���A���8:Mʳ�r��j[p�Pr�^Y��{i�~��g(=��Al�L�@����/��ٞ�N����t�C	;hB���T��?
���ڐ,��8�5$�z�ښ9�W��JK`�U#�<ʣ�xz%���7]L(��<�TJ�7�~OU/���{��� �� )f4�0�_�y>w�银S���s���)�r�Jmmj�a��)�px���p,&U�Gǡ2�.�Y5�� wW�HFا��~���>LN5�m�����' Ro%���<�9O���Yd�p]�@`t��+_�/fp}n��,Y��k��(��`�"��bM�P�Ĕ�cd���H0]����@%R���aeHk��ڪ^,�*�E�7tm���W�����֎L�VQ�Șr��6#���c�0-~�K>;�����4��<|�)�H�@�?A�[L���#�X<�zt%m�B�ce� ���ɥP�
�g󶈍�EW��O���C&�O�B��nT�v�	�)��F�Ɂ�d Ɔ�7"�����=g���L����"L����$�b.��:�y��� W��%Gn���i] ���F-WRJc�i�t���+%���q��d?�bp]Q��r�v!����>8���[��Q���e�h]u��;5�N$�ރ|u�S���D.�b�z_��e�@��C ���v�[lM��M�%h$������������p�������\.�z��]��-��/ /��c
0���o�����>D2nlC֍9��\��Ơ�{���ār�?s�=��G�q�y^")[�;{r���q��f0Z�h��>���^�/�T��<<��l�jD��XcVC�Ϩ�zt�����aoM�a.�S<�j����Ͽ�J�8�����S�*�)�,�	����R�۷o��A�1��$y��Cu+Dk��+F��6�f��H�ʀ+�� r!�|�����"����~����o�W'����20ʡ&cV�X
��)��x`�n�Y��?go馱��f��bUu\#9E����0Z��js$*�%5r���b@���U��׬��6�%�>��r��l� �AC瞯�TR���s#�5ҷ,u5.���#�tv��z�]u���}�ĉ�Bo[�u�34�Z�-���s�0��>���³�R"������u�pb.Đ�n�Q�촟����*��u"y��i���eU�Ԉ�������o$��8)����:�a��1%.�/<��(���)��OM�j�F̣��"^D���4�1��d�N��,K�"��s��L������.�C���>��~���6�z�äd�a 2�j��1b���1\�B��cg9�ͅp�F0�����|�����?��e���Y���-��Ӟ��v1�����|_����A>�\~�+kަ�^�2e��
=VH��=r�//���z��{b^����I��<��P�V+����G����Ebg�p�\v;M �妒�r�VY|hU	#n[Y��G�Vp$٦P���#-ZS�ݤ^X��S�Cv�f���׭<� }�^!�y�k�E*�l� �r�$�8�&�e"w��H�B(3���()��s=h%�}�C�˰
ef����)Ujh�Z���@8x�ʼ���Y��$%9ud�|X5�����R�Wv�S�1����,���p�Z���vR���l$��UzB���Q[�����h,k``\L����cS ��9�����6�L�)).)�Lb9����1n}m{TvE�(�LRR>mE��(ZK핈����Ƃ>����3ʫ�K]�"�F���f��p����}Cp��Ͻq4�u��#��Xw�f�k!Qm�p�r�?���<r������K�6����Ke����=���L$��m�zͤj�6y���=����#���%�B�y.�n�=k5F"a�Փ˙�[Z�ʄ��������iZ��c��+�ݪ�)d�+-�V��V�M{GK;���zև+6�� #b6Ugz�֩X�h,�cC����K7Ts�N�f������Z�o�dm��7"+K��=��P����RMH��>��-��D�\}���?K������7J��E�0i�Gbs�ӈ�����*��Qq�QS�8���9ϕr[)�/J+k@J�hk�LɆ�F�QSV�^:dL6���h���wr���aewf)<j��10	�v���0��3�E����y}Qn���28�`�a�,9%G�7�4ZMY9��F�a����#����K#������ʐ��K0V��9Ȉ���-U�&["�"$<��ڋ|R�ܤ���9��[�5�a�m��e�r�b��iLڤ�q�8g�o��b�jա<���0��5�����ULAtN9C��B����_��].kR�)�I9E���fK6�Ξz
۷���$窒[�� �Lqcs�+UF[?g�%د�������b������tS���,��s���;_˖��W�n�`A��S��>��AJ1��LX�
��x��j��i�Q�SG�#~ڼ�y�-����g� ��I�a�o7sÿfj!�SY[�r%��W$~ƅ�h>�K��^�E�6{B��&Q+(*�q��r���X5�:Ǥ�s|o��9�X�I*���������T��/�U.� �"��削���w����n�+T�������v��9�7�A����6�aY̓�Ht��Vm1˭�}L�9� �}�X���!���K Lȁ���ꂹ�^M`l(�>1	�<�=�~y�t剋�C�?���*W���:�9���7]�A*��o�Ħ]:C�hs櫈��-���^F�$�n�{j�.B⣂��ਕ��A�J��@�3<_%,g����2�o�Z�y���1>�еl��n%i�� θeL�F�Rי�Ž�\nϛ���[i��U	��N�,x~0P�Lq}}+_��[s�!89��c���V�=*��}H7Pq�x�WS�G�`N����@���-��m�`:�r��I}�&qN���e�$��~�}\����4�o���r��g�a�T�Z�eW���D�Y}dE��f�48M�<�Nc�豩�"[�ڄzDBV��Y~�ITS�Q 1e"T���Y���Y�Y!�M�\���~�4�ؾ܃�{
����~r�|d�,���_j!�B�c�$�0tS�����Ƭ��y7�����9�N�|��r����L:|�.Gת��V�[mt:���rɩ��TKuI��X���:U$��q'�k p�a^>xI�.m��+���#"Nl�jl}D����޿R*��u|/���e�*��f�r��~�{�2�I|O�Ƃ@:��7�zrţ��92�F��y����Wg�3㛋Y�v����6�c8kkH��$�Q"��ʘC,���<ɉ�����P���Lke�}V����;��Z�չ�<*9��6��G_l>�y]�ܧ����3�J;�2E۝x5&1c8p�/�փ>����Wr���kG�ߩ��X��Dw�f�'K���(�JTp>i	ꭑ6���T405��x�/o����qlʈTЈODݜ�����EN��!���9�JT3�AYt�8����kf�lF�,����X�Ю��[s}��k�o��x�G���s�{uB('����ڋ++���UZ��h�������T��� .�[w��ma�a�TR�l��\'&u��]���e7��H�ܮͥ��Ǯ/��\Q��9���$�F�Tw��ʁ���>�uY���g�<���F��&��iU4t���[�Wx����	F�m�B���M�G��Nr���p���E�`�ʪmz��?ފ�O�O݁�
mN�q˓�әl��x�����T��{�����y;ϧQ�u�q��Jٸ�:f�a�3cf�Ģ�l���K�?��hB��kQ�JUc��a��%����i���kW�3�tS�-)���c�����sg���������o����4��)�yBi��CnͰ#����v�H��-��5sݨ�'f,�c���1�^�dv1�t����-%�q� Zg�m��B���}"[L5�K�����c�$�e�=����|Q�f�@����s�\&r�M�.�X��!�A����sO�d�eVU��M��jY���.3�+L�k����I�Qj�	U��ţ�I�$f4���6�5x���D3����ҋ��ɢy��5"@����)?Hs������\t;i 97����{?�d��2��s���ÎWuRϠ��to�J�Y"XRsR=�E`%��hp�>�#�\%�l#/2��Q��!��}����׋�)6XU�*a%qR�_{�µUP��)F��/K�j1x��!c������R���EC�;�'��Z����n�>�%�dUHv ܶ["�~������ 4�1FM�k�V=w^|���t�?�z����|Ľ�}F�s����� ������m#���$�˲c���g��('���l3N��8sm̥mRd�C� �����}�ٌ���Ik'�����R�b�}�4__�뺷"�#���^���!����$k;S X�dEE�o�+}ȟ��9��'T�q����9 ��)��D˝�p�i���0�\����n�ٺ"�s�������1+�s�̯Xr�8��?k�M����U;?����}u`������:!� �d����Ր�*(׬Ι+����ށ�$����3Fͼ�*_���F^^7���<ゝ>p}M����잎�}�a�0��^̰�XO��,˲��Y���(�̪�ooL���*E}����Մ��5�8J���h5��͆MҢZB�F��>�k�B.�ʸ��1>�w�,PCk����=��!Z�\�b������T�NӨ���g�¬b�b͟^!�|�b'�i����[�Э��&�������,r8��{�=x����Z�뇚������%����H��0^�����KY̐�OO��wp�_Y��-���9�@��62,�i�|�RUˌ��R��?uD�]{�Kb��jT�1�.X��斋ϫc�>x���9���G�V�f�:���kt|6^��D�uC�)�q���\S��f�cD��I����\��XV6R�e��X6����D����j�Uu�	�ߎ]�Xp�Q����ϳ�H r���$�.1J,���0��@Hu�Z��[Y��?�#�F��J���At�JE�ߚ�)����z���`�ַ4�V�Õ�K���	1M'Ķ��dٌ1�O
�����5
��S�	��I�4��O�g5x}hTs�#��R�5.;Ng�����hNz�1� �#��i�?my ���j�:�3�yy~en�މ�A(X)�13B(�����KL3��,饚,����Tq����>$��}��+�pPn %����мћ0��@3PIb�{�B�%�!K� �TX�R�"l4)in��դ:����*-�#��F�_:���.B6ׁ(?y#�Gw9�@j �L�j��{���[���^������F�.�=#���}�%�Ĭ{���X_����=�HCһo��#}�u!��b+�俇lqϳ�6ʣmO�7�l����Gh�C�ww��0���� �Q�U;c�4�C�=�zX��+SG�e��blke<�şOￏpџ<B��:�Ƕ9Ӱ�g����( �$6��^hF�]�̚hԡ~��/77ryy��+�3RZO	v�\�~�������S�0:�������U7���oεg�R"mӮ��wC�rL�͙mչ�K1��VJ�����f��x�հCKֳ�yft�9�/�6����x:�ް�Wm/U�1ä��N����Q�` �'�?S,1ɐ7[s`�A5!�漽��4����2\^\�xsMʋ�5ܬ/d���f��Q<Ҁ�#����蝁��J���8��sz$�p��s'� :̹������{������<��.���^"��-�鴰����ˆ:���'�"�|��j:��N��j����g��ͳ�x�,8>?��s�Ʀ^!8���P���пc�rZ^~�,�̌�%��Qqw�0�?���h�u��|y��5����|r�~p�ζ\��ؙ��ՁI�z��J�=.M۰����EJp)e�[���V[��y��x#�0�b��5����Xq�OFo0iIv�*>�1���#
�H�B(˯���Dh"q0��
0�kz��uX�/���7��LӰ�S.J��G�񲅗ɬ&�$������Wx���= Q�DAѱ����m��$@�g���dYt��]��k�s�gr�{m�9pNS�(�#~�&��O��4`n�K���{�V\���4�@��+a81��cA>f�w�R�]���<My�$ɛ�������3˙?� ��mO�i2�|���})�6�&�����T�VpӤ�Թ�,��Y�/>�`���ZA�54��P� ��}�5���C�qO�G_Ofh�"��(Z� ��w��cq�'�����,`���}��R������b��ֱ�Y��@���k����*�gy{���RǎH;���j�����p����C����/�IN�jN�r���������N��/�bI1t99�>�hWx(�~���F��j��iyC��Ԕ��!���M�M�ԯd�Cg�"w����J���\{�k.��������ovߔ�z,���O��4!u�{����nxc��i_<�H�}�Æ����(�\%�8?���+r���*Ѱ#e\k�{NL����'7;�w����R*���>7|��0�2�z�{���I
fj�ܛ�:��jp�6���q.�w'yZ�Q�NP�Q<��c�g��������'y�ft2�iXJyT_�칌𔮪r���7���w$o�~�ղ�MD�6�e��2��6t<��^J1x�p}'|�wQ=�Y:�p����v�a�V�Z}F,r(N��_IG��#����c�Sl�Ǥv����߱�TM=���}W[V������X�Su�#�0�����G�U�]b�ö�����[�����k�b)�RUY-OS���Π?��w$�4nW��S5�m;
z���Ϡ�?z�k�����C����n���Űl�����ⲕ.��R�!Oa3R�����n�,x�hAT��6��U[-R+��M�a����N�6#�Z�*b13E�;���������|�dV�Ί���>+[��?���͙1g#K&*��z,w\m�l����ҋ��Jg��Dh��.�ռX
�7��{dPa����2'U�{�	�@���K���T�dH�(�Z�~�����1�M:*
��j뫳��/iRW��hI�6b�A����@`���>/ �
��v]�X�DҪ�����F��7-+/�Y����¼F4�9H�z�A���Yڢ�Ԙ�'�%,{.x6���l?=.�WE�ȍ�Tk,;}T�R?{�ȻÍdP�l" Nx�#��6+��<��t�oem��+gz��[e�DjC��n���Z+!�iY��WXD߹�RD���<Y���,��K��x���̣Z!8����1Iչ���1�T���UuC]�8\,����C�,��4�.:�@��vy�O�G���U��g���ǧ��X�o�>��z~H<zD������)�a:��wd����s-�>cƠ����yfr��Yb��m2V��T�a�Ndh׭�t̷���|o�b��|l��&v��ql�iN}�:=Y�g��r�J��ո�yok�/�� ��P�>�� y�g�s�R^��s��� �✣���ٲ�)�iU���vT�i�%7}p����3�L�mu����a�[=ܽ�(fr��;�kk�>�hR\���cmi��t�GV��t�]�9�Eg��_� ��_����8�^�lr^u�uVԃ��:�����^+q*��~�(d8lQys���U߳fd�1D�HZ�+h�����Ņ��Zb]��G��V>�Cn7��gk)���F�m�ǝW�-ڬ���8_��6\|�c�,Ω�Zz�sỶj�?�c��hn���
O��8��v�����Z�t�T���C�\���ZO��ո0y��vX�z�y�ɫ�f����Zq�0u��n�����c�x=r�,�|�s�����]\���T���g�{�X���ƿ�k>����n�R�ޅ8'ے[�ѣ��ˋ��xւ�ZO3Y�b�+�e/>"Z�u�:��Y��^:����3���YgT�O=}�V�����A�!��Gr�w�-�Q��{��
{$�Rf��c�TM��~ῧ�yi@�^Q���(jy"�;�f��_\�%�zZG�Q}��A�dI|n�ݚ�SmdX렦ṕ�G���Xyʰ5'o�Y�l5��v��{.�f�A8)R��>1��"�1��?��>��\���E�n�f��w�P�0�h�}�+�`M�f+y�X��+��/�ˍ��Ro|�L2�ΡRq����:a3�,�����W��IɃ\s�]=>=���3!޲�Uf��?S�U7p���^�:��M:T2�}�py꼙,_�ɗ���s6h����>(I
�*x��_���0>�U�!�;Q��t��'I�-©o�#I�YϱZN/��)Շ;u|��9��A\y���X��~Z����&�����������+gyǸ�W��J)Ic�h�d�GV��=rW>Ҳm�;��ko��L�r������9WݤƯ�k�b�^D��w�K�$�;��??��q
��nk+�
Y���a��g��kB|c�v~=_�I��#~���9��[<Wmt�+�d�J� )[�ZO�H�]��w����`T�yL�����?�3�������r�f�^�?�d���������W��cFFe��Ռo�/���U>/Hv۱R�^����>�l��˭��˽8 A�h6v�'�܌��Oown_6��ɕ��Z�|��J~S���`�Y�t�ǶN,eNGF�"R�NV�v�5��Έ�}�l���/������V�8b��xU7�V�K�IX��*m�#��nk;��Og�F ��5�v�� #Jq�p�3S�&���"����U�C�#SS�b�S���D$�j�op��vޜ�W��흏dF%�br����s�#�����͕�R�v쨯��j�G�~�S?�'R����]Fq�����M���m��k�Qև	?��*j�'U/��c�t���K�ŉ���?q,���Q�E���޺l�bi䓿��h� j�S�cۧ^�7�ʢ���,��o��<�=)V@�s~~)��w��� �)�hRg<��=h)�{2;Ì�l	�xqy%��7�5����u��ӫ��g�ؠϥ���R����XCi��a@@It��)k l�0p|��X��l.x�Q���E�=�MX�h_)�E`~�e�F�\��rE-�����j��<����k�ʭ�6>X�P
Fie���kUK�W�:�!�u�Fև1�S�ȍ�wH�B͍�g�#�Ql��'$�©�~� �s�\�\8��/�[eq��%�AEg��
".$,:�OZ}m���-+*|��.����o�����h��}�h��V��Wl'B�Y�l����-�dy޹m�j���R�&�1jo�E�s����'(�{��;���r��,�Pzss��6�xؕM��}��s�$`��ty}Fk��'Gb�3�	1��qv�żD2�a�s!}���mޟk��?����L���≿%,�C ��_��z����Õ���\�Y��(���z�fM�ܠ��x7��?�����I��G�Qlg����Ds�!�w/�J���"1.a�M��
�~�XԚ���y���e0h�y��.��+�9���ǲ	�K���w����x?;-�Bs�c ��;Nҫ5zKw/�H�$��w�3c����ۜ�s�D�e^E��h�c݇��!Ǉ�@Z�p�5��Z�o�m)�%Ur�VMj��O�7>$�/XS�m-����wV�G�^�2"�#Q1A�$W �{>>�T��0Y+GS�lID�:��χ�x������3��۫���o/�s,f>����̈��xj�Q�)�8i%�՚
���ϊ�A=�^]��M'�����-���J��"u��r��G4ߣG~��t��#rY�čB�6N����'�����w�������3�X�IG?i�+G-O��?�u��͑��O��.��(F�����m���!�}���G������p`��߈�ڰ#t�[@�~�},��c���x�����N���-�O�^���/�_�/��*="�}m���Q69��aF�s��lһ����syq-߾�$?��Y�+yy|���A�v�����J�3��Ӝ.�&��=w �n�P�|���Q��$��W7s���4v�����=+�����Y��h!mJP%�?�M�Հ)Y��ƽ�mt� ��D�+V��畗m^���QQ>�@��z�0�z�!��'G��!)��t<x?:�h��hKaQښJ��=zRP���mq�y�7��*�X�'W�� ���s�����dF������P�r�)Ujث��ڍ#�1 {9e�N�����v�lvJ�C��?��������8��bQ:�|�NV�������H$OS(��=�h3��ZΣV$a�=7`Zd�3�ϗB�د��J�*D��sT�@�5*`�{zqy6Ͽ3�!�iּN�\,� Y4�X$����:���)m��s����]-B-{������O���u|�{��~nJF9?��+�J��ݓ�7{�(9�����Ǖ��ޝ}���~����=��MKB@��yLU�hѝu2i@&�@�-S\�YbXBi��/��5�^PAR�~T�h�`q�ڷ�4�&�3��j_b����:l���#O��_:�4~�[M�[�"�������2��w�b�f]ZF�*��^�=@����E��$:'�c+��<_�l1��m_�38�]���f3�Un���ib�$���<�����|_x_���܉j���g��%�9!�����E)'J//|����W�Rg�Z�F�e���7Y�U�=g�B�b��2`��,���T���AC��̫��:�Ӌ�qFdaΛ���t"Bxb��6�f*0jc�𛬑�	�e<Y������Z:��􈛨1P2Y� �}��٩5:��b�׋�+�g#.�j9�j�AͨƝ�JAT�r�B�+X���88�*��f��	�4�{�n�rg�NbZ4�����[�5:�voy.$��ZWD���8�q,�2�����f��ʗ��s��yXi��G��|��������h���yt5f�S��`�bl&�-^Ul8�ׯ�*J�����F��q9u����"r�zӷ.,i���2�<��B�a��L���bt��=f�>P
IR��V7�RP�p�z����Ō�v���O�ܲB�"��VܹX�QY��4� �`�2�gp1_���
"��,�:8�=l(Al���KB��QV,�4�t��i�h�)a���g-��t�T���������Ԯ#�~�����0�Nղb�ݯ�03���\�
��5��UB8�02��Ov��.������1!�]`М~� P�Y��G��L��#����8pwÔ�m����y�,`v5}|��#��Ru�/ʑ����(8jn�}Kfb����`x�=:]'$�} #�	o��Щ�P�R� ���;�y�sl����A��7s�;�lQ����fG)21Kff�����A�~�f���v�ZVz��\#��rJ��Mk�]�(U!��ӏc��t�],
�E@�������
;^d.�j
t�YoI��Ysjs��jyW+������;���-���/l�v��l� $�e�Ĵ�@��K�Д�$�#�vw�9�fҊ㕎q�wig�h�!���Ob,炝�X_	.���}VAt^���V�r�,󳵸p�}.W�#3���0:��I%(�!����H�Ä�ܬ�sa"����^.��tL�D�Ϗg(z���d�*C��4�)Ԋ�?����DN��.�A�����sʻ%5(�1�Ԁ�
���wq`k�cF@�ͪe�0�i�h�� ����O�"
�i�&���d��<7�h�M���d��곟X�ֵA�

�Z�V��u�� ���ԧ��b�8�<_Uܢ<����Ʉ�i�d:���:W��A��i��9�M�8���DZף�Fpu��/]��N�����:�Iei�����k}�z�bWt?F�jt1�#����l�I���x�H3D��)�gf�m�@�ś[ .x� ��w���
y:�@g�]��w� (�qA��67�M��!W(lڸ�ZH�+�ࣃ�h��� ���G��l�i�G�N5�_�.y�Ek�'�0:/u� �c(�s%�ΕĒ�p_ӊ�2�[%8ݫkw>R�W�)?���.�	\
Ϊ,*<�����28�6G��G0��u
s0��E=���]�y��)KS�˔�[t�/etJg�OA�e����?ֻ#��3�L�.�F��@�Ypg�C�=�9�@3{u�r$(^T�����CʙC������[m�p�mH�CQW�),fN�$�Q����W���7X\,:����w��)��Ztr\;�X8-����vUMZ����UG�7�;�;��k����/a�Y��<|��m��%�Z���5Py�X7�=(������:[�[nJ�$�Ϥ"W$��������bEگC�Pzau�R�aw��1�EE�a�*�����M& �1��B��sJ;�m��|C�~�����v�M^��-�X0`�甝���.��K}BԷ.���'�� DES{'L���q���p�5Y^�W	�J� �&o��K�u-O$#�ZAy�1�B�h��O
����hһ�l(h2�&#�@�Ъ!P{ ����ӷCe\Ȓ��#�� e|W47ƀژ�s����y��H��0Á��M(�e�yT�zm�G�2l�b��O����9L���#Uw5l'��q<,�>��#*ϭ�zJ�=��)��K)��s/�8)c�o�:7��>�L�����mήɬ���JL@K8.@�e��(�":���i�A4zʝ�j��'�*w�x�mw'M�Ι�i���?��d�UA�B;�{�·��{zju��5N"}���:>��u�v/��Q ��������Īw�Tq�\�Q��ӌ��F�=��IW2�pʠlߖ�nh Dli�x��g@/��7�9[£ q�p?V̫]�1����ߙ�vNk�?*v�A�(|yB��WvC��5}���p3o�҈��,���w(�Wz.�.���j�d�Rl'��;�U8i�I�|�ՍE��d�'�e�M��D9���0�t^p��O�zX�ްų**����^�ߡ��5�t���,y�-d�L:��(?�{+��`^���G
mAH՚�f�X-8TS�ƌ]�i��|�yb����Jk��^�V4Bo��L�|y>D.�ዣ��DP��q�f�]ϳ&z�a)` 3 ��xs�,�]_,�������Sv�;�>����o�o�z�'�J	�P�f�hD��d?z�IՇM"��>=�#�IF�D�f�[M�`q	�v�:�NN\�'p��vrb�9Lh�	?��\-�`��w���E���S��N&�^t��r{G�tM��́ј� �i��e��c�N~��&�(�*�u��6�<nֵ��e�-�t�Y7�/���A�xͮ�7�ޮ�q�HD���nn����{�x�E��Jf>���8 ��F���`�_e1a�CZ������1�1�`�8	��n{���5�F��W)�Qa��ɄSD-v\���p�.*?lS��J�����f�2���qZX��(8��6�l���1S0��r����6�<�+=�]�0��3w,�7[Vܠr}ʟw��<�kIAnL���
͙�P�28�ns�oW��1A�I.�ӖӔw�c0����w�v�h�� �r��;q���KG �w�v��k�e�ǧ�wӭ#r�/)��i6.R�L��A�3j�5)�Z���1H�u�/C"���
��)RJ���=�f�{�AI�3�w�&Q���c\��
�x{=c-�^c�Ɗ��zp��*y�����A�|�� ֭�����j�`a>��	�ຜ
��W�@�,\b�Q��Ej�����X�Gj����d-�O�HH8Ή��?�:)v��A���Rb�F�B��Av����c���x]��z[j �܌����5.����_|�A�o��-�E�ܑ��d7<�h~��N�[��0r���'
���0���VF�����҃���8 �Jd �7V �W�욞˖*��"�F�&|x�lW�x�HV��m#�8�g���=�(�16��:�`�D�*k��5ڔ�X@�c8c���0"!��Q�B��:���%K'�+�~+���9�Nvp��ה2_M$�Lg%W�pj�}B�˷��;�`h�sJ���|P�����Ya��f�k~ /�i�?�����E���+ʻB��7'U�ϕ:�����Z�ud����&��:�����{�9N-P��i'�]/�ӇUwݶ�j�A�;Z���a�.W���v0���Ew�rqW����v�l��}�]�1��9�p!�'���ݽ�.�2y��@薊(LMC�j(61���� /Ѹ#V��{R^#9P(.�G�������}�����W�����#�j�5H�_����4YJH���8 �D����	q."�P瓝�)��g����	�Ӗ�t������]m�Dn��\>� �!��vn�x�)��F���>�����]�J��/m��^隡��e����{��yP��.̪�-ܞ)tv�n�24��̐7�=E� �j��>{��8��v��h��,@��U��p�j��t�@�R���od)�x�`�	�U�(�Y5�+�A�Y9��V*�+����c@h4�F�C�ٵ}�X����%�Ngu7�pف���v��=��x?Y�����.fK8�a��E
�O�w��#��2�U�K�;�ꃱ�q$�ч��-�"k��}|ג�*�w��"��'"�@�=��3�}�U�9�F8�8�v�ebpQ�,\�@,Ud'����s�b�;�*Q4�L�.v�U�:���z��c0��$������U�cټUZ�<�x���Ov�klW��٪��ׂ�D[�S�$1;<O]�<Y�J���0�'O'���잗7p:[H\����.��''������+(N�PO��aPW_U����'s���g����%s�a,�T�$�S�,~d�*�pة�$�*)�p���Hb�L&2�yF^hI�P:�F6��N8h�7*w�o���$;��]�g�b<�J�NC-*Yd��<IR��e4*c�·�lJ�4#r�>�L�4�Ewf��g���~�٬��9*j�{�l.��r|'��I��4~ ���h�7�ԝ�?�a5�iF�@�iӱ�	N��[��"�R�}EJ�N��4���3��h�N��pInLϟ�-�8!-o=��8�z�eG�u����`=����;�\�O^�@�ʐ7��q^�Y�H�>�ˋ\_O���%|����O'��X?>���.:9AE:*a:��*��t7�k�x�	��:M'w6����ɨ���0#���)�*g5_�U�w�:Yq��n:��la�����s�AT�K[Y6�Θh�'A�� 2/\�\��T�`�����3�~�
���O��x�.���G���o�X�������0�tO�h�(r4�ICt�8�a데����������Q�M �E�!#p����}�o��>��5Ĕ�qLhz�ş��#1�-jL��f��`����)���d4��E�l�֨ᗭ�Ƀ�����\�����u��	m�O����`|��I��3���k�Wp�K&�bb�i�޽{׍��L���?aӁ3ڍ�qr���=�~�sJ�4k��"����3�7O��}��$����G5X�t>������@C�Opw{����A���R���ݮ�^s�)���JZ��T*5V��z����̯^�$�xA�&s�|�w��KB��?
l_�$4Ǟ����_'̮W�(�_!T�9��0�2=l�&���>뛤�ӝ3�R��� �ś,s<[� f}�TA�\.�Z���*��{�X"k|L \5hS�p�O����aʷ\�M�bE�����zF��&"�k,�Ԅ���Kv�9^�
�Lfޕe*�'�),�sʀ�Z-(5�*SV��F�ս
슉 �釲__ v����\����]�������R�x��>���6BKP��d&u����m-v��C�W���8;�Y�S�;J�A�9h�#n֘����ӕo8V�z���t��t���R\&�Җ��;�&�P����<����"M9紂�[���c�vq�I������FJ����G�lG���g��wsm%e����W��t��R�ה�w6�Ӝ�vq�bIѵo���C�O�L�Ը�y�s�ܒ���cwd�bF��l�R�p��sJ��ޮ���ZǙ��վD�{��ܳaM'�����R.���XF�����3���st�=X(�B���q��y/��#�C��:'ݯ0�q�}������~7��w5��y�:���ߒ"����y�ѫE'K��������li�4��ê۠�g�}�����h�:ڸ�p�����᷏�����d5��|zx������yEXH�v4�^�X���M�~*�q/��9�̮k�a������ma>]»���'���0`��3م��C�&��cKR>o�n�p���X�d��a�g�v�R���q����P[7�r����}­
PS'�H���Y�"
�~`��,����9&xٮ��d'�О�=���
���& kg���mÆ��驒�Ǔ	J)S�2� 8�.�( jR��t�=���N��f߾�n{G�p0nA�� ���w�,��~�����jtQ�C�$f���x���gz����>���GR�\\\B�lh�a�eT,!HZo8b0i$��VO%@t�������{	���t#��;r������9|�nz��!_{���d�}N�AG�Yܑ�/*�2'������A ��*��r���X��bv)�D��3�T����o]@f��0Z촁�pBU���E�����d}V}��ʡ�/�t��m?Z\�+S3Hv����K.�6�٘���{�x��&�����5KV�V�7��m(���k��=md�
h�$C�6�:rrØdl��������Q2����A45q^�
�L-v ���x��C���\�I��ޑ?{�����|#�����;;r�G�rT�*��g�Ix+f����ύJ Ź��n9a��� �UVD�b	ߡ�ͥN�9̨�������{R+��^?q"�N�ĝ��=ۃlXM�]}E������-f�������Dl��;��S��K>[7�M+�QƽB��9�$.d?�T��%k~���r}�2t�}�s^O�����!["�V�8�(npH�q�{���p,'͡�UʸP�Rj���ى�T����l��'[2lbǵDr�c�n��3��UGsn��;
�>oK�Hs�e�>��%�5��b����h�}J�~&�	L����a��Һ�����9||�>���o��%*��6<u��e��Q�r^��J6�T͓��;Q�V��2�i�( ��ϬE�>�N E�ه�G�����{N��>�ؑm<eFqn*��AP��(��*�o-���IV�xҮ���K��lJn���.��v,��	!<{a�w���]��`]���u0���	m�,v��QZ�rG��\�W�m� (u�W\�9!��� ��m��>�ǡz[��r��:��0���K,w23�pp �:������۱�΅�d�~�?: ����B���|�������A;X`0+��o����Ѧr!c��u�6�<�#F��bEZ�,��9L�)�0L�����͎�K�* �&��O9�����9k�(0է��?��ؚ������	f:
��[�ܱ<'�G��HPn��WhY�pd4�C�jf$|�A܅r����۲���1�M�`]{��.�i�̗��nx0���
t=�j"nT(oV��s�Qqᜍ��� h��]	n�lP$�8�	ZHЮ �O�G"�hH�3�x��.��H~��K�#f�*����V`�_��K��k�rgB� SH�P&���BΪ82xH7��(P���T�����|�)g�:�q�v?�b�^�S�����w��c�x���5x�dB���(���MѾV�	/�ɚ)D��,[���=Y������Z��ɥ�KƗÞ�V��#�1�t�<�����.X0�b��>��8�*�P�3�/(n$Z�l��P��Bρ��!K\0�r.{�%]�e��&�/{�R�����UXF��m�ǵJ,v�5��.M����/Ч�~����%X��i9��[iV�ղ�XS�g�:	�Ír�C�Ҽ�����x�@�kRu��=|��<�����X�'DCJz����.��P��s��nΗ�%�W���;~ps���w��Ҝ#}k�d	�.�kr��Pf.ʬE��r`]S^���N�z&�V��(xp�rƢ5l����ۮ	55���ڙv�5�z��HwZ���l$B��(5�
Av��2�͊+=>�3#���.�������y#^�g�,�
�=�NA�#ES0
��;�u�*,l�>��fȡodb:&��
�k�c�W�t�0�j�	n�
<r�׃��q��Jz#��.�zO�}ɾ��@��e��~��;\^ݐ9�ryA)<��O���@fw�Ƈ�P�����E�s2K�1�E��2�K�YV�! 2f�B�eJ9�=	�E���������_���PM��[�����fZ?W1V�3.F�n!Q����H������N��{t:�Ǻ�ɘQ�$�xV��ևeS�d��f�Sl ��@ڦu���p��w���o�T�x�V�p�M֬J6������R�*d��	��ܞ�� �)�ޔ�
��͆��nd���F�+|W|»l�Ej�'�\R���J��c/�t<[rȦ��`���iڐ��ݲ�6�A�4�J��|�f1�Jˊ�۶q>��4
����'9�(��#ѭyR�b��@:5�W��r_Q�m��RDŨ�`�łePRo������J�o�Pk��d���߶a��P��]�[��VQy����;8,v�#��@SÚ������:t�$KRf�6ƾ�q�W���biv}z�8qE#>9�PM��k@��J�*��-k��;�����vu��0*�I������p�C`�;��O�=sLc���;VBo�	,x%���z8���ʑ;f1������Y5���� ��0��<������)�¼�����s�`Y�M�R���^�1 �'�a�� gĂ�]��J6B4�A뚎�=�� O�u$����?��/�>=�n��?�SP����l���BM�i��'�5�(�c+XM�P�|�����^^^vr�,�s���㱓ѳ�9p�Mp(���i�(�_��I:Ę����4�A`x-�"�4	�-�{�{�`ƅ�f�9L�	�΢o�B�ff�5i�Q�Fi[�N�j7��2�S��7{8:;��K�QkH������cB�	���a�+u|ax���)VM�%�A��f�0g�ִ�Ιo_�����؛�?��e1Ъ�%�
7F������Nw����Cc��(� xA��a��#�5�*ͺ���o0����ydu�{�h�ܮdz\I���v g&x`Ek�p���p�q��)N�kW�+�WG�.�ǻ;�4��_��@0�ㆾ��_���6g>��S?:o�Q�������y孠���}���@���_s��EEIiv�J�z��N��wX
w���fdôtuj�YJ*ec�S��b&5eN.��+������@���BP�cm�5����x�>��ϸ2xgzر�4���P����Eb/t����FD1}��!�7��탤�h8���v�K�!���S��d�I݅v���P')����o�V�E�c�K���?�Oˇ-w� s�_����r��R��\^���l����zQ�ŀڲ*T6���ϕX3�rwB�jp�ЋV���x��b�²\O+���S_��Θ��J�I� ju�}˱u4��1�$�;�gJ$$��;�{����
�Ɗ0g��� �偔.$0��𡢝�	e�b�5ϳq�jڜ����#�3���s��B��ap���|�𻸁�dɳ��������(ץf1��<��;=맓��x���W.�rb�����_�:M8�1��1bQ�3T��w��>��g��B�S&����=�h���o� +�$'�5����W�q�*V총��i��}}��-��5|��w��'��م���0_L;���G����|J�W��;�gJ$bՉTi���V�0���B���8l݋ ]��{��'7�)vv$��6I!��W��N�:7�gC�՞�C��d�b��GV �*�.ݧ��-.��D�@]2O%m�i�-q���r���k��1N�ն�J#R;V�]��e�t�C�ｒhu\�|�O!�J,Ŧ�8
C��7��/)���|5�Bý:DT3�0�B�NF������uK���+��%Y�  Beͻw8�Z���-i���5k�1 [��)����byA��)yP���n���?���wr�B@��%�U3Pⵣ**��Z�c�A�CUvR��(����3�:?�S�'!G��K�CV!qF��#}��gj��5�:^T"���\j�C�����n��ˇUu1F��,u�,X��l��R[Z`ֲ*�QU�h�&��y��U�$�U">��P�X��-��ʶ#�
�ɻ�"I��]|H���}�`H.;?PrkPMXK>�k����F2�%V+2kQ2y��R�a4��.*��+$��k�zg.P���b}�vIĤ֒�\ `�ʜ��=X�z9(w,}���d�����R�WR�iP�8g�ź�/�!���G�[%1Ѝf��W=N��"������$x��#�Nx�Dp��{�2
1փ��(���{�B�*��Q�9�Kt�z|x���~�]ϻֈi�ɜ>���pE�@辀�[r��0�U����{�C�1����<�4�üF?��y�)U���5v��]~&���>�������M�m�tG��[��N8�4ʃ��S�Qy�sR����x.�#jZ�*5�!�C��H��V:��}�����á��������@6ϙ�k�b�%��0T��5�c�~�F1P�U���Ļr����~:'�T��1tM'+�n�?�װŘ>M'
�av�c�<W�[�C\�0�ѳf \�n���Wi�zr/�o�p�T9� uŮ#�V���0�9��t�^��ـD�i4�е�I�)?��s̠���i{&�sf��_g��3J�����g��	-����WG
M���]�/~&�>���	}��\\b:��a�{��3H�	^��`��z] 9��C�h�S� B+��w_������~��_����I�_v��P�0{E����U@���RN�#滮��՞��������\�7Jި9�ɲ��
�U��8Q;^ss��R ����W�r$�ld��}�a���~���p��6����T;G�7FH��I\���ݯֵ��ʅ��5X[5����<U|w��BP�(��t����G$M��fZR}* �=�[j���9��Z I+��F-�$Ùo!�Ae�����]�0��Iʇ��9	�SS��k*�p�چ٤ڨp�)m��O�)y_�~y1}Ƕ�g7����J���N2ú���!K���]mz'��4� ��-�R�p��}w�6�%5`6_���{��~OV(,=<>����9+���X�eʂ���i�0�w=p�/\�V�V32W,w�YeP'��5�lέ^��z��l{]Ა��W+�o��*��k��-X�^Ku��Zcŉ7�BkgDc�Y��l�#xw�d��7�l�t$kh���
�gl��8uhQ��2�sS�X����[M��[���n]�2Hm!�߆�Ç��=<��z���X�~�VF��q�Y�[�1�,�M�$���6�i�X�<A�Ř�S ؎У��|��<fW��;���|�rA.��*#$�|�X{T{ Ѥ00��Z�+�>�J�4��* .�2@��I�-���yN�ů����yC�+07Yӷ�p&C���wvw�(u|��oQn�3����+��{_��=P���lɽ	�l���@.S��b���}�4��x�����nQ?tD����0��R��Ɠ���q@i��ف��tA�S����Od����g�����C?O"^5�k�R�Ҭ[�ꏽ�
ё�u�/V(�.�L^�~t�h�ܩ���?xC#޼���/oA`aF�s̊�u�aw����w�H����im�t�73닡�V����z+���� �B�������5����9���V8q�Q�!�D���L�=�l�V)�Rǁnı{O����"���ͳ]�F������0W�):�v4�r�h�M:QB�p����u�/T��@U��!Ȳ�DQ�[HXF�6�+�������?�8G���n��Rm��յS	�X��̰96���d�T�F�����A�0�������y�iKq*|'���ͬ���=e�����9ae��%�Č`��K 6�/��uPVX�.`�XQ{P�;ٷ�w��a(�)|��yLB�W�@��$f����1!:;�'�����Sb�$+���u��_F�ȹT@�2͎�FO���/U�t��M�cѓ@K�&�S����\�8����g�L����$��V��pB����w5�B��/�J�޸.��V8�֊4�'�~���л2Om=���x:~��1"��|���\�cpO>�&̸TUa	M�!�c���Va��1�]C���~C1?\���\�����5i��I�>��ȝ+O�v��M����dd^�+K�Q7��S�N�j������Y�
p��������l�w�r@�g]�z_@��-��КjX&ug�Q+���]�_��M� v�/��s��f�5���KF*\�!������\��ݢ�; 4%��ZcӮ�5햑rGͷ%�Q]��w+�T�P!ḽ��o_?��/_��ᎂ%S�4��ğ�NM�iC��(1�k��_��_���翺O����R)o��)u98�q�z^�"}�rLA���N�;?� <���Ĝc��6,�4 -A>��[�Y��	)+��֍�/?�xx��b�@FkƵ�X���M�踑���3�wtl�:b$/��j��Ǌ	H\��V�b'��������
��Z8�߶����敭��4Ȃ3���J�����C�q%	m��7]�x�ƿ��M7d:��I��@5e�'q�F!�b��$�Be�.6���.�!�N��5.πR�TF�
���z��Z�ϻ��k�y�߽ǖ0�b�b��)�*yhi�	�́Ҟ(��2{^���l��;�-��S�Y�uP�!DJ�Z�=�=b.N�r��/M��vc3�'g�I7ly��/C�|�~?@��Z~��Hn�����ſ~	T?S�ܳ#ʓ��38�������}$�r�k�}8������9LY>�:zԝ�<�v�}G󦰘/H�zT�S���j@yu�Bd�BAu$�$ٷ0���@4�,�PiMJ��ֶ�,!k%�Iwnʩs��J1|�G�%+"��-T��m���ph���Q^+D����z�K5u��3UŸ#�&=���o�$a��O�8P�a���g���k59�8���Cf��)^�1��.Lmġ�ETq�쾲+��!��˵�.�h�n"(�@�ӆ�F5���}�Jʖ���.1!��b���s��3�{����hE�����-r�����Z��:��b�	�=�0�������9�J\�_��T���K���_�睡gϩ�WFN�Y��'�ZO$�b���]�W�	���%����s�W�.>ʅx�ZHew��'O���ϲ�O~��yW���Uv>�Lv�R7#v�⾡���X�pp�h)��U�Z����Bn�LEH�uS��R?�w����?�%�Hz&V5I�.뎕!A�^���Q1�`7�8�$?6b����p��e4�&���t�=42����T���xJ}>�(�Ք�S�o�[r��Ѵ���ccbF2�.�b�L�{�����D��kIӋ6�E��]=��K��~O��Q@�g�:<����OO���7
F���I�kΆ�XID;�-w�{�@���?�ZA_�3J��A-�������2av�_M��f�����
'v|���E�aTZ-O�9��WF�%�bx�$�B�/e�
��
���|��E� a�ѡ��t���@-��eG�&�DZބ�X~O�c� ED�t}}M�̟���L�%�ZM1(������a�H1�Z�p��X�,C��~��*I>7NU�<����7���
�U��&frd9(@2�;�k�D.0��~���B��2<T�c�:Ef"�;�mqD�s.�y�4��+��vCud�־�o,U0�-�1�L�A��>\���t�B!g:/`��:����5*3�7�Û�|٭�����0K*d�u�|�Zt�f�-j$���������c�� ����U\�O��y��ދ��Y����(����总i�y�I�h"������D�����O,�UF�O.`1T���<UDZgz3A��Ji���B?�ČF�8��f� �%*wTYslLc@\y�lBD+�##e/y�A��bD0����ʅ�����@�7i�Ћ�\���!��&�Ry�i�\�3���&qZ'Hs��+�덿3B�\�}p[��Qɓ�-����:�J}��q�4Σ6��w�.ZѢ�C�~��MJ��;������
MǏ���m�X���˛eԱ�1R<�g�bk"���AWr��Ê����\tB�ǀ���T�R]�f3�����y6�r*`��y�;�9����b������p�-�~�#W���#g �8��a�x�<7MP �9[(n��ە>�=�ޚ�k���)C1a8�Q�$4tLy�E���`�����K���ܒ�E�4u�	-�?rȋ鴂�b������ﰼ�N�j���+<޽�IG�;��o��|:���ط����1��<p�iG�n��a5_��~��	>v����`uyA1|Ȓc�t|c^;���z��ۇ{h�`��OA���H��W`L@�X�_)~���^�YR�-���o:���a�iO/�R�����F�w��<����:g�Ms�:��2Z��2M'�2J�Ԭ��
���a�?��94T�ODicj�m��D���x�:鏡�V��q���b��/'f��.���g�n���9�YU���5�}��J�/.��1�L�-�n���Q��5��o��[		�5�/� ǸX�O��k��-IS9Ի֠&����N5̠�&�yQz����30���aŴ�q��� ��:��k��̜��ʕO��������:Ok�s��[��p��oJ�����wů�T�g������5vVQ�\.����>��~ja��:W��uE�N�Qls,J�@�Y����=��K,�p�彪,H�-�6������j��晡=Z=��/��%���?o�XIcDۢ"@K���"�=�s�����T�ߨ�q�[E��3O�m�ך� �|*��]���/�T���i�:�8Œy[E����]�Ex@A1)�?h�duO�\fxs$�1Usql⛁��J���<-��|ڙ5G�Ϗ���ƣ��c'�t�c������5+l��.��ӂ3�y���M%u�&�N]ӆ.n|�C����[�/�^�i�O�p��)� �1�J.Q�����"
cFm��1H�������{�%Y�|��,M�S�C,��b!^izw_����8C����2�L�yg�����l�+5����~]��7svL!���_$P)�kz�-ڝ&�v�?y���1=R�]����`lkoQ������J�[�n�&N�V�*�-ͫ	nt�&UC��٣.��n�a9[���(v*XL��C)��������$����)Z86�6.�on`y��LW����u[X,�X-i3�i]^^»w����x��V����W��м�mH;�B��������D��w*�@@���!G�:�0# 掯;�Ty?�>]'�/	8��Z +o!(w@�<4v�b���[%N��ݟ)	s�֞_���<�����-NثvN�aV�'b�?�^�(:�-�ϟ3V�)W�ٙ�&%�f���S�9��
�U ne�CY�;��A̘��u~ٓ��[��(�"ؓ �d;/'�C;Ml��>�:���O�}.s\�Y%�|B�8�NC�w8����� )� (3�#[�8*��״*uDU�_J�3 �ck�g7�[�c6����c%��^3Nd����9���2=���=5�����e�?˔.*�c;l�
��{�J����U�z�#F��C��Xq,+�����x�ؓ��v�KoK�{��!>Û� 
&�Z��J���EH�.7r���O��]Ye4%Ʒ�y�='p3�H1[F�O�;㺑�RAnڞ��B��}���}���<Z�����Z6T�9HdH��@).b���U�C�i���x���U���*�d��o��#Z�"�5QT"_�i��ӹ�k6���q����(� ������Z���n�B:o�`����S*.�,�"5C�SƮ��v���=��<>�B�ƲNn�ݐ ���;���؁2�tC�^�U��5nL=Qj�������\�p�
-�0�'��A-��1w�"���=	cC�qOCV�l�~��%�M�γ<$�(}�8po�S=�<)����@��^�<���>&�m�9�^�����X�S�NoԜ�!�����Z�%5T�srqr�h��ݐT^�	��S~N�lm�p�*g��(�L�q���.�-�}S^«'Z��m�ǉ��Wb�BJ�(wՌh�tڐ�b�Ѹ��[hѳh�ZL���
f�z�a����6;�m N���#|D�f t���]w��@�KTy�࿿������?�O�'x��>��	��?��,/���#���t�`��dN����:v�B%O�<h�p�Ɣ�������a�	Ͼg�VY9���rG�kM�N¯��BR��;q`�Rg�������D ŉ� �Q!�YB��u!��Lb��}�"�W$Jy����ܒ�c��eJ4�����# �����Œ7d�u�����*B#�Jד~o�`�S����f��q{N�7uy�[&�� ���뜒�&-�y_���]��� ��/~��翉Uw���éS)�
�7�|��Ww���o7x�'l����9�:��7~Y��M+]�H�sp�3P��F��m_T���D Fa����G��̵D�5��8D�Q)��+u����u�(5^D	fSU.~������9&QEEe�=����ò \v�7��nX�zN�50�~,m.��{ ח.*��Xm��+|?����^Y{�`ށ�Sk����5VRW�*�M�0�Uа��8ƍq�j`1[�[�i�*j�f����f������߾~��0P��Tm�0Ņ��c�&�q��ň�E�Z�ɮ�m�:ր.G
�$pN�Cz��#�qH��'��E�0HG�H�G����_˳�F�	���γ�([��ye��m�0�WK���h��?r��"}9����e�=���?��#D����S�Ո��f8�<)z�� ���G����;�|Vu4������+���"+�i�O��)�4ps��&�Q�t��s��F�?�������ۯ��
�]�&������b777p� �w���>�eP�;����<AbTP%������	���^&�+��z:�l<���N����G9$~oK�I�wh5������/^�\"�� ����kM�U��F�?�ʥtǶ>�~���N>d��!��(�®lF��j��_�#
��5���|��Ee��I�O6�a~�[�~E`���q\�H��U�;r���E�G�������W,��Ճ�kn������;�/)A�(���bi� ��#�`�8psB����,�)R��7����aa�i�����s
Q�Jv楃*�x�S�1�G�R�{�e^��bBc�XW�X��O�D�����CW�M)I'�r�y�5���|���x�ݹ�T�$�, ukb}��v�#�3XͦSڭ���V��;��<�
� ���v��1zx&[�h�'t�R>�MB� �}��L3��V�9�/~1橊�{��7�=c�Z�u6�b�
z�E�$8�s/�/WFy���I�~��K�*=���~��JԕEy)uJݛ��(�ݩ��/Z^�T;8�z�+h녯ǲ��m����<ޯ��<v����m�i����>|��o���c��7��eY� fAZH��*O
��_��?�|�������O��Ǐ�'�>�`��;�����!׫��/Ws�;�c�L�~���
�(��}��9�$�h͏��Nna���Hj2s�P�a�i�mÀj5�� EH���J;��z�h)~3p~�<�<��/Z�
��G�'�_	�KZZ����{�M�������� �}v�dA�*t�h�9T���YBJ��5�='A��R�2�g*����Rqخ��%��^(P,�^�YX^��
�ʱ�q��<{�_��=���)?��vae]���1z;>��;���^�x�o�:���K<�������9��_�pG.γ2]X}�+��^xө�ZR���EJ�%��x]+;!n��wJzd�0J��=i�� �6��x�G����1�t"�.&����o@h���']z�=������Jo��7X��� ;�i	�� �Vp��.�F\����J
���	�T��.S���@�RLi�b@-ٮ�9���E���%�5r�.X8�}U��s&O��g�u�R�g>ؿ�eLR6+eK*��s^���u_����P���]4�	�ݫ���$�B;�X���;v�8�W-Ĺ2�ғm�\a�mQ�$~�0�<N�G�}��(��aڊJ�i=��vM��Ȣ�XOwO�Ѿ�����R\���+���`L������+�^��hAK�͖㤢��{��հX,�ju	��%Y��cM��5e��k�ΨUЂf[�;y'e�Ȃ��~�3d�@�Eb�K�kd��)y6x�4^B�Ĥ�-z�q���Z�Dd��2iʁ_�X�~�k�v�0�Ӿ0�\R:v�)#�9wqz��]����(�u�C?��Yw� 2$���9����	bI�����P�%%��	C�!�b�=o�{����s�֏@�?m֙����ޏ���yJo�X���R޳��2�*��l@PhQ1�y/���+w��S	 �G�;�]SҊ儶��[�?*j��H�X�W�zŊ��=��1��*T��7 ���ª�Bs\�|���4>`N�|��U�����[ڌ�(�.���)���P��%˔|������I)�Օ�GC)��h�C1u<�T���̛��A���p�Úh)�VM�T�	X�n$���#W��1�3�7\I4���
��C؉� ��(m���J&�h���e��JE�:Q	`���Ց���ō���)�n��	�߁�<�j?rt�b�*u�G2AD��&0�8�:��MU�.]A�݅��*���x��^7��صح����W���l��f�Z]�b>1i=z1��8�9Z-�g��R���t	�����(sw��Ί3o�:z��i+��_X�<��70=�`�N�@���DU�|8���o�`�+�2��9������Ա���TE��+�(h����x �h)���Ç��@�h��LR�s��1�N���XQ��*����8�JJ�tE��S�:{:�<�������?U�᎜*�M�΁_A�tn^��� ��N6Fc茗���Ov}��2uz�gE�V�(C�BC�}9�J��H��+q끌��J�jР����+�"7	X[��fJ�{�����5��Xym�b+��5�"�����y��8獖���_�����*o�FɊ͠hRrHj��]`���ś�5�NUyQ�4a�`��]0���Xq̋�2xJݔ������xOj��A�C�R�Vp��"}�i�ϙw!v(0�����f>$�`Řl��Ղ%�o�~��XR�D���2cl�����U�͆�X�n���>�I�� QD��9��ب��)��M���M-Qꠎ�=�7����H����F-����0���LC���
y>)e�=<�7���W��?��vX��o���a��;mEY�.�.�f��O���Y���:�l�m����D���=�-.��g{���jE|�,AbC��ġ�������1vT�LI�N�b��:g��o�p�;JF>m�D��*w�G��u��	`ߑr������2���N&�'�/W�<�Y�gI��?#��/_�qS&�'�!֎���kJ���q�19hw���雂�:�5|���rŝq~l�<W��u�[bm�S��|�9���~�2{~D�C��n-�<!�����aT^��L��;��O�

+g�5�*Z��[!�6��_	���JD�N�k�<&Z�f�|�'�D��,�8�P�n+�+�Gd��� �\���&U�c��C����{�מ�<y9H���Y��\@�^,�f��--������S33��$tԴ�MȆ�kG2VQ e�>� VֶM+�:+����1�j0Y����y�Ep�P��Q8.Z���T�&a)��M'�m�>��i����QX4�q�\P�����[�!��(K���cn�]M�E�}�]1Y_j�:y�׵�qG�OT�,���sB�>��+gb�9R��i=1A��J��j�?,`�r0_�&�epsq��|R����Y������&�f:���������)\v�q�6��c��3p�)ջ5�� �/�*�0�2*yP�s���+gQ��[T�,�3�M��l�[�����ua�HS����:��@^M����O=g/���>0]W=��a��m��q��`����#�<�M�ʓ8�m�Ր�\;Cn黫��y$�<��"!*t��t�������cm����M��a�Q �aUj%ꅞ�$Em��,��OS܍��i���d*�|��B\�Mp�T�Y����(�qv�������},<� bd�Ǐ^��|��|��Ҋ����ͥ���yu�O��a)��#o�����5�'��dq��Z����G@��@�.������X9�7T����ĞU\E�oU��.['��ʷ<��X_�֮��N�9�� WY��l%UjH�M´������݁,�;mL���(iɓ�x�~;A��+%�0�
9m�)^�5ȏ��c��s)����Q
*�~k5��/\��I�w�U��.�KF��_��d�U���ʆ��V6y���=G�-��$.FLHt���u��q���:�K�T��!����HyN{Ţ�V�d`EN��:s�n����C�W,��z�������P<M^߰Y�7�&f���L8��AIk���Hl�dW~��	�V{��w�$<�4�:� W�	F8��������9�N�=���N����9��0�;z5�h�l�����pu3����]]�r2�մ;�X�XW�S�0������� ��)��/��byI�\]^����)f����K���I�;hc�Q{;�ؐ�U��ڑr�^C����Z�7�*̵�ة� )�%�Jsb�Y�����9�n�la������-yP�Sͻϒs�Of��Aш�XC�zPAP b>] �]�q�)�Z���'�<s(�2a��:w��8�X���0�DEV$r���[��r'.og���t�.����Z}t��8�I�/)�*��oە^�Z���?c�zg���Y�k���< �Pt򣲩���b!��{�X���v�9��\�o8d������O�]下Qq�u��T���2Cg�>�#C�l��Iw��Nk�S��H,ש�|�����u��*�4�U����|��*8T�Kfܣ������S����&�(�kZ�;K?��.P�U[�d�0��Q>̝gl�3&�ɼ:2����7"E�b��N	3���o�R�IcI/���o�xc�d�(O+-]]�6n����Ӝ��h�q�ϋ�/9F%�A6y�,�0�yA�+�iY�Zb��t1�[���|�W!P�zl+��q9if=�ޗj��O|S�I�3��{F+}yM�Fq��ȈZ���xT3~��_��벛+F���7@�˽�@�6��Cʝ�Un�0�m�3���@�����&�����Zb���-d�sG�&��]�0�o������v�	ܾ�[��@���{��n���&�������ܧ.�+X�V���)vμ;�����֛'��T�b9z���C˿I��հ&��3x	�t��w�R׏� p��yb��M,�d�v���&��T!?\���9�4�UO�$5��ķ:9
�	�x�h�޴8 -tO�y)�\��~��z�S��U*�p� CP_0SГO��K'�K&���C����t>����ǿ.�����nq?j�<�2a畊�V�;C�S� ��R�ť�7)��f��9��<���»��b|�^̄�J{���+7!zb��� :误>=�K��3t��9�U������X\�"9i-��
sR�Ш�X�R�!��Z���-�m�zΖ��?��>LxK��z���r�<~n;6��9e\lw=ٮ��	���h�k�?M��bf��TQ^�����|+[�뱸�;��G���S�s������e������������^#7��li��iI�J�1Q��P�Τ��G��?±�FǕ|�_�t#W���&�y��'�E��A�:�7Ʊ:4p�e����Tm���Na6E���I�}Z�PZ�	L�T���������u�滻��_��ڣ+�>~��o`9��|1�w��w��X;k�۸����h#i}�����r�ZLA�����p�B�<�wX���f�H;̮�u�!_W�����/M0��v�r�i��TC��=t��t��5`q�%����2=�Λ�C�sTxq�����?����ݫ%8�����JI|�O�`:�3~��R�'����KT��kP�[�؉��Jh������F�5��~�ٿ?e�R��tU��R�C��h7����
c8���������搁��^p�^2�fWx�V{�*�V����*"�����m��;V��֑?ݒ	��Q��U�&q>��n$h͠�G|��h�m�!/�Y����ɚk�����(⪔�<��U��7�y�.�3������~9N'#��&��H��̡d�6���P����7^C$��9c�k�����*>���v��F)d"�����fC2S����/|;��0�_X� Җ�����h�&��h��s�̇�(V�"{��g�gt�r$���Vo�c�u�0�߾��9Xo<m&��L0�/X�1i�k>�ì�C�����%,VK�6�������a���n����h:������T�kv0[�`�ݐ������-Y.��p�� U�g�R�*v	Y
��<<Y@6}U��\�T�L�S6���u�B՞b�;��\:���`�ظZt��*c�3�+|̢f%����\q�K�^E�� �����_>�#��yúB�K%��J�ړ�yV)Hk:��R��ucS����8�[Hr�8�˲?@�;ʴ���<
2Dz}Yt9��z���m�i��"Ш���흱z� ��\f�C�o�|v�+#�a�sK���h�2-Zx@8���u�����=<M9ܣn���=OwDQ��m�|�ndw\�uެ��	ݵ}���Њ��=�)<��ñ��/'��2�~�����"a
�%��&w��Z0�v�[��:)$�p��ګ*��k|;_���6<ǅ�����-�mʱ9:Ԧ��J�4#��%��}ے�l7r��r�{�%J���aŢX>��D�0�y�+�!�h�'WF�F3؄����?6�q��Vk�׼:�8`:�b�(1r�7:���e4�����o�?a-�y�^��*�=�7��}�a����PQ��͘>��C
���a��I�2�;v�l���ܦ�Q�C�|:�鬻f��md�s��������;|�����
�]�(~��M���\���F�)����cr���z��e��v����w���'����>�`�_����#)�(�`��v����'�O�p�.��N2b�e��?��$S���)g[O~���&���Ԥԩ����>ȟ�&D�p$�D��.���a�o�GP]�MN�wh���7>QC�(8i{�H�ÆNy!��
G]�e@��V@*��Z%>�U�e-�o�Yr����K �:j��(���
�=~<�<��+s*���^�m�*=~f��������LA�0���q�j� Vc�r���|AI�y�Wy^��<<:}�`HQ��4m3EF�
�����Kx�O+�{d�d����3�	v���J�X��5>�-	áP>h��x��ы`)b?'������q6��P�1p�г
�:��ьX5fêk3�Ȏ��k��i��a]1)�r�L���)�9�\ἧ椝+�<�!�{�51d�=�=9�Z��z;�Õnh�d�n'�S�����K#�c�5Q�-��ҊN����n����q.�>-i����$`|��1�9B����g<�$�����<����}Jr�D��"���* U�)��w줇缽��Ij�E����2H�$&�9�:�����,7 ��-ُ�]�Uh�	וD���2dP!HF)���T��&�nYMZ�F�������}h`򹅛�xs��%\�p��ՍG�`�K��>B5Fw��=>ݓ�Z�<m6���|F�X7�W���n�^?���=���[ء�`֬%P0eR�� XL�}��dA<����Lb�Ƅ��qD������>����<�=A�[�jyr��G'�B�-��H���JFI�&L"*wl��ۿ���s�yy. ۃ�SU��BD�3V��E	�=4 X	��:N��,2�;�L"S<�d��d7�KW�}l�Z�!HX�9��H��D�O���e�����/=�y#���������yQ�q�+�h׫"Q���g=��8�,�?�#���Ù� ?e���o��T?����^��:=�[V'+؎ܓ�;Ѓ�`��f��z�����/��?W`��(��V���j�rap۳��_��OȎF��e4>��=U�c�?�@r\���6
�bߒ�oRqu��9�#ﹱ�҅5�_���@����E��CC��}=ޠx8c��m�����j,P��JBB
��ܡ��q[���m���z�S��);�9�
d�B�&��\[�����'+J�-�D�Sɺj��+�g�M�,�����u�LF��b5�o\���*�b�,9������* v��_�aEܳC6^����;�������m0�����[�!���<�Dz��E���B4}�j��M]w��}��<�@J�鷧'K(�v�|I�3���!ti���
+�%r��x�o������v����a����[�|�}�Op�y _y��|��
�� ���)�LՎ2ea��W�kV�����b���k��0�xw=��龣5^�qw�]G���C�
�\Y.f��	aq�Ŏ7o���GM$��YߴX�T;�z�j
ͬ��];���a�Oս���2�]�X�C�4of�O��y� � ��Y��t�e(ϑ����Q��!�G���4RA�y1;��Y� |&���=�%S߯����,
c�V���(�.���f*�������P�O� �w�Y�m�JK�,���'��y� Q��� �W����'�dl���<ﱣ���0��N��nr������0��S*�3D�EW����Ⱦ���K��KJ��͓��(���K�3P�&2����]�!s���#�!G)����<��)�DZ�T6�g�����ci�qXͅ���%��`�]2�7ތk����`�ø�0��ͰB�����y仱�V�2&h�\+aH�<��J�Xi�o�+̄�PU�KHV+�J6��8;��/a�Z2f������)�]�G�1���BX?\�����	�t<�=n�1��FDqIi�����X^��gU>���Dp�����^B�K
�@as��kg�'�qw��s��S�f~�*�����Ч���ǌs����`'���]�y�iv��=N�*R�����
��ϛ�5��k{V�0;G�>��Xg�����9��Hhp�ܷ<5�(e���st��<�D�:%vFP�$���3k_}�<c����3��wqn%ǹ���'��P������z��ۻ,ۤ�1p �y/�d���c_VxZ��]ʨ��Ió����?�֧)�ۂ�cz��|��~a�'��o�;���Mw+��Sf���xܮ�n�HI��z���7R�L�9L�3�&T�������Φ<��{�_tעAZ�td�@�B[�P yl��x�R��@��'pp�١��EV�B>0J=@���\���z����&���Ω�e��ן`6�������{�
�|���/{x���o.%N��<�X��t)a'�į]�La�U37t~p�`6f��{��VN�Y�!�m;sRm��9<5c g
 ��\w�.�G��VC��U���L+	���j-���NK5q4ƪLkNq��If�m��~������%t�Ytbj*��� ��Z��h�1@��H�&R�)0��{=����u6���n���
@��1Ad����Ocm�T	�2��@��=?�GLe"��W�jܽ�����~�����Pݶ*�r?b����}^���1ф�Τ�U?U�g���� .�� T+���?z?�9Tu��m�)+.����u�u�a�����%4��lڇԡ���d�~@��m��+%�2s��)��w��:�x\��;��AM���sA M�	H/P.�Xi}^�H�}p��:�*K��Q!z
fxƹ�(t,nca,w Z�����#+��D� ��X~qDh6-Pz�vI�4w���&�$��{��K_h��T�}�d��������<&�صe�ܚ��!/^_���BZL��분oDs��8�w3�En�f��uVWD�)f�(�x�h}�X��MB�3��B�(3�f
��uD���:�1�$��Q*��3g]`CЂ�6��
��Y���
�L�>-*;R����$��MY�}T��#w���!Q�o��/�X��R�@���bɊ]!u|��>YW|�畳�E�B� ���]ϙ��<3�|v�q��6��qR0���z�����0�� ��5�!��i��Ww�s��5�y��	>S�C��Kp�{Bؓ�B����ҩ��cc]��|�d3<��ž�o��[-G�����~���Aa��{^�5�z	< ���q�ħ�|z&b?����-{A	��W��^�3^��C�3������~
yE>�X�9�"���ƎӰ��r��Oo�<7���Qi������]�r-6[7�b��ŧJ�����H�O��h�tF�4�FU���?�*��'��r�%�S�9H~�vW`����	Y��c_����ێ�0?[��#]3��4�g2��NI����;l���W8�{X������$�t����o_��ᎂ)#v�^#wm��1^O����m�N8`��D�'\�u%
�e��sf�)Y�L}�}>��lp�͘�by�}n`6{��r	����x��&��;�#�l���&Ð��(V�����7uN >)��OTH�w����_��j��!�b�*u��Lv2�`��<"��2lb�N,
���F�;"Tԉ�ڴ;�����l��" ��Ϭk6Wk��<v��
E�fK?�����m�S�����5(g����A6�B��̂��+�  �>�:��9W�7%��%�=���]�P��=��V��¤�*4e�K�TT�$�ÜS��%8����U�a@WQ�C��0��4��Ut�C�Tqv;4D��c��r�֬� �k�;�N0*������t��!)Kp�jV�U�u;�md<�2���V�P�(~�ʱOi��.����	2�LF�Lv<b����&kQ�h�c��Њ+�q25�T�n-���H��'�O(p�/�U�hR���c�eJQ�;�eo�%}�O�8���=[�E1(�2o��4���@Y�-�.�C ��o�+w�ۧd�tA
&�e��.΂�؀\y��6�׎��V��<#;��Ky�t��t
�g����6i_��O�1�����L[9剆c!�Z6� h�l�U+�����J�鷸��J�+$�^3^���e��6�b*aQ�0:&k�׊��ę�w�?���X�%;Wүz���Q�����]�9��ǐ/��h֢V�t�s�w�6(Fp��n9tvD�V��>vul���+�3e*]��(yd.��e(rb!b��5�v��X�4�*�nۄDs�>Gؗ�]��w�0wJN��_��N,囕�X�'4:T�(�	��~�n���4G&a�P�&nX���3�t���Ob����-�� j��^�#�x� <��P�<���ڂr�>�YE�����^�� �Vᔐr1�K�̞U�&�u�y��%S����_gfa �]�|Y�7@���J�o��  ��IDAT���+�4nd���0����:�T�~���S9�wMxFznT�v�8����i��z��~�֘sр _���͎K��9d��gzf��ˌyQ�ac��Z̾�MG�*�Cm�����v�MW��L�ԑ9�ڡM���;siO�<�n���������od��Z�t��̗K
��֋�e�v�	��n��d � kq��Ɋ/b᫢�樀�(��g�\������Ng@�#<��c�6͆��y�<��a���>���6kWi�+�>�<����̒��ƨ4)f&4/ L�F�˸sI
��7�2�&\�c	f�]-�:�Y$�XmIə�7�ߧfŔo'��+�L齻1V ҍ9�a
����<?�*���1"�� ��*`q�@F��r,�U�.��e*�s�&m?�V%@��0

���^bD�w�p"
7Vt4q�,�`^v��m����/c��B|*��wj�,��7�@Ĕ���PIG��
�tQ�[+'�bJ!P�p
Bf���ՠ�9j��ʎ=VSE���=:'�WD���0,ʤ�(+,Iͣ�Y���2�J-Q��4�H�g�qb8QL��Tʭ�J&�H�y_���9���V8V�S�c�{�{Y���*���b �
ע�T�V�b[���M��|��&�JP~� <��N�8�➄7�)�՛��pq�a�Fۛ�3��I���������V+
=�&U�H��(�-�]����`��e� XZ���^�^�^��yF-
���z\��5������g�O����X�ʳ�Nۡ�RiY����I�7-n|X�<������F2��Nj��֭�FٿBjA�+R�7%�c;"��{(�i
�SCZ�7Ǌ�VC������'9�8�Յ%�W��&la�}�
�� ��A��L��7\�0ywǧǿ��7cyz�Z���Lb�ஊAr��m��J�������Q�-Cc��	}CGH�D�<N�tș�<ަ(�q*g�����:�êЉ��L���Q9��6�/��kE���c�Vc�!��ВsN����&�q#I��9�8II�YUݽ������N�V��+.>��r$��Y���@ ���ٳ�v�j�{_�s��¨�r���:���Q�Mo5���#N�����������E�.<�E7��������9Й����͍ԗ����>C�Lߟ�����R����mM-�T���_.�wG���>}޲�5���	M���t6����f�c@h���6��'VQ�Hs-~m�Y'��h���B���s�;Ȃ�A��Z	��G	�g}��H�ˉ�����c�A����Rp��c30\p����pk�ܔbd"�	��웼�*��:p�Wc���\%	�f�{S�9{�*���<vjpb�Tj���)Z�q�<e�L&H�!����!�u���y~ j�Dw���(��j@�m#4@Q5Iy�-�޺���_��@��  �u�������V�r,G&�*"9����iJ�W���3�&�m�T�Ӻ4w<wx�O�@�9�X
,�M��I�+U���NΩc��<��N�D�����"��yk[�qT���9��VLץ`�n�cڰ�^q���/IY`V�b��5A>���s�
��a�!ʾ��~|�X�"�����K7u� ӌ��� ^Ԫ�}$o[�����]Q*���ȑX������C�c��'>�J$�tB(�s�;*5��{�J��T��.6@Fת��9Z���ޱ��-M���u�p�ÉbqO))�c��յ��k�,=����r�vf �8�k�m%�?L5����7�g-W��+o/�̻�q��M(�S�m.~�?'Y:3��w�w/[~��xٿj,it(�G9�w��P��ab�='���R6��$]����t�o�/Yь`�UT�j��O�\�Td��`��c�{���X��M�5�����ӫ��(/��EJ�f�a:2�$N�5b~�~��b��}լ`��F��3Z9��yp��G��x$�{�(��B�؜�쿊uݼ�*-��Ryj�h�����Ȱw�\at'�ѹ\�H�օ�`���+,������m��~ro���)��
ͣQ�d�Q��Q�<O)w����s�&Tk�X\$����r��ɘR�)�U�[Jp�|�X�����N�O�P�
%|�1����砘1O���?
it������\?*����:\0�}��/c��ߖBN���n;)Y�_:�\�y�l�j�H� vZ�	"Pp��� �̈ԩd��M�r�Q�#�>bT���%y�֪����Sk;�C'�^��o�#໧o���o�;��i�Y�G�2�-�C�Ȯ���|���@������ �7�@��熞_�K0�U�Rr�`DWS�}��O���{���^A�F�ZB��qf���w��޼��a���A"\8k_���RpAIu�[/d�N�v}\Ha��� w4���>���2�}�m���;M�������N�����Ŕ�b|�$�E�T����Z*�H7����*M}������_6���~ݍ�yw\�Oˡ6 .h�d���/��� �8Ls^=;�_J
a�e�u���7�:Ē�Ѷu��y��r�� J$���7�n��qb3*�����э��I����
��a�x6�&��J�KII�`�ˬ�pp|��h�:4�!7����Nq,�D�(�oS0����$��d2 �2u8\͉�਌�*_�Rm��BR6Ǎ��7ɢ���m�(̈́�{����F�q�n��'�����s��b��8��]����S׬/��#���f�ҫ=�.>��|�U����_���-y��4�_}��S��f,��[G	8����o ��o/�^���W�:�y����z,m���r
t�w�o���o��g0z�@���_��'�L� ��lm�Һ8W�,�����P��5:��O�����淦m��/M�os��o�<�����"z��sK?,)�De���n�g�WTfe�`I��Y�\�G>��C}^�w��}݋z0ξS��F��-^0]��]9�"���2�G��5]"_h���&{W)�gsĦ��������#P(8�t��-O����4�9� ����p��硁�T��܇����}ļv����8��R�C9^Yw+n�e����{�bO���r��V�������~�7�(ϟ�cw�S�ǻuN�{��X����E����p[��9��Q���u��Cej�:�������o�Z	��V`�R�|H�%̛uCm��zck�Ɗ�x8�a73F��m��5�լi�~n���ݖV�ե�~|�A��`��j���^��M_�m`����Y�h����-�q�f��.���D��ONyB6��������!���ys,'v����bZ���w�E�����-r~©V�4�m-�Yl4�r��S#�i"�`�^�0�A	YI�a�0RA#O�<�s���\5LX�' g,@#Y��Sʿ���ȼ�������4�(*�e�ڥڽEj
w�Jc˳wA	��ؤ���	+k�~?�9�G���,�6j ���Ԏ�� Z�D��(G��w�#��p`3��:*�p��`�:��D�d�%���'T��[i�J牅a{?M�6��W�b	��7K�*5$�ٺɪ����x��SF��`� ����|2%\7�@�c���ߕ�X\��X������B�j|L���l�{y�d�ф�uGr�Ox&F���5*���d����K
�e��;�͏��~i�\�4\�ɼ����V|����{��e<�Ɣ�ȌS�)�-�rf����o��Oo�s�h�sS��k[(�}u��e?��ؽ�t�G&����Röf�����9ǒ���k�;��V��~��;�l~�K��1u��ː����-]�\����g��;_{�{���Nt(;Є�o�$�At>W�c�+*�X���F�9��o˟�d��p�����bw[蛨ki�����Q�+�����@?�BT���a�g�܏�4�o0���YDƍ����Z����O9u�2Yo��x=o��N|���t�d{� �b�
��;Ӈb��ғ~}g�)�]�߈�/2�Z~��)k������]�éD��sk�Nǐ���11���&W����kZ��_��?o5P��VN������c����UpT'����PYl����� ��6:�3ٸd�D�����ϡ�gS'�H��:�����ꔏ�[Y^.����Xإ��V❿?p����
���Ȭ�Tw��;M��z�l�v-U���0���~m�m��W�!��R�ﻗ˅�B%鸛���=����呾|�Jۇ=����ӝ��s�T�)r�y{}� vB~�B�+�l�MX>�6Z 9�+�/�:p�����0oK��%_�<��İ��hi+q�Y�<|s�Me����U`s��s�n�R��*��i?�� �t�����S'e��Q_��	�ɀrh���5�Q&ͺ\$D��� �(���12��~�n!�*�rIxp��P^\�@L�QD�x������������R X����&�
9�H[j �@yQ��s��%��S��g�ok�p�Jt%QJ^������5G�����Wqj�E�4d�M,��T�L9l�b#i]��{�O5s5Pǁ�����}�*7꠩W&�����-^r���������9���|��vEn��흘1HD�3��3W*ly�0��X�T[���c�����7Q�ƮW0,�7�ϡ�5�ǪjEY��!f�m�VS��FC�w#Z��o
�)����{��x�|=^{1fP��{��Q
�p�q�בG�T��ֻU�
Ed�+�f6�����{DA��mI�rA�_~�g*�>�c�k3�d)�c~���ɒ�q[�����)I���N|]����ZD��p����]�9�#�P�b���3`����������3�����{A�~����+G�.�����^m�'��)R�Ӣ %����ʇ�&#�e�[��J����T�e��QY��B�qzW��f�`���w�JI�����sc^���k���v�)����9��Σ�}'��d�g��H�����1�1�k[�[�T}��(X5k���'����J�<d�G�vͦS�Gfy�_���� ��77Ι9O��"OA*dl�H�:���%㘩��{��S^3�忤��xn^��2�ʹ@y�#Ʒ9�\�S����_<�Q,~O[;��MNй�M��Q%�Z�i�s���x,��ߟam������D�Y�W[W:�|g�e����md.���s:��y��R�6st����Zv��/�3�AR8c��W�2�C:�OplWic�җ�{���#�w;��w��T��& x ��f O��a3ȡi\�^n ʚ��}z=�×GZm74�Bp�J�m*�v�����d���݉�)�b��S����Bh q/n�$�8-�.��:8c��x<�K��K�F�*[F/�+�e4�|�ޙx�$����RY1�#��S���V�I�u�Ӌ����_�q�p��s���N��v>]�N�[P����v��lyP�hL�t:Q}�"4�{: �f�JM6�¨�,��$jAȟs�J�H$UB��Ĝ����K��F�$)7�Ҍ�T��f��}�JZ[���R�쨢ȥtǲ��n��?� ���!#5s5��6��@V)��,��HY��!�<?`�R��>7�$ѧ�$۞Q�8:@`ݑ�D���`p-� ��G,2H�cK��kԄP&�Ż�l�鹪�DIgb�c��Ue�Lt��熃B�G� [���;}G��aնƐ��p�� J\�S�41�e�Ҳ��4�!�oU��x�t���Dc�M˲Ja"�M������Y$V��j�Z�4&�F3C
�Z�P9��-�S�~�X���FLL����fdT�9�φqt�,S����u5�31J��{6��x���ɏ�����U���x�����8�hy��:���o~++pb�_I֛��{&]uY9��(V���E���W.�e�Ę��R;��{���:!GZFߚ���7�[�h�)ˮ��A���������
� T�4e��S����-���r�e�G*z�vsjg4H�֞�w��昳:*�	d%r��}�-�c+SB�#����c�X����O��9ov8e��0�g�������~��a"�g�⮅<-򑌿�+�U��S�0�#�+���	���I���E�Z\o�lm(�0���q�������x��/���w���i7Ep[�� ����V�szy6�l�^r�1�!�����&��B)�m]VS�����Q
���1���2{�IN�a��p}��Y˾����WϢ{�U��s��q�1hs���Qۻ�x��/�8�+��}�>�,�\����)�WG�c�7El~��>�S:��dD�I�j��D�CT+����OS���J*�}��cr��F���ŭ�MnT Y�X ���ŉ-��ø���_�?��7���}�����Z9v83!�M�c��wp��ο\�<��������;&Mnr��TE��d�N�/ޕܴy����S��;���{��`���VJ���S�z;�;
��V�5u�H�Y+Zp��=:!�]5\�(�!/�{������|>��/�Wp�X�0P��U��vC��v;�6Zm*q7�u����^��}�gzam6�ǎ��Z�C���ãT#�:x{;�s��(aRA����&i��0C�[��������63��Iܮ��6��V���ra����������,�K�И��L�
[M�~D$ .�?\o�E/h���@���ta��A.y�zqʹ �,�4n�݆���g�<ʛp`��r��UK��y�*����3)�<�|��������B!Y �ܐ�s"�@<_��S[��W��ċ�f�HN�UHu]U�\ ��E�Ԋm��~̆aA*-�L��Ֆ*y��k[|�N6Q(��N�+xIs�k����<���f���-T[A+W���#C�9\2L��;���$"���/�j��AIV ~��D{' 42JiFd"5���p����̤��Ufu���}�Ώ�������E�/cm$�+ѶE�F��9��{U�my�����y�p{-C� �>bF"b����-*���x�M]ϟ�2�a�VRs���$zG�B�/����ѽü���݋p�{�2��n{6m��>/J�^�XѮ���}+�nI5 7�J����;���j􏂫�?
`�5�y���׏R�UD7Ϛʝ�!W�4��x�D��K�"K#�2؞��qkr�g+�120��E���C�"��^����Q�N��.�-&�$��
T7ųA9��Ғ�M��J{x�����t�*��}qj0헩�X��B�`^����ڳ��i�1�`u\���?gj)��=�!U�p���ʜRcV�!�P<3C%GVR�6*5�����Ę����Jd�U��8��=u�c��,*8��M%[�}�e����y{�?-"��I��0��r�όRb:˩B��{x����cL�i,u� R�z	��Ο��n�� �v���V��)`rm�Q��p^����#QM���4��D�ϛB�F�Z�j"�zx7����)0y\ק�!.�L� ���Z�3̉YLߩ��N��|��r�O������
t�73%�îU��F��q-���0���	���>�qp�m�G]�dQ�l��u�"&ݽǬRA��n�q�@��w����U�~+2(XΧ�d��~�cV�&ꚁD�p��]�d�Vl?�玞������?~|���Iߺ${�>�Nu>WcY�o���v|d�~1w�)�&P�3]���n_��vx��W�m�{ݲ��私�$H�N�T��x,f\�H��~eSq�#O�qtt�m�����<�9�f��B��H�CW��Z�r�pBl��ӑ.'������v��G\w�ᇂM@^���>��-�ͦěr2Uv�o#��=1��tDm7"�����m��x����s��qS���>�2�y�J{Bֆ���!�ŭm��D� �j�r�~xxD_?�Cz����vl��t�z:�~y~~�a<�|cS% �� J�~}L���זh���4o.?j�
� �q�(��9���� u]o6d)�ә|��v�<-.3<YR��6�#�#�
���v<�"W��R����/�C�Y�� �7^1SN��5jԜ�F�db>b.!er���
�T����/j�w2�І�����፮1��f��zIuj[IA<�
)�;Qve>p�a5Q��;��t>�>=W�&n��K����*5V*M������~(GDF��P'r�^8�HI��%�)ԑjʠ3�A����Q"�C�m���2=��>�H2."ۯ��j�]�̜LVu�"�DQ��8I+E�����y�5s0<�Fr:C\y���d��
4�ΪF�q�\ΗD�.F�Ӥ_�~�������O"7
�膢���z�yϔ3���;ѝ�W%l��?sv5��4yV�闏����t�9���T��)��'���H�Y�|����T��dc` ,�Z��L*޽����RQ��4�eE�\y���>)���O��Y!�|�R�d��W�� ˍA��Q�TBϣVH�([��9�g�E�<�'��h��7� L�ח���垛ϩ������u8p���c�v!�4-b��!=��ŨrNS��h��;9�S8���\Yv�˳�S/w��9
�*l��Cn��I���c\�+G!�G(�W��m�ڕo`)��Zv1�J��*Ģu����9�B�+��vp�Zg�Q�+�cBt�R���#m�� z�'��N���F�s�#R,:;#)#䜇W_��:vylM6�q	�/-\�?,"3J���1��?I�kh���t����m��V)_�@�` ��=��2�IF�P�0���Kz���D5yW�+���}� A�򂨌 �ɐ;C?wx��J�>�p}��Wg���t��l���]2�=�\q�l�*XI�5i�o�=���ӷ���Y�V^���):MSN�/U�8}�O�N�]��	{c����O����������e��Q��������Eiڜ���"v�:�?�� �(^޷�g��^�_��鉣p��������cKcWQ?JId�Q� �ʃ��m��	��C�
D&\�8�
+��AH�~���+�ސh���.LFꂔQ�� +F�Ö.��b���+��gc�kC��0�c�rOT�0ܼ���Md*>�MM"v6� �ao�h�DK��#z�1$�N�*(�n�J{y�b����TT�PRV�D���Ö�<�i��3�f�ְ�^#vN'T`;�$g\�畢�J�Cm�3�w��ڨ����H��[�����"T�]Swb��Z����_��V�����| ���Ǖ*]������}��+��%m �������s:5<_L��J}%J79g��eɗ���F�rP�������1Њ���������'k!�Q������ۋ��1 �W��!���(&%/<v^`����jY��"Ɛq��vD��1y���Q5�>�^1X�H-�1�B����� s��L�m��1����S��7��������������~:f�ΠkĔ���pb��	$�����ݰi4��_MNw���v�UӃ�_�s�
��K���㵃�g����V}�PJώ�':�}�t.����{��Ǐ�wλ~Ol�R@.($U'���dZ��
X���vn�W�h���ny�d
6&�m�Y��O:��3��w�$����;�.RϬ���ύ"�n���vf����j����\l!�N#i�Ʊ��@�|�+��5�5+�Dn��'��5e�@N�N���� ��>�sNy�Җ_�r�q�f�{��)�N5`�TK��|���:�<�kU��`#⚿�;o��ƫh0Z�TO�ٹ��$����V1��<d�"mT�)vT��5��856Ǩ.�@��4YTj	�R��c��:�5t�e�o?��<dg(�b���U�*"�JA�ge�0��ĩ���^U���cA��'��({����J�|�iE@b�9d�H恲��S�RP�ZW������y�y	�P���G.7f�������\�G��6㮎��}�_{̥��~�J���G>3��|�b_Q}k�7O�y�.�QU�N�O�B�Ɇ�	E�]A�>��~��=���4ry���;�W�:�W���!ך���sۘ,}:Aѯ��ɖM���(����T`�*�u�C�^�z�h�$3·#=����tO�#�����YKf�f���Wζa�W���樝��"Ȍ��ܽ$�����Ĵ+�Zd����
�;9�O"dC��F�c�	yL&�%M��̋��/ݙ������vYz-�?a���]N��Q ��ܑ��$���)ys��
���&��|�K�����9�bm6L��٬�P�W���D�
��YD��	<L��P� ��N��g+%͵hIuaRZ:�	@�Bŭa�s��,&�\ɓ14��(kA#�lM8��rhň �g��'�eд�V��cvK�%h�q��S'ݿ��a���!Dפ�F_Yx4ȫ�«���sZh�4�"{�$�Ј��S@���+�V�x�j��i�5�s5��A(�ذ�J#OL�8_:�t>6��Nx�������?���M�<@��e%�=[�[��U��ަ~>���֑�V�y.�Z��d!��y9s�x�e��P n�ڴy�Q�)�۩B!FYH=�<u�IK���~��]�W��/!��\y��4f�Kk(m`�3@�� y�^C��*��#y��.?����mJo��UqFjU+ !���Z����c~#����Q�������%ћ3,��a��h���i�e�s#e1'1��^��K��d2�T���f?����V��@^y�*�������v7J�n$�R�/��Z� �=��
i��:ߢ�Eb�D�&�n��@r��5���{�q!�=�R �| ���8���9:�v�
ƍ�˟d�dr1̯\�ˬ�戝P|��ם	���_��)�v�|��Ɨҳ���'����.��y�����z��Q���8��2��֣w�P\�h|i>.fp���5F���I�^�$�-���Fy>Y{���AU0�A�Yi���Nv4�IȂ^�~�Q��6B����3��}�?�i�E�:�~6dt�7b�$�����.��ժ����U�Yoc��ʚ_��!-8��r��W��_����{r����������#Y4s`�9N�8�K�9U	����,����m�b%�l�b�р�����џ��)��A�H����l�ǵ��Z�5��6��F#�jI�5'��l��� ���@��J#�i?�雁��΀�ц�&[G�pJ���E�R]�+�=r$r�kfDG����������R=(�9A!��W���X:n��FE7���SFr`(���S������ș���"A��G��V���^� ����]��/�b�8v0��1'k��l��kLx���e����ؾ�����y;s�[�<w�ݱXT�}��|ݙ7��ns!m��U��4st����;�2b"���n�t?n8�����vL�B#���Ӈ�߷J���Ι�A�O���噳)����ܥm�b������xa'��п1��C��_h����Meֈ��S"v:�ex���>���@�&Cz��I9���ΕN�
*�Ũ��\헕nǁ�h�״�}���c2���(�&C���o��R�KNǧ��b���Ц�`�qe�T�)o����1�y�gU�6B�M��=���|>$e��/��,<1 '���F��	<6�pfAA� �q���=1�k�+C����(�~Zc`���O�h��j��$bBCG����]��tI�@U3|�\|\��~hy�̊���-/F�P݃s)e*�.ۤ><l��a�)S�|➈�@*��4�4�C�g@;��E"= s��$�A/�ՔD@V��)A�Ҵ�Z�}��"Տ`�K�#)s:��Jc�s���m��7ɉ̼,9����	ω�>)�;(�-��_p���
B��V^�Dr
TQ�½:4vF�����N��ԶkzM�P�����!J"L$5t	���� ���/]�s�ޖ�mЪoC���~���I�����r8���ҕ��qT�qP�A�#J��\V���|*IvjR� :��������x1Jڜ:�%bl�;��ہ�5}Ε�:�>d~4���vi�2�f��o�_�fx�F��ڈ���S�_нr4/�U�P0Z��R�o��7�]�n�aN[J����!��|�0ٻy�e���"����i�E�ˊ:��T�ۙ���� ���s��D��!M����;i7��Z?N�f�w��ܺw��\�rPǽ1ֆۚ�TΊ+K����L)�����B��%ō��g*_�6At�vZ��+��K���4C +��$�?u�8�����m�O/j4�� ��>���F���_��#]A�[��h�q���jt[����^��䈝�T�dPG�0Bnt=��������H��� L��W�aB���m��z�@�/'�$IqU�W}<�Z�S�n�Y�/|�#%z6^��^�C{W��Á�^����Ռ����U�G��\9�lV�=���^U�ɵ�WIY����N�/^ �{.�Ј3g��Ⱦm��qHD�8����_�6hZ�<W(�}yn���rh�;^�;�i��)+\-��Z"�{#���Ry�O�uQۿD/�C����xaٸ���;�v�W%4c\g�Ue�M�s_�
�����
��^�g"��̸����{qv�^T���}Ie}�r$_Ǌ�L"W|/�d��f� ���k�tIs�,o���ȇQ�Ri^�=F�*��F�n�H�����}7�}�S��"��S,�&��5^�E��L��yy�%�{�}�x�i���;_Z���/m؇ߟ�n�[s�ҋ���{щ7�-��TUئ����׿�ׯ�h�adڜ��~fG��ź���5��:<��ҵ�T�dO���$�|�dc%D�l�;Z%�y~}a;	{y͕�+O���6��UĎO�9�StB��p�hD�K�� �lC7�II���B�?�����6���ZT�:�9B#�
����V�D����c�=��\3��Â���#(���!�:��&��5�<07ROH=5�d �/,�I���  |Lދ4���` �7���X��B�~�|)n�l:f���x9��V]����s�k����tDܮ������}((��Y�:�M�dA\��DHVb:+��!p�������,V�6�I����Iǣ�h3Fw���\8�.H��"��%�"��O�E��cj�(��	K.��J�戓GU�[A/���֥�n�����!Ph��(����%�	)�jU��t" lu۸�Ɣ!wV�/')�����f�|δ؄v���1
7vLz�m-�ՠ|50P�	{x(���>H�Y�2��5P���A��FB�1�����"�ń��e�.�I���+g�Y��S��>l�1���߿2��i�i~2> 1��)a�~.R�7=m�k�08kڢ�@��A�X�w<Ww�{;T���-m?�!�����|_�,>��Y���BBьc���#@�n�q�&&���ъd,t̫�y��c2����/�D����I�S�D�S�r$H�%��;�+Wټ��e��F_�)�Oo�aޗ��ߧ�°��ғ�#	�y������Ǐ>Ҡ9dFLTٞ� ��~��^�^4&3|'�1��`�g�EW��A�?	�s�էـ�7���>�����wk\{Ls��`�t.6a��h��F�y,��l����ȹ��2'D��!g6ۖ���!M�A�u����iDT+����JM-��ҥ�Ga�Og���}�r�Ǿ�r�Uh�� ���?'9sR�(�l�G*}N#�t�gs��"S�%
i�e ������d�W�W ��+�t�+�6>D�H1N�>�l�!ȆCԾ�����(��xm��ΊȞv<��w+�`z
�9)Q�R&w�ƫ�h]�`��E  �H�|��v���$�\�T�<��,�P��u��Yw�:B������XI�2@=8Q̙���AR�g��s ׻l}K@��X�^�t����=�h�����BV���9k��\��:������˄	��U]8��srT����e��͞��}K6L7S�#;���G���-�$܈Z���`�~�B���7Q�=M�]�Jc� p���,�{%Eo���#����O���+�38w�=��Eb��Q�P,t0Q����k]!G��$).Pv���<ω�����~�(?��U���͐&�����W��Ӌ�\͍_���}�!�ѹ�Q�e�����%Em]����m���v�=�^v����߾$��砇����pP|���m}-г9j�=��� �qT܀����2�H}��ʡ�����s����˱̱�fo��<%���@``'�k@���7��������a��8Rc��#��N"8$}B�mD�/xf&�ƒ��I}��a�%�ة5��<C~y{���Wz{~`��i��ܳ0e�=�N�ѫEH��&}���c������,A	`�G�!�����Pd�y���U�
��«v�~��)BdK:��ZIV�8:�&�I=���c�ן�n���%�0)�I۫��,N������ŐJ���9��2XD����i���;_�T�J�Y%���W͢um"\:XD�Vn`�yX4Mi�܋
|Mj�>�J�t�i�F� i	Z;�uU��G�D���#����v}p/���_�9�6���v�}=j��G�Q�LQ�� ���˞��?8j�*!��nHr�vD�(�ӯz�c6]wJ�D�3 �A" ��jA���=/5^�:���Y
�A�D�ӊ�����h:e��$�|�:���h�"7q/ �h'�f��2p>�
�h�����4w��T�̶_.����MY�����ri��ծ�J��SdPmKc�g��Z+�♕9�f�v5��s��霷t���/��:I���]Qx.&`������T��)�g�!{���5TbSH�',��=~�6�'�l��s�z�q��WH˰y9uG�:��\y��v��[�)۾�;y����Z! ��գ�(�lc\hE��M[�~C��tm���6�w���D�X�#�y�{�C���K])��y��VT�U{j�J�K��>��h�Z��"6�#�t��<PB�~^�y��h�JR?�5G}�j�#�A� ��eU�����r� ���k�I�ݶ�Ӈ��߾��7�HR�@Ȑ��c��l'�P�,"d��޴\�-Z�Fu�U�H�T��V]������;�/�D>�(�M�^����#E�۪l�Z����g_,%*���;�4'�h$2
�Vr$�U�GM�S�r��0C��i=�$Rg�kّ	}���xh�z[C0���
�l\Oǃ��W`G�<H7�CD)�9ޓVj���gBn3�2�����8j�N�U�]��Y��<�[
��;3���=jLN��]�Z����z�W�c�Y����^1*x��9�!�K��"!Wg00zL���QƑ��Zx���&��V�Zꏸp��,m����_�b��Y[􎌏��E��;�N�e���@��}:��s�l�)dnn��k���z)����±����)�K�8R�I���;�)��(渨��k{��v�;�_��(u�RR�^%�$(�׋�sD~�6��/k���5���^5�}t-B�l�#'���_2g�:�gc_E�d- ���4,��!�s���������PR��d�T^���؋l���,,�$�,i���ʱ1H�.���c��v�u���<<��Ю��� �pҍHҊh�U&��C,���T�K�4̯sK��"$��Q��� (80~Q��U�u^_t8�Q����eE@�rL��B�¨�p���[.n��f!Zԉ�a�W>�N}7������gЪH3�WSx�p� m�PA0RO��c�.����]�'�ORE(*� 6aN/j��x��͛�wR���v~�x���ޞ�2�d�e~��b%[z͂����"ʜE~H(�xl�l=OJ�x�j�dT6�hY�*hE�A���R$�0g���qԏ�D�p�j*˒ba��,{�����íJ�x�P>Qa/\E߇r�[f%i	P�DQ�"fA�3Z�c����;O�V����܌��S��:������SNq0Y	Sa�a֭��o(4�<���VR�#u��""�J���7��k%<t�J/&�+M���i|��&�:u.�*�`FV&���4��jܑ(����J��[����F��;-=!� "�@�h�T� T
�:&L9Pũȅ_<j�D;�6�х�U��IZ~��S��k%�5��P�Y Ew��_�`P��4.�
�:L���R�b���?��؏4�j�����٨�l�^�4��\�˰@��xd�V�!��x��o��������?W2gʿ�#�ۚr��54��'w|L��X\�l`�,NZ{So+@����傖��@/��|�f�ۿX�ŝ
c��Q*�v����F���R�fk���x��D�f���fr�Ԁ���˪x�aQ���Mk���MWZ�e@瑣u�Z0�Ʒۏ��ȗ�����W�CM����SD 1�K���R3���?�fi�U9,�3F���Y�~�~�7�y���sJ�00��iMǴ/����k��1A���u2Gӥ(�~���ʙ��!bR ��3nD��o�"�����~y1�$��pg��q��U"G?�KC���ۭ��D*�c�xn\���9}�i�)��r������k�8>b1/M��9e��8	��!��1� ��D���q[��|5-������������q���: .N-v������6G����)������L��BN�he-Xt�+����IGv42�8�"�� "ð {�s;��,g婦k	شR��5���ə���FDA��4\�d{	 H�5�9�dε���ZdA��Z*�y��8��t���.ٮ�:�}p&ߣ�\�#����E�4�&��'���b�x��#F9�I{'<Z�m��t��&�c�4KST���tL���@
��\/(t�) 8��ȋ�����r�i?Oe��ͫ?>vLTM�,���y�w��,�|q���tO��s�ڦR7��<�����Z�i��b?|H�ַ�;���.�ot>��~�/���`��' ^�=%f�r�+���A4�V���/�k���P
*YZ� ��mat����U�H2@�7}��p�3�U���`� �	����������7�����:�e�#��iQ=�M�JpH&�,��
g�*y�+�~~n|���\2v�L7׬P� in�	#ަ��'�����F���6�b�(���P1ɫĤJ6-�R[��f�a�~���E\��WN�2ZCB�\`o��%W��<���M!���|�`�!�/]�iS��&�m,jg���9]��MM<%���iF۸+UE�X�eLd�⚕��q��'�U곁sο�����wz��D�O�"�6�Zp��_�pD�#�3��wߟ��ȩ��'��u���/G!�r'�T�j"͋
Sq/�	 ;n*v�����n�Fq��@�+J��D`�ޕ
r3`z:�7"���;�M"Z	sh.<m�]ǂ�B:Q�ˏ����Z�Z��+�˥�#oL\���%�/�2�LB�{�5tJ}��<(�؅g�5̦�=��ۉsO{VJ%�7)��:����Q=ؘ�D;]�U��T�qE�����c^�=�hn��C��i��h0"]|������+���sʤD���5�����wDJ�Qͽ5�y>2�w��W�N4@9F�l���1��S�>wx���A+�E!���3�4^�5���0Qn�����*F�H�`9M��+֛�D� �e���P��zI��X�Z���b!��rX� �Q}�R|�֕��E�����U�2b�2H������_���wM�X��6��T*QW�2��2U����aA�����Y:�h�J�L��(���1�x�!�7�형�X<
_2W��!1e��ϔ�;��=�hQs3�//;!����e?�`u���q�6�a檁�a���t��Lj��x�bZʼ�s��J"7o�brs���l�y��j�������T5�&7 ����i���	�m�x`�,�/=��|�SɌ�_�&��bPڣE9%'�E84,J��r{T,'N�;�� IIyu0 �N��r�<2G�%GB�{lm`�l-�h�����*8T�iV��9���}��h\?���G/��w ��� v�d��yW�8#����̉�wZD��8	Dv���"�@xx�	��v̀�D#��8��o�t8D���|�78W8cc�S��(��:U�/<����'�#̍�v]Î ��� � ��F�6���_�����yZ	�����+#��PW.�0�t��������r4\p������4A
Y)��������ڈ��?��C��3��.5��P�1�����l��
��̋Yv*����8�ϲ#d#�T+�.�]
E����/n�d�%�I�C�����F�4^�,�������Z���^9p+'3(��+"��2�n��. X́�	[;��`������~L�#�+���#Dy1��6<'�~��� ��p�Fzz�x��g��+���u:YY���{Q�C5����C)=Kt;�Yث6\eh�ث���CxYՙ'Т���C=%��$�Q4��M�4IdUX���&t�*��"�n����P%�e��kW��Ӳ̘W�{��U\��;%�OY��:>rO*�麄}6A�>p��un\w֭ea!�YՒv�{C>�C��}�n�3hev�>'}60��v*2n.gd1Ǹ���P`M��d��lY�27* ��:��rH�i蒽�a�>_��#��&m9=Tțk�����?3�)�&2yr�5�����F �QY�E����W���o����_��#	�'�3	�K2�`�u]ͯ�ߧ�h-uޫ|�c�9��Ι�2�=���35<�C��d�XxhA��w`��	���- �1�b�p���$��h�s����OU`$�Q��a4YM1�O�3+r�d �s+-79����Q§�52�Q�G:V��VD� D����&�,���:}i�0�$��E%m�p��B��1?=�П��!�n�oL��*yՙ��r� ���R�`A�ҹ��<P��X�����)�)����ۉ=.2��?����S��8���@�*��-�&	[AQ�t�j:d��H��5�TĚ�ZS��+x�l��!%��L ��I��`pG�ohˏ�g�.�ꯁ"����_���E�.Zm��&mj��id�N����KKY[1%;m#UF��Vc��tf Ӏ��=�����+�+q�tд��� ��z���u�.E�Z��X��N�{d�	�-|F��u��Ui��7㾓px�8�	��OJ�����mE��N�fRz�\���;�K�d�q��c%���i�n�()[�`黳Q(ͥ��(ا��M���ܦܠ�����I6C�%���Gke���0xx@�	!��e�̀���Ú.i>� �.{7.��VLZ�^�F -���Q����94����g�=yF��{���H}��=Lչс�˗?�䑣*f�m�w�p����Y�K��{I��E����ca�N(���������[败�n߰���6&yR߻sP`�R�4=����s��������3�s�(�y�"bg�M��;�*e����r	5�C�m�d���-��^vY�J�/J�\̛��Um	ΊA�\-��V�XY�!M��#��m�0��5n^sWu�JHO��HZ﨩�G�C�Ȕq�@-*��ua?��P��Kf�Rg%sz���Qǎ8�/l��X�"	s���Cƅ0��7\E���Z�7��=��P���c����G	�Rs8���->!�G���)A��_K�,G�������}�ml����^�(�¢<,��V[���Ұ�y�D���.i� �i��E7�-*�""+ʆ��1�X1W��&h3@B��5�g�\,c��^q��y��(Q�1(�M�`�8�$Z�ܥEJ8� FS�gKc|"l�_1H�)WzTG�rE�x||L�}K;+.`�:��c���D֣ϡW��9�z^Vm"\HV��l+�`�21��RnL��y���a�D8����2��ѵe�X�3%��R�4��K���SW�' #Dqh9�{�S����.�=I��u���l=��-AtN���1��I�HA���������hD|Ui#G�d�o����rcd��B�!�	WO�펬O;RQ�����)�w!C!,g&��?���},�xF��Ё��4T���Cq�����Ͻݓ�
����)V%��Q��y��+���̣�o�ǜu�K ��H��4�K�s��>��pv`�D��OO�����pw2߰fq`x,Q1�l�	�V8&;a�?���@Gn��i��ZN��u�Z|h����D�P9��R�Y_� ]�l&q]���+������Ƅp���?���@���O��A�a�JF���e�������YC>sD�ԑ���7�(!N�T��V}�����n��JI|1��=�P�$�������0kX�AD<CS�#3���
��Α�Yk�/�8J�TU Ch�Ի�v#�r��4Nб��� �����ʈ�:�a�����Fh�D� y�p:U��]�.�U<�2YRD��V�Ψ��<KY��Ə�P� � �녎�� �"l��Q��NM�-��W<%�2D� ��M(���!m�6����"��=��G��
��J@>���h�A�B���Ȅ���W�'��B&��&�^a޽���+�H���ĒR�#�:z��p�,TW���H_��Ư�7z{;r?p?�D�@����?~�]�����%kj6G�y���g�[�A��d�0Ob���D�55/�~'�Q�jR��6i��뫆n���"?^��LPD�}���G
҇\�K�/�����Y�q6TԈ�=ǁ
U��*4���QM���U8���:u_.0�Z�/y&(��[Li\G-u/������'@�xʘ������q20e��7!kt�,���B�#7LA	�8�U)�ǼCz�L�v���?)���
�N,�U��ߐ�q�c1�����ڦ@�p��i�)va���ø�,����2��oa�W�����L�~���y�WWP0*�o�	���;�Yn�f �Ҁ�\��F��k��ƹ�$J
�/"dex>I
"#���d�k���Ӯ{s��������-����7�"�srO-*��������u��uH8��O��4[��#��y��OI���mQ0$ۆ���`�����D	�@��¿Yq*ﯵȫs2F%:�d�dLV�y(�9�O����\hc��)� 2T����d�/u���c�t��)+�sw}T��I#\�yG/��=2a�Dt���b�I�o�e&=�8R��i|"WeN#�`C �)hD7����
��t��h[+�c��H��rCO�:M��g��2?T#�ɐ�%��Au���S�R=.���D�u%=���=�;��C��h��/F�h��Ze��"�D��+M�� ȿAg��4Du�Z�Qμ�C	�	���3�a�h\�@�.<�"�Z���J�]Y'�^,Z��1ލ��EycI��1�]P�֨6��u��m�'q�F:'��*��h�g`GS�%*qT*�Oj_"r���N�3��
B���-,�t.�0��Q��ͯ����vC�FY��G0xU�m���a��wn�ri�������C��k����4��L�f��MNRl{��2"�%�\�������_�?������%���^|������?���d� �@
j��`���6yb���W�oi��i��1���i&C��RY�Υ�������^�i%�G&O��n:�,��6w崓eCZ�~���4 �}=�џ��d�K2~�U�6b����I����6�P���c!I3��t>�=����H�A$�P����n$ch�/��ç�^�\�>�ߓ���-A�����s��)K
����h�b�D|CTR��=v�@RK�����!�\0t����I"Q\����C�I�H*ef�vF�*��_'5�%�]Rʐ[�>;$�s�=pt�Tf"��TJ�Vk9�Z+�� ������p�pU�x!��ap�5R����F�|���.�(d��!�co��d�Wڗk���F#iyZb�n��0'���s8^�f���g�F*{�!0d��{��EGo�3�J�y�%r�Ր�m�N�]�BV+)�b|�����#mЇ� e�GU���(����-��/P(�z�k`�>(� ���J"�%��*�ծ HzAÀ  G �FYv��H�{EՑ�i#~�9È�(� 5�V�o��T:��m�V�Г��l�a��V
�~``�h%b{߄'������s���ǩg��-�sTR땐��UI�
J\�J���p;���E�{�s�<b��B�[�r�{R����N�~ﹱ�ZQl�$G*7�~����T�@�=�����c�^���Û���q�[q��vz����v����n����>�>����d���Ȕk�&�E����w�[������P���7���6��K�>՛p�rv�h��w!���6��Z��4�ǿ�Og-3�S�����V�c[I	�HȑӌA&�>EM{^ĩ���_IC��?)�]�+U3��.���q'����t2	e��ƝT֊|�t%sDT�2˾�C�b�[����%e]<j8�裪:O�*��Z�s�
�jz����Y�)n�"lE6*��m�{I�*�y�;m�*RQmҨ�DA��1��~e�CY��%�Η3;��j6%ί���$x��>p2�h ��t�ݎ#`�C��D�����8��+�pp��^��H��عX�(S�����CL`�z���!u]�,s�Y���X�ԇ=�n��@#)A��Ϧ)˕V��4Xk��ِ����ƴ��FW�$�kXe0{�n�F��G�R�<���	ΟF#��g��)vQu�1Z*Q�H���y����Q�����z��1LMx�c�}���l��^���C__��޲�%J3"4+`�i�.�b�j��J}����E�J�����:T�S�Q��ҟ��`E:(H��΢x.�1=��A�$L�x�C��J�fY�������",� ��O|���b�I(��S�'4������ᗓ�[��cR_����i�N�-۝����'G[�����lOpN�B�~挊�u붑��Qm]Q�*��:����$"�@O����g�> J��q�V�Zb�z=Mdi͵��M�"B�*�I^�yM[���ˆ,�j͑�vŠ����� ���tq�/�p��>m��si��T�DjJ�a�i<2����]���$�B�|�����G��z#1ߌ8����LB�C��r%p��zB�dY�%�T{Z�iM'��%�#��+���9�9�L�a��~/m�B���[U4_)b8��j=����Ip9�pЈ��D�tL>�rcC���G�w�Ց� �Pɞ����o@�����a��x΄D�"�	�B�8b�<}C��D� ��k4��PY)𦃱�e��&��{6pIqzabb�������~�X���� ���qD{W �^�]��Qr�ٛ$����{SB+���M�޽���^����x��G�e}a��X��c]�9���1T-14"�P٫��?�~�p��FATw{;�R�Ԯ��z���xJp���#���?�t��M�\U��5�����wV-��i~g%K�Q��1�X���E�l��oj��1"��XO9�R�P����)eO/O���������zݷ��=s�։�w������+�>#吉9L3&E���Q�K�3�:
����XES-��]�:9�%��z�py�W������Te�a�P�;D)���������ؽ��v�ȭ����Lc���F�V5^��?��ש_��|8
@�bQ�*�N�C�a����|�I�\�%Y!Y�V�}n).����}��L���SnE��F��OO����V�37���|��'.U��X aڷa�;e�UV�����YD����.�I���md����{�{�]�6����8��\n����!D�Ty� +@����6�+I�$Z�5����������6pٽ�<N�s�  ;�*��5%���a�dDU�����ǡ�Yu�*�,j�c鄁���P�@%�K��a�
�LÑ�£1��I��N�� �9��0��}c���0���!N��}�R����~���7z~~f��P%���a��<G�0@��ތh�F�YT+��`IQ��Ϋ6�k�jtL�T�B����S%
W�9�8�K���
�0�`�\��g���4%^tíV��=�DQH�F+�ˡ�a���ypɩw����(��2Q_LR�t�m�zK�t����m�u.��|��}.�����Ƀ+��5�zy�ރ��0��u�F���]Q�O:W���\;�贽��3��Z�tT�.9��q����i �v�$ߣ��h��GRV�C1�X��T�����m"sR5MZ��1�*�>���@�n�ٮd����3,��a4�d�0�6�ƸG%ϕ8�$���q�j�^�T�FunI7��_�eHlg0O��N2.���(�<��S�m��;���d�;o
tc���lԕΰ�
K׽��b/�yB,NT���$k���Ý��P��E4���% ����\��Ȁf�����Æ sI�B��͎�;OI���!���A����}.(��=�I�e}`J���W:���	�"ϼ7�1G�e��2���	
/�>Id,�,�#����)�Xh��k�(e���4����9��U�gHKw�d!Ġ	��u��*�X<��|Ĳ�����sN~��:��*�n�O>(�'@F�B8̇B����v�i�u���"@����ߑ��^���' S��]��f�ҰXZ������%��El@ ���+��}�|�b��V���;�^�H�N�y�d�fZn<J�)߷�r�|N�P�H� 0�o(?�Mv�,�E�Ԝ�x��$���Eb@�a�eD��0"9�h���n%Ό�A�^͠$���"�yL�S{��^&&#T�Ec9ǹ��)ٛ2�|��jC�/$Z��y�w�r�4Bs����)c0��;�<�I}����ӅF[��ގ�����vU�ܖ�|�/�&l`��>s;� P�`A�| �)�uOJ'�E����^^�)~���2�1Zi弍���:�*�I(�U�^n����n������W�{cC Ԋ�x��o�r������pJ��7�3�yg�I�<���=��{/��,��d�A�	���5^E��o�d��3�<�=/���ݣ�����z�񚌋$p^O$�td� ���5]g���z����w��Js��4/�4����=�=�4��j+��l{���E�-Ejw�w�QD��?"PJYarq~�|6	��|��?s���ӊ�����rĥ�Z ������R�6_U�KN��}8��y7�ٺ�lG_υ)��7�˗�U|M�2g�4X%���ܩ�P�)��Z��D8�������X���SB^Vђ�+��#U�������p�FyJ,z�KGAb�fi>��P<��*��娩X��f� �^_p��F"-����lc����ш����v�ɠھ/ͳ�
.��ȑ8u�� ��Ȯ��I:qX\�#�VH�*X�:~���F�w���%\��r�ב	���"�ӕ�'��ra}2���
�����/�Q>C6ątֺ_�?�O���F;)��2A�88��eN'n+"KG��BFC&1��ĠR9r��	���5��y̩��Zq�<�U���~J�us�H*_	Ioج$�|���h@V�� ��~<�q[���~�ty-��d�(`�O݃Kq�Ԥc�����`��eH�{V�$�M�劣[~m�I'��T�Xe���@�U>g�d�n��b0�����K��s��b�DB���^9J�gz��ksnx���[�P�}�c{�����I�ڶR�ѻ;l1�r�� :Z�� ��dN=L�:�B�8M.����n,��X�s��LI��I���I�^��u�\]�ޟ	N����3`�'�?���wT�H��w-�?��n���V���;������)�U���z��׌Q�y:D���("����.@R�m��o�}��ޕF����
�=<�S��>}w(� �hD�c�kul�mZ�ăX�F4I�����&�3�RI0%��#�Ζ���+R�~p�mv���I�W����2F	w: qI�"��ϟ:�~��� �s�Ж�iIIY�P���~"�e�D�E[ffkN�}���e��D��	�ܾ�V�b��ͩ�|o�z���{~'��z�y�$�ǀ�`Aa;��h�#|�	�Q�0�Yq���Ӱbf�Q��t�j��:Zޔ�P�BN���j��R�teKs��lk�Pَ�wԬԠͫ��3���ēۂ����I�t-@C���(.Q`���$�����&�S�pQ&�4��H��g�?� 2�t\T�@��g\&�`F!��T��F-�>ᔚQ�� �*���A5�4�l����6���%��X�@.h�6ȗ�S;`�"�U"/Vԃ(*�(�=�o<�̳զ^s��*��Z9��Z@��Y�@��j5��$��5ϱ�db=�5��R]�s�C�,�T 
�4���c�"����1F�9<2pE��#��xv���EA�h��l
�D'�1��~����Oܗ�R��ii��?!frFxC����s����G�ңj�@Y;a'D���ZBI�N��/��z D��6E��3A>�s0W1V�4����re�t/D�P�WC�����6����K�|j�gu���*�q��dT�t"�Օ?����Nq�X4k���)o;?�N3���K�~Q|.��d��7π���>��(Q�'�punK荙�%@�;̜��UL�'��!7K�0SM��p�=S�*�T�!Q��`\y�.ͩ�1P�}�j�b� �+]���bz�//�,��8�VSd��q�u:������J:nƈ��$�y괼�EPsE�Q�VY�'�v�<�ޅ1k�>d�Tަ���GKSE̙4��A��ߙ�{2W����|��;*K�5�|�)c[��iYO�����?�������6`g�F�j�:?����-Gow+�9T �
7+q�dd�� ��r�5;C��� J�n%��D�_��_�aGD��5x���#�|-�\�;��)�t����fo����9��b#�V��3�����Jq�+�^\�������1�}���(��#���ռ& ���|���n2(��ʹ]1��1�/sH��A�>�
rVuc�u�7 �<^��p�` �~������g���Rz�����'�<����X�ZЅ��A�O����JZ��3	|T��\�=s�hn-��m�:��(����������|珚�=W���x��_�1���~�7��l�\�ޯ�Wo\����������/�:�ȱ�E��f��Q �VH��:�+�^��n��	Xi5��k6��"|��d�lA���tI���Z�-�0o���nQ��h��12�)�����>�^ЩӾ]G��L�<+�)�Run�.��2�I7{���/.��3!�v�X�����q��I��\�)���ة�D��Mb��P�Θ����s�ԕ��wF�;���?��!���n�s�d�\�k6bIA�Ȅ�gA�Tj�S yţG���ìu���Ʋ�3s��E�'�A�\�ِ.��`�ܣ;�~�vH������K% G��tQx(I%*C>� OTq���a��I�
��D�0_����)4j��,H��(j��V\ �5^W� �nסt��j�����[ 9=2�;M�ó�p�.U�5u�H�@h���'-5/��P	�C�/�*S�׭�ZY�:aJ+�@W� e J 80���Z ��2#��.����$�Q��F�,m�t���^Da�ĳ��'�n��D5.I�k�n#ɰ��|�H��)�� �y�U��S	�f��̑Q�۠�&s
Rּ�k);�IItMy�q���ܖ~.R��%j�?����ّ�$�5Re7��{���o��+�\��˕Ӿ?s�����`c�S`
�� �{c��tE��46���;��'y���p�̓f�"o��Wl鰹�i��̕j`�>��/�S�%�R8&���R�K���o�XϿ���ּ,�s�I��u,�3#��#���2��b;Q�\PE��r)Y���V��8��L��DW/X.2 m�{��n���8h���ޘ��1=���wϺq�>��5��{���0���K�1�E�EEyΆ�Ѩ׎ViE��m���h�������+D²�-����nPދՈ�.��
&�c��p���K4,��Ōj�"!��>K*P[��LiNyZ	�#��e/t�؉����U=�^eJ%E%\��T��<?�T������_r�stׅ��N�t5Bg�*o�85�ڮ�i�Z"��G��jA	�>�B\��#%�mE���6�C��GFwަZ�����Ui��k)"�����u�a��ѱ�����V3B�@�/��Gk���h}$�3�i�m����r�Z2�����EVtB���A��*i!6�*���9�|Z@ї�F�s�S5���>���p��#� w��^.Ԟ[��sP�v�_����v�U������%���3��®pRo����0�ӻ�^�F���hԋ,���@��Ǳ�4y����D�/���À}-�>T ��%����m�ΩG�	 ��ԃ�\z��.�V��9
�N�PI*:�]�i>�y	n�C��&�粰C,wO�zu_,����Ө��P�2��^g=�,K��?��1˴�Y�Nn_DE.6�H�T7\����u������V�x��=��x;����σ�]�-_f�:sQI��?�����'ݸ;t����b�*v.�}�(:��C���^�۷�$� �H�Ş�4&(2�@�2�=^"�,p�uw̦Q���A�
@F>�f�#�=D�/
^��?~�"�&J d�9�A�@��T,����YUD��IE�#<USt�Q����.�����X��@�.
�m���:�ƭi3�-ih��^w������=]8=��,$�A���tL2�mC�%�9�H��^��(�y�TBq3j*ދ��lq
HA.�*'�EE�X#R�^%8���P%%H.��M�pU1�I�[����X��'jx� �/����V�m\:/H�1�ye�U�!�g�y&���W�v3���|�P�~�E�Z�G �G���V��؁�0JXo'�!�u��Н9�(��Q��2`q<:YvU�M�6{ni%��P�@��:ETW%�(��`Cy}y�y@�[�?��5J��D-�.��	��5�kWU������IȽV�NgQ�,�˲��j�j�Ix��#!!����a�׉��K@1��vJ������{08 �`΍
�V\�;f�3��28����~`%��1�y�(ۻަ��e�l��<��)ݻK������ն�%_��C��'�^��$�E<�Pƭj�$Oڌ���{YՁ�Z�ƞ��ޔ`���7���-XC���WC|s`"8��?���<?~�r�A��!��(�hwŝ7r��|_����]�)nHohrJa�$�|TjT;o`�R�N�r��'N�[�Z�rF�ͼ�c!��~�Z��I�/��)8S�su����1�x���JhV���]����������EwQ�Ѫ����̽��#9�$��Ï��쬮���;��[;���̈����a!"� �Έ���~;�b���4�� ������@iؽ��}���1���v��L�F���+�,�D�2D0*�@���yYO� ��_0��^��Y���ܾ��쏾¯�B�rĲw��m9����b�ʁ� �@�`��ש�]���}��x�Sv�+XN,]�)�����,�N�Go5%�<[wC��xX��|��sj� ]��nV��,�J�n^�O:�ј��Zم��6�7c@�H�ű��z�]Cnګ�� U	��$�7;[Y�D���E��<�4��v�U��&^ۅ��Ů�Gi�����z�ܷ�'{���C��>i�/%	3�)�Ĕ����_��J�m�:��n��V�R��d�/2uᛐ�+?��ڰ��Ö�T ��'�ϳ�����=P�gw���>�L�v?���Z~�m�>�[�i|���T{c�-{��q�N�h��lV��8��T�+���P�<�6����!hw������;6^�����b���9�V¸�'��)�v�^vי&�#��ډ�ݗϿ��������y
�v�D�G�3��l����+I6�v���#pf>��b��l�����v$�rn�����v�R�S���;�u��,���x��h� ��;�1?���z}�<���_ ��rX�U�`��?�������I[���47���W�xe�W���Ȕ=�1W퐅�W�Cư~���[�������osQ�_@��l{�{�·y�G�V��K�<��9��>.�~��^�Bn�������1�/C�Kă����|�f�Hn�M��������+<�=���<��S��|������;� �*h�B�nZoB{���O�K����]��#����aJv �s�ꆩ��6�p�t�uhwC��\��꼅�:s>z~�LOł+:��! ��@0�T#���,�,$w��3>]2޶R��=���EZM�;��w�B�S�MY�
v`L�AA�!�S�Ll��0�	2���aVH�1&��aw)`��TJ)
��E�[���?-����Į�K�j����f�-�#�:�<q��l"c�;��׆cQ$��0=���Al�`s������s�9D[fMa/q�d�S,��D��|���n(Jmn�9�р�Ũ�}a���5�)��6�=�PX9��Q�7dr ���������z2k�,b����c܌ց���~K�Y���T�I �i1����f8��S񳗂M���5���_|�����kQg����[V�Jߚn]�&�(�1kG��@���(�tf�U�X���8F�#ʤ�Ǽ��~~� j�O��'vA;��Q�b�R�E-a]I�"����*�-ㅵ�r�1?c����w&�[Z@����>sf�*�Z"���X^�h$�N�=���H��jAlg[|+��fmWV����z/�D���q�4W`�w���f�hs�ϳ��p�(+S'0iA?*Nb�i.,r�����T����.�Q���_��E�ۇ;x+A��Gr�A�:���GRM=��㛏�5s�ʸ�4���~�<�J˾�Glsv�!#���-z��on������/o_�Θ�s�e jv��Z�6Tƃ���6뛎�ϒ(i�bs��4k��F
Ƅ��r6o�����#����#]��n��ɱ�jۂz���o�G���׾��=zО�q�fkB�,g���屣.J����3)��[j�TE�R��V�Y��<}ݘ`m�k�6��f��1������3؉LР��n����α�ιw�i���נ��FeS�q���Sj��k��1��-禮_>^�T��˙]7=q	��k�3_�2�x�MB��N,jh�8���/,�A6�j�i��#��ߩ��V��"ܖ@�/`�ٺ&��{pB����/�<�E[0�_r��#�0A�G�C�J9�&_�΂���\'��/���0�C'��Z��'E2���U ;�'��c�1L��C�������S<cj��������s@�p&D�j�g������e��.n��|ua�)��N�R;��?�XS��� i	^�zީ$0��S �-c���EC*��]ۥ�����`�OI��-k�%��{Bgq#��tK�,y�f*'�4�xy��z/�0�kִ���mh����ȧ�n.��]w��0�����k[�1�j!�ۆ��;Ŏ��7�a^�r#�g,�����/K���Y?�JJ�E�^�m����딁:�;e�	�+��'r��7N�q��j����2[��b��m�WU��1�*$���mMw���WvT��~�>�0�y�WI�N�=�tm���b�D�K��F�	B��W K<h:=^���ܳ��Ʌ�|lKZ{�}��x/;�`�&\��)��	;�(@BƝ�r�Xُ?���p��E
���a�IPn�mdl�2��2w�&���Gn�`?���6pކJ�DPƤ3z��jW�&HP2�]�<���я�a���pP�f�Ԓ�����iC��_��{�qm5���.�X��^����RP���:׷�,Kh�ʰMr�\�Y�Cm�f�V�ث{x(Kp�^}�J9RX,#l�WY[כ�!6Nk{��Ǽxٔ�we���}Pf�,���  x��Y�Z���m��sP@��R:��͈�{���O �4���:Ⱦ0����0��2}�5m6޶�� ����no�v���V�M�r�-��T�k*�oͨ�����![��`��b�e)�xf2G_Z5�2:�,�N���.�l�`�-�,���S���_�5�Y�7��>��t����u�k]����4��Ʈ�
v^��tw9�<'0q0�ہN��wV.���iH�Q�'ZPd����ڞI�=d'bkN���3\����
S`�;��������X�_-��3��(�6��E�~J�������p�I��y���=s��]Ks8�����/�֘���4тl�*%S\�h��6ԍ���遼n����s��'>��?H	`mE.��hռ�v@�eyկ��Y5��j��p�寡sy�� ��Lg�,�	:;i��g�N6�Kޝ�����Z��O�[3幔u�:`Q�N4�3�2|�����߾���7�/y|kδν��#��d!w�7�ˑS*��K�Д`��v�Gjg�R:s)�A����==�H�`�AO�m�9�p/����+zkn�ڥ	A������}� Ye.�m���{^3�M�J�E�G�X���w�/�fq<vl��)���.1�ƍJh�=zi�4�K'�Jp���W�"2j�?h��=HP�w��7���,e_l��&꒪�(�SV�����r� V/J��s�l@�3p8�d:���õ:7�w�N�J�I/p�w�{���h�լ��}�����K��׌<��q`D�٦�2��G�fO?��4��y}�ݏ�
���������ĜmnvL��FK>��N�t��� �|&WM*��B�z���b�}��K�@�?y����pn�y��sO��n���t`,�'���c�%.��c)�F�a�ڑJ��c��ɚ�p���l�"|��"�8�)���v�ߏ���}��=�a`I(�bIB��5������ssq�w&p�G�q���v�F*Q��lg�D|~~�f��ˁ[�I8���tB#�� ZQj���kZ�n�i����!��u��]_�s��=V�o��^sٰS�x_�Zs�+?(}�+�V����?/&�����i6�:�i)�N-���6��
�/��ړwA��IT��\`��T��S�g�v��ә� C����<�vU(�>�����\�ݽ���4��lf�1�i����tv.y&%�e[�q�ˎ�^	Jp��p?��(�����H�/�l$�"�աhJ�"X��XI�ݩ�=��	Qj���[��-�R�u�,�_��>���!=><�xbV���u,wA��؛i����	�_�(S���o�V�q��Όp`�7��@{3�,:j����h���t���d�'^d#����)�-J^zׇ�4V1G���i���y�	ǿ.(k��B!�-�� A��^۪�7��[	�!Ӏ ��Kd=7;d�}����U�?Y�TDwvS2�gTX��{Pk��C��zۚ-���I,r�R�Ũҁc��l0�:�R�1OFv�B�=ڐb���G	�nQ���g�ˁv�;s���mB�c*q#�;˪9�Y��U��^̈́�LB;/��^jץJ	Ӭ�g��Cݓ��#Af��j����љ���^���͈v�:cL�2J�&�{�S�o��q�:�ŃEE��.*9@aYoָZ{u�. _{:Wwe����p/�k���J�:2|��+م�:��fam��2��Iݥ d�{ti��-T����ʶ��:m���-`M�H7�X۸���Y�!-�m�L��2��I-��l����`"Z����l�~Cw��3ߩ���ܱyj�n�9�
��w���vg���9[�|��H7�E�8��;_W�ch���X���n�;�^�x(�k}��<����`�T��H���ߴ>��>(���e�zg�S25{��u��
.���شL�N~ɴ�����%��v��G�G^��~0G��������qȴsEz�>���cI�d��-B��B<�q���E	%0�y���I�~����6����	,�ѡ����R]/�B´�LEe�Ryŏj5�=Ch~7�	��ד|9�?�X�H<�����ש����3���O��T4��}|�bP��3���T��=�+�c=J�bp!h�6����	O��j�.%~�r_.��2)Y�r��q���rw+�'�c1v�	��]po��7�w��!���?����U.�Mm��v&ژ���.�{ wi�b#���a�:Gg��Ԇ�slQ���=֊��%�e���d?G�;:����:��sN�:�+*Z��Xb�7�L��b>%	;o������A�2@�ҁu�$����v�,���������j����(_��H&21�f%FTz�R7[�_���b.��^,*&V���� �`�/cБ�| 0����m�I�c�~W����j����:�+�_��fe��w�'
`Z��H�+u��Ϥ��v�c�� �HP��(�i2��5̍�1�N��=�F�b��M�މ]dQ�ɪ�Y�r�Q�2]�ᫍ����O�Ŷ��e�����UI�w����o�ý��g�����w/K��G�5���D,s��T�Nu�mX�e��q=��Y������܆%��BRI\��.t���~
wc���᷿�-�=߿��}�ovzB_��0ʮ/J\�����	R `��c�y>XEF��x�mhX���Vwѥ���E�JO��vn�F8�fmk�R�������{tg�˿o�J��>Q���4iU�8��Xf����wk�/�&�k7�˓�Y�ys�H��!J�ϓЫ�|����&�$p��qT=�b�ln�.�Z�{���1 K����g��8��mi����\'w�h�s�ή�մ�&P�@
cg�T-���M��da1�Y 3w8��M��-#2�戮g�54����4���(����O1�]�����17�lq���»M� �����̱R v�b�!e(�d)�Xd��2���>��)�L/bd!�7�ח�7��	nͅrM��v�V�[š�R�+}�au:o8�Ѐ9�Mr�d)nzqx}rP?	���,`ل1v8+���q��iR��o䎜s~X���6#��U���lx;�h���V��\��C�����ZLpq>�k����1��MWK���o���N�B����-ܻ{+1��=������&;	y�>l�?0�EQ�I6h>�������&���m�"�D��*b�ee��i|��N��IMpl���'3^�L��3Խi9~2�z��κsv��A81u�<�-���W����5<@��_�䖌I(�`�T[FB	�Z�εs�K��ѿ6z��V`�ng�՞�����9��C��;j��t��R���̴Q�g�ci��K5[�rX�9���Z���,�_oAu�t-�[ �e�Q=]ߦ�>�`����[�e�����Ew���Y{�?��U�VG�}O��Us��-����yo���B�	t�9Ԟa{�Ѳ�A1�-J� Ң9�@�䁀�C��0�h���B�t;�4�����&1�OV�L@?t8�C��#J�_�I�D�3C4��A�v�W##s��͎A�@u.��K���L`߫d�\��hC��`X�X��X�B�6	0��Q��^I$j���t��wr+ V#r!bR��3��g���o���u�:;��:H�.jԛ��\~���9t���bY����}~���y��Ʈ#P2{�<t��n0Q�#�<~'�|}!�"�B
<�%y�K��%v�ة���;��|r���Ȉ�j Vb_Y; '�! ���e,qb�s)�w�m�V.������� XE������W�4\�|�Ǚ%��tQ�R�+�珘K���sC����&B�`c�+cD=,���ѝ���-EP[�[i)Y�-]��kP��xxS3�M)b)��}c	+����v�^�!�:6D4|� �nWXpx��`AK畍D��Y��4���X4'C���9}����H�����P��ZVo��_�:5ŉh�����{qeS��9�o2�\i�S��x�޷����;��w��?p�B��~J7y��9~s�N讎`q�
���,�v5�]���UM��'�̻f�}?t��� ����	`�Bv`^s` �����Ç��~	��c����?�r��l�_<�?�{��Л�9Y��`1��k�=Dg�]��=�ڎ�u�U���t�j�V��}w�`��ܒጄ8	J=����Uvn�36��M�,ec�M���9��������S����?�����Γ�R��C>�Ǽ�e��xRȷ��]��O��tߚv߸���4�w���Z6`Á�$��Y����, �� ��[�L;I�$ngǄu��y~��Ak?2P��M�8aa�m]�n3�c�ج������#7 ܀���^�0���t��ҙ�w-#@3k�@� �ۑ����}��NZ�|\��c�4��f�P,�7�FR�8�N6F����A#h�LA|I�H�$CKY����xff��Д�-���`�r����8�I�^�36�m��>}bV&�9��1|���0(���E�:4�:��qy��Ǧ�5:[���Ȉ���qڈ)�O �����$�i{�r(�]��S���)s�P�c3U�Y5, /�M|���֭pD�I"�u+�rvf�m��d͚����iNѠZ�H쒡̊o��53����59ZM�.�Y����/E�����ȼ�9�����1Ƕr|�K/!�h !@�;�Bp�@�Wp�:K~��N��1��&fN�e\�%^�n�����������S��s�ףu�PM����_�����!s���� G��8ub�غ��ֱ����ʰH��m��)5� (Ė����֡H�?�pӮ�oywg��������]95W~ZkkC���@������]�m���������̄�@ͭ?��//����~�w5�6�0�P֧���+��6�e�Q����'_v���fY�= �e�S'Bu2Y�����pu��k��{��������i�"���E��3f��i�<CpJ�)�]h��P�ּ�ntS�w*�L����b�"0f��,����� nΔ@�y�s���&k~s^�0����T�1���>
y �o<�R ����e0�}{41Y<���:d�'�c�}u6V�ִ;���~�ي��*U���E����^�E.v�^=Yy>��  ����d�xc |v"�؏���ⷝ1�ňI���3��q_k�|��2�/~#ٹ{���\�޲�s�bw�qp�eR���=Z��z0��<�<�`��4_&� ��dWtۘ՞��[/V�7����貙�����(���J�}�2�!�T�2@��y `��K�z��R�h=W�BR��5��S�̎gyX!(�����NɐR2�}B�ց��rV�ִ�6��!BN�r/6���dzM*�b7�Kg N��T
o/��������푥�1�� �����i��X�j�K R���O�5z��?@�V� ����!�ہ����-��,i9^�ҙ�.�7;��\L�OH�ɿ�q�Րc�O�r)ag����~+V�d��	��vm����O��^�r�}�~����o�a�9�6��wi_OW �w��*�����*�\��(>�Σ ��'���B��i��o��H�0V�{�U޷.'�ڪ�i0�Hd�m�5��>?����%��w��:#�PPw��oڹH�S�h�籖e�Ji�u��N�l3����/$ʀ��m�͓��`睳W��T�''jx�T�i/�Bp����ْe�7���%l�m���
��s����1+��h��_���lx����`��m����k�%0������?�����x�cY�B.�c�F��"�q`�)1+ ᯇǻ�/K$���Y�F���ӧOl&�$Ҟ�Me{ˆ��ޏm#Lӭ	�6�Y��F�#���6�';`� x��3g�w�(۹�:�e��9��{{}f0d{s���#7��'���	I�/�7��T+?�8�(�`���1]��tvcht6���AF�K����W/#��3��씁��S������g�)l�Z���%s���������Ǽ�������������$8<��P?��ae�d}���{��r��	��G��3	�[v�=C����7
��P������z8S(��)Kf[:������n���,c���,�}�2(�:5H���R�=��Fu�@&�E�eH;��-��`NM��6�^�L���h�c[uS�����KT�C�N������o��o�����8�˳��v&�2^HFJ�h����fv�~�J��^�_�<����fV7��%r=��BԺ���H� �*˂��� �_ ���`s��,ή1�p��Mb���S��l�v��qь��$�wȌur�fЖϋis�֯iY�"�q�<�lm��V�����i$V_}�y���_��wP��5��#ß�G//�}���S(�9�:��a�"�,�r�`�<�kG�/���Π�Χ�=&�h�����g�e��fJ9N.Dh�cȬK��#S�D�)u��q��O(=�߱��j��f�A�5��{�Bwj�nB���HunJ�@k�3�%�-)�0�g؍�Y&j������eN���i��V�˱���f���-���#�7x�>�oyO���_W�����W�4T���>R��9�NU-9���>�ivv���B����ϟ� h�)w[24^__�@�n: N���yLhZy�Dꂗ6�/�/���^L�d�㋒$���k���?Z�r&�_��YL�E22G��%�Ff"�wV��}0�Gu8J�L�%�-Ax���y�ؠ��v�-����jL�ӟ\�OkV�Ө2�ݖ�b��{y������ip�س���{3�5�&Rv e=��;z�	��oy�ؙ��۟;�fLX����}&+��!��n��<�<��3��z�HPivE�'$=����w|b��y��d���z����p� :~��	�tL�w�1�o��Rǋ�H�����9YgR��g�^)0�B �����%_?�M�� �ױ4�Nw*�S|�+���;�u�ξw��;{v���P0�:�"���l|�h#��rP��>j"�v`Ki��� �HJ�>�W�O,�.��[�N��f��-.S;����6Z]#[_�j�[!NM�;I}s\V�pT��-+|u}����l}��#�?T�zI�~�|�]��k�^_q����� ������9�Aw�����Ľ���{kfC6�¸D����+�9��L6�MO�k�s�=��L7mVS�N>ؕ`��5	m�S���~�=��o��LP����#�X�{������R`;����������7�c��?^(�v��վn T����� ��1� �k*�ZX���y����d_Q��͂���j�U1Z��*��R:�A`� -[5� ^��2>}��h�hbH��Y�~��lPK�,��H�U}9�!6m��g�bgH��`MAB{n8l������7�&/�J��4oCzH&:��\G]{�%KO(.��Hzڱe8�)n R?~,��������q��A0�7��V��͐�bs�^�/`�n+ ]L4�<u�&8�'^6⧯��� ���`[%V#ep"� �Èn�0�a3��3X�纩�⎹��q���ۙ�h!��ީ6�ʛ��C r����:r#�OS�<?y���&���=5�u��3��eoyF�I%��q�t�^'�D�.Ԉ���v�����R���q�Z�9�v��_�DZ��#�7r�7�ʮ� ��ݣ� X5���v�l��_~��3bؠ�;�&
�E:�[n�Q�u�i1'0�M8� ���S,%�`�P6�Q�s���i�Zt��XS�l�vB�,�9@䎨Q�{�<:W8��r�V�);��܉�M�L�"�Y��8�c�|��2G�+C��d0�Yr 2g�:�NZ��{�y�g*e��1�^����d����7����b9i�	Б~Ӆ�����ݱr�^�{6_�G��9��J*�l���u^�W�d:;eo����G�8r'����y�~��M`d����1��E��u��;����ؙ/%���ބ=g?J0a��J0�^,�R��J�
瀮L�j�R-�u��V������y7?tc�)h�%�Gw�Cq�=��K��Z��oY\,��c�=���-��?�;W�7�����������
e<�$��)��$m��q7�L�X�}��ԫ���髕i���� ���AC���Qs�:� �d7H�W[���l��g@<���$�{����`�������Ǎ�vq=:�*-G�q߅��̹̀�K������"V��T��b��m�g��!�ӕ�K�J�P��kW�q��
�+�Eb��خd��H��!���a.X+q�5�����+�y�d|��t)	�$�spݡ�K`G2�|o|����u�jg�e�.�58�=q�%�f�mth������p��i\��07z	}���?��d�ŏZ����m�Ʋ?5��%�����R�N�'���w_b(P��<�
׀����1v��,QO�;�����F�Yi@nY&9s郞��	l�u����������p��lfO v�t�jVhͷ� �����u�9%��(;�]�����b��b�����W-В�?�J� w2֯����lNd�bj���J�yW{e
Ί���P�▱�Q����;5��'Jp�l��S�}-9[������|����yM1d�_%+o�d��֔x3Xپk��s�yzRu6 ZǪ���]��<�{�\S�p�x#9����:�.��)��]�m�Xt}o���=�8���T+����9ө<�cw|�tWS�uJ��9��f�t�`�T�y�f@گ������������I ��g�}Ѹ,�Ԏ�h�]�.8c���e�{݈u-_5v��?h�BI�<�|���i�'���~����C�s0DT+��i��&ڿ�����jh��2�CY7�U�ᩝןIק~�X��\6z��h�ze1�Da6F��jĭʛ��k��{������=>���a�S*��)^��tu��h����ܲ�X-�8�ф�:��l��`���s�ɋl?h��b]�?;;e�������GP�A�t��ג�E�!hk�?�����e�	G`{Φ5'Fw�D;%%�9e���v��M��|�L�ф���y߬l+�n�������9<}SM-:俿�BȺ�KGtt"��,P��~f6��ޞ����7a%|g�زt��&�M�c�x��n�h��'.�x��u��I�ؠ��3�>�|N�x`���{l)���J����#s��	FϦ.&�(�+�v��K����7��'��b�������~)�u�J	 Io���xX�8��?by�@˒���u�[�Е�������$��ڻl$�H�|�>>���Ȕ��zf����A��r~�i/�����\N�Ψ:���u@��w*mZ&��]&�h�3�8�F1��Vt��}��J��3_���Q�</l]>���������3|܉v�vB2�&2S�ZZr�3�G�#Y �g�f��ՙ�(k�/�mq��\Y���[Y���A�J9��	�t��n�I��5_�f{��Ţ2=/7��~ݝ���gn��FS���Uǣ���B*�i�/�]��S!g�sHo]�;�ՙ�	�T�\����|Qg�k�!Xx�fc����*�4N�yK�ag]\T�9ѱ�>�p��hB��{��Żnx��@n�=)tk��7��{�c^U=�jf����,��Wy����ld4@ �M̶�X�r�d-�6f]�c�ٗ��|��>&r�!�(Ⱟ�*����:��D�b�(���P@�%uz�bs'k�Б�R�/�7&X��i%��k��� ���> )j|`l∲E�n�؛�Q{�l�a�fvw�~	�	�&�.�\�*}�����O��쳽��t�5��D�<� Xc�sꚤ���dʓ|��m�����m�@(5����:� c���d��Av]��:�-b�q�{�0ZC�]m��~������e���S�슇�ǟM	$���K�G�e޷ݠ0�R~%�k���}���ꠟ��
��I�x2��!MDb�D�[�L�g2��;:��+v� !�=8Ȟ�u��4�χEZ�������d���P�AO��.�ٌ*�8�L�mF�t4�U&�cJ�A���~g�0h.d��p�6�嬤WO�zO��J��Svb;_Ĉf�5	�a�od��jg���'���0[�[)ے���^F�c��8���`<.˯԰!{��v�]�d�4�l^��̍�w�<}�˳��h�=���f�*Ʉ���^!��q��81��&�˸r0�l����>wo׸�u�M+���~��z��~=�_Ct?��9|��N��#�gb��PƔ�d�	5�w<+Y�y�����UR�<%��N>�ʂ�#P��q�p*Mnp\&� �d[�N��y㞰	Ld�fB�A�>?�~��_(�������v����꾱��r�=�#�5���{7�J��`���iQx������)|~�~��9|y}*,B�!�:��XR����g�ɕ���w:�����Q=���(UB���	4��&�:�s�p�M�n���:������gvՙ�z����	�M�٠�x5���!�|I{�B(��B�/�_�s�ÇGf#F�kV�PQ2�3k6g���H*s�f��2b�jQ�捌ul��}4� 7[w���z3����;-(���x-�����dx���bjz��:�P�:	�F�I6�z6Fb��D� ܫ�B�����w���D`�;-9���'3hm87d��ݝ�"��(�)/��,����6�]߇� ��0�v�fҏc�o��*�;0���l��y� n�����ݾ�Kv���Y�A����>��r�� '���ܳ�n�1���X�2�6�.�7�P�{~~c=1�/�19�Ɲ��ϼ�
:e���ԪF���؜1�����ϝ1�lD"P�L��2R�m�%�s���{J���6�ł�N�ܛŘ-`%-Q?Ơ�<g�5���[���J��k-.ړB�1�/�b�����l"�I�bYK�tzϯ:���!�:0(�&>L`ł�~#(�Ֆ����0�x2�W��3 ��`�3��:=b�`lco�4`'Q�he �9�|/�i*A���O�x0'>� (K����l̬h�Fo�y2�Ҕw�u
K�2�d�
�5���8��F�F���ƻ8H��u�?5p=�*�c���y{�L�l�
-�پ�|>���,��·젔�5x��? v��j�Z�� �����L�w���I���v�ά�?~Kil�΂���sf�ˑ@lT^|�����'T��k���S �Yf=�S��c�K�q��_�zw�pM��Qc�>��}�37��[c�>���ʼ�q��>��+�0��*5���ٚ���1����7���w3Z�C�>G��@���VS�c7x�V�� �q2���a�Ը5$��o8~tT�vV�YK���	\�M7/��DQF�	?��9���_�5�$���S;���ω�� � ��A���J�'���r �Α���zTsg���U^��w>$���\���yp�O��ƣ�*O8�AQ�`n���b���>��U��٩ ��\F��mc���[�TL�� mP�vO��	�
���%� ��1A"�?���'	��aU��)5+�2z��L��˲	�[��q��umi��E��IƎ�kF�����~p�[k�F�'?��ݯ4���3�F`ɘU/���x�Llt�Dv����*�2y�2��\��DL�4�I��Y���sM1ݿn~/�^��pP믙TE/�Z�Ɏ1���H��
�Ϧ��O�G����&.m������P, ��e�<�6��u�m�gэ�7�c�?��$c���e���_K�u�������Q�8j*�έ�yw;�}�����>�Ѿ�;X�B����ԪL�=n� �`�꒚�yf������U�o qVT'��DK��A��р��l> �z�����-�Fn�r<�Ϳ���.s�3awfU�[�J��u�9�he]'/l��&%������v���y�~��
O��C��j��䍔����Y���W�K��Ȍ�� ��篿��������O�>�#˱^_fC�[��y���~�;�h�M,��xT��	[����Q�z�������,�A����k���а�Y(�u`b��A�z�/�a�����:7D{%�&��lu����u�R��q���A�c�ƂǓ@˿�u��w���#�q���WDd������۳Nv"���p�`0&8���N@l� � �aӇ��k�0���D�l8��"�Y)L0&RqB�Α�0Řs�����zż0�7�ٜecX�
�y[�����b4d�2|�zܤp�0�߷�Z��jw��~^�Ԙ/*I�8w�aD)�͑!s �%�5�y���}~yOO�v5h�ΐ��`�(YP')9�#>�d]��&+�� "��Ŕ-
�~�����X6�}�:v��T�^���od�tƲ�A�B�?��gd����"��kG�Z8���c�1_w�����C�嗟U�I���uҊt\�^�,����ק����ewK풆k9�5xy:��ġ�Y0
{ۦ
�>?1W�����������e;:� u�Y�^9�-��5�=�V$ѴY�o�Q�X'n����L��ӧ���\Lgf�����hY�.�p1���dP3׎��auVK��L�t���:��y�C*@����[�����-�TbE�mA��@�l1�%���˼��9��_��jߣ1���`&x�@n�	� a0O'f�1Ê���"���������>��Ǻ��� ?8 �pŕCi���-�!� \h���4'su~+2��I�@�Y;�$�3�H��N:�r^�L'��x��~�ڙ����Î�/w`b�B��\;6ǒ������,���HܕD����M�$6�P�k,,��X�>��6��Y�}i'L�l��un��x����QLվ7\#��*sEr�{� �{�$֥T�e
b�	UϡY:v9���Q[ �`�/�S��-;6b�[8�f6�8)��zx�c+ef附��>�H~D�e��}��aa	ș��
^޴�o�f������(;�b����8lL���d��x�E��R��&��=pJ���ڶT��y����׼�=��ׅ���� ���=�x�>}d @@4���C0�3�g��v�K�	���E
z.Hh���k�����ث��u��0�}��4pV��&�� o
�o�L� x��&��;����,�DZ,x+a���PK��~G�Ԯ��6A���(f��� �0�]w�%m���$}K�%���}L�3ǎMX��x��2�i�{>�|ɢ��,6b5��=�����4 6B�Ó�Ո:zn�T��Y�����>�]t�IH��|o����2&颞
P�z$�y�%�)&�ʻ���f)��u��n��%����1ݽ(N�#�n�(@N1���n�/�,����yl���U4=[S����dRۄ��g(�չ}�T�@���n�}EكJ@
{4����˹h��{2}�:ȝ�x���7A�?�H#�
�hڙ(�X)���Bݭr�&_ʀ�[�0К��i��l��|��c����_3W�����i�:�&�,�t����Yr_�~6[}$����:�3`
1�q�{t���F�`�8�ܸ/H����N�}�:�4߂���<o�7 �z=��R��B �#�%k���N���-�q}S�}ʩ�+w��L�W�`��}��b�V;��b��U��G�o9h<Gu�.�l�%�|���	��#r���o�!*�h�fs�';��%��:7irv�\x~�I��դf�ڰ��b��X-4����$���pCU��,�OǍ٩lo&:~0�w[@��	��˜�3A�!�6��#v�J�|MQק����`@�` �mr����H�Y�ߓ�a����K���`�u#�9�ؓ�1���{��K°YO��%��t��F�M8G�FЖ�Ϫ[�X�����L�q-'��\֍�����m��z��ckbq�8Ȑ
���2:�2BfP�A
�Zs����v�bF1ϝa��M���l�Q�cb?��|����׸�	A�����ב	ܪ�ڒ��r��A��P8�Ƞ�t���N �pQ'	7E��v�I�����Cz	��#5tp��������䆰�^���Y��*P�`����&��e��ߝ'�N2:	����mdF���n?����*�:}eL��]��r��L�-ᬪ+۲�<���JwAF<�V�� w�y�ne��;�:e����AX��\���l��k��E��v�`�P҈�}*�cK(L5�Oцz��\�{�W�ǻϧoV��R����7�Ljn��8N?�'���T�r���uf�[;�;콗�*[V@j�iT�{ʁ��e[Μ�sZ���w򞥊뱎�s���1w="�~�7�mx��Jѵ�C{"���[��m&��ɕ5�l�����F:y.~�6�����`��~
\���<{����h�X�a��wwګ�mKM/cF??��hO��,q�I��S�m�:�\z���Qmam�ca4odKd�����3A96V£e���b�E�V� A�߆���7,�V�)�/��D�@%a
|ML�V�g�C���P|X���k!̋� �_�jأ.g��?�T��Rm��옯�8��}ʾ�9ܝ/a� 6N=s�k]/p��r �`\�o��nxg)�>��64�<��h����Y�%xo<��%�9��5��_)����p�ce���O|gR��l }ah��=�US���w߳�������qV��X6���&+a&c
L�%3�B?x	U���ؑ�L���6�Y%vԖz��N�v�%*��|^ty���ː�l1 ����ؾX�lkMR��TRP}�l�ct�<���y�y�A{Ѿ󸡗UB;�e���ݮ�LDW�=�ý����`N(�Բ.Cpvps�h�����>��a�V�W���u�����[�z3�{6��hYX�|f�����4�A��XZ��ߚ��/y��_������X_��Jb��?w}�է�g`��>x�K,R�o+%�$ݲ挣4�\��A}?�딅YD���;�����1^\� �V+�Ҩeb9�Lm�%�s�9���
�'����aXx��(�,&E&m��\ew�^����ܿ��۴ɿ��\���5����S�+6����C�پ�A~&�2[	�J@�1���c`'}�EZ� �2d�L�	=J+��d�ͤ�7d!�<PS�T���;'�o�1n��G;��]�i4-29��MG ��eϬ�Γ�h�N�l땭�z6 �� �gp��)���zȋ(�D���1�.F� u�BƿVL����49���
F�3q%���F,g�kǷ|=/j�}��t]���^}A�Ig�?bcA}�n�m-,�CM�#:.�*̲�ǁ	Kr���N�vD6(��q؎&xW���G;�`��q(b�h	�v�$uN��l���2V�	��J\��MP2�uf�� pf��u��Y�3�^�h�~���}N!��a��i���������l��%h�{�k�G�U�j-��@�0��^X0ش����4>^deb8(��J�|/�;��� �� ΋�{ ����i��N�dٕ9I�[ݵ�s[�Eg!��Bc����a~��Cxxx$Ps��2 D��N	�0��|,�*����׹Irx a���)�n��o�� �`h�9�L(8�op��&"(��nw��֞�����k^���p�zǵO����ۋc�zQT1�o�x様���vw>~������j����Ō;��pޢ�1��t�-���8�f���b���.��9h�"��*͸gv�gd|
�{���E��dA4���Gp0�>�bfX6t��	`��9�Z��=Ho��=����=��\J��\2��c�٢��������z�N���� ї��aZ��Uz�s�[b�G?��ܽ������#XGo���XM	�U���~Hd
p̓�<!3u���Ќo=��?$�kJ)�H����o�c������� ;�g*��й���9j�F�4'�����WeTy/���~Wʅ\0e���:�҉Q;�yR�����}H.�s���b��%������܇od�\�-M��3d�4��6mHVF��5h�(�``G�� Y(��K�G *��*�lݛ�p	%�o�xx��Q�[QL�q��&J��<|x`�:��!�Qv�Xq,�};ѧ�ޅ�V�X[�|%�[�ɣ�fGc4��c�R��������;��|�}��w�#Cg]�6V��, �s�s�f�ڛ3F֖�	�*N-`gR`�Up'���sy��*	~F�`đl�3�^¨�ٚ��V;g��Bk��\0M�� 0�D�S˂'Y�X�9�$����B	����!<0q����G�p�!p|��:ۄ�<g���Rx/���h���{��Kpu���a�u�:��<�;;e���h>���v�`�:�#M�s���7Z5b��/�� Լ�k�Qw1ʹ?�o�<X�21Y��K�E�-7�U��z�K+ԡ�g���9V.��ՠ��Nl��?�y��
PV�P��2���ƈ�P�q9X-�,"H_k���R�յ��������w���ў�Lm�$�N���۟�ukISުdl8�����d�%�Ȩ�[֗c�ݓ����le�xx��nY�lI�`�)�}��5�A&���,<IGǺꡡ
;H;�����9���ݭc���v�Bi-�2�u���2��$]6i+����7L�矰�ࢰ.1�`���z�3��C�+v��ЃeD�`�9�S��-:g�X������X�޵�Z�o��D�:���P�Y���U�efB����]8���g���x�������Y�e+��}e|�!.�U<9Rf� ���
U�쎤�	=7��lhO��"e��`��y������"+��+�ȝ���9/�*�!1�q�M�N��(��P&"���V��6�`��s���k���_�R�l�(���ƢJ����1��s3�-�����n���y/E<�����6)�}���8�S���nH1-�T�F!�ie�od�TϩyHx*p��{��<�c%E�,����2T�|�cQ�َ��ـ)ьgr&����S���y���:����eJ/Fɝg�1qq5�j�l?�t$�vD�*yc�#,�j�@ej����1J{g]�\O�l���Ԥ�^$^�gm�x}��u. �ub&�)����u�ߍ�ʏЯ��'C%ot//�,��պ�t�: @����F}�y��!1b�����J=����/��Ӄծw����򽜤����Fݞ��H`T΂�ʌ5�����ӐsS�M��7A�4��lF�]ј^,�	@�rV��z&�"�Y[T����r h,0K���"�3��8*�7�e��(���[�l�4��u�~��#7��e������r��'��;vV\	�S���2+���q+V���8e�j��6����rϐ;�d%�V�_��[�o��l+�������}yP����J�>���=��~��7;������Ą@��@���J6�YG�NvJ$�]�f�`�h_���յ���3��i��Nl�)�0x�N��"�w�����+���Ns��L�>Vc�z�z���V�V��}|nx��'}c�T��W��{u�IǞ��L o] �M�fx��P5�\sMeދ��̍}8ޟD�2i�]8��ڨJ���Cah�z��1X���h��` z�0��k�{��FטBިb���r�!�1pg����;��J\͚g���s������4fb��J�2r�_����|��=���D&�����uϊ }����1��{�l~�woT)���u�Y�5M�1~d{o�[��/Зžw����:=Z�lBbl�λŽz�:�Y�e�/W��9K	�w�qv�l�XZ^�Σ����t��Ƽc^Z�pel
b�9���= �-�"`%��X��(,�@�ҝʺ�].�>�뫸���L�>�v����v:�k��#ɳ5�n��Y ����'T����+������jY��oC�L0�I������_N�HWJZSXoG����q�oRz�~u��c�dY���Z����Pac�K��*6k�[
�+M�zW�B1˩�C�769N�%46���.ML�\����~��z���G�S�;v��q=g��!������W�Ɩ�vI�i	�2?M�@���+��Oc1�����t�Eڗ���"5 Ƀ9�a�V�mho�R��	j"a8�Pv�m��@�x
o�7b�)���1|��	����a�f;?�5�2c���J��/a�<Y�+�@���*��l]aB�+|����W���:s$�C�>$�>2����y]z���ؗ���]�a`'U�Uof���T6eyta�6���dfSz	���	Y��"��nj�X���T�?f�Z��Ci��w��ČXL`uC��Ͽ���C f�����.O�p¢|UM��"un�
V���#���f#H���d��f�(�b{MXm
R�g[Ds�T��|�(
�
��8�����_��/���!Z�� Ke,e?帅8R�/�:���$��,�	S�c�B|���Bl5������Ȏ�c뙘�4:vB��<�l�\��I�"���td�k���Æ�	3�Հ��Wv��N*ِa�Z~���#Qᾀ:v���k&C�Kw�AN���j,q���IB�d�0[z.�N�~�3'� w0��+^����`5��ʥt�E����U`�]nvH5��DV�̹����v�Y�茪�G)���s�q�iJjb�����L�X��eW;*����ƚp���{H� ��<��%��@��ّ����˗�C<�[D��5�*�z]k��+�H��{�<��;f'E�jG�/1�X��6P�;:+�K2��N�܃eC�E�R��ۑ��w&vg��!x*N����J��<�_��F�lg��\�[�}	C�:NM&�� +ȞH�N�V�~������^���s��_���O\G�iE"�����7��O0T��Ц���xW%�n.��R�rE��{L�����C���Mk�Ϳ�*���A�<»ϩӌ;��@'g��>�}{���g�p�.��p=JR� ���>W|�f�0 �b�j��<ꠃ�F�o��p��Й����	�L��Г�`�ֵ�X��;юz�����U�[P�}WM��b\�qZQ�=WڐDc* �>� ]�������vp�L�PW�4�e2ڰ.�4�k���wt'i@��<�vdmJ��,G-L�J�C��ͱ27���ͻ>����{�aU�b*s��� ICfɒ���%�]<s_�.�
&��J>њ��s��;��%���E�q�Y����,�I+��8.�
���ԕ��Ҭ�Kف3�p�F@=rOW#��I�Ԁɲ����q-�$�l��s���y��QS�K��[�:I7N󯲹=��a���\���"4�N�])�Z��(5۶����m�%��yB�Hh��Ⱦ�!��qK����w��O�EdrJ�����♺Pg%�pO/JG��8�koKx�L�=��8b�ky��NT��y��6aw��n�o%V���Ԙ�ƺ4�,�ZF��֬ �OH�~��@_dT�E}��H��]��&���1�=[��R{R���Qc���(����^v�e~u~����jR����~���~\���&�ZouAm��0`g:��o]UݿY'\R9vR�zH��S��6��}'��p�7b����]gZ����,��UR�E���T���Gu_`��X�2	+������'Kؚ��v�;��&�\D�b��"l�;j���T����ݣ����><�}i��9��r�4�����-�_X>�N_ ��(�~�@ʑ1σ���Ljo�@(��-����#[�wO}p���E%Ѥg��>�1�c+����Jv���R�0 W�;딇�;|�M����H®�MR�ݱ����({kK���K]zlOt���L�w�V'1���)��nIdg��6�lc�y*f���D�����I���=l�eb��?^�=[y�6HI`�U�K%Qq���UFK�ؕĺ���h�"Kt��am����>)���:k�M���:�L��$�g�
� �@��}�󑌘/��R8��;���(�i!�>8�}�X�6���mԦsJ�^Y
�O��k��L�i�����l��y��t������@s1Q^��ٸ�~Q o���%�{��s��(�7Q�É"w�>�f�F��X[l���&2�%L�96����� 3�9%�(��ѹ��g���92�}Py0�
��:g�u̼��h{��Y�h�S�q�`�$o�Zl�\v8�0T�́�����2_b�h�޲�Ȏs�ًYk���k��cq��p�+��@̢�,k$(��1����}~����)z�3ڈb=oI�fW�b��|�����]i�j`ke��g��5S��T���֕�<u�	hF��������E�#�UM�E��5j����R�qxe�X�
H8��Ff�z��Դ�t=��͛򸽜��<'�S
��s ����s���^m���Wx��˞U����̦�nX��.�E7u�x�r����L���W��s����)j_�E��|����lbُBa-y�^%�[��>��sM��ٕ�U��y�!���ʱ�kW{������Yv��ډ�9���+�C��4�F �P���O%���co��iK$�kd_t����e��1V� �)����	�Zv�1��s]��+����a��3�\7�}=F����AN��"���fUW[�3[�r/��{kR��]�g�mX���P�4cD���Ae�b�S��w�]wf�1Ly��e��%x�V���}��.�֑��b���l��gg��.U�It��y"�G��Y����/���m��o�C�ص�-��b�KF9U>��N&��Gtz;��#�J-�7�s��e+t��Hڎ~�&~����3�j\�28��&Y�`֡K�L=�:�*:l@��L݋Za�����`�^������=	g�����j�;�%��1��;�����v��їf,k����k�`V��[*3O�X��5 Zx��=��Ԑ[Ԫ~B���ם'��g�/q��1�.�Dd���tyϼ���c���+�OlO�u���/G�>���.�A@��{��ㆽo���X���q��͟}�/�Q��0�IR^U�'����t[�+[g�@l��﹘�s��F�����͗PE��c���#ؑ�;��jnI]m ;Ѐ��u�~�ҳ=�w@���7]R�[%��kpGS������=��N�NR���m8꾋z 	��qc�F������T��H�c����E׉���-WW\l���7/-T`���tY�8w�`�8�#���3		��� ����oiRc��x���1�@� 㠄-5=�b<%�O�>�>N�Y �sl���pʾ��������˯�{A>}�9���g��O���^���������o�J�9JV$z�Pav�{5i���1������ќ�t/���1�I�;�H��-�ٝ�?��i��_���9c��Щ<��"��\a���9�9b�U�:f�G��Sk���i^��E\��C���\N���L�k庒����&�*6��qf��fK���n��yU�E���p�.&�*j02@��E�l����+�� ,D?����V� ��I��Q�y�X<X�2OV���iP�Z/��36{�L��Svn��K���(Ԫ�K�������9�-/�׷�hp:�M�`g-��ř(w[e��'�4۩�5�p���!lc��@��֣[Jm��d��^lJ����ꎧ������ �C��R;O,|.��J�n"����(�)8`����]B���?�1#�'ä��!y�P�s��O|sG@m�/�Z>瘍a��XZfΤ��H��$em��^]3�,e± �y�p/Z���� r}�T�͂�Eb ��; ΋4��d�/ڇ&���ǔ�{�q�/Z=�c�����~���ҕ;���'3.�G8�XO�~�~��2gd�{��O�%��5��+);+a'{P��AO�ӳf���^[j����:kL֪]�>����T�R𒄆m���^���3��j�p�3mgk��{q�v�"�p�cIk������_�]�����ib���]�|���n�~|| ���E-�e>~x�}��u0���H�A��`no߃�����_�L G��U�zu�8PЙ��L{R���ƪU/��$];m��=���Tjg���6>Xi�uJ�V�s/�J�2�u�&Ѽ�=�(������P>u�؎~���o+�'�3��,���Kl�y�mtX�qѤ�� �0MVN�R,�� �?� lq��DuY4Y�6ؙ���ߌ)�k��;����b�Դ,�z�ܙ�,���{��u,�NJ�C�w�@ٜ9c�ؐB��j����f4vBo���U��v�0���6�Q����q)����f�7�d�奱�������h��09I��3��u��:�8nw��'`����m�x��=�ALY��i����^]H�N�qG��EF@����>dew����*�����H���&�5���v�~��tt�-3�8[���
Nh�W�L]0����DK� ��������g�Fd�Gc��$��Ÿ�i&�\(z(�/��?ľB��AuA%cg�<dp68�cYd[�s���O��ƙ�т��WH%�OMP^K����s�~�r�.Q�Tk�N�Y�A�|���D\�X�Ią� y�_�t\k��#z���s��\��(�$ʐ��﷒�dϐLr�]�S�p��A����}���2I����z`r���$i���$qn	���8��,T�w�?��#��bצ���a1&JvuO�����#r�21h�������`�J��`��`z�D�ǲ��3����u�[e�R�*H���CHn�C������L8�%%��r�X����֬%(ۍ��:m�Mw���KqRvH+_ #A1��Wŭ]�u�jܪӲJ�8�=��r>�Ǖ���2��B���(�S�|/�����e!���>�L�v1���y���bB����:h�G8;P]^V ��W\6i�	���	��=;:��3�ؙ��m���6���3A�9mï��l�_�/��9��rd7��;]?���/�+��oUÃ�]�ߌ:�Iqۼ�J�=����v����p���M^7h������ގ�9����gjH�h�.�xus���W��`NO��VẸ(�c�r3�y����]��A�&a��	n^T;� ���PI_�{����L�sJe�0����Y�u`_��O��g�C�YLԅ�@��.��;�z�����5�F�E��lY�7��_t^ ���^�
(>˿�;	:$�����%H8����O^�j���N�-��4�Q�k��/s�|B�Ǝ4��6t��,d� ��c��b_��`�Z2^��^�'@n%\'�G�U4pX.���3'���m�����t�>�/ڀ�~'���/��Lҍ��a4�~��W�i��`-�#ul���-%S�{ڐq����}��}0� ��&�'�&�$cb�M�\s,�(sQegs��4���]P��MKD�J�X "ڄ7uก� }"c������+L�F��Cvd�q��=��/�Ǽ�TG,�8|��>~�@痚>�j�Q�t�\ �gf�;:7/���h�̳�/w���c���j��NC+���,qW��.0삌��*��Fk��q)�}�fK��fxG��d�5��I�I,P�Evhʓ���"�d}���b7�^� f�M��ooy�����n�y������ޮ8Y�+�Xf��[`m�T�����١��
!���	��^���z�I�5���Rmq�@�Ʒ��-YE/Ӵ[cN��,���(#֢��y��-���{����J������8�+�L+`�+�:~�R��Z�fn���={�C��-bnX;��d�	W?���ǃ�N���*��J]p���2�نPcG��!9���,�dx��;�6w�MɅ�j��_O�������G����V [p��i����3_nR�Y槐)K��	)�*=�{g�����X@jd���@fli9�8��=;�2y�)Л��$ �i�'װ���ö��k�9�So����77:%������+Ƶ�5�m)��M�-� X�אh��M����f^���nZ�� t4a32���^G��Cv�ߎG5�� 3��=�=޸W�s����I�݁�6T_��s�,_c.&W��4S�{"��˟��mI�D���Q	{3�{01��Db�K#$D��l�v�V]6K�����dqN�:g6�@��e����,����9�-O%��7Q�G%�*���׺f�,{_*��QB2�%�Lnm��H��Wz i(9�#�$���J��g�y2`�}_m_�m�5�Q ��A��ׇs���q@������!���'�\��ه9^ʵk�*��1�(�r)��S�+0��T0C��h9}i�Q�b�5^������3��#ΦLl�eZ,����8���D��7��v�M�
ƜL}��1���4b,v���K%`-s�;�E�}u��X�m��z����A�R��%�1�b����u"kd�o�M�[B`_���8j���mcҲ/4��d1�X�JB��l���`{^As��H�jDP�I�߿�x��X�������'ސ�%Yc����D�M����0��p{rF�b���l��b4�-K�����5��0��u���4O,�!^��J�6���YD����U�^�7�:���b\2���Bbz�م痧���������T$Wf$��%L�hr�5p�LS3����A��zx	O���rF�̉>���K�[�0����#2�C!����;e~��-�֍��Iݎ8		��A�ҧ.��@c�9pL�Y�q�],l�@sC����2��\���:K�8Pu�ޞ��.����G7gˑ^N��(�&ҠZ78����������ѱf$�w k$�Q�XNr2�Vt�� ���bGF��<�-�\'nb��I� ��'�13�X�5���.q���XT�I@B�1 �os�@*�p�ub#�0�"�C���Á��Z�� ��K)��`]�� ��휍��Hx��G}��Y�F�yq�E��3`�`� �1(�S�D�������G��"�BnP[��BڝR�.�P��8�p��3͂�l^_��2ZW+;�:�eO�����;
�<��Qs�%R 1��J�A5� ځ����K�I�X��*�B�L0v � ��2,��֣;����k����ҩ��ʪF2�6���N��Q5�*����Ç�����:�;�ȩ��)��
4~�ٖ�����a-��l�@����?ڽ��=�=(kB�C
j�e��H�9˩QGd0� �:�� �<�bʳ;�QVͫ��_��U�c)��ڎ&�)��e-�����B����hsfЦ�Ĝ�ɲ`��C��N�~{�?�1�H�h�Puʻ& c)\�r���)��,T(�'x!ZG��N�9d�y�CV���>n?��a1?,ph:qy�P[�:FHX��E ����)��}b��.υ%�)4I8t��0�[�@��Ҳp`G6�-���wAEw�<K�	��\ok!]$�kA��S7��be���<�l������{�.�q$I ))�����{�������n�TueF�CO�X��; *��=�笪��(������F$܎���t����Q�mi0.�����A��w�vG��H�2_����m�i�����{�"����)�I�̥
�ϴv��;��q�tZ�դoC�*�_���1a�w�{��O��
�p��(��'�#�mdw�=���u�$`c�|�
��N��Y��s����@��T�^����Y4�`��K�eϫ�������~������~`��>X�(c8��������#(G�́93ĝ�	E��:���1<>>)L����`/¼@�dM����k!�[�]i �|��� �E�+�������/\{��%}5��H}���G��dv8(���j}�.aV�=O%Y�|�ɴ��:X)'�x�찂	飈L�o��ac��yrAS�u���ӥ$��z(vۓ /�@au���f��J��%��B�_�������J,��=K2����nk:c��$�eс����A}����P@��H�}�Q���:Z��ҩ��#}��'�B?�?�3<5�����Xk��� ۂ�g��iI��׼��A�_\�S{�4�����߇�RvcN���``���繏u
UHڷ���`ҡq�/���}�3n:4jUu�Er��$���_1NP[�H@@��ϒ���o��[�P���'��ѹ���S���4�8�Ou��N��i	�w����#z ^Ƴ��Mt��|����6S_��y��ڟ��ӟ ?v���:\n�X�	C�̊��v&KTZ��h:`��- ��^��3`'ɗ�c���>@0mF�e�^�E}B����_ވq@��
�������.z��������d2 ���vf��vyϙ�덡�^�%��7'aL��r]�����؇��{�:���$�~`�-�yP���DW��n��7���|�-Hd�k���!�)N�!fɄ�׫|3���p���7���҇+g}�)���#|cg$���r�!�[��;�so F?a������Nk~esm�����O:��ysG�����9C�B��l�A�l.7���Y�\�d��e��`Acu`�
t�2I�U��@!��`�Ħ�EO�FT��l���?�X���=vC����(���!߼;�'`���Q�RoNT������xzz�ח� ,��7}e���-A�Y��=K������/C|��lD(��\k^�ƫ�^�L�0 ����^�a��8U t�N��	�Dӓ�q�t4PF��bA��댙��3b��}��R,�:,�
��H�Q��^���Z���E@�@ }�\�o9���qs}���H�)����e������cgMJ$��e��ŉ����jeZ8�J��?�#���9|�t��v���R�S>nȯ?�D�5��.��1�y��C]�L�YB=K6PF�����mx�v��v6 ��`T���7*��
 �!.���{6��ʯ�1	�(\�k�p{�߇�с�Qr~<6�} �no�(���=D4��>N;�T�;�ق �Y�8Xi�g\�3Z��`�v_��Ē�u�Vr��^���:�(��b�Fd��z�2%�Kȶ�T�0X�y����d5ǵ�Nb�@���+�a]���m��k?@P�@=��qo�D�E9H�?�;�t���){M�����t^���ٶ�����f������Q/����%����;�JQ<��ND����|&??�)�;�ka��8���55�Y6qs����
�6
�y%��+.����{�i3ZV�bT魵�^�0f��zl�ũ ;��΀.e眱�~e����j�jnk	K�bL�8L�$S��ч���#��-��t�c�@ȝ�U��Ȱ�[�����v�'����a<����Y�d�N��h
? 2X��$0�p��>g�'m#}f��Rj�$/k�_X�7�s0�O�ҩ��H��!Ml�D��j���kR$�XZu��؁/Am�|��ۦ=�xJ�+mdz%�#�JS��m.�^�li{|2��"�^v������t-)q���L�%��A�X�=�$���u>�q&�x���X�㢤�̡ق`����zC�?�tP*���.�!���PB��PrQ����˰������!�p��T���:�M����R��1�N�X�퀋:��Zal$1ަyӉ�s�W�A7t�K��/V�7+�:�WJ��je�
�681ъ�>�n�k����.��vǒ���6���Zx� �5���Z����J����$��	n�����a�|Y�&M�2���1�<	��#'�ժ�P*��l����W��@�(���M ��x�T�btJx��fÖ���Ϣ,�q��a����Q\W��;�Q~�h��,�_i�lB�	�|^5��>Ls4����ȣ���K��B�`U�V�����c���b|<�U�5�=�|��ظ���ު�f�
ln�BP��0��' Z��4	���a%�R�Jd�`lc��|86'J�<��q�6�rQ�|��jo�5m��� �<�5h�n�\]
����6�N������wb8	�q�7;�g��X��1������T�v�5���c����k8����=^�T��O�o=l÷����s��6���$c�q@�qO��.�	�ܜ:� ��
@��cO�k6�����찾�u�
�(���D-Rc�R'-���h���! ���!���
�c��LNwt�N�Wţ�ߋX��b��Z_�������C�����]�Aw�-�����o3�]/�GY� `��.4C�{^̢PO���'�:�
J�N��!���X�>�D,6v�!���x��j�o�1J����q�x���bFc ��P�h����}4��#�<���>���l�U'�a~F3����YY@K�e~�B��d���N4�d���U�,6�G'��l�AO[r�a���-p�C��u�్�-���!<]���G�&�?Z�[D��5�_�pB7 �q3��臇������|�;=�z{�� ���>��9c�ߒv��a	pτ������x�pJP���J�J�5�.&���s�g�:X���t��m�iQZd̓�h�]���FN��� "��d5?&�����`Sj�\c�k_��U��G�-�g��������3P�Av~��1���: u�a"�ssՇ/��ٜ����6�W������qs)�o��2�_��c�g�9��贊V�>�؀J<��	�� ���3���1�`܃1ϐ-�?�P�X��c��8�t2 �V�:Z�����J��7G`g+��(g�(�9Ұ����A�*ug���AL*�J������<�<��q,�ۈ��b��$�Y�b .�磺nN��NtƄBy��U^�[���Ue�Sf�8�wo��9�:a+���8�����Q]��5=�����>�3W���v�"��T����v
�J�xy.4�T (��s�^�6����$�=u^J�}2�S/��?5�<���ҢT�ޖ�	��l�
���8b~���/n�;������d��N���E�U�. rr�w�+�G��n��3@rg*.�^#S;���So��3��"/����h/wD�j��# ����h���i���`�@�TAgl�}���.�<����vaemf�ĠI����?��u��{�J�������쩄_�!]M��곃}���:>�@���ͷ�q;9���e���v]�i�M`#�^�9s�ip��䥡�T�+�E���!��D
�_�����D&-��#J�7�0C��RA�5�w
(Gf��0�;��8*u��s(�����ցR��X�jbqD yw���#�䨱�.*�iևl�'5��R�`@�7Y_��,�c�gX6�} �9�d�2�?R[��Ԍ����#ֱ��,����djU�j���o&r�X�丏)A���'k3�l���c�1��4%�U��T��ٚF@s��t�tn�9j��dNP�6�yVGȕ�X�`c�<�m�ĐP�h�c8�'^��/�Noe�*��C�� ���ǐV��9>??�����p�(v����ҹG����C�o�=^���B�Ǔ���\���'���u���^��b'St��suҽ��Ȏڔ���*�os���c��N�t���9A�ǆ�旯�z)���81���������+�R���D�O��kځ�Iz��`1Iz��Z��=�j�k��9��@���4=��� �lHb�D����9T��[$o�"3@2mJ��dׯ.l�
+	��=6'p�d+�+�9��k��v�(yE�?�Oݣ
#�_Zl��B\�m4(��nd�Gg/tw]QCu.oV���)|��1|@�*tG��cw���'���v��@̜M��?}�LV����� .���{���_�w?p���n`b�Ĉ;��Ӣ���/���[�iЅx���`�Pt'6�!�D��)lX�A�3����h����!�.T*A/��f��@_{?�R���]u���"Q-�ʟYv����@z=���;-��|�p�s������K~�@�̃��?�����7��'�]\�fg!��!3���0�9���T�W�ΥAW��[|q_t��W�!���w%Q�`����V���IA0D�C�~�D;���E 6r>L��6uu����h�z�f��'�6]-6i
t]Z�_4�ׁ��sC�����r�
�')W�Ͷ��+�-��`�@��R�+`�M���{]t5�p`���bg�ɞm��I`��I��ْ�p$����o�(b����y��Uvn��;Ȳ�|�	N�4�j��cI���q+�io	81=pC��C��N��-:I끛�8�vt��N"Ǹ8d�!י�(G���h����~��@%dvh�����P�kQ(x�&�QI�ћ��pVkCكh��yw�������(�Dp1������pOx>A8Y��d��A�x���K6�*�*�\���F�Ú[�_]��#*�6�/�T���'c/�̪�<NV��e�&Q�;��ɺ�c�f����83� C'߿|�Vph�~�k�� ���0�S���:;��Pf�u��I�(,�̜���y�Wwّ�3�u����X8pܓ�Φo ��v84ZcY_�_�dii����V��.%��5����kC�rs}���Z�t��n'fF�B2��ttt���J$X��N{lv�ʳj�T�*���������P�M�3�%�K.ǁ|ucf��WcW3�KZ6� 8@P��N�����"���+�A�!?A�[0��J�x�(�y6�Y�W��s�����ؼ5-��Ũ��p��d����SIP�r�j0���빊�/`'Z�B2zc.� Gs�[��V��+��`C7�^u�U�����R0��u2��
���!T���S�ښL.~�Ɏo@N�;T
N�Me�&Oj����ȣ&sd/O���zf�/���:]  WY3�D�����A��%i���@���������>��P��R�@,�5�,��#sd${0Gg��,A7}5L�  ��̙ f*@�� (w���h{$|<��]0�Q��l�+m�Z����Ě6{@rj-���|��q&@��E[f�O�OCP'0��dL�#(�E��w0$��J٢�����S��|�(�ɜ�2u1�.�ot[i"�B�����i}�`8���F�>x�$�i��6��'ul���� a~�+�u��
�!y>U_�e��,/���S�wq��s�	�
��֐�B�Z��`���^q� ����{�H�Α�o."�2ͻ֏ֹ#�J��X's� Z`E��|@��AM��5��!��H;�\s,c�u0���A�.|�qTY��K�1> ��SO0}s9 �Iɮ^z�L�4���j2��m*�X�t�2����g�����פ��n�=��>>���ٺ�E�i2�J�p&l�#�K濣�G��^�q�R�~P�~��
�V��53���</�F�B��[y�`Mk��l�)se���Ϙ�]���\l_j_��P�Oej�����e�M>�R�2��߮��:��sq`=��_�}���]���T~oY�������^yp�	X,$ �xzα�S�:�s�{��|�-����3�\��C^C�	=I��6�v���%�l�!��1����ٮ��Ow"D"D��Oy(Q�qn>��M���o����%�W���7g�X�7R�`�3��tyWHVz\\��d�O?�>��3�r��
�\d��=�P����Q�ws�ו���w�|y�����Xvcl��#���D������������f���7ypS:�P�0����Oԍ���,k����N��T '����uaS����-�Z[84ħ�A=�6Z���2����2�~�A��O���:   �� ��0�ґ��m]��05қ�FYo�N.��'�e��
��Sw<���"vb�@�f[t:G59��ϧ�k�r�a�/���	����X��  ��IDATa���E�X�2`< ƻ�T���K26hw:�s�Ȱm@��`�8`�N�݂)����D'����a��L�%�QA;�.d�F^s`gu���5��i�ڸ�	���s����&���-����cO`��L� ��k8$Ev.B�\�,�
Fg���H�2����s�[죊jJ�I�B�����(�����s��e���>��F��߰LP�|����/����dh��Q�wVɔm��A �C/=.S�?�@������u4����:hL�ē�?̘�������� -=���S��V�>n���X�hيR�ׯ�Z4�0ju!���;Φ>�T�NO|���g�qt^��N���	�oxΘC�q,�$s���:�/�%k���4:Lt�Mh�;�s�n+�j�O�� v�����+��bpy���#�q�n�ח�>.7V�<�e�����1{8����&gST���yTp�:C��H�~.�*�RR����Qw�X��j>�����eݼ��ح���^.A�>��S1y3��06�XuCf�Yz�-^L];l)��ȻcՌ�g���Cg'�=��>)��;���S*�^W���g0}�ɤ�h�]тJV��ץ��+Gy��jG1w$�y��'��`F�=8�|C�������,KA�cYr�q̓P�S?��/p�$��K�"��w���9�/-���0�܅[a�egOر�3JlV�K7�%v��X��Q2.Ʃ���#�su˒��숑!`'R{�狮= ��wh"1pߓ�B�1���U����u��<�����:��<#�k�q6�1�� ��#c��6�ʫʬ�Hhu��sy���ʩg⽭�8�ʼzw���tA��/y���C��k�/"�6O��y��5h�9�C���˞7�����@�&��5S��+��	��(8���1IeY؛�JWbh�ћ@�,��c��9���2�;c�YK�%�9��_�mv&��'�1�\��s�٘�^_�%��dS����|�A<�_c��l>ɖi;:�<�
f� p���W�0��$J Zn�N����ݳl=�ٍ㍧��2���L������F�A�L���D�`�^�9��-I7V`fB?��u*��Wh�M6^Ν����`Vש�)�rF�� �y:J�h<q��j��זx���3���ؼd&cM���
��Y���u�&'�S��׀���SJ����������g`O����٬�]��9~wp(��eM���R3�m�*I	�/����Q���gl߉�o0����;Ԙpb ���c�	���l�s�sܙ^́�l�}$����C���
��A���c­� e{b�bެ��E��o���qD����Ly��%�ԟ�:����#b�|�ǩ�Ҝ˳�d�������Xf%�vdR���X���D��RBয়~	���	_����&Qn	"�Tq^�\C*���T�$����pt��T��;Ë[����a^�������l�.n��7�!JC�>o4��cxx>�o�� 쨧�d�o�~w9q�*�/>�%ua�v>.��{^}��D�@�Ӝ�r��������C`b�?����V���ac�(*��;�-���2G����TMB�xal���+޻�iN��جL���K�.
w
��<����|R��q�YuZ��-i��]-���=a�LH
���bԍ�K���t.h�4�J��q��l+��Wg%�\�3�s}Q�C��,���9<�L��6�=�&w�l�L`���	r��IXǫ��Ĳ*dyе聥C�B�����&Ӓ�����}�F�6U�9���x��O@�}�u���:���E���i � aD )�3�.��c����=�:�P0y;��3@�#�I0(t.�K��� ~M��ё�:Q� ��.BҪ�u�3�K�t/`�1�)ڛ??�hh�D��RgSPeJe]� '�h���L����@q^�n,HPi�j�1���{{O���; ʠ\�D������mI��V�ʡ²$3;��|>��d��8)h�9~�3I>��`)�[�}����б���"���`{g��N '�-J	I����U�{}K`h�ن�|�W P��$c���O���D�u��(o|~~���5<�q��uoZ7&>I�2xAZm�/C_l&o����ϭ�v���X�C�6�਒6�4n]�S����������Й��}^��pj@�d�W���+�ڵ��{]p;ٿ[�d�Aq�X�9-���q>l���8{C����`l�`I��+�{ڂm����%U��m��e'i� 9��'94�D��'�g'��ԔX;x|>��)��`�[O|%��
��e���[��lW�/�K��u�ǑVTo�4�5�ˀ"�oy�~dw��a?B�0�qe[ܟ(�ne0�P�̻�G�x���PD(��ˋk�*s�%��f/�K��n�I�g�fv�����4M��R{�T�b�K�3Յ�)�#��X��r��e��v���2<h;���Ot����\�#�������;$�����-s�%*?ӯ�̑?�c�.` �P�r���t͒��J�]��!|��
w7e	�IeC�#9��w�}�v=�M���ᘃ#i׈�Â�?��>�}����B��?���}���8��@���W��[,��N�^h������g\������C����^�7��}�[\+�/�?��Sa��^Z��woʱAW*�|�kM�>1r ��,�ˠRo�T�9�6�L��_M8�m��q1A+)���wg�����t[n������>bhO�F��,Ok�_�Y���J�M�2u+k��d������������䉮�%>�ion6���}��J�F �M)��*J�o`P;R��!�&�>�F��'K���X�d	�(�#f�``�3l��f��v�1��6d�����X�C�8��~�!DE�ڃ7;��aH��Z�Wl��'%2U-��y����b��P��_U&�2����}1:�BsW�G��"2��ol�L#��$syr��MB#�e��E"�}���K�ķ��|������������g�c����9����=?��!���� @�Oأ_��}Ϋ�K�/hU�� 7��`ː:�y�k$����u���5�u��_�#�OXQ����x��K?0ߵF��Ak(���F ��e,1t�oVw�Lh�5T���O�ß��/�<��Cl�'�G�3؊���zE��'����F��R�L,�|�x�����q}�/=Q没��[C�ǋ��"��m����H�#Д�b��8D%��Q2���hp�Ʈ��h������E�Q�/yF�2���*�8���*	����n8u_����/�0݁h���B"��M^����w�ቿ!�'���j0�fL`�8���>��9Ì����+��MҮPV,��Pi��.��8� vv����aM�fa=��,a0���&P��$�Eq��I(��4V�L��,E���UA��ik��f��&sF��N��%7,��v���k!�����P�%�'�Q�̗{��t�L�Y�^2$��hY�@�-
�tzp��iHj�t�)�H@���Q!1�%ūᘡ�,�� �|�8����l�J���c����S��D�b��lA}<
=1���ֳE���W��5ۃz�ߛ�k��:(I<&9���,���۝XP�r�G;�d��"�2h�9���ژˠ���"���W脰�|�I�=Y���5���B/�5�� l���\�)E��5�G�:e0�A�&���ʄW�ms0�.:��'�9}BFa��%uhJ�l�Pdf	8�`g�k����� �� �IT��u�@	"2�WU �P��+�%�	�s��,�������4�
5��K���0�#��Q���M�� ����(��tt�Ew�I�e�L�#��d�u��7G�N�wk��E�M/T��S���dIy�!�:�Za֭|�2��׳��(��YC��m:O��q���wASZ������Q�k�B�Ǵ�N]�x���o��4h�]�Ыl`~�&2k��@���Hf�'G��9���K���V/ ���w�%�W��.�K���i
g��Sԗ�:�5�f<���u�M��ew_�dY���Cu�y.�_�9U�"&�Ņ�&םZ�|(X����S`@�:��
SLZv���k8c�):��٤���Lk1Ap���f}=ήedZJ���$� s�A���^-m�J� OV�G݃(�v�����d�#l�鸖�A]�q�dۇ��s4g�ɽ}�u��΄�a[)TT�40!@@_��E� ��K��b�m��4+L�eҝ:��� �J�Qb�cb�eYV��$�b �� ��9��������Y­d:�5A$4�>���G�Q��d}��ĉ]���p:Y�D{���#�����\��N�K?��V���>�@�%#����ں7^҇�򠽵	f������^���=X��u�:�P٠�I�ch��v&�rsq~�6�����5����.�O;2�Ym����m��`�fv�E��L�8ݚ:}(
����f�GlH���̟��q�Р ����8��=v�L�sb%�7�3ٛVgr�~�����+��KHg�FI�P׷�UdX�����5��K�鍝�һ�i0�	�h��~5�W��`�^_	��+vUVX��Q%��,5�R��c�T}�� ��[P~�.聦%��| �\�ua��>��@�h�I-�J��&�w������M����������B��� I���%�GgY9X�+�<������vI�#����y� ����_~��l�`�9��������
s�fP�g����&���H^�{_~�=L@J���ں?ϝ�6��]��T�I�y��έeS�]C��\�����Di���|9��6����/�3c ��_�~��ȟAq^�c�r�3�1���^}c�[�6z�+��7����˷����������><|y�9���O1������Ex�9��E?��;@ngt��Be�������y5���*����?�pG�W����)=�d����	��֛�%f;e;�ذ�頦�3Y4��h%�����~O�Z��Fvc��b�r#gY�A
���I�F��48&�$�d	h���#����j��'kۛ'}������%o���A��`4&�2��R�X��.<��8#����J����`A�h�L
��ٟ$Nm`��E��	����!�Q� �ЩU�~˘�cs~�sl����v*��(�mpe��� �5��C���
@?<܇o ��;2�p=K������4u��(�\A�́.]�L`R�����R�R�͛TʏfkE����������U��ƹ
2�D���8��TW%�\�`��9�r���,nP6�3�yG�T]<�H?�� ֏t-�u9ٜ���:	��Ϣ�;s	G�����l뒲�K23����ި�y�0Ow��{���gFR�pʶ��k!�K8�hQ�9М,��M���JT��{�%\W���4"$�� j��B�6���(��'����9_,@N��5�)�p��`�K+贰�.Z��Fӫ@v%����t��1=���m��j��3#�I?l�C(v~aڍY�z]E<��}&��Tl���*b��f�.�ʕ�߳�6H�ynĕ��v����Q�Ǿٴ��?����ڀ�w^/��Gg��[����֣�54p�3�Zbjz�^(�M��,��>g�ov���v#Yqd�:OL�8L�����6c���~�`g�8����=�U���W6�Q�ťcw~~RZt��Q{�ӳu�|��qW&><�-���S:
R�m�f<�F�a���<��]<�:�p�]p�]EoB`4Gfg�5�N�.�8��9%`^`��3?����FtL�H�Le:����ٲ�uR6�9�{�v�
������Y�0`���¾qi%g,S�"�$���$�?�Ǖ� 2��L��د�?$�oBK�@ h�z���0p���Lg��r�|M�e����<�QD`yc��N�=��s��	k�쏣|jf̳�]�l�e��� �K�4�<1����fc���=�RgۧՐde@�ؙj�0ҏ��#s��d�F'7
`wF��W�M�o��w�/H�����������=N���%��8'�Y
�#�1������f�d>y߹��dk���w�ru�"ڔk�=�M�Ji�3�Js�
P}��<�6l�	8�L�p2�0��ղ����?����'�>߽�x��ʞ����으[`�rI�F�2!z�:+e�.Ԭ�4TAx�@�FH ����(�Q�IL����ƖSc���T7&�` c����n�(�\�+p.qd�]�*��*�fu�P�v~�b���cp���%�q:7���Tw�R���(�X������"v�UO��S�~_�Z�bX,���鑭�$����zs���^��;%�/�H`�^���J�΀<R���{���W;o���� .�D�w�;�g������� ��	���G\?H0sӛ�<c.%��3���������.u4��7ļp%�����J0�g�������� ;��g�[�o�������������p�>�������STl.�X}Ӆ��l���[�jQWB��U��T\��.�o�]�%���2X8���4�ԅ�f����A1Y%ѳ0��%�v��^C�g�Je=�!���!�����7��r�E3�NS���D���何fg�x������,T��`"YPV��J���1k���=�@��b#!�3N�]p�;�š��4Jt&c�`\�p���쎪7?�	V�M�-X,��K�w�͈���K dm	.�I`�P�eٞ\�+���}����o���7�t 4-�k6<1�4ن�-yq߷�	ʒy����7�=�F�8w�%BP��Mk�6��BcXm�=T�p��1*ٙ��>vܳ��2�.���گ�����xWj���K����
6p��\ �tmw��~�Q�
C�h�+]�S0tO�z���*4���	�ٜ�X��`���N���(�n6���>�h#��� �3��1E���b�dׁ"���a=�MT��3d��#�Mㅟ7����y�yn �AQ@k0�# �?��ȝ�6�~�q-�9T`���T����t�U�
�V���lD��e =۷�R��\ �N�Ip�|�%���J�B�8���1Q��2�N��W�xia�|$go5o-{��i�����;�u�P�sp'��`�P6��=��g���-F�߫�}I��7�e������[��W6�S|��k��~���b�A�p'b����֟^:��.:P���T��ܙ��;�e���>:�E���;�����������WK����]-�����Ͽ��4�N�ipA�mc�&c�@X~�Pg���@\����ʰ�L�h��A�ٯ��X�}�h��T��`�/%�2.�.  �;ũ��˅V�
 ����X�[:rF�6�_0FI��x�'Q�×�&T�I�[c�a���%��(I�    u��`�QC�2��+�}���1�B%�6�`9����+�W�W<>��da�t氧��\@�l��{v��}�O����Jw���'!'�Kߋ���6P��d:=d�t��R�$x�&0� y0PI�	e��.[����n|���:0��+���1���1a$����X�յ� �y%v��ol����(���iG6�8h.�Li��SIV�t�a�c�IR1ו�#`�+��-Z�7b#�8U������t{:i=�������eU.0M�'���k�u�i�9�:��3}��Y���$����O��<�����c���T��Z��#��z��6K��P�%���XcjM<O��w n83Z�\��F�V�NVt3�#;��p�����2�s�s�����D_��9sDC������+v��t�Ny��Z���J�c}k2[��w�[����_�n�	Œ�jO��s��^YS�����r����3���-�ʿd{z|��Tt�N{})�k�@_���#��>χ��s8��;l�!�?k�߁s�w�(�8K��.�6�Pⅲ�O�	�4���ƚ�(���J(>��Ɣ���H�<��l ��I��2+��w&l�V�H��u��i|Cx�{͌(��*5�N�w	l �Pp��#j�<�N�K��(�{�7������;��Q�� ���](R5�EتqVX6>^��Kn>��x�i��6�m�W�*����Xy�hFڍW2A]w��8DG]#��̂m��q���t�>U�J�d�=��t���]��U�� �vƓM"M��B���ڞ��-�L��ْ���h��2��;�.�n�[{��{ӌ��9�V�;Z�n.��61�L�xr#�܄�������ڔnV��	���`P;�|Ϗ;�&{'�h��`���NV�������X�ݧ]6F���Tý��t�*�ܷ��4M��'�G����
�U��fyC[iNLu�}F9ԓ���)O�a�W��4h��ԛX��a���5<=��6��>����gG0�@�>Ek��<ʹ�j���=��e;����U�bґ
��LXz_~�J�a�	N�U�Z��1DO�[;��˗���큎�w�����IN-XH��=�������V�g6k�{#�?r�&��z d�m�}l�kB�pf9�f����1�3�b}f{�cr�U����kmZ��b�1� l`�*ة\���Ї�%+����A�2�Bk�b��������?�(F�`����-��\�%5�g�ˉ�ׂ�ZV��KC��S�м7��;�����w��#�(����d+�m��$���s�)ȝl���8��e؆ؚV��?c��J	%K����_�z��_�O�{��oG���{&��``�'�4W��-�Pg(ر�X�t�O&]lx��m��p��KOv��_@��K��=_e.��[�P6F	�
���b�ǌ&����)qJ��hI �Vµf�6�vV���g�]*��6�@M5����Y�u����jR9� �����B�n`��24B �#���������{��U�{+}Vi6���a�{TYpoZ�8)����8a�yz~��ݤK���]�!�sby���Z�z�zo(?2�
����²���.X-�\��f+��������𻘯����^�G��,�o��B�6Xȸ�ـs�
E�c��)���2�=ȎG[�|�c
rh�:x��8�T�0�I�����}������k�a�����!�1]�N�T�9�Cw'��36���O�L�����ⱉ,[T`��L̻�n.fco�B�;�Z�q`���E�7xlU�|���|Ώ[��{���X�`e��tT��D»�sQ�x�"ݰF'� f��-uNS��b�*_�����]����Ѓ��NGp�y{w��ŗ��"ʞ�"5�jWY��E�����\����[���
4���������Qb�zi�_�+�����u���A��d2 �[�C��b����	��>���3��7Щ��_S[k5�!$�nL�w�w�O������{09�%�й���.�\�\���X���r�H<�y|��)����������k����j���׿�-���_���H�|I�Ѥ�@ȹh>�2�c�1�b��P�"_w���ù�w��Uڳ�<�	�8`�u��Ҩ�������S^ܿ[��|�0��]�ae4���,J�FUS)�*��N�\�����?��b9�����%�ۏ Z-8�q'� !!h�P��Y���`��gy��M�btѬ����u+۫���yI���d͈&RgF�;�=�ͺ���	�㛴g�*�g�N��n�B����u�H�l'�����y���C�1=�x����SKZ�B@G�-�X�~z}�����}G3ĵ���Q�%f̅�
.ڋ���Uv'�;�	b��/H޳H���QjkI
z�v�N���q4�<_cr8�$ɲ�I��<���f)mw��s�\e�۩��N�D���bshʌ�|��R�ztT�,��G�٠l�./���s�y"Ci�y9��H]s���^�S��`�A@ݤ@ʪ9p����q�
G���2����j�	� 3�,a*��O��߾<�� b*��9t6{X?S�匘_����1Z*��d���af9�wt"c)�ӎ��̩���7v?];Kck�B<g0�W��#��m<�	c�L�:���Hj}>��gQ�wFk��p;�ng3�A6�|�X�Zu�tO��t���/A��}(,�";�?ܩ.�����i�ג��&@���м���=�^/�z����w���!y9����S����b������7�)C��YeGd��]o{�;Cʶv�H���� ��i���Qz���cY����b����+���pi��d,b6� 8�,�Ց�!�B
�3X2��#���(���v��줺T��:z���䏖��)�gr�c
 ћ�y��5UP��/�tM3��d��f���[��,�U:�Y��i��.�m C7ڭsf��7L��<&�z7�q�R���>G	���b��ԙ�P��%�b��<��C|��ݾB�@�zg�vj�P�Rh\YJu�8��g�hyV�X+����_�#�:'y9��j!@F{��j3�}MW� O����eE1A�1szq0��Ā���K�f2��� ��� ʏQ����̞"�L�:(i -���s��`�𞉏9�q-�q��g�FN��O�LKq$�����>*�8YE0�B�$;+�;���&��#�ap�1�u ,�襨�S�s����i��W��!e&�H6߲8X٧D�����&t!��r���L�6������8�=!�XQ!�_0U��$=�|��ں��j5��:�m.��(�N��:Lbq���J��q+�=@�� �vT�ؠ��f��g1XP��rH�?�>[g�+��Z�Xi���=g�Nt�4���jt���n������ٮi���p��Xg����,��8��������$���M��Ϗ�w���-�&��)���Յd�P�;��L�a1e����(���κ��xs{#=�y*`�l�e���I/szq��~�%|�1��jc�� ���6��+�ѯ��G�$�m�Q�"�V�3�!�$α�3_K̖K$��$���v��ZX�z������N��՗���,��Y]�Ѓ�hb�9�AiL�&����P?b��kvA"U�}���8�e�*T��y���.�?��;iv\��7"T4�0�vJs�B�\��/L�T����:(���jn����<�v|<]���ӳ�X�)��̿�B:Z�s������ˆ��f\LY߷��ʒ����b�VϮ���P%s*g�-k�Гد=���:)L�Q��kڬz}�lGbY�h��:Ɲm��p<��+�5XF�d��6¢29�}b�pL�d(8��[�v����S5��;vi|E�v�.��z���h� �;���W7w�}�	����e�4�E��	8MD�̚��.��lnn��g���M�^i����%��ge���a�=g\w���B�*]�R��Y����Z�k2 m���D`��lM>L�o��6��C�^m���|9c����Eg�9�h4���^�#���IC:�zU�	o�끛nC�Z���F�dX?�@gk�Ʊ�'3ɖtV�������E5�n]�?>=�Mp�b�`��JK��?���w v@m%�tT�)�}m>��-@r��2��2���}������j6ᢵS#��!e�6x'�`�酰����p��G��t����{��s>ʞ�`�2o����?��
Úc�n�KRH>Ce&R/%�W��:��;���ž���.��Ϥ��ܑ�����[�E�m.B�d���&����	�����-�nb	
K�˧(� �<t��x�P��s�v��v�^:Pt/��q$�{P6�zJ"ygS��
�{�)�I��T�JQҍ���V&����1�`��a��)x���ޘ�3�J>p��`e-�?0)�=<g���2Zt�bY�'?��{�`���{鞭��w=F�֖�d�$�?O�R��vǿ������,��7�XX5� `������3̰��<A�\^h���4e�\�,S���b�aJ��Y�4�'�#� ��5\Ds��Bc1�q���F�v�z��t ��!�պ�>�EM��V�7n4�1����*��AG�Hf���ɕ�Le�/e@��U�j�>��Ov^��UZԅ�NL�ap@t�K�:F��@uqE���رkf�9s�.@�
�z����zF�q�=4^��Q�E�����y��-�����V�ٽ���#�D��p��d�KT.�����x.'��R76G1�'�9�^>��t��uv��G&�c(������h{��|}(>�'f�c�ʼ}�d�<�u��������k"�ؾ�x�������c���x�R���;n��~�Yu� ���c����>����m��Wl�4��% ��� c�>��㣆Ύ��D�I7�7�P���S��x~��{�ݞ�_���V��p�Ζ5u�ގ�H����!gS¨�`���m��Pg�g�<�է�~��`)�V��3�Ye��|�85���*�Wp^\�7k9cR�����}�:��z�f�AwH�d�0�J�W��u�BZ��,M�0�d��p����֮�@�\�e���x��/^Jg�%��fƾr��ԆP3v�	h@vN��Ͼ�ǲH����ԕ�^�N� (�p1a��u8O���]g�NXR�W��eaT��0��c*N�^�^8I����Q�e�1����5\�0F7\�}S��l�8��8�z-ZM�X[xS�o5c��Pf����ݠ
2�:'MV�f�3o�.(���|�S,��sq���9�T��N5΀3�}��D�=�3�4�/�#V��t|t~C�.T����b��� 6�O�ࢷ��!��)����X�8;|��n!�kv��F�uٚL�̵*k�YS!X hUJ���.Z���V���r:ڦX֥� �!M{w��������75��n�6&^
J�4�Zy��e�W�v=�	a���_;g������4\�A�!�]
t�vz@����Ǿ#\��o�!H Ԁ���h2F�I�_�"�	Yt7���xV��D�w����I��P�i4�
m�Ԡb����})���v'm�-X���~�1ʏԼ��v6�K��u~jg��H��}�;]�6�߹�J�nf�:`?��#��;L�����+�_K��2L�vtg��Q6&�3N��J��29Me�:L���yZ��u�*�1�z���������=[���Ⱦ���W�죍�����}�U�*���T�@�����q_ ��6�5��Cp��-�P��fhc8;ۓv�	G��ڬ}�0�F���@��{��83�/������հ1({�9��|Ϝ�88 �׎`w��ʧ�gjܜN��Lvs��[Дؠ4�{>�eO ��5uS"�0ZEiX���׭�x���i>��lP�dR�Ku�\�~
>q�&4uP
]�����n���|���`��ʓQ?��@  k�$���8���Zg�S��;��y�{Z	 i)a,�;��K�7Hh�p���Yǅq�I0Mց�Qɛ���2�+�^�u�SmLV!9�[%� ���&�74����L_�cu~��#A|c)u��Ʈ��Eͷ�s��K�_�,k%Ҭ4��U��ŵ�ώ`�p��?rNy��ɵ����2��e>�X�����K�p���Z����  ϻds���%���ƚ���3a��`86�נ����W��Z"�K�*(�ڇ	�C�����	��O�	��ڌ��1/�i²��D�5�{�,�s\���Ϣ���^���l��&�oW��j����/���^ D�wtv��c%�.ųww¿��������]�!i���S��`�8a�����������o�))���6�>~wW�d`������:\��PR �,tƂ�f�`�! �(��D��'��$z�f� a��6��o��x陭	C\���/�	��_y��ki�q��u)���a]�.0���<^��zѵӘ����c�>�7�ţ�и� >fw�����n$�.o����*���7׷���.���|��y3ț�s~���p�M�-8��3��S/ʝ�R/̱3#�6�L���+/�,Ql�B��!����2�Ƀs6<���t�Gnm� ��+�3M��uش|A/J��|��މ��Y�O�ve٢D'�)�|�V�¨�r�vk������d����;�v��kc1J�&�M�F`��2����z�1�_�ɦ�6N�i�LhZ����VMe�X	
?A���E=Oxq�!V��R���%�R�>-6�����P��Gu�7���t���;t]x���Xk��D�hc�;�~���c��|�:Y�ɳ�w������C�%hl�z:ٵvd�D��0#�M��.x�S�A�+k�k�H����1������. ��`�Q�w���U�g��1z"G*��.KKϏ��:�9@J��Ńm,�����d�0S��ݼl}UA��O��G_i�rCy�D��!Z���j��EP�3	^:�l������/@�N�|;��j��F�{l��~^P�7yP�ݯ������z�e�����¡m�}����W����)�Z޺�~ݓ�4�fc���Zg�~P'6�E����ŷ/(�~��6o;w�y��>���|��}��;ox��h�<b˓uG4&0��OP�D-t2��8G%��C�s��'w��,���!;�C��'�Ű��'���٘�� ��:8���VϿ�����?�u��^۹�B�f*��$�{<l��Ǯ��T ���_Uڃr�#s��@	[�I[��x9�I˾ؕ�6�M��h�V�:���}`�ù�c�p򱰄�ʙ{�J ��O�ǰ1�D�p;68Q�U��m9Yr�Da�h�O��ȣ�'�*;��w� U�<����G�ɦ0��A����=}>���kt��!�x��/cl �(�P�P~���u�U�^�Z�$E1`�s����;l��D��Y�f�X0�ӞR��0�0n�ݖ]��}RM?:�C�8��<��օ�q���Ѓ&������J换Of�ӣt���;�U3p[뾯X��5I3K^AGr'�f L � :�'k�`�Mߘ���x�>�'!��b���(@��@G>����)\^���=
����$���C'���AL�<� ���F�7v��8�A�z&� ��L��k,�K*�b)�=�ctV�6��l#/���d �7}i�%9Si�},>R�����b�{2�.��!�lE��`	��ĥ� ��k����������s��iЧ�[�K���!^�#cZ�{[������I�M�Sew�/Q�Op��!-^���k�[�.zoɇ��h�w�=�9��W�=Y���=�X�x#�r��7w���Ĭ��c��w�n�E[�,E�̼�~����?�������u��Ͽp= �M}4H(tb��(����M7�E�ss��,��`�޾Y�F����d��j����˼��l�y�n�O?����d�Q�"J'X�di$֒*����h�۟xwmOa�c(�-!t��h��=�n��7;��O[�N�?��%Fp}��S3��L�?0\���2�^~W��p�A-�%��t�*<_!ߋ��2 [c]2̅5�ŷq��>.�<�L���+/B}�Ż�o�k&,`*����Z�0ߊ�2��)�`�MHK���z�;@�K�r��Qr��2N��:^m����)�E���/�aY���r�3&�F�BM�P�5Q,g�xF�?D	���
��l����"Xي_�3z���B����h�R�zsB�8�*ݪ�8-3Vy06�kt��6�T7�`�O�VC6�"�����(�E�~���~�1��񝠢�4�;fIK46N�{Yj���Z,���ݑ�3g�΂�io�m0x�iO��)`��LՍܝwg<�s��כU�ԙM�i�`�7���u3۪f9dR�߆`N��	f*���l� �1x��������g���r���C�8r�j$$f�ݦ�z��j�����O����"�l�	g�(g��4cu)8q�0+�'�����_Dc�� ��[9�cez��?�k���/��_��Q�2�M�;�1�M��n���ٛ��T��m�5�\�zϒ4&��!~9�s�A�b>c(bɭ=�{O*���X��h���z|WC�����i������oŽTfxJ��2�zữ�xPp�.�U�bl�o�n�_C����u�<��R��T�)�!{��q�����o�2��O����nl�[g�K��f��;�� �dE��ԧ��,�#�� �aםN��08�(0[�q AY�0:�ck��չ�Vz�i���d������\V"�66��v�l,����b7�^s@�dW[k�m�ij�#5�^��A~�[�Z�o�ղ��̧�j�A�ў�urJ-��\�g�ǖ�=��b��E��K�Y���Z'@�胳�m)Ms)���W��;'k&їD�X��i�O)���l��Y	��&�W����Te����<M�?i (zl�b���ːER���L�~<�]��v�t�rm���_Q[j�L�\5b�˂ t�f�لf�d-�K)Ywlj�{��l�.�d-�� P;�����>l.v���w_��-���ɺ��`�l�����ZA['�A�KtE=����-U�gem�W�o�k�?Xsꖅ�gcM��p{%ۓJS���d������aV6 |�����d�Ҵ	Y��۬�&�u3�)w����Z�	@g������� �P�皑�rP��~�ͨ�6v����Ƨ咗o*[e�x���l�7��g%�:�b7S��S�����KP��s�R���ɷ)6�&$��G�x=�[�V�ݻu�[r���� �E&
Ʈ"�
�c>���-�Tv[�>,�K��Z2�W�o�����A6�
%X�Wǖ�: .s�;��'Y{�y l���c>w<�f\����_�~���d�u�?y�J��ČI_�}��ђ��w���ÿ%u�þ�P�U�����l��<��V� �9�~�D4�bs�67�������s��g;cY����~_�N���c� ��:+&r�ι����M��)XM���������"��%s��jXk٪���>�0,|���5}y�C��{W��Z��Vz�U�5������M,l��!�f%l�$u���-2��Z8ϕ=����i7�K���r�c��}�&�����������la^����I�'��2�̰�\ש	*�qR+�\3�
`�L�x��mv���kf�ư�C6�d3[O�L]�,�Є��S�zn
��6C�M�뱷N1:�T��`�JW�6�Y�9�[F�H��jQ^2�g�l��|�׿�T���n"��=�-�U�w�7,��b֡u��r�6W��/���Ҭm�S_}��ꬴ� �^A���1m�k,���s����c,cW�Kq��<Z�J��2�Q	�Dq�n|���{���w�n��Q�ێ�+��{����=��fs���w/�;<���c���W�.�9|��Y�^^>ʑc����I��������������E��m��o��7��\�[׾,�oFQ{4�_̞�7�k2]@0	{K$�x�&�B��^�S�z� u�fp�jPu�ĩ�y_h�P����#���c�	��UKn%���Cp�k"�,�c�����݅��J80��dl�م�C냼|�=3Z�1\�_8[�ſ�K��f���8Uy�V��s�e;O��T��T����f�P'�Ŝg�	�z�Ud��L<����e����2����Az�۵��,������+#�w
�q"��S��c���xk�mG�L�+8;��ƥĐ�u���I|fw����3�sݾ�(���gR�g��akrӕQ�'��(��ua��ʹ�V��/��%��{�k�_c�Z�K�*��Wu��	�m��<y�!F�u�ٸ �08�.���.��sM��tT1]���{�l]��v�΁j�%3���T�hܤ&Fm7$c]����z���L(9c���Oi��-C��6�Ye sW��}��S}��D[�?����m�6������Q���������5���V�'�c 0 (�������d��k̑������/�3�`R��
�>&��G��1� ����aX���<���>P����a+���V%Z`�J,W�֙8�ب �	�\]���ׯ_�a������,�B��e~���/���Ӗko85,gKt���'%��`L=�4�&[�H~��J�l0���f�+oJD�\�jg����fݾ���π6��&��_~	7W����&|��>���c6h���i�{�Q�#Q�ֶɀ���n�K�?��?��c��o���E�_}�;j�����OS�&.3�
�[����os�g��zV/��ы�ή!�5;#�>�\s �*(5��7A�;�QP{CW���o��\���b�	�&���7�di�b"��Y#1�^��d����k�?σ;�z'fy�13�}�|�ͮjJ��'�g�̃�����@j�/� ���:�Zk!)[�%��u{�m��͋�/X^ͮ�R-�RR6�s+�y�c���=�����:<�ӊ��R��֩s;4N��{0݋��ܮ/4΀_jYͤ(NC{m��'�վ)�+gK�h��V�G{��c���〯��|o�րˎ�����)��->S�1�;x����.�o[
����/�Y��٥VJѠ�d��~�ߎ�S�����2�p��!��;N�?���`��r����
�,���4c3�_|�}ٺ�!-C�ol~_̗xk��@���2�R�4�|,�C^��߹w����7gf�'V�#+��^�N�a��^b�-ǧ8��������l�jGc�9Qt���@�2�4�gcn��A�����}�T�g}��~�^��Ӛ����*����>LrM������Sb8�֠���k��j׌9��9�����A����Fܮk�z���T-�,�����̦��7Ѱ�ݓh����R^�v��:�QBs���`H~L�Jʏ:E�+���d�㤎N�	��E�1��ĉ0/��K��T�^۷�7�H��,�/_��R(��7�4 E���\~|��NhM0���΍���C̥���$i��I/}���]�r��BR��;�^.��\�R�N�s(���������̊�r���P��澵�B��Wu�Eb�Y	�cT�O���D�������Yh��b��Gll���}���}���'����������v���+�5Y��j�Xn�f�E��$�Mt�Ck�?�ۛ[���-�:	�~���rlt�$K'?.��Xru��0��r/����2���OG��uC���R���n�H�y[�e I��fA�'�B.�ګ�oO��Ai���J��*�?1��kI�p���M�f��{7��ـS� �]��oJ�������լ�E�]�U��u��v��yͅj�bk�/;B�o���1�-����1\]\���-��~V�Z��u6׽�$�-��sO�v\��'s����<��m��+r搹̹�JF���f{6�<�X��e�����ᮙ^�p:ݮ�;�+5�|�]&r]���)N���:T�@,���N�sၮ���L��Y��=�~��+;�4ۭ�w�paBw"�&5�񹽽q��\+/�8�b��xh�̍�� ��)מ����h�*�x��l4^:f1D?��$'��g+q�Ͷ:T>f��x*No�{X￾�,��r����_�QHe�k:ҝ�vN/��\^���_�O-�쎬;]*���Tɜ��t��/,�����J�dH�ژ�+i����X�]�.^Cs���!C�:#Ni�OX@2�ά��L
�5�h���}�I�r�
D�����<�u�m.i�J[v�3u\�2�:��<W��|+0�L�ZBWʊݏ�R��~��������$_������7;x�w� k����P�lw�pOL'����΄W]K#��������oX����?��֭y��M�?;�^b��5��>^vi��^|�&n��r���n�Z�q �Ef��y��/>_� h��������z��=J��o���=Ȧ�v����2�g�.f�^k�ɍB�6=��e6�]s�o�6��CP��$�5�M�-b��T��ߤq4��w*�3/3�=0��FG�2d�mm��B�/���-�S����B6犿�����C��Z+>HWW���n��&Ra:y�ic-�9� �uΔ�nc�sj�ŋ�D	'/'�;o�l�i}����{:c��Л��e�b����?��Y�����3�� ���r3��Ɋ�[~��|j� 6�ۖ���bS��CG4p>������E�ރ�/�lƣ`,1{|Ѕũ��h�b�GcL�$�iΥ�G*@�sȵ3�s��^�-���[S��b�uZ[��3	�2���+n/�|Uv�<�~������d`��b���T�6���v�4��j8�v��׽J|�y����>\t}�(j�Ji��M���Tƥ 4:����/��Y$SpMl7��l��1O��ָ�l�����#���#;��6}��1L7�! �9%
Fχ1tSd~�4�l���5�%!��8���ǰ�֡�i��!4O�l�M_��1��ܬ�G*�Sx�����������sخ���r�.����m~������Fo�����)/-k\�9�'���?����Mx�Gz��v�t��!�c^��噴G=w��x�X�5d�.���[��qjί����	�>��A��Q�Ϧ�+��1���1�_bq�d�i����8/E�)j�ƙƱyOjv?��~nM�gZ��V�g�v;�iS�������?_d�cXP�q�9doh�����pc=��S <����L��n�F�Hu=�����Qx��ܝ�˭x�X���M(���-���Q�]F�A���W���������:������2G�� t�����Ks)�k��5�N[��8I��6�ȵҬ�vRs��c^�Z|'���-c����~�Q��hk�=&c�4��08����}�Kn��Yf5�}6�����[�b���_<��<˭�:*���.����9�G����	?x��{�-��g�[Ϯ���V�@��΋��;�أ5E1�;b~��zbxa:J6���~�.�OX�]�7M?�oz��"+����>���T���g� ��{��ץ�ړ���R���g�e{ Z�j�5ݖh�;`gq=�%7~�7׏��w�B���4�ڭ]������J0kk�Sv��+������&x=��Z�ӷq[S��W`'��܃� 4]�W<��y3�P�9��qe�S�?����X�� �Σf�7�I
���N��ƌ���C�e����&���͡�q(���E�/��y��6��T�X�������?��"x픉�����F�f����d�O��y5�]�e����;��᫲ھW�F��de���ŵ&�G�9;R��'���v-*_e��3�b�7��a�~X��cs��G���ml�*���-�����u�����3��U��)�o�iE뼋�����_��?��au8��	�wv]��ʞ�����V�^,�#���tT5��Jy�P�5zWL���qs�	q��.�8�� ܀��ԝ�p�S����1<m�(�]%#�:_9]�~��P���~�..Y���~7�v�0�v�,�������|	��-ޯV<��I�.L�}m�Q��K{���~އߎb��R6<��ak�F��{�f)�b�@E�C�R�-��
5o��<���)��܅�돼 (͏�!L�!�e8M+�\7�C2Eꔪv��}���H����m{�}� ��͸e"�+v�ܷ��P;�����h7�����x�2����Ȼ��Q;�R�u�%��:�'/��ܙ�S2!Y�5;^��P7�h@�\�v[�L���ה�k��<�����I7�W���Ek{��ٺ������|yV���bw��Zr���g��W�����&�:k4BwZ����*r��1�4���
��T����|�<����LiE�p��v�rD|~�d����Q�rG�@lsȥ�`+f�J�yw.|�� >鼢��8H^��6��y;a1G�܊�@Ua�إj,�%�w�>��&�=��F�.A u)�-��f���h�}c�6��� Y25�UD �YE���Ew��*�����d��J�PZ�����������ҥ��0ŕt7^�G�x�]G�����w4C����6��y�5'�Z�=2}���jC���9
�mq�����Fi1�.���~�be�G����P�4O�yLO�QrFD0���������}�V�"�4|5�US>xD<w�.�^Ό��ӯ���'�|R�r�=s�N�ܝ�ٺ�Jy�gQnZ1HtfR�}	��{��^��<C��F��a���o��R�����7Ѯ�$ia����Y���w|��"���O��q�m���Ǡ��^"�e=�\�m{݄Ӯ��K
@��T�q�a~$�\����O�~b��x�Z>˾�:zN�d��z����^�eQ�4{�9�qTl[�w���v!y��
}o��e\���oT�y��\n��7��Y��E�B��7��Y���۩P�·�yϨa�'�#�(�rN)h���̫�|7Qy�ӡ�&��SJh��kmq�aad�O�hMW��٣��l��������{t9%�>E)�;œ��Hr����&���zM���6{z�$ԓEf����h�``g��D��V�5�BT�nI����x�n�;���<QVЍ�V�z~y��nM�Ö���Ġ/��=ɕ��x<FIa�hh'�W��?�H׫L �&\!s"y��~�\��o��ww��^�߹���b���2EC��1��A���}q��*� ������C�s�d��̑_j2���ꌭ���|WS�E�S|�Ɇ0a9ʜs���q�#j)�sFȐ�>C��Eȧ�� 	�ޒ�{�{$Q�1�L������y�gő��7�]�
&{!�� D(�y�$�~�?':C�MzV�)B�~\<���5r�wC�.�J����;�����@!�t�S^�6n<��a.��b��}�J8m�u&P�g�#�)���"��l`C1Ƀ�	.�[ ��*ۖ�X�s�҅T�X8L��4}G�rY� V��T����7��Y�Z�$��}�_6�������ڿ��02��0|�X��>�ު ���t�. ��'�a��x�h([j�@v9t� �u?�6_��er�k���*�so���^�
�'|/S�S�V�P=fl�ȿ�[��\�~:��"��K�4z����~]ă�^�P�c�ה�OV|B��K!p�}%��/�h���/0�K�/{����Yp�}�����(=��Q��/i�n�B�%�"��W�u��G(>��F��P.������j�:��!�|�Go,�1��,�\xU��\�;N����7�����^ص�r���NW�i[�W��y���m���qI����r0B��끌z�?��d���ә��־SZ������w���������2�'C��T��{kbyQ�o���w���*���d!Vs�4�*ӊ�����]����"B��8'R)w���P���r(�xH����K-ܧ��T�po���$�<I5<�6V���g��oك�*��g4(ڽ֖���X�s��ϧB�}�kY����rL1�,ǘ��%�Ӆ�tcd�����F^|L3��q��y��R��w�rK)���E�����s��Dq]&�n0��b�����}��P�D����� W~��z~x��tNW�%��K�^�����9OOO��f��P�j#<�YH�}s{�	�����ߧ�[�t\]]�
��V+n'����H����D����ẃs����Ż�cH)O83 ������=�� t�ה����;��$� � 
a�-�W��A�ȃ|DxplT��$�g��C^Nqq�i��+"Q}�\=(�S�i/k�S:�%��P:{-w���=��?�� 9Y�¡@�1Vv[�j������E��.R�t�2�*w�&Gܶ"M���`���C�M��a�^����⏚�� �[�=]��,�^΁bV{��� 8��Be�ȗ�(�>�[���#gj����9��ޯV��L�<�FZ	��������O,�W)�d��>�B�#��CΉS��c'�$�.���w���G�.�4��R� �:Ԟ�� [�U�r��ȱR���T� ޿,�����K�ǺK�fw�BO�b�Ld��������f�s��uջ��>*ex�Gѯb�ǭ]k5&%��S��<����V$��x�XI�~.��wc.�}8Z�$c�*"W�%Ya(��*�>�顠2 r�*�h�7� �ѢV��
~@Zʾ��	���NT��5�e&j{/�W��7��g�O�t1[�n�0`5ڎ��B�+���H�A7Lڒy��0UKԀ
�^$�#�ʵl��Ź��W�t�����*{-e�k(����M&`Z������2>��k�0��7S��^Ɔe�.��p��x��N�ca:}�.�:�	�<��x���q^R^i{/'t>�b�h�/�lE瘟��fi���*���ڮf��K#u��3@dl�b5b��sc��p~��0�{-���N�����P�1�F���N����)dUt�\O�BcF�9.��̺����Y��<*Txl�s����U�Z���kyФR�� 嬸6lѷ��6�,#��u5�ͯ����q}�D���ΐ�,�W�gN `T{c���1>o��Sok��h�h��	�%�O�&O��y�ٱ)ƾ�?�&��T �Ç��){Ud�8h�$�檬a��������[�����E���]�ey���1�g��;�{���6�1�/{:��}��}T=ǉa�u�o��?�K;Nn-ˣ�ſ��3WuE��w7����;���D�����v��9�j��l�����K���juE˫%��k�{�@��������? w��9�V^P0#lZ:�5�G�4$[�����4^6H�U>C�w/���LZZ�%I2@!��<�M"�wӃO��#N��N�3Z���lA��>|ǞG�8l�t؋��7[,P2���q�
%,V�����OҤ���C ��I1��X�U�N�'��{��&������N��Dm�СfBsM��=<wZ!\��8�A�4�]��aJ�\?ju8�ֱZ 8����*�e�b܌��k�����0-��w�E��J�*�V�u��qr�֡�����R�+����F��7�&�opݧ�S�d��S�$��[ȭ�Bݘ��g�t��T>� |�D�7y�QE_f˶T˲�-�®M��}��΀�z���P������d���2���7������5ʀ��dώ��g�,�@0Xrei��b�](.n��p��8��mI�;T?�׊ba̸+��u{�+�w��OW]�&�=>@d"3��^�-��>���1���0Tל '�G~�%�T��	7����Xܯ q���<d �	�R^���2�8�]�e�Ǧ���r��.��U7ʕ��s�-uP_�6����j�����-��+�a���7�=�_{��aK���B�ol�?^����18z_�p���ڄ�R�q����^ח^Q����ʗ�SxB+������k��N����n�P>�m�֟����R�򜔯=�����$ꌡ�rʂjQ���hEA�l��׺}����!��J.3���e[N���kB-{�}���8� �<��e,����Zڷh�����r����;�o5#�5Fm�ȩpS��g�x߇cZ�h[�C�����3�k�O[#ŋ�~��wc}�+�QyU����!����� �������g�r�'^�Se����{�b>cy"�����\3���Mi�̼��Ӭ��\7*/r^�G�ws.p'w 	0�9�9sPn���O�Y�>�l�r���r��/��t6�5=�5�����%�,!
h���`α�����sw�ޱ��~�s�� 2�>����4(�*PD�L��{���4��I�[�L��1�q�sZ�0J�Cx�a�֜�F�^��X�+R�!�� �0N������?�]G��)�$խ��/�:�Os�8��,;y�Qk*Ǜ�A�G������A��4��i�&��H�DR~�FĘ��[���w��0�/������1���D�0�Ά�wP�j�H�#i�Ac�����1Be�:f��`��ʶgy$�23��
�*�]�k��ï�l�|�F˃K���[&#o�sW�r��(�]_frϖ;�TB�&�	�\gp��P�%ǉ!��=�:�Ϝ����s�~��1�J�Y��L�m�5 dO�Pf�CP����h���Q_�J��,�?!P�5�k���}�n����9&��M�B�.�X6כ}Jj1�$��`~%����E�L��%�O���:��;����uH�,:��,�s晤<�S��1�3�8~n���G[uW.��ą�v������Yკd/)�n6^�?�~[g�	��9��Oo
�k=���K!�r�~����w3 hH�%�t-��|�������e����2���������[�`("_q�x�Ċ�8�Z�ONĚ��dĖX�p�:�H9{Cն��⥾�[x��\�.��N�w��Px�4��H���p�U��x�<���Wu5\� �|��vkf�A6���ٯ�p�y��w?����._��<8���0/�����M_�E���ȼ�sVrb�a��������g�G��(�b݆|I�E�����(B��-a�� �l���rIWW7tu}�iZ�C����kZ���p<v�er}u� J���^s�r��i9D����޽�>�iu�b��+c�G �����O��A��~K?��r�`���L���c`[��0H�T���p���;{�L'��I���9��}c@@!�i^���f�^C�傦�)�:�V�*b����N�s��������6	��ң8"�1
쌊XTn-)����-�^�m��7h�-��(�-�:2*��q����LG!�f�E[��f~�˅�;.W(�:7D�"��w��ߙK�	�/��/�,�s���,��k,bysN�������'煰<gu��߂t7�x�׼���~e4�]q��)����A��к#�J6�@���!����m��]U��m�|rà�5���g�����h�4*�
��լ=Ѫ��5�U�d����揈���ח$G�a��_���ڈ�#�[�q1?���s�+,��\�>C���~�	?_Om3�V�j�]98��W�F�y��R����R8�����`������g������?��L���̺�z��!�k�w�_{�K���L����:9�[W��^���a|_��w��]��|%v���Ev��7�䂲�%_�Q��U�/=8~���R��W���L�H��4c��yy���@�����y���Wa1{��|_ѪX���Է�������1zz�'rI���gpSᵝ���_2��Q��J?ټÿG����o���@�{���r���B�i^i�1���L?p��\Ծu᫒[��-��%�Y�j �����\0�˒�U�T�?d�sSP���i3�B�.��V�Txz��=����C���Ϗ��@�0�y;����G6�s��ٜ&����V��g�J���rI�7�t}}͹t�ͳ�nh���J�\y{>��jyE�Ŝ��\ʈ���8�����/���}zz���g���m9����Ҳ�J���v\������n� �o?���3�:�����a�|�d��I������������%�E�>�6'�yy�*V>����� aSGQ�2����.}ڦ���s��b,�pb��ubj����`ʑq�3?!Rxu��G�>�Г���J��?F�*�x����v,h������P��Gz�֝t$���U����nr��������Q�c���q/�v��0<�j�%ץ���P �j�8~h�-�L��p�\x�q	#�D>þ>e-�U�o%ǥ�n{XAKl�ݝe ��KE�K�7�
���~���~p-���б���}K�G6��(jf�k�b0`�Y1%G�ы�z���	#ߌp�_ _8�i�rj��	�S
ҥ�2��Ͼ|F�v�~K�����yN@����	�c�����7�{h�e�D��ѪS���7FyI������q4o����U��_>�Ic���~m�Tww��W�l��L��a��J3ܷr��j;=����+��R�0~~�P��8C����_k�%S^]����-��,�\��ڳ�����/:�����+�kw��ap���g����o���s#�{��9.o�5&)�9��vL�<ft�J>Sʥ�� }������1��O�g��E�_e>V�x8��F�ʡ�&W?M��_�?�k�����3�?��Ѯy:�Z���������I7�kZ�W��������h��ˆ��-�����w���Ռ�����[�ٔeh�(H��R�-�ᆓ/�o8 �������H��x��owlLEhV ��3ϧ��D�k���o?�L������mj7���&��A�<x-�����-�|xO�O���_�����{���"�?�",�I�g�ئ1z\?���a`�A�t@�P�xI��x3�3z���Wn��]�U����Z'��ܥܮ����4������2���f_e��ľa��MX=�>!����e���C��֩���I�U�DA�k����G!zА�*ǫ �oj��� ���y���*����[GE~ׅ``Bӂ]_�Ig_�e��Z�@���w�l��[�ǁ�1��<?�s�y��RvȽ�Jgs2Q<~ve�n
$g٘/ד��R(^����c�sʞ_,���C��L�GN���Ǐfm�#�E��G��XN�j�HY(���&���OЫ�������O!:F��N�u��-���:]��J@*��i�^�������)��_��J6�K
�庴��Fǣ�I�P������1l�J��*v����NN���v[�}
F冂��^����P��_�`n���_}�c�c��k��U�-��8	8ǸG�U�r6G���v�������\mc׽�̱��B����9y�n�E�}ӍE�FZ�F�/e֒���K<�he=��<Y�u��^1}��j������th�N)��X�\#��di��΅�U�_'�.N��g	ܸ���ڿ��Py�?��0��8����s�����}w���_����W�z��3=���U���MHNׁ)СɌh����}�%�����ꊁ3z�Й�R�����v��T��NZ���"-�}��4}��J(W[�!p/B�����B�>}��fM�͆f�9�zY�,�4�ł^��9/�.�aw�qb�ǗgzZ����9{�sg��8����7���a{��aC�ɒz8�Rȡgp�D��d���x�-c��F"�e�@��:�:�'KhO��Sw@Vj<wZ<�wf���a��_�܎v��Tx�5��q��tY.�f�h��ms"�t���\"�����;��.=�tAƘ	i)I\T���͞�:@�76f�4J�M�y�\���:�S�6�6T/���������J?�7m�氶�5j��M��c_�pfdz����b��V6�+�W�T���?����Ԙ��3g����O��cB����EI��m�����J�=ɘ�z���
����������s��`_��AƊ{8���������TZ�J�B���C���6�{U�*^���8�ة�����z�����k�)�t�x���Q����M}�w��G��︀3�<�
{.�K����u?0]�s�}�#��{4b�PЮ�M����U��t�=�c%h�z:��g[^2y�<�;.���QY�z��&f�v6{>�︿�a^��7�g���{��pr���Y�������k��kǥ�`�z0��_iZ�Ď�G��җ�a)O�܎z��c<=��QR~��W�b2G������9�����OE<��{lY�<,08����C'��Rw��K�&7�F_�O�հ�kJ�����0�����U��{���e:�q�����}Omh�����y�4x� �鈊�ݑ�WW��g�۲�̔�7MzX���=v&��=�ݞ�{C!�����,V�<�h�Oi�}��ˎ�pƂ啒y��3���������E׷7t�������n�n�o��o�������������̐'��ܡ3��9��\�WC�]�����[$p֐2L7�ݡY����u�֮3��S��}�dE�$Q�E���+6g(�/����{������9��X4��>�ӗE^���e���n��#������!�G@��'�dQe�氬�#�ŗ�cˀ�<>y48���p��iY�8��s: ���f�(_n�M̄�J�0�s��^��&���Щ�,�e���ZLs�ƭ�Ÿq;�:�W�k���T������6���';��y�xI,۫��O_���iC�֌�)�G_б��M��%S�����E��\Һvt��hI�C�>Y79L�T���=\XK|����
���,'	��B,�����J_��w=m�˷�NX���fZ[έ5zp��T���`x�/OԁxN�C��z���HU�t��3�t�.���b�����uox_��e9̼h,眞5���N5Ge���g��1zM,샡~G��.���֣����'��F8������r�����_Q�Q�k�������G�,�وj�|�s�睟&[4#�7�CI�_;n*ƣxD�V��1ђ(f:Y*7N�y��*�XƎ̧u����H���A�Ǫq ��\�~{X�"�/x�����/��������3M.s�1�Q���痡��F (R��`Ȉ�����}�`M�A�D\��Q��k��[��j������`\'�B-�� mL�-��� �x�Z)圐�t�/��uq/�M��
��k*�km?Q��|�d�|"��d�	�O��|Z��k��9���3�S�0F��䕾��r�i����*?�5.R(�~0/�4��`9]�q���L���g�
���������|��%*)�\|���9!�u��/p��#�|QҾ�4�dmx� ,j=[�r�`@�-H�<k'��l��3���AT�J�!��r��$�h��r���3��<�I��Kոf�^ C�ق6�91F� NE?�h3=c��0�c�!^pB�B'�`�,�mɉ���z��=�O����6�k�g���"��N4j�����	u�.\�r��:�s|(�񊖆�����e��jFM d7�L��O���� #Q��ߜ�C\�vB��<M̜�)j�w�Qb�~�,�x�I��}[��A��tɎ�3��@�L����=쫏X��_��;%��pЖ#�L<D*�҈b�D*E���-,g�T1Yh2>�W��w�d:cQt����J�����Fmk���G�'J q����P?�/��Bϫ�>&�{,��^�s�B����-�3<i�3�bR�_��O5WFs��}_�J��\-&}��=�(#@�#Ƽ�~� �z��j=�U�/J�!4��Q ����쑂��w��i��}Z %��0*m{Yk2��g���&�I��������8fhN~ݒy0Gm&L��V*+tGI�B�r���:�{�4��Q�����u?�|K實P裖y��ތ�?��{�»	*`7�.z�"��
$�l~���<?eB�z�Q�It�iMT�P������7�q�v�
���z�1��LxC8�٣��|�J�ă�<n�z��l7��� �¹=��l�UR @�D1Þ��C��J�z��=ln��k꤃����SǕA��l]��L��ڳ�cv�����oX����`�N���g�R~��}����颿Hަ�eZ(D����w�GX�3��x������9���oӷ?�~��y��a�t4���[��$�X�M[��^��k��x<\�L�H9��)�����*�H~������cεԵ$��T._R�r�e�AFN�z}��
Q��`ȳ���ȁR�W�Hz���U�Jq��JC�N�u�~�*4��Y�Өa�.]p��D}՗,oIU��f�lr[�2X�{U�a��"d��bM�C��Wp��vTY�	M�2�bd��
��j��kt��}.k2guη-��TXu�R����F�D]�<��:�1�8�.�6Y��D��������&���\`[�\�v�^��f��q���s�s���[l����L��F&�z���*3�F9>.���"�"?�R7*��h�_����ƫN��G�:����k���<��\V|�8÷���>�sf����5=<<Я��J�݁�/[
�f��V�{��6��3@yaN�t�~���x�����p8��j�_t&t�=�fSId�ɋ�[NҞ���v*	�g3z��66E�I"o���2J�|�h����C����^B�S������ѻwwtww�^=�͎P�{�t\��]!o�|��c:,'�f��NP��&jt��=��n�s��h�|S��M4�8����UVݨ���Q�!�Q擵�r�+M��1��炦7�{:��|1e���� M��Ū�
��*ſ�ߞ�tʴ3#�P�G���G&��æ9�!¡	��Ɍ���6	wu�@�
�d������)1Q�+���I}��]!%�@(��3�T�� k�̗��L��Ɏ
7�K�j�+�6�=��ѨB�KQG't.P{��bF{�DBp=L����}t�!��U%� 3�~"M1�Q�[ж3&
@�����"���#�袂PPpB��Mg��SPkUv�m�x`|�zE����f��d�{�;�ېg�v�����R
t�81�!��b�P!Y��O�_���Ͽ����ļz�GdA�	B$� ��X�����72��{�H��̻3� Wnc[��z5* �b=� 
�'ay��[��>�7���-�f�m3~��3r����d�Dy/�+�{��K'�Š�3"���|lt[a~L!�;�d��r벥.�������MQ���N�P���&������Bm���Onbh,A��uY ��;\k޷�\�74OU��r<ƎAۭ�՘�Q�4�5hF�o
/ۘ??��l�n-DWDe���a�;ɝ���hm~��k�l������.�|w���Q�y��%oW��1x�c�a R�h�:��o�u�a��ط��T%�& ���g�~��h,YPf^�	O���������j`c^��al�����4�y�,�s �u�4ZE�i ��̐=�P�PxT��l�8�8޶TPUo�T�$w��N�ɴݔN_ޗj�}��ї4G���@��q6i���-�$�JK=�D��W�m�hԋ�gF��d?��-�x�l ���~�71���������d�F����@~t�.��ظr�F��z��*��?t0
�h_}_(��f�x��s2�0�Ǯ
�O���R�0zi����J,�>�|�[c�����C*��A;�E��1Is��|��Ӟ�F�Α5esK,Wwd���
�'�wY���G���� ���~��jW���3�ǧ�'N�<��i�>�o�n߱�4_-�by����h�~�m�q^�k����6���Ah�{����ދ�6�͆? ���9{����9�5�C+��� M��0�|>���/������ҏ�� �Nm[Ηt����������:^���iJZ�@+r}4G�a��yā�Q�_��(��?�'D����W�8�T�gD����q_گE�F��֗��d ¹�F����_pT��Җ���3A|�"e���pkZ��o�Wtu}C�*����9}^�2�w�T��*}�-{\A�B"*�t��ڶS�h�i���sb^@�F����v|?�k���N�"}�)�6>8Y��BC��"�F�$���W���0��`��B@�!v�ݢ��$p�Y���>����2~�N@�����R-D��#a�e��r<�x\8fu:����6�5����M���� u�O�$O�������H����/�@a���{{UuϙX���$�
֣�Y��,D����D����m��X��ЅqR!�a^�������.�}Ѧ�̑��&,Y��r�D^S�,_O��y�k��a�0���@Ξ���,���X��oX�bf��HLQaX�1�i���'�sW'_C2��e���N��� �̭X��F �\d�ȮXK��H�݊��٨��Ls�uG�F���a�����rK��A�E���e�Y��	����� ":��ϰ���&Pz�X��2�s`���6�n���4i��߱;��p��C����A`\�mV><�wY����ҕ]�߼2��&]���Vј,��G�m���)�����j��o*GP���zޟ��áSB�L�?(
����ɀ�xO�0�72�����9��o�"��{X��Ǌ��A�N�{�=r;V8��'�~�CX�'��7O2O�!^�M�FF"nk���)�b�ɟ�Qx� �b�k�:Q.�/I1�ԫ䘞���ȼ���4���;'0G�)��4�(*c���u�{Q:|Ϟ�1T:�]�J��u^{T��?jr57,U���������BP��x@�c�6�\�v���6,�u<�:j��^��|�X�/�k%��x/+�*7��U����ju=(x��'���U���c��7���>d�_�RZdn]�X�h�w^L77��������T��ĳJgyݹܪ�^Ǆ��;�^i���$�_%Y�*�%�-A���G�J6�u�Cs�g����i6O���A_�b��ޞ5��`��H�y����>�s(�|��۫��������������ݾc����I��-�������ӧ���|M�������E_Mh��z�W=[{���}��H?��w�t{�>�[.y�c��q+���P/!h)�H�w�ȡ��7O/,g!���������2��8���!����{z||�Y+������a"�M��V��=eD�98��(ߵ��%�;�} �5�Y~N�m�'��3�36��&^,7�[T��0�=h�)n.d�Rm�����G�;�w�|Sˆ�}3�]��Fg�/�g���"�%��@�A�I������\���w$��=M'ba�g�G% x鑄׃����D�%�B2*af���fIy�?hr٦b���T��+��G�!��@+��f��k��l�E���OQ���`��7��p��N"� D� H�a�&��.�q�Z�`xXG���ج�JƠ�Ag�6͏$����x��eM[R̻:Wc���Ez��z%��%L�:J,Y'��s��)#-BR��z�@@�{:���X$bzs{�g�٥vw��u��'�X��
k`ҝ(�m��>&\@ ���7�+P4�A�(�)���5Ԉ �"�X��;;�2s��³ׁſ��9���3;m#�e��Q=k�4W��S�v;)+(J��ޫ�,���#��0�g0*���L¤E�!7춭:vO*|J+<rLl�~
�#�+	g�����¿D�A<o�MW|w�.(߷_�ľ��-��8*�8[V�+s2p]��
M4��G��h��^8���@��0*֨�*&\	;5�@Ka5t�<�U�3�gA�g`w�1��Q��Q��6�_s�X$G�����������ʗ�����LS�)�5�|ߘ�D�7i��X-R*�����R�7{^n:�2B��@�[�q�����{hU�E7��i0$ė������yf60�u�]����a�G�k��9l�h@��`�I�7�D������ ����S%��XQ|g咃�]��Jy��Ԥ�!C:&}�;�O��r��Q�.�9Q/�!빓cf�i.���^�͌m���Fu���k�ڤ�!�i(�,�7�Z�I�]�T��n���>�g�=O��4���Z��d�ee�z��տT^���	�
���Hxg�x\Y���ɺFΫX|o���o4���W)8�Vz��J��Q�^�j�I�1�͡�r0��0��!t�N��n�͗�L_��]��jU�4zQHr�t���*�r�n�t�9��>��;0���-؇b䛈�҈+�-�Wm�cFy��J��0���a�t8�q��`�z��P���6}^���$c��{�C`!�=2��և-��pO��3��g-ui|���;�~�/�7����೔�k:�o�;zxy���~>t*Nq�h����p�s5��\��q;v޿{O?����/�m�{�{pvIo���G���_����=���y?O}��ӈ{����>ǲ�kEC�����c`܄(wʅ���dgT1R�<T�w�FJZ��o��~�)��Z������O9$m#��Soi%Մ(�7�|m��<'�t�[<d��iQ,҂�f����ݰ�sS(��O�g���n}�'�D�ł�2���j�.q��<x�,l,����T�%�� yu�Xp'�.[���3Hg��z��=���U��̵��" �*��j�bW=(�8#	b��P���O|��UD5�pf���2��j��LB�'L`�y?���^�>���[�gK�l>aP	��r�d���n ��^���{ɵ��p�̈́�n���_�匟-�"��c�L!\]/i�XH�#@����ꅱ�M�|1Ӵ>V� k�e�B���s��Gf��W�&�4���/hc�������pd`瘈��͑L�n���yΦ�L#�(8.�pF��J�a�$Cy��ApϽT(���N"�`� �\��=���1]��V�~{��4���f	� �����AȎ$N�Q����g�����wy^V~T��E�W��>�"��d*�e�Efݑ0ʝX�Z�z�$�$Sa�l}�|}tڅT��ea��=�"���Pp���&�Sl,GD8��bj%�^���+��([Q!�E�>fY@+�����|UU��O��l]� �=Or8��CA�=@ɉ�s��wr�|
 5mS���%�y�g�N�B:���j8)瑹�����n��@�ʽ�fa�k+.^�vW�����A�ߕ�)F��l;�k�YI�<�s��0ًw/h�d��O�ye�u��@#`��Ԋ"�����U�	���S�����C@�q ��#Ѿ�Dɽ�g�2a����l5W�3a�-��r����N���^(Qý�ҫ,.�k�RjX��m���%fUO�
m�n��1lY��}���9#�*�:�� #�������t&A�X��@[�|˽�(:`ߨdF���kH�mT�����ex��-<_����J`�����u���p���U�o�V�)�eKm_����|9j�jD`dQ�h�S��-��s>���z	��M�k$���E��Y�����>͝d|MAx���Kus�~(k*IRfE~���g�ltmi0c:��w�����R�7V��|�F�rέ��Wp�c2��], sR�z���g�t�%�L'�]���{z��L�$��5423�91o;�c����?��$�L���'L�'�u)뚁�ny�ϳ{����Y�Sb'�r=aG�I2���)��/�%�^������&�:��� �~{�D�$紋)qo����}�_�?�.���ֻ�x:I�LM)K���s ���m��h/� |���(����;��ܜ�mOO�/������O�?�p��EO8�"-,<��0��G_�r�ӞdG��#|�vk�(���Iy��:.� �ѯ2�9���#�]^	,�	߲Y
�Ae�b�Č�vay�M�gBV 9 V<���=}�I���b�zd@V��39+-Jlv�{��{{M������-�}wCA=�yy~f0������bS.V B������K�a��ؒ���0��v�a[�C�҈b>���A��K�91j���$���B!�����%!�7	\�Pv`�j����l�e�^����9g���t��~x:T����YS�~T�E����Od9�  -��\]]q��n¸?==�w\xw�-�#�K��L�6K����5�̐�Q�	QŻnҵ�/^���)3��H�Pk6`���U��h+�pOdA���<���v�j�l��Fn�3�I�?�+�Bw[q��� V�t��_����V׌�7���5�(�euuͿc<������������})��l*�� <s2���(��7�kΩ�|
��Χi~ox����zU ���T=`l�;��		�G���ߊыK;���0.��X�ԇ]�	�� ��t�c2�+�m�����n�y� �#!<��rk��2DE}���#��pf�c�Q!^���h���ny�`R�؆ �I��|��R�����Mi!	zm��JL,l�<�k@���I��O���Lii4n�e��+L���� pL��ջ�}�<)�s�@�t���O�+ߛ���o9enmrEɍ�Cٻ��x��{���V���{�����'�ۺݦ_��A��	6�PT^+�7{�w��q��1�o��$��qeٕ�]��pBJ������(!��������{K�Q89���,�z_��7�R�S�2e�]��li�UN����@Rx\Di��X�.#�p*�lI$��׹�3��Wp�y-���A���@��-�)�m�> G�s8Өq@]d�$�+:��A}^m��E蚠��*�X1p�����<�b$Q#�n�}aeV=��v	�o�k6v��FW��$��S\�Rx��U�u)�fb��y'�-N�����2��Mב�9�5JaH�f��*����1��s�W���Q��<��׍�7���c���� ��pr>��NMM�0@��1�Hs�qV<�A ٰI2;��!�h�y�����'@[%�cņ����5��1���s���\"@�����n,0��B=}�a�n��dܼc9rD6�*��O{|�n����'���;9	g�z�~��qK��$Q��t)�5�|~��W�+���xO��X��<�� �<<>pD	r��Ж�<��.=��IGEN�� '�L��/级�<���!��3<�����O��I���ᙦ�z� �K�4�C�5<#��$[|J��֢������`.ޖ<yx��bA|�,��6՛�޸�L�t�&O���mc�����6��P�{��bͮ76�����~���j�؂ ;PT��j �fI����r � X��^<�a nh�7���`���E���3g4gUg�1�f"4TgΛ���(�_8F\CF @)8�L�
\W�.-8[2Vb�P�%�#7@\û$��(H-w�iL����&�	%���Kb�-�K����>���a:�< ��7P���_߬�8�rR/���*)~z�vw�9y"�^�e-�v�HmX�~"Q�?Oc�����	\3AC m��w ��M�6�=��">�Z�4�x���{�@T�!���t�����KP����������;b%P F�HG���':�.��Ԭ�X��M )���͒�{"�s�O�>|'`�|�e��{k���e��W�5t�B�޽���J��<n\����8��)��'Fӱ/��!����r:����ql�X
1 am@���������ߦ���53�w��&���u�y\�[Z?7��"�Wք��u&<�Y��V���.Ә���ᵀ=,%$�li^�:�9u�P����������<\(�&�]�p�F�*Mxo���Y���MכK���:�j�=ߪ���Y�L��"H��^��W���Z��^�p�aE�`�o��#C���V�o>���?�Cz�<iHm+��o^�IokFm�)d�����8���#Ϫ	� ����4�X� �"LT�H�y&�+��L,MƮ(&'������Ge�+I����A��bt�xG���*XBg��s�	���������jpn�<��B��.���L�7�y��f�9�!��Ъ�b�Z8a'�Ys;t��p�0��K��0@&��/��&���1�c�}���|�F�E��ܐg��ah�y�0�%�R�P�(e�s1	5V�� �u�ϳ�W�dP����C��d�YF9�<��K0�JL�F^A�'W�ëtcp���s�1.Q�/��	�%Մ��0y�5��W��s�J<]��f���T%0��=�J�&��!6��]��˕��� ҿ��>i�<�S���C��t֋mG�ozt`�	t�)�g��1v�T��������������vE�>�џ��g���ʲ0�������o��L�>�Jk�<�w,�b]N�2h��E>+���0/GKs �Ҫ~I,DK@�cs���_�}��$U�8�ꌯ��xO���{������@k?2�|p+�QD���_��XTԺ��.��k�r�퓬-�zy8O{�1�)�
&s���"OQz��gI�Jz��e�:����>}�ǧ��y����)龟�U�@�㒽+����󖛊4�S�v<lR����AiW��VLE�+�va�L��G�觡�
�f+��Y��i�3�a�ۡBv	v�/O�W�|����0���u�`�ٕѻyf��:�F���gC�C�8ï��}�ȱ��)�;I���5{���w�}��1	���2#��^X���?�J	���r�	B� P4�_�,�� ���t놈:g�f�Ý�e���:�6"I2��x���76�A�x���!!�"�#�p�ق���y0���a�I�-��[㔮���0��>͵{��p4i%?��A�`�c��]�;@��5�^BIپ�Y�R���:�g��GF�"`� t��� ��Sk0��l���{�y�Ҁl]<���bŠ�	�������>X>I Y%b��>��v��ь]�"I�8��X�|�S$B�>[�
[���͈�E{wk��F�6% �l0Δ��,��o�a]]P�d��Ֆ��/ 1�ǵ�lFϭC�ϫt��߽O�vC��X8� us��i~~܋G�?2맱@��,@�������-x�5$�C{,��$�q��wwi`V������}o��9� =�'�F��QJBG(��F+%�a��:{������9�4x��'onh��v�9�e���~I���s��z)^���ȵ}������E����DC��T-�%�� w��O4�؜X���P���{M�6�.�kP�I�Y� �G.t�U�G�6��l[���zѓp��^;S�*$ECr!H��&��P���z[8��.��KS<2N�JV���Y~Me�U}�b|�J}Ӆ��_+�T������B����*�V�5
9��������5�N��r����F3~���T�0��K&vx��?�cy�A<n���(�,�x5�/�5���'�zE1�M��	����(��\���]��������޲G�]#¶*�M0��^�bI��J+"��ri� P��B5RJR�Õ�G��,��s���_xM%��Q�
�gF1Ή<"�V��HrJ��%V�u.�@Ǟ ��<'j�j\�byp��0����R �|�fe��P c�b�V�r��w���<3 � ܑ�InJ2�,�ѣ& �\�{I����1m�N�ʓ�<X���Bp�G
}D���pi�{� �a�f��}�<�C��A����Nl��W �^���+	���9�qNP(�ǩ�Ų�&)��򶆁��3>��k�h�7ކ2�I��j>3�����`�z_5���uY��.F�$,ؤ�P��r�=���@�i�����:.���:9@D�G�ᛪW�Y�aD���'(�7�Ќ��L@�b�4��R��Qjj)9���d^sV؂˅ﶜ����>g�P�	�{yO���Q�4ՙD'O�ޗS|�G���#��=�yK˴�=Ը.��`/��VԒ�1��(xdb�%z�=�<��ݩ $�}��	��4�/!���m/�R��cT��=���C!���t��QC��D���4�I���!}�~�O?���$O�[��P��3�{Ag@4M<�? �9)�QC���cǿ��Y�K�뚵=Fl�%\���R���S�QW� �E>�����Q��E7� �CO�5�b�_�����'/��X�<z�I��%zy�]\$DT��8�R��..1B\#;�! R�n��Ƴ���ιNn�{%^)���N���!���&���A�@KV�E�/��&<@��﬜��Þ*Z�J���
6;O@��;��R������<>
Z��!�*!�[�7Ŧ�H�ʚ�$��U�./~JQ��ss{G7׷�;�~�����c�~��ǘ�l�9ԧg�=��e�|���Zi0~I�c�i�*�	bB�y�s�dk�v��}��V�(ó
�S/Ϗ��9��Q�V;)��p
��%?S��Cs�B Q� ˒�i�W۲<9�/i��Е�����X�ƴ��߮ۂT����A����fu�p�9�NI�bh��oӸ��
�
�\�{�*��}�����j&�c�g/X-bǖ�����������c ��w��!p���Z�9��̳Y`O( f�6��9�]q	���������8I��]Zc�k_ ʴ�� �p��u�s�� �?=��#��y��K��G���ᅎ��l�p.�h=b��*�1ޥ5����]��;�+o7��x-���"��T�� �;��������r8���-Nx���CL���Zrm��bU���CBsH �u��Խ���Qy�U_�!�L��LX9�i�c698��{�j��kH].S/}��$�� OP��ǐ`�cZ���KK����YӚ�>�N&j5�� �wr�Uנ������c0v������]K��� �����k��,��$C��Z3Y%QY���Η���S^kو`L�o����b��^�C	���þ�<����i��׍����⊉f��H�I�x�4���շo#˕��K���������O�tOG���Z]�CXϳD��nVL�m?K�]R����9m����S�gC�4^B��D��&��>0=ٷ��-�RT�Q��{ZȔ�Tu=���,w�%������~���x	B3�K8���$�=kH������g��o�4��v�+�0[	�r@i��[����c u $]�#���CC��"�y���)�!�M�՘ĳg�^��w�Һ��Ո�ף�0\ �x#���/o������JW'�(��	;N�#x#T�ث'��DP�S�j��?���I�3˺I�0�+Y׬�(0�4]=v�"��Q�]��c�3ȇ�Y(t�9��V��4�ւm\��~��{�^�6<�����{`����",����A���[�)0�a OH�U Upo*E@���Cs`�7�ڤa��0V���`�-��hpT��,3���k���\����э1x�Ћ�_��"�?B�?�i0\�+dۗƾ]��S���g�/ ��9�Z���YdP�T Dj<����`���'��Os����K	o��g�{`
���9˥(kJ
E_#d���<=FА������.�i����/�<� ��|�F#:!M�.��a��[��P��~����w�=184e�2�d� �_l����ثA\<>A3��8�Ա���V o��}�	_���)�,i.������o����7}~��������	H<c�t��Ւs��H���.��!qNm_o����� ���Jبw�K`gD�I9O�1)��!� eJfe�+cB�h+��S7V�T��3�*n[�{cȯ��m~% P�Ɖ$�iZV�Feu���ší�9�cG�]mW(\�b���
t~p�k9/��f�.��H�i�?#PK}���(×M�����470���'F�%�x��M!a3�p(^�Y�%�`
�D����&�b�Y�z���gi_,r�����R�T���4�m�_����ԗgf"��(�Ԛ��U9l����Sd�����Rlܪ kW�O��	�i=��>??q��F��`�M?�9x���^ �$�l�K�J��L|�[��k���c�m7Ҿc'�Ŕ_EW�4)�������V��Af�*愽i&R}k����������;'��+B� �@��:�#� '�U���x~o$B��{�Nk�Ձ�5�Jo�z0�̔��H�o<I�'䍺���9Z��Q���cOa"3���A�J����� j������	P2V�u�]��|V�Dr6���mj',���l
������e�V�K���qhݜC�6�׋W�^�t`��`G_}�r��� 6Mғ��ѻX���\b�5]=���RRShKx�-�D���-�E�H_��B�3O5~T�cp0�QO��W���ۦ��k�(M��i�	�/ͧf���(�8'	Yضd��[TKta���d�r|Ο<��RF:���	j����2ھ�b�V�)�sq�Bцz�umL*r��+w���PǎJ褬��h %WJ�jXs.:�b�	�O)�0c:���x]���%z`ɡ�+zww��]�Ȃ���D�GH:W#԰+E$�E��LsL?��"혗v&���6��m�r2D�'��P��'�7��n�� p��5��CQ@kx��0` �"%Ć��	{NK��+mQ������{zv��e��J�-���@�� ;ө� En�C
 ����x�lX�"���Z�^�77w���6��D��d�uyIr	����OJ�[�n���<�G �ꨕ8�<y"�r�4�k���L��`����KUǑ�)��8�m��}���$4Z�3`��'xZ������S!� lbOM]� �y�Aj��Cj8��b��D��緘_z�D��Z�/'�]����=�I��㈜4��K����|N��<�"�`���W���G�b� A������" �ωlQ>��e�Y���
zBjʽG���S���LQ@�d����e�C֩%��Z,�o�׶�*��6|␴=��ȑ*�ʧC���&hoTw;x.˼6�&���r��[y
�?4�	�}�����0���<3 ����A(����{+�Qh�uC��cz��Y�s"0F�}�)<�^�A�$ lA
��A��0	�!#��Г?~���/J��^6��������G��y٭�]�}�z��Y�;�eҧ�Vr��`�7�O��[+�`�����y4��s�g߿,1��%<�=����Q%T[3j��E#��1������Iݘ4+�3�l��nu%F���o�9�;#gP�&�,��o�0�io�iu��Ҏ.x~~���s���,��� I������*N��۶��0yHd���]�.]'�~L�R�	�9�
̀K}�Z��E�~�zm��9GJٳ���!���2�T�jb�Z9�bdfGv�����펅ƶ�n�dp��Z��~�V2���ٱ��۳�I/n���qh���@OO��Im����������2w�-O ! �H�v�D��3���B�UI0@e)0��2�m�.4�1�T�1_\־O�ێ�)C����c�;��b2f�O?rBc��}"�����w���޾c����#�U��%��-��bb%Q�$��ߒ$NB� �â�ɛ�N [ �셢8N �\F�wM�n��%֒�����G���9� ���%	�W��ө�`	󳩎�x?L�M�J|��y,0� �X�2����R�`v�$�\�n�-���<y�]+���V��阗���X1��;��*�Õ��������i���!�
*e+��R�"���v�~u06��X�o?'�S��ܴ�j�X3G��9��Ǩ�<��w�@H0�4��ôf����)QB0D�H���ڈ��[�U2vH��Z���L��G��θ���Ko����x�{�`��˳��zU�b_��_�����7oy�(WʳIC�z���C��H���:�3��2E�e�p���2�x?x.Bv����� �����z	��3�v�B,][N�8��(�ea"9n�^�lԒ�j�]�v�+�42���֌0 ��6�kN$:�k����F�M���}^$
 �D�E���o�h4_��B������	�1c��+�����c`�+|�����Ia��� `hd��a��9T�D^��gQ�L�dC�fP�"�@H��8�#!e�9��]z׌�OO����^����F�9���E��K�W<����߽b�
Z��a�B5O}�il��P<����˶ (���p���u����<�`��s~( PV*�\����Z��H����r�)`�ToJ����1�_$$2
��Dš(�I��@�*�M��Z���W.��A����I�}��!?�˙�~j�r�$�w���5a�3`՛WPk�t��@r�e��0 ���jk�?[N���^[T��(
M6�~�!r���M�����[�$Ao(��sx�qd!5m+���5dm�@�$��%���%����,:��i%����^��LۂW�t(��XD�|��$��9��{�����}�S?�?���*���ų}�H[�����f���4�}��_��A���-��Ig��km�܃\����\9V�-�y��$�='9�8�1�w{��|����o�^�|>С��v�l^D�j�I�C� �<*O��6� �G0��\>�¡[*���gO7��d��}~�qĲ_�u�cF��}��wL*��_��/���~2���N<[C���wȳ�����ӡ�r*¸u��|� � �o���K�_N�F>�%�M�<;��� B)�"�&�:Z�V<18����1O����Ӂ��cZ�O��^bOi�Sr9�ۘ�|�z�,Ț��+� �{�z%-���x��+����"���y�jՆ���v����c��f����³��Jnk�@>�ݔ����ܒ��8�l"��������v�U�0� �@^��au�Y�30�x���E��X��,� ��d*�����i�� ~��4����p�o�^B�<v,lc�����0$�9<O��1��S+e�u�yc�~�yNB\F�!����'Az�dA`�4�+G���9�u/x�I	��@'�w�P@��(�������+���쥨)ċ�(�!��='��. 6I�����Ez¢0� Ů��iLWbՃGO���-����
9t'��P�9}j�0r��$g���s������Ԗ3�1&��B��$&�������	��H�	I�L����/�Ϲ����M<D�eZb<no�/V��c�\j�9��ʥ[���sնF8�����5B;��37^v��=�'��c�P^m��_~����������>��^�q�j8%[��G�c�e�(ex���_{�n�p��?y��P��!�ҫ���;��W?K���Q���	���ȒJ	�[����F��o������{��P��2�,8�P�>�>��z�b:�e�[s)x+<SxyL9�h�m�T5qN��L�(��i\����[QL�7ڮ�U0��=������5ob	�T�\��B��oU�Ɋ��(�{$�<V�.6�!�%ț�0���{��� 竫)�H��H< ��#Dp�x�"\(H��̼�s�)i�U�!��;F
?\3_|�7f���T�~�m4U𾛳!ϓж�>�** �܁�VCg;h̳G ,�zR �Ue����`���haq��F��.�
hHHB�`�aM<v5�0{k��V@��~��ɜs���VAM*���ZM��Pnx�H�����2c�Ϣyj�& 9��̀Z��}A�މ��Sd�F �	���%=�@�-�3p���΂�㼅�C,�)���[Z��Ε|8�$j�;7h"��v�r	r,�~VYX��MT<����S���i4�(1�xsw�2���-:�0J��JfX�d��xT���(W*/(�����Z��A�L��wۣ�wN�١�6��C/�ǰ �E;���&�p��2;��NkbƉ���@��?��^��e-��t���^�����un���=��o
�D�eC���_��zIzt��zK�� P��=8������ԢD��B����}��>|Gw7Hw�$C���%��i��m\���{�l�޵~�g^y2�U�ah��R��Ćg�?���J�ک8o6��a��_[��9���aK������tL�ϴж��A6�dɓ�1JQ�	�o2�˓uE��1�J|�R>�ǄB6p)d�Q�>���&���<�J G�٣'�ч� 5��D
�JA�������Rl�tT�|CF̂l>o0[E��)F�r�ui �|��41Ձ����
�Fv}�c��
HE���;	����� ǡ'�����AC����U���u锸�N-"3h=۾%2�`4a%�\����:�a��8>�l]!]c��A��A�Zbp�}��% "�Ƃ��������ʶ#�bI��L����JW�ċ�.	�iL���uЬ�P��� ,6�d�>��Q�\sI �R��6��C{ϛ;��$�"O�Ɖ!�2g��g�q��[�����ٲ�G,$v�N��݀!�J|��u������< c��@|��3�.�r\b��Af��g���`Q�82�����I���ğ�CH���~�u�y"1ӘL�b�l��\qRb���g��1�W�`=<|&��u�jU,L��ap�:oo�I(;����c�`�"s�n^W�z� e��|��"�����5x����@$3n�焂�Μ�3D���^s	����X��J���;7@���{�駟���O��t{w��#y�mZ+��i8wЫ���yý濓�<�){3�Q_��զ��Qe�$�'�R��6��>\�!o��e��e�mkh)��A����󹱕Lݏ�*x����y����M�ۉK�,W��⮅9v^�م���u\�D�T�o$1a~U�qq#o*�x�ϋ_ָVf%kS!�t�Y7������)&�����z�Jg�����hX�$��ri��B�ksƊ���x /�,��ӑTACG���RxE�Iom>������%���P.��a���� �x<���_ ��Ͻ �
�o�dy���U~d%�;���q��n8�l�
�A�ݻ�Vsh�ab���qn��)�{J|~bUP�@���z~N��ݹ{�$~�_3�"��Tc/�[���^'G�I:��jk��Ef�Dʨ|3��stjyb�����E>�sA 4��{���	��L�ꪦ���A�2�&�؇2�� ;ȓtOWT,M�!T���Hbp����Sگ�Lt�������I�3i��A��c���-h����#B�7S��;��ІE�Nu8�P����ݕ'����8_ڑ��i��$7��SL���ؑ�E�r�ǋ�=�왦�!\]C� ���k��O۩�'�3��In�+��*!4��c�!��]�-"r�X~��,<��.W���0p��p\s�ؐ��-�Ƌ9���d��J��ϴ��o��M��U Se_��{�R	>��� ]������f�r�cC�YȺ/i̞�;�*�Cq�������?�����?��M�� ��U$�$�Qt(����[^%�2���r50�����d��8�w���=|��y����#}j?z���L,'"��&�ʞ����wI���w?������ۛ[�u�`�T���I��K��zZ������/���E�J��� E�C��6�]N���<e ��>�)��V�\�������~��Hq����O���pزWR�,oW�9t�s(����Z�����g��D�2�|�Z��u�$_��މ>V�M���8&��0l���룰�y�M�W!ɘ�?��X����sQI�*�0�??.�!L�^ [6T�
�W��\
Ǎ�:������0>09x
pH�D@�uZYjF5J�T���=B��#E�l%�3	�	�U`ak$O�����7���Z��i-$l�x�0p�Ѭ*�f�ʀ�<���R�����yI����M�Gvx5Ȼ,)mV�{V�l"	��Dn����ӎZ}A=u��Nc��s�`�r���$J|xo�3�I�"�C1k�Ax�$CL힉7UT�U|�d������d����H���<���2�}/n�"x�xM��
n�.geI�o|˱3����"�m��)��������[bn�Ӛ�%`�<�!}h��� ۝�ox�|��GR'�^�I�|$�pJv~\�ꊫg@����/@=p���6p1�r�:2�0	B�g+�d:ѱ���jn�.{,,�&�Xx''�BC $�=���a���Ġ'�^.�5VkN�׉%���^8[H�#X:97Qx����	^i�j�Cb�97������~��
Z��u��]�.{F��S]�d��c^m����Y��뤹o?<��*�����P�)�hj\>���_ <ȕ��@V$?�y����9+���^��@h��
�۬s�]bi������G�FwC���R�����4A(�~���K�/(�dDe`� �]��܃'��G��K��m��f>/Mte�-�$�T�X��3U���W_�8���=��pܲB~���ZU�g��Y�?�w��!���C� �[g��sR\%R�3xN����3�YtKF��c|L���^%͑\}K�,���T�n\��C�ɉ���s���A*@���B��ϑ+�n��m�����m�� MTn�����`���{�%9�$IP���� ����i��h�v��'v��f�a������ ��f���"���Y��=4��	 ���5Uf���oT9WQp.��������9ٶj˳�V�4�r���b�5�Yۜ(������pB"��w��P��Yya
�Q�E��t���YPy�\]^Y�0��c�3�>`��1�ŵ���i<��簱��E��ĮD�v0e
,F ��Yj(�̽��S���J7����|17�aKW�;�b݀����}̍�U��k�iٱ֤k�"ь?'��L)���D��u��K�A�Y/�����6��~&b�4SNmw=�7S0��=�ن���
��m���\��L��`F3�J��R��~!���N�uQqB�qs����+7�`�}�\��򟤖# ��f-GĻ`	��-G��r����Ux}E��O0�Q��������"��Ys�)ѐ�p����	�Q��d;��2ǩ�y^�����gJ�ݗgd��倈wK������CX�r�C^	EY��&��J-�ij����!�#��O%/�����?o�49�C�|	��Z�?��З�
��&��S�x�&Nǰi2S�d�kW��D��"�o���T����h�L|��R�/%()�n‣�����*Vq��>�J�_^�^I��d�t����P��N����7n�_}�^_��_${�[^��o<�����o��!E�IX�͜6�VU����H�e���`ɿ~?2�FE������'k��F7�`��I�]nݪO]�(9�4�`��C��W^"D�p��rK Ǘ4� 4�.Ų&��ۭ���0���$�aX��Q�U��`˽��*m9�(�S�dķY.�^����zq�6��ʁ߱~ڄ�j���a�v�Ȋ�\<��X^p�C��d>�(�l�M[�͝9 )��>S��.���'�Ö��l�>yLT������d�P�"P,���׊����z���1��?��_�@�cN����x��� �"0�(��� ����Rr���P�`\
<�5/�7wu��ժ�����T(�?~�k�`+V���/������-���[�����[�G� nS�#���/������89xX�u73�6��KT����f�Tc�;���&���́�777��ϟ���CN�D��X���S�_���m�,�k����5-����7�1�Y�U��Yw���ҴZU����G��ˢ�_��q겻�8� ���΀�H�H$�ln�=�\mw��+��/s:f(�W�� O8�5��:���zܩ���.��+l5IzR��+�N����ys���[x���=�+5B����
vG~WH�������?�sL�֏�ʒ͡0���2�0G��.���BT�V�y�dtn��������a'A�<���Di�,�|R��5V������0�>�����k�Q���M�Y�/L�fN�^��N~�0v�]����v�Y�g>��.��qP�u L��`��a�1�) Ē�\����b ZrB�u���.�ɜ����ڶe��=�0��e��cs�g�3c�d3���<x���	�� ��K�HE:���v|dcO��LN"��A�XP��4w�"�� 
I w��]�Z��	��9��[4��i"^ y��k@���M{���P��vj���l���SuS+�>D��ٜ�Bt�a�˔���E�5���O��^,�(!�ɾ�YK*��X�I�l#��O��,��Ș,0�I.iC���s� �h�+G�Tzn�hz�&���L�(�g���l���0����<_R�������˾Ke��l(�!�3��6?Ks8w�O�K�?������K�^�8�����m���s���'����j�`��ͨ�t����cK%v�(��E(��`\/ƀ��'���Y������b��{�:�|+ �����?����!;�j�0�A��ġQ��yͻ��5'�^�"��_��
�O+P�=`?Y`�g�a�Yx�r�A�nj��y�1�z� }fs��ɻNvy>��י��zF�^@v��?����-�-����1�\?H4���I`�R�G�X_э�ᵭ]h��^�2-���vZ��������B��&$6�Qϓ�ف�M�+K[A��w����W��+��K��{�4���j����o����P+g�+������)f�	T4�.L���YK�@ӑ�b����d��z�umF�VH�C=��.8�`A���'^��Q{������
e�H��~�у�xr���� �!�D���		~>����T3Цru�>/.98��e��ڧ��Qf gNPCצ7��9m����O������+^W|�����
���0�3'��#����ޙ������좉��ꌀ������F�3 ����������E ���|�/���dQz�@�I�7�̥��;9Q p��N�����=�=�!�`0v .�]�Xd�s֚��*�������m
��b�,��8ZjgU��l�'s��Q�O�>��Y?�5��k���O�O���@(�;�V�0=>t�fj��3�������u�`:(�sm$�)��Aa������ufB̲a]0�I�?>������y�Hx~��' ��E�j���4u���>�����pq�w�4�+��\�xa6*̓XY �&�_���~#��(s�T���xW�i��� _���:� �BS�;�b��}��;O�|5�,k�1�s��PǞ�2�6b���[������T�u�x��ގ���窬��d������t͂=�w�bSy���dg/�=�$ұ�(a��<)?�[��=��U�x$}�C�PFNl���I����kjV�ZGl��)�1�i�)<�N��g�]��Y�����!_~kSIӞc�lycs�e9kl�_Z��90l>�9Ϸ7�C�xǊ)�<��� ���$}�E��������o�|�q�*� xN��t����0{�Ȧ�L�g�@����M��gbV><J_�����oǁ�ˬ�vlh�B����c%��r�R�p��c6�h!�5�9��v���b�Q�b��.�O��_ٚ8ґs�<����;��Љ��L�Ld>�5��l�ؠ�w���#vB��2���k�������0�6����+'�7O�?�� |@W�s�`0����-���X5Z���Z�粕.�����4�<n��Fbʀ��t)[r�v��y���B�f�8-�N(�a�-s3�X���}
��&�x�`�
n98�8�B� �� ���d13�B���� њDV�㚅��[��l�Eq��'���2v�b+
��{�G�1���V���:Z�Pܘ-��ѹ���4&1��/X>#^C��x�m� c�JgǑ
d[��:�0�4F`)���P��~�	?�h����a�B�00�XP�5��G �|��3ׂ��e�Dy>��yJL�!��Z���x���̀��A4�\c\��L��L��׿�h	���,�Y�<�i����������&_��O2�,���黽�k"����=zN?�cȀ��w�<���y���G�w��2���bU..�"���]@o�J��`� �D�r{wGI�V覛�L�n:�9��@�!�����Y~>W�p����3Ԁ��L���l��v߂����R9.[�&����,�ґ�r/s+E(���<#��￣��|�	r�;&���ci#5y�j�2�pR�q�o�Q�q2��i#��,8����DGa�E�Յv!4�ݐe�y�g�]"��a0����*���J�e�ƫ% �#t�4�'�������W��7��W~O������uU����y��� �ui��zoL���h�V)#�1�9q`�a�h�G�F,6ź2��1��n��e?��'���c�/"������{��1�n;��9�z����m���P*��>���?8d\��_�1^s᡽4Ze �����E� ��RU�1lɰ�A��ͧ<	?p�=��x��!V6س)�Gl2M�P��k���9y����cW%�"/�x>P]B ���G��V )�Q�Boֱ�>\{�bC�� ���>�W� ���-��iO��yl }�"��b�֣��\���o
�":[��Mf���@��1p\r������@?��V����S���#��q�pΨZb�Gۡ,����:�7���p���4�X���kbp�g{���=��a�zq1#�ݝ��/��oz>#p#C ����5�7Z���P~х��"�B�p�>�� ���F�#/JO�]q�����}G�����M��o��cR���˕���B[�͗{ѧ�lQ�K{1�I�4�����B�y��G�?mA�泧鹳��6�-Fp�'����d&� ���]����d��΂�`��+1Lu���r�S{X��q���Y���9�U�N�c�P{������Y��1� y�����!��C���y����uh�x[]�s���DOv߸��+�X/�p����8�}Uv���|�}�{�1c��R !5_قA�L�)x��ݧ��F	�C�� �wVlā�:�E1US���k�Rt�g��?E����_��rj�����: o𘃍�$�ꂁ>> ������h�m�@ |'m�÷_�����>���Cp[u�g�9������W�Խ@�X�=p� �Π�b"�`�n�]a�zwV/��!���o�$�>_2�~	X68���'&c��l�_s����Z�{'�wy=�Kb���D��t!�	�{ЗC�s$���8$X�o�n)2���-�l��[�k΢K��b$�y�!�i�^��]���^^\q]�Mw����y.�v�W��(f���d����cal��8�� �@ӄB� s� y{��Į@��s��"����۫�������HPl�;/U�A�����"H���%
[�e��}�������:��.����ء6�R��+��}�u`N���h^_ˤ�ڐ���0�R�w���}�10Ԛ�x���`����F��O0���(6w�s|����%������q�b!���?_ϐ�<R� H' ��0�=GRKyhx���8�k�֢~�c���>�߇�������r� �tP�a�8V�t�{�Y���� ���hw���2�Ֆ��J^�1�dE�=[�Vg=�?~������ �߄���������|���ux*ڍ�܌hj�tT�����$@���Ƹ"S�ѡ<�tq�y1!��^����u�8�s��Q ��i'p� v0�s,���Ǜ������>Ƨw{��PH;��*r�m����������?S;p���w��z���tX�~|Xθv�(����R��I����r�������Q�]�Z�b�Dctfm�ύ����.���W^�����C�����?�c�c��c��
�:�y��~������S�r��t���r��;�q���wG+�I�w�٠w�ё������-��h?��>~�yk	�|���oV|�_���V�뉖���'�*�k��	�u_�5��E��zvn=���j�䠾�+	B���\.�9�u��)����N��x�����h��%�`tF?�NA�q��2�)V3:c踶�#Y��I�@�E*`��`i�H���3<Mr����x�@����	Q��	L&F��B��K�XA�U?���ң	,��@
�+�@�	�}�ފ��We��0��W6[В��Fi=�Ml0JL�д� �Bt��^y ܤ@� �4��D� �''�^�K[��o�fk�=�O+s��	��Ĕ�S姳
&�׆������J�z*ϱ��c5�)��+�VI$�yx
�k����d?�n���}��8ۛ�lg�2H���%&��u_�e'g��Y/|�qho �''>'T'��E���)���ĺI�+�7Wҟ�T���W^�iS<�J�~�1�i���ы�����v�|�@/�3h{i��ק�7X1~���䳭��06�����g,?�Oj2۰G�
׷�::����N���֬r���Mq�&�{�˂v>�y��w���x:'~���y��ƨh��7,O������y������P��d�Ml��k[JeȨ��j�(ѳ��㼹#]?���{�w��N
���C������HU��*��>����~����)PW <4�.�:V闡����u��l�AA`+��ڧ�>x0�͆���cq�1
 ����ie��[;ƕ�YB �ல�1ZV���i�xF�P��^�gWM�~�]:%���Ԍ�֛�&x	�I"�b̃-1iv�u��9-��tN BN4�-Yh�������D�a[��[�<���.��I��6z;~)���C~f�b��n!�����1K��c�ۥ,W�1&���Ҟ���l7ZlQ��j��7��I�{8_�tçq��`Bx�g�|hm����[�Z�kMߐQ��!��,�U�ђ4�q�����Ą�/�3h�8������_vT���C�~(�9�1�;a��õq\�D}���:�%M:z�M�rJ����h��w*k���n��ce��$ Wl�'�A���1�u*q����!�S�M��,����׶�?v�Rs���:��4�A��)�'�j�Iy|F�N�h.� h�hB�R�퓴3g3�)]]]��*����֏|��o��KA�SPCpʫ[|��߸q���Y5UkN��6��'0����.����%��ԋqp����/�<�89�u ������y������!�o�:�I��=��	������=W2؎�I�.ۮl�z����C�TH��Ep+Q�+5:��BQB�B#�I����y�� �Y�٢CW�!���<��E>��e>�}���|��9M�+��+���S����- �V���O�s��$�D*��h_�:F���x;V��6����z=ȧV�R'i��Kќ�A΋�L�]|�`�/������V:Jz���1	��0,��0�:�$�����ba���*�܀�rj������q�X�A4e|�mJ�yq����=�m��W�B]tWUc[��PB�yE�MG���Z�hA(�hY�|�>��~GV :!�Q�(v<jّx/{+���G�'V|Eg�+Z���5����a{��: �`NϾ[Nt�t�v%X�5�$�	��"�2�:JY�Z(F*��m�gF+�k&�Zض;- ����zR+�nE�ǙKl#r1��L��/�������0��xnK%�3,jy��]d�Dz�x��D��	l���h��:�L�o�x�� ��W��Q��Me��0[bN�$�^1�Ejo�
�r�TyQ5����o�܌�TK�3R1MC�����|1bg����rr�i�����@�\�����m��ِ-,RO�u��e�[s���t�<���[s���y�-�����w+�lO�/��}�d]��7��k�˖jrX֙f��:��8�ԃ�#����L`�~�b�S{�N�u��W�;h� ��mo�v'��׷�����nA����{cuc�f�m�A�}e8:Hӂ0'_����s15�=��}'�N{*ؽ���liB�����ґA
g!��W��~{�+�ؐ��yHru�:��Yr��D��x\�B�2v��ߟ�T�`���]�]���-���y&����Q���]%ʩ���Eb�	�v� ��v�b]#$�w��r�����#���%ʿT�q`�dр�����h�nYtEK�d}*?�'���E�C��s��Dg��x?AM<
C��ѽ�:!N���'�(r��̨��!�TBHqb�� vd����c���DnY ���e�'5̜���<�u�HT�#�(���v"�_��X�F19*�����xţX�6�L�`P��\�1��E�y�KI���e��c���u��1{��5��� �i�D��܉}y�]�!������I��q-m
��w��8�=�w]�t�s�?K�pMs�c��������w�E�ʮ������Jo���cV-�]�����cI ���~�p|g m?�)��p�sY�������aL����`�A0p�n������v؆y����>v�&������C�.NZ/W������»/�����Z�� Η���	��}x�?���7����
-Z��Y��U'MMP���"����eI
�� -f^h�/�y�g{�|�����`7�:�!7	�32�ä��y�>���~�6�!�-(xx��kE�v#��I'/{�^�N��M_5�����&�$>Q�9)�S8
���f?/S]P<@��ꮄ�&J/�ʷmVj@��Z�������fO��1{Ԋ�o�Vs�A�g�9t�ɚv��@�j0Z�_�1���2��ު]yb�-s�B�d7�n�.�d��[����W_�R�W�{����A�&�s������ ��u���vd��Hs�@��:\]\��M�����ܲ �h����9�jM�!���Aᑌ���%X��'�H��!�۔�r�	jY�+���*�� g���h	 ŇY�P��	@*܃��ÕaS{g���@�tg~�@&���ȋ��1�ԋ��탕���[�/��'�-��Q�%�%$gv�~N�"2���d��*��t����ʁҸg�>��� w����R�$���vf6��~�d��9\4��dU����b8X���)�[U����!�/ �����Q�d[ �R!t��i��,y�cY8�9���:��/��e�+���]��3���Q����S�y���`
�]�:g/</G[i�(�~��o���}�p,������������֑��t9��۷S<���������@};���U�����ccV�W�����X-Uݕ�b�/f:s��Hd��^2`hz�����P�g�⿎�/Elԗ��؜�k��`��5맍%���=yl���~���u=�fǩ�G��Nc��Y�%�!�:�3y�=�����X=�XV�SV��"U��F�v���ݬk��7�[��h�r�s�sa+���H��THf��+���x��Q����	A6#g\V�;�[�&�6��){[�pj�9�9M��T��mxynb���@^�7�sPL:PO��A�B�-bb��Ԗ����3 :̢��+fc��$؋��z%�dPgH�+m�:h�����!זX��hZ�6B��$j�CoCa�]_��?Њ�:*v�܊P(���=ӊ=��Z��y�$��9���las&�4	P8��8 �Ø�X0�R
x~���s)@g�&=�r�8�ۑS�5Eal��X��6�c��sP�=��]L��4�@O�F&��c� 8F�8����K+� !�� 7U���V�U�c�Ih$�s*ϫ�jz���x'���{��\H7��XNG`��U7uP[�\:�'^�(Q뵭Wo��b��rK�-�nyx��i����l~��|/�=�,�s|��Ɠ���5�Њ���BG|N����w�QsN0�{�Qp\�������}c>_C�7&w>N徺�yhќ������tg7��c�W$'���'����|�@��ap2��|�b~�<&σhi�t�9|y�O�u�3vX�4��aX4�&�n���D�Ў� ����� ��9 S�k!�.��,zG@~�Z��c��FyL ���8��F�^�����Zl��0H�������qe2�7��!��;��bC.��Q�yit�ˆ�8Y����+#+�Ÿ�����L/|<�r��9������	PsP�T����%�K_O�]������z	��h��3��.�s��Uk2
�,�e����=��9#��F���`���<�$t�~�?����$^,�n���m��^چ� �g��������L���-�����5��0�=�K�����x3�*V��*4M�@���ǻ��p�S��s��#� �2�3�Z� ��=f0!�!�;%W.z�ɸ�8��	�t��(����Ђ��h-8��ɶt���J�%�ŦY�B-uh[���� 8�N@R��F���� �-O���/z^��3{s�"}�US� �ң/b꽧�ŕlJl]�I�1/~O�ua��B��K� ���k2J���ڍSa� ��~�`�m�3���R0��6��������r�+&N4���~f9p���Y'��:��r�
=�����#@Q�\�BU�ari������a���K�_����!�[
�6�q�KL(�kԳ��|�c`y���-��`�ɪ��*~�k���T1�ꦥ��~SN����a��&���fͱ��K��ԛX3�'`�g��,����c����گ؉_[�~�MAQ,�5n|K���~���&�Ǧ�䰙 ��j�ԋ, �c�\")B����|��m.�@�Pu�_f_��t�R%U&����w�e�BGף�A-��!����{^^t!BQ c�ZV��c^��2Uh2��� IO�Z�r���qKdo@�/*�CF��k�Y����΁��6d��V^�'�S��Bj���z��t0GI85A7�2��X������L��k�;֓%�"g�n�an6{��X� �@�v��}��<��B�Ijusvm�El,q-.����ao1 �Q�~���a�/����k�B����|Y@�=����V̢`)+�uT���L���uH���6&�Ɗ%� 6g;�����ȃvxU�m,�b{o���\ӡ7m��d!:������v�kY���h?SK=�vH���A>�㝵E�M�~<�2�@;��@���zrGc6Y�g�#�Y�9�r9��8&%�rJ�V�O�����{��x{k��f�1U����ul��;lvm&[�].���4������=��Ū3�؊0iY-��9_�XI�8�t=�������
����.8����l�Q������t�m���_Av�<[�e��8�Uc�ἓ��s�	j��=�x�&)��s-C�BJ��|hgy^;G.����o�܀�s�9�<݅͘����I �Haz�8i�sͨ�ZG"�5,��Y��Xf8~��g�2O3�k?��aX��U-�Y_�Ѿ6�?&�!�����c����Pz>�q�`��E0��{T���{�/��ϣ�֮��-(�/-n%q0zkATO�����4Zy~�-m��c<�V�N����a;���������������9s���_�E)��Ej�K���԰=������ȯ��y��A�L���pD[-O��L���q�i˄�,ޕ��ܣ���W����l�`��i/1B�F>�,�'b�0�5�kp��d	:g0�>L : a�=X��O����n��D-0�X�"�Lս�n�
`R%�߫�o> ��'(Yۍa�6-��@�+}���@�k���n͒���V�	�:	
�.�`f����,�EVX[���{����nP���8+�{�q�ָ^{ӔQD�	Z���J�//ﯧ('���_p��i�:��'��f+^'*�ӁBqd<EV��y5��]Qo]��XU��"��Aml��Q�4v��(����9�B�s��&_�l}ۛ����$��j�H�f�LF<F6�*���B�+��[Y{%)AB�r��8c��+���y�2>�h��$��/���s���/<��[��K�O~�[�؟�;�n�թ����de�r��x�
o���Ku��5�>^�*���'P���x(�2gݞ� �i^)�6�oM�Z�d-t�z:X�OÀJ�����6�|��V� ��}'AJ8>�o9aֳp�b���U)�A�π!$���e�_9�j�Y������Պ|��rnR�������?�g35/{[lƾ�q�s��5a�`�Z֩ @p`k����$�C��Ik-/d�L�w&��.rQ®vV�R�B-��� T�{Ҩ�������D�̑���|X�D��,R!�@2}�P�u��~oF;7���yh�:�`��X;P�{��XAdo�oMğ�bM�U���̝d��]/��Yq�"a"l�4��G�e�DT Dߓ����P���x��y��E�i��J�R�A��t*�uzo
j�w�ve:c��]�iU��`�0�]?0�S7#����� �$�s8���
/^(KA,&��%�1 ۡ ���|�uf��h̚ќQHR��A���_��xt?����Ma�dV�Ҧr�h�!훩ٴ��z,s
����5:��͝7�6�2������t�'~D�^B�"�!mĩ(���^Ty\	0��IS���������5� x�ặ:_�����_�b�E�$7�˹�rl���w�2�6z7�Q��n�)��@-bV���?�����,��� �(O���V��h�k¼G�G���=<��'� B��<�}*��ڔʵ�m�b� �8�b+%l�� ξ:S+=r�ɀ+�h�Kg��ll�gwy��02��Oy~�r=�����XјJֶ��]�j��o{��٪sRe�B�g����ڭ���_o+B|��h���g��������� ?�<�������
����k嗦�����	�cbs͒_���$'�Б�2_&�ry����J���\�G�r���(�E�h��x1�H(L$Yo?�<�� M�H� ���k.���"��H��e�)=�T��Tu(A�����4P��P$pnL�<i^^�����*Z}������Mvon�-�d�`�꬗U��-L�U�<�3�O�Bg�)���T���J��J&@pO�EoZ?�{�%�&\����U��X�H��s��[�;��8jJ<��?'�SeM���R<&`0z���e8��
�T�8g���y��#?�qqss#7�3��:�V+\�~P.,N���t\?�����D���XM]���8��e�8�8)�P�X�J��A
���[K�֥�н�+�y؛ˊ*��>y��ș,y6�+��M�R �-㺲=���8��U��g;�|a�A�r,	�	u[�h�\�^EO����+[I��h����~�~ʇ~P��y�SC��W{��~�5+:����K�o�;T�$��ho�����4�8Ъ}��8U��Ǌ��1(����͗��a�s��ޅ���k_�J��p�'G���qk�-��6'璎?�������:y{�+xL��5�#�� �%x�=���?M�MR���a�h�bȷa|�\�r���놳hy�S��<�}�����u��[��Mm+�
�%�I����U�>��m49A�U �gװ$'��R;���eV)�N���yc����m�=��������a'�B3�����'Y���h��c$�`�@|�=�V���n*�c�@u��i�����lm$��F(뿀%� 2{�_S��`(ly��H��36���g�/�%�x?X�α��E�-a�x�BI0�@��8�5}���x��!Ƃ4Gk�����l=肏���M.���6A{��/G�V҉��`��`����3.B�y�D����+���?��⭜H�I Ng���wq�:���d���]쨈�6}�0�q�,���"c/���%B��)���%A^�h5��f#��k�m��XZo	(b������_��y�[S@Y-�� ���`Ym`����Z��9څ(|�Χk�ou��(�I��}�3�ܻ�o��B�|9W�/̽V��i�R[1>�ô��o�7��'~7 k4��>ޅO_��ۇ�<'>�B|��]/K�tp6�c��µc+�X�E��.߅�y����C���}���G���Ϭs��m��w]�?�����#'���)�6 h�#<ދQ��8�0�>0��"/p�	�)�`���lCu�1q+C�IE�Ƞ,D���75�Щ� ���*�:Z��kpp�n���+�����T���@���X�hƙ�}  ��IDATEg�S3����T����	��Р)߇r|�j�A���|�k��4)�/(AQ���Sج�a��أM�	��a���}xW�-.bL�e�5�xԎ��Wq�%�*.hx���OdQodJ5I�]{g���U!T��s>�%��N	z
�@y�X��vJd}��k�N[�i* �����L=�lau6#M{���ن֊ww�e�jA�@�C�np5 -t?����ڂ��u\̢Q£Q�q]1�b�9�ч#�ޘ%��O=�a�q���c��C�Q6�h���bK����a���{�#�K:9���1y��#B��h���ٗK�|�(��x(��a0� ���1�U�ڌE�R�޽��7����I &�G�V�� x���;�c�
^]_���)__X�c��eh�����}���.ߣ��"�̚���,�'�F�$��%��>�Ŗ'>K�}��;;�)�I�VE��b�<����W� ���������@'7�xct�B�Y,'��g� ����D`�X�Ƴ
����Az(��"^�,i� Z���/��{�Xd"���K���R�U��T��0ѷ	��N_�N۴�*tmծ$ֈvTX��������ȝ�<e�@��Q�������� �ɱreos�T���iS����0�9����B�cf@�9�`��$�j�R`("�b�Y��u�c�@L��l�V����/������}:�����z,Yc͙.�k�`:X~OC���O�^�Z������!%rpP���>�\��
��=�Mu�+��9���&.+�E8���&!<j�OG:;W�x̹�cO�ч�`��[sm9?������9M��pM�4���A&���?����3��
�.V�jFj?Ӽ����h�Lr&-�Hb�3���g�ui*�/mS-�CHt�uk�:��������5�fXeo�`��Ζ�U��.Vō
����#c؈#��m[�;�����Ĥ���?]���1�6 ���i����*�VB��L�ի��)� ��?��v���q�|�|��<ǽ(�(�
Vq��΀�
dK*?NV�d촟lmH�	'���י��n�Ӧ�E�8Bя����ۡ:�������6k��m�N�%�Yu׮s4!�֪d`e��̱��
M�M�t�t����EG�5�p����0zѱ��+���v/�֝�bѮ��aQ�ژ=�8�ȉg�s8�ς��Ĝw5�:�D^�Ͽ�yr{2���J�y����ya����q/p��>��P�s����8p�_���nZ�s{���!�7���)�=�{���m���S~����;����8��cڠ,�ϱ�bМu����[[�����!�����mc���]���9���@~]PFaU��w���bVu/..�s��ʡ�u \4K��)���<!!Ag��sv���y��j����t�r�v�"�!g�ru.rN�]h=��j��j���-��9��
v�|?�9�g!Y��N]���������ݷ`N����j�r�=3�nBvu�J+���^;2�<��zP��!f>:�l݄P�
���5	������fM�OX���l�иԿ��4i	�9r2���K�xrP����@�uhL-&]�V�g�������|Z��9�-��{ʤ��g��?��1#�A&�;O�P��������]љ1���,�F�Γe>}�q W&������5ۇF9J=��po�H�Yg��;9�V�9�)���T���;��0M.�X�OVũm0���r5gH�E��l�91��~��lHA������p�3,�$����0����ϼ�h�^A�(E��,�?]q2Z��J��l��cL�E�mC�;4��P���i-
g;�#2��n H@@��~-�1�w��b�U�|\�cpm�ы���`���=�wg���[V|����v�L?�µ&[� B,x wB<�9 �I��Ç�������緙�l4�h��f�g{1l`���Ƃ�5����+���ĳq�c�F���a&z3[��;޳���%����0v0�Zs������+s��؎� �h%׮vƦ��P�_ u <-�E%W�q���Ԏ,�ĵ<�����&�E��(��g�/xSIB����&|};�P��#��CY��|�o��;
S8b4M��+�����Sy�t�r�9i��-�� H�_����U���Dk��1葻�*Y�ޜ��p�>�x0��{��P� B�w oy]	B9��^ե�d�e�/��� �K�o�(����/ښq��8�c}���yY�29������(��7���_҂�@�y_*1سs@���e�@<�iN�A����l/��k[Mt��ϛ�z�|g�vͿ�N�*�I�hT2�ś�!����D���#���.d���
��D2A���rު(�(��U;�D���*���G\ �ei��%�3c�<�d-��
���U\���%J����9���ߓ�sq���3w���:;���f�<��.��i��q|T[���;e|2��V�0�o���V9�V��Et�
>���3!���q}E|�d��ti4������9x,*"F2еN�J�4.%�H�5Pܵ]��� jg.6�N=B�ź{sH3�z����43ez��caWh>�*ԬUD��`�#'-�#�ٵ4�/Z��{�?�(�]�Td���Zx1Aa�z.Q�E�������-��*�?(R�,Ɣ,��-AMܿ(Ab\��%�S�&��]VS(�Z��,,__Դk��ѩ��O��	���{N�Ί]�J�+ћW6�1}��k'����EFtv���l�O�HB[���іŶ�|?@��z�nG����>l�>�u~����X����N>���_�|
77_�3�f<����O��Ɋ��b9�x�_�؜���Q�e�tgv�h�������w��Q�eΌb�^:9��.����$�%	�����:����yx6+�  ?Xfs��f@vf��z.��cnS]Wm�U@9��g�X�c�a�g���2\.���|�c�B�� g�E��{��I@�;31��������1�\��}`~9� Mm�C��^���� W���H+η�
b��^�|�.����("$V�����0��؁�Iޫ�]N�R?/[��!�΂�J�?I���--E�'�TPic���r-�o�Ց�_:����fE��ߗ���_�t�5�&``�44�}����� 1f֏>�+,�s�#K�Ըճf��Ȫ�$�������݈�r��j�dtǚ�Ux�<����qCK�ۛ;2$��@-��o>[���`�O�� ���TL���#O�������A�e}ऺX��{J{j�l��p�.���L�����^XH��@���ft��m;;R��	�	*��A�~ �F�d]X�����lD5z�Ae9�"r��
[ �۝U�TmZ�7���:V�P3��/�@
E��A�~�6v�w����fKޯظ�P�:@`f��2�`;�Dڵ�j
���1��6�>�X(pFp��؟W������k����GX�
l�S����qg6�^�t]�R�E0��1ﱰ��Ta� ��tox�]�W;r��r�+�H��Zb��X���&�X]4�����u-���^t�jmtP��	��	�b7=ܷd��ɘW8��	w�"b�JB���6�6��7��;�_���#h�D��jSa�^Mp_M�=�.�N�?��ᠿ�fB����V�����4'�]���ܪ5���
b.z^]�w�h�s���ae&k��~1�n�s���Bȯ�e�M��_���H%�}��oxy\_�	�d��(�t�hA�]�֊ok� :���,R=��wJ�#��]N�:6��	���w����T��6�4�2x��a�v�R�l�`��3
��M��mH	�n�4?/h�pV۳�|�Z�%��9Jno���s��jst}��9F�`B�rӈ�wPYn����5>bl�	�_�WT:��Fk��\\���1o��u����	���#�u4(Q+�XXo��(�B�8���DX�Fэ��]���V�^�B��`�Z;O�ԚϢ1,�q�'%1��X�_��}Y�5A��Z���7���ڇfr��AZ�Ww��L�m/s�������z�2b��^tV4�&<�(����wd����yu���B�N��upl���b�$۴d��X�u�o�C���}iˏ�LƤ���
�My}��5�P�bA��Q���Ӫ2��y��Դ2��yNV7�W\�X u�$o���aȑ���%י���M,XnH�[��۾�:3y�e�2����ކq�m�)!���l!Q@�)?��9�����y����3��"�4�0!p��}���@�8�N'�w�(��1�bj���zkr���W�����_����p�s����,�'�5���P1�Y���[i(��B0L�N�]�ZM8��g�~
?���B�^�g��E΅��δ6��){��e�xO���۟O�~��ρ�o<�������>�|��s�������H���	�b[i������w���&?o��d�v2(r�)U츒���p�}��y9����M`�b�2������ �3_�B�d���o�ָ�V�ꇯ쐰H�E��21�-�l�I�֟�t�*��#.��)	Fj�alȚ�ĩAg���,�M͟'�ۺ/�ŵ�&��6x�E����'�7B���X@tpR��hЌ	����hqP+��ۢ�Hb$`qD`A[�|d9��> 6����0� �`�(��.��8����Vv���~}8�ǃU�������؇;�f�[UGm>z�����r� �HV��𞡊Գ�i�$-����֞�h�3����c%Lէ���tL�Y�}��8n��]H�1���ƨ�E���;�%�[����!�b��lg���0�VY�{Ӝ��A��6�y�ߓAۧ��C�����8V���t�*Td T�yR� ���~�`{ɹ��,�sn}�ʑ��Ȍ�p2�b4��rx�hxv��^��
}(��\����1����=� k�,�AR��K��zo{K��p��%W����p��ސ���}����ǁ#9�	$��&�76Q7�����"���` �����'�����c�y�s�C�J��fK�_ϊ ���KQzyf=Z�K`�&�'��jd�9�[�Cp}�6p':�tz(Au��>��I�&n:R���wǯQ�]#�Iq��U�~R�&TݴFC�;�w�����2�}���-�y�7�X�p�V�K���5r�����0[*���<���� |u�5<��}lb�:�R�w}���D9��h��1����%1�x?@�d�	9�(�iCA�<��%к暋u�܄�'D*j4 �1���V����L�7����C#�?3Q�ΒlKT��kuo��P�)I��[4��"�a��4Ƌ���Z��Y�>����y���y|x`���Xc���R'Z�W�7 �<u9A��r6,>;�ܭ�Z�� ;cb�
�#�C��|��fV��p	.�k:z�e=���K�g,k�YA�gԙ��@�>t��;b���Pe�Y�۞	����?���F�8�3���l���_-�}���w+�=s)Ll9�$�"+�����e��ca�%�W�I%t5G��>Z`��|���C(V��-ȥ�g.���,�Ɏ^���a��"��Cj^��J�݁�1��I1�V_�+Vp3�hNR���d6H;1���t.j~(�>g������-�>S�%���&�V[#4O5���@(9�{��8�~Rd�Ÿc{��S�ۿ|�#�j5�1o�����-�d`�-2��҅��m�<��:����nk�
I��:>~�����-L
��y0��aw�8Y��d�ޝNw&��Y\|~!� BԷ�[g����?���_û�+��䱁By����:�x~HC�Z#'^����$3��@b:1��3:<�o�����o�o���&p������Ga�?����Ύ�ISX]���I�M^o��5����,����i�1�S�ym����>��"�����˜��c"��}�g>�)�W�́�f�M��f�*���+��H�v;�vLv#�*e��3����VjC3[���R�k���gϮO:Z���\��������Z�}b{,��X<�|�c�p=���m� ��0'�����-a4o-.���{��nÂ�˫wj���a!0��l�G���/�p�>s�ƍVu@⍄��ֻ�!�H^Dg�m�Xܠ&��`�PO6� o�/ނ���E�9ہVK�����T������ˀ������g����"]��1��_pR��-k�3��� �$�3&g��`�,�vv��N�{|��q�:�����d�-cg��l�Ǿc@��%G�Y)Z-�`�qG^H�>@$�h�d�ڽ�{��FA��J�3{��-s�A�W��0�� {0>�C ��X�X�4A8���Z�9ZZ���7�	`_g��/��]��7b��(�<Y��6/"`���� ����<�����0� fGP�O�?�Ȓ ��/��s
������ӓ,�-�d�V��[�����"������%G�\��v<��Vh�,c��`@�~?���6�bű}v~V��<b��\� ��b�
�K ����ϓ����J\~ϭ�۾�L�_��v� 8���ņ��VDc_���n���5�C�!����BF:Z���  ᔟS�7�6Y"<��H�����!@�(�ʒ9�Ů��t]u`�K�9�Mu# ��]��p۷�<��bx/b�%1)`���L��}�5{����	��Q2���7v^��~��oY��
�+Ew2���k�O ��ի�}�Tw�X�T�'G	jJ����ŮUӞ�@D^/���\θƃe��ǎ D�amMA��i��r����|\gĊ?�;�ޢ2�����
�"�Abfr
\�T16�{	Ɔ�M5�v�sI�V��p*��VR*%r���<'M�û��<�/�?>ܒu�Hg�'�@Š6b�{l6�.���r��]N��������`)m��F�B�v����4��t�g�< t�u�Ҧ�5��VC�y"��!T7��c	�h�Fb��m��ro����nOmev i0Sӥ����ig��>�[�b0g3��ս1�+p0�=i�tb�/'�e0;k�v�c'89�	����
K�y�f�A/S
�j��6�I-��=bh����i�_;�w�Cr8tl����@m!�g�;^k�&įz��9P��ƖkN��
άƤG�>��eDm��0J�mt!�B�Ѵ������e>	��m��R��m�s��`�t���k,g���@k;,z^�%�<c�߉��ΰ�V�f�{lXo5���pF@���^Ӕ�����Μ�d��yQ{&����D�\�]�����G�sep��,>�Y|�����[S�c�F��7۱r^����	�"�&IHSG��=:�(��:RZ�^c|���gU-��8R�=�{o (���vjg+:�%�Opu6Oa��F�sH0x�G�gh���i��q��ư�s�- ��;�u�{�<\dm�@n��Ӕ�؅14��C:�+�k����=�<�ynw~���gs���h�<l��.��aI��fحa7u��`'�	� �z5�Lѐ���EG�}R��)Q��q�cm��8WP�jp�7�6�2!�*��3�pE�[ޞ`R8чh��*�X��p|���D���x<c2�Ņ�~�s���	Pϙ-H�睊m�]��E.+lfl_ɉ���߅�
ܾ�N@�X���Ar�v4&�+�CGegL����ҙ��Czw���s����EG��S{�M ��c�8�
Z�S8S{��D�.:NAt�왽Dkq�ڢ?�y�q��Ђ��hfTA\������z��} zq�ۥ��`���#xP-7�<�K���RQ����ݚ��5��gO-P{gb�
j�w� &D^{�n��ݛ�6zR�G��I����|�2Q��޳��G�w�Cye��.����#��6f�*�� V�F��O6k��Y�� �c�+d+�I����f���O�Z9�!d��%q,@y��Y�NtJ[�tnd���`&YES�K���s�c_�]-??�L�t�³?x�Ā�i�����Uk~��d ��re����ؙ3�Yo���f��:g��F�y���]rx`<C��5
8'UD%d]m���G��Y��Vv/^�|A�m@�o��c=�7��m�R��f�-��k
x��>��'��R~^��ʰ�օ��G�}��"N黧�l�����|���EfC�|!Pq䜽g���cq�{���.��,����<)]�����o����\u���\���i��_S�\�=P,c��.~�yϵ��g��`������Zac���IH�ЊBEh�ݜ�W�kՎh����`Y�c3+,��1������fN)4��1�K�˰�(\ ��z� �&z,g�N2W�� #�t��:GL^u$��b���o
�ә�A��Bł<'�nX���KE�X'�FC�����!�[�R���E8��d`%��y޾��
ﯯ���k�.X��ur�� ������;	sv%( ]_���c��k
<�;���;�����ߝYjf'�p�b�l�P�U��;L4�.��`�rŝ��`-����9�%����3ŭt�@���!Ơ�i��&��G,�?��Pи�u���)�;��i܋�ܹ��C�
>G���LF튆	�7�A��C�J���Q[��2�������V"�����D��\��Cv�t"���g��;�A���Tf����0Ikm!7)2�w*p��K6AM�_u�~�R�P���5v���7:����"p�G�g���}R�")�s�E~P�C���И���0qS�&	������9��w;I����������
Hh߉��,�N�����Y������[�ZP=x��B�x
���U5�#R���x�Ȝ�-υ}��$SLWf�3�W��m�/}'�o�,nB��sr.=��"�7r���y�H�A.CR�b�%B��8e������`2��a�
ꨙSb$С���!��ކ�r|���lA��]���넳�;���s&�91�xr��b sz��{�o�������U�_[LΖ+����:��̦����͵�O5�-a9L%X/?7�.�(7=�vE���s���'g�4����f_ǃU�.�"���7�Lho^���&�����vq�;�(<,��cN�/����H����JL���aaA��s���w��0��sk�򖨁@����|�X$�s�$�`~<�1i�.��^��E��b�-�����\�<�t��F���v���}ꅍ��r.s�@� )�j;;��B�#u�dGVĽ���U��{>�l����l�,.6�`�n�D�b�i�
{t��	~�L�q� �m��{wt��c��PMB\�e�œv�h*��R*�X\@i$�m2�BL��O]舼Ԙ�T��r�tk�;�'�{�	� �\y���*A��4��ܒވ{�k�Z�c�"��k������w ήܳ=p�+4N�1b�B����9H�7a��@�A A��/W�������$��p��kEY@�̪n�l(±�ހ���}��ड�ڕ��`���� �v/��c���&[w�Q��0�(pl��]�R�"��s�2�Ŵ�EO�Ag���5�m��h-������sd�3�'���NT/n>W��^����o���ׯ/{�3�	�o,���5�V���=9`Ӱ����M�.�n@Sǡz�]L}nA����7�����ү��cn�c�W��׀X��TƉ�;�-S��� /�f?�B8�3m���1O���qVL}��8�W�l6��2L{��=$%�U̞��I*���� ���_xUI�M�B�v�݊�1@	�ߌm��M������&L�l��.�u`[�:]k�Z���L֤��%{_k��g��t����E�-�-@[�'�>���d��� Q|  ���￻�!�x�5/�0�n�V�ȄR�C#[� �춲����+�F=����k�綋�]8$�>�����8��u,@��=i	���k���KM�ouo�1:�˩  j��x}q)�.><<����p����9�\�[����a�c��_^H������q����s��m�,k߮�N�<��P��sk/�5L�?T Y莌�u:��b�Pu��������ZF�?��!�?w�/U��o�~���6굙�+`�Κ�Ǫ���ye�p{bG *wt:��s�־���l!�A�K��(^so4`��-��m��<��P41�݆ p#LN�&�@b��M..8��^�H|�gKZ���5m�ZO���l��f9/�%?G�e�W �,���׏*BRv yc7���5Tu�\�^:XC1!a� �i�DH�C���#������	v�in�xF2҇�e�X�+b7�خF�u�W<���� )3XK�$P�.�I8�"��U�i�m�G�y��e���?#ۧ�&;a��>���P��}q����2�ڼJ����y�|ou$&C�w��Rv��Z�t��@��^鐓�]
���m[�9���=g�6M��s�씣p��&��B��L^*<�BJ<��W��dD��9���]}8�s��H9��k����s��~�

��74�n��[	�, +�S��o�o҆-X!����F��C��Q�����(΋��C��%��Ph���@@
���-Mf�i=N�@p(��R�ʠ�s�~�cp�z��>����b	c�� $ދk	H�f���)tKiPrUz����{~qɞN ���E�+��T|�� @�fG�%��"�/���f�D^�T�%}]pE{UUa�O{s�I�̀j�}W���Z.b��:� �{��Ӄ�2��/��8�p ��@׎�B�s����=�lˋ�� �`�U�fI����1�D�=$�:���Z�`�����k[�����
��L��!��j$�U�ks��Y5N�5���`��o_�&��`�Z�\(Fs�(z
Se��I�������w��<�Dx^Ȁ3֔�ֹx�����q�UGi&6����)��� �S� wë��t阝R~�F����'�U�������Ѐ���
�>?�:���H�e�cy!9g]?J8���ź�G�ol�{�ꉄ��g4p���<M�$��A���4�Cӎ�
�8+-#-�#��t<l���M���s��z��x��t� �P�}��05S��]���o���R�o�e���	��5�@�il�>����JbC:�i����שj�2���H� �?�������,%Dkb?���Z�����#�L 2J������9�E���mv����Y9`]Y�pジ���\���ߏb�4R�`���m�p�
ShwbkI���[��T�V[�e�����s�S�3�0= ���8��u=��B�?�ۋ;�i&2@hS���k���`�zRu�Da\z�V7V�-I���W���7,Fk�Q|ɸ�6�������5�[���ak8b%��oo���O_�}��x�1ʸ	�uU���ɡ0�tL0�]!]!��l��j@@�0~&��h]LE�ҵ���7am����ċw�
�{�P�Rꧩ�B�>fcɓjK�ک�����n��;o�������F�!����y��v�E�h��@:�lB,ǧ�>w���D��u��ˎ,#����� Y��\F������Sl&q�N{�����G��d�G���@^���*�%6d$1s�� a������`l���.
4�+��G�B�M�f�����.a,�x�Θ�y��ߢ๛�Fg�� By�<L�<6G�@�:7�C��,��?1���?�%|����0�j��
�19��.y�z�i���i(ס+���#��1�8�v�� 3��(P�@���F9���X*�a�i���L��s���ǲ
��Y���g���4q� ������� K�X�5�G$�IY��'�����N���*|��`���U������n�ͧ�1�d�OL��0B�dK�zsq��C��̎��HK<�~�c�6U��\���/�]UX�h�?�A;�����~�_���7�� �'Ѕ��k2
�y�Qe��F�#�V� {�C7��� �M&ؤDt2%&η7_��m>�����uH����pssn�ܑ�́gN�P`U�1�CM�P/u�>}������	��q�B�!�ʨ�^�3N�-�X�;�d0�������Ȑ��;��ʠ@�@�����p͉ȏ;�B	`�B�t����n$�`(�`�L#�����9t�k�`�Cwyr���Ƿ�x�؇˳�8��$�Ŝ��7��A��@@�6��z.2�������x]�9����Q���J�+	�������TW����4�?����*�+�c^��&�)����y� �;���D���?�d�E��i��oG&Η/7�����~|�Em8�P���|����C��=ZϏ����������{��xG��i�U0Lƺ_�
�0c�����=l�kE��x������u1���5�.�v&���j��&1���F �˒0��5�����Ꞃ� ���8�I�m����}��]�k�E [o:W���I�` @�g��Fg)��e<V��hB!9 o�E���5��vG�ګ�f��y���%񴄮�-��=��臮�O���т�h���=��d�\:��$i>��W7�8f;[�?T}�t�96|lִx�?��%D�2�y��{�����g �ֶ-3'�x?<�x��.�����|m����'�ڎ��1�tYbhA��*e==�[Og�ײ��k4�NtfdQc�xnu>�q뛷H:���,���b���˔@�|G�Rl z����޾>GW��Ak#�ǂ��M
��Um�ͣR�v��L�'�~�9��6C0��.��� �48BQ/.��� �K����%����� H
`���<�s���J� �����kbC��.�j��$dk6�j1�Kk	�53I]x���N����g~/� a�0�`�b]_����k:�ď:}�2��A��f��<�Cx�A��l~��Õ	k�C\�^k�~D�9\�Vj%^Ď��K�מ,@wc��hšd�¢�=�A[J�����fs��������r'����6��g]p-�{0[��d����h��J���{��G v�c6���>����A�K`Oy�`�F��|���<�k�_���7�l�P�X���8�*����'i�\Jd��Ӝ���(|�7�����KG����3�1H���� �zkqc�����a:c�֛+�q���x�Fmq(��}�-i+����t���<��V`N,�Kk�Nds�S����I�b���3�D�,ڭ��Һ�8?�%���+����Co�jrƣ�t�g�xm�:���յD�Nl���J-V�L���1+:oU���։NM5,�Lq�iG�9���7�0��(�Ĝ�}�H���Me]�ƕ�+o+�U��&�?�������»�w�*����.���wa�\L��ښ0f��C�����<ǌ�E� �ǧ�f|��	�G���Y�(HZ5�c0�Q����iI0?���<Y~C��b&��&dP-�
h��2aĺ�b7t6�ܺ}�I�BslN�J�<�8�/��ƽ9�� Gdڡ�l
�p �H��:�G#T�D�mL_�1�zoX����/��uNp����G� dz&="Q짣�{[���^�]��}�m6�gY��v
��>,�7"fI�P|��֠�܈Xk��!1B>�m�� :�W�D _��ɕ,	G3	��x��0�-א�jz��!�`_K��Ahql�ZK�vs�!����,����;��o?T�Ԟ!l�813q��.jq%v���[��0w,ֲ��G�]a��ٟ<H�ZL&����QUIwf(��G��pN�g?o2�c�ۚ�/R�jXf���:��j����i�̊�2�_���?�Դ*��졤��?�֣�ϟ�����4 79�zܐ�!�,%`��O�U9��'AgQұ�d�&ydi������ z�IYϋ6��x� Z�1go��!�������cK���l�]A�_��_»���i�@	 ��-[��(䈅�2����Z����b�����C����'&�E׈�y�֏b~��G���~���t_��*��������?��	W�ˡ�^�d���`�s�����W<3R���ϝ�0TR)���~/�w����įj��gF��������^��v�=�sF����)���c���dc� k���|�����pi�M�W!���ZA�n����o���t��-ǙXl�ڴOѴ��ND��Ma_��(yC��Q��$�����ߘ$ү�6�R	'�{P�^��
����X��՛�c��-e�v�g;����������)�l��O���@�d>�.�����^B����|9>~����V�]ף}���c̫B^��ʴ�%^m��}��1�5�V��c,���g��{���( .d��
�������B8b��K/�k{�o]����m��6қ(�Irӂ;�GvʿS�њ%x�I�؝i��mj�6��IZ� ���Ns����vd�"!�&��~�>��3��8C�cl���\��0U������C4=BͧՅr�5B�����
��u��+ڽ	��C$G0��D��_��j$(� ̚���I�#�MG���6�qY\�gp���:�U�	X����9�Y��Ăz}��~����[�Ua)h=d�K�měC^��|�qK��`�\	8���t���9Yգ�V�a�����i�Qx*-�gg�p������{h9�$W��P���z�C�}��I���=ܥvwU
$t�?���=HQ-f�dt��B�4m�u��y_�`�3������یf ��c��i�S���d�}f9|cƘ�j�����s���!�,^���J%5I�\U�k��ۅ�1�y�����֫|�"=u�~�U��z��K�$�zk
Ɠ#V_�����Y��� ̞H��D��'�'�ʂVմ?�>�3���&��
|���6x$�d"��Q<(w}sé,����9jZ�k;��+��ը~�øq�e���e�=G�i�Eaw*F��-�{��vM%:-�1C�הmQ�nPҫbA��t��h�Q4�s4���~���ߙ�~����9����=-g�{b���[�/07���^�� �\����-ɷX'�?����Y��)�;�
0�_������bf#�^%�e�X.T�.9��@x�Q�� ���G�
���Vݛ���9
r<UV���n�=�Nz���B��g��љi��\,E�h�c�¨V3���y%cE�RB��1KN\fK�gjd!UQ�p�V,e�`���WYz^mӵ{>�A�8%Z^����_d^ yy8���A�&��ػ| b�������+�a�"��=�5��G�_o�I��.��R)�x��nb%�)k2�����Jp�s����#�VJ�Q/�^
�?�s�]0���S� Ex+ʱ�2�05��!�#�H�j=R ��M�=R���⿆�A��d�]6���3�I`!���z�v`L�ػre��5���g4b�Aaɝ(�#gb���U��CD�.��˸K��2;�|<%	d�O�$FFJ��C#F3&r��U�4$@��D2����AX��v\R]�+���ۖ����(F��G@a�F�D�!D��j�ZGj �')�j�T0N!�T�G�\�(����o���W�E�x����y��<��T�Yxa�Ϩ���O_�uy�B�=$ax()���ɀ�a�����(9� �~d�,�G}H׮�1�aI��s��~�!��H,�
��z����n�*X��|p�"�F1PeP�����i)jr�"B��˾�K�TV�J%���_E#���Y1��J����Po|���}G8��m�2X�]#��Y��i��\�f���r�����[��z�0����~3�	����m�V���]Y�F��=>���1d^Z�=k0�RF�)�������F�,�Q�[�1��{���#W;��k.� �G�r*�a/E 4�2�����T��M
�S�Ä��U���e�z���g���h��HE�M��1�,	�Tm��(.5��'^��O���ZE&\d��1Ӹ �T�A�VMh��f��Pz�m#|�����<<�2` jfZ�A\<�cy�H�Ft�t��Β��R��a�W��r:4�3%LԈ������7�N+�Nm�����h�84He�N�w0ǝa/��E��p�������,���j[�$`��2Ge�)"g/���,g��P��.G"�e-�GG{��G͙�q��n������sDk
��M';�.�x+r�n!㴌Gx�ױ!/4��BG��a�2⬕��^|b`�X�z��h�2�T����^䄣�!��#��W;���GzW��8�gy!rj']:U�m.�j���r��;�a�\<c���$\y��2.���Uk�L�_�-ŗ~x�jNY�����  �Mtca%6�h�e7�[
��)�,��a,Tg�V�ca"J�xt�O.���)1�k��"r�D��0����c���֕�T��E9�.uOm#����˕lwb�g�r���Ma��曻;ZΖ\ɬ�^9F�puKA���<��O?p�N$�
Ɲ���D���M�?~��$�Hno��������C(2>`���{���zC���~<8*�Q�1;m���y��|S��<s�F3�0�jؑI5 2�4��]?ڄ���Vl��&�17SE��`i�Y!�ef���.T�P�qF:G��05�=i�9��d���g�N|K���E'���1mD��A+�44K�[յG{'��)H�
j2l�=, ��F����Gd/`��`�WD uE�Ð�?fu<h����1�g�~O�z��D!�4�z�)�<xʈ���H��k�T9������r%�Q,Z��t}r�b�s#��B�yi��qP� ��QCS����WF����EY���3�1����(��ew���#�1��zS?��qP�U6���8?�-��.�`�R�L*d5[����-�s^?G%�0L� v�c|�x�� �!� �!���
;��� ���ׯd���g`���k4&(+.Q�Ѩa��a�|X���/��9��~i���q�(3�D\� k�h ���� ��O{ d�O���vN�iο`c��<u$@o�)��J*H#X}@�]���+�K']�Ps������2@�RɭZ-_�H�℘q]i����R�)�������T4P���e��)^��e�瀞�s��ve6��-�~���Ө���9#��k�tk����_�����<��<]c�A"���>��ߋ���'_#�ڊ�mkld�z'�����W��!�3�U�y�͌�!FY�V�)���N<y;?4�,����#��="W�k�W�Z�Y*�s$��p�ѩ��T�,vĨL���_菌�7cp����n�C����踨`�]�$���	�6j�^�T�Ã1�.��T��b, )��|�y�IpC�^���Ɯ�J*���Ѩ[���4'|/�BW$Q�R `���@� "t�#����ӝ8c�yĉT��x���@�Q������/��O�	���sZ.~I���Y�D�b�9j�XFvH^�5W3�}`8�L�vvb��l{O��T��樆��($����>~��2�?�㏁p=e^+G��Tn>H�;*l`�H���j�DU0�n���9&c$���N_\M1JD�dl��hcsa�j�C$��&wL9:
��%�*�Qp6{�ek4��掍a����x1�# :����B��$���p�mΌ�B�29LZ�Ӳ
��/x�ڛ��l�9{������b���2r;�vN�J���5AoT��J��P�te��0��B	4�8�^����y3Q3��h!�k$�A�,0� �K�z�����Z����2n؀�������Fg�����?|�D�n>҇�-ub��|}qIX�;v�����4��K��vyũ�KDw�6t��ֻ�[�A����uCp�`���	�{y�tc����}����OTX�l�B�Y%����	�;̰a�\d��T~Ua�j�"~ -��1X�v{d����j<�ߤ�{��hR���x Bi�5̐8���%�ٍ�#�&�g/T�m�!w%�M�Ŀ:s���T?�2�!�M��D�Q'�CYpy�pi2�}���yY�d�r�qh�j�Ī��kT�0�0h�<$3+N��R帇U�A��QrI{M������gnU)�s-Q6Y1E��h�Z.+��ID.z�;���n�ʨ���ɿD�z�HЩ�wA,c�s��@{��Һ��[��� ��Q��x����V�L�A�z�@���P���&�I{-wV@!��^;��e�� &�/�/@P,xt"|-��+����0A~�a�P�T!h�}4#`$��5$����7 {�8�����
���s4@gS���XZƛ	���A*J�8��n��!���1�-\Z3Z�E���h(!��/��g#���wAB��M��-/V·E*T�L�E�ا� "��<�f�1�[+����3	�}����p���fo"鲰#
�#5�Q*�I��8UQm0��J��5�[V���D�0���=d����N+�.��dʶ?7�\�k_��E�y�U�g}�B�+����v�=�&J|�sT������ϣ�^���*��|���כ��������V)Ƭ1����s�Gm��&	i��9�Nq�Z��?�r������0�P��\��\�W(�0�M���5{5!Hsj�lH;z�J4mφp6���IGd�0>/x0D�i0I����~��'>�
��#F��mE�s�����s(ը������Qm@��)�i\�� ��~m�\���6�`�h��� {!�f�J=�'q�ʶ�۹F_0fbDe#���-�^�K�G���u���ȲR{��9u78�P��\��<O��v�f9���ۊ��"���R�$�C���mb�pP�f�æ�"�hq]jϴ�to8�0���<��X��k��'�8��c�c�#5����Y���.)t8m	�538"�@<�G.�p��-CY';^뵤�o�#FI`q0�2�Y�����0c�G��^�v����C�9���Z����ǆ#�w�.��5$��v]�Q�.v�0n�b��Ǆ�Ep0>�I��[��$��i��ݬa��&A�F�
;��Ҕ#���(T��!�B�͖ZXG V�H_6�9�8C58Ed����/yI_&��uJٸw<�~�R�����,ʺ����W��p}��=�� 	 ���t)}��(����Y�H]=�Y!���f?�hD9�/f��,�������<�.$rҰ�����C��aZ��߉A@R�%jՉ�|�L������#Q�'��?�im-�9���`���|l�a@��.�j�4-���h��N#��!E8�IL��9R��=����8]݁۽�c�
.�t�?p��:)�*U�������x%b��`_JT4��W��#�UF~h ��V��=���uL,�����L�h�
�y���a��Z�f����WOj��p����u��}�K��B18�bwY�X�9۱p�+���y�ԂU���cTp�ڸs��s�?����%�eʳ�!�X��L��z����]��ЫPQ�{���rc����j��O��gYkCS�7�	��PJ�c��p�J�������o�y^�!��b9�Z��#4T�tQFj]9#@!�Ō��y��|g�x:O&j��|%��c"��\�ܘ�a#�Ήa�#1���	Q�+����9c�Eĉ׆ۨ�>��,:i��4��� U�z5bI��٩@¸��k�&��`�$���ic�CK&�k�U�m&�K�I���f�j0x�=4���Tj!�M�G�؋�=�n�'ϥm�K�rT��sIho�4|<j�� BG��E�gjZO������8:^���C2�_ܸ�VC16�ܖ��N'�>��!��w�.�j%���Nq{f����܂Q��QܜB1J�G�L��h�(.n`(i�����RMI'��Rp�}������P�e�{A��7���g��=�x��c�'��<���k��c�̣RxB���:���g�����+��-n�_���F�3�����s�\E��έ�	��7bv���2Q%]i"�c����Fxj���$���x���WE	1��TX�>�K�1`���p�@�x��p�(� �M�bs����Z��(\ITr��`:�F
�2"Pv\�p��z���Ǎ����i��XbVb	�i=	���|�?:�
���&��#K�������w�
�ۚ���Ŏ�;R�
bH�/<�lD��k�oI����)��q=�z��B�������BS���B�}�-4�u�b���b�0� .����U)U��U�DY�a9o� �;�s&S�G$2�gg$��z'ц=M�`,i,�a0Rq�zO��F4
A��C`cΞ!+�����0T��KK�#�/��gN��"X{��h�5R�s?�>˺�L��s6p�k��[w��p�W�2�a6l�����d#)t��4�#�cP׫|���[�G��,[�QG�k���g�vl@��@�@E(��;℟��Fa�]�߁ǝ��f7g�F����W,w[уXQ�7��R9����iՅ4jߪ�fe�}�(/�Ɣ�\ax�t�{�eQy��X���C�F4?���}���l��Լ�f�M�s���JrU�Q��n������Ւ���������{��3��`�aݿAd��u2�U�~����O>�w�����a¤Y�G�1h�Ӳp��rɘ;x5�,k�Uf�Ha�?
TI$�������6��y��t3D�3�s�є�ĳ�i���O�9#���1�X�1�#v�>�dƙ�b�Fo����o���+�?@a�5�إI��dP{���ܡBO�*>
�L�==�2��5�<����0�-R<�l''�?*��F��]^��X�{f��I+c����<����[��	�,8K�i4j���F(���#�qfl� жs��HD������򆛵5h�Gj�8�B{�2��R�icpEOXsM�ǲ4 p%q���5�2a�c�B}���餚���+��g�3��J"�����׌�]Z1�p���O�o������/G��L��*�֡�5�'K9����(�2�b��|~xHx��M7Ĺ�q��n-�:��*�&&��a`��zɓfR����2�VjT����T�^��kq�#�H�
C'�	��I�Tj��zA�A�ZƎ�h"/��~0f)
��Y�P+�*�A�h���dcS��!QWb��֚���z��[S�����h Æ`�Cө,�K""sU0�2��<<�0�����vy}�g@�\��2M6̖�E8�����d��0xweX��J���7�d��F �C�}��}|�Q��w����w��u��۶�Oe���SC����ʹu�52Dx�,r6����N�������) �0���uǘ}4��h��QӣD�i���"�2�փV��p���� ����!����>�����`�%G(t��J���;拇}�,0nO7�w[�b��ıfX��*Q����\�`���qo��b��Š6I��p�d���laB8��("R8b��Pҗ�r�S{� �����W�Ih�@052�f�	d�5��pT\�^Ҹ�Nҟ�f+id��VW���ʍDY��}��{M��⪞�Y'�
�1 �J�I���# ,�t\0"��7md��L�権g�btT�IK�£`���T#��f�>3��.��6i�Η�jM��L�X3����:df�}8q`�q<>j�P%r	g��:��k���}��½a��~�ÛSx�:t0IJ^ۮ�bߩ�eǆS��X�(��T5DUA�C��8횜�6�8F[2���1��X��D����q�+�0�n�;�C����YfmQ)8ĩ*%�okD�H�/W�ô6�x����:���Χ�6�MT���pυJ��D�Ӛa<&*�B�,y�T���ZL��=vυU��3�N�������k���W'ߓ$�Ǵ����8�U^�5�Ӣ)����I��
���*�R|*j�DVOU7��o����0����� ݂A'����6+�4�4
TM� �� u��2 �X=5�����_Z�Aʁ"�dwo��&m��#�Ѹ��;��2���D��ܦ��&��D�b|
8m�|Q�!�"Hœ8�ɛX\J4s���nմ�zl?�TS?����K��I�H��k}��;rTmK� ��1��<���~f�RiM��6dFAI�3Xj��W#�W<ǖ]T�+��QË=f#�0�[�z���(��N�&t4���`Ԓ�&h��WF��
�](�G��%�Ӕ�|���n���
^��"9�V�F�iɫ�w-�mU<̨�_*��1Y[{�,�����<?2��y%F4�O����࿆���[;��4ה�V-��=iܠ����Giy4��l�y�-��oclQH����R�
z`��� 2�C�{�	��p��R�rĎ4�sA�j9�����2��D��lA�ƌL2O�V%�����;�h�	�Je�jؙ�!-c�c��e��q,���=#F�&�%g%��?�ը�T���R�����)�K�_�%���1�N,��F�.&ۻ���.�HÔ!k�9jE|X�B�������%���/�@#c�ΣP���g������O-�5��~�ȹƽ6@��'m��ŗƒt=���6ƵaG�}q-����ܼ�^���6:��T�.�\
q��_��k�����!�#�H���9���S��;����\p �7ϒ� ��9R��i���9X+Gg��I
jGV6�1�`�I�$�/��Q%����
�%����<��P�Ƅ�3��ȸY��h��A/ֆE5��ˣr)G��RN�2����S��,��r��X�v��يҭcg�&hJv��&$K~�P����Ж�/2���`�*?��[�+ �V8b�`��F�]�gg��%ܔyM�'"K��"��Q��E<�FWw�	�W�Њ��c δT}�Z����5�V��F)vѡ�2�b�kɊ] ����
�{6�I寃���S_DI�5�=紶'6�p� �U�8�S�xF�\�DI*x`#R����z��O�:� �N��`�H�(F$���jò�&]'UC��)�u���ꧨP*�z��],�"��?�>#�Q�!�~��|1���d�2��6���0�;fP���(����#�~Vг��ƃ�d��#R��r�c�4d ���k���.�#?�<�dk=!��",�N�bؙM%�x���z�������A�Aѳ�hH��a�ա!D�S�@�#��߳���Zp
*�w�g!
���7t7�-*�Ew59h5������&HG&�s��%;�9[�P�]��fX�(��(W�j�j?�qY
�pU����׸�P�
�B��ݚ��-�؏�_?��?�X?�#�3�qX����L�OD�-�dr�S�@�|[Lt�탁Fn������ W��C�چ�7K:�� �d�O�����\��^�%_��Imp\�
Q�+A�Z(G_�do�0��,lilА����XO]����R3o�e)���/
p�0K����`hʖ�]	C�ZB�T(�H,OT�X5�ћ����r���(֋~e��!�43F��?E���Xf'�r:p��`a
�����ө@`ϵ�)ySp[�݀��Dj8皅lb�1��vҸ���:5T��+�3�,����\lT���6zhu^�jQ%��(�3�{T���1,!���;/�%<z�t��c���T����e�N8�K6��6�7.�R��eaL��G��\�����6пŢ�ƛj�
9�������i��mӪ0k�& ��s��Z���"�Jc`�c����TGX�W��k�j�iōt�<�Nk����h4J+����L�!�Ky٩T�u�%i��HŅ:�#:}�����f��aA�L�v�qA��W�o �ՠ\��̼c�ҭ�D����}�m�qG�uoI89*]R.g�-:�!oopPa�V�� �JO�|Rl��?�g�������`L_Tu��s乕["o���z���mB���Pݴ^��ܱ�4��|8}?�M%m�X�*ϴ���fm3�o-K�i,:gG��2v�h�э�FC�w9��B4*a;���˅���\d�_��d�1�� ��Fiq�q�,�u}N��)�"/�}�2�1�k�8�b@�{�����̙� ���ʘ.lx8dޣN	�Q�(	���@t��;�o���E�reCuN]�L��Ե%���Rv-U�	�f�/���L���dҳ���Ǫt����ee�e#�̠^e`D�F�J�A�mZM�C�E3���mN��
�D�z�4o�?����|b,�(�S=*[�=G>i�H|�Q�=�+�.SW�n�vG�ق�'%�����SÀ�(�M�:V��t�z$���H1�Z��#u��O�r�DC�j�����CS�%:A�e�e�u��l�SC���Y���Y��Ձ0�0���0�ɪ%I�p�،.��u>�F7`�:0�(�q	���QeziG���.�4Q
��3����g�BT�],�bX�Ho�@#�i�c�+�:v���4�Yk6Ĕ&����Ht��Tͤ��?'e��W$�g\�B7IƛTZC��.(oȬE[c=���O�y�����Z;�c-���'l���uⲄ�kgv1����������U���V��B��8�U1�����*>�x'Xh��{��j�L��V��P��)�"�Wh��~��G�<�i�n��%i�~����ݞ.�K6�aN�E�_D�!�y���h~y��ROO���~���n2��}H�sl��-��R��l��N���a�F���1�C���&�9)&�Xk1�-{a���lGd��䱌:���hŞ�=�=�]�vNE��Dy���y��|I�v�a�m\VGͼ�	�D���r{�)�3���s��_%ps�]X)�;�w�����ƭ<��ʝ��@��Ȅ,d��jcĥ������qXy@7�(�,�|Ǯ���Bqhu���C�]HM+i
O�=BX��Xlr^S�<mSU~3#J�^6���r�X�\�|�`�􆷢���Q���(� ��hiU��FKU*5�F�͓�5!�w�lu&��պ@��N�
�?d��J4T]�L��y����c�I��P�F	i���pS2_IZ����^�ymk��y*S�XYvr��x,$k&�?��I�Sy�7F������,�'�ѳ�C.��Z�I�^��z��*B���R1�´�T1y���*c�JU��U�B�m-��((8���d� U�L�ר����L7�a��@�`�B�'մ��$:���f�F����k6�x N����\�|�2��k��o9jI�v\��q�C������ѷ��D[�A;�!���5�P5�q�w�oa@�(��Z��	/�>��������mu�
<�6"�udƝ���|N�؀���g�hB�o�Ɓ��i�Ҽ���}k����(���#�|
���]��:�B�5_���)����iU�*��OFK�V�R�/x['���FS�:��ﵖz�cem>�̲�P����nh�V<@ӝېƍ8�D Q9��+y�=�G=	�B*�Q�Oco�0&����Hq	sb���n�~�E����H��v5�27�k��>g��Cpe��cN����:a�-��|��Nmc�-"�+C6�ktl�-�Y��}Gr9�;��N0�6��Q�mcARr��F:�Uvt<n��V�Gڒ��ͱI�
O�<3bX904����$j��T���-�_�y���bš,�?[WGU굢����>e����Iՙ�U�Y�2?v��PۙFL�
Î��s���8�OsĠɼ�w�=��"�}��m�]���KO���,�V�p9�~x)��{1:m�9��9~�0����v��N��ШS5G�sό�hr�`�X ǿ1p��%p <�(C�cV)�B����nvw���\i7��,�h�>�x��;��TֻV{�,��y�����=p��=��F��(�^_f�]ޥ5�h����g�����(�����5}n�06�>��E���+jg��ڭ���ot�z�U��>C���cmP���)h
�L�Ɵ�8�:^f�y�F1v������6�!�Ԫ�`c�2��zM�'Z,�hqqE��0�\$e�:5tI�YG���Ƞd��n!���<�K8�	�����z�T9c�d!WF��7kN ����`e���"������(:=ׅ���3ej�[�3��1zDB9wM�L<[��B,	���jI0�h�D�ȋs��Y5l�m$��nX�Lj�Q'zd�
= �jQ�!-7���N� ���<	�����b�Ze0-�/���Y��O��`����ܩV�@�R�V+@G[iׄ��Q,�c�0��n)W5*��
�<^V%+YƐ����������O�ߕD����Yf�k{TJ�Ҭʶ;�V�2��4a�f�^��~�5N��5G��U�"%�M!�>�H[2�6"�������{D��n0�����k�F�J]���|�X�;��T�]�I�~Þ�F�B����Kkv�ӵ$��
!��J��xo>�����-S�^�;���?��;7�~Sή�0e(��F�_����qyg�����7u��4�I_!;(�W4b����׾��@`J����T�ΜQ��^�]�ee��DsD�e��C)�ŏa�
#�����\T�zQR�'�Y!RcI�"��Tq����觮`
Ц�,n�@�J�o�z�xG:�����y��؊��*�ձS�6D߄�E�֡?#��HW�C��6n(^P=�::j4�F��0r_��>��f��h�GqR�
�>֮W>A�p���6�ՠ{#J�H1��<���\�[0���tq�r�@l�2�9�
j��i\��?ik��v��Ϊl�n�T�3��Ə�%雾q�b�d��ʜ|g��9�����'ZE�Σ�y���/�r0JC�k��v��޾�K�f��SY3$��!��X�S�)��{1
!�mRܰJh��0N�^e�k�C�me�?)e��>��~�����ӫ��8R�#�ɜ�6pl5j��0����������ߜ�ĸ��S�����{^�Ǵ`'3Z\_�y�h��#ox6дH�`|��1j��n�x5�V��O��i��+���Z������	 �ݶ�h��	~">�>���5=v�������6ѮY�1��?�!��y����+�����wt���>"���iņ����|I<�G6x�..�n0f��C�u�c�����M5성/F�J�4�	́sq�.����k������M��:��4�4'�Ԁ=u���[�ǌ$�*��LIRc���-��*�@V��@�/=![�2�9���a�D�
K�|߬��ݚV[У��a�\�p���QA�1�}��eeɈ��nxj�_h��
Uڧ&�ԍ#QC����c(�^�jc�y�1ڑ�'����WcW�h9s:�h
MSlL�h��/��aXj�W:
�%�O�
����YtǉvH�
�"G���G~!g���[&Fs9G���,�
}<�&l�`dQM<�Y�E]���Hi�?��}5W?�@��cx�pM��������^7֐�����b]�%��9NRt��C�������/������^�>3�^�*@D�~��fe"r�o�E����PL6-ـ�m
��~����<����acT+x���+�28i�0ߝ���865e?��52���#��Uy���#��=o�fz��J= g:{F/��-�W�<���݂�M��_�%�%����ƻ"Z���ǐ��Y���>�L�
#��sδ�E��=ֲBU>�����)�X�0TL
�A�JY'�A����Q�|�l��ߝ+�""I�7�V��:8���a����M� Q����s�l\�#`FIk��$5'G���/�-0Q��[��h���b�@��_���ۉ�0�W�Ρ����g��������a�:W��:���*�Z@��L�n�N�` ���Ǎ�"��ʦWO0r�?�q�m�2��Q�T����htK�Z�=�F<��c����F�H�vYX��/���lG�-��S�m���s�Ǎ�;�^���>W�M�&�rzIr?��}W����yu��Og��>K�`+:\�� ϭ/�����#I4�P�*;�ީ9�ҿ����5����*���޶�4�I�>��=�1O�D*�������7�gAz�z�LO�����
p8��"J��h�{�c��p`�|[=���W���bZp4K?�(٧I�l�2 ��	�He�tGN�����W ����+���y���(<��^1v�X�*��Q}H�u�4	���F�Q��[��:LJ�(5������;e��e�g�*͖�gx,Q+{�x��*։�PЁ�
����z�@m�����L�f�����,i�^�I���|��s/���!�Q����Q�O��}5Q*��'��1��~).�PqO2O��=
�	%�3��>���]{�M+�F��{S�O�0��X,!fa��$y֍���H
�Ss$���z|#���;��=��ʑ'��O��j�.�s���f<e�>p�\��ł���!@Ix�Q)�;vj\�32c��[�{�f��#z�vRe}��|,�8"����� �!����]p	>ƌ�r��S�	@!{��C:�<O���xS�-Jk��6-��ʞ�l�I3 �u�T�:�%�5�X=y���p5��{)$�}�G6À��^&��EHi�7�0�ue#�9�R\e�u�*��}�c���A�1m
��߱�ӍeAS�r|_{Ț�Ө�w�����dÂk�αZ���RZMx��)�ʁ=7�q���˂@40�J��%̊�������
��1���?J!���-f�?���g�$�PN�'Kh}����[��ANr&)��� �ޣ�c�=���S`���w{���ܣ��[k|�bl}i$�/m�g�|.E�����E��$d
���^ӾӴ�F��{ʩ�&�$�rc�&~2�#iZ!��Bu�?%���R���yv����1��ʏέ���)SzI��>���N��irɐxO�TA�ݱ��̫&R6ݕ�B��}��u&�)�F)�ݐٓȞ"�_��Q�d�*OT��:��X��1Mڢb���zI��XY���	�(�yT�՜Puɾ�h���'9<�A*�*\Tϻ�o^:���6����FF�:g5-��)e����r���o8��T��{����BN/����*_˽���ڼB���
�M/���e�ӱpT�T�*�C���,����}}�0�������U��2����W��/����0����2j�c{�#W#m�9��;[�:���*�q��y������M�����~W_��<[�X~�`|M�C%����٠��O�A�:���NABv�aC�㞿�uZ�Q4�-c+�#�~O����/�ן����hLY!Г�'�f��8�P1�}�ώ &~f�����tpUf������)�<�1��:(������i��y1������H��%�/?��b� �w?�<݃��%o�x����w6�>�h�Գ$;`�'����4Mr|��#�A��(@6�p]��3ʟ��/��4��1��A�0�L��㇏�?R�׫4�ω���ѭx���*�����N1�/���=jI;)\��a{�̹�Ύ���ę�H�7�,b@"x��	
�	�oO��	S�Pp�N�@�LAH��$cC>n���T�EiN=Hb}�u~t,`h�H�6OĻsd���K	J+e����s���]\�PD���	-s���g� Y{�8 �?����!����q��ϼf@�G��x�y_�r���A����	�x��5��|mj�`�̦��1tA@[,f2� �e��G� t�4��yK���1��i�0Yv`@	�rMQ��Y�Z�Ρ���
�K���Nz�ON�Wu�)>�������.�'�˩��G�=,Z����!�}��}���|���D�+|оr?��jX�̺��&�rΊ���V��b�v�,�4鯴�¨s2_1���FK������'Wm;j:ls��Q����2����S�5�t��<X����V����wF_b�)��8|K��������^:c-��Σ���e?�۰i�����;�x%��F?X�[y��<b���Ѿ�.�Xˍ �BG��H'+�ί��Z`�(��0zMM)-�6�M���Q�N(�����|_ǂF���+M^	�c��f���q�T,yA��N磋mf�1,(����Rf[<�\�S1����/X���g:m�|/d���3*�Г��`$Q	��R{а��}�O�V�G��;b�^ճq��	��{�P
}��M��Q��8����s���ﺶ;3j�xv��i2�6�cH��Q��E�VP~��ȗ�r^'՚8=����F����Q�m��%m��c�f*ӥ-��(�dǜ?n��q��<�\�/���Ӯ��6ԧ��?����j��a��Q�4��d��eߗ^�Yfc�/s�����?h|��_�S��+dE�W�� ����I&#k�w�LK���nJ�ϖ��m�k������L��Q�`��"]��)���aÆj���E
�W��1�/��;kc��Fa
��5�vjXNژ�}�%oM��T���f�W�q6��ǻ;��_�ag��w}��Jޠ�77�X^���!.L��H������M��sX�&�lM�nHBA�)6Aq����ڄ8���1��./8�m�|��>�K�
��h9��ӇOt}�:�:�ӿ}���KJ�11�>1�e�蒎�����h��c��^e@h�.�X{��)kekM��ǜ
����yڒ�m!x()cw������t����	�]�3��8L���J<T�P�i�aa<jf�#M�E#�5-X�d��;���|H��x^���� �{D�|��s���G~ߠ��j�6j��n'�!��)��ẓ��"X2�VjO�W7A�H^ш�oy���ͻ�L�Ɯ0~6�l��
�<OR�P�m�ֹD-���q���w�7WLh��*눃v�XLӺO}���Y?�!��R��ق�@N��
�|���Q\��0~�,s?����	2�G6��>��*DŤr���0������]'��P�"r�����<v��U�=�K&ЅBAr��.�w�u�����hFzMm�7�R�4�ޑ=�ގ����p~��E1;��|��[�%{���
.]�&(}�%GU��B�&K�[;l��V�� 4�7�D��6	x!��Oki� ��_����*�����t�0"�?�ȊNgN'��HCݭ��ŗ�S^V_СM>r��e	��xm��Bzڇ0�1U[y�D~f[; 2ק�ޓ�HZr7��k8ݻ��fwC:���hD�T c�D�� �-G���N��Ւ� �_]��.)Wv�p3�M��)؏�e�H
�D�	>��m;�� tos��O�"�H��>{�D�w)�e���/�� ��9�̆He�Ũx0�A��c��2�܁��'������
A���x>JeK�X���aƚ���b�~��?<%� &������<�9���n��c �S.p��K�4;5��@N�*d]��"cSv8�x�:���_+�}uဵꕮ]����%���e目��y�T�)E�b,�cDq<{(5�3�/ż<J񗴥�y~��e�N���r%=,L>�h��I�hE<P%�^��]�~����zI��� ���{z^+;l�t�~bU���&���S��'M�v�6���J�O��h�/H�"x�����ū�f��S�B�z5§s0�5�{F��-��^n�[����O��Z�5��!����^e}�Ip��鴼�/��k4�ol{�5���턠�qyuM7�����R��������:)��5�_%&x� �m���Uy!��i{�a�͢>�����,�rU�[2󡰑��1^H7����:x��vJ�

������0R�U����}��V_��
OqKW|ˋ<�Ki���+�R=�=�DEdId��J(����)�����l֦��+j�m&$L�7\Em��LB��k�)@.���cRc��5�n4$O��6A�#�J�"��۵~,����D�6�`��f��2��4].4�O��W���m2��
Jx��1�R� �F�RώE9Q�*,/��X��r���[��>�r����A����_q/\W�Q��[���ճ� P�#�j~��5��14 �~�VC���NGɟ�m)��t`dt�}=����{�*tt��1|-ߩq�/���{�o~��BuZP�A�4�`7W[�{�*��ѣX�ڴ�.����<L�%RVEh ��%��כ��1E���{��C~���b��q�PFz�7GKY;wpQ���o�0T���uD5��^"�m�F�f���$���_|�#98�)�=�gp)�!�W9cl�~�a�ՙ���w��E���8e���>8�'��kl�d���ˬz�7'G�m��hi^%]�y�='?����� %�a�E!�цe��\�:I������k�����rI2����8eS.3�
�;�w�S١m�w�Ɲ#�[���B���a�T��(�v��٘ÎW��K���3�M 2Q�r� ���F"��"ZZ�N��F���t���0}���46P��;�p�P���t!U[���<��|���Ȭm&��QI�57\��5���`C���}�B�ãj9�P�K�?�k=e"/�E�G�)V�d�ꑦ� �9����c���h~݌L�K�.�5 �A�Z<�:1��y
펴X�?x�N)/�8׉0<�>#����G��14/8��"��̓�E�����hj���ڻQFDr
R$f�hEůb�m��.��z}�i�^+/���Z�* ´N��\�80~챗`T�B�-".'I����H8�4�M:.��:�ikp�$�Mz%-���[Z<-i�]�{�H� vw�;��/1z�Cf+ɼ�e��I�h�����@$�!)���s{}��현��?���~���m�}j|b�I"C�|��i ZKyh.MM�G����^ ����P�'��߲�-+��׎�@oDPY�����G�<��/�Œ�֨'a�(w[f:��(w^;��T����[�=O<�DʛX�kn����D6ˢdF�o"��bS�`�� �2�6b_@�@��
�������i�޲��n�f�$"4(!T�?��)�d�4�ĳ� �*LV^��(#��\�H(<'
�s��U/`iݦ��I��3=?n��j��@��ݔ_0� �QI׷W�������Da�H��a	smCY��<���?tMg�]����)=8����3_Ez�8�NO��e���sp�5_
 !YY "�˴Y��2��)�?�\~S6�QD�F??cU
�*�k9m�;�~b�>�`f�<6�<1"I��`�	/k_#M�~W����7��U ���eIC������ό�v�+u�6e����zE*�5���)����s,s�ϩ�,��Fő�G��]xp�u��VQN֮���[sP��p2���J�Nt�nS����Ǐ����Q��qň��l�1�Ǥ�wH�]&asA�d�<\FPxM�k΢�C��>�PD*���`ղ�����[W�σ��/�p�4���G��o�]B���c���(Y�i�W-�Y�{_�ʚGԠ�`
b_V��9�6���al����{��� ���	\\ ��#�}��Lد��\�������o#�W��0~�T��Rd�J�E��:]��@���Sd�qf<	(;�f�7�4��`3L��������aD�,/��]^����= :E��z�d�́+�"BG�+d1�ԴN�v��!��y�s���a��x:���|�㮝��V��p.�k��9��lۗ��C��7���k�$��k<*���;��yr.����z����!��(�}Rfq�E���w��Rޟ���р�~y�����<���g��˭|c�̟�B�������X��ˣ�Ȁ�4<V�:ʇC!;�Y6`~���1�q���������Dc:u�?=>&}�э���*XZ-М{�Έ�q�����B�Աv�3�ZUY�OT��ptp���"��Ri
���1��.0,��F��O�h4�r6�-���L�m�k��MI[�A�"�`�q�p8��'^R5lJW��^�;��_��zJ�͎���!�.�T�)xB߳rwa�^��W«)-tn�<�g��h2< Z'&�&r�Y`�а�Bs��Ȗ�����N��©ҫo�d��~l �� ��^�M'��ޮ����kay�,�hP�ڕ��P�Bw)e�t~+�J��bsj{�T���*�@>2AC�N�F%�� >��J��m/��@�Tv6H�2��H?{��,�$T\^.���]]_�&0���G�<?��K�t��z��#��>�:�QTAC���![�x.l<p�bf�AB'6Ly>M�o����"Ād��8D Cd���kD�=�0����"	u�\^��)]_�|N����~E{�>B(!�<S�f��v�-���!�����Ic�KL�zi��;G���B�������V�7�Is��ɗw�>R}A�N�_|�k0G����	�h����xzDy~�����w����.�#��\=�y�_leEV�cB^Ԅ�P�t�O\(��_2�1%q����'�h����c�?W�~�Q�q!ꎆ�^(:o�y7��,�eŇ�^玷�|�� p���C
>46��>c�p��ْ_�/�i�qi��OB�!�z�#Y��n���:�/��>3��bN��2�{�z����ר�0� N�>f%�4N�{6����~;�VeK*�J�_���ڎ6
��Gޮs泚Rv��F�`;��b�പi���WW����'��^,�L��_��s�	pl�G.�����!�|�Y+�D�[��e�]ف���0pPnz_v45�Sŧ��C���qg敷��0�<�黋�e%�<I�X���bA��5���������@�Zc��F+�ᾼ�,-��5�s��)�at)����ް�ҍ̹*?�.h�[� AË����#m�獭�#���Lé��=�B&"Ta�I=�����S�x�փ���jL�p���>�Lv��9P8�{!���M曎Ɍ��ܼ�쩥Q��#9X`��=�/g~�gD����Q��Otw��>$�ػ�����`գ���L�N�\^&��.�״\\�?\�n#;�U�%��s ���J�R-���@h'�l��]��"H�:�`Uܪ ��l� ��~0zt��+��xO��l�Ay��T�fl1����$��<ֈ�L|`�պ�l���������L�9��!`�~3���F�/Ou�>��򦲋BIP��ן�e�(�`�1���1#��.g���'���\rZη���y��X����?c�:.Q���d�D�i�䢋��ȳ��T{h(2�� �Aõ�+(s��+�vU{l����8�A-�k�0��L+�hB6�U��<���H����3��pM�w����$�,�۷{���'z^=��c�~lMj8�^�<��%��ii��P���{�
���a���c䲟̍F�����&�@�Fdpo���&	{�b�`諛�a_�\��}C�����R_�a�����o��(\D�l7�l���\kX�+���.����k���N~���H���5�pV;����m(JE}o�we�J���5�<�5��J��(\eۆ_���K������6���N���
c��e�£EU��h����c��2LY��5x�h��T�2�����d�*���T����v���ZjD�
|�u�e:�J=n�BB36.#-�m�H9��/�����d�q��]�DY"M��EfX,���
�T*�V�� ������ r�E����m�_H_?Ɣ�P��_vBZ�[�ZS8�
�m|pd�(j���1��Ɏ;H˞/�n5�(d���>}LJ�G�V6�8�ִ֖�@8���m�)��A1{D��3B��a�����jM�è�aJ@Vj4u�� aā�a���FO�%@�R��i߳�h>��S��jK�����?�N���E*{2l��:2��b����r}���JW^Z���0��^}��~���EןS��zm|��SanxD�m�%`���Idߟ�'M�8o���?��u%���:��yx�a���2q���g��?З�_�z�h��?���D���t�U��1�X�K��7���������r 6�E�jE$�2}�,4��,4�	�sj�6ѯ�zE�Ϗ�Z�i�����dc�h�_w��Q���뤓qfJz4,
$>Ε'3~."s��Q9URV;@;@�ٰ���t?�Q
��+g���;@��D��3�*��ɰ������T�j�@^orqJ��lb@]
���(��X��-^Q�B��(@ O��*��0ȈGӜ*o���ގ�9���jSJ[�m`kU�W�E����DS���x�{Ep9����p����߳"5z]��egW�cpgW,û-�Oj�q.[L;.Y��)c�$���x�t{w�@�HU
\�{G�߾��j�յ�>h�-�
���YI����]D:��Е+�@�'S
��G�iXm�=UU�1rp@�:�|���$�9ͳ���Os��ǂ��յ`E��em�{_O}q���E?^��sKg(��woc�/ܳ�sl������p�qr���3���S_��}�'�$�������t��iە���ε{l�����3��$�ʓe
T��7܅��eN|
:PB�s���S��fg($�ԉx����V%��|�M�;��F��=n���t,�Ŷ��M,z�]�[�^X	���z@���z��b����
��i,�ke�k�i���m��m/0̡b���{��F9�4�C�Z�����{��T�9�a�|9m���������c�4�7-~�q�����j��\Fp{\O4!(�p�p�
�=�Y��{�w�dMn�z����;ت�'���6M�)�VӔ��G�ŝ �'��/��Ņ�%��KM�
�t.�ж��D(�Tzg'���-�m8�c��h{��p�J����D���d��7߰��x�}�*����F����P~xm�ҋ�
#߄3?����'�Y�������|*J�o88���Я!��/h�ۏ�f3�J�M�т�@ul�w�k�]�b�t����9;`]���SI�s�Y�Ї����}���&��mD����
Q0i��9��N"uإ�Q�t���G��8yH�
�j� ��$9�Zh��}vI�}"ڦϽ!L� ����,��y������1���#vҫU=�2Q%|�,E�ء�H*ye�Bmt���?�����"�N���$f��`"�����%#��������;�tu}�$�L႕\��ÝP�h�v��*\W~/�~k���S@��x3Ȭ-4��!FW�L��n��O�4I�n2_DC�Yj,����������WP^ی�+��� ��u����wca�t�[)nbX7�pTӄ�P�c��\������ac@��-='�F�k`��V��A@�=v�!:�.��N�<e���,��B���ID��0��.pI8vĒ*k�L��?��I�\1b�A�S��t}}ǿ!\�Ç;^ӓ���_���۽�hfD�"�Q$��R�r�\,��Fhyi:YZc��[C|�a=A	��v���{�l��Ɲܶ������j���o+�1:ھ�����1)M����q��b;(Ӱr���Jr�w���Q��pS�FiH���B;ۢ�`0n1��E�MwI�=��_��2d~M(i������Y���p��G�����?Z�Nȑ��o�"W�)��.D��)G��Q�����\��h�?������㎬�"����!�*N�s��`q9���Y5%�����&,� 3O
@,ٙ	������N��WOt���:��0�G.!J'{s��&IZ�����+��ReF*f�#���(�ŉ�Td�D���<Y��η"���������a���1S������Mj_��M��ᐂ�
ʊ��f|PI�v95� >6'c�w0őF���#V�`6�Է=9~)o��{#0�h����*?���H�񵑲}�o^z�Ҽ�?�\�d�t2���)�l�u�'��,����-JY�ݍ)���%��<zO��;ɸuX��k�4I�G)��\�^&3�häkOL*��(twyMW�ez���7w���h�n���b��`�חl��w\�O��"���s�p���V$�[2F�l�T��.k_�}�{v���3�s1H�n�eY�0��P4F���R��2�j�@�
x�z4E6���s͠�;t�N��j+{��uy��������9L�:*�5��Y�T��a��ek�O6�=aз�&�%<��08��(�؉N�L���n��66'͎��0.����Ύ
/lc���$���W��NӾN1s��y{��~V�����J�h�b��4}E`��ޢU�7�]/���noo�j��"���%6!�X�'rF��O5Ì.��CƼN(eβ��R�G�^��[51 ��8�ԫ/��D]��x�İI[���!؝�ou&,���������]��$^��E��C�h����Z�c¹�}�FǨ�RT´����O/��^����C��5a���9?#�������w����.�]���[�>�������d���lc����9>��h��o�f6b�-h�������P4M8,���PѦ2�خ-S�*/��U�K�ʢp����(��1��_�-��S��;�a�����)w#��C�U��cw�P<�βe���Ί{Ø��;��̄BKD�,Ÿ�F>m�9"k�����4��O�g�P���[��3>{5���?�CV#W��$�"
x��
��9�~��[�}X�bq��8��re����}�p���v�Q5�u��p�2hEg�V�yM�i%�S�o;>��ed�1���ɊExU%�p��X���0� �1�.�,�	&OHr�5G*=�V�Zs�9��M�T,�m�R}�:(�k�F(~�qV�i�>�}��*�A��а��Gr�G8�]|�����ލ'3��m�ΧWϚ�[��+?tXse(6�/����������Ц��W����T��#�R���k9[��f_߱�F2GD��0��"�7Id��� ��:"0P�B�,�q�yt�����ԧ	͗��������2�2�%	v/��N�w}� �B�JZj�\��jl�w���ȟ&8�V!q��'����k�P�H#D-y��oVVE�S�7��>���򒜽T�t�*PN��+I��^��7��"1 t�O�ڸv�%Ύ��A���iB� .���%ˎ�b�hys�
RQ��*%7V��+�Eb�l2��4�������K0dR[==�Pv�
f��G���Ƞ+����%$�W�?{ԿULξ����W�
G�a�Q#U8�n�����/�7�\]^2X�÷o��R��^������
#Zr��y���f�ϹjIыP!!�Rb��~�7�sԋ)y^)��=*t��.�A�e��\D�H��$c��s�u�4j{���=��?�o�a�6�\,/��_ت����H�`��~ˀ�LDD;Ȓ95��PY���W=�-6�ׄ��d�иc��K�Q��)WgN�0x�jzޚR����Oe�)S�T��0�f���1*���>?�ةt�":/��B{�	�l���}�+L�e��~��b�;d�'�G�������fԼ7�=��d1���q�mIׂa�a�V���񚏅�ƕ,���#bŻ�m^�~Dp�m*�9�\sa)�|R���
~X7H�Q<�մ��C���{ǧ$*VFVN�c������ݑ`6R�5�電e�g����lؙ��Ɯ����ҷ�?s�q%@�\|B�&�_PU��J�����v�/t������3.�k���p�b,j[7b��e7�ǝ�����J�9�n�I�ل1w.R_/��z�Uz�\��m��<)a�kz|z����&ӕT���8�l|�ֳ3"h�,3g��� ��#:�;��[���]Əz�Ӏ����/�~!���<	).����xp@)��
k^����+�\;��vH�}~/xc���� zO���bI��-�W}����ɳDw�Y�݃����㣤1%�[�i=[	Kz<�y���;m��S�� �2ѻ�I��l��鲠�(-�0�,-Q�]$7��jd��:�ă�3��3T�k �r�(O�W68!|�#x&/�#���D�!4����.�1tB6`�@��C�V���Ł}��x4Bo@��0;�n�	�*�R��� ��s��;)i� �J���.h�t'6�p�hZ;�z۷_���/f��a�P!Em�΁��<�p��,%�G�M�)��w4M�	����6^��h���A���C������]Q2�TN|ÞX��6�|��@�C��	9"&x���'��"g�A�K|.&l����s�9���g��˿~�J�O��T<I�j�&��k�=ߍ�������E���Z�D�z�A>7!�ʤ�V�T\8���3`&�Ji�
AXod�$������?��Ơu"6?����?��J��o�Oҿ+��?�ٰ�s�aFŤ���ܒ0}�����{"S����s�wy=��z-);ޠ���*���Ef�|��
��$ul_�;��;����K{G��f�zI�.m~΄bU%�ϵ����C�ϣ\�⛻~��������0|���<U
b�+����1�ލ�M��C�5r:V�j��=����*�n�	�Q�$��T`!�l`�Y����S��*4��O�)����Orc�z5�ֱ�Z X͙n����8)�Iz�$Z"&��=h������y��X6�H�n\�f�Q��^��X_)��z�^�{�$+���9�H6_mH2��Bb�@���%:�/gc�)Ն�n~�p�U
c�k�66m�Q��>^^.hyu�8�w�uyu�0�GD�@��������$Ⱦ��=F"t��C+��$���XЭAۋxq=W&$��V�-Z�P���9�˥?"�����N�^�t�b灋X�Z�3$�l�1D� m벿dVh��4KJ�󖞟ִ�Y�������M^��,sEOb��/6�q�WRzd�4�0��K6��l	�6bY�*���F�#HGe���S�h�*�ƻe��A�C����w���)/�����a����@j�]�O?��{�T�9��I{�/o�΅X�Z�׎�3����꺲=1�>.,��9�U���B�86V'�F`�L&\Ij1��t袙�Ǜ;�r�Q��'d�t���hO����<H��؊�ӨH�W��@����W�<?'z��j��0�u��Z("t���)s»�&���/��W�TV�6�7��	lpR�6���v6Q�s���h�0hc�g�%1���$�����jP��6L8F��M��C� �q��F:�����*�t&Bf��O&�E'�n� �Z�BE�#@��4`P�|v��k���@�Na!ę(K,�X{�]-��	�"T.X��F����l���֧	�՘]�oV�^K�E�D!7�4����5��/}A��݅�󻪚�s�J��w6b��'F��mu�e)#"p� ���//Ũ�S�W
���}��T�`\�)n8!� ��C �Z0����Y�;�Bc�֔��E��җR�|+�Q�(ʥ3{*�,ճ�c�Q6���G��.�wV�|E��FD�ʡv �^?pu����S�О�[ J��<\������q�҆� in.���eBc�\1�J��Ka���2�ŋt�D�y}��A��Gvj�;�~YUW�Y:�D�g�"傩��8�w��-z�SNnikL12"���C%Xh1y"�����Z�e�������{�����Fk[���(�O�s�㋏����Ǻ�<�2�ڮ������u�?Sc�G���~W�������^���F�a��I�ר�yI}��n�əVR�����܏�m�_�87�>�1G����1m��3�r�ŉ�C�渺c����ͮ�6��q�6��g�e��2@��@mH�y����<� ��H1>1�-�Â�#X�3Qu�9n�NH�	�T���H���v�ɝ�;��G��`2N�|fb'�fyn��Ҙ3�����Äϛ�
��S�h��9���9]]_����]s� 	��n�e@N�4��������3��V_y, �/�rV��Ά4:h��*Y;��ؒ�M�!
����Ш�e��p
���ު�!]0JeҰ�h�|>=�>-/.X���I�
����eR���@m�~z�)Z\Ɲ_�E]���=�+����	�19��q�y�ɶ��~�[,���K�Б�>]�
�Zޏ�ʜs;���l3WvE���q�/���X~�@�����d�s7�F�r��`z�ўs�(:��w��;W�=�G��o��k��������µ}[��e����`���A�������?r���_����9�HH'0\,��~9_R�h?�sFN�tt�H4��#W��4K�ͦRJ�J�#ڧ׊�3�t��-T_�(�f"�����[�A�7�N����^8�r;��Jנ�.�HM�,��`�Q��<��:u�� �n8*��BRH���̓:�;��Q�3���	�H}G���4��{:Gai��ƕ�|WJVK��F�`��$�iT4��<ٙ0��o�~�c8
�v���˫%�8�x�q9&PR�]`�'I���i<[ �� ��_sS�Ϋ�H�l��\E�S�V,N+����~ˇ7,� � 4J���(K����%���M�6�����̂�}�A/��d���C��}X2�G�;�^鿘`��0zE�e��Z�VJ�*_.�\��1 �p�Ξ��=<<2��q�4���>��Th1@���Ԅ����b����P���a�CI����r�ɼ4�� ��N�\��@u�+ޏ(�* ��̄G��#J����ω�X`�����(�ʠ�
�b}<��z�޸z���iƳg�"T�2�[��@Y���:��@6uޯ�'Ɲ�zvA;���k8�r�����p�3�����/!�.(��9�sˇ�}����|0�����~�޹��է�y�&��7}>�RcJf%��m��W�Ao��(��V�V���ׅ����Rk~(�d�N^��WaԱ�͈�I}���[m�M5�c:�(�Y���w,w�M4��ETmW���D���r��(�����Ј���[X���>��4/��ji|���a2��.C���bi�)�Ba��Ԫ���e�-h�&�.�vK��`�,�Td�k\S����;Wơ��,�hb�6���������Z~%��ӏ��ϽVS�<�CG�ײ����r�F���k���cG"x�d���i�^�MR ���*��vE5��x�#�"8fW���Wc�l��b��@�Q����o��`�`y��J�D)�`����Kku��*^����W���$�lA�ɂ�u����1��t��c�Lkz��S�H�#Ts^7,��O���)�ꔨ��g��B�v��o4�����N_�?{�%ɑ$���OZU �=������y�{�m��6HU�Ƞ�vMDU�̃de( =����'�FTEEE{qD�W���5l�z��z�O��c��Ο(0[/Q�/<
���:!:���c��5�s���o���'�%���zu�[*��֧�x��M����>�ɭ
��rK�By���*�{��� 1ʐ�$���F���<��~o��-3��������ӗ��q h󬒯	��%ʇ�6ry}%�~'���>><ѷ�sC���d�o�G�t�ip�uј�$:�{
-o}�P�x�ԯ4Ov`�ĎD��2�
x����[\^�K��w�i}I��f�����r)��� ����NsS���?��s�e�ԗUf�"���J4�V�h�N��Z��,ݸ5����z�J��%mu�x/?���,�Bؑ���u���B&�F.@w]̨�4n�od�Z��P��q�Lt��w��u�2��g�ז';_���}�����6��ݡ�����-"j���B1�cS5?����k$�̢�-��n�YY����ơ�����JN	/i:�:�T`��A�`6I��b���T�..���B���?�}����s�`PAGW�2'�L��`5}���C�Z��0q<f�3Ө[o���H8~�l4�,ʗ�>� �F������
����d&θ���[���O}���ҭp/`� �`����YFw{�B����_9E����jc�s�p��)zOцա����3��4�ϧ�N�-���
��K?pң�Jj�C�����/c`�U^I�����}�����o��{�����S�pI��}~h�����a�?�Q̶�Wr�)Ft>ƙg^G���|�wiN;�vk<�V#�be��r��.ڽT�)�^��@�Y8����[��P���k���7g���b��`Ѹ����7���^�k�<{�[���l����>��^fKģQo��P��A=���WS^A��*c'�x}V��y1�}Y�B�Oau�)��L'�b�xjf����z��I>��Q�ᎃ_�g��e-�T[�g��x��l1��+T����?X�&�y{w/��>����j���cS�&h�t��dly{˟�?�l�؊���|����ps;�Bψte/��<B�] ���v�����?���yT��u#��s�G��⢧}�
ա�nCf�����ܳ���l�7l�̨����Y,?�>�T�3�x�|Q�\KN���m!M�lT�����S9����Sl���ye�$`�Y�C}�浵,x�� EG���Yg��Oc�u���Z|3�����_;�/m�X�����]�ס�W�ϔ���� z,���x�h�Q#˧��?N�Ǐ?��ý��n-����v��9<Ӆ%�//	�߅l"T#�9��*��F�(X�w��$�r�"�,�ϴ�|z�����R��Y��;%� 5L��3�z�`���K�-��J}K�Oi� �s{�^>|��<>?����K���z�֔��������N.ҽa�}��̖�ˋ|J�ˏ?�H�z<�O[���e� �"#���M8rԿiB�+�i���s�ȕ�f]���ܚ�J���@����4���˖�TR
�:�X@���7	�����{yy�D�!��߯���+d����J>v)���B2��N^A%�W�e
`���T�!�z�!�eZ�v���e�^3O|�N�Ԑ�~�hh4?.G��a �-�u�_y!��*�a�b�7s�O/�C��~����Q�B+���Q��R�N������"��R����JO��c�|H��@�ƨ�N�+���M���ƭW�j2�*�kg�xj��3������!54԰�M)�E0�-Z��Ө�Fxt�L�r0�K�㿾OϰW4��->}}{�y�1�c}��(L���Jw16@�^�l�__ceQ{5$�/4m"�!�<�s�$DsXh�Y��UɬOh��$����~��3gǠ��)�Z�Y}5G�bu�?`{�1O��E�rKT��̾�����!���qC3��Mq�,���`vx��>�e�d�*�)e����l^O�߽?�%d�is������}�O~?����~�a�~�	I�_<8ơ��l��{�����=������5O��,����(܈��P�z��Q�WJ��.j��;�e(�[9��N�ׂ���J�h�u�wڹ���V�*�Ě=#x��|�� �dg-߀�`��0rl����{u{�7)�~;�gy0_�Cߪ+1�wZ�z����d�\ĸ��N����f�=���9�P BY�Q5#C���8ÔO�u�đ}>����v���@����b���@#��U��`���!��h6%�����4b�4{����k��Z�0��1_\��>�k��}�r��v�{���Ʈ��.2H���Y��v<��|�<e?��P��i{�ON�;F���G��+��ޖ�P�;��y���E�Ơ*��,zWgL�W��`����Z�vw,�cy �ĳ����4>�&ۗؽ1V��>�����oC�#����
����cƏ}PP�c���k�)�>�)s�&��颩Qx{G}�-}Bl(��t�N���כ��� ��y�M+�\q��vH_�2R����I_&?�����֮,���R>=~�03X���g��S��ty��\�WsqE�{�u�(cTD�h��S��忻|'�������C��VSxG��S��N����#��7���ne��a�BS'�/K��i�)�<A�[>1�m`�D�"N�uƎM���ڗ��'H�x@�C5�a��R� @�����r�;�d�����ϯ,+ ϏO�!�m�ر8&��VR�d�=�*��R��Ţ�~�}as�����l"�f���F�Zq���B.�>P�nD��vD#u*4�wb�/��cBWƈ�sp�`�P�<cק�x}?7X/�k��͖���c�3"���m�ݔ�4�P1�����`���x~�w�r��^��`��X��f�����=���k 8�Ǩs��ĉ�'��ʐ7<6��ez����d��V�6�s#���T�=�5��}��>��6+�N��^�^7o��d6V֫���/i�;�<X�@ͻ���E2*C�%B�6Ay= ���ѓ��8jJ�^�)�Ȝ���a���n��6�f���g +Z��>3��}��+Ŀ�He]'4Fk�`Mct�FN����Ț�
[x�[�;��J�V�1]�"�6����#�ult��/��C�����n�g�{~a�n�@g0(�f)*�gڋƨ�~�`}ؿ��HՇep}��(Y:����qkúj���+cg��/�u����S�"�|�s��k�����ql��l+}��)�����V����� rp�sk�0<{Jי�Kre��fE��.;݅]��O���:xҕ�˕�W��i�q��o[�/-�r#K���,��;ZoǲM��t��)��ln�!(��(���Z��8:,��X�m�d�1H��x�h0��Q��o���=��j��2�Ox=���<�d2K�&&]Cc�v%�Ƶp]5[dpa~ltcV�������f���C����^\W�ݧה\�x� y�\m[����Q�H8T����&pyy-�C�fL�W�Gm$�� w�.ȸ��W��<O�Ϯի��;�[�ln7���,�ʍ�{�8�C55y�|]xe�ScK�}����2 5��J�w���)V��G����w��"{�ѡa�����C��������~��yR��/�^�u�#��C�=�mW{fG��Rl<� ��{`Ш ��������ݕ|B0_�CӘ6*@�%��q��X��Y>?�A��]�58���p8�Z|��ﾓ�|Na{�8Ǣ������������s�_3�F%V,Hߚ����������,�3�!'�
���R^^�2M����B��c��Hv�n����oFnxVMU1]���kM�S3=�������=�OS]�2N�1���	U�Wd7�>�hH�V�qP�a�v�A'��ʩ�g��i\��lƎ�ؐ�z7�m[�<��9�j�Ra*H�N;��p2zv�6=�wr}s+/�5�3K����;=L��74���N��݌z+1&�T�~�P�
Y����Q���x]fZ9)���*!�9��n�saD� ���)���hDp�0��f]�����)���dl�)s��BH�G�<�X;���f���gH��q#M�a�b��F�isZs�A64d0 ���q)kT�JѰy�̑�2��~��,�Y(V9��5�b(Q�~K g�I�*s!=�6��.�>1��l���&��3��ݮc
UT'A������*E�mR� �?
4G�F�p�@��eB�
�@��tu( ���򑦆Ե�^�:�������q�d�dI�)���7�mv�r�ϟ�*+;����׀N6#8��8|e�5��O �5C���Sՙ���N��vs�޵���^8aȱ�r�3 D�!: �z:�x��P�#o1*�9���_#�9�>wUמ���곷?���ٽ��S���a=� �յ�)Y� �/�g~���#�g���Ur��μwd������6����g@#��y=�a@��#�7�"�::;	��!� �,c��  ����
�M� �3�]��}<T�N�j_����z��f�u��=4�Ƙ�S����PA�ps�7�Fe�Ԗ��kc�햝���[�6�;B����ļ�o|F�^��ڋܨF�`� �r}u-W�7�h��;xY��ԁM��l��X��<A����@��`�~�%2De�m���T�(�ǘmgs�!�@L��,���:��:�U()�;3�Ey M{���N+�t
���֖�N��5�p�%ك(E�yrFr	�x����V ����Wۤzα>�����~���V1?F��õt8��Z$�&�6�"��W9�ъZh�7�M�o΢��~�����'�ڒ�v��m�b�f��(Vu��򝾄�K|��G'ze���l胝�����J�S��PeK}5o�}����s�JI�Fp�6����q�9n��d�  �Ud�`^�ƙ���'-��|p�����$�K���fϏ�N>�2��O/�4��R�`X���d2����H]..d>���d!�4/��𸹗�tb�A=5����NG�^\�ZdHqf
vO�*]a�����}�$�6ͮ��߬ewy��w!q:�k�A�����)��� �r+�~��Fu
P�+��K��^/vQbq�9d��� L�kL��'�|GP��ƞ���٢
V����Dno>P�p~���߫.Ϗ?����;j�`��EƳ@c	�;�q����>�w5N�=脶@ ��}����zvZ���B�d:"�%�e6�J�8�ҵ�7��i��.O�(��4�<���l��rm�w1&�9ZC+�J?�ϳS7����k7�54�.��4z��Wm�Z2(y��!,�2��izF-�ٻO��Ӄl7Z2�������t>�	4�rE /���Y"z:!=,�������A�	�XBEtg�	�,�Y�L��Q�E��h\S�o	��_q��}���u�y�����K9��J��Hf�	i ���p�	bD����%Yj52zFJ�����dL�..�=A՛h6�����He�%7,k#��y�0Y����~s���X�K�;{����������Zy��q $ԧ�]�_k@�9�A0u�P�9��Ȉ쨔V��W�+�H>��U�[���P���1X����'2�:0G�F�uǒ�P���������!7�R�!�f0��)�� �̵���RP�!(s��Z��, U�x�t�϶���S��S��̖�V��s�u{ �O�������X�^˲"�
��sZ���2z�2��,.�g��wӪ�2v��ǚ�C�L�
���S��^1؝J����֖f���y�<�*	ʬ�,��k�uo���Ê���Bi������۫Z����Ҝ!�n �`8Њ�/.�s���|� t  �cZǑ^�^oY"_K�B ��3@V��TI���2��(����\Ϣ��	�wÞ����gn?3����e����i��ɗ�4�`���:���"�k��$�3���!�|?}�M�s���gy��T4C<9��+L	Hq��:j�܆�_4F2�B�����/-f�6�=���_Ot,��1Y��W��X����Y�:u�{����ϕ�r�U�;���lEg����_�qb��d%�DJ?{ӱ
�Ͼ��W=����vAET�H1�vpi�
��\6:'��&�l�4/��7��S i<�ps22��G���|���[��ʜT�/��d,W��Okڦ���f)�gh�m2���o�7�D|�A�K>�M��"�ST.�Gyz���!ց����Q�0ɷ�k�3iGd� ��Pg�Ļ��6�e�����QV�e�a-��^F���<�,Ir�.K��'e6J0��g=2q����:t���W/>��At=h��eң֛ɉާ�[�l�K�1���-�PO�������{�(�>�%G���G]XJ;]�t��f�쨽��X��x������֔��)ٹ`�\KG|�X��Ս����:ڧ�?K�Y��=SP��L>���(j����s��s�!v6{��Ӈl������H{�\jg��#�X�e���k�@�c���h`Ǯ'�4t6K��|�ҵ\�\q���l@W~&�t�~�@�f����7(h?���@X�$݋�}�8�
�S`�Z&�L�1��L�FftO����3�F���;ՏB[���b�4Y�Zd�g�]gy�b��?ːZ��`k����Y���BU�@�d܌��5ʢ\�B���&?��`,�_��2[����	P��^ШzIcGK�*������GJq��N���q��"V"�Une��靹�
���3�Ϝ��
��@̻��b���'�m4*y�u�Χxm������1�s[[���� .�2�a{�Uא�����Ha}-R,{Ƕ`n��HQ%��}���Up��i�b|l��o��ݼ����_=�i8q^��x�j@�6b�{�Cџ�>Sw|u�2ǗJ���8[>X5�Ji0���Q&�3&tl�N��nmv�Ji��=���?�����ֶ
"����3Mnؗm��W���F�/�<�^7�p�Ds�̹hXK�c)�Mx�/)����ȴm�4����+��W>����zD�����WJ�j�g�� ?��V2<jB��X[hE
�WT�N`�5RW]:n����)2�u�T�~���X�˹}Č]�t�̀�XxA��(X�y�l :��%�mD��]��⧟��Wk��v�QT�[0E�3�YX;��b���`�9P�;�&�"���!^ekz���(}K����M'4<2�).�^ZFSc���˺��6Y��a�g���,^�K2�_,%��)�X��9(����k]����N�2��/^��`f}��C�QҔK?k��<����8�cH۩�L�Sln������n�x��B3��<p�q[��r�`�"[��8^���W���7�c�]zc�ev����l�71ےy��e.�L_��%ڱ�M��W�7l���>�E�?se��}������;�}����۩�S���g[2hF��ei̽I��d���L)�Ό��Wiq�)o�g�Ё�9"H�R|�Rm�E?$.��8��-+A��4!�����4��AS1w��s�(�>�8��+͘����:zc�qN�H&#˕��A��2y�65�j���Q����\%?�:����%�)�7�)��a�$�x�)�J��C��5i$�l�Vn���l�">@����R5���E��t&>���q�'c��YK)���{�{`�<��;�\�Ũݰ��Yr.̽ҡDF�6^�+�;�QQd|w2��)�ͷ�������k3��z�H�:l"�t&sD9FyFO�S#Ek�;Jo��-b�0����� �!����T%�,��T���r<��A[���KE'B��'4��Q0:�Z��:����;2v�ء#C�)X u6,�-F�]��2u��+�L�S-=h�i���g�2���R��`��lo��1�w�W��X� ��bF�i��o>�!�2��g�0����&<�B��Dt���f��LjX��8atjB���r���;S2��`khL�vx:~w���/�B]�=sJ��@�G�
���P
}�ڦ���q�&���Xe�&O��|Z�
Ñ��|�A�������\ž�ab�R��
p����'6�L|�*�d�2C��L�Z�*�5ud�f��-�� E�����W����;��6\�zAKt�iǥO�0jdDy��DFR;`�A��t6'X@G�źo�g�y��f<�xt��h>#H�b�Q��J��s`�E�c����>ɡ�b��|�������5U-�s輦�UfA5�9=��O�W�@NKQ�F3���2�Z\�5bTVӑ������H�	kԝ�V�.�;��p�U=�s}T�m�[y17�߶�$s���q��ma0�u��������jjd�v��ȋ�8�gS�]K @�^0`�l�--5� �;u:��b�@�/�A��q�B��W�ҁ.`��;2��HM9����H?B�loU���z����ˊb�=S����Ʃ�Wu0�w^�>�3��֦n�����Mw�{����`]Wf�4��r�jn��Y�v	��u�>�l���a��!��Z���ʠo֛d���]4�=8oY�H�;݇�w�⟘�[�+@�H�V�o�נּ������!ol`�6T�(�C1uP��bOe�������&�&�~��՞�7��B���'��LA[Ŕ����5�e�� $z�q���˾bH����̡�����	Y7
��6#z��Ԑ����^��]4���)��� Tp�B8���RMx#O}�����r�];��l@κL�پ�R>��,1�����z���&V�0�1�)[�u���M�~�*��/y���٪	�؎
�xC�l�Hi��i��1U;
侲e��0@Č'Z�<�F�qQ: L[�<Hq� ��bzc�2+#ͻ���;X�c�sd�����Bi�6��Y�(�O؄��r@[�+�4�\��]����:,��@y�-ʷ�p���D`'j�TA(!��o����N���{VH�=@�f�|��E�U��-����ۙ],r�[�'��j�����5��,��y��D�`4�G�)H�o�R���6Z�br�͒����t�Ւ@����O�i!M��v�~ÈA��.���|L3��k_ ����,V�H�w�3�Aڐ:�P���ɘ��%��#@���al��Z�B#gJ}���	(�,�sٯۼ�!�=Ġ�t���x~u��l[�wNN'�j��hr�p*�_&�JA�*x�H�{���K��� � �F���Љ2nhD�(6��g��F~�����(Q�b�0��cm�Q�T���"f�0`g2�Q��(��GBH���#)lWUYWu#��AT�QP7|ܙ�:s�L������DӱƓ�'
\����m�c�R�j�U�h���z����YL�=�B8�/I���7��ɤ��se�w������gݬZW�/Te���ڟ:�k�瘬�ɩntt~r�];+3��B.��83/�	���ļ��k,ze||ni���ѐ=���d���Ͼ7�o�C1� N���"��&����qb�WU�����u��i�K������p'NB�w�?;~��g�be@Q����Cf^����r0A����wQ��:��s�K�f��!�p��g�W�o<$2d���;�,`/uB��}O#n�:v�ԩ�pG _���b���h��T�w�њf�g �;��0c,b�5���C�"�-��N�9V���R]�h�5��O	���=����G�w|ރ�����p{�xZ;o�,+����1}uyM�,��z���;���e2�aú�s��cT����K;�����j�����t�(��rx�р^]��!X�g%�-fz���?��LyWQR����G�Є�����>�&��h n<1���>��z�ض�ə6�D���M" `��x��/�m7a[�Fƞڒ�t�k���DO9��(y��j�[(q����Nn��g�NIa.	n�Gg��4�n5��[��\ A�9d ��X�ǥnU�|6�`Yc�d/����
Z��UŊ�_�꽪;&�xM��r[��I��aW�נ2�9��W�R'��u�1� 8`��k������Om�4��������r�kڄ������([M�+�,���#���Z���P�S�&� ��"����d?<=������x���lW���)��Z�$�k+�q�R\b��z�B���4��� 	�S�;Oc�qȄ �=�� Ƒ�i�$�t�|�ť��=�F���fs��ع��,!�������ݝ<�d;t��uA�m�c �6u����
�9P�,���pw}5��\h��v��4r$V|��.e�~�sH6Cr�A���Z�25���E�w���<��z���<���|o�(� ����i[{��1Ұ'mt4��ᤅ|��EZ�780�B�w��泴ȢzdyG��}�gtԤ> �>h����J%����¬@�}UD�-�S_<+������G��=A ���dp�����P}\��;8�.� _A��r��oU`�j�#�A�m<'����|�5J�o��$O4\��G�A[�Ϧd[� �P0�)]:&�NA�����v�A���:S�c��SiG4RX��u|N7�����k5.��M��=�`B��F���㋦+�s�_!��F��m1�/r5/..)���U���iU9�����(���������1���,��h1ej���1P���{#ڝ2 �0��mw��A�7��9�\�ѫ^d���s{9ԯ�}v8�n��[k-m[��P�o�N�%-W7�r�^Wi�GU ���D,������P�`"G�;�Թ0�|� \����[��C��?��$��}4�����s�sh��cWG��w'�×7����x���I=g�x�	y����_�ec��-�[v6ҒZ�uLo;u�o���e�ޔ��)5���V}����.�b�lc�Y����X�4� �Vr�s��`댘:�y�i7����!D�"��-UI�RO��S��o+�]r��f��F���u7_�%�f"nz���z`)X���A
�:��n���c�e����O�~��q]`�#X�[]͓M��3c�k��oh�3�}�D�i��ڐ8	�9�^\N�9. �!��C@'��x1���JoZ�uP��sY��5�ARK�W&��F�$35{悎 ����>c��hiӘ�"�(��i��#�I�*kɮ�P;�E;�,<��Ů
fԕ�|8� 1��it��f��	vKeD������8�:.�y���q-s�0���>R��4���$BS���1�����K�y��Gk��p˸��ﴔs:���|_�����K2���$�6R����
Tddq`���y���8l�?��D}6eLx5�s[�>��[��d, 
!�٩�:$9��Y<L��µ~"} k[�30�Fc]?{��)�y���A~��'���#�Q�{�WdQ������E��c��d��i^�����"@O�F0_4�ce�Y-X�X3�8׍��fi[�֙��r5����ǸL~�e�_o��\%��J.d)XGS�y|~�Ow��/|�|�'V�z�\�L�+ڇE��H���c`��BW%~K��:��`H9Px�#թ	�w���u�+:4V���qK����Rܾ{O��25�����j��bM$ȿO���$��*5w9�!���X�~�"�Ur�H���b,�~�I�{ߒͱߧ�hz�7�,�L�ުSt�~(L�⵶�	X���m���rԥ�vK5PÎo/�t��!u~�h,�Dj�=g뀭��f�f�7�ǁ��XL��z���9�O��#�e���ӎ����5�4�v���=X[`zu9ʆ�Ftn^�13`�Bɴ�A��F��}�ވ�ÍF#V�[0d���2��'���^�jF�8�F��OФ�3�`���!������~���7S��}�ф`�]�<�U�_�r�5�D� ��`9M���Έ��5��^b:	����`�ZH��.}�k '�>�1��u����-l�nU�����׺\oU�T@Z��
�����AG���5cZ ۼ�G6�s_�:[x����GN��#�g�vuJ8���E8���x��G_C� P%�=W/�~�T�������;��?�Z���h��|��s[({n�=sǜ0��[Ѱ�2>��lh^��K��"S���y�>h���H.����g�ē�W�;���rLؾ���g�n|��y���K������#F�Q�ྜྷi�tV%��YYkT	���h�F��|땚��O��{6�sM�Մ�T::����CM;��5��iO%1ք:�j�+3�Sd�^��e7tL�7M�X�P]~��؟��mLg�<U�i��v�i��! @����[��2�j�)F��yJ=,�!H����:9׷W��zs�U��� �,+6�ɰ��h�  BZ:�nn��km�#ôϖ,~�����H�XЮ@z7��>�r�89C`��|B 	6Æ��aL���:(1�W�m�r�nL�+[o-��4�p��Rp�Vs��G+�� 8΅���Ǘt�����y ��,�Y����dߠ��8�3XX����?��u��h0j��M�a�ݪ\��������ms��Y��w�L��b9��o���\������ �@���z�:d������*؆�-����*���������@���Wb�Ǧ�WS�?�������˞�3�/�� ��	S�m��Q��S���\�Y���=�E9��@eߘ!6v\&;��;y?s�O $cUܥ�BT�kJ�#������o�S�O��d6�&��M�e�BD}��?�_�BA�k���yl�6�������q�Nd1����RP��&}/|�rsy�,��U�Bژ��|��v����C?.����A�𺗗�Z�ض9�]a��>�#`'V�N���ߛs����A�uRR����8���lv�S��1�6���**�v}y#n?��y�:P�����a3�������TViE������tiۮd�~��*9�Js����p7fO�o��Ӓ�/6 �c�M���}�P�-JЖ��^�
 o�%i�H�r����at�_�i;5�3��Y�{�L���p�m�+R�@]Ctd���,.g�`����j1���Y�}'3���� Y�Xb�,Sw�(���{h�Ъ����FKk�i!�b1����jz���<�ԸA����_^��*�_��yo�ySCD�ˍ,w_�B3����w�o���o6Q�l����fc2���V�l�W��?�?��!��7RQ�m2Y�YPQXgT�ý���F�}^@���W���fu��}�w�lt�%��^] ,k��Z��&xi�>���G概I�4q�԰��qDs��L�n���2���{�H�h}���`����sVCӈ-ƅ�=NҸђ�vr�td��ʶ�꼯7N��E�q��� Q�.%��:�����*�.ֻ��N,��;~��xE[f`�3"
�4d;Ę!I��\c�_� 17��ܹ��x����}�:j�`���k�#P�3[��S���s>��TP�����|�i����g��c��Tw�� �;�:Xb.,6Gs��EC{�)�w�KƲ)P��zV�2�b�{�ʉ�+!)L�r��=� � ep�	
�Y��?���CZ�����66h�L��,�[1�Ooh��M��,V�<��[$=�x�iN��us�b���������2�� ���ˇo�S�@��V�r�\@+��+�����E�^���0���c�ce7C����2���h���R _���$�I2�^]NN��6劎�
�`evh�HOn��������[yw{C;f>�á�M���Z��
A�,ݧ	K�#��ղ�c���j/2�נZG]@��;2�e ����Ԫ2�O�'���ƨ����4��=3�z8p
�fX}��4lJ��]I�:`;(��1n���G������:��b�����w�#� 7#���1��B�@�R����/ع�[�*v��;��i��oIn9��5W���nd���)p�Ė�lwo�N�6`�ur>�^�這_pu� �v=�V0��2j�,�ML�G6P�5����4/��f����}�h��"�7��ͻwL[��������A�~�m��1�ԙI��f�@=�X�;8� &Wc�P�����̯rq{�Z���m���N��ŵ;�+��.rjkΈ�c������?��ӏ�3XF`
��^-� {�-3�$0-n���~�z*��H��\~��܂x�6�eQw|���+!����qq����,��˂J�"!i�$u�������!�N5�=�[�"J۪�g�˟��/(�{1���LƳ	���=��c��˴�B�h.R�j5����ܛq$ybt�GoH�WoPvS��J,����i=��jF�0��ic�!��M�j`�FT=*���U� ������4�&Q/��#J[VeP��;��3)�u2��_�� �����6?/��2�����n�4�w���vc��a���� �lq�S���gӑ��߈:==.�u�ta�wm *�̌"�4}���9�&�Y�r������q������k���1��� mu��L$��LD���#K�__o��$�y��bV�85�h���G)n�8m�0u�������d����9X����xb,�f�9��ܰw�����tJ�1oJ/�fV�w�\��;��_8�=}����>gQ�m�GQ������qp
> 21K���o�I}s�*X`�al P_#ڰ~I}j�Zc���ĽS,m��\}���.i���l�H()E��t���ų�S�ow���8s�I�ZI5�R�K=�]e��M�/|R=�̸�����-J������ۤ!�6����v۹����+_t*\����-&Fv�dl�E�C�m��U8p�8H�Š�u`�rfŽtc9ۯo�vM�{S�aw��ƥ�PK
�k�J��}��Pk�L넲���93
��j��jv���e[�d^����<��)��d���R[�O,e���1&�G���Y\�&E@g����\e��1#�HP�\Y,�Q����Ʈq�j�s�w���XB#�e�F�}�j7i`i�*�����+(^��͙�2�2�2��\�^�mͿ��Ύے/ f�`!��@���	��o5@�6"�y\����	�������,���<�lEJ�WV1_O-`�ߺ�BӚ���q����U���\���05�NGV�(�PS�����{�Jk�w�~�B3� X8�R��{c���l̖�`^v��%�E]%aàr�ڶX �١�~�k�������%���;���ܦ�!��K������6���l����n̿u��,/c�lC����G�!i.�J��*S�_t�q�d�^������	Ԥs�&3�����5]'[sR�P����Q��VK�#����%�s��6��ʹL}t�X5ɇ��_���i�cǋ�}`5_�?�6��'�_V/$-`��SX92D��z: s��ܦ5�Çz/�!���p��!8��BpY���&�,��Ʀ�h����O/�Kg���=�@Ӟ@O�3���@�Yzq[�"�B��ň�+�O���*VV^�@&j��ub=�hхԯ�;W�U�@B�CD%&��񒢼W�Wrus-߬���i�_���&u��i�jR�D&��k����sD��ԕdL1�Zr�~w�yDm���?j��hQ斥�[���A����hr-o�gkQ���`O�KY�l�3F������;S>��l�����VD�;Wg�vdk��Y t[�X2�]��;V� {h��B�V�3 ��2O�	�?�A'�	��m�N]J��bB�m��&D���ya���T@�%�߽<<���Ӄ9;�f]kTn2%�q��{u��~2U�*N $�j@����� @m���6!�Nr�P�i�(���Q�����%�u_
S'��Y)v�i�˫J��S=J�s#��^�Q�G9��	s�(�Y]o0
���"������'�S��Dyۺzfs;�v|�R�<ܧ��:���b.�T�ohl�6kwV�����C��1Q�^��W\]�;uz����;�#sg���o�a^o\�b%N�_���._�1� ��F�X���\����Oa�����lȅ;�-��>���b��t�A	�M��9��V��.�*n5�#��E�b?L� ج�O@$,g5���.j��v�ݱ�����1��\p� T���j�Ko�KY*4��t|帕W��_��j��S��O�m38{5GL�����ulL�Rv`'{��I5����v(��[e� ���x?�6��m�)�x�T/�,���dÌ�6Q|�>�@�dPG+y�cb��Za`Q){�t�d��>�V�06S��#�|���n��z��O��ӫ�d������U�bDD8
NjX�Pb6�
�h,2�B{�z`��=�iL�w�0|~����x�c��1�y��ujc��6��SVVH[�2��;�nD`�E���Gҵ�d:�}Ús8�8v��:�����U�F��u��>�h�d��,���'߱���Yn��:�m��/�r��,e�*�e�#��7���}6�����{��@�_�_�R]!L0u�͏�X���u0��A�4wBn�i@{
�=����05�*h �d:�\w{[G��ڛ����zv1'@�����0�s�����T�qL~�S��:#��4�����g��i�m�3�����J�T�s�;���Wv����];�fc���������5�p��傂���-S:��g�x�k��]4���X�ۨ5� ˄y,1`�)D�y��[�IU�,M{j�+���v�����r��Z3F�������;��f<"	ﮮ��Fw;O�;�@6e*{�ˑsD*���
�E�0�(C����RF�SҲ:,� &�.ܘ�����R�ש�^��S��y�n(h%���:�h�h[Q˶�b��h�X���2����Q����2����z5�q(ʀ�5].Oh3�
��l�����kJ_(.ڑg�j]�	�Lf
M�����B���j��9�Lƽ�&��\��t�5ʕ
#�Z�U
� �Y�8%+z4d����aF�*D��ߧ��5Є��c���LwL�b>�kg�Y4�B�'�1�p�(���h��
RM�5��ز�V:�V˧�<�/���� ����<��je9���c�;�^��B?�L����9�Ĉ �'C�v�RSw�k%eUI_\�dt�&���[��ȦCY�0he1u�j��@�� D��A�o���ў��i��xDHh���i�{ע��RE�KOfl�̔:���g�̃&:!�M��ۜ�P��)+�#	�c
,E�.�"  R��-�U�J�AaF	H���
#ү%�,0��("�o��"����v�%U#�l�\bb�xXgI�/�7� 菀�S�=�z>�_��2��-�_X>o�w�	Wo!����z��o�)r��X}�mh�]���z�=� 7+~������T�~�sWP��9?����W��W/��K2�7�[������e{2���4V�ҽ�"�)�o2�c2������Aȓ�Nv��,|�gV����W_f)���Fbv�ū��}D]����R:M���8�t�'T	5��\}������O����7�C�9���_�f;Ҁ�O�h�����o`���?l�z_���j �mX��ַ�Km֏2` 
>�Y��un� ���z%jo@Kgn��#��-��c2�<����<}���k�~�:0���leh�'Z����+yws#�L�<��[���b���GBe����"��-�} ��}w��!H������L6����jI�XZ���ͫ��K��LV ��C��̚7�*�ta{Mr1d ��$�od�<ygZ2���M�c��VԊl��4��e�5���$�/�%,�;Ӌ�zM�)Z%�}tO�������{�f�a;~~;<F��
5�8�C���^�:�	r�gО����y�'`Q�K�U�'-�A��j��9G�����y�V�e����T��.bm�ze����e����z�vQ����kϗ��_�.;��T]?屳��򾚑�iD���#�qk� 9�'�W�0�4|��I�b��_�T}t���f�_赁��`d)�(zԌU�Z��G��2�\��v-�l�^��ϲ���ZUJ{�Ƥ���� ,؟������\�����~���`b�H�`����c�]��i-w��t��Y���W�U�����,H$7n����z(�t-`�>���w����@�����l��+U� ���1d\��6H�ء �vc��t��~#��>9�ir��m2L�*�j��M����r�h�3E�� D�j�x�BT�թ��K't���+�S�{�J���.�d�0 ����if�u=���*�?O���t�N� zr�;�����殫b�}��8��hfX ��S��Ns��ћ6��X𑗽�æ��������\�l베�>oO�"r��G��u�{d��΄��W��V2,�	�	�ܞW�p��fi�n�}�)Fbj��r'�h�B�.{@ۈW!�A Z5F5t�ҺM�5��v�9����ӝ��?c{�.�0.�&[,.Sے��������"bۑ�\�h���0���5e��F/�s�*����E�?=ke�t��˥�}�����]����^`�)X2�8�>�x�(^0���Ѱ�����43�؏�޴UL8���)���U	
;��AC��=��|�`^������iGnHsh
��M��i��q�RKI9
V��tMl�73�|LQy�A���N�Q������߲�������w<z�һ��4��܊�(R��m��)�v�� ��zm��_����{0��ޞߣ�W�y������kIf�Ӓ���܇�mn�rL��N4}e.Ԡ�9!X�;�S�����t#9�iZ�Onf������[ȝ��˥��0�Y=~��,������;o:����"�j����l��:z�3�[�y�T�<��}�[���l��A$=�����i��u�?kN�n��j3[ :x����\7G4pU�M��,ME@t>�V�q�hT^)Sq��;լ'S#Ci�r�v-���23�_<����1��G���X/�F
�`Kf��ʭ�`�$T!�R�h�\^�9��
��렻�AP������@喥�DP��?N$�0�{�Y�xR!�5 �g%�ٜ�_'$j�6�� !أug:{�(�LN�H���P�'T�o�l�t�V���M�gb�` �B�j��~t��vh��V����#��$���v���v�m�3�l��;z�S` /Z ��[���xՕ�Z�`5ޱ�-��1v�X�N��N�y�n��m��Q����b�ڪS���y;b?����YL��iG���c���s��2��_�x)�Gc�-[�^�_B�陒�R/�O33����B0̙�py��:خ�
�O;�"^D��_{e\k|u�s�À\<�X��&9:��(��	g�:�䴭)��<�-��_ �]�Y<��������խù��a��#}��F%<|���r:0R���/��`T�z�v�u*���@�l�%�y<0#_Vd��y�4�.�:��9S�������E�`�l����Go&i�[P� �ˢ8��6|���}�|yc�Ը�t�|�Sg#��ϛ��������������4�dE�N�`j	��\_\p�������w����I�R;�ɦ�d;���3�9�����H��{E�/v:azޘ���ғ���*@ԥ��)}�����<�|��_e��s���"��9�{�ʣ�&�O?�ǟ~��z�GiI �4\0%fc�.��zj �H�{ �3��"o!�$����,�ϲZ�XZ�ǿ� ��\���Mr����Y�\��������c�K5sqa���3j[)Q�@��*c)8�n7�⥝E"��V1xj
?�e8Ǭ�0��lA�tZt���{�K�&#]�m�j~�hJ�h��)����B0�ᗲN��$��k��ǟyF,�͖��.8�t�%咓���"i֝��\�>�1�L`z�T��\�T����Q�,y�갼���R���5jhh4mմ�}��="]ٖ��~I������#��y��BW�gu��wl�5�Tc�Sq =��Q��OZ�xo�©h�3c2x����t���&G�Z�t9 �'0wĥL����3zMG( k��~�i�;�j�#
�1��QR��ZZ���f�m�n��*�����O���_XK�� +�^J@>�����R���Vi�I��"�Su3�>py�����R�ČԨ ��j�:�r����<�ny�!�`�ᔝ,7���4�,_ܳ3ب��3W�1����#���hX��?ST>�r�d�V�
�=�����'�B�?޸��������:;u � ��V3��w8�:�oU_?bO�nf�U��j5����Gs���ׯlmwv���1��k.�ן|��5����)��fLAB@�1�:��*��_8 X&K�l��J�Ϣb��R�1�\_߲�l$J�� �l�?���h �9��^'���vl�����
Ʀ�����W��5�A<h �f�GN�*�W;��D��a�d��������;أ�}Lǃ�7(ӵ�����'�:�'�?��X����?�L��lu�^��<� ������H�(s����,ߔ�ܕ �~���G��}-���]B^_|�����p5�U}b�h���K��u�*r=���]���3�ڇ�Q.";�L(����J|�7jL�`�AIW�0=Q�]��q6g�9�o_��v�پ���2ܷ�T������Z�!`T�j6[|��ͻ]$n�[  ��IDAT�_��~/�6T����AR�@���>םIK�gh4��	��s �,ӜJ]�톌�����k����c��\��>I��(s��m�1�g�م��
�4����?���2�q(b�#C���N�U�� ������l
-����?��;�Q�jK`g����R��������"؏:���!h�����K����?����r�FE�1_A����[_���~b��{�ɋ�=a,�*f�K�6��h��S�
M�X��>�i3ģW��,W[�l_be�)^���/��U��_�]non���F��S��C:��pSc=?<je��GN��a����Ki1�^OW�}eˎ�`W˯N�s�.l��L�Xܖk���t vP�hJ�`���  �8]J?b��}��>˓�c�4�XX.^,{=�!���D���М���� }�!�����vTL�@�A{I��>u��OwZ�4K.�&h%*��,�Em�|��W\�c�`*�F��U�)j��b���
0�had	탖K7`���!��:<#���/k]ȗ�=5�Y��q�L&9�y�V�ˢ)� 1J?ޒ�`+�niz���'�@�*л�� �ӊa@n�z�����<�\*322��-';�QT���y�5��[X3���#K�/Tc��j��D�$c��VM��:zB.]ܤ�w�����<h��}kQ�M6�p�=�8c��Α���3Dۯ�U0t�<W=X?Rv�+�#R��p��)������d�=�uD��$C��6v�!*��Ů7`~p�h�C�K���ӟ��v�i��&Q�k��}9V��>
�H.��A����ܼ�h#.h�)�������+c�7HfQ��?�?��v�J����6���eԶ�|���vp�s��	���[.�:u$c5ٞ�xV8���ED��T�E���K������_0�������ht��Oe�N�x�|�+b��@�]	�*����؟:=<<��~`��3m��w����f�Y��|�;��*�^4���e�� �î�1q�; �T["2%{�n��=Y�|�.��nMX�BK�7V-�)�6����� �i@������Ɂ�����;ZA�f����=;N���rE'6.�*%f'N"���KN?�C���e{y�����cTr��s�Dr�h귦a�����@]�SF�	M7uj=��f��X��ƕْ�y��&�Ϡf0ygl����U��[E<�B�O9�i���������U�vȶ[����ڼ`���LhW.. �����Ec=��:9ev
R)�z�-�����]��S�W�OلzZ��K�ʆn4�tZ^��c��+7��.̦�hcSzg��C�b����ys+R�V�O����~�Q~��'�������Ԛ$�ӴV���@ [��]Z������s�t�Q~��(?}�Hƌ��ݩ��f���݋��xZ1k�Ώ�S�x0Y3h��߳h0������Z�
�?��t�[�P��������Y[�E��j��������Ս�O{���O���A����㧟d���� e/%��kI����s���N�'��K�~Q٧*7��\ǂ�H��R�/�ɻ�;Y��C��uZ>a1M�y�p]�p](Y����-����N֝�-c���:�ц�(�`B(Ld��t���UK��	����N�����+���fi�tO�cg*�ϝ</�C�m����=���R�7.F�5&*ʾ����}�[ny���q�y��a�өu�:l�J,+G��e 0ھ�Nby�t��� X�L�u{�j�M��0X7���	6��WS��(��i�Me����dZ�S}�7`�����b�f�ܓ���d��̛]���"
�Q+�E���:VP!Fk��Q�&�z���R���5/>�dp�\K.�i�3 ���!0�/F�z��6t�ҿz�y���U���a�9���[:�^߷fh G_��J�/�� �vUܶ_v c�2
�d��5h�v-�h��ĪʪFK�#�]��T��9���XU�
?��ҹ�!T��=���k�$�-@%ET���w
��gU��~n������^B9��{J�Z��_� u�&�ύ[�|el�L3�Z�;?�3[���Vl�mAr$8W��-
�Mq$WԊ�h堧��J^\�Dl�}����R�ެ*������Ϟ/�R">�he� �lk-ҋ�-lM���!�1�p�ӆ@D���ʩv$�7���>>��*��prVk��Z��;7&�2��I*]d��<R���[�}7���F�- � 8����as	��a�+�g�&���NB��)죐�Os�&M̆�C������H���k=�ѵ�B�����s��o���%/{�'�C�$37ʃ��L6�UM��s���C�s� A��8��v�iܗ?Z6㷬��-��LSl�RI�0��o4]?xt"��e����^��Q�\��sz؅���aƈs���a�rX�,eד9f:HY�UB5��9��o�����pvʂ8���6�Zt����� ���O�����)���c����D�}G��Ͼ_3�0xN�x�#h�9�L}��; B�Z �K?�ϒ�[�X�ECҹ�D �A���F�Q�&��wkV�ڮvu�ݣ��7�ŝ�vp;�d��,�����9����>s���T�}���gzA.���׵Z��s�	����4��^6��ӝ|�#	����-��)�͒�̏��Ԧ��{���i��\$�X߈>w����Q=��+Gڳ�P��\�);���"�h��|#����7%/MqR��i�H-�+V$ �Sғ4���� /��"c[�;v��p,��$=0��aL"u�ҳFd�����1!!���R!���������4؛4����ݧu��Pzx��XP�6Q4h�>fP��2m�,P4��+6t�q��_��1*�8[Za`L�z㆘6fo�-l�P1"�鹄�}R��8�R��BCcZ=�{�l,Zm�\nw|�f�
s��q.�7��5��@Z��Jw�Nz���B^ŭS��Ӻ��١��fR��J�V½�!�OK��4b�9}�>ߣ?k�/e���O� ��Q5��FqQ��������W�P/��a�h��:���{��T'����[��H���)L��~�l�fP�W���s�膔h�C�긿v�M��Y�Ό�T�,�Ȓ�V*5X	t>wT�k��g�y�RǏF���/3/�|�Vc,�����/��/ʁ�o��1nF��;,B它���On��l3��k��5}�W�<��+�5zu7�'y��;�v�W�Gaѯ��8�7�H@��t=�j>,N���erǂ#�����>V ����8�WF���qj;R�����<qd�|n�n�:�/���V�?QIj�#@�=aԳR�� ��2 F����3k��Yi������R\�Zō�ٲ��hX22M�q�ڴ�Q�� ;h���e+� $�����h_"P\R�|m���������v;�����P3"�9����Wƽ3�����>���i�YJ��d{�ˍC���;��޴�X8����"�� -��r��Fr��Œ3�R�F1���9	D�����W��b�x����v�f�7���~��I5��9_�)�Dr��q�X�Wׂ0�����������d{ۃST�-��jQ��.�:1�oڎ5�a�l��Js� $
g���?��3���7�k �T����4�(�U����r_�Jf���{jҫ��;aL��Qu�P	{:���K�������t�+��a0��+eЈpg�A:D��i�^n�鵒�n�ߟWϲG�ɈLqT���tS��P-�מ~o ��*`wO���dMM����
�X�2��Ɍ�������4��y�����^VO���i����p��1A&�7�qP�,#���؋�eWa^Ĭt���'#.�j��kۘr�	^�nk�/&�Ŵ(vk蹗�����V�Գ�m�*��Z���R^6/�])us��x�O~ō�HK�v�t�����X���l�Z^�&]V�VF+҃�=����2��ￓw�������k��>�〇Aiq�J�oZ�:-�MP�"0x2���.Qg= ����m8����&�X�3o{�š(��4]�51�h�%�"E�$�y��#�x�%5�E��7��u$�`nT��+����ۄ��m�h�^b=;I�(��9����&��-H����Ĥ�ߴ}�?�ʴ�1��FQ�3��q�����Q,�Q��8e�
����
<rJ26�������t;3x���j���f�x۔��#_���疴^dc���j�?FFŁw?N��ldvN�˼�EW�֟a���K��Ա�SH�:���O2�i��a�_�&I�: ўK���T�:W%���5o���X�9���䥖��/��Ao��h@c��1��͵��a}��9z�?���[�#��Z�Cm����+�yO��|�(gM���� ��;�:�hk<�`p���\׌�b�ux�u?��⎨�\�ߧ��ʝV����"p��zI&����,�ϻ�rk���h��E��Z�~$�G���1F�A#̅�ی@���1�]�>Ё��b_��2�m��5��֋��\���j�҂DbG���3�lc6�>�Oc�훫+���@U��q
�]�ݜ�U:C�j�ݖ�,tG����h_ꊐ��
��؆����`�>4��4e�&�F�^���j0�~W'��W��)k<f2���ZY�m/�D�����u��+@�e��=�/�� ���5��ꛯv�5�?��;��g𬽫c���t�-#w����g�fz}H�5R��ƟPMو \��,��e��������7f��B��_�~fU��6����sd2�U��)1?ue�k4]W+T�9m+a��>4� |��h*���)�$ǜv"�#-P�l��=bX_������ ܹF�E�_^��.x�74X\^�M����-�rC�g�)sG���b%?D�o՗��8�6�!b�n�u5��^hU�Jɽ�C��Üh�@�n5Y���F�����U�֛�N����	�4D&cj��:6��V���3s�l���Ss��i\hx
�X�:9���,n�������[Sx��)I{�hL��2���vZ�X%����(U��6����dk6^!����<�C�ǝ�z�ư5'�K��A� }f��ʔhT�B��I�a�FKVS� IK��hQS�ׂs�36�"hۍ
À��]����!]pb�x%Ըi�1�N���h�bd�q����}߅�����X�Pw,���Dk�ň��mwԅ�R�̃���@ iv/b}dgƃ���h���Y���6�"$�����NU��_�,�
rf�󜭲�Z�K���.�J,֐�xRs�+g]ۺ,���U�Orj���6I����~���� Uv_���Q<{�g��F�5�Ƭf,/���;O�"_��R�;܎�W�L�����1Oy|��^.�Y|�_p��;_�J�nje�~~�k����sC���_g{[�1�k�f��Hrm_��s���F>t`����5�i*�/��
��y���3<���b��X_E�M}�U�tMk2�^��=�-I�¼�;ו�3<��]{M]�:q9�d/����[����,���&�Wv�E���Z} c�7�n�XpV=�>!,�`:CX_�V�->a��}K���bε�E�w�gl���2��*�,bav��|�Qy���a}�Cv�:+;�`[U�~o[\��ךQ�^�8+҂I����S@�����]���}ݢ�݉�Y�n7��I�M|zb�=�	+���x=Ԭ�_�{���f[�GpfT�
j��l�^�W+<x<�J!�db��]�ur0m��]�����~����k"\���-��6����������m�m�Q�V��a������TR���_��r��Ս�E�]�h�,ʧO����'cVL�w�ru����H�w2{��U�9������i&�i��D�9� �^Ќ��(p��������+��H�BQ'd�\~I����Fߪ��bP��O�3��4���c����r�~��[٤��f�30��,(ɾYN�>X�G>8}��Ιk����q��#�:�hP|�v���� �8�~�x�qrE�s l�^���8}bnc�x��j�cF�(�b�smց�e����˄yb�$թ�~4���.;-�<j������������I�λ�w��N��\�2uHO��v��z��5�D���Z��d/A]�'ډ��΄�*B-��y��wj~�<�m��bA1G�qMj@t�����.E���NŌ�YA�@���MK6��Z�B�J�tN�>�������6�S�k��|�.Z��a�A#{vD�K@����]1f�!�.e�2x����(�t��ȁ�=�X��VAN}І�"]	3��B؊ɨP,���
l��L��H��"R��+o��[��ƶE��9�%�S������՘᚟���4խ�dK����6촙AD#XJ�;;I�֒\�\}dC��2�}"���)}m$�����H��H<��J�\�V��7�_b�3��"���[ϑ,�a������Ym���T����s��q8� �J��O�c�.�j�ƃ��ȿT�s���J#Yj�#T����(tYO��똿�v�k��K�Tw`�����J;��m��-3�N��{,g�E T���~�'�|�*]d�W�!(�5/�����ꤾ���W;���n�t�����od]�*��T����[�����j�gp�a0,�E���_�O�u�U&O��qf��t.%'��3M��@�y� /�!{��Z���i!��ՠ�4���
�Z;�!0C���Sma�nDh+m���4�\ͩ)�oLϵF�X�J�(�ڣ:IZ1*3�@'K�p���:�1�T����V�o,��Vk�H<P�Hn��h�T�x�J���Nm
K���ݶ�Q䥂m�+N~&�`���U����9��XJ��ML�)�vMn�d��׊����.����>�a��+���D��y_>�V�^#������W:u(}����'�m76y0i��p�Y�n���o�-�~�B"��,.�M��<�{Cf�?�����3UZ��~�-���A��p���\��3�
��lo�n��687�����Cu�m������I���Y�f�|gT�EE@ݟx����R~����K�c^�.��兼۾�6ͥ��9qV$L~X��9�u�ǜ=�ONi�S�t�EL=�<KT�?���5 J�4�ᗱ���d�	�]����� H�`�,$ Q�ApA�̧s2~���b�����7hT�`��>/S�z��T�i���2GT��R�H�[�N�[�ΐV��5:<_T�0���}��Չt�(/��?{o�$���z ȳ�n6ɑL�'=��������L�9��<����� YW�����D�8<����5�8_�O8�m��_J�é3k�� C?ڀR��(`��_	�5��QG^=�U�:[X"P �5�3�+1�#"M<L������?ѿ�˿r�`U�{O?|���7tu}���x��,M�I�p;f���kEl����p�� ��`������8;���&��8V�&�΋�
�~�x�����;��$WfH�U `����3�B���c/'9z�� у�3_N��\rU�v��K�� ��9��VS��L�F:{1���h�����"l>��@ƼA��l:O���u�䙨cE�DqdO��-l'Q(T��I%�b��vN�WUV9
�MkUX�w��ԏ?�s$6���:��@(�h�_+3)��.F������@�U��K�mV�+U��j����,ρc����(�:P8�iƲ)GQy�J]�[����0\�)w�N���xۦ��X�FQ��]!��k�]���������Z�	!����$E#ZK��ͩn�z�fGS!��xx���MֿG9G���rO��S��������O�0�����*�Dq�X��-.�@�W9B1���w2%�lܫ��������`F���7mKykܫ+�㑱0�{s�`���^�1e��G�.��z䄋���s�U�f�z���m�px�PʟX��V������{Z_��c-N�Nm�P�+KǎTX�hRF�6��mEz�ט�7ƥ��W2XF+[�tÎqr?3�~�Ðݢ:K�}��y��ڢ�=�N{z@4ڂo1j���.�J�HCyp�8���ѪrFE1�AA�y�̹���x~��Z���� �ܒ��EIoG��C��#q]� G
i��.�s�ƫ����#�+�Q�[XA��b��:��tV��Hc���&�o��9ݞ�'V�h�~t��|���}p��0�A�m��e��s��y�+�T5Rd��T2]U�~ɪ�3rQ��r�}1�h��Qwe:O��B!7z��IBY��zދ�Y����=u(s�g���;�žh�J̫��uOY49���d#�T��?_q�����b/ ��2[����>_]���ر�D�`�%�lW������-QI���%����Щ��UOŶ�3oi��R�h��9<e"yd�V��RQuw��%M$����9�lE�pMfsZ�F2�/8������=�~'%ѫ�a�_�Z���ڼg"z��B��/�T
c����[�D#$�&h-lB��~�8.sr�A���@Ԭ覾��oޥWL~N�'��,f�؞����Vۍ�#1�0:i�r��Fum6Jt��$�Y����Ȅgtn�J��I�5����)���Gf�F	JܨY��?���/���F�ԓe 8�P~lA��9r��*}(�C)���ڟ��x�E˩0��	�%T��+<�֞��d��u�Q��9��Ƈ9O��n�L�F���
G�8R�:��	;����h6[H4(�=8:֓5o-�\u.Xy���P��Qo+��T�v�=#_�8=9efubA����S.w�"?�ͥ�7��ixF�?�]�lq�Q�NZ�1�S���5?�(
���^���k!'yB��x�+�piϮ�ԛ�R���;��m��� Ϧu��ܐ�����Z�yF���\1�g�)��-)/N�e�s�U��ŪN.�tP�s:��e�/��p<�y$s8ҷn�۠���_�pLΙ��/G������6�k[(���������_;��o4�~����������|Kɓ3�e�(����.�������9a����Q�W�p���'�7Uiʁ�J�{I/�0�X������:Pv\�]�|7�"��0�{D�6#�t��9tD���]+Y����5t_5��N��Z+���E>�y�g?#s�%=���̓�ʩKh8G�c��X:.	"["��l5T��J4Vyu`\���o/��m�J��5=p��#\��i��&�� ��������P�<KT����j�����5�.�A7����!`��00w����vr�ՠ��%�JǱܟMnSb���7�y�\4�͙l�<�J�Ü;/���e@�Nlxs�rzd�D׹jZZw�s�,�VSb��Q` ^�g�G@�@���Cszvƨș5*P�����}w4O2�<���c�N�}9M�8���~�H ��]%hņ����x��O��N��#Şⶥ��^$�v��SS�X��-m˨,�C��v<��)�>�&�{�=�N����5}���m>.���f�ZI}<v4��)�T�(���TVn+�:,��1����~E��[>������%͚95�)-�i�]���qd'���[,N�$�Mz@�M)���Z�N��Q�ف"�Ш�I�Fv�S����J��7��/��S�?��?�A/�f�&�t�):@]����@�Խ�-�c�i}f��6}Znx�=ⳅ���+��5�j�N��fcojv� ^g�$R{q촜(�2D�p!@װ0��9�衯��u���oIs�oZ�p���x1dr��6vx�P;%Re�|6B��N^X3��;u%䁓IjӴb&r\|���p*�[&Tl�w��a$�����9��5꼚�|����2���$�f��HӊQJ�AIj��i�"�+8�(&¡�ٖ;R���x،�;B�!�SB���ҡkʗi��|�JJ���"�ј��:lc��U�gQ�#��[��S��qD/��ǳ�;߾	��ז��*Cđd�E_�ʺv�:� ��-��[����������v�Z���Ͽ�W9�3&�ߏ?�a�ϋG������W����Sc��*��e��,3�� �#ssil��c��Y1R^�fh��g�	A~����a�l�=[8��V�P�Cd\Î0Tr�s�;��� p�p��=��h_8u�w�<0~����IG�o����Z􅕣6�_�#m�:����9a�/8GT���{Ak�Ƀ���R��#�k��"iLBG�{�����-G��(���[!�݈�HXuRd�Vv<t�ۘ~�)�C� q[�/Qբ�1���V4�s��c:���˞׆s]�����.�4���H���u��KeE���kq��7Q&��%�iH2���(�0:�Ly�M�Z�썝��@\�\je^L2�Zݩ�U^�te[s2aN̣Ny�P)ky�䟰C���~���U�����T'�yzy�ȹ]�i77DW��A��%��k�����K���t��'P7p���������>�셋6ʺ`�L�Cz���sZ, (���3	��N��˧Ǵ6V��@)}���N.,�������!�?�娊/QO��y�򙖋��iFxe���[����I���çS�l�&Rv��G*ެ��A��KZ���f�R���z'�W�++�-:��A�1���3HmS��
'$#�
F���~�_���Ͽ��~��t��3׈:�e�)��wIP�	'�Qfl�a9'@����;�>Q���7]�}��0x
t��Q����,j%Fy��Z�)�m�tt�s��<�f��+'878�Kj�3Jn
�@᳕z3n���3�
"aZ���6p"qNx�δQV�ٜ?kX�@aQN��B���=��ݤ���p��!6���v  �,}�$�\)��	�qIx̻�z�w�䏠l�s�VK�#:�g�KTL�1F�����!h�pB�!R�<����E��'���$<�jO}MG,6a�H�&Y�����o��A�o��59�9Q��*��zN���~)���/?�Qf�����~�\vo�}`�F��o�ſ�������;�{p��7vڀ�.���jy�����q�<��<��Lx���o}Q�R��㍐�8�y�����:x\F��X��y����o��E`�ss���=��g��ʯ!�}��3�b���p�?%2�Fw�z�Wz"Kł�`߱��k�����󋳴o��βۀ��!�i���������)�d�Q�R<�ʚ�yM�J�/R�d!�'Kv�4Z(b�z^L�	^Ľ8]�yz}��ZA���p;�&B�̙ܕ���Q:��lJ�'I�[�� (�&)���=
�k�W��*:�́�G�V!�|���;e�3Ya���ʜ�� �cEJG�!�e��t;����'XAgVҸ��S��e9%˪����:�o���^gN�?������P�6@��\׷���/�!Rq�V��z����X���=�s�p��>c��g/���Sz����
�=�׋�d/B�qy��މVƂ3�̶�k�h���$e�b�q����2���I6�# �4/q��3�I�=l��珬��ݞ��{����_O���_����tAMhV'��^V�m�c� @�2��~�N��5�!���;��*��2����-ćS��]j���3�mV���r�RHՆ2��p䛬���:��1�4y摉cB1R!�ºz�e��g)~�P���SZ���tɇ�.OM����VB�h���_<�:�T6���!qQ<���g\��V����~�����/���g&O���u2�qdݞ'�~�E�.`��*N�
]����"YM����=_iǄf� �&i�ߌu��Ay�X*R !؝��d�H��qR��+�Hx���X2�H���?�=�A�08l�R��$0ܘs�[m�zMZlW%�q��>͡�Э��$)F3&,4"e��tBj�P:��4G�k�@����t;ʱ[�8�
�*�-#v��L���U������ڋ9�߲r#}�c�����J��T�Be��BJ�2��h(�V��'Uj$��myt��5�h)Uo���^\�8p�(,J��F��o�����L�Ѧ'��	e嫨
��D�=ˀWE��e�c��{[ˑJ���WԿv�u8n�<֎��|�$��Xhs�N��(���O�5�p07�7]
�|�ï�ޝГ��@G��O������)�8��h_�)�oѨ�_�0�N������$�#2��1����O_q��[���i�ķePR��j��Ux����Ӆ&I狎zi݅S�9ݤ�5Siu�&p�V<'Iol��͒޾=���6j��p{��no�r^����P	B�a��ns���4]��(�.0�It�]�5H����
_��jYm�"y-wZ^*�r�0�=��E�0�t�n�n<�7?H�|���n�6nI��^����c��Y"rf#���.1~��ԩ�*����4��$y��ʆ��(�|N7�Tr8<��s�檔����}�����x���9�G��A8��2C;�iq�\A�pRy��������=d��	SxnƮ�{�Wԟ�`V�X��d����w�L�r'c//� ���;� `��̘�SGx�T^����5~=[�<�*��B���R�P�U���rm��ճS���Y��wsw%�.��������bqJ�7{N�z�{{�B�v�V/��1Rc�{� ��I�+^!��r&����~��2�����~MRv����St��A�GݓпU�8(���z�fi��|��L*=�����;���[��zF�d�>��d��L�d�<_\���މ�y���Dy)6�r>��ԫ_�7�Die����(e�	�E����mCz6o&*w՜g�uR����g�8�)�GD(^#+�x�cf��?z������`��a6�,;��C���1!\ҫ��7��#�u���ײl��&�b.���Gb�r� ���Zα�����?���_���Қu5�H����q2�ni�kh����C�s�:ƾ�y�Δ�s�٩�1�������j�e�n�z����ZI��=D�*���;g��I��b9K��1#<��1��
��F`rŚ��q>��.,tA%�S��H��{��z�H�ʮ+6�������r������s�����C�>%��>O,��M���q��Z��*@(~VT"\~�>(^=��9ux6D1�^��{�9�b�v�K�a��ް5B�;WJG��K���i�ߏ��G���SD��KR��o�oh����u_�d�v>k*���(+6E�AuU��l8I���a�(߀�7�5���0<P�a���p-�d�=���9�����yz]�*�$�q#M�9����$�ˈi�\_�W��9;[2x)�D-����:1�!Sll�Ļ��3��"9U���t���<����}{��][��r��V	�R�B��������cv$#�<:̎*&-�R�1C�y%����;Q�+����N���9M/+&Ĩ������/$��J�; �U�W6L�����;�'�+�Jȝ"�1���DG��U	���{X~jE�V�Av�Ѕ>J����:h�����ibG�J�S�X[0(��nـr~����>���8_ G������f͌�R=!)�$��"r�E��u-��2��q�p��^姦�U,+)�C��}���{��yk�j pt�^�L�RyP2��/�i�d	m��Z�����vb�n��6���$�u�p�T�Suu����+��W�Lg��nϙ"�M�ӋS�N���Q�[�}�ono�\�O~�H�&^�px4U��J�gV�ms�ىZ�<����h��-�pSkja���oF���!G�����b>�� ��3Q"�~Caؔ���W��H��Y^h6F+�#������}8��;&�8vN�2Eݠ��ai:�WN���&��m���ye��N.;{�����3����%ܩ�{E}���oV�5�A�g��b)Np���Ѱv���S���"]�9l���l��2�vC) ;:r�?_��,�F��b4K8��E��vT��<��T҆Y��.$��Nã(�<��b$N+�\���D��
gd3��f�NMq���L����V��wR>��ѨƵ Y��f-����C�gP�� ��5����*_-Ĉ�i�0�{ogCT�x���!���b�{���B"��y�ű��k�(��U�[Y��y,��؝�(ځB�r!����*�D�%�uʍ��
Z�BB��y��p����mߣ�pj�g�<�1X�3Ԍ޺�X��]���-���QF�p]�R���z��딑���=��|N��Tq!�՘k;��ۖ�� J��{��*���vrG�'ö����/�L9�Oc���9���G���6�i��_�xj5��V�/�:�f������X�B�C��P>�^?e8�b��k�^^���] �+ڸh;mp�����Z~�d?�R������<��*� A�(_�Nw�Oo4�bĞ�!Q̱/C�A/���K�\���o'�h�*$T�]A�VqR��iX�N��u
�.��L@a��d'�����钃iUȑm�U��I���p���{���=�xA]��ͅ�IEΎNN���<]b�k��C׫R��L�6~��4�6��W�w��Y�?WF�=f8R�3;�(;:+�Se�㪅�S�SǌI_�Q�"i�9r�u��M�/7B��(%
�GG�d��ԓGeVϠ�Wa�-^�u��h�av�x��V�����.�R%*�����| Ө����zʋ�;�(���2F���3����z{H�6i�|�� �+����Z=��Cℸ_=���5}���yk���B�:م�Ņh��g�@?��^�:��3n]�ϕ��xY��L����ǝdT�h�Y�*SPn����r��T�vپ��(k�̠id?�l�Pb����{���ػH���N9P�HS��YJ����,E�K�I���g�`�����3l�l�y���>��uswG��e}�N|T�
L�Fg��qD!U�;CE)k��$�m0	��V�a��u�Ӧ�Al�h��d6I�0������kDt�-�����O��Գ��!���jq�i��n�����ŠY$G�W*ި�:��.t$�0p������"|�҂��ΛU�S�yxDY���\��úQ͡W��08Y_3rFV� =���J��P��_-�E,&�zC�P�
���|�iMȏD�	����5�V
a�=0vȁ���\iP����g���2-����V��m�<�q5�I$#n�hm(>�ڌr�pL�/8�@�\�R���ZU��i��\rV��k2M���G��L?�*ͯ���$"˷PP��Rjcw�5-;�������=M}�p��v۲�k��vxT� �"Hy����;���Q!},�v�2��I����#v9�}U�(�hfl��Ĩ8�_�Df�3���s���kN ��W��b��[U	��r_V�mQ����Z-�+\Q叔$l��2��(���Ʋ���)����Ɇe��/�u5\_a��c֜Kr�J_�Յ��J$]l4ӉG��;��=��U�~��j�X
���[��b��v���W�a���L�)��37�/�V����9ɜ�]��z�G.,d��N,Gc���q�J�H���Wjo��g\MF�K��3�/T��SL���W��ILB��e{���{���_{�Z�oS6<rkm���v(��HY�:�6��9*2�~���y
d���l�kԜ��fcd���)�ޱ��婑�0�k!�E�{�uϐ&wr��y�;z����Ϟ{3X_�AP�O�{��!�AYi�X��V���d���OV%뤳�L�׊V�ݜ��GO�������������Q�{5Yj�r��  R��a��{/��Ҟ��6��S��L-Ġ�ɔ��`nN����nq�����]��'Hs�c��pd�c��T��5-O�x_�$�+���`�yV�kv�@��z/)���D� |V������-G�̺K}�bf�:�H&#�M$x���"NaR5��T����+�ǑƤ2�1����
f�TV5�2�HP�}d�у���4�0#u�D�"�*u4TP�>T�i���s�N��C3�G{�x�P�qZ�Cm�@�9tl�ĩ%f��krjts��o%�`W�YO,����>E�o?r��$���]c���o��Q8��gq�=Ѵr�C�>Y�\���׵���[~����l��������W��ƕ�k�'���YJUe�֎�xD�5�h�r�c�_�=�r%�v�����K�n�$��kv��A�ܩ0զ������j7�$�'R����,
k;)i����� 9$ �N�cT���=�e�ƜOvb�3���$ׅ.rN���w�����g�S>�Lq�f"L^*�oW������kf�v^.<"�T�m���Mh��F*6�=�I�:o$��j�9���X�g'4YLeq��H*Lf�mk��D�I�=~�3D� v� ����5���A��TVZ��\s.L*C@����ɛ�b��R�)6{/�r �-�X�/�W����'��r��";����ee~���΋EZ��k�?;U�yD;����gKq R���Y��Q���aC77wt����d�Q')M%�=��, �6y�ٙ�Ip� M)*�n:E�muN�f�0�%9�6mۊ���V��J�r�3�3��D��mR�;ut�J�Ϙ�'�VF�b����iX+V��~!��$M�0�N�`��}��f��2fļS�!pWSh,��RsdL6	)�jeG)G C�>R}yE5iLi:���<���umM�w��Vy�N���ΫƜW�n�Uf]��<�?�兑�ȟ��ga�d��<1?{��h��#نd�%�h.���86Y�(o[�����:�-+Uu�GzD��Pȿ�a��{���R	-�h�-Sx��mD�g���Wu��S�J-��fйVd ����iW/���Cb{��֧o�^�K��V�#<~���G>�?g,�c79~�W}��xf_eFvQ��,�(�L��sB��N��X�b��zW%[x��:��8�y�����)]�5�<z�ȵ�⎦F�_�����z��0YCq^�nM	�*��X�K#On�i�`>�9mV+Z!�;� ;Z-]%pŝ�ͺJ��6�褢�������`��`�H8���~�t��d&59���O���;�(�gI�
]�(g�C;�;���d��b. �A\�4#�Wp���ML��
���x��9W�J�<��B"��;.�Ѷu$Iu����_u-zWHe�Ί�a{�D6��_��\�A�o�Ugu�B�P7������9"�牙�A4�	��1G��K�9W(�8�"�������J��u=⚍���"�F��������p���7ƗǳCݖ�)BjxA���WG����g�:� F�]�eTP3Q�F�/U�m�"�pà�y���e1Vn�d�7��6Ku/�Z0�x�s1�ۻ�acb��)�E����F��������ncp�P1(����ض�91Q��i��I��}�T#�2Z�;{	��("vTC~w���Yi@����Lu�*Mz�x%��Z�K�m}#�k��f��_��ng�4I��lyF(�_*W%s����Ev�ٹY��ܳR�c�)�RU��ҕ��)ą��sq���8ı���� �Jh^EqjW��x6mb�q�!���zź�(bfA�� �uc���A�D���q�KT�
��M��7�L ��n���Fا��!��}2�뙔�<�jE���~Ҏ1ا��D�PI?w%�E�P�t(y�|�UjÖ��[�9k�&�@P�� �+�@MNi�P�S�3���&�n�d!"���K/���/Q�N|�S:Xh�?v� *�O����N����4dTǥ�wkJK��QM��l�TMZ ȳ�z�S���.-����3��=��"��c�1���&dQ(@� u+Tp(�I=�b9gG��r.�sf�W�D~�ù��4[�V��^�i�6 6�n�m����v�m�׵i�Z��������=לf��������x�-��ɜs;Q"�-R�n��놑L;� ;�e7�s��?̈��AE
%�3b��J�׍��3�X�92���]������F�d���R����Cn}�7-S��bV�1�jfA�f�۪�<S`����|Ve5�PO>���3VK���͘�ȑm���������E5	�(Pz@5��Z�/�tR��0_�_[���9:$cT�ԃ�t���q��Ì��#猽��&�,���͏��c��=vk�u��G`�1�N��y�����3���e��o��O=ܨ#ξ����U9Y�޾��e��b��}�����S'�\��)��d�}�y���Z��H!��Q∤��{���I��3:9=�=�&h9ZAawZ\a����1��=�'�0�n����0ܱ���>���D��Ip&��.��t�i���Y���4I8��i�YIz;#µ���V��J��)�����-���܇�o�{mú:�'�B� ��Y'��OS�ˬ8�M�X����r:9���J"�H���R��ឋS`?3d��]�H��h9=X�TA�"�wò	$f+��YΒ�=K	��Gv���b%G�;u<�ձ������KYc#m'��FF�Q�V����r���	�#�d ����U�\,O��Z�;����e���8�-�nmH�`�� ��Lw ��	�1L�F��>/��(�΅���2�P9�s��D����߯��[��O�a����^�� =���/�J��� �:r�pf|��Q�p(�g�~�ZH2�Q�p�����L�l�ۍ�$r���Ew�V����
e��V$M�j�6E婚+"
��"��n��������M���N������Oϸb�������`x�r�Ӳ�����Oܬ��7��N�#j�)u��`�A�a��ܹO�3l���[ZoWL��2È�k��<6?P���2����R���I#6^�\҄d����NYӑ��*	/߼�8󎥿������'
�=�� ��M�Ͽ����d`#N�ެ����B��0�������H��������J	:(��i��Y��Z#�A0���٦L����h����R�����yvU�2�5�D~��k!+J���S�!�i�!2��XIX�}�VR�҆���?�w��o�ةs�<eE"-��_��\	���u���3�T)� 5e3fe���0�X��R�n�Ԧ�D�o��l���-�"΁\����,�	�#`\-��\{�,�|T�e��f�U��Oǈ��ՆS��94�F��Bz�{���n�o��N�J����qvyJg��uΕ�P�A	E�`a#�X"�v��,{!�vT��xE#UN:�YJY�U��(<C�hU4��Ǧ^/�K�L�r�u��U��Ȇ_i��w@�7
�d�tW�TZŅ�i�1s��ˣ47���AA����������|d}g#�.b�=v���G�y��Y6a=N�*su�f�NN�����Ђ'U�L?xa��z�ƣ"���/W��F�?s�G��G���'�nX�fXD�k]�O9hm�%9��ӷ>^��@���%���y���@{ĵ�jg������Kl� �חL����n=ђX�{���	������?rB�ɞ�	���Ze��������A�6�XA��pA)j Y��tO�rJ��Y�b(�N+��&6�M�� ^Ƈ��4��^P��/�@?� v6�=ԛ�C���9��.�]��r2�eǩW�=�I�A(�XЧ���L�>0���FIG�v��(����	u�	*�r)Q����5L%-�N��d�2��̓��Uoű=A���n?w[�D��V�S'*F�M���s�x�X�6�����KgP$r}D���rsRfk��4_J�R� �{\
��}ϖ@h��ꆼu�!�U�i�˨_�N������*Z�)M��o�^gNu��>&)�����2]�v����;�f�۟y'�m<�w�K�#� $��o���1hN��J�<��?Ze��5����\Uh#�E��E8t]o���S�S�3[9�lMa-5�;`3�^�xζ'�X�k���t��;h�	N�١���Iv�jp}ɃQ�e=�ǰy@�䷧�t{˶�)ȓ�����^����F NFuh�Im���v��B�����t�X ����YR�P"�02`��-�%A���#G#�_~9'�	�ޠQ��0�!�&\^tQ��ج�Ք�SI��g���Mꀇ��<����TwG�W7t�7m"�@Ģ�̡P��)�9|0@�BȠl�"�s��j]U�i[Oyp+6*=!�prr�{�Y�S�E�X�'��"�v�i8H�a���s������U�o��!Y|Y`G���O!�{�&���)�_��	�L����)�	����YI�4�W����!T��`����vH���M�F�8c�O�8�(޾��]�)�4cQC{����^���AS,j-[�1f%��2�p� &ѰVs~+�8F!�唰-�c�h����2}��ԋ,d��(��ah3����==M������./�p1��usK���;u�α-G����`\N{��1|1�;J�4�R��~��"$�Vu�,�b��\l��֡r�r��{Ut��1?�ߋ��QE�:z1젊�|��D��@e%:mANy�ږ�;�߳�e�����}{62>����n���o��\�r�p/�/�j0�{=��v��-��uV~o`��`z}�3ǋ�H� 粁�U9��񮯔��Pol ��c�傠�)F�hnx�C�l')��mf&�ݣ����=��j���Z�����Y��j0�t��q��H�I��S����X��ŧc�iYOػ�{/���� ���u�ۛ+n?�W@��/{���ћ�?2�0����V'�3z{�mڷ�o���������)FVJ�Ĕg�����4���[Z�,���������PZp�����A@�#M�K:=?����.��/TI׊tM���mk��f��PT[�>r������>a�գ�@����⪞@#�l��JIHɟ2�����Q�($�ʷ@ٯ�W���<>���R�u�y":
�,)�ε�m���`h���>��0�����kK:J����Pe��'�"iju:ϙW�r���Q@��T~�R3�U���ݵ�=��շYD��;�����a���,ч�ܩ�F'I�s��J�@��j\���q2�҂ ��^K�	��-�9��j�k��t�X��9_���{;l4��u�q�9*^/O�SO<�:�K�#C�cvWN�o`�%9�H�\���?��?��?��@��Ӧ$V쮆��du�ڵ�mx�p�tu�K�������ݢ2�~��]���-3]�p�@�u[�[��z�����_���>�%��g��T��I���������7�L!�V��/W����3�0G[:2���uIe@Kk4hT���9���d�6HŝṰƄ��QV5�s����&��ˏ���y>:!���Ɯ�N�<{��Fyrz�^ˤ�֬p��`�TR� K�nr��*Ԝ�&+dI��F�&|����n�`m-�Mb���s���^Ӱ�,N'@u)�A������HyH�J/�̚�AF�at��^]��k����/�	�6�n�A**p�K�����=;T C��B��i_l�0I
�&���u��[���&���ٱ�ΞQlnM��J��Y��V�U<���֜�H{f���^t�Li=,=����"�r��6VR�%�ʖ;uLI�|��|�6x�⦳����5�ܯV�m����������xsI��I��ӳSZ�{?��t�������H#6Iم4�0�qƊ��Т#u�r�0�WǕ{m�)X������f����qb��#U.e$=ߌ� #�L�F�*4����WiT �2�����N�2��x�~JV|�z,�0��k�G�сi;��|�ߴ�qEMF��ݥuT[�C����|P#������%�:��ˋ��6��a�f��>u��o�'}�Ô~S�s��lޱ��=��5�袠�!����Z�;�ޤ��6���W�ġ������G���s�����z�+�5����>���Xnً�0f�N$s�9)��~��16iF�c��H�{����Y�t�����_,�[&�e�tD^�h(P��ۛk��B�0��s@�Bw��@)��K�A�ަ��3�0P��m]��
��
	%%�|m8�a����T�rN��Վ��nYW99�t��Ұ%��w�>o&+!D&-=]<0��-�;I�@_�p��?�Z�t_��#��#�zss� t���QRh&D��i�4�������f ����I���Pƣ�sG��P:�ԘQ�������ߋ��0E� �������#{zPv&�W<5'���*���03i/�O�Ϋ��ET q�?�s}Z
���X[���~{����"��u����: l��0P �I燱��ݱ#�U�+-��v:�U~�$�ȷ�{�4���s�=�����v�R7.�'�}��+H�:<!�8�G���λ��rqJ'���s�)8]�_���x^����_~��>1� ���B��o���;v���4R8v�&�y+U��p�7�V��pCˏ��;��
���թ��fdFw�I��f+2�(�}��	�
Y�Eq�b�_��;���'z趴J�ϫ�x�A���{ՉI
��kr h�� �w8�P�O�"NT�~�Ǣ1��|В!>t6�ǾmF3X�?�1�BOѨ�|Io.��Oo�qǓ��rǋӝRG-��������qu}M?}��_6t��A�_ؤ��\����#W0tU��W2c!R�) �"j54͑T ��-熞 �$��k�������:]vS�j�?�z�2��
M�Kh.���P K{8"`i"���%A�	�掉X3q���ÉD��1]F��@x��$&^�r�}?r$�D�mV��-�k*F7��e�S�q�U�bH�:�<�$YP7����T4@K���i����U�euzp�-M1���CN�J�uzvΊ���9G��>D� ��|}G�>|d�X�Ǫ!M����K�R����X!�0%K�8r��񹠋x�(A�8�r�%S�Y��T ���?C�pT��ǰ�CR�r���Si�'�3G��N����Ƞ��K����E�]�Y����s���*�A�U�_�Y�)�;��@��O�̑4��lܶ��]>���+�64ڿ�L�]u�C�9G���^jve�T���,�D*�V�G�x�<:�c��]k���l>��ݫ�7�?���x��ח9��QvؔF��\��1��({��17�iYK�{�8i��K��$J��K�O��0�kU�✸���p������x_�\ul@�oE���V�_�V:M�ug�#�{�<aDF�o2�d�DM��Or�#��I�:�:o��a�F���7�bv@���I��^(@a�BA�Λy�Z�s�PEҵ�Y,���@qV�;��m7@����z��u��-�M߬8�zXkڍ:HP�d�*2��~A�U0rc��� ���o���y�`e�Kyj{kv��.!���sP�eb�G��.�9�Ю��.�=��o�Q/h&���YC�m����:�_���e��������t]�JI{���`���R�� �:V��e���0�.��R��H/�:#��i��k��P��X|��e��?�a�U�~��윟����?����Qh?8���F+ 'y���m	y�%��U���<@u*�B��+
�ȝG҅�HvN�n#�_¦L���"L�:R��0����nn����Y6�����"yTO����Y��1�n#�<hp$�x�����4=_0���;j�B��"#ZЪ��(R[O��O`��oa1]�T
c�SV��-RG��\�z-C^q�!����d�"�i0./�����8v�B���I6�3f�F�aq`��U?L.o$�{��ߘ�]�Ł�ˮV_g�XdjD<�N�LL���;��a�J��`4���T�3iiR��Yv"��#��7�Cn��%FT���7�/�3󸫕ś�y�a��q�b �}����dɈ�����cSc��^�dr�L&�� y��h̥��#s�V�=1k*��F� [?T0��Q�-�2�z'ʊ8_�����eB�Nc?����8m	���^��8C�T��K~���,����A1B�0g��_]�q���{V��9�p�ՔUT�\������D�p�/XĩUԝ�8J�q�Uz��R%�P�C�:K3)f�8�t1�)e�(�uJQ�?6���������6Uw�|4�X�����t�ͻI;Y���3^�d�XIWf�߷�++txJ�uű9�8���Sz�T��E)(E,����B�����G�sjYV^�w��%7�Δ}����O�h0O<��>Vpw�Ur�rnħ�Bǿ�m8~�ɗ�=��f����<<vs��#<u�z�p�}"�(Cϴ���,�����܁�e�Q�Ey�B>=䗣�oK��unP�87.�#ܹSw�����ȑ����;%���z�)�B�2�0db�u0������ao�����}e�P7�{�P<@�Gd�p��c)�Z��W��=���$�ڒs��\�D�b}$���?���J�ņ�{�h:)�8uV h�b$�N�;lD�C��B@o{��x� m�Zˆu]<8������9�'��M�|�'H�?;c�P�HAap>#5�d��@�;s��<I>m+�i���4Z��̊
%��M9u��V�<�
vGM]�}�/��i՝*�ʐ5!���Q��Y�yOб��O>��ݽe~��x��8|_� Ϗ���q���E6�u���XϞ��p=���W�����Qi\L�X���T�=��h_}�ί?��;:2_�x���s�9M�dR��^���ӟ8c�4��\�p��w�3v�lο������?�B��Y�Z���7�U�}�k��0lS8�����D�sp�̫9Wq�̂��V���Й�\�r���<]�J�ؘ�g��^����R*�����oU6c�R��,�+�
�N��*�ǵ�Mh9kI J5�U�z���hZ*I��z�i�-��z�6@��-�'�û���#����荴ql֪ ���n�y�ito:������0���ҹ��C鄢Qd��%[U���Xb�G�/ߦ�z��$����0�-P;<���I*�fhn�6ۭ�S��#%.��I����ܱ���VR�������	A�^�q��B$VQ�V�{�N���(��Ԧ�T�Ҹ��v��P��b0e�i�mb�k�MGVx*��Op��M)��i���8$-�4���f����T�:Um�d�@��`#S�a��1c�JQ*�`JO/��Q��EZo%�����c�MճP�
Q: ���4��1�?og����\����$�-�x������I�u���3KI���%�'�i�h �hUמ�.�F��nJZ��V �d����	��R�;_�鉨������Gޢ��ڴ����~3���k{��!h9ᘉ������� 
:�āg��o[A��P��$6�P�_�{�W�?�O���q�s���c^�Q��1#4ݠ�HD�Љ�O��	���;]�_P�"X� j�42�Dst�����2�(�����l�ܖ(ϲ
�������ȉ!<q��w�H�$~�!��E��A^< ��9T(�GPP��9�pN��Q<��v��M��gc溧�y�֨�Xdn�\�Tր�������^"��	����K>�}_��ﱼ^�y\;_��6�'N�v$�{'*�ԵD4�]��Ke�hp��D3�n��
��A���t����pz�� ��!&�R���-�9��S���DZj@T=A�~2�Ah}�v>�Y��Y���ۤ5��z����x�<_�uvYW��2
E��*A���i�*�Z��==H�aLМ�_����r[���z'�I�����3�q�u��0�`JP�*�f�]��V^�t1���0�+�S6_�1P[��k���$����/7���{�t)�~\�g���5�c�n��#��1ΐB�ܰ�*������q w�#��ֻVe�b(/��xv̹�龤��x�LK��)[6�Эm���ǾwL���-�T���������/Q�|�}+��S�mV�Y �s|9����A1��3:�-h
&ɣ��2�˝dN$���p�k6W}J2h�d���_vu�D�;�A�֌�IٲSUa�c����i�t��rF]C�=�d�Ռ�Wd狡jjE�q��hr�@*�����Ssl��v���t}��%ه��EQ���ʞ�S����a:��8�Z��5��aHq\���;1�����h�-�GZ�Fm\^қ�o�m2dW7R�y���^4c�y�+�=+!����䔣1�̤��.�R8�"������5I���d)%�HJ�as�$�|���Ҹ<t�jR�/&Nn�i�G�t٘}Wp�$��52e������hGđ_��U=lX�b���.g�D�T���K��j���^ӱN�i��o0�_^T|J}���E�9���n
~����(F3��v�,{�U5��
~q:E'����YBh�L�ik����n����fl'̛=�	D ���z��;��������~]��vu}��ҖV�-�'��W� ���
9��9�(���{��'&�ß���EK��W�'-��E>�:H������%E�(�ĕ!��z�.U{)T��9"����}��,���Ǐ^y�s�p��^U�P�m	�![f����rK���jT �
e�T$rt����zҲ��ژ�A"]������V<6N��Ǡ�z'ƬH��0\vÌƱ��wqC���ڼ�l#�N�*�:>��^�Qꯅ��?�h��5ƎR��_��;�ǯL�K�]��_8Ǿ�rj��R:w��� ���+�1��pp�c�}�Sm{o��5��yt���s(�L(����_ÔZ��ϣ��7����P�1�w���M)O|����|�mþ�Q�U_J�r_����=��6��ߋ%�Gq�F�DF�±}�)5p͸����9�R�#��`)��j�.jŬ�����hp,���� OR�vH�Zo��k�DnظTd��w��ƳմlC�p!
#�:�6.eL��Ao^L��b#�s����Z0B�S��S:���&�Z*�2DO_����t3�7�@����"��� :�UX�L5a:)Q�=8e�sF�Z��,��Lv�����-W�yUp?���G9_'�o�z�Fǡ8~t�#[l�����Q�R�Ϙ.�gZ�~L':0�;uF�R���Sؿ�?8��a[�mߋ��F�@G0�'���Vt���s�ug�Ũ0#�rrG�$���dWwl[�d���<�;����&���!{����h���фڋM�@Z>����}�nK�fF�$7&�'�;7��tw����cg�U�?�T;#������L�o(f�tXv���9T���t�k�@!¿�ua�&I�IMo���Ux��U_��m�=��D~4Y���MU{5Y�A
������7\�gyzJ������?3�>�J� 	0����;�>m�]{ǐV����,�@|h|����g�P�S ��Ҁ�y:�h Z�v{&l�M���ϟ�sz� A�H�\�z��ӋԾ�4�P��h�)Hڞ���}�����"Pe�?#A�E����@� ߇�#oꧧKf/?==ce
��(�����&�"B�[�;��XU��OL��
�qG�j@��hi(���F"�D�Ba�iʊ��Dpp>%o8��M]��s���^=��Lg���N�m��8tN���s�{�����N�M�U��{F� ��D�j�y��
��\_���v��Hv�"��|S�lL�LBYT�*�`����;�S��:�ܘ�V�wSNCq��e� ���[7�n$"�%�ԑ�ȕ-�z���-����̗^�5N���.����D�^Z娒�s,�@:'�C�$N��H�m��u��gt�^S��X��N=��8���C-�f_:vJ�\�_ƕ�P�\=b�����y���s�g8���j��è@襂r��&��wzT�_~��}`�(֯9w��2T���u�������w:L{�L�h���,�F�QX=��d��p�%��yA�	��!--Fҡ"�F ��CM3�ƍ�;DүX_0�!�& ��&��Q�-W$I�t*	�&NR^���{A&[��ʷ�N��2�D�����'�q���	zד�ٱ�oT6�I�G�Ą��/.Ϲ�*�����~E?���͞+�v���J9R�$�i��g}˜'�
D�7���� ��{��R�!_�xEE��5�M@�!t��&fiԻ�"����8���A3{��:K����z�S�Ͽ�,���9:�պ�m�,K����i0�+��ǎcz�ˤv$��뒆v�ѯ���>�w�Q�D2�c�������;l��[�����;���K2vN���9ˀ�a�W
��X;He]�s,�\it q��8�SC	���z^'�.Z�1�q��PWG��w�'v�0:g�=(Z���1]%�;�_/�/���+�y���������oAxj5�u��P�
H��n��C[1�L�� G���b�Gwb;19v�6���G�<��h|��(9~��+���R�%��`�G�<h?��ÚKM�d��oؓ�F�p2�1@�x
2%�U���f�Xu��n��ݏ������ާ	�~��(�v}C7��VI�@J'�� �K�ri6�p^���1�w�X�$K����/z��|jL��p��!���QDZ���R���<m,���!����|2��>��F.�y#�"Z���Kd
���H%����h`�X���ȋ����-���i@�isg���Z��yH-�Aj�y�^�9n�w��ǎ"�[(E��	���.�P@�j#����g\�a/2�#{3mq���@�Ҏ�l�oD=�_�~W��YE��Ү����OOI7c�\�}0(����æR��k����s��8�sŹ���z�2�×��ý�y�ѣ�\���-�f沰5(i�p�������UeS"��V�D�Μ:�u>|���r�hsp⋔�q�%jI��N�h�5h�n����#�.כv*�3t?o�F�)Q��@I5������f.��)�;C��Y�Л�Cg�7>��I���o�	e�V�|�Q�:��S�z��ƍ����s��4g�V�ToW~�ex���l�F�}AO��������N�i�NE�

G�����x
��=��@]�%�`� �.�V��}hB{AǮ�]���&��Rĕ~'��|@^&[:�x��*�p�U� �p�{�~!1��"$���abN��_��,:W�=f:m��|�P����߃��z����&#H�j���e��լ�@���'w�[Qt@�M\6�>��V���W�]��@��"Ʊ���}f��uR�S╿)�m����vK0��R�A�x�A䛁͉�G>z<���N�sNH�WLv{�eo��"����$��H�zz��_bp~�#}�{�r_�3��vv<綁� 9���MK�$���	yjE�`�!߫i��W8ܓ����`%ӵ̦<O�Ǽ��\<���>\|�dQ��M��f���nG�݊�iMm�!��{�����6�k�U��Y#�I�?��]�}C?��O�����g'�B�ɆE�p���!�3�;Bu��^p��4��˜�9�� *�c������q�sU.u�r�ߖ�¨L��r!��Ay��|��2I��7o��,8I�Vw<�H���-�Q<m��rJ��[���ч��ٹs�:��4��o/����xx;���eيy���i(i ֛U2�o9J�ݧ��S��ڵ�������ڭ��)RXR����B�DjMj۾�
P���]Z(^�{ʂ�0���2�M��M�>��c�Źcv��+Ht
=rP�7�o�w x>}�H޿���1۽TrP��EO�Y���lU������T���:(�>�c��7g%���e'�+�Q�e<�=��C�~�i�~N��5L<Tшtr6�w?�a'�y��x8u������*��MA��Dy�+�}ge����MQ ���纼}��_�UpTY�h+ {��0��^�U��������"�W�(�y���oG�d�)�SZ�E-M*K�f������l�_I�A}5(���@A�*+�~z_p�0�h��̎�j�]�TC����q���P�$�K������+_[����?}lsU>+I�cDwJz�(�[d�|E?���i��l�{7���x�>����S�g3��~�����G�F�֥�1�s��Oy��*��P�N��w��5�m�p]蹽b_��c�B��BȤ��� �q�zuI�8��B9�{�Y�'Z�hȳ�K>6�$�eB�W�9*%���@�p�P�j�V�#
:W�&��uB\�Q�c�*9� �D9��G���Ǿ�Q�	Qu����DW�4��,-:��ͺ+�Jm��Y���ܖI����tFoޞ%}���Մ��}����;��|ˎ��S���i���9���/Z�OR�'Hln�h�b���42�R��ry��xȺI�*u��R���W�OMK�l/�>G�~�
�T��߲�]rJ�8?������֗���Ȏ��,U���f{���Ƿ������(T��{9����l��l� ���5����L�ʸ�#����Ked�v&�	��b}/N��������<jQ%�^��Hw�W�
+8p#v6�M���i��D&W�� y>�:���9gAN�SF���?����\}����dǲ�*��@�		���v��²z�k�;�OZ�
Z�'r��|V��ˠ�A���ٻ�p66f6�<��#��ّ���l������<����e�V3m�3�a�dйH}ځE���xT�����"-ϖ��.�$Z괚k�[*L������G(KC`8k#yi����4�v�� �dM��bR
�^��z88
��, cOШz�N('�I�;���}��F34��';vԴa'D��D������778����E�Y_\��^+e�Z�F�ߵ�d��a���JP���/C7h�l�ϧ����J'3�TԲ�������FgJ�F���ڗ�$���0�Qb:i��s~~��ȷ;�W�⒏�C1���-��>Hix�7H��h�r�	.�UD���-�R#k5�!�5�F��>l�ZT�Lq*���t���AŜ)��ý:dC9�z�-��P�z�%����]�_Źsp��]'�[U}����q,ۘ��#r.������!������C�e��#c~n�T���:Gr��p���T�~���9�G���ا�d�7�ܹ�瑹~�r���oOqM]ʝ(ds��T�o���>��@��D������r#�}�Z	�?��j�VȊnoޔh�8 Y���srj��G	�Ћֳ�ݢݱST�t���q]�s�������@gAy�	���K!	N:�ٙ(�\vw�r5��F~�?�I�BW9��H���=o�f2�P�uo�4������Y+Q(�zUMB���C�H?G:�vb�Z�>LN9k6m��d9�{B�A�#P<��n����5;u6��r�~h���`P�F��HY���3R���J����s�%B7�VH:V�~W��m`{�E����æΎ��.�:r�pO���vy_.E�����u���x<�E�����Q�;+�_�c|�a��ˮ��3��s�e}���ȍ��,z��߷9���8z�1C�N�1�p߲ã� @ڀw��_�{&�������TĆ�6#75��8��l�~��o�k�#+��S��$�������v z33l� ~vjw�pp���T"�
YD7�p���6e~�$׸,;ʹO'�Û���{ �ϻkw�^���ʓ�ٚ0�%�g>�Q?�9��D��=w����MIS�{�s'�oڲ8AI1��,�d��rN�����͍4�
R�R��=�s��o�6��d�ߥ��3�^䜷9wR��6�lQԀs�X'��ᳮ����Q�P�6�f��7L"��ۮ���N�ņ�9}��+�4��A�@yC=�����z��M�z��-�֊��"�?-q�E��e��T�_�5)B����?��Q�����X�����h)�z�{����^rw����Ar)�i+�>R���N��*2�"��T��')��M�N*BH�JKܑ� E�!ٴ$�e���q��Ӱ�v�\�9��y�X̘���s��P����O\bN+� �Z�&BT��B5��8���Th=c3 ~r�""��K�
�@��*Z��4���tC����94jPF_�e*�z*�k��W���\i/�����(5��#X���+� ��Ąڕ�C��w
{��u�ѭ�(�!ĩ�,�#H>�t0{/�ν�C����F���w&�����s�������}�pRe����!���@ź����ԗv��� ~z{�~�7=X⒥=>�a������Y�3"G؏-�r��׹���D/8\F䇏�XMyF�^��1<kޓ��1�.�S�:=���ɜNOϹ�e�ĺt���~}��+�T�cy� ^�-9��78ض�h�8�:5	B�;�I�v���s*-^�!W8��|@�U��`蘖�;%L�}� �Ym�ȠA���w��!��(4�L����9����:F﶑�l�݉\g����a{��m,��D�9�j��7Y.��'j&��G&��ʼ�8ez����x(-P!�e�6��s~e�k������R{��АDE����c���~���W>�.,Ob�WQ*�I�x����"�������2�P`F���=̐,u�g~�>e\�a;0���8j����N�3Z&9��X8r�4ɔsMs�j�+|��+&�j��u
�d��p�#�?�.5��I&�\%����@����$�Q&����L�ܜ�P��S	��N�#ɖ��������{�M4G�'4������K���������=A���/����r���������m}��x�K�k��eո<��Ԟ%�RYΏ�̈��0�
V_$�R2��+��������.�(���"��0��)��㒊Վ�=^<x��;������oN����YaL�?þPB�U!B�vZ��##fh�F�9�dn����\����~�[$gly�+fLgoLz�3�;�Kέ�c0�G��Q�Fk>���R���AQ���`�xwd��8�������J���ӤYIe�L��ک�����JڷA��G�����?3�Qv�~DU�,���6��=���Y�32��T	����77���H9�kZ^"�
��
i>���I��Y�ЬX���k��f%߱o5P �+��^Ʒ@Z
�g�p
����vY���c2��V���/7������k���tVEqU�|Π��[3*wFO��c�o��'��T�>��3�RD��oҨ�D�D�G#p�+�D�Ȫ�;\���f�v��s^��;Ͽ��G�M6�Jr�ew�N�3C.�ʱ��]4k`�䴳Ǟ�x�/�-B~����g��8���`j�U1&fm�������K�{��_�zdTF�w�(<�{=��/E�d�ad����х�04�#;�F>[_�o{Ս�[�|x��s�,?c'yȁ!������
g�1��*b��6S���S�= կ���֓�?n�o�!����ac�nY�2O�b�E;���'g�r��"����+	lY:��������B�Y�1tmq��XG;;=e^@�e�m�N&D�����'s逛���.��:��G&u����y`{�\(h� ��D��Ja-h�ά.�a��4�h{|���{r{�+�������d�:�rZ��DYK�wN����3������&C����u�:���X��o���8�q��������0�{�8�F�����ԕ[b��3Ƥ|�yxŐ63�˞����q�A!t��T�'���5MP@)�'��+�(/XF�0������h쪶��o Y!�?~��h������թF�>TN��HBJK���J����N��.l�b�߷R=5��­ّ[�Euo�x��Lv-=��Wן��no������K��8�+݊�c�g!������F:{�o9������p%��t^u|pN�v6�5J1Fb$�8x�؀���{��.�1��}�S�i�Ӑ��sB���	{������;@��0`ؤM��Y]~\%�͐wq1�
R_�� ��[v*qy�錿���
��6���_G'Y�U�ܫ�>.Ҧi[pJ�n�D��L6���GF"fˆ�>���/��>#���.�_��]d�D�K�S��a#��>
ϥp������޼��>��TҗXy8?���~1z�~%p>��- GeAa�η�Jus���gC���,�ssRU�$7R���̝���Vx��Z�Sg��&=��Q¶��ی��O鹷{�b�#C����6E��\j$w ��U��t%��Nb�_��Ÿy��v]�@)q��|m2�V��|G	?v\i��fQ������f�)Si�a�T�WK-��z.��KG�=q�p��b��j�)we7<�ߨPL�p���_�
S�^(�Rѝ�~��rJʘ+��8�����q�#�cΘ�L��Sj�>*�c�xB��
��4"�����e4cn��i5���5�P�P�ºF|�G/-��'zJ�}m�Z;�_�i��FG���S��/\�/:���s���0RIP8e���=�ha���
K��SIVV�	Ye��ٹ1柶f{�	Z��9����y�TqO��z�0&�5J��<-�0Zu6s�y�r����� T'�����a�A�o����lq���ٶc���H�����ڻe�-�Ֆ:�4cG*W	��3u+�f��W��&t�P* E�@�v��꺵�\�ځZ �����O$}<0�NN��5�"�{�S@�ZQo�o��E2V��l�t��3׬�YQP	pG�:����D#/b]Z.��yl��:U�J�;�t���'��\F݊
PG;�R1�pÉ>���xjZjV���\T�����w!��i��L���1���]������e0:1��Pl���˯u��|v�VG�H؉^��(�vDwS��8� ��Ot ��dz�a�L�uz��/����/}[�X�#;='K����@��=���_9�2����nonDM�R8i>K�#7�2��$َ�����{v�̗:�<�	�-'�)tH��#U��fc��1��	Q�-�̩�g���L���v}}E�U�Soo�׿�J?����^o��@?��3W�~��o�������O2]�s��{ ji����ꆜ�bvkg� �kq��]�G4�����J`�����-:�|C���Z�Y	<�<�������ruw�eb�$�џ�b�ͥm��TU�!Q���R(6޼�=u�0�
d9�0d�u#9�`�fFn!2�H���/@�N�7�\�|�U��-sj�A7�����	G�^G�n8��ؙ�eY�o΀��4G����L*���6<~+T�Io@���3V�����^.�[yB��[^� 6��6�$A�L*I�o�\S8�ȕ���N+-X�J����YyPcg���k&G��8p"�Y��@N�JJ����6piԝT�@:��直�W�W��R1Õ^��éJ��@�xb�{���AU�b�
w$��K��"�^]��#��s	�gc(o�;j�uUX��I� u�������}����r̕�±��YO�C�X�]�\���X��0Y���<��0�L��*�/4����wO߳vơ!��@���a�zll�\.W�
�qq 3:T��ȼL���c[_�x�����~�����G�5wx�A0��j;�������#/dH�#7~2bz��G����r#��/�!-�ں͆I���[UD>����{�7�$� hD�r�3�������K����骒�h��y�e)�i3�-�U�HH���8q"��]|?�^�XJ���9V��\� �{Ooi�־E��k��T 
����<O{���Y���j8zg��[&I����ȕA�L�Yթݫ��
�|1�E�F��D�S<h{&�?�3�n3�Ҷ��J����F�B��fSr���|´	��<�ΓA5�"0>&L2h�^�g�4r�L �ڬ���Aoo3���6W���S��>�LO�`~v���@e�8Q�l���+�U,JF��S�l�7@�\���쫡?�jl�\�FY�
�{��C
�h����8�Աu�8h��x����x��q,�S_o���D?=������gفy���|xd�e�-N��ຯ�9�[5�j�V���G��{ȡ���6�÷���(5{�λJ��s��${@�4��Lm1���Nt��� (4��Zeh�ň��
��*u�Y?��*#��[��$��!t�H��!�Ś�������)����4����D� ���BH��l����*p�A$��L������D4�3���F�L��xxm�������iI�?���>�g��}zp<{�Ax�(�AU�5�<Cd69�|�0�@qE��g�3J�Em����FCT�{2BO _�]G.6�ĠE�t��윮o�p�%�oAZ
��NF}5Mm )p�v�k��==>H�Y��\��P����{�2��
�RI,�3�UR����jL�s�fm�<�����1I�8��%)	�~V^%	��Պ7���:�'����?.�Nˋ����T���0�̇� �݈�a2�T���"4�Oh4/L��I��i��Z.W��(���{Z-� ��[�9�?!n.�r���5����͇E@@Z*Vz	�����jkQNDU�/�f��x���h��0��`��}��Ŧ��ko�Q��FP�^���)5��[���Sx������R�1C����<��Q 7n����3�?��Q��/��`�Fʨ�:���Wd�S��?W�����mm�>�ю�7�*�#K�X�a��������P��hC�{��}34��6��ֽ�7�  �.�̿���u����<K:ʜywb�L�x̻���pJ��~��\��*I�v	=��w�_
���zUe�VY6Z5/ ;H�N���G��V�d�Яf�9�1b@I����ez�s��k�끼bR���S�P�
\:���k���N���ڝS��3�ˡ9qd�E��:d�~��'���_D� p�ӓk�ym�Ƌ�:7OQ�����u�x���Ι�w'�	}�8	k���wm��Ќ�.wh��1�����ɑ��o}��ϗ�;�dį}�����gqpJ��wh�7��T��x=R'k�,��0���cr�r	|5W�Wt�X�z�{I�{���E�?fZ�Q|v++A<�DH�B����+kA6�|���t�f���{�i$ c�<r��a��؋�VT��!��lV���@��H1�8�����w>p�*!?.�h���S�'�|����,�n�h�.���|S���>>��=D+�课���!]�~\>P���D���ٙ�!��l�� 6Nt��Ⓔ�-oB��sި���U��&�H8	s��?jD�Am��!��#8ȕ�մ��o�џ��/t��O�֑�uO�Yz��6��6��{����6��� ���u� {�7=l�� ������ ��1|+��8�au��� �����}R4:�$b&-�j��3e0�y:Fq1w�V�b�!�wN�ze�XD�} n�z��V�3�X$��:�t�2��#)��/�v�J�6��� v�<X�i����G�-�ͪ(WICq��|��9|ol<^B�U|�ѭ�����VAxU�:)��A�𽇂�q�ף!��2�c�*]�����G�A#�H�W�������+�.z��i=64v�����a{�o��g}U7|g-hdq�:8�s�cs���Ϋ����{�L�8Pzܰ���"e���3���&��5Rd^~��=���P��G�S^FWѯ�����G(B�� m��-t��#�5B�ĺq`��pQ�8M|^�b��L�_��'���������+�����)��px�~ԝ���i�O����u��g���9K��&�,�\ ts5�Tg�.�Z���f�zOԴk)\ ��%DZʼ���*W�<!W�B�3G�+馥^��BǑ��L}. �� ܁G{6��W�Ҕk�.H�����q�տ����m�@Nw��LF:L�2�W"�t��q�2��Zŭ��DߊRP#�Y��I�Ui�.d�'��L�p
���'���������)$�8a��t����_����~;�?��}����_s�+���o٫F�_�����z|��p�O�������OL)�*MC�T�NJ}�s��{�T͒���Q%2��\΄�<��FD��7�Y�gw�����q�9ʠW¹;O��E�k��^(ҴC�$�7��q��U����\y�H����+�R;t,�͊������i��҇~�w�����9Xh3(;�ws�f;�U���VW�������?���� �⫃l9Gg��頪!bz����{
� ��2ۭ��!�a�k�6=����n���}��g@�&ɨ�\�M����������M��y��%� 4y��R���.#Mv�٢����QrcF�;~��٢���s��������7����(�|�eܧӳ�|�&%>��#�9u� ӳ6�4����9���p��\����Qrp������v��U;���ɋrr����Xpe)	f�c2Ո��ÞAT�zX5!E	��kr	l5� �D���Ȑ"D��2�Jɀ9�`�9�T��J�$�<c s���*]�� ��j�9�B�ز���
��-��H�^���H����'p��J�� r'h(����|.�n�v�CIc�Y��;��^�-rՆ���U�*An��Q������T�=}�*z�4�ػ]-�1e�A��ߠ�6l�FǱ�07%cV\3�eq�c�(p�˲\-+�������-�t������k�S��dU�|:��:�.]�������9ht�҃t3�sb�xbA�<$'�2r�d6O����(�P��������7�ǓK�0�} ����N*�s0��U��'�K� v����s��
�T�l8�\���|��&]�4ry��V�g@�n:ݓ�x��^�"�7i���#q������֚�Sk�G�pjy`�@�@Oma��OЯy�>�3"�co������|LmZq�U���%B�dxť���K������A3U<�LGJ*o�2.���D�I�j�wj�@ֳ&�j?6K�Nh}n�C�t��8qP6�~b P���e��� �b#���X��^<�Bq8 �K}�p}�Q�b}��}�Q>[迾�l��^6�%d�yp˱�����f\�����'p��,�E�9X��q~���Le��.!�M��jZ�Ap�CF_�T�)�I��ө��*�l��m�~���b9����"�����jI�Ow�,BzZ>$1+N��{�Z�� 2�׏���4�a�J��>���G�)�����$79������N7�o8�ђgɶ��d��o[���id"L$=�69E�Zs�	�YzM���9�1����'���|�)=6�*hK�sD�0��n���#p�%�[D�lw�>#��g6�A��h��|�H���=�+j����{�O�����e���tZr���9����oD� �û����-�K �Z&}NF|2ާS��!bg���*mȁQÎ�1W������o|���~�eEC�IC�x��4T���. ɖ�)B����6i��
Ŕ��(-f\1h"����GNixy޳�~����i��4u��C
>� @��[�����:���o%kϕ0����V�e��ڣ�H٣FU��WY�~�H������u[."w5Z�ͪ���l��҇�oB���S{%��<�!���h��?���R�*<����%���x�=3���r�t82���/�3H4Ӡ�.X���G8|�P'R/
vpX��<F������%�t�5��k�1a�E&�|�}�6����<J~Pż�"��;6��@����n��s���x�k[���.�?����Po�"�`��|.��� o�젂n�)�:#�I��9<ы3�>o8�w�Q;�3ƨ��N
T�Z���+VEI�����;,I"�'Mr��M� ���\�3��N�����r� O��8z^	~N��x�*��,�g���������=</�Q���v��Dg��%��V���T���V����5b�LԂ���?��TuӃ@��_y�q���:�J"���O*�t�cGp������v�G��\q������.3d�^��/�#z�?�Q��C ް��:E1�]d��38�$��?����R� �h.k{��D�8��!� S[�׉ZAk�d"R��SMk&`^�����5�/��Q����	X<4�����x*C]������t; P�.dq�~�nV��#�������%mR� <��D༣��33��E��:l2��DW.���qy���9uc�mx��0�/on�6�J�Qa��;�3A����k���H�vG�����ځLR�75��:+�L;����u[y����w`�Û&��k��Ï���Җ ���i�=���� �c����yz���r�%ی��$���t�zC$���`8��E@�y]��;����ȇq�l9m�Q ��:�����L�p2����Ü�����a[���O ���Ĥ�J�,�^�nI���JDWkM��y�J�rF9:G�>�QiiS��+���ņ^z������N;;�f�t���#d/�ȝ�Q:gU��-E�۟����9�����H�X�~�3_N��������^I��X���3��1&�g���|c ��Y�Q����;I�`N	���!^c�S��+���p���3~�a��wXz���r:�b���1�~F����?�Q�n0�7�I��������s�'�ѱ���k�W6�zE�[ʥ�0�8FÑ;pV��r��zU3 ���(Cq�R� ��׋nϼ��mU�`�H��΋^ �믞��O+u�J��M��ʆ�|���
� ��r�����A��=G�K���󊉞��0��pZ��t�+t�0`��]��|��jetT���?��w^q���2g�a+`�V����q,�`�8�<���=��t����f�do܍R�ƌ����2�N%��Ks�ݰ��ră�^��F�5x�<���#%��>�ؓQ]@��8����m��t��r젽f54�N�+�)V�>}f`�ۉ��FZ( r8��o�������2�j�J��'��i�!Q)�DK�-�=<?0�4t�HjT�!�<�� ��J�lj���&49����9È9��<x�����?л�����_߾yˤ˟>~�ۻ[zH�/�»"f�vZ�W�*w�,3�%2o���h|����N�u<�y=����R����7��'.��^����T�wk5���`3Kƌ�Ɉ�&y{O�w�IL���+~.e�n��@T���fwJ^����2���?J����<if��q��`dm��t˓���˚II멖w����H�!�6F�$;C�K ̰�PnP/_����������E���yܱ0����X	v�S+��jm��=Doa�W��4W�Js���Z"y&�k����@";��A��N�@�(�� ;� r��K�5���}ə����(g�Aԑ �I�c�@+�)�LV^�`���$��R�sP��nS���/l������bӇm����D,I^l�Y�wK��j�������B�*X�Ҙ�]�B=|�XXu��1O�T� ����zy/�o E������F(+���!]��͋V9�#JpGʓ-�/K����n2G������1�E�ۼ5Y=�F��0�Q��� X,�����o��1@ɮq0o���H!~[�Q���\Oe�U=�4�Rc*�k�w!>��;���K�?^3;B�-1��_����h��~��7tΙ\��o���nA�`�ʉZM���Z��p�j1E:���
er;G0d�46>��`�����4@�9[��(��@w=��E��3'Xj��v�i�i;�����:�&)��O���M�	�9�٧�/��d�W7��5j����줂�6�]��tZ,MٞFJ�ޚ�T�.����v�Q�E�*8���/����F6�B��0w,��,�Ys�s���fH�W;>NŇ�#����$���,EXl�ά��� #_���>�d|��v����l�@��0G��ʥ�TCIy�2/"�C��ܹ.Rwxѡj�Rו�G��?s��ʎ���_}��O(�X^�dʸ���P��5��sp�a�U����.�������ᫎ���6�;:�Ŋ��.#��~5�Tl�'��WɆ�H�Ֆ��O�8Z�6����T�U����hȢ������+>����-A�?�5�h8�	go�.�.��z���fIm�ge���[ium�ψ|`̆����kɤ��rԉC�M^���Ҋ(�O�?r�v���oV�Y8����5�����晖�Ot��H��z|�h%���Q�*W�m�y__SZ�eu���_��^~���N6�!zz���?��Q6T �bيô&|l.��m���°>�N���K�YqN[��&����r�Q.F�
wf��n��Qiŀ���Ї�1d�l9,,� `ܖ	���* K������b�N�JҤ��@n�e��U��,�g��m��`BH�}��M՗���ò��hS�;{�-\M9����I%� ��kd���Sp��^tqq��f�y�P�$݊���l�2�,��\I8'Gpɏ����ʃ��p�(eM�G	�1�8􏄰���Δ�v�jU��KX� wD���R]}��7(�B�4��S��d��A'C?�)B� �)4�B}�@p�cq\�7~1Ju:'���c�6�U�R��gp^��:�!�\����󤑡�?G��k�2`��7m�=ӵ0/ cWJRkza����T�#���D$��y�>V������G&������ʅu�Տi����9:�yN�M3?��cccs?t���%�54k�#�苺�2c�UC�8�d��B���ck��w�[]?�ݯk�~�ol����L��T�����v����7nyʜ��Gb|w=[���QU�sr�G�,v�W�}KA����Z��CzG��-[�%O7c�����������g�
��L<<m���#q��$�S��m\g�tL ������gbep"�z&�]�&���T�VS�3wN��L>ǆ{(��t-*�k[4t�j����qD� �A4��-��N���G��j����<Y�q���h�E��*(�u��(�,�֍>��7`&��rN���[vK�������K��1�-�|~t�/;��_�D�e�䉯�r̢�qg�>8�jc}���맗�����`�}���:uJ�R��/�.��-V�����%�<���>Fe�h7���t-{\.�p���~t�T胟2��l�.٫l��96�y��f�]?�'���h���O��:�b���L��� A��5���f� ��J�OW�W� ��bkU|��77��ٮi���s��z������d�HQ'�&��>&��I($��)�tB	��ڕf	�>��7�U0���$�+D��l�#<0�0���'d��㈝��ڹyC?�}Ϡ<hg����/?��>�B��[�����I�� �TX�6U�����5n6Ĵ��	fsA�.��<��'�7���^JS�S�Q9��aN������G.6a�,����)�=���be�`L#�S/���]��*G�<#�$J�u�L^ D;&=��T y/�@b��`<<=	R2���B_�r��v��i��'�mjÜ�4J�`���TX��AaX��fF0E�T])���+�߷��Xav�mzͶd��)=���U�˛n��t�#Yd�օ���D�0�:-��WWk'��i����)E[�\�ҥx�C�iI��F7�(�N�����%�ԘRݶ�X麶�'���.ɿ�+��nW�GG���'�ٺ�د#�)����7o��_	�dojV��=��9�D��9⇰4�T�����ٽ�H�H����bF�0�T6��9��tt}��\wݗ�Y�sp�Y��6�������e>���{3���.�^}����~�3E �>Y�
l@,c�ϰ��v��MS����o:�7Ģ����qd,~�����{���/�B�f	&�����W2@ �cI4��c�}�@L��0�sc؜z������9�`����xDh���jቓ��.tey�S
{����Ń4'0\�v %y#�P!����@�'*5�̘4��0<z:�:Z8�J�n,�X\���q�O�o��J]���w����F%����M����)�Fĉ��'�������X�U�Y
������^y��@�H���u2�B��@GWU�{{Ď�]<tB/W/������3�;��P(��~��1�g/R:���o��V������_.;	�<h�C~�!�j8�GN�#�b��9���{�v�P�3���t� �R�loT�ނ�
���	s�.���>���M��� sA�>2 = M��۷o�݇������@4�8"(@3*����� (������y�����v�Q4��*]�Y��6���E�k	�����h��۰�<�ޥ���]Ra�Ebj���&�f�J�咣� Z��e������|A���|v&ՙ�w*������Rc��pðWc����P��QF�Ҹ��7�x�c��4,g�O�"�����o��ԶB��!� v4b�C�H��8?�p�P�ׇ#�Gfp�A�;+%>B�����!:�9K%5J��������	�Eu2�'I�O� x�=� ����anU���K��՘8�!��%����F�"��y{���҂׊ť���2�PE�î�vQӥ�GR�txtG�G"9j���dU�J��QO�F�x���w�c��#J�XUKd��J�4�/�l�Z�J�QhJ!�?"�}�;�*��^���kܾ:ݯ�b���P�2�z�p�z�(������)#t��'K��Z	�<'<��#�ڽ�Z��#�b�w��<J�A�Bb��ﻥ�R(e�"����f��`d�N�j��?O&�r��\�sa��zf8�������.6C�D��c	E�������j<��=�A��{�79�J����o=�H�E,����W�ʰ)������H��vL�ʺ����|���`��G��k�@l_���(Y��~S��C�{b"�؊�|�D�Rx��q"U��ZI�%�F�
)
�3vN�?��B0V�z�##:�'�.z�ɶG�Ӯ�s�ZqN���sUK���~�=Q]�3�#�:]���afI�/&Q̝�"�~9r��>��9����H�u�r�A	��뺣����\yQ�Q����Cu�ʢ��K�t$9_R6��@�7���O�{{�+{���V-w]wl��6��_��^��k{lN����CEw|	��M7��x�;b^g/�7 pG"U���-\}z���u�i��77���W���3M�3��sz��s����7}�����o�Ï?л�o9����Iʦϥ�t�RkuA I v~��w�x��yu@�`g�$�Q��r,��ES��>����^���X	����5�����BdI����>�ׇ��đ����-�{�3𴡈"<'Sv��6�N�g��;/R�Ĕ��'_��f9�f0�u���<���>�}u��NR|'	T�)ՁK��X	���<�@Q0�(�-JB6Uc��y�]��($���:^7N��)�&a�9l�0��D�LfS.I� p��s�Z �j�D5��NJ]���N��.�H{9'�3u#��AT�n8گ�(����lј���k��F����.��|���dƞ��D�XT�U,��d���ZU4ԑ�;
��]G0��X��AS���i�Ǯ�CGٳ��U�}��<�i���ܬ>`���,Y*��Kmh0��`�2��A���@x�g��F^H�]��� D�c��_�f�!!���HrE���e�ll~v���K�O"�L1�.�,_�Ý��P�KT���%�펞B�2��4TzF'�
��2yM\���CE��ӻ���Π ���AS�Q�?^���,�������E6G2��e�c���2GZ=�yK�7W��8��Ԧ�qdͿԜ�ˆ��Y��3|�_��W�+C}V�T�6	�
��Գ���6�m��׼!/>��ET맷V�:xL�0]O��b.�<����rw)�.���'�:z&y����(n��&F%ul{�8f��~�m��[�w�����2}Od�u��h4��r�����D�L4�HF�,��]�#)G`��@ؔ�����\�R�s�u���U�<��k����fg�|���a$Z,�M_7*����w�~y���s��"��7ʜP���F�'��b��. ߵ4���XeGW�|GF�̩�
�I�VK}p�t�U<��%�s)?�=��ѱ���b�����߱a9���TY������r_�R��w-0S�'�#�;��x�B_m�}b�����_|p�i�3�M��n�<Zo9��+L,??cP`W�J��&D����ϟo�`�����l�b���W�0N���;.r�M�s�B2T��L$	���6(�nG=U�nH�=2��̛��V����t��x�R"��G�Ѵ�[<o����'�{|^���K��H_{N�O�#�$�� [ъF�d��:��\;2�rM��P@����<X�g���-�n�b$q�����l�`�������He���H�	�Tkqv���U:��H�B���b8���yA�:��e
{7^c���}&XJ��ł&��T��&	n��UjK	C^mP^������?3Y��53�|���W;J�.��=�.1|�������`�/eT/]���vP��
pGu>D�I�� :�R�Ĝ'D�U��貅�b�VdUS�4'��صj���2�C�5e�ց��kGB���43PǑV��
8?���VL� J)`Nm�\3j�3�S-c��%؉2|��P�/�
)�R(\}���*K��?f1�k�q޸�tq�WuIˍ�\�`��:~���ԋ����#���p�N�Q��k۠�=��I~;7E؛M�^S�$��~B����7�����qt=4��+fs�<R�KR�L.��!�GF�w��c���m	�g�Eu�
���(��:?�f �Ƹ|.��Nӡ���=x�xp�/�����fD�Ǐ��=����-/1����ޝj���A6�D�px���<�>3�`N
Xi��r�2�U�Xw��T���pb��07޾��(�8���R?��$�؊���5y�"��À����c;Ti�82DJ��w���,�s�^� G�����:/
4b����_���3;ZL��j�N�$�꡵�k��$O/����pQ�V1=#j*�#�`A0�&~��GV$Eg(n�啦(��gPCڝ�A��8F���ٴ��y-Wn8��z�f�>��������^�G���r��zUٗ������AW��ߞ����#롯���UA� g'�̝/��C��͘���"(ޥb�~��DfTa_��@��m���PY�k ����5m�7���9f2�8i|� �Y:o:���HK���\��ȻN(7�������@�i��9���ȇ���|��:��Av������;�C�N�X�mH�]g�.I���?���42��V�F�U�T;�p��S]����Ě�38�(}�+�7;�{����3���g&�F����:�����sT
�㽒=P\�G#A��m �����U6���Hx�:l�;��Vc�C:!�Z����x6_���I�t��t���R a�-G6����
%H�w���F'�n�P�M@/�i���\5�|z$�i5�G�̰�4.��dL���;h��f)�4J��dl�=o B�,�^�Z!�u�������P�
\cv��T<�7Y�/����X"�۽���l�^JiW�|��� -�R���kR���)�J#0��f"S=?��N�UIc�8���̆�ܔ�Y'�x����M9���[�V��{����r�׹��~O	������4��C��*���1W���r�uT�#��[�7�"of���F�reVtl���3����d� �Bx��oo/�*��xkȶy��B��m�'��V,A��JV�!��)�9B�=��t���ĕ��E�����8swdE�`���s���yZ`�pzr�n\N�2bʸ2�pk�^Ɗu�GU4n,�}1���r�}S���_C��_�?�ҫ=rS��U	��j�c7;Fw������瘱u�Q�AQ�%�'C9<�&��g�, �6�W�+w ��*sޕQ�M+��cx����q�7�QҕZ`�y��&�4���d�wx��������@6~����? ��*�)��N�+1'�F|� ���R�Z��� :�]��_�3A#b�r�I�о7�F���=`�7|��0�DY;tN�ы67��!�rEJ'u(ޗ"F�
y�h*�59T�n�׳��KC:w�}1�x12�_����I���@)�
�jZE���3���5ӧC���1�s9ǆ�G6'\K���Ӣ:Fzs¯3X�6�]�Тo�5��8���]�q�l�RF�~�������u��?Ҕ�&3�x�5_ЛG�\���K ���;_�����}��4�����^�aRy#B����Ӌe�^�88����#��M6�9�ի�+����ղ��gs������f��M�e��O8�e��h�[�z�Lw���^ɾ��M�;Hn���Z��+خ�z�4L�U�tRs���$f�8��i�i�J�6
7�&=wmN�:0��j� �M�z�\@����:d�Q�h���N�e3��\ު7��
���}���p�t�s\�@��h�d�t�Yj�s���e�ߑք�w�E�򥢒=�mvPD!t[��̈�v.ϑ�6g�	��a�ьł�?j���� <=>���OW��\[^���pNy����$���R�n�U��vʀ�t�0����$��Z�&[>L��y�
�=�b�Az��J�T1oAͥ �yR�,]Ɓ\����V²�iܤV|��%5�H5p�ICe�6�Cf��>	8��z�l���Nw ��Y�6� O�D) a,��ļ�6�!X�`�LFPU*�#����m<ў!?_���#� o�7�n(�9y����ȐYn4�蒦M:��7��0d�Oގ�ӭ�~7���j�k��{!�ߨj�1���G�)[F�cS1�D�8x�K�3�u|1��6ws�[�~�zJ����F訌��5�c����h6�Qm=�B�o�͠�oqx�u��\�tu4���#���@����R��- ]�k�{�G�xau�!a`Sԡ�˝��{����������|�#�"G�Vp@e�����C��cS��忸�E����OԢ����gE�����_���K�yWQ+ݘ�S����}+��Q��[]������kU�D�����2@`��$��ϣWNQ �C��io�鹡+@����j�|����E
*u�hĈ�ƺ絯�5�{�V��I�瑽�J�����e�}f�Z�d���W�m϶g�΢Ju�Աr�A��`\U�4�<Ƣ�5~n/�+��4[1�i%0�8B��c��t�[�-,���ʮ���5���"���e۬�rS��ЃB��E+���9�� �,.\��v͹�K0��� ���8����r]bЕc�.0�r:x�טx#�������$�ǁ�#�| kL0�$�ܼ����?g�9�M�4k��^�8u>{������+�Y�����-��H���W�U���w�-�u��\���ryq���I�ߣ�L�-3
����>~���w�>S���)'+G��j߳�8����^� s8b���E6���&��]�-��U�����1ĲW`�@�IaRi�=8j��3K?�O��3l���{ht�ml�LЫ��Q�U]��汯��/���}\��l��z�f����bBd���1V.[�P��p�X��.��6�qvvv��[��s�$qçvy��} 0G�fU�U.�H����#t*=�Q��S�N�<4�i7{�,�V6�ǟ4ɨ�&���UD���Bg���eC�us�9V�n�ڹfԖB4�Z��Y�ȁB!7O�����)����e},�'r���Ez�{Vj$�3TU~��Э0�����zX�ѣyD��ZAm��Y��W�WhXo�
J/e�����	��V�U����#�$�C6>�����)���!�K��jQ�w��j�.w���;6oJ���.�E�CXg5��eDU.7�}h���/����Ɣ?UXai�b8A@��sg�a}��$ �tUl8�
��w�٩<�r?0��I���B�9������zB�V�J	ڄ��ʩ
�m}��4�n
���-�I4P�ee�$g�(�Y(@b�'<GFTyv8�ɑ#~�)6nyl�*�Ak�I����$�ScgD�����ȱ�@S�;{^OH3��	�'�1!^G�j�k��Iܳ� X�d��L��'O��.(�ĨX�z�o���Q>�ĐI:��sdQv�RW�2-�� r���J�g䆪���P�m�s�O�����G��|��u�WX ��Oǿ�3kIB�����e��c�f1�E��yqp����T�MHW��i��5Y����̿"Vz��@��cU���rW���ͲkػnH(�������#c246��Ғc��\R� f�Ջ��C�=�	}�]��!�}�m�Q}�r]��;zB�n�z���;���.��
���#$ծ20as2��vk��r��S�G&���:����-�;v��LZf��%�G�+Ǉ�/�`�ޚu�Χ��7��/����ԙ,`�:тx��7p�~�2]�@�>�Յ����#��q�y��"��Ws^{�{#�dU�*�����1��,R�sǝ��F������z�DQ)j�n��(z�t>��*^
��{.�����9�$)ŸnV�Z>f,3��4����������b�9'_��a��ю����s�N8�dq~�9o޾�w�߱�N̜}+;��ۓ�*��gtq���gN�F(Y����S���(�|Q�����0�'I_��{Γ���ޯyM,��4m&�KU�.�I�)�-��M����)<a������A��"�G��9��3�FSOX�A�l6W��<���S��v�N�-;�S{V�g�hڣ�{�u[�o�L��{�-�Qk�Om�CA,OTNҏ$z��O��r#�*>|^+h�.u4|�8���.��tsu��Qq�9uT�l����t�F���I�FT� Uֵ� ;�G:Xn�Ǽ�d�������:Q{���;M2�͔� �ꙄD��������g?�A �gOr���1��Ya��X�,l)�ola*V��̀�%��!��虢���ϼ#�[ƝL9� @�J�|9��.oh�v)	`'!kB������5Q�ӂ��
�=Bg>�W�W��Jz=���CI:���d�S�:=/�^Ev��{�+U������<��!�l�29�;q ��fEm,"gz�^(�j#�y�V�G��-R��.ݯ�"D\y��yu%����,�?�L` ��^a�)�6�(�Y��mh��{Ie;�?3-i
��ۄ��)d�+jv�BI8&�;�ni����oh�I��س�Q��k[c���|��d"\?j�B�Jn;�@ڮic�r߸��*e4�T�2�����]��6 ��?c�~�������H}�l��f�zsYV^/����t�P���Z����XK����<�����r�EU�1�ZƮ�\���ls��-%����s;+�*��R�d�2�_�4<GS5�����|Yd^Gf䧽H�'S��]��M�Y\��|�V�<�y��%��_��h���ON�4�ӶdN_�ȃ՜���{�+S)���������糏�=���(kP�Ru׃Q�i�{v��lѷjCt���f��y0*�qڑ�&��S���i��[�Tm��o1 O|ף��_�}�����!oޅ3�e�t�e��T�V�1_2���E)0��~���#�.b_S���+�/u�S�~�Ե���p���f��=���!I�P=�������NA#�Mw,n] ��8��m���{�۱�;���O���Q��Օ =��z�$m�#�����5W�c���}"�W�t1��SE�����I#�+ӇM�#{��(��֊#��]^x�h��T��s�1c�eb1�y���k��/�H���6�ȴQ1�����Z����.^��K�p3����_4"��̲�E�#_[cm�ϩ'�������r��(�U�Q/��A�
����/�6txu�RP�B���ƝT�S.Ц@f���9�  Aл�YC��i��q�j$A=���s{�U���ӆ	�[1C�>��S[��@��_��+f#E���_�����ATPZ��U��vK9�2�y1I�~�QD�]-���
��]�Cܥ��3���3���=/���=��6���f��Ύ�v��ݔ�ft��	��g�4� JL�����aRQ���Պ�SC1q��"�
��d!�3���w{2i��bQ�k�4	��ܼ�w��@���9�t�	�(ʧO�Z��N�� d�#�q��aB�ˋ+�&J����=>>���
�<�M�ė�|l�)�l�Jj��R�nmw�h,deW_���g��B<y�j��<��Rb����ľ�)ƺ�j��)DM�����K��ۦچ��Ć�0?�V�0_�hy#W�B�iv���ݔ7���i�WU5�[����CSt����r�5J0E����ف��se�o�F7�w��!�:<����I�����2z�ؿ�`�h��0y{ms�q�kiE��)'�� ���%���Ȟ����"m��Ç7i�a<�̵#=Ţ!#�P�������X�Bz��O��N�c#���[�*��<�`n���\>q����e�=��� �,mf��<��b�������%Y�6(��~V�M���e�v���.�9�����(u��a�ױ}"�w����b�g����x��L\�=d�����A1H�c")���%�i�y��Ұ�N9�J.��2QEc]Qy���7P�S���NדE��]~��Q��$�DT����T��P�c�j�t�#͏�$y�}�;k��12O�}�����G|�{_y�J��|���ɬ_�J;�Js�-U8�m1�}�A~���^)�1���Տ$�k�_c���F��[�mf@�]�����1�������`s8�����_;/�O���#�{Qu��X^�gz��R�5#ǘ�=���, N�֪	�b�N�	[f
G�\��7u�e�I��UwJ�5U_�,s!��	�6
�o�@����ߐ?2YI�͙�:{���0N�M�T�͊H��8b5�S������P b�����`m@b�߰�|���j1l�e3K�8���nsK�}>����$V�̕a�YH���#f׍���dV�-�<f�3���H���o�m�m��?��n.���_��S.��m�����}�EfgR��?��ur�e���l1g�կ|I���l!��I�g~�<O�O��eC�v�Dī]zo����;�t��>�~�R�8؉j8�{�~�`�l9����3��w�9�}����zKq�)�<a0ρ����Ï�V��޾E�O.L� ���Fq�6J�̣GJj�*=�Y�yi��L����O��D�z�hy4>�F��&Q��F���f+<����@�4��Ւ@�%��Wk+�he�d�Q1�O������1VkA��+�c�����!t~�zjY���<5=M�Ֆ��T,��^]^�ۛ7���-����i:���ӳ�+�Y����Oҽk��_?�n{G˰�(ʨ�6L�D��J���(���W�
��m��D1���v����f� 6�ap~~OrE�ȥ������#�a*zX�O&.l�3�Ӟ�-��2�U���S�a&rE�ɱge�0�jxs۴:%O�Wʟr�!�7��`U�%���Z5ZiA�xys�Ab'(z"��⯣R8}���̩c�]�Q�3Oǅ�Z����p�1Y����V�"��Q�c�4��cY�����|O���?��Y���9��u�ŬD���e����~����р���?�d�0H��v��V�VW�ػ��m	-�l�|��M��wwt�@�В�v{�./����w����
�E o�I^Uyj9|�M�
e����1�w�d�^zJ��+�{��E|�2��+�+>�ZT�6���Q�9T�.b�$��� ;]V�q%�Riѯ��v�v0��Ք:�Vb b}�˥���-���( "�����#���(2O�R�\���I
�[�l����o=_�x�&,�:Zoօ��V��
E�����%�Q, �Qv��=��n�?�Na�řSf�wf�!���2�*���r�H��|��E�Jq54�~ǹ6�Z�����w�7b��U��L����o�� ?���wm�+���c�9����<u-��=����BA�hC�b/�A�=�rl�>�"�9�pX�F�t�)�'����=>�9�x/\NƵ���J��l��rH�ї����/j�DsWW�D��P�BA��4���O��B"�ᬪ-JTK�+9�v��hV�p�o`_���k�NuuK���Ca���>'����}Ł�b]G���(��Qu�/O�--�>�[DG#}�-�GmHO�+�uGv�(���<hŹ�P���u"Q���\����'NK�6Ӥ��H����/�߿0�
gɤ��Y��/��₣d�����]@�g\��I��i��R��� Ҽnnnh�f����h��]Q9?��������h�^2y�6C�ѡ�5�F�X7���iW�����m�-?�$��iM��~C��tyvAO��D.�S�,�p�,�K�X�9��ß�/����?	q�E�[`A��3,�m�{�����Mmۦ~|��ݥg���WN's`���j���-�;��&��(����G�SO*�!ȋ7O��Rd��*@&ڔ�6-�-e&�>��h�ԙ(��G5r)4a� dͶm�T��E� e����s1���Dgi`�M���ɐK�yt��q=��C���(�\�BS�0@�L��2b�f��V.ʜBP�Y�Y�����k^�Y��a�%����K	G�_��J���p
⡬Ө�N�c;�+�G�K�WS��~��V))�]G�$ؓ��[[�Kۈ��ny�;	���S������+Ai����$^
G�'�n �f�Ю?�5�b����㦊��}���ȩh�s�*¯�b�s���
�B���Ε*甲G�_�L�F��W�m�N燔?��kbvBt�H�iRk&v�2�^=�ZX�e
He|������>��p��p"bh2AZ`�
K��Bb�e+Z�h��]���#vj��!�ٛen |�OV�V�k�@O]�=^�&��ѯ�ǯ3���Qr��8�8����� �C�����CiwòA*br0�?�K�bY���,���D�U�{�߲ ��x��c��EW5�/E��M��g�n<�g�ȵ��%�dWIʍ9�2�g�X�K�{�S�2����_��N��-��o��8������S|W
�Y�#'����{t�ߗ����NW�]D�XTg���`���G��{W4���B�=�K���v !zՄ8z���>��S6l����XYG�6��W�����5s��|*��K���`��3��'�#�e��{�c˓�_�}{�=K�N �V�#�?bh���Ǳ�[���%�� V:�K���g����[�(h��R��`v����e�t��#L
4,���=��W��)	;kř1 ���=��l��Ƌ���8���F������v�����c�y�~Пۖ����`u�/�,�M���D�*�X�Y2B�\�:�����%m���,)8z��>n�����ˍ��I
z+zrHLsd�����T���kN5�xsé� iV�5����J��l�e>f2�c~R�+�,�6���Oi/���9]�������7t�l��dBW�nhvyF��?-�����ǖ�6O ��հ�El�m��K�py��h1Kי�h"�]�{*��w��	�/�L�|q�A+��gz~|�j^�BD���F�͖�P�i��/&����6�=.��sv�`�t��$��U����X�n�n����e�BM��v@�4m��ɬ���}���n�>����Z9	5&9�00��SM�R�:N��)or4���7\�x�9�x5����V��m�LX֒2%joe��.���D���c�� IQ�7P�}��J@XƬ��L͊�Du��v/�I���l�
��s��8ؔO��%k�|#�ڏ�0��P��G�9˵����8"3r�R	t���!cW/��N+�����j������s.�VA��	p��NԿKO~��k��y�*+�cj���j�7��X '���S���)E_	�xU�9Ԙ�$F#
;)ϐHV�@-U�`��5��-Y%:%��5^3oF��W>7#9zη����s����oBo@�$%d����6����K��1Ҷ:�rYۍ�N2�=�yZ�S)��.0���Ճ�݃y�gl`�yB˧47b�� �c��Z�u%��IN��HBMu�np3̬߳�>4ȊN=z|�L9u�:@�G wX�ԪX�s�{��8Ԗ��k�p@�^d��D��ƏTN�l#����L�����ו�v/�n	
!Jl�|sZ��xU���595KxQ�_�؟��A ;�0�[C�!�Q��pz������P��o��g�hVVW�N~�Pė�7�;ɖ�,�Pwo��u��� �5(�'pYV�ԓ�N�{���K��^>/"Y�NΉ��Kzq?8�/��9q�x��tx��P$
���ڈ>v�)�l�g��IQo��Q�m~��;z�c����s�ڧ�͗�HY�������=J��Ҝ��-��F�UT�d��*g�G��>�{��Y%�e]3��b��ic�9B[������T�i�ɺ���Jrl���"�g��W�6�����kځ�#]c���bFW�tqq�e�a O�&C������g�����b�t`�Jm�<Ԧ��G����(��(u�"T���#$WO�͘���E�R��Q��H��Y���5,�PNG��ߌB���A�eN ���;痗�<ͩ󛫤'�(>�����*��t��~K;�����瞦�F�2Z������_8UiZWWW�ޮi�����;N{��uZ'�7�4I�z�t����/Ҟ� 9��b�DY��uD6O�lz��(a,���S74t����Wiͤ�2� �O�.3��ؤDA'<���[zx|�1��z��xu*�9^���~sC��7�go v�5d���O�AĎ�Uh��۳�v��0����ǚC�?�~���ϴٮx�����Yd�5'�ft1��[�h�B�	�B.���pW�(T6.�[�\�+�2�IQ+H�0�kMLZ-ܭ���n�nY�aC��zcm�~��}�I��Ҁ=3)4of��*[�!�ډ���T�e<*�I_$�J%+����>�����"3á���pv�1B��b�3�p@dէ����{Ze�|ԕ�X�[4c%��\�|�Ȁ���x���[R�@�U�ب�\JV7CV��^Ct�SH7���Ī"�F�W*!q.�S�Q�GI�����u�be��;��>[?�{
���T2���Ke��u�,�����3{�0�U�K��@l��G;p ��iW�VIWs�c�x�ڮͤ�Xw�(ߒ�E��!"�nH���;�W1ƥti��l���Ӵ�:�i���	��қ�KV�H	x�Z\�/�K=a�h�;sF�Efiu��Q�\{�Y���,`��la,���yة8��� '<d3��h~�[m�S��:�l�#���̰h�30��F��yn�Q@DH8��O]��L �V��) ��(<"���A2�HM��Ӕ+��Z˳��g��-艹&�΅h�y�t����lL�����n�z�6��.J$�C���i��)�j�w�~˼�}%��eͩ��c�X�{��v��Q�$p��,%X����[�P���T���F�P*�6���!&{D��]����M:�ȏjD�_��=�Dwڲ�.�^hS��(X1v�~q�N�h�#��~3�N1V�T;���w��A;F8Kʶ��Q�C��H�B�����pZ���F`���鰓��|��e=)(����r�x��Q�H)�R+�@޳��+�����b=��b���Jt�bQ"�@܌+N�γ���� ;��Wթ�{�����d祟ͬ����pc���؛:�[�L�S`���_%��йh�	4�!1�J���ka��d
e�& �}�E�UB�|�ތ��=3��7�X�j�ꌂ]=�<�W\L��x���f�^���9K�|G�|���I/{x|��?�����P�#wj����7������&�i�Y�r�L�vCmZW���CO�ZK�d����gi����'����8�]K��V�-�I�w)Y m�9��yô��T.���r'�� }f�� �@��� ~^����
н���pT\C�Z�����5/ >�~|xz`a ������6k�G�1�sDƕ�9�I�U/�-�2_�������4H���6F&�!�-����@)�
J��'�S!i�F$�2��*-�<lg�h�F��DS"�`�t����$ @�H��rE�>}��~����#���z�KB�Kj&���z|��f�O���#ڨ&3h;�|v}��C���X���i�G8�����߁���M��hV�b�*�@�k�/&��1ᡛVg�J�?bXkL��#�7Q��j�Y�E�T��#����3��e�YR,�9z*�kk�({�+)�(�,s�pi�"�+�<���E��@{5R�VrޚT����t�N�,��0-S�,e?���2�s�	�8<̶ؤpb�*��9~��ܛ�R������VI��5�Xp���a�W���@���3R^P!��yOk������ˎf��N���2(^3�g,p�OH)E�y���]`�r�o����-i�z]G6��z���Y+iZ���2�=x��dO�,d��AZ�Ct՘D��*�F��U�<~�)G�R
���M䜲�=j&蚕^l:�����[$*�W����Y(+e�;%�+ykk���I�~��p��ۮ�s�D�'��ryu�$~1v��u���a�s��T"r�w�ڪ�;��;�>�B�D�2�z�$��R��H�wsZ�ǥ�13�ʳ^��_����G��~MЯ{�;���O�RcO<��Q<V�ԕ�he����<�+��C�Ϩn�F�(fA����SY̩ﳮ(� �\
��.�=�����\���U�C����������޾�{��#G`�B��r-�=ő�7��zW9�rN��#{������o>�	חHN�a�6?-%��_��˱~eM�>k�<_Mם�W (�c�M�BV�t�}����� xB%�����9��9KZ��a�Ԛ3:u��#��y	,��v�5BR�Wˆ�Õy���{
.�f>�$�f��d'H+����<�;����d��٦����i�*+�az�@�����jy\Ʀ�`����m�yqi�NQ���T��:�ꢼ���)g�ۦ����Rp#�:$�q���|�l)z�h��7�S4�:n�w�6Adq3�3�-��2Ϗ\�-��AR�g�����L|���`��;�N2!)^�V�5���.�T�j�dvD�"B��	M�3��u� ��^�چ����T�ŏ�G:K�qsuM����/�]p���Q��U��%�[�U��+z||��%�&#�f8��9J	�~N������=;p\����9�Ȏ����+p:��[y���TL*�G2�6]w�θ~�Sj�v�L;�JT��e�SRa�i����"V��W�i�'�"���Zj�riQ;_ �rrGɷ�)��V�,�� j��D�͞#>}�L���-�U\�q���:M\�<F�y!���fT�9D����(���Jig�W��=���*�8�MH �N�E�)�0ki9K=�h(��i�O��R��Ϋ1���=�nU*�(Vl cSFhk�9�{��  �R�BLY���A�1xx�TO
G~q�h���m�cZA�Ƌ��:��'3pL����͊�D���.{�y>k%93��sn½S�R����u��M��5dV�u���l���2A��t,��n��#�#��\}̼����F�{UWI�0��Z�J����cޡP��(O�]DY<���)�Ѻ����ԚGSb�Po���1��A�=zªȐ���:�4�u�Q�^K�*b�Saџp�M�~f,�A���;�r
)3���H���4�Y9Ţ�L�R��g��FB[U!�9���	�X�-鳕��L�����RN�,��g����hۍ���+?˷jG&��^���<��]v��e ��U�x�%��3�Pg���	!L6��E� �IZK%��F�F-�ZI�bb�I&S7e*�$e�+�E�
�:�>I�����}��pE�4�����8�X�u����f��r���p!^�x�!o� �x�� ��NP"�Fˬ��9�������B��f	&p�Gb�L��ZU̬D�,�Q海��I�r�ӱ��G��O�Gx�3ϓW�&�7��G��_�8�k���I����Nǎy��UDp1�/��qYa��N�W-ͽtҘ��AOe���'�F��#�\c����%j�|�h�RV�A�h���e~�V2g�VxJx�|"ǭ����(Z�������Dו�(�>�_��~�Vm����qgJ�}���?�S�c�l�yѵ��^��Z�}�e��Ѽ�j�Bs	p�EE���>׼�r-N��g�}x T��r�kȰv1�J�H1Ȣ?p䱔էQ�>��6�#�s��8��s��^���xL�ߩN��S!���B�O�����me�~�7s}n9��ʯ�SS�
��X�<�s3HE�p��q�\����^8	�X5�v���Ez]�GF%���!-Į������V�P ��ʹO��b��4�$�g�ӧ��*�}���O=P��Φ��1�z98/и���HR�"t��c7{�����cic��低|	�����:��y8���]ܯU�����m�o�-Rꂵ��v�c�b��"��&���q]��O��ן����:F�~��g�|wK�Պ��T��T�ڨ����gZ|N���^T�B�s� �~�m���\]_r��4�ҵ?}�DOK��Y�l�i��{~��Zֻp].촗BH���?=-������5���ޯw���S���h�޵�{U̇su~�:л7�D�����6�Nt���|�����}�����6۵�	��>N��5�[������򵜅����Z,�U���<��Ph��-s�l}CĎ>P*�<� �|�1�Ft%�2�1hU#�@ ���pC#$eҨ��H�]���#u
���4p���2ɟ?���`�@��-�>;�h��e��u&�c��i��=�-��!z[���fx���-I53����[S2*�A1=�6^��]:����&**S����LTc_ƈ�BU�\�����u��}��J��F�k1��jc!x�L�'��
���YQ��Is���<��~���)y�rWH��5`��p�r_IzL�^��S	��yj�	":�B����x?+�"��Ti��V.s#*�?#�!"���t7�7HyM�� NDR�)�
�h�T��(G�&��i�(�G-����y���6STx��TJ�Z�]U�o/���e12%��M29�"F���f�I%���p�h�m�Ĥ�,)!��5�X66S�,'�Ӟ�SE�ei�l��I5\z��f���9�-Τ�N�k,�7;�J���גKOr�k@��N�OS�����x.�W�Aژ��0�SJ�Т����F�}MG��ݷ���r/8}���R>������2/G�/���{���e��	�n��uQ��N���c����Y�����]�7T����Q� v��Ӷm3~I�jÆ�ĸ�>�S2�N�F;N������:T��1Ŝ˺�J	��T�O}�K�Cɰჼ�h��vP��U�
�&� =М0X��H��>*ab�jh��~c �n�cX���9T�k�xd���1�}�j~}��9����5<
��2g���'�_�G̿�<�m���_��F��yBNC��Ɯ9�_O�Κ#�*u^���J~��d��q/�<0c�EP��4O%W��i��?* Ib�h�e�����{|>��k������q� g�:H���Jc�;틞.ڸ���h-r�v6?C��3�0� E 8At_���F�߳�UITW׊�e��D����6@��򞒽��GKO-R:��.,J�ҹ$f@�0�=I�z�l��sP'G�G1V;�^ZYߺ��=?���\ �tv��a�l��<.)b��DU�e4u����E��#f �@^k6� ܱ��Ď�0����r��w܉B#y\7�:�;�ׅ�M<��u<1�q��S����8�k��f�����^<�������#�Fn�a����ػ��qҰ�;߂3�fG[�iNu���1D��[����.k��:�N���ɮR���)I�c->�?�?r	�v1��`q)�_Edu\�,k8%��u�@�4	��лCiۓ��A�c��9t:o_��8Hs җv�TZx��Nٿ��'Z&�@��O����.��	�p�F����E�O�����g�vD�ow5� �����4�ل�DˏO��|�6�s?b�v
�˜���j��5�.إ��y��Y������k���%�U3K���q�ѫ�%]^\�38IZw�|i�8G3�pd�>��czƻՒ#��? `�|���tL��*���s�M���jK�Ҕ[��gg��*�A�^�$�&g3n4��E��m��/S0�� .�9:�]�(v��9lW��D��G��Rg������W� {�3���
o^$ʾ.v):I���MbH�����&Oo=ż���K_|����4z&ru��
������/�!z����#=��牉��`������K3b�9(U��$奙 z2u��G��7o�iq��Mg���S\y�7����2��J�j�-h�邋	*6Zz1-hx9ڝ��u�����z���8d4m�(Q��푰V�pf!_�����ej�G�p�+i�d[OO�]w��!�؂X��^���Y�����6Q`ǧ_~����C�Ĕn޾���>����M�9m�O鹟Ӝ�!�	����4TL�u}�ɺ*�j!�q����B������� 藏�ԎO���1�"�{(���� p�rι48��y�e#L���s������� ���ais��T��(.{��QV�X�d��� �P	p�1a��9K����8LI�lv�F��='?ifLz���Oi�>����� ����9pH�T)!��s"
�-ϡ�p��D)��F�H�"B�9ʦ�k��}�;����m:G�s$���T�8��������jK��V&)�F�m�:5(پ�y��0��4pX|g2_3co�
D��KZ�w9t(m�h)�G���������)y�9�IPc�b�i�yN�1ɟ�V2A9JD>Ǹ ܛrĖlD�a5�G��xT����IJ�DNX^L����K��U���n��П��g�Lk�͠Kkܙe3e�"x`����k���1�!�7�~U�q��`���e=����A��Ɋ���${�{F#�7�[�#�e#�V���r�v�`i
-W���Z�oL�����;f��7�^\2����G�gOsDǢv��Uꂤ��娫Lȝ�q�gX*�;iz^�r)ze�)��tL�\�#¢P���t�Hx}��٭rJ�UM1�P���Fנ���V 
7Э8Y#ᦑ!u�{4i�i���GI@^����!9��k]	�,G�Q^O�{���=-d�1���#7�M\�)R梥�>α�p���p��k�<�T��6�#0�\��(Uh��w��j�q�f�Q4q�'�%JX�D"��![�<VG�u�*G��R�d�|s�$��Y�mCzR%Q�����@J��4 ���_/�{k&@�QH��!Z���}��l|A>TEt���9U�'U���?E�iR��0�´���l��-Ҝ��:[.�(H���[py�Y�Q�4ZQQ�,U:��C<��K�4�٠!
}���tӷo�8�G�x:�$a 3V�&����9��,�\����֒EF餗.�y0v��l��1�Z��{ʃ��ƴ�/����Q���c!�O]�������a�Sk��&��v/���S��Qѯ�K���пq��U�.���GlJ���Y �u�|W���`/X�@�d;4
z�;Ӝ�����u�w��������{�.G�$9���qǙ�U�u�r�����p�q�ٙ���+.?lMDT�qUvϐ�KT�#8����TEEE�..�����1|����	|����  ��IDATS'lڤZ����r�9_.)���q}��ђ�2�oM<�k�j���^d{�x��f9���"I'���܄����bM4����j��D�ݮ��w{��A�RI���M�	���&,����TYV7����$�Ks�9Yx���9������<}����t�,�� (�H�ȰV�2��S���{��ip'2���2�-X�f����}zv�%x��s{�&
�
�Vf"�`��g&"zQ43:� `4�}9��!�"���.�i��ǫ/�������Au����ݻp��}�������txn��W�y=;?���֤$���}ǎ��ӄ+o����puu޽�f�D ��x���������ܛ�+���ۻ��ӗ��|�������C!�5�4.26A�NP)��S���_~�����	:���M�NO(���<ˋ��2ody\.�!Y��sp��ׯ_y|0�Z��9(��履~�钀 |O�!~��7{�S����+�0�>��G���w3N3�{1F��3�3��B1��� Ȃ����p�:@���}���=r�U
���n�Q�dOgcT�3�}ך��``G���.���ז�4�	�< ,w���!��~����A����=�`m0D|���%:0�-��_���<7�
�*j�� v��6�t(kg
��� /.QӾ${�6�맏���<�0���j� 8�Q�U�އuv|.��B�/�����t<[4�X� �並�s�@l�@V⻗趗bqvS������ �[�tܐ���b�+�6j��bM��'��h����JJm�ܖ��$�9�����>�g���Y�=~�@y�1�d�4�,�YWG���,�ba�@��p���S�`HE�����(���:O��{�?�}le,-8&�W=�9�dZ��y}�V�����?���޿/��l�n��8..έ;��ðx`�AfK�:��6��k:[	e�x��o����?:� d��g��)�=��b�u*�ItT*�/�&ۿ<�S��)��o�T���ey��u C-�ƻ!�A1����Dr�i�G�3���yuvO����1�/ =�V���	��lF�c:v<Pp��~LA�i�L�7_����,�Wc^�!���q����~(z��09������]s����˄�L	(쉃��C���+�Rc��?�m.����ɽ����PD���9��)���=�`�ԩ�f(yaZE~�h#\�k8&&��33q��K���{z�v�C>���9�!R�k���1tDk1X�#���t���V<�/���,{�y��r�����u�gU@���qy��Xχ�����ǀl�`RP�.U3�deu�����#Cei/!�q!p�{�!�z-��e=LV�db��=Y�ӗGA�89���IRYG:,��! DGMh�,W3%x��'UW]�!���:�%ݘ��j! �V�l�ٜm&�K�� /;�a�[��q��,�|�.���;>)���<d�/^��Cpͻ�&�<��WBk1B;Ͼ#��u|Ȥ?&��ط4>x�1�)����o��1���c��:1wd�L�n�nJ����a���q���c:���Ce���b��v+��i�	6|�1]Km��o����1K�@�V�Q�F��}(�W�?�̿,�|�$6��/&~gV�`�|ܳK���O���;����߲�~�XÒ�~-A�|�싯rl��q+b��9�d�l�R�m�PF��ށ��*=����eu�UY)�
�'z/U�� b0jn�ބ���1���P�����m�w�W�puy���B��M�3f�쳟�u{�9��o�uއ�aǛ���.�΄����OMx�!���,q}�w��U�`�J#e4�f�_�me������ܸ#b:��1���q}�8<X<m�d
�����4n�mee%� ^ߵ�!�޳3ؼ��uű<���/�,�rZ�P���&a�����eu%D�/�>����2�֗�Y+N¼8�Y �1��
� ��<;cg��Z��&.���20�Z>b�X.0�fZ��i��q�� A����C��{`��S8
 !b��=���h N[UxM�qv{#�t�'���2�� 	@֚��fV����x�}�Y �`�Dc!�K�:�Y8C�H�jW1���c�d�;���^mL���d��A�"�G�`��_����B�����A5ؽ�i:�MT�>�aB6�x�lKDu�r�r����������;*��Tw锉��Q�	YL8d��|̑!��̶ҵ:�a5�]:$�SW�艴�*�c�!�5���r�մ�+6�~����h[n"��a�?�q@�o��s���p�gvD�Zv��m��7X=рeh:�Ȃ��V>��� ���!l�;i���r�Fg�r~ݠk@@-�@@ 1eGܖ����QEgЩ�^�<�^���#:�ͭE]Oj��9�g�!���mrv�;���������xF�����5��V�(0�c ������(�_�8����|�3�k؋��}x�=]f�(4Y��o�g�=^������'�m!��hʭ%!�y^�g\{�}�]�~wMG ����A@ckg,����'����k`Ɔ0.���&����2�
�;�й��q[��a+a[�v �'$�g�Vh��O�؊M����Ӻ��Y�K�:kY?�X�5(�~� �a{�G4�J���rg�OX_n7�0�'��A�h6��qyrB�u4� "^��F��?�^�[�Yz���)[���t
"=OZ���o�;#�����WRp�6kNqͲ�(l�dm�Se���}�iD�G�n>[��Ʉ]����F�PtK!�o��.Bm~����j6몰%�����[�MVY�ю�-4l�>^~25��x#sk1�8\+>Ӳ���]a���gC��,,���V�MF����B��Z%��Œc��,�a�|��4�מ�Y�0�H I�P ��P-�m��1y�q��x܅4�z^��>	A���7���y��k'g.y,`�W`�?#�>(�+K����Ŀ	6s��`� ~x<�����z�8���a�*�ӎC���o�>i�s������[&#��Lb���
�L*���Axu���d��d+Ą�=#�9g
�v6�T��q��$ @#׀$V�'c[&���}�B�s�a��[���K~�=α˼�Y6��~7��~bc�$�|�`a�}��Ow��asBSZ�*m�<wwR�����^�O��^ni���N�dm����1x�`��J�l�˩����X��a���rʪ/e�d�NJ�gֳ<\�=���Lǫj�OM�qV����M�;�ckr���m�j>�(����C��ǟr�v�s,�2��@���a���ى����9�\,���>?�s9��ي��,k��p	[�Q���Q�v��QH�H0��%j�`�g��:�:63}rĨif�>|ތ��^�����<v܎�{��G/�����6�=��̃�T�WMi\�O����A{�>Y\��c:�*������_͍�#|�mM����y�?tuJ�Ļ~�d��jU�����:�9yq����8̉oBP̾,�2)�F({Ö��2�T���M��`7y1�w�7~��ł��H�G�-���(qu���f˼)$t,ʋ:�M��3b����^�	@h�jsD&�����"��`%UtrR�������31��������1p6�k9�� 0t���ݠ �L�byL(0(�V�'U%����E�v�8a����҃�hs��X.�@���v:��f��z�N
Fi$��A�!�	�̑t��	XV�{�r:��m8F�_�Q{; iQΖ�ǅ����@m�Zu�h23I&�9}�,C̹6[1:q�S�h%%���춵`7?��4a�}%���}ާ�0�ގN���Y�9��0�@-�[�Ě�{fO sV���m��w��9�ʂ%0(�ĩ�y��Y���Ζ��e�TU%�N؛uԦg�vq�����9�^.�l������Ppm�Kc��G��a�<�M3#�nnmJד��z�6��<{��Ԯю��~z̷��g��]9��
����HM� ��e��zI���a���v{��=�����93�7Y���GID��x�6a�W\	��u�p$���B`���d� ��Q���*��y`I�c��|(��ڻK���L&�rr@�]B�X� �~@=�>n�p��9���WAnYF �ꡀ�
zHb]{T��8�C��O(��c��;�֗{�5�h?���]��7��\����*���_9F���t�K�ʝ��`�|y��D�0648R���Ǩ39�b��c�2~W<�Go:4g�Ψ�3�Jޗm��G�~  	)���7�LP�g -T�ڇ��@f�Eů�PqO��6�c�{ȁŌ��]��߻`�,ث��Z�r=&Θ�3f �������1d��z��y�%c������'Pr��g�f>绛�y?��^��ƾ����&����Ƥ�9����mP�' �]�{��R<��oа�zn�	 KƠ�����M��|$����E ����P赠E��L��JwL�	.� g��Gj���O���NQ������po������� O+����|*�妶�Y	�B�m!P��*m+�z;߆p{viG[�l�S8wo���IL�t�t�r�U1���<����@��:���d�O���	�%ޘO�	v{IHa.Tb@��}�@$�#�ٌ_����4`�4Y�
+�(�}V�P�Kb��m���x.ԕ7�XPw���Ǝ'+~����������_~��H��|��?��k� �Ĕ�n��lg�ג�(�9<aN�5�E��$�$'31Hlԍ��YP\U<,�O��z���Q�Ǿ���%S��֮�jc\J��둾k�A|�٠,{?�v^Cg�tеE�
q�-C�/��I6k!~qy�y��3�W�2*|(R�wæ�Z���3A��"�u����m�/� 9� c�[��f&��1?g�nl�.�d_v��3�7�t��ix,�/���~P�n�� �+c,+���C%^��﬇�󽍴��Gi������	��\~�1qx�5�I� ��'��79��벧NQ��]*���Ʈ9S}���a��<nx傦8J2�����9�^_^)�����Sg,PI�y�^�Ih�,l%��`����`�����4�2�%c���h���4��LK����|{��D%�f^j�Q��'�e��Ϻ�����5���`ڳ����4�tn0�t��A!� !,�� ����*o�ؤ�f�x@?�1�����d�W�x?X8��d��Reu�<>����,�����f}�r����t���{����t��(bL��m����T���>Pl��?ܱU2d Y~q�u�тs �!�fļ�xcq-�t�U�5 ����l���\�]8��	Q���\xP`6{���4��B`�� �s�&�QZ:�N%�tف�C&1T�;�����<�_���LAǣ�x=�$��a����A`N���.|��zbJ��2+*a�&Ĉ�,���[�+2�GpH��$��p.��L�5��R#�j���C�͉��s��^�G1'�F����X��K�� ��:��̠!+G�ӎ-"�iA�KFp,X�n�JY�S����u3��S1��'�ʲBno^���{�p�������ڹ<�DJ�%G�L�m�}���a�'t=��?栏��F��₝J`Z/Հ���Y��('{�`��hv&���r(��y��Xą�C�p��!���_�5|�������Tpl���,��%??��8цg'%!���Lm-�^B��흑��p�p�/�.��؁�x��fC���n`,Xsnɏ�;����ią^>G�%�B��N��������Lн*�Ex}#�0ePx}I�@B6��_�11�uxDs�ˤ�.�q�z�f_:a��Di�j+�Fa��L#���?�����dT���M1Z�eH�`�b_ �?̸6����# $m�������/C�U,��;����:������0@`�g�-�(����� ��q4�17Q���_�s�h8T&ap����L�qmu���_]_�E�@�ݣ���㵴�__^�5�� �f�:������<l�3���v�Y	v6�~�
~�ܫ��<�D���.����,a.p�e�g�G(�/���gT����~55�^ �p=`"���t A�sC� �}�Q�}��߆��-�&����� �����'̬�2َg��\:�geG���b�m��n�TJ]�T_%O!<<h�t�:+�VWUVBg�W(@�&�U$[���_���zq�[1����y?j8���jG�7zb���`i����.Z��Ǳ0N8�����d���@�������x!C_�4��`�7�m����:c�j��zx)7!�߂�J��"]5�ێ���}v�[�p�_|�ɟO $�7ԉ��Z�� �S� ���B(&{�E�dtp����&c�#����G�4f�_�k�l��C	���|:.U�7"AqF_*l��	���a�לs���s}Q�e�_R�����c�a���a��T">cg���p��f���:�&�O�}%� �W�Q��Z�;$�u�m�Ͽ�5�/�º^2�_��w�㽕���Ş�u�7=: ��b
&�/�P�/ჵ���0_6���*:ۗ��� tƞUx�	�ĉ��lɋ�8�h��1a-�w?ɑ�����4�x����d{��8�*�RЫ�m8=s;��0�Hjq�7�!P������@p$}lFq2 ;)��i-��.)~v�g�]�F��0�&��V��Y�b�������42^��Y�Z�Ū�����l�9�z�V� �����#7G�S�W�Cц�u��(���p��DHe��P��׫�e��ق`&/<6�%7���	��N�<'�bF�H�b��2e�7gp�Tc	�P[�=b'�1��-�� ���.�72�?$uY`��'�7���2�
��%Z�TǲW u�~��~�l�}W|=��r@��8\��g�yϪ���AƋ��%������w,���qqC7�B�{s2X|~aeb�O`�P��:y�¦���,d>�C�{�����������DoN=�K��%[�
:����J& ��jF&�4�I&l��RͯlÕ!Hez�]%N��ԡN@H�øZ̓�f_P�lE�ͼY�cם�����w�)��,z���Y{���e*%o�^�`"o;�[�ѹE�����"g-CE����ҹ�!;v���i
jm"V�ֻcIk�}��#�������Ix�kؔ��x�i��S+�٬1�{��[0��1��牧3� �4���l!����I�c�ى��e�;��9�VX�y���>�s�.�u�Ӛ	0�vl�D�vg�٦.�����;�Vj�y�v��1���1��׿��>|*92���K�`����ӧ���
[�8�}��K�� Yr�*ch�'2��le�?n%�G�����?|���݂���D���W<�1bрN<�	6V
R9�gɑژMS�ן���`(l�u��,;X�q��݉�r��6�<�q���7=����!�o���x�4a"M�L
' ���)g�p��௰kҸ��A��]��0'NZI��y�Ǒ�3|���UL���Z���%u��-2�-����%��`3Y������:]��6�t�o2b���4Ya[�$������}��	v�y�36g��ݮa��&�u���5�D��)�NN�0��W�@I�\���Mؓ��V�~�;f9Y��9�?7g(�W=2`ؙL V����1ܳC�:���C	���Xڛ"M [X�ݵk���d  �C(�ܫ�ނA<�p���@�v ��|ܪ�����*�1C ��������`C��I��2������J��ˍ��h	�b�O��@�DO_���ƍ.�w�ƞ"����*�Y��p�P�&���g����!��O��!X�q�V���dA!|���7 ��L��;��I�`�[�4W6+��,��_�+�)I]!�=(#߬{3��?xbȆ��#�'b��Ŷh����O�|���K����XO�4�P��O��)+S��^m.�i|Ûf��'q�*��Z�9��b�GV��pjuC��K��3��R&M�1��+׏���b�6I�=�C�P�R����0����4��^���Z'ൔgoTq��M����ߣ1�1�p-�s�l��E��R�6y�4�0�S�ɔ|b��!ܨ�H��B����>�A�a����,�ʔ|�?��K�\_�e�˯6L�iM���n�j�i�Z����nz�
���Qp_�����K�<\:-;�8Ι�e�OMys��<O�ى'a�y� ˺K�����A��q�ߦǟ����!%�]3,����]~���0�r����x� &E6jCv��)Ć�:= <��Y��l4�-)��ˎ3Zw�<�f���m�����R�!Z�[�_�c���$�*%�/O���~�,@�MA�cXL9�Z3�]��t�8k �[�*Prb�gЦ�f�g0`aƀg>S;�Y�JJ���󈀶R��Q4_��ؼ���Q�:��9Xy`j���y^�;��B�(�I��-�T�/X�%-[s�3p��K�� �5�U��c+�5�>*	2G6�%�2.Ȋ��k��_J��:�y���Ih���NV��T��>��_�}����-����2����	t-Kv���S�h��>����}�L�����G�:�!�53[F���5�F�c'X�D��#[(2;	0j���s������iC��D��_���}\����{��4���"	I�0�D`�[xe�J�|�u��tM�,8K��CF�Ʌ��r�fst����y��:=�f���3�ڊv<7l(dgDi�P��3�r0Ї� �Rۑe6q0P�UKF�
T��w*(��zm�<�F-���F��z&�Y0[J@l"�[[�d蝹eB���I�U���揠�����^J�@�k㓗v�x\�e���<��I�&6�_'�� �S����i����ɂ�J�B�b��>R�v�7�af�&��~\^^q�2�����C�<;��wU��$@�MZ� ����y�ٙP��𗿄���#�
�n�ސ1��B� ���C��xJY0��E]Dq#:�Q��'�"��c��=�����O?�ϐ����OK�b��8�=�wa���@(��� ���U�y�
'ʉc��5����^]�9nman�MX�! ��_?k0P��Ux�	�׿4/�����k/O��o��Ҧ=y���.�=��P&��L���V�ɒ����o�.�c�	~zƕ%���ί�^���6�ٛ�<�V���Ӫ��|:�����T�����ZL��Jm�׀9�z}�]����cO[
f &x0]���S-K~��h�KpH{ƌ	o�O;=XY.��Þ{�&�e/Ծ3oTbT��\��X=C�r�d>�c�Q�eM��f��W�:��������Ō��e��g�������(Q�d[�n6��������L�U~��񼼐�0�ɽ�.�Mõ�1$�c��X���왑����8~�I�%C�G,�1�m�?S�{=�������E���Q�>�=�ȃ���5�(�ǽ=?0}�m'�
oLo��������H��]�T���jE�$Qw�'`W,)L��4��1q0.�=����n��ܖ� `�@���l���q�DuD�O,�*vG�;cި#R��ż(g��WH���:�ύ���hؙ̚L��ǽ�>�kz����%����}kr�®���Q�g`�T�`>fG��5�q/���Vᮓzb#Ɲ>���u3�#ҳߞ?
�{j��J��o{�m���{�Δ���T�	�'1}�D�j�I�>x9VeJ�*f��"h�oh��<YJ ����h�����n\ Db��f���&]�a����+s��o����}�n�?�¤�w��b�.����|�}du\����l�,]�yЫq�s�Nz��Xkv�Y������7
&����"ۼe8��
;׺�E]Z�{EN,��*�(�G{������]�p���3�`� �
6>Q�,�P�?p�3��?��L�������J�R��Jv��PO&h�)����)XO�� �08��t�.�u�ʙ��щ��x�(c���|���ߤV~��Y<�j'��}?����e���f/8���kPs |h�� -l�7���� lU7�"`�dP�P�]a4JL�F��Q�/�Vb�W
�ah��#�sq�a�����<���8����"{�29R�7�j� �j�a�V����ɩ���p�~���@�uƇ���y!އ��;R�v�������:�`ӯ�9�N�(M����p������Z��D���P�$M�\��-"�K=���;�EG�* .0x��tn���8.fk��c7�]vns vG�!�i�|T� �5�<XЋ�CK�Otj=�(��l������KtfZ�:`��,��f�n^�H�Wɘʒ�U��R� �f���Q�b���{��|a���/<�/��\,P�qf�~/�
ej��;g�ca��k����Y�Μ�W3�m��Aݴj3�*@B`'?����U��+u�ٚ���NCv�C \���rOe�PN�n����F�U��9kc�%	I��/Vj�
S �r4�Jd]S���T�)�!uӈ���k�Q�
��:]�8.(n,��2'�L�!�R����0�Z}�U�&�̏%���L���#���ʺ��(G����Շ�~��L�/#=���G�ɜ�W��/]|�Qf�-�@�B��;���+megl��~���s�8��{p��A�����giAu�c (��vm���{f�� d���?��yܹh���CQ�$=���e�r�j��4��gӝ��&�ͧOt���z' ^U�[`#��i��1t��=e����f B)X˅2P��|?��q�X���8T�/������Ʊ\���+]|����^���ox�8�Y����)����[�x��GfLq!��[pA�/_r�?i\�^?���($?V5��,�k�+Cl�~�$��G@׳�6N���H��}f|?���&�<#2��ٶ��r�$�`l. ڦQ���jWl2ِ)�f�+�O��F߆�!{��%�RRzo��lr���\�����9�jQ]YS����)�����@�i鉉�\���Hh�Tt��4�uO=��m,�����E��3�j�A�v���=,���,���Z��d��Ȑ���3�6�e��w��h�L]@�w�r]��D`
� �s����5�=�Dl�N�j5c�{7��M��Xu%9���5Ah%")v�>����h)����32�([��k�T���|��D�Y��է ��:�O���ژ縁~��hK�_6�-�8�m/��3qX��%���ԆK�k^���b[�� 59#����a��LB���6���c'q��A�����~5;:c"q?R3�hq��7C%=�X[0:��L�Jy����tj*�.��=3�,��8kҹ�|�� ����|�������;]��'�g���%X%;ؠ�4�Pn׀{�D6���ep�b/kj*No��:���:��`uVgb~�}�]{IVc|K�iCfb���7f�~�О�Ӹv;���ԏ?��ǿ��S8lwa���>~	�W���.�����ԉ��W)cn��ue1AG� l����]�����ZzMU�*<�p~�l�Y(-��X~��
�F����#s'��KT��7M*m��ޡ�ē��Te��@�F��|P1@<��w�����'���5kO�����a���2'�LQWmx>`/|��ܞ|�A��msP����3[l-���S��J����y2��FfQ�,�L΀V���ʧ�d�X�?}�~(S\������G3y!!�t���4%��A祾�M�hA�i��b�gF]�H� o����S�1Ci˞�S���[�x�� @�s�:ﺮˆiۚ��zDA�٥6M!�po�����st�9�AA��r ��ym�n������2*�K���Ѻ	����q5U�ek��*�X.�����U�~r/m�7�@ą�ύq��bz��`4�g���;���Y���ٜ�F���/��۰��UN�JC@� ��#��1���ʌ��SE}��Ȣe"KVBm��1 �֌gM~S�	@Ŭ���dz�EwbMa�ݮ͆��N�="�a}٢��wdЩF�P�>��k���w������<�NF}��: "��z ���SO�����W,�g�T4��:�&�և��"���х#���K]�lӦ}�Y��6ޱUoR@�%�z�ȷ��6�-��M�s:?���KLC�-=^~L���@ٯ��ף�Z%ê�1 h���5-(�����&6X8U�� .��?J�b�'H�θ&V̠b�>�����&Ⱥ]��;V>T+X#X2ڎ@g��Fj�Q҈2���*g����3g�H�ӏOV'*L�Y���P��v��l
�
�ː��wigH��ֿ�ho̎���E�Nb�%�O����^��r^�b��qc7?>�Q $��.�ޒI�(���Ĳ��$��"����Bqa\��vm��� c�:}��),<9�]�h����;�?���<�9}}⸕��œgi0�`A��ؐg�s->�$�4I�y+�W�J�sq�����x-��ńQ��!#��2!�v���i������l&K�S_�&�w3:�֡��DO60d�fd���`�VW_ؐ��Q�ܛ�>���f:!�O�s�S;\ub�q2�+k`#�@� J1�:2�a{�Ek�,����]��^b��q�*��e^�U~�������ȑ�$�8�oo�޿��� X��d�|�	����{��S���N �e�q�]�<XR���~��¿So��&(Lo�V�D �2��@�0�+v[���xh��`Km�GE �z��������aǴG���t]M��0�� �U�ts�$I�L,����,�@s0=8�Y,p%�����@���݊��l��y���=���Dc�w���d{@t���H��%����+�^��d&�=��_�!U
t��#� �4������"�k�X��)��Ĕ�~6����S�R�:���%M���~z��]���xt�N�K&�'�4�@s�!p�m6s(9&x�B_
���^����#�׫�ww���&�LZ8zQR���� IƪZ�9��t؍��
���{��h;�1JLX��Ͷ�  ����)���
�v�
�d���b�R?2�I���c�=Ǆ<���|����]�'�jA���c�$�v��6)_h�K�A'���y���E����io������H�Rb��6�˧���~]3V9^=��:o�0�=��XM�:X���c�sz��q�u$󪞈�'�怖����sNF��tZ��xr��_���d�Yj�[�	֝�r��<Y�Ϝ{}zr)�?���N��>�2�*��P�ʺ���|�I����C�Ɂv���7w��I�p���Ҍ]%,{� O�t���[�����T�6�]�����ZZ��f�o{˰�S�Y2Bft��8�=���|�qT�K��aS�XU�!�ױlIL�`���@efֱHY�I��m�l�8��3�pFa�L$Q����u�p�R#�{�k�wz��c�9��1�>pnZ�y���[MeG��1XQ�n:b�I���S�(��U���lE�H�t�,�*;�u�(t,�m�� '�AQ�G�$e��tm� v�24�L���	b�b�4AI��R�:�]>�:G�ًUU���nevL��Tf���Y]jf,���Zp�0�(�=ٕn��{]e�����/�������c��P��!E�RtvC�#9ؘՕkL$qQ	�u�����E��}���K��I����`y�X���|�D�0��Y]����
-g�%�+0p�k��X�X�k�W���h�OdS 8Y2�vo|~4x,+�P�u8I��˖���zY�4�{�F|b�N�/�Efڲ!�6��O~!�	��U��7�a���#����-�(��h�q�jŠ�tjZ��ޓ�'P�x4�s<Ƕ��x;喁f��6�����	��`k���6W�ys�y}�s}���ޟ���֎# ��p�nr��K����}�^ �H��G:������W�Ta�Bw���";Eg��(IΏ��_�Y$	\Y�`���ب�9Y�KX?Й��{G��+�����
�C�e����}��ba}OU7�h�1.���@S"���oW�_����?�����(�YC�Bз��%�Q�=y� �Mw�d���=:�1����NA%_/����.1���QY���uT�0� <�68����3e�8�����ˡ-z6���Q���`���av��=C���J��C���R�+�^��[[B
`-ŅQv����]!�uc=������%� |k��-�U)� ��Yj��� Vh���6���.M,��*�뽉����g]K߇����_�?�`B,����Z��\�af>�#��l;��I@BcM,t��L{d0�A��M��2�jP�������@¯,����AZJ uؾ�V�t{x@��v�z���^\>�f��6d��Tx��T�)�S��U4��^�"ɻ������|~����@c�{�A�(��-�v`JնĢ���� ����t���`��54ѵ�����4�a@&�gg��Ղ�
��&�p�6��~����>uқP:<�r��p@��#HE��J���!��Ǚ�%M��bc��w�Q߲� N�g��P�~nw'�?d�"A^$��6K�)3���s*��{���R�¯��>��޽{���gb�5�,�"`�h��lG�E�S��dlV{��;ČYF�xMq�vǝ��ƻ&�O��&����]�.�ߋj|�` x)��mƇ���G;�H]�9Ja���H�X�I�J�ۥ��H���=J���P�nn�T��f�hT�ٚ0����-�9�n|���pB�q��/�M�C�&\��������0ڂ��);0��B�sڭ�%�F2D�pJB�@=f3��O�O4�O��c��w� �����Ӵ� 3⮔o�~���ӳ�����.3��o/(<�̛`ț�6o_?����po�dOfA�l=�6�M�Uh�u�(�1��������VO��A��R�ק��?��&9�,9� �G��2Ƥ�ùfH%��sA�N�%o�����3`*�
2��e�R�(��?�m�eV=��K�x��}#)��;uԓM5��n��ٟ0\�x���蘩� i�Y�P��lEGC0��������V�0_H�P�uɄ9� �YT�*�`so��@��N�J�����XB���7w!\"۾��e���4�����%K�:������&������a�R(5�m��g��jIC/!Ն�ۙ�w���PK��Z�5P�si�X�x<т���C
�:haF�h��P5v���r�z�@��m�l��۵ZʮT'��e���%���87���܄�����߮��B=&��!} �p�1�Qb�6���z>�r���/�1�1p�Z=����2s�X^�TF�[�\-(�Ζb�ƚ:�%�It�6�9�K����˸���s
��l!�l�!��Lm(�J�9V#M[0���P�J%yx k�Ƀ�۲s��L�{��M��V��[���it�'�kb�bZ�>��G��~���Y�e
���B����
���0X�\Z(뤳j��v�@�'��l�,�`��q�n�Ԣf�hc-���puŒ,��7�>�>~��x#��2����k	�;�pl,�0��:��
�`o,$ԛ_^^dG�.|��(���ڗ���!�?���C���/d����|q�|� p���I����Dȁ�'����MF ��LU�v�Q�I'��@�������0f:X�T�9��i����I��3X�h�'����!��q��}����Ƌ:-�
Ž���A��6r�N��RY�b�2���J��ii=��?�n��?
,k%d젽8:�A�����w�*8�w�t�'����i���3I�����&A������%{+2+rݓ�Kw{�����b����}:?�.T
 �i��U�ظ_����9K��&D��d߂��[Kjd��3��
���>2`�ÌyM��=Jn��P�Щ.����(���}`GO1��?�>�sc�{<K���x�UyȊ{&\�JaG[��)�΁�����P3���m#-؜�j�`�R��JL����i�x!�s�}7�wLP����,�Ն�PQG�/�/�e3�g&�[p�`��勶*o6=����-��5������$�R�6��h4 ���&�7��IL�QQ7Q��.2>)g%��pJyH4&��[��ܒ�*?��u�kf����.L5j�T���x�����'��`�FIQOm�I�����LEE��)���_<�WrJ�������.�D����6wYp�����*ź�Z�}H�|x�>�������|�~q�c�#�����A	����>���C-�����u��3Z�\�x�?�<׹���lj�Ix�g�ݍqd/U�a%� ����߬z�� @���y�ߚ�]l�fF���|�sdI�� v�O8#� ����
�9Hϯ�>�B���P>�<{�qn�"r�=�%�q/0f���?�Y�����{2�/7��Qh��wŪ�����I��h�:���|D�c�y�/k��C��tm��y
�'��N�(C^t���)�ߜ�&p�=���8O� w��܁�,�PZ�����7`j��`�Ԣ�h���o��~>~�����tP{��X&�����p.����-ˢ�6�l�枎�4���R�uzQk����ғ4IzRf��0���s O����.�[F�8��!�/�ٯB?��%}O8��ŕyMw�	3�7�Mp�u��L'bV�œ���0
��� �g�����*)AOkۭV#��#3F�T����B��]Z���\]�t*�19
%�Bg��2|�  ��-��C;p��̆��6���LkgY4b$>m���g��h�� +��Ƽd������^��l/�IA_�,�1X��}�VT[XUt )
��/��xD�Ʋ��16'tECD(��������*�-t�V�pqu..�s�a�uE��CƖ��(��ya��h[io얤]��X3�,KB&lP� �����F�Z(7������P�'��e�-k������>��-��`6���_�G��6�j��I��;����L�ʲu��]ºdUkfx�1fffF�{�
J���1Pǆ��Z�k]�Sم��b� �|��QCH���Ų��1v�a����f�^H����$��/�	�9}�4,���,�b3�g`��v���=�u��ҭ���A[v:1L�Vi��҅�TU� �ejhG�1k�e��5pFe����z:���{�3�v���� q��#����n�X �\�/#��,!�-m�[��<m֙�����}h>~�Ny+��.��ÿ-��R�95]��V6Y8��b�@ю�(f��\$����gە�:H����b��Î`<�3h���I,��͍�橗\<�=oM�^����c�(M��mG���1�~^{��jB�K<�-P���㩹�@��o3�(�4M>��������Vf�.U^�ҫ�5�A��(����R����c�|V���G0j��2K~�����D�r�/A��Y��DQsl�A�p}�rt���`�����*�X���(S�S	"�!�=�7���g�eГ$��L��)�Y�Dt:`Ub�+�)�)p����f�ݐ �</��� �h�ת�qP'�|�n.�Eܕm��YR�/� ���w{�l�a~ւ�O�ֺ5�G�󅱔{�w�����@�|#��b����a6 �/K�&s� �0-���
裗���hMT�>���)ݱ4�`���e�R>
;��Q��:�����B�k1��D����-@o@RYR��8P����~���=�s��fUY򜀧�&h�L�N�/�k5�k�;��~G��#�����x����o'M����	�aC_L����g����{/�;�����s��H�}��"p�V�W ���P�\��r��c/�D9X�ލɁ�7�/��a�w�P��XOH�������$�����tM|�氃�����G��%�����{&��7g�o �b��QN�T|�1��`r��H�AmC0MH�$�CZe]�ꨍ���^���:=�Z��I����P�%F��n���縲FAS ����y,?����<8�2����w�(��c5��˗ح��.#ݻ'ܝ	^`�e�7�/#7'�����֪x����*��kS'j*��-��X���_\h9-c�*;C���>���Ro������Ob^0���-��Y㲥����lpތ���O�����
r����Ք���
o�o�����Qb&ˍ���4��hj��N�Q	=�Όƒ���i&��(�e�=�!�(~?R��N�kGN��k�&ȩ���A�0�h�p�����JԖ�:���F]���n,���Eb��v�є�-�n�t{:�RQ�z�"�;��i�G�K�ӱ�<+{s,��0R��5�����=?�1���n�K��q��$i�$T��.���U�m`+�=����<�o�{��� ����܎TD9��9�z�h�j[僚��Xޱ�EOב2[Q�j�2[A-f{��|d�Xv$p�`ܯ��H�Ӊ��`7 �WW��bi��s�#����ǹ%m�)4�����.��u�Y:X�dYb1��w���)x�k���1؜�n�(�� N!sDYJ{$pH��.o֕�ﺦ/ &w�x�#O��i q[f)�
/�U07��]�L����b�`�v�ڸ"�&03�&�8�H1~��脫�P�~d��j�@�T�QPp���(8|R�!�����i���hO�k`k���halAcg�+�c�he��t�b�u�S��~1��3r�% ?�U�C�����u�@;J팔Jm5m+p@2�+������z���E{AedQ��v_��]��)X���3��P�i}(����]�>��r��A6�l!��z5�l�X�~��9���o���ٚsk���a 9f����0���~ g*��8?��2�t��׋�>��7�>'�%��G������'D�a@!�9���VG���/#T8 ��u�������F�\����	���;��1�˿���4���e@Ib��C�'�o��+�^d�z�.F���Z6|A��Q%��������,m{c+`�%�;�����	0c��֏��Q�>ij�`~�b���|+�ϙB k x�=�:`���	d�LY�����Vn��	��L���-�H�X*O���I�ˑk%��=�[��6��7C	�J���J70�E)�7�Jk��,	섨�Ԥ�Zq�'9�7�Q	����A�0�|��`soMݱD{�#�͟��.�X)m��B�ߧO���c�%�J��&^\�}H�@��1}G�(A@�o)�}�$���rf��*1���Rڈ�o�S�%PO(��uC�-�K^I�`�;���'�=��r{#�?�n�oC�0v�P�h@p�<Ha*"��w�<�]�%�×S0?m�<z��ҟ^4QO^Lo��7zn��<9�ٯ�@�ۂ�op�dz��d ey�Zs�c'�}X̗�[;幂������.������O��ϊ��ݸ̟=�����OŮ���9(�O���B�O�#�%�s�W�������w߇�w�J"LzL*'�ެ ��,��J�[��CR���������_��,���K�����1X��&�D��Cݳ�-޷��g�PkR��D��&9��|�b���%`�1�燣	�{EIur�}_ږHH��M׵c�Y�w-� 4Jǐ&��c�k�4�yj�
�S�k�э#��=E��&>L̈<�*���[�xq�cڄ�c�x�q/���mi��N���X'����u� �}���h�|����6
�;Jٕ��ۑ�o�铀R(�����W��Nm�H8���@�����r�� ��IA����	��(Z��9$3Ӏi�JL����n��C;v�*�s+Hcc#DQYm�Nw���B3 B�4 ��9��l.G��P͢߻�t�Hv�ib�ȶ��7+���7�8vĉU��O~��N[*SC@�4Q>83f����2���Z�u2�M4i��Fc����Fr��@�`�&
���1_� j�̤��٨QG������F�KU�c>.@Jv��%��;d�,g4V^bʎcQ5�n���TBᎠicP�et�%�i,%����׽Ƈ���邨:[Ҫ�-@ 8�ip�J ��d#��rn�j?~$k+ϛe��5P���V	��tv�dJBv�:;�R���X4�]$ㆱ�PK�� G�'����Е2���(�Gr���bb,`�D��F�Ne.%Υ�1��{�7ۆ�S�߅��(ƣ2�UT�vtvS�Oˍ�̝�:l��ԑŲ�\�[��ɲ�Z#����M-j��ŖOY;�)JeK���9W�F�*��d�F?N�?��퓳mfKp{&�rծ��;��ك �`6ޏZ�.E5��&��E�Ft�Bi�� ) �mK�V�'p��=��-���x�1j-@�i%�)�2�Ћ +b� �)b�R�W�L ��Gv����+��gO(���} 2hX[sӽ��媵9* ](B�Wc±�.�u±����y>�;t���% �[���oQ�1� �޿�hk>Ηϟ�?��?s��_H=���K�zx�t! T=���jyf���}��!�ft��ƿ�#���Oo!�lvE�DW����:Ɵф�G����X��������	�:9��S67s*����}3��ӟ���6&��F��f��8���!�dݓLs@�U�ɽh,����K���J��RAuT��O�!x��uk�'8LJ����� ��ӽ�?3�����Z~7�Q�V�ߩo�}�:�{>����k^�`��T�[�E5JF��,��!}( 5���q�2�����XQ��@�i��,UE�˚3��^���H�����1k���� =�ZM?f�W����0\�mأ��������G�������@b�8��LJ���4�Q8iB�O!�o�6�K֭�P�DQ��3`��Ԙ.���TYgYuRa���۾��}΀���d8s
أ�./#Kf@Q"���||c|��y�5C�;,���ӽ��TC�2:�FqPPk��H����ro�X�l��|��Gs�f�|�����#�ό�,��A��O��'�����>�/M�8o4"�G*�T6S�>�&�M���U�/ aj|d�1��t�����p-h�=G'<�`\�-��k<��`�,q:�΄9]������j�{d\�,5�:%�Ă?鶑�e�T� � +�3��w��'�:�1���6�@���NU���K첍Cc�;�΄�mM��`��<C��uX��Ù�7G�ր"Ə!����'0Ҏ�z�IO��� �ּ'�ՙ�*�A�uQ�s���szX�:�
A'Kp��u�Ӌ�I'�y�3��ٴk�+b� ��t2A�?��O����x
�OI���������i/rr�Oab�+�e%�p��l係j�>g�j��"\�EV��o�����^R�X6Ѕc����c5v\`M���0^�?���A��Yh/@{׸��9�~y�l�_��ǳMm�
��h3Q����ćǩ1�ӫ$A�e^!���L��2=/��k:^��5�j	
Vʽ!�Ǳ�ɲw(��� j?괋�L��^��*��)$�LA�p0t�lL|n&�9<a �80H��x>�T���q,N��cocamSCoea�5�6/���3�H�7@���  �&��c��d�l�6��{dy���dtӚ/"ۣ�1��Ї��u�{G8�
cG-��u��ܫ��Z"�j?޲+��,8�&���α�S��9<nu���Z�X[Ag2�D��Z-���:���:s��o�b.�eCd�;ꊑ�t��Ve7�C����lV���Q��+�l�3��8œ��U	��FAc�x�0���4v��g씵��(!��^���x(� ֐�I���jY�4t�U������8���>(�����ׅC���d�cW�j����o�m�92���43�֔��v���	hBt�Ǿ��X��@�'�w�2�ᗦ��1�~�n�l`�dH0o�:N���A��l&�wstӁ��E�����.)����9,��#IZ�������s�N�B�3�VF�׺��(hN�V�2��w��	X��	����Z�����	l @dq	��1�����e{Э*_�U���EaA�N}��%4�QJ��]?��c����{e�@���{�t����;���������i�	�H���pUK���J�ؗ��3}F�\�li����/�_	��O�D�`��c�L�ckZϭd��Ԩ����Ԗw��[TWȧ���»���7���=��P�ѓ�UBU�o� �ૃ;�+
˻`z�c%}>y���'�i��>M�!T�ɲ�����f��3���@?�X�Gߓl5
�#i�y�=�]���tG�A򩖟�f��`��ZE��Qk�j���g�h1�������1����Q��5_�J"l����vC�x�#��r�!h�B��!]��-�oҖVJ����Gڌ��lG?��a&'���#Q�M�t$��d��̀s+�$J�h�7i�95���Q��;�Qs�p(�A���4���}T{fO��]r&,�g���>�J`[�Π:D�]�P��qO��F�.!�@J];ci���1f[T�;^��2��3��q=t0�s����9�s�!�vyu~��{�_ $�a��()�7G+������'kAa���l�����+�;���nG0��0�a�$��RI�u�w
�M'�y?3�x]|;��ǣ�o�� xZn�l<ds������ĖE���2D:�9�-i��v�`I�ʴ��N�{c��1j&f}��y�P�4��Y���ctp���0�x,z��Ȥ���KO�d��Ė�%:V�_�8�'��zTU��3��@$y@:�1�߅�?��[�c �̤\#��������������>{)�H�5�(��z9�9����>��5���§��e��"ǵ�� ��s i�2�G�����&��F��j�s��=;�0Ƃorsw�D� �O|�ryq�Gy)���Dpg�υM$��pnaB�9���yX���%�[{v������=��6�>P�Yku]w��,6D���+�̭\������S����j�WB�%��g߫5}k�B4��h���)U���t{�����u�f
8<�����z2QN�t�\����LM�{��+�^��R[v�q��̔��v����b��S��#D�n��G:�����8X��Jv�y@e��30L�5��^x2���n����A����X�td�&���6�.��J�}�Z�C�:�D�m|�=H`6@�]y��/����5vfY��c0@@i�`ASGfw����t;Ws7�yЦs2��-�d���3�Jy@o���j����5���:���k�%}g-)nZ�x��� 0/`�� ������Y-)߫zE`� �{������!�*�p���W�Z-�g�@��[v��[ߋ��ZXP!l�٢F�}���	�>Rl& ��s#B�;;M��t�V��	
�}�k6Q#��p�삅l?΋"��!����7_�.��F'kY��2K,ㆲC/�벓��� �zNGK@ cM&OU����6�4�Z-b;�p�-�����=ڂ�e�xպ���pza[�a�Z�̴����"5����D]3:�ut�E�K���rд6M"�7�;�4�:n9��_Ԅ�P����c3tfEp�p A��^��x���l��&�o2��e��������9F�`�q��0�Tְg,��ڔq�CGf��4\��dש��&��M��pw��MBP������9������:�?v=d{�a�,3�jˎAh��MdOpvJ/d�5������E�"��hzyyE�n�RG2v���V��
�:����zq�c~Y��rn��vf��uwj�띏=�Y�P��t�#5{(��P�E�GJ8�M�:��Uw�-�m��	v)��ĉg���H\�}��w$,*{_�x�o�MK/O���t��ct�F_�]g1�����-�+�v脑I����F�1�F�����g�����	��'�����E~Vi�k�?G��wd�&HJu���e�x&�i�� ����[��X���'�`P�k��ON�x��L/k}&���)������A���y7�����u���j��;�#ӻ���L,�[yq�C=�Ūt��ɻ�}� LCp`ĳ�~���s��Z]M��%G�� �]I�j(]��!�I��#�ܑ�|Q��C����Z��ٓ��X��x�:��^a63Du�9R�󣱍i�ؽ*__�[�Q�[�Z~��^�d��{����PC`�� ������^�����lz�' �h.�@�%�ݮ�j^A0����~]��v}��|z㤚��7)6P'��I@�`B���_͠=������68���b�Z�%�^r�8�}Xm��i��6�Ω����ސ����M�[v�s��K�W��u4���D�ww����I7jAz��Z6n���~z<vb����I�݅�OLܓ�g�PǐJ��X��#��m�����q`c���Js+ϗ=f��|�Hm��pqv�����+��� ���d\�%��V�iq�v���6���˝���a�d� �_8|�<�ٶ��)���k��B궖��6>p^��ۿ�kߗ?�fs����/�~]�^V9&��˱պp?��/b�l�cx��Z��`3{J��X:#�Vd̗�e�//�b'{����_ �{��Bqf���(A'<
K�hQ��w񸤿��/7����Q�c� 0��Ĵ{%1=2w���<�H�h��flT�	�b�������0�;��	��IH�MZ�(���}�Fı�����Gh��`��!PjԸ���?~&�ڤPYu7�v^�i:���I�^l���Ke�
���0��m����hU�(�?�`9� �G�X^�k1���6�c��� �)�e�gl��,-f��h��S���YݢDt�p.�h�m'V�ȭe�q���` �s���m����w�<��D�U-�w���d{:��l"�	����Yv�9���]_�nX��_s�������Dq���U6��<`�\<�I�%S�z����n��pL��+�\�6Jc ;��I�`B�`V0��^ο����Y���C��}D�ɶ��0,j��%� �U�C���2�R�*E!>���g ���U#F�oќy�uMd06,A��<����/�K�Pn���z1F ~��CD:Y@�I]I�y�B֎]��X����|;J �ы9O� ֵܩ�8F���2@J�� *��-(p
-�LG3�Njs�4vj+�3lk���-����,�[8�Q� ˧.θ>��L���������н`�(�����{��Y�/�� �}u�	g�Y,��u������<FK21�����v�bK�X;ev�����OYS�_ڍ��Tv�/���_��ԛ�9��K�4��������s�� ��:��no���=�O}g��J�G����To�I�DQ��e�{�T�MN�J���q�!>�ϐ)g�G���$d��Hر�����|�򕉃��L_�J���ў������>|��l���0#�	���������7�/��u�ܰ�|��/�{��}x��C���x��&?~�(���d�u8� �8���nU���ԁ�	P3�1���'��+�#���������/�%������A���Ե
1�s/�Uf����>�)�b��O�x4��Ϗ���pJ����Ig�>�%�W�/�'<_�q����r��Rjb�'[d�#;Z���}뒁PԷV�Z���M���m)�dצ�:�Lu�K�8@��F�=蝶�R�ש/�و�٩�Q�/�R�D������S0�� �5�ϵ����yWƻ6QPԖ��}>�zc����6/�:�ďM ��{��.�T�+�w��� w�Yv��4���;&����D�{�+�C��'(�>����crf�$h�n��G&u��ofg#���u%����]/p9xcq9�H��Q�R!��T��αQ6kP��٤�㋀�`�D������_^]��2zh��s�����5�j ~VW2�W��C(e�C�΁�!Wp^��F�Q;��W�V̍%�*c���`8gR��Z[>�'��Y2�����j#��2r�}��;�e��*}ji�HS��]�%i�8#赡/LM�<����)J�������H�)��Z������=� ���s�H����ks�]o,m�/��#��*�V#;���+�E�g�h�Ԝ�"9�NT�ب�ހ�~8��`9��ϭ�dS)�3��/?�B�*���qO������Tu�<]���q$��^f���?�����ty�����>���O���zr��K&��Y�6����m�y�<������6��@FM
����K~.��r	-���K���p5Gc	�T�_f1RH��J�(Wm{����"۴Uc��l�9���#E��k����U��}s�_�>���� C���@;8�t�~�����k��Vb$$&po�>�C��w����&6�e� �ON#6J^{���hJ�eɰ�#�N�t:�OP�q���F�,Г�����`�_�<;��h�7���Q���x*51(24T���v�ORY����3���h�y�<���U~^�����wOH��t�K}g+�R���?�'&�e�G��W�J����`�������Rԕu�6����%Χ:p�}�둓`Ƴ'S�4�8��E�:� �g`�A7}�ˁ���6w�-��az��ߟ��Lc��J�`Y��Y�4�t�!�C�]��# �v2tV��l�c��V&���d�ʵ�x�.	佪6#�����Ke�W;a�KO�	zf�嬱�|մ�]@ژMp�	�5�	�A��ˊ��$5x,B�k�e�X�``�guSa���uz�%h�p��C�6l�0�R�?�\��G �L�2~}�WO���+���as0�p��.;���7;�'��V�L�I1E*�L��O[��)0�4b�T}ь�IsB�6�C�[��y����*�%j��ʴ�
 l
����ǳ�
if����On���^��$/�Cf���;�uw �|������n��79��y X�5|~�С��K�&}��5��1
Ŗ��V=���8/"�0�~8cg/�|�p�����y������ϟ���T|�l3�"X ��FNM��h � ���^�ad������k�ram� x�Ei@��wZ'X,��_�2N�M8� VG��朁�r�ޅ��ߓ�6��:���33��U�{���X����oh����ѶH�
6W-��J�,R�1K�r��[=E�on���Q��՞��vli���t�a�૛�P􎨕1�[W���u%�㏶����<衵�E�X3	b�[��=���2o����8���f[ۉ��Xa>�ϟ>�s� ��Ap��bǥ�#�晥P:��~���Ӆ��tRG/{��&n<�c^��7Q�
VzP��Η+/�
&B�����*[�=��'�#�XA*�QFT����J�~�su�C�TJpKiG�����ů�{�$���O�+>��%�`M,��� G�zYH� 8�������)�>�߃wϱ�K��Z�����אtj,ӽ0�9j
R�U���,�Zl�J�@t����̯p=�����(P�����]�u�D
#����k�+�;Q��"�G���L'r��U�79�F�x$������[``�1�Pv�D����o����� ��k��6`�-Đfb�qgs�|h,�䕘��Ic��8���%��*��t�E�����dSD`�A{c�L��J�F��)o�u=>�nc�[�%p+�F�����`-���e�Zki�i���)�b'���8����~� �B��'[��m��s�iom�7�����
o۾��޴��$It� ��wefeMWu��~���OveEVd���:3����_WU3wɗ�5�#ҨB���fjjj��`���.��a�Fie�[$&��$쨽����L�b�2)�dh�7 4�����'�l� �\/?7�`��@��9�F�M�y���k�#���.i? ���1�g�K�ł~-R :{1^?>�Cl��0<�?r�,�_�@<��\�riLz�Ӑ���;k$�lƱL,�2�)����Sxح���Ṟ^,��נ���nX
T_1��,��}�]`�#K��#u�V �g~����.1�
��~��[��2�Q��
��tՔj]�!��^�ęk���*������i.
Ͼ����mfq] �p9|�p l@M��N��C�<��dʛ\���x���u&��֔���d�'Z�f��5�������y߇4�֟��v_o0! ݳ�v(8\6@Ys��0�B�����2��~��G4$�&mT�<OՉ	�E�m�.���ԅ�o�:���>/>0O��`s$Z"p�W����Mup���}��5�8^R�Gm4[�m6֎9X��k��G����q���]#;�����!�uyuN-
����w�>R�aa�Å�5�� jL���X�-���T�q�_ʎ}*���-�����K�"�.�\.@E^�0��77{9T�%D�1f"����	aj�S^ҩm���������B-*X����l����m� 1T>u�߷�dp- _��S�1���"0(�A�ީ��{1�p/��\[{Rlޖ��@��#ՎN:e㼑@sߩ􊎸	����%�&Ց�C���9��MVn�4|�ǽ7��:��)��m�L̱	�as�>eg ���/�q�qW`��Z�C�&�:����֙ �\�i6U�h�����������D� ��$(;*|�<��h��13t�#u����Ae�Nav��o.��TJx)�j�FZ���]
�MJ�/�B�~�kP��ZTf�/��_>��2;gCxs�
Gg+�#C'��� ��1o��u��G y:�����b-�r D���ɦo��~���.0�X�A�?�i���������1�}�@mgA#؟��������Z�>��gg����p��
�4k𽰫Q�X�����0
�zdg��]5�֎�8l X��p��w�wr>�ب��`L9�a�$b��B+��-�N`�\}�a��=Z�.ɳ�;�w��ȵ�b��A��\�O϶����?�o�항,�
 �֑[PG�M,�+���3vV�o�s�����s%�.����m�/�I?�W��P�i@�uRt�h��4���b��m��挫<O����P��}�\=�*նN/�]i�X�J�g����k�����A��#VR;���P��� ��Qk�x|0b'K�x�?��K���q8˶���v�D{�o�65�y��Z�0�aS���'�:+�i��IgKZM*7ߩ��hZ@��Č6^�q�ǧG%�U���%!g���D�t�f�dL���~*I5O,9G��� +�&0�6F��i�$���9�	8��2�;��/�Z��h�,u8�l ��S%�l���5�!�^����]����^�W��ٛ��
��R٪�Ӝ7�����TƷ?ILh���M�\@�!��ĕk2YZ�:̸nOo�W�ŅѿԘQ�q�f�T��߰�!hB��\{6?8��g����[]��f��Lry��a�?��0�}H�#�&8�.��
f�X��^+�-��o��q��D7x�w=(�F��9�H����0��Mj�!H��~��ɦ� ���#�cO��c&���o�,eD���:̮	B<���A��
�X$�-=<���ʂ��.)�\�QK�|�[0�N�a���<(��O�?d�ONٶ=Pdy�?�E	�����d�nY�OL��K"��t�]���|-�O�a�v�l�Y:����T+ͮ%�����)��'(���%.�Ǿ{�GN$�㉝� Hm����� �ڤ��ʶ�k\b�ܟ�u�M���A�j�	W��D�8��➚`�-�4�/C��m5:�76�g�9����~�R�m��OS*��Z���Bk26-H��C�����l�*; l��:h��+��~��w������I>C��<�&P�bxz@WЯF��(c����'����&
� ���U:�\���
x�2�����j�!j�A�ͧ�mx|���H6�j�gf[��MސWÄ5�u�]YĘ[ ?��E�[b$,\�f �F�bmI�"���1*�6���T��qv��.�T�7P�7o�r xaZ���;(_�A��ç�굝��KW*���Sٻ|��f��܏��	a����a �V�ڂ��`�jIJ6i�
���)P�H�����j\C�+���[c�]�􋹤�o*��$����l8d�05w��I&ȋ�������瑥*� ��R[���d!6�<W��pYY�Yc)���/�b����q�R��z�����f��,�(#���.�X�XmA� F@/���CW:t�~a�Qv�}	�H����z����\��|��L6�ɺ�-ʓ�_��p�HߵN#���~�:�nkz�s�e>&>(MI�!�� �ڰ��n�R��/�YAX<c`?+s-��b�q� M�k���:_ʲ-Y|}�K1������4+h?Mbۡ�R6Kٮ��O�������~� i����;�P��6ޝ�c���ovd�F�7{���A����NU�NN�eK�b7hs�It�z�vǳ��%�;�����?Pg�Ç�d���?��G�������[��n��>��)�d�ޅ�dJ]��EoA����/۱����1�䬩$t��
v�������&�4ʰ�w�]t�F�Kyh@��:Kb_����m������(��o���iC��[��g_a�o1ͩdA�������%�戉i~��]��'{��mgԗg����t���o(� �kG�}wv,��]�QH��sRgG2BL��j<Tb8*��ӂ�2?�XY9ʎ��@�p��T��N �ݔ�s��8��	�gpCf��AL̺�s�\��R�;�=K���g�irڛ/-=2f��hy���]�:؝�v�d�n����(�{�T����Jda��뱭4@�`#IPY@��@w Ge�Х����K����j��U1-�3ߌ�#}�a8"��7�U�����'.&��c�K�j�Tb�[�u���=�^0{tV�K��d���ylӲ��S�~L �ͩ���_��C)>�#�M֎]I^I1�e���^���Ag�$P����b�ڡZa��'�G��"8M?�(@��
�k����"�|��iv�е*�����C_�g�֩�a�/S|��������o>��U��e-��'H&��j��D��|�B���iwX#xo�1��[�Vv�1�1M�ܗ���|���o��Z㲿�Z��'�eC?a*Zbl�5��v	���U,%�$F;�?��w���������=)�d�}��$T�sC�����X;�(�ڲ��̞�q�sgq��
���s��2�l��*�L�nqx��(����1]H�[���?܅u>�}��G��&�ޓ����`����9Ge4�vGJ�[�%���)�z�5u�% �*�_�ǘ 6ƻOŧNe��1,��&Ղ���<b�]����~ӗ*��/%=2("=�T��z#^��g��rrȔ�Ը�F�=�ӕ����5��}�=�cd?�D�� :�%�Ԧ�u�Xn�&�NN����� �K�{@���;tL�(�팡�W���2K��.����V���tV~ p��� r���>�6��V���AX�&�����5K�	{�(�������yw勂V��5<�-�o��^j �J�C	'����o����ll�dT<��ۛ���&ϵ��&g�èZ��0os�ֲ���N@`D�j7��Bz�S���g<O��0߀�j�2P�ۙ��}�܎�NhPU��%0F�fѕ`�7u{�pD�]9g-\q|�I���[�Q���@Щ�� ���K~}V6Nk�f?*sC�"�{�z��k��8vZ۫�����&���f��Q��k�h!FW���寂P|/�K%0��$��ex�E��=D�IY>R��_%<;c<LV�5�	�M1�G�g5��H�)Vːr>�a��[���ս����GC��3���{�Pfw6�S��&@����%X#�<���A	b
�`���v�+�v�����i��ޘc�o�`Qy��I-^d����>\[�_�tR��y�7_P�����S��˿��ԣ/�+��!�z}��!�� P8���$3��_��Oky��g'��g��5�Oz��9�ӥk�o�υs���#K^��Ŝ���FZ<�?}&kǻ(1n
,_���>�����O���R����w����g���S��z��
��{����Y��t��@�� 18����nee,�\�υ�f���&�L�T�6>_1����O�[j���/�}g�����  [rj��>yP�����E��{�#��K��k��eX�Zsb%�m^�?���f<|s}��?ߺfݓ��:��,~�"�J��LKJb�c�\�#P˺�즢� ܳ�n��X8^Qa/o�!Ůqz�
�,P��#���k�U���\�ϳ�t�OM�׮9ĭM����vm�L3�r������wyퟓ�7�����;u��S�m��q&�hkt� ��3vya��EY��w�1w�M?s���FZ@�M�� :��n���@�r�=��a�Ъx�d�"��)�
�}���T#mg�D�e)|W�P_�$%4ܮ�[�o��4����	ؚx�?��h�局� �@���ZttrF]��$����fl�=�)v�4B��A��f����}̏0�$-����2H���f��hZa���a�@ܷ�hby;��})�����7�G��nV#�nQƕ�{IL�{�������;5� {8�{c�s�cҖ�z�9W���n`�q�쨛�����^��7���J0�f��*f+�G^/��&&�-P��K�����i��h�v�{# '�i�m��X"�c�Ė�A�D8.�	���|�.�fķ.\��w~n�uF��� 1�g�~�q������n���d�B+���)`k�T��c����'3e��o�e?�}��율�/b��R1lEꄼ�_�;�/1�C�wn�ׇ��m������h��	eMꨳU 3p7n��Jv������乎}� Y����XjbOၘ �V����:$B����LwϾ���������,9ܚ�δ�J2����y¯��m��w���k�v�� �v�]aݦF�����M���/Gw~�	�>V�k���k<�l��P̣~O�$�G�a���g�۳l�Ap�9 `�	,PP�iN[��"Czqu~��D���1�g�'�S�X�9Qd7��韈v��l>���uogH�xd�|����cs��������Й����%@�,B,�^��=k+�#��\�G��3��N6�J?[b���.:�Ѳ��`�T��-�y:��t����Pt����R��66�d8=+2Y�f�
��Nl����pz~�Ύ�ƻ`��~�����@����:ʙ���`K������!��t�y|P������l�{*� ���i����j�j>ԁr>����g�C�
��W,��f� '6	ӧ3�3bD��Y0�gh��V����Ѝ[��{`�G�.%^Ax���fUK'T+�-c�8SƁ�`���(�;�~n�#ۗ�I<�DCU;{����r�^�xe�h{�S��j�6Øe3";��_$dK�$U|i�j7��alԚ֜�h�p��zR5��K��KVf[�u8�;�GiA�r�Mm`�8����X(٢��?�t[�u���5����vb����e�>tym蔡�  ����ͤ�{�5/�}%l�ra�3������y�zh%�k�P^�.����<K�W&~�>~� �9\�Ӂ�� �2�ǒ�uX?�Sܓ���S;���ɼ��]��d[Xt�ų`����=6�S8�w��ğ#!
����媰M���Uch�?���׿�5|��B�6ݳ����;�*��ߚ�ݮ�zI�X6~j59B��i�u�!f�1t���(�\���U�-6M������V6��X�-�cY�y)��ƁT/=������1��Z�����b���16N�7��+�����!U߭e�ٖc�Ij���"0i��CČ�k@O(܍g�x�)I����7��1��|Mv���_�T}Eג�\(-@�4�\#&Zy;��5��q��P�}/yU�C5+P.l���I��4I��El-�i;#�;�4�s�����N�PX�!�ksM�(��K�u޼�R�)h�� �!�4\/�jQ*=Y�L����y���3*�kb�����1�҉d�ӽ%���?����w�[�Þ��!j"��V�)�L|��]L7p� �%���؂�E	!�~>�u���x�vq��d]��;�'B2����+���Ҥ�m�j�Lk�x�N��J���M/	{��k����UI,�Rُb���֥�2��Q��N�q����y��G+��B���Ѻ�%�H����e ]��N*��2Y@}��?�2䄏\��p�b��D�P�\�@՜��,�z�Gx���V:ǐ�m%�ZBߕ��a1OE�n���ձzc�w�Ӗ�*���8�=�4ϡZ��&��M���XnHc����ÁB��ΧR�EKǿ$6�8 �U+j.lo��v�v㖾�}0C���{tB�q���H���㡷�#N�= L�ٮ��r�t��'X�b�M&�!��]�\���Gċ�I
b�{ι@M�%&�XW+X�.U��4�Uג��V�(��ځ8vo%�@C1f�>��� K�S�Oc�����r<H6�#�����T���yz؄��;��b0V^��E�����-;�D�\^Y�^��NR����5�>kr�i~ F�h�GR�M$}(UH�I/t�0i5�S�:W:w��J���:[�ɰ��ϵ�D{��_+�,���g��XVO�A��Q�|p\�JE�%���n*:W�]��C9���)˯���?�M�o���[�=B�{�o������7i�RO�	2�bbʱC�^����1MV_���װ�呾������4�(���x�v�|���/����$���5�^�Rڲ��� ��p p�LR[N}�����'����b�Zu���.S!�{6O66f�e���fˠ �ݸv#u$���m�V�GЦ��1�GL!����|��k�a��� S��p�)x P��+�A���5���Ё`8�d�鬀%fم���i���8v����:��{�9:>#�L��O�l�����AG`Ewu2[���s����p]��C6XK֋_�ӳ������F	YS��@J��%Nh�ݛ^�Z^�+'TNLg�j\��3�,;���#�i������x-�����E7��E+ɠ�?i갆=� ��T�kXi��O袾�a?��"4��?_�p���%K8��>�]@�>��(�K��)A:$p$���s��:31�-�gJ�@����@Mv7[@3a�~o�*��L�:�Z��w�V�H�+��D
x��_o���� xpzzNN�XW}}��_���ZN�<rL�}I��$��T6�
"\n����cA{oJ^��-�Sq�������|G�?$ |��aI�:87�:�}=�ɜb�s�^�?��튥}D'38��4cx/���T�WI�؀MQ�V�8�H(���%`"����Q�����PtN�p!��Sd����:�.~��1���O촅�߼{�."ԨAf+)����1�k�I�{�9Cx�=����M�-r
�>#H�0�be��NK�n/	&0j�8{	S;��]��=���\4���I��,a[�3�%s;�"3�Sp�@�����(�ԯ��?9XY։��vK$�9�I΁<;?�ᗵlaH�B�Ɠ5�䟍�4~��,�t&�7/��n��6&x9,�P���fc�a�EO��񖬼�,���S����W����b��<Vr�ۙ��`ϩ��h>���f�L0L�����B����`AgT�Dɯ9����8S�>����:z(%???e �NY�mx��_�?��!d��6�'@�
�Հ�첕�N�}L�Ь�:��T�d	��1����Ĳ�E��V�)˓��K�����Z�2g�~�}ɲ��S�E��a��\;��Q�w��U�ո*�E����3�Y��옝�pL
�o����7O<�ζA�l����י�A�[t~�C�4t!�qO�2}�D鳴*%_`:9&�%�b{+�ҥH�K�'+��)�dIG A3Ť�^��0�dU+%�RYI!E�S���9	�V[�V�O%�^T��"������5��R�)9k2��%,�Q�ؽ����N $@T0��N��5n${�>��L�X�_<�<8���ڜJS�B0p��+�����ʢ��M��/狕���o�o\��c%��� C��u��}za�a)�2���p��� /������pc � 2d�3����-�����S�?�\|���I0��8��cwP�Y���X���K8����L�n�#;Nud� I�1��>�Ogv�Bb��9�2VR�`�0Ǎ����GӐCy8ħG5�A-���i+�C�NR���<�}�=�� �C�J/^���b�<��Mڂ��� �}��g�_��l�G,>�EtP�t.l,5��}(v#��5F�7dQ��.�����5=s^}4~I�Q6�ε|3�"�W��;8�g����N����&�>�(�����1c�� nV7�ٴ)�^�y޿{/�����h���O?����mߡ�%��q?X�1���O�8N�r-�Q��`AL�g�V�pSU��]n?��?c�4�'Z�T�MH%0�Q���{\7�����Ur�Q���Jd��I���8c%t՘�b0�:����<��jƩN�f*��-�3*�V�W��XP��� �g��,Z?cӉF�F��\�ki]�����Od�d����e����~?�����P憚-��ٽ���c���q=��'Y5�#���o��$���[ם�!8�?{GhCP�қ�rM���j.�Q��&��ZgV�L����$�]���1��g��iꝜ�d��*�=��)�%��
#��5/�B�Qk��SOt�Cp�~0�*X�!�Mgz��?��׬r�$�e���Iٱ=;V� vY
�:z
G�<6�]��}�ne��	�Ǝ)s��ߖe1�1Z]/AzC��C�Ɔ���w B�d���Ԟ���&cG��nfq�q6�������7�f��==�N��>	�[o��
�qƎk.4>Q<���v[�w�p@����H4,�Q�c.x0���S��h���H0d tPfaN>�f2��i�L�����*b�P��Θp�&N�N"�E۬�$N��E��V�:*�4;Sr*)Φ�>�t�ǽ�bW �,��w���O����?�)|Eg+�����[��=V�Rw/�8�<���u㠎��4K8%���p�v�<f+�0�[֭/�I!힝���ݍyߕX�n/�{2���&��^_��]v��/�����6ۿ��ۀ�7��t��4���z��^ ��>]�d���|���=���gye\�������ܑ)7-����𓾿�i�^M��-��k��3&��ă�͸/'�vf�OKIr�~i�Eg�������:�I7p,8uFI�yr���|��o0{���=�n`���@;�������:*7I��@���e�Cd�è�t*J�^�T]#��I��='{:��piR��|Z�s+kE>����L��o�{d?�������Qj������d	4|��μ%�@]� o7Pv�������Nk ' ���l��S�(�!�F�\�/MI�s�gt������3lM�	b�[t>�eG�	�E!��c���ƽuګ�'�ӓ����쨿�S�d���[k�}cGy��4�`nJ��3M�Ƣ������Oz�@�\G���	��l� �Ӯ�3�`�ٱ�~�'�\�%����canw�'j��X�?�W������d�����^��S���~ДI��=���ہ�j����.�\$U���L�R�*�U��{. �D��ک�;�<��cOh�M��S`l�l�Ѿ���6�u�~|�2��7״'HР�H,�Qځ �lx[zd1��.����%����~~��\��c��NMj��ʲ \����ʱ��⟺��$}{G<2p�CI6���0Br�w"��iW��VV�.=!��]��v�,\�ۉ`͍�$f���x�g��*4��Ω97�
��;�e��!'5���#�?e;�e9}1��F
%@}�Ǘ���R�+ ��FL����E	�
8T�Mm��9�.�(�
�q�ni�hDt!:	%o(z�m+t���O����\}�I.a�E����n���(��Ϧ��ڪ����1��9�Ӂg1Y�'2k,��oNK��Xdv��-L�{���cb\���@=+�Էдb��QFq�B���B����hc�;��g?�9��'�ގ�˥���g������13^Ȝ!�c��':~�l99��>�Z'N��ՖL-�?xX倘5�g#�� 7FctZ�k�p#��e'֋/XQR�}�FY7h���{��]$?i�{�ko�;f���҅��n���93)j��ষ���E*$���Se�.�ކ�6[�O%X2�N�;�//�fyn��UJ���~�1L��u>��6�](})<��E1�����$�}��F±�hi��%�,��:[/4r�De�ܠ6�Ƴt0J�te~�&��ݓ��4��m6hM�Ǜm�"�+��vV�R�ln�p,��F.�IO��7�_7�v�Xa��A����}]1�b�X�x��4�j�#^��u`�ۘ���6�r�ct����X��?���;���Gt����P���}Y�b����_�B'e�����V�́�yP;��Rf�C��;5��褌��)�eZ�T˒ )��MeI�V�N��AJ���;vv�S_���^Lm�n�`���{�:yd;|�n��f��T뻇{� ��2���<���y.Y}|�j�
��P �"6#���W�lӎ�,wP\�c�������n�ِ	���':9��y����}���(G�3��K��W��F�0�ɇ������Es����Y$��3���ژ�gO�K�o�a�P>��ơ�[y��SA6R�!�؅!�AY4pg����x�n�j)�{Ä�Ȥ��"��C���k՟"�"�v�' .�i,���:1BO���O]e�ՠ��c=	�"��@���$5.`&;�3t���,:�jxw�5?o�^i3�fh���tu��g���E��u��v�#˩�}a��ݢ�W�K���-{�[ߩtH���ʹ�N� �J�c$���wb����-��K`��ڢ_�����d��dV3�e�D�a�k��Q%�,mξБ:.I��ub-�ԇ
�Y�PJ�J�0�c�V +��ґӂ�d��SIlh ��� ��,YYV)��O�k$rl��*	|Ds9:�鬐�� �-΄X���'�qq��B�g�>[�N��+���T�J'D�'�bˇ����Qu�ܓ��F���t~l�����7���T]c�}�.���4�s�=���ϓQ�x� N���ة����s<���s�R�cZ�t +��T�AY+t�a���=YKw���5~N>Gb�����βw~zF�gaZy����r�E��c=�Gd���{��]��d�����ط�`�P��]����2��֎T�Y����K�7@7�|���������CX�L����̣�l�m���]��>���c��~đـg�1�G��й`v�l�l3~?  Z�3�ɶZ:�9��{�0��
2?-��(ǑG���L�k�q�� ز8�eL̐�n�L�	C�d�l`Ƕ�(�H�����P+ �ĸ�R�朁�/���xN��㊅w���Y����K�!�Mm��t���g�Q���"�.��a��x��"z��R�d�Y�'�Y^o޼e�������񗿆�~�)|���Y��QZ�"Z���m�����l=�g%�Hd��Q~>�:�+�M��
�f!�˓�D� =ɣCsH-�عj�k�� �ixd,x]ra�A�X�)&i����Rn@������/.�� ��4�BW`C7{��P�k�I_����/���!d�1�`v>����	���/�� ���\@����XY��y�1�+e���a�F+�`t�7���\.�n~��2�vf��;Q(�bf,��H~b��<[�����}OyS8�q��1��F�Z��<Y�)j�?1Ӄ������E�$�4�B'�
���فz|\������Y7�&T�Z�z(���d춢������ѩ
��v|}�N#{�&! ��N���+�	�d�V��p���;��>8$�w �Ľ'M:�;! �%�|On�Ã4T�;��8(�,��Q4z}��� 4�g��w��u.w��u�9�����wdRe�t�|�&�b���	e�l���➝��q�{|9N�.��A�@Q�~�`5�Oc�ҳ7���90�
P�~�����8�M��5��WK�� X�����z�S��DP/���̭]���6N�1�{\�ʞ�I;XɅ��T�\�΂IC���Ea��l'��.�@������M{�o;> ���uK�Jj'+5�� �>���5���þ
��4� D.��9��HyOPZ�~t1��j���hui�zp���-H���G��?U�sP�p����~m%XI�OjO�m��|�|�����`.���=��~�:����GA\^���xH��>=Ib6��ű�2(�'�O�(���V}���/t���	|`YU {2Q�yI�I?�����SW��+��n��F�2� ��'
��OF�ֆ�	��Y&N���Ym�:Z���ɺ�&o%(0�p ƺSv�q�d���o*��̒��1��%lCl�{�����l�,��	�옸��铉:�_��}H`Q��V�2�vV��7�4K�QFޡ<큠5�/Mߣ��}�K.�~�����5��η���Ň���>�e�����=�����-ԓ�b�$X��-�ucU�0[�v%̶v׸�����X��nib�}F8Q��q� �ܳ�k�8㫰v�酏��]�m��b��^���p���h}�v���\�!%�Z*�NUX�����DI�����%��v��:{W@; Ǯ�͎��߯o���᭬���B���+���ղ�VAX�%a��аy�}Sk�=>��^:2�����y�I�ٮ���}�k�6�J��/���(D�q�پ(�Ě�wW��ws���N�`�`�Aɦ�;,�d���FLT�(��xb�F I�4�Q��/�Y������"\e�	%]�w��1يw�HS
D�&Y�f���16��68%�Ԫ�6�%\;���뵄���� >���6��!Q2��|/�~�7uO�n��Ť+
�2b���c�M[ŊZ��L>m�7��:c�dG� ����S��`�`R����mv��?�Rp���͘V�NPPG���rTyu���8$z���&3�!���~�+��.���<A~����/���_����vNM|+��
E�;��wzSY�"��m�n�RL���v�	l���U�づ�;��!���X]}�"ڌ�a)�s���*�܁6��Ѩ�h�H 
N�arP��I:�S'M2�໊[��"�������X)#��3 9*�Pӱu�89=#P��I8(P�Slh3�8�'d� �?:�Άg
wwt�`\��߱9g�3�7g ����A���� �#��X�a�a���s�F+c��6jc�8����Z�L�6��mb�9R�hF=+�>��@V,;:��@�4�h�<�iK�N��f����]\&��\��ĸ�����O,���;Ӿ>�A��h4�����	$~����$�D�� ½�@�7����S~��uM'��J诠noX��Q��D���.�����b�-m�(�@Z `T��u�*�	�����ݸ�	�.r��$�0vV�î�%f�ZLU��s�e-G�S��4���L�t^�w��w]$�09��5�5����U�w�����u��.?y�߲6�9ı�Sc���,��%��������:�o"���9�s����&����o�`G%*�R�����v���u�B�^Sg��g���!�pD���v��iӝ��-P�YZ��{��'b@ubw	�+�s��S��؂Z;t����.� ��lr���^�k�\4�>^��V�n#�.e
��I��{���̕� ��H�\=�٪�FY$����zo��Ɗ���:��O����5��?��b�z���t^��ɚ�H�g�X䵯�Ϯ�_�ձz��*y=T��������jN���y�r*& �z�}���9�=��K��\��:*Fc�)�l L�-��`M�`��9���΀H��x|�ry�}t��5����"�:kN��Ǿ�����d�����:peB�Eۥ3�)�Ġ��^�&�ֱ����ZJ���EMl��h]�5l����7SK����#����gä�<��W�qʛlL�TJ�T~�Pp�I$~��/9x���ZDvQB�f��ׇ7�@�&0I\E��m@"#*pJ�=9{*�?J�1�مkP��з���:�u=X%}q
�Sl�������B���9�m�$�����-�Ĉ�jW��l���O��n�U6��� v�t̒�� v~W��͹�h�J^��e�51�Q]Qi�cmD�wl�F�b_��~;[59��}6�~�},ړ���5�j�{�i�%���3D��!��~�y
F��v�M&c����[5��8�vv��sh�,BI��<��_�����`�s!x9No�<}�����1�5�aXϋf��`�P���0+F��E���\^RV�4ۊ#��A�<$J�n86 7#9�i�}��|��|��Ev�X�� �T��@�
������>�ܺ7`v��Bl��3�vi@�Nu ��jw�dc��8X���7����n�&������p��7|yت͞����-�'ť�����)۲���o>�㟤�?��O��������)2VC|ǒ8�ͻ1|��n}�~1��S�y�b�%a�	�#`��ue�r��ꇼE����jD��%ډz8��+?g����F�|-������� :t��q@�Pfo�V���`SzU����j��,�EQ�}����=�ۢ�5&���/���,�z���F��n�pR�����. �կ�A��0g�=S�A0d�^p^�Y��(CS��� 9��9�Rl%!,C��6�v^K6jFB_�{�Ivƅa>b�@�8)P&f%`z��E�x��;F�Қ6���8����0�v�j�]�Z�$2Gv���=J��ίةaO��-���iA������|`a@���q�1��]q2��yNVK��n����ܻ�������?��������:ӆ�H4K8�`���
ݏ�zu9a|�&�#�� `��w�$aق��N/G�Se��S�d��h���C��X�R�f�}��n%����,���:�w6}d�VG�il�Rg�⠴S�D޾v*��)5A���1[�b���0.��ɂ��,�u��L��l���VU���,Y{���8'w<�Acŧ��/Z-ŋ2uz�
�A7�d+-%��`��!��*(I����(ݠ'n�jm9�����gb���*	�ԉ��Q�m*˲ھ���%c����lH9���s^�ccIuљs��<�T?�6NNs4��]:��ϵKLh�,���b����˯���u��fn ���v`}�M6j��a6v���� �]�]74��\���Z��r��񘣕$��Nq��wV�d�g��y Sk�����S'��$��F��{���۝��b+�G��)JJ=�l���Y��;b��?ybh<����k�����k_����3��7��M�p.s�y�Z����<`i�������Y���W{��o�������Rg�4�dzX�U2O�s%�$4��h@�Jg�`�|21Eߥ�>:��7����*�t���yQ�)5�5<w������E&�w4{���o�5����R�
�z���s��X2���|E�l;��0l 5|��8�%6��+��������|"Hv�@M	�/�B�Q�4�\���{�������Ob5�^�\�OVr�&�E65l	J���cG���%%+v<�{ N`��D��y\����ȥE,b~�{�2q}]pg2 gn��P�"��~E����x����}I)�o���܍�7_���l��
�CP{�}lİd;�u~(���I�f2o���G0��R�~�2��1��I����R��ggcGc�ȉ���$ �'��������%ƽ�` d�{}/�woȬ�gL���h����������"���`R$u��נ-��ĢM�`�ڳ����3�1��v_��#�Lƛ;5�nш56�YA���5�L�W ����:O|ob'���8<m^�֘.�f���%�^��D�d18^�u;K�w ���4��wއ�>�wWo���mX�?�|��IO?�(�W��Q)��IQ�"o8	��6N� $D�q��6Hl��o�*��6PӖ��]H�
`�kFB7���a�td��)S�)������M���?��c���%/P��Z�I�gj~��R�C�U�����&�d�m_�<�� ��i�S~% �d�����s6�������hN�F�]@��0vΜBm�L����=0Gd"���_>}"�s�o,)e��0x��XN�;𓪀t;n�ů��c�޿5��+�|���VO��䂛R��Щ��~�b�',x5�o�@��ͨ���Fr�e�0�{�`���S�pֳ�)��Ǻ��\�oz]�~�ދ]�MOd�=�̨�(����:X}~� 1=�	�#R��
V��Oe�'6����=��p*��3�s�j��>x{t	�i^��|ޅ��5�	�NO���9Pg�!�K�Mό�hG�[2�� �lkO X;OO訵c�3��b�scI��>�?�ϟ��ɴ��@v0X`Y�wXS��o��X-��札�^�h�p����D���-Ez���Y����>^���X@]P]s�s+��^��a�NQ�p���,Z��۾ DґI��3t����.�v�ݴX�t�Ҙ-�Q�R�u�CG��` F[Oɑ� [�R�^����_�Ѥ��Y�~I_JY������(�i߂���[�&_�$�z�q��gW�)�����H�ޅ��,�}�q�A�����_{�>b�!â�L4�.�5�~N�e�Z������:��`)�֞�D(%sVzs���Z��K�o��1�i�0ϲ�UX>�Rq�[�,�<@���_Ǻ���`�
H��x�L��Ӏ5��7���6I\�4�^b?��#@m�A�l�sr�si� �A��z~���k�-C?�^f���15<[m��Q��:c�и`k�%�ꊑ\@�&�ٻʅ�%��%��Q���ɨ|i���!���:Ǽ<�ߟ�%�|i6�mj����J��z_+ݷ��>��3����P�t���I�\�
��&?c��r�ζx?����<�&
ġ���}�ug��0��;S�@ƀJ=�l�D��S�BJ+�R�nz|�p�SS[lǃ�����J̱�N��~������M�6kWM"�#�0�*lc���i*�ʃy�g%�|=كd�ȳ�>���jo��+c=�RJ>Z�.&� ���cGꍨ�:@ڣ(�R��z��
6�xtzz����F�d�W����K_-1k����A�����&�lv�Y�P�&BW���k��m�G��hX7N�8CP'υi���KT5�L�FX� ��� ��۸̮�#���n���C�����1j��VB�y�����(U�k�#r=����K�'QY�i�$i�8��:��Ʋ��KP�@���I�%��D�,8gOX����y~�6��Q���7|N��i��i��4iI����<� m^����Q����Bq|���B���[;G+���7`'9 b:Qs�9S>b��B*	�4��6�F|p��P  ��;�dՀ�@��I~	�l���˅�p�3	jG�y N�Ϩa�Ï?��1��������Ż(c]��|�~)J��?����>�J�}��l���D�������~�k>��S�S����u
O�v�ܦ��������<|?
P�������}��I,�e��r[d�,Q6�XG�Y$op䮀:i7r����m�/�rjq;����Ʌ��B3�aEt�bS�>�<����L�hA��[Wh�T����=
'����4	|�#h���<�&����x���Ƅ�p��U6�G*�ʐ=hۖ��'y�8W\YK�x�X�ߵ�	��2�<�5��V�ڻP��H�f�x�u8`4vD��T��A�f�K��[^j{���gN�껅�ъ��'nh� �;��8O�v_������z������� ٙ>���.�z���R��J�"�0��j^ ˸q<zm^ɯ�oxD�CX(�������qn[�wNt�І��a���k~�S^��&���|o]:�c���`<�u��q�v}ѵF�NP���Ke���\ta���(���Ε`�`��	�Η<�e$`dQ{�~Xө� � ��?�&X� �@t�pAl9�=a�!��5;w���ޮY��p�f[o�������Y-�]5�>ea��)	f��o����#�ۿ��5#�w^"��Tz��8a��Mj�+gPŧ��8j��7��_o���b��bM��~83�m���K·�,%4��ݏ��H���E	�w��+�O8�O�6�&7,��S��R��4�TJ�fAC����/�uQA0�,��w�yݘ�x��Q���| �qu�N�W�1J�\�Iqڼ���<�� ��������;�z2Ր��M���Wj}�k�سP@@�B�1x�V�Jw�|��ؔ~�YWy�o됽���Ľj4���w:�$ ��/��]/�3S�dg*8��(�L�v_�e% ]�Y�+E�ab���p�+��|O���NEܲ2�\����}��d�Z`����,|���a��Ͷ8�S��6۾�lV�J����`�@R�V��Q�]��<gR��&�i�ݩ]�^��{E�110� 2��裡����%�TW�� [�����<קd]����mօW���z���QXh����]�}W�;�-���>i"V
����S2vUdI�!��ɳ��[������=<�
l��Jp�R_�%5�T�C��wPg�^�,�����Ʈ�� �&E��b�-�#�1}H$KT��l�%�u��P����,�脟�^	K���f7�$�������zB�G��~�\��v�Ű�>ߨR�R})#RRn��:I�kf}��}|q����[]��ec��de�A��d��"�;1i����ZN�)�~�^&��{o��q�H@7��S�8G�s ĉ��D��:�x��d�Ԟ6d���'�:�(����2�K s�"�8M1��x-�+G�	����?z�}T�@�2c�w�ݟ^�:B�y�*'W�cE6Ղ�������(63@�T(w��NF��!��P�Q�`��:>�$�����Q)m�Y꽕��		�qة�X4�7�!Β�P����k�@��	�K�K�xr��ƦIb���ь�K��㼤\����M=�CO���|�Z$&�<���  w�d^���h�� fPg^���VT?<��=����T]�����;����_�c	����R�}�R�`M�l{X�{<�|OA,�˿��u�c���&z��qwǵ���$q!1����i�{�:N�ر���`$	�%.�c�a�������j�䶒m�F|O���:�||��'1�}��]@��$|����?�!|x���)��䋛���X���w�7���͗���Z��<�N��Bu)�q`cҐz��;�4���Ο��>ކ��C�L�|�m�f���(������<��U�آ�U���2�<� �]����Y��j��.��ϳ@��n޳E:H��ɒ�a.먳R;?��%ʭٌ� ���M){s݋�Y�JS�����J��C�o#�M0p���|����l���R��^OFNkv=�p��|ȃu�'.�w��H��:����	���nk_��2��A��F�iV0 Ò�`ǧ� \(��i�D��iT��BOc�r��HS}.��qU�7�kf��AY���@Y�%�f�i8x�gF&���=
�y��66�;3U�V�a�(����w���:!�Z�=������/l��R	 c�T�I� d�й	�<@�������C�����%�2K9�2$_Y�p� ��w��nM*$�킮�EH�����D����ތ���@�zsW���^�Vk��ՔV��ư�<ۅ���b��N��Ztz�6���P�7,3��
6��,�ݯn����ҙM�	�q��ڿ�{�c�j���W�{�H��,��
��c��Y��� e_��`���t�7�O��]�,�	���~��p���J��R���;Z3T�9jx�Z��0���Z�G;���~�@��}�O�* p�D�f\u���١�2��9iڋ�����D��D��uo�Ό=��?��{�����ݣe8�
�����r>|�}��>�m�ּ�N  ���[
%c��䝞B[�����������?��ݪ3���,�׹��/L_�v��|8U۟]�gm ���0��Y�J4�w���T{	۝g۬z�������(��������/&��RU�&��l�rBn�giIa��YzO�I��1���	�M	:��n=��=xȎ�Qa�tjH�g�q6����!���d��7
r�%����?�/77�1;~�u��Ćgk%.�T����b��O�T���~��I������n,��h :��l��R�f���z��
{ Pj�yic�*"���1	t��1t��������,�Rˊ_�0�?���߁�<q��M>��ן� gĜ�֑Lq�B�-�c[���B6{?���>��o�;ퟃ���	>�cY��k�]|8Yp��+Υ��V-��� pf�f{���1z�yN*�D%{%�������Ya�~SH�(�IZ�	� "�n� �=����w�&"���n7�Ϝ�oX|�(�ή���߯r�c0&���Y�����҆Q���l��|04��hc%VR�뻆 :�Ã�W���a| T�ȁ��*eA�$�����n�S��mlR�UM{3�]�eD�-��Z�5����zo������$�����cq�m�`{�q��\�$ �B ܙFj��l"��-��Y�	�D=�����rf\
�`e�1�s�d�4KNN�	�`<w�{hW��"�t��l�X#1T��=��#�Vh� C:~���g���a%1� � D��J�w���mF��`�����c!���R$̛u�� �T�K�op�6�د=������}/��_� Z20k�$�w�\X���B�%ƈ�$@G3������ki��%�?�ߗ�o��%Ŧj}�X���L������Q5���f&P���C�*Wa�Cڶ��U����X���Ǐ�����?��O/�i�B�Lt�at�BS$�1�p��|�n�\�M^`��My�)��Ǝ�_���}?�6kv`}����uy�}���]���11���~��C_�_��Y2��.�y�.����������)�����׏��ۙ {�Y�#`��xp������������NX��|��<����=����z��}��������Ï��@�Z����{��_
?}�~�z�$Ŕ���;��G%f�T�}Q��m�	�#����j�%W�`P*��Ç���[���}������?��?�S��?��%�h��������}�ވE��\��D,��ns`S,Y�.��~7lN�Ԗ=8!�C�d���^3f釦���"JG�v|AEl�z
1��t'��K�Dnk�A�R~P�߽{KE�ӳ�t~|�7��AX>�z֣E�-Ͼ� m�Lc�ȟ�J��ZQ3�eB���$��3L���&U�;�rF��ʢd�bբ S���X��������\ ��\����_�������c=��;	�d�";ٹ7���8@ќs������(?�)O5�+�������B8��/�����av�]�G�QH.�jnή(�s0�l�u�3���dN���D�����q.�V�[�дfO�ظ��_\�6l��\��ư_l��it1圊k�i��&d�g�kN���|�C�91���Φ8����f��wI�8Y&ca͑)��,���{�e%tt]k''��û �'@�����Ɗ��4*7���ZJ;x��t��Xj��U����k��8/R�ҩ�[u��=����<�¹'uy0�m���_��Mv���d9��-�9�Б�n:GhkZ�]{ �t.�6��DY������q�v_]�̓��y���+;���[���ue҆��t:O)�����E���;0)��˯nU?׀�u�,Q���2��Po�,��������N�Yp6U�@�`�N]RN~g�}���W����`2���l)�[k ��
Wy��:��}�ӧ���6�n*�����Cc�'h&�3�e��!� GJ}M�h@�Bv�v���k��M���ɀՁ �n��}i�j�B*4qwv�������R^��ig��,��
�š�' �t��}� ���k����Z(C(e�6�پ3�ln@��m+����}�ubVb|}����/�V�a*O~����	�D~UMV�3��D��g����9N�Z�7�y� ఑p�֗���湲Z1��ws󕚊X�m��9�y���Na����K:�\��c��,x���4s?1��)�����u��2�9i,��Z�!ܞ������ݓʞ�;�u�t�ق������ނ�5��H򭍥�{l��Y�<��½:g�3�!�Ef���	�oHDqt�����C�D�2& � ����U�$�<�|�߭!>� �
A���g���1Q�$����c����j�ൕ�-,�����4���M�/X+�>��{����-!a�T��  y��(3ԙ��7���4�>L�,��,x��!震	"��-��} �^���{<m���O�wU[�Ɗ��nr ���l�R�����Y"���'������,�4�����$NUև�q��u�%6�WS����փUV��U(�MY��������a�s���2�R�[�'��ߋԛ�_�I���Ƥ5������ͭ|���@_Px��93�Q���T%va�\*1jYzk� ��;q��@cRŪQ\����It��p�i"����Y:��>�H������/���C��6�a�@M2^6�@�8+��B:�y�'�w���<���E͎VǔǘF	I?����6<��6�[���]R<���}��U8>;�Wo�<�/�ݯ�� ;�'�c�����Ix{v��g�8��gW�b?�u${��^ z�P�C����2=#���R<������>LxN�Itr��HBD��1�gO.���U�ȃ|~zf{���3Qϼh��`��R*�lS�/$�U��"&2'��K�����	��|�`?���](�7��*{a)H/��73��1H̃|�<
�.�0 A����X *���ɺ([�7�g���k]��P��>�朕.A�=��k�֯#;�~ĺQ��~uc���_=��o����B��W��������s�7�|kQ�J�M൧
��(cqBg��xt��LJ�݇�|L��L�[8/Kzq�1�|��W�����~�b�,��?|s}�����h�ns��!�������]�O���5�_R�����X&}�Z>ki4��^���SNm��ن� ��Ǡ��B���)��`�M�0�W�Q	o���eVB���r��i�|��Q( �� ;N�sJ�]'vz1�M`P�~}$xC��h��c�h,���<om�,�YX��N��;�|���߅� 2(�y��t� �9o�`��?�W���eX���l���Cb���'����d��0�k~�}���'�7Bg��8�9г�Gt��L$�GӃ��Uou�S[�d%^�Hb��p(؃�d F_.E`��L��听�gW�Ή�b���������v�� ��ꧽJ�d���'f,�L�V��]6R��kߗ@�%S&��Ln00:X{�D�7t,��!�b#������S1%�X����
>@��0�$�:���e��98�C��~g%���6Gv��=���/����~�E�<�>�P:��g��t]�Х�����啞�n���N,n	������o�"M &[n��<Q�ŉv0Ƨl���ܓm�e�7  7� �j��+��P6H?:u��	������i-�E�B�ۗrdɽ���^"R��}��5H�;q_0S�3���{�K�~0?X���&���~�Ze�ç��g�����!�3f�̧~�Rq <�-�r���v(������(�|ژx���>�d���VF�c�Ei���N;�c�ܧ�y�m��%�Dv��]%h�Q �p�K�&c4F}���})W�L�[�N�fD��Fa��	��z�?���y��j�P��I�@̩XXI�1����Z�/Tf�X��}��q4V���Vr8#e����Ҽ����L`$ĩg2Π��"8Oz΅��ˎ�U�#���/Z�s�?�o;&�v����d؄{�X�	&,��i0��X=!�l;`����-�f5�庪�UZ�[&%�ӥ�|�&��+ Y��\^:���ْK͛St�1��/u������&aW��o��O`<9=�R�'2�>g-��L�a�2ܥt�4g��R��]�vYk�iT22H�]d	��)��&$B���F�!�����r��*�p���N$ۇ J��\�/��E�i~Ͽ�뿆������*����,�r�Y���
�:
��V�L;@tO�k�$�o���	X�'���۞��ur��~�K>�)~l��ٽ`���<��Wy-��<ʫv�6e{���?�wa����tRޛ����s�.��eb$ 9�GE]��+�ہ�lM��$TXB���o�5pG��m=>����;/��Y@�,�ŁM���,�'u|r޾�ޜ�o.ކ#Կ�ƪ�E�����]p�ء8֜?'�뀶�0�A��"��E�iQ�}���P����T�A���?=�&�N��eC�����C��|�cR�h��z�wm������^U8ԤPl��_u{�8`���<��m��~i4@����/�W�� �=�,���w��g�;��s���YG�3:蒌^�W���ӳs(ca[�6*%%��I&ЬԆı4)§Ϯ��9\j���w(A�ab��&�1ܩ9�����-�{63��A�P% ����__/'�� �
�Ng�h9�'�h�r��P�T�ּ5���#�hm����E��Sm����M��5�����èYGu��6H�R0�B���b	��1e#G�L0�(�gR��ioz0�^���pL�����A
�����٬i�p,�%��x����Z�X�-�Ӏ�Lh���p�@��K
�́;�u/�Z�ct�[�o�͜��k�lb/?tp.��=�6�j�!�����Ky����}y��Ҥ��b<�g��.\k�~Z�(�����H�s
��/"� ��bUJ��?	I8b�V����\�N���RvXԵ*X�f�d��Q���%g�(�@��9l=r�'��8?B+��oɾ�l��4[�+�Z,��Y�(��3�b�쭤��S�\�~����ߊ��$��4��k�%�8ۮ/`.�1$��>֙qs�s����_�}�5��αeS��Z���;����:&�������ۣ���׬@9��&+Bsީ�.�+A��Q*���=Of����{��,?K�-�M�r�2����`��=���Z
-ۜ��e���U3�}PBVmW�ڙ?&���?"� ����#�0�8�tNL�.��LX�C�x~V2Iؙ����쬤63.��������cټiY��͵����i�KGH �{�9���Xy�JAG+i���'�f��B��#��-`zo��q,��lu�\���D�V�Zʋ|i���ymZ���s�v'�q�<��Y:z@f�,s\�Rc3F%\�K�KYNW�Of������6f��p����w���.�ʼ�����H٦��H`���G�1�1?�~�6�pxp_��c;i�/u�ݍ3�aСb'�I݁��t�*�D,�����0_H��$��l�i���Dҙ�7�|?Ć/lo�QS�� Y��\B�UU��?c��o�������j��J¤�]
�ڥ}��lœw3K��'�[�,� �ڞ J�S/�8��ӎ)�GK+U�|e�(����b�S�����T�uօV�Ǐy0� Q��Q����K����MX��r�~��1\��P���[�OC���8��u���c��%Ⱗ��hR��H��Л����
oN��Y�;'&�����>���6���6c����&"�w������Ex��-u��u��H'd�@�:l`�A�fX�|7̄Q���;
�4ևc�\���n/��(�#^�(;Ű��s�e͡�}�.<C(s��㡗h˿�]s��eu?!�>Z���1��|�^���-�͖%왵Cд
�BJ���.~�M?K'f��]	�fT5����ة��B���&��$'�@׏��������9���o&�	դ<�,���x��t]���TW������3�#�B�eCm��_�dh�v�_����Gwx�t0��I{~�� ���|�o�ָ&�!���M����g=�ᗿ�oH˱y��ˏ�Cj\'+;�3��U�j�#�_[UϦB�������6�)�8ۯ������y96����X�����"��
��fko9eǣ�9h��]i&6+����A�bס�YI��ZM�k�G�%�^���
vok��;/��7A��gQ˻�ښ� ��E+}�8-J��V��`��ҙ���Z�:�@�ug B����@�;�rѦ�da�a���F����I�������9�B�f�����h]T<��6�9��Cn�-��K���	�Z����8ߗ�-�T���h�_����*h;�W��#XP��\���s��V�K,l.][g��t�R�M~���6܃1��F�m�r�F�:�b�y_�y���7G��uQ���';����_���]v��>q����;
���	Ka��ߑIk��Ɨ���,VT��^^o T�����Y3��6����F�'k�W��&;i�yuj�M<�R>3���%��O&(	V���}�Yk�����P{#���:>%��_}��4L��Yv�vߎ^J���ͩ�V���z����!�(�N��~�}���sah�d����:�������e�m6V��#��n���T+{�,ϸ��� �z7�4���Dc�J����le@�cw&���NKB��3��ϴ7WЁ0gf��Θ���r����%
������}��ns�r-m�;>�Vh�{dZ�UȽ:%��	�I��{�����[YG��x�j;DwK4��G�i{)�m»*S�ʻ��Q�f�G@.�r�5Ɲ����Х߹���m*�	p���+��9?���yh�+XG�yr��`¨u�$�]�^�H�B1�8������ֽLI5�P�N�$��a��V v�c���֚\]wf�f��<	�c�[��Ǯڎ��*��Z��%c���Z���H[g��\tf;��o�G'���I|�<?���$�k�^s��=�[�~�W�@Pd�ޥ����:���#R,�ߴ����ŗ��碋��F�XL�># ӟ5�F��/�� 7r��$T6�%�<�b�c>Rw��$|��C��8�NvJ����EZyj)��	��ͩt�s� D�E�o��(A��P:2�Ce�ؐʷ�Q]3Z�	��篟�۷��J��GU��N��Ey>��:CO^�3�NC |���m���y�ߜ^�����*ϥ#2�N7����,=���$R�^6�{� ݯ�@?�8ϱ��|��+b(a}�_��
�#t/�|E��J`�~��e�Eo�:u-C<ξ[<a�-�h9g�?]|��6�l��+��B�v�8(4���;�g>���1��՛7�����Oh �F8]{Qfq�P5�h]�9ɘ++yqv�z9�P���&�g�2 c�jX���s^�V7����эw*(��
�M����UY>�0�A=�<WOW ���{���$[42��vٮ��Mϼy�����3�]�mm��ȗ'�Lp�eWu���D�@"�Ȉ'���zz�H�T&��o�V	��;VPNC:��j���0��p�/�>9~�ÿ����A�����$�Іp����DG�N���@o���4�J���v��3�"Wϵhʋ{�x�t/��>��V�ٕ�#m��N���n�6��T)��c[>r6�����ct�R"��T�g&U`,<4�`2N"9E�t�w���?�yq�-_Qrn��@�YK���jwC	j����4�=U}(�/e
����2X���%
��A���8g��+h���/����&f��RSϩjwn�R��ɽά����s�Z G�6�����s�*7�/�6;z�/����~�̼=���X�����m�?ê1�ѭ�(x�n�Y�r�=���S�J�&F�s��@M���()LI�U@dm�12�.8���H0��I�q/�}'s�G�5�'�X1Y��~�fX1uQ*xuY��c��9;ͳRu"/���(֧�G��h�+)!l�6��  ���:W	���Wd�!�P\���{�U��t�����JR��<�$$ȃ�����9��Px��y�s�@�����7��cJk:��|1��V�?�G����P�_�XD���m��Z�M�~%髃-��|?#E]����R-�V��#YDO��|��|�B���RG�TO�{k�?����"B�ݸ�ʴ!��pK�'KSKAɌk'LQz9����eOS��ʮF��J��Ԫ{១<� ��V=��a� )'�zXH��A�8��R����\�F�8�Iڕw�ӃD�X��G:(ئo3���0(�9�x\��� ���{8�㈡Œe^ �P>iY���� Չ�/�%��2��a�i^f�ʑ���DVM ʂ����1�XG�^
W �����k�*��|�wǜ�M���F����-�4��
HH�Y�+�*�\�&� ̺*tu��Q&� ���|��|�t�	W�����Cj��!�?���Ʉ>������������;I%��$�	�^��L4=u��AM�f��T���A���V���cn����xxD�*�=�#��#:����#L#�lA��0 �$҃��q�_0�AT��Q��H4 g���/)��`aI5H'RZQ��_�j�Ҟ�>�������ў���㙛�ʖA �[�����X��F

�j��j�܊�8,zț�;��G�4��V�m�^9 �d����©�-@�$�S�ՆS���v��U�� W����q��o�nhu����Δ�2p��}w{�:8w��J�3Q���.z�9�l�N+vTmD�Q~Q��M�H�#s���b�0�� H2�Q�����} ��x�!���/�FHs�d�%���"n<�y��������Ǹ��'�ꌤ![Ll,0v� �����8�?�W�W�"A�[F%����]�]���5���I����;9��!�:!��=Bc5/^~_ꇋϘ���>�x���\h��5�Ώ�ҁ����H��=�Tu��������'&��PX'(����<�~?[G:V��1^�vP�t>�7���k0�����[��@Ǟ��a�C6��Y�L=6"\�x��C���5bQK����'	�#ԝ`���;C����j������뭉���@T�Q	UB4��Uti�Y�?��H��$3N�xf%�n`�2#M8eiwIӔ$$99�W~r����v��/QCSƹCZ�$l��	E�"�C���p�Ϥa��x�'J�ۊ�5>?J9Ԭh���2��=�8�T�8Z���jT�r0����=ܯ]�0���j�����ak� <����4o��i�%l�`?��=ڔ=(�g&�%���Q�l����do�����.���z���j�,c�XE3�k�4�aE�+pr�H�B�2�T�)r�ݒ�6��d��Ĵ�fE{���Ѱ����MY[A�0�~�
^��錫fH�U*2O��m�j��\�'+Y k�"Cx߽{ǥץ�d���+�O?�>?�ДIa�;_���UU�$rF�A����w�C������G1(�kF>+�������ZyC�l<PB��te��P�^Y��<����Nۀ{%��q5rrV�K���q%2�W H��Y�׀�Xtx��5F�%��d�W	�v�㘜�?k�THw2��Z�fz/��3eA�{�D��~��j�Mv�&�'c�{G3h�`���BY`���>�Y꺎E����N��"�s�DZ�Be�*;����?M;�g�x�h"�w�tW�C,�}�lZ�M4�+%���s�F�XI6���zG]�����qZ3�W6θjP3a'AqJ���Ș�R#2vͰ�B0T왴��e��9`.T�bl%��u.��T�߲]�����������^K����_�@XT*
i{��ْ��q�̉-����NRڙ+�QJ`�ɺ�Y6h�۞�S�պPͮ��;�
�8z��A
h��؋v���P��)W C�)7d)Xa-��]��\Z)�t��n���p�;iPR�Bn���o�z�DA�@9���H[���Ӵ%�Z�φM��0�Z�V*~%o�o;��U2��$�Sz�gy���Ǒ9�TK�r�H[��E��9͑8K�;���:��;)qp���m��E��n�TV�%3���8��W���u�s�9���l��020�זPKunm�(Ց�<�*s�v�6i��mCg�^xնY���@�ՊA�u�{���K~�Ǡ�!����-mn��:���X/�j��{�!b�A{����9�iD�_���oX/�����A��A��8��2�;��U����sjN���@e%�W��w b�#p5p�+X�/�̋���_~���雙�[�d����	�Q�����k:sZvk�_>�ǇO���D�/��<�{n�9�Iۓ#@m�#K����8w�c��M/%h{#�̋��3M�V�p�N7e#�e+��Rdػ�F �aG��8
o8��h�ݘ���mM��C�E]�U?�M4�;'�Syycu�T�ܒ:#�� ��G��뜆%�-��x.b�OK���^c7���{{����O��������@��a�,Sp��<v��4��|. eW�[��+^ߺx��U�R��!o�<�o�p6��>�Q9�,�C�!�)�Ed�����G����8+�Pcu�[}���M�p�A�Eb�ά
n�c"d�%7Z��zT�j�Jʃ�IV1ԫ�t�k&����?L�x��R�<2�<�ޟY�����>q����� ���(���Q�P�?���۾`o����T��ӵ\ϕr_�s�z�;,]G�1)y��p1w�9�� �< �� �����+��)�)KAʰIJp4 B�͗�����U엃���l]�.�J�!���c�^����,/��+�@Ij�dc �1�^=UZ�+��1pU²�ko�b�%���#\A��k�8&�X$~T�@��/��Q�#W��>�����Ӗ,�¹��>����9�kA�7(0�@��(�,�N�U��+�9�o�VLVLO&�N�#��dސ�<w���y���l�9��:�\�kmR�d��D��Q��L����Y*[఑��q�PP/�<x1�>`�n���b\�pAz��#�:��R٥0W#"�LJnP[ʯ��=�z��B@/��:�#[_��>��x?r�yD�f�,;J�"�S����D�M}is�Z��"y�F���>a\���l�T`�K�F��ы	0�R�0ʑ��	�]��"�X�6�G���2��7��� ٳ�O�ka����ksU��8�40NsC�+(��r)vFl8�E�9�TG4h��*�� ��,_7�ew۬��Ge�T`aU�X�1S"l$I\��"��pR���������a���S	T��|M6U�����}���M�R�{o�NI�ۧ���5�ܒD\��#�Ӛ� P���9�|�����K�3��TK�N٩�̕N����m>��Q`'�`n��~��_w�����\L�&�Dc�@�$ED����.�b��X�z�H����dn�Z�]���<rK�#�Ǫ�ҭ��?{̶s�h:'���2'.�Z��	R�%�g���q6Bgp��y�2b mr�\�ߡW����6&\1�7�8�@��Pf$��L�ȻN�)����?���vE�'���o|M ���EֻV,YzW��T듧�s���}T�'Tn#�<:D�%�P�M����+�!M�,�/�(�4�����[m���"�׭T4}����)�+h�j)u�%�o0���V�򌀝���|�}#P�&z7bx��I�%�<&���=}��7����_��w�0�;�":D^�=���/+^p�״��B]n����j��[<<Ȥ�2y�ł���j6�bR^=N��$p.��<��M��(һV��.��$�v���?��rq��y�M>HOϑ@b8�2F*!��4ݐ�)�s�z�\�R�B5!ҩ�f�:���i���Uݘ*�ޞ=�Q��qp��:W=1�b�o�B\R�ȕ�D����V�U��?
ǀ�+�b��MR<�T��c�:�hWF�M#}�T�eu��=��.@���U�/Tߕ0N�(�ZUjke������_ �a�yP���(4�y9eN鳺RoZ}Y9rF��Q�'���l�D�\��ۨqX�U@C�1;�;K��Iڒq&��_��u��54j0��"�.�85Ҥ�����r�R�<(�3�S�Ť�F�5MC'�+d%�-�&fy=�����n���[�r���D�������Y#�jp����V��������2^ף�����5��̧�D�Z�xuM�0e[?���á�A�W_7I�����B�1��ݚ�ĥBqZ�=zg	8j4߲g+�p�m�}�h@���,��6!��0��@J���KA�+@��J���c2������߁�g�`�F�88�L�c�Ijvl<�*&���Y�:������_���?�y�H^��A`T��tJ��CyT����5��#���E�t�i���U��*�ج<�}5���ʘA�I�<*?����N
��Ы����͜��`�����ñ(2C@��4�hH�#}����+���B*~#�zi��vG�U�04�]����/ě۠{����`����6�ʸ�j/�&Ϙ/H�X%F �d}�j`��}�9�ߓh���1��R��I��r�#t-QB�����Ye��_�^tpyF)�BY$�r�d������A(�^4 �z��[�E��:��3T<9��Ƣ�jt��*cA�Q�s�u�a�NA��!5��JȌ�a]���u�0%�Jǅ��^�*'5N�F�ɐ
ǔ�>�T�WD#����F�
 �n��'m��K�^�َ����Y�et�w�~��s��N���qFdȒyr�xF���k��jm�l;�|B�D5����^F�-r_�r�\�3 c!�/�R��D[���:�H��g:��wC_$u�[vb�Ⱥ���h+��۶�!b����;����=;Axo���	 e���3����BҒ���:��)?d�9Y��;�y�p��0|��LR�d��;p�Q/J�� I�:�Q���@D��Ϥ��[/.��8o��тk.$����6<&H��)Y;��Y9*���Bw���Hg�ԯ��N��To8���#���,�Z��"R��8;;v:��1�y���+���e%�Z�O�6����HJ��1?�s�/ H�:?@U���8&�kǖ�O��jr�#�(��ьRiU�6�+{��b[��cS��#"���(��bA�%_�C�C��3��
�;¯��c�O�c��x����J2�o{I��Z^+�Ze )P�k_����}�ƓR�~W��:��e)�CΤ�y�=~����#��ϴDe�4�����Y��
l����p����[�0������Q[�A��a^D�<"�488R�{�P}Ȁ��sTƜW���^���n�Q��~��Hd���7��W
��8�V��p���@���ʐ~�(m0o��X�z�������M���]�Q����J�O�2��t	X
Q�ʦ8�(J�N}9&	�PP���)�֚�3���<I�l��)X�T���^y<H #���"Ug&Uf���QJ�{���x��!�7�@Ւ^` �r�0��g4�W&Ui���T$��11eh9:�VA0U<��u�޳�z�c{�L[����8>_��T���be���o5U�D�T�rY���=��`Uh�zSP�N���2G��[�\;�$|?�����;W1p��:�w��4��.���I���Dj�Z���0�ħ`!��8'��d(�)WM/����(�T�
Lh*�RbZ+XɁ2�F��	�Hc��y�gX�Q��!���P���?&�����Get��{�����T���k߽��t�����u^�$~fo��|��S;N�Q�I�vTK��A9��~z�4:� �@�S*��jމ�WI@�� ƸtWz�FKx����7�>�����1Fo_I�*���s�	(�{�=�<�U��5��|�H��9Oce�U�@�t�
	q*{�����14��ɯ}�$}.��(�����z��cf�ݠ������{�ϜK_�*������0�Qc����c:��{� sH���P��)G+HP�{6%t6�O�H#}&��݁���k8�5�������1�L��|��G��.�-�D�y?Yr��r���3��*�\�R�����I�3p
��W!���f����k$��I�+����2W���+�C����@��6��$���K
�p�� N�E�Z�fo � N�^��F�dΞ��3Iݓ����quu�k`��0l(������W�@$�y	9���[T<����W�tӣJ��J�\;\��GgqM�2��o�E��Q�,V��ϵ*�FU�eX ?��⑦�	#Ӈ���ld� �.�V�T��fY�M�D �AE���9G�4��ϦgtsyE���s$>�K*zK*�T7$�%ۻ�9��_�B��`���@����%]�_�{]pŭ��[��0���Ź��C�c�6��#vt^��z�(2,`�Rf����4�Uf�F�U�I��F��-x9L��K.50؃Y��}o���署�W(#:b�0�njZkH�1�0ф#�j�R*�*�L%�Ba.��}T�2O��&�y�(sx'��B�q?yycvJ�I	��d#4���pV|�񕗭m�d^���k��`)LQ�,l�N(ۿP�^���EpQ�
p*���:�y8�C[�A�D��.�~,d=Ug��x�|uɷv��Q��Wvo;t)�N���wZ�n�+��8�$��͡�5a)="��i����B�j2�͕]�r�)YyS%QN� ���]D�YAs�ŠX���Z�#*�l��K������(B5�Yb\-hqe�¿`�O>�m]_4p�"�~m����]�%O��bl'S�O��@��Ƃ��QF�����y�q��wG�b��'���T�)��<0�oo������_����g%>��|؉Z�L��)MEc�IˆS�0o[PBPv����s:��_df:���c�!� �tC'�К��p$LGDe��5����Pd����BҰg���.	1-W�w-��� )'�������l�JŔ�M
	`GRh��q��n'�Z�KR���}�N���;�P��Uӑ}B�\H%��������+��#��?��ف�������tL����0Y�G��{�Α��R�r�M4/��*A�boѠV}s����3�;0�A��Mv�T���%���R� %/i��;�zj�P@[�E�늬���$���#�I�����L�,p^�*M��  ��IDAT��=�k	�O2�ϪuG�F�j��� *��Fr�y��%F��1����9\�73W;ѢVm�{�=+����@�d������U{Q�:����*��l���DoD��{~ԝ�3]���H~�=�W���IzM�g�|�,��~K5�e��,%�^��1w�l�o���h�gRb�ޣ��V���d=0�P����YmUl��"��[�f����c�R��VnJT�:�˼mf�����o���P���3(`�*��_�Z9�l�j	td��e��61 a�#W�j�IH���ET���+����H�N�\�wD�</��|���Ĥ}���.}Ñ�I����DZ�}>�#��k��(Cs�.��R�Us����r!�>��sj�&�4BDy=-�R��˴o9�8��M�Dչ揚�/����S� ��U�3�N�� ��}��>�h�s���`.,������J�\�W� �1�����ib��L�f�u�J^�����%�e�^�w7w��-�??r��a������y��_ O���C��B*��p�/���K.���^c9#���NJ�h��ԅ�x~�{.����ES���,�d!!��I��$����\�lE�F�%NjU�<�3Y.픟s��҂A(�M8cg;�PEV�䐪���B��3����M�=��c��Z�}|�ѕ܃�y��Z�]�ea�^�v�~ݤ��|f��]��M�i*�ٽ��U�<c:r��H����p���?9�{n�Th����|��u^�)�d���=+��*��m<b*?��`�I��V����P�kаy��ȕ+���U�����4R�XTm�n1TG�3i^�)�z]��M�P�g%Q��݁#�ī8��*B^�o��F��ʃ!�d��H���Q�����h	�������%�ę ��D#�S"<���D���R�*C�~3�d�Ċ��2��4u��wu�����VRR�\��×b�"xU�ua� ��z�,T[s8dp�*c4��%�r:�l[NM���\�`��8V��#?{�h2A>����\�*3�p �7\?���)g�;��4Z-Q�ef-co6�p��j��|��R�ܙNك�pi�����$����~�?���@{^U��ҝ�3}�U�P�A�0d��~���AE���V��`	�V��oJ%��0	 a�N#����P�I��-�5�d�����F�\�?cq(�D��E�#w	���&\�kc�ҫR)`�;g׽�PT��#�,�,w��lyViJ�P�Ocmx
����d��kT��XsZ:,A%���&��l_��T���?X�J�2�(����?[��9|�����:�CVQ��?��ճP(��Χ�p!�([s~�s�6�b�*�]ܻ�=��U���GV˾�QL�������̤`̸��O�� d���ojd��:
��I������[�--_�u&��h+�y� �u���/d��F����ʺ�T�>b�������
��-]9�&Q#��F^U�e~�H ?F�wZ�*Q��"P���c��!M�K�#r��x���^�
���ȑ18�$ɇ�0�Fx�l>����V�Z0����9�����*ڟh%�N��Dx8+f���iA,L8\��$��A�jc�D�i��1�v	�xy]�#�����j�b�����)~A$���;������w?H��]��9wW7tuqũV�c�C>�%Jɣ(�(�1�Þ�L~<���"*9v���B���o��:�f�%/�U;�x�v���0���~^޺i�:����g�������t,�*{J	�Z&��#�2����ȝrv~A�ٙ�+I��Ԍ��$CRҋ8�	e՘�e�w�\���^��Mt�N.T�/��b
���C1�;�ù�yl�`��o/s;4G�܌�+�hhW5r��-� �[D��&�sr�}}�yM�>�������0� ���.�
jğ�{�\�[y�n�!�F��Εr�ʓ��Jl�����J[1T)u�����{���ұO���/,/��8��[#��L���M�G�N=�^�#e�t�N
T��<�Q�*erx��5�`'�:�]�`oHij�N�,���0�9��\�A�lZ�D��S����m�c��0b0WetK���â=���zu�0VT딝`$�(S	���N��a$C��wZ=}�襹5DW��w�fU��U���Kض),��5d䊦М:x,�����W��/�k���j���#�W��5��(4�k�A�d�e3�
��י�Z9f`g� U0�{H'�A�?c�/m#�w���Z�J��rĎ��N=�Ρ�ݑg��?����6W� �%����j1������AHW+���S��)��7��?���#uB�ɢ��Q�[�}�b�%5�m�������Td)UJ|n\�vX��7����6$�%��z)��h���ǘ�	��5�2*2.*w��Z��Unq>�^�{�闩���r"d(}ˌ`MK�_��JWk�n�!d�MnT�'��T���x;���y�� ��,Ըg�P���qYTA/e�-�~�W�0+�͡P�/c1�5����h��W����o[��T���>3����T�[�����h�J�7'��np�?�o�
j���ᨬ(��d@F�d��Wz�-�����kz���u�0�ʥ)����{����	��jK�7�{�j�����Rm-��*ں��C���m��os�K"��g�h6�9�@ƅ�t&|o��T���kt�T�«�K��:&�WD����Z7��m�����&!�t!�ea�׊�أ9F���e�����M���]�:1�+pP���؜N��X&�����m���V������g'խ/on�?I�j�4�(���y5������g뽗�k��;@GPNQpH��n� ;����?����_��&81v5����KD�A�]�������8�<>>�O�ݼ��̣܏��Aԟ������f����|=�up�]^v�@c��WQ*��Tbؗ����#vl�'[���9n�=�rC]|Q��/��.+i�����.�����M��u�q96���cd�5k8|�J�C�rb�*O�ʝ#�{�Z0�-�wǉ��S��2syD+��?��+��繳M�M�����Y� p&L�3���"��>��a@f�:���T�H��8���m�cp���c�&��m��$��rΉ?}�Ѝ���緑�$-ݧ�D*tR��<��<��`�&��m_9/��#�S�G��֊J}�~v`�o�G��Ł5�]~��Q��*-i�['�Ѹ~����&��J ��ǈ,��r�J�I���Ai�'��ѕF~/�A�h@�����T��DR�� ��7 
%����S!Е(��퐨�3'���o�R�jo��H0��ʚ���MJ�u]���ĕ|�q�h��=d��
Je�w�ե�S�wF��f������t}0룃閎�].9V=��Q��$8��%��kd'��V���\C�W�4'�1�j[�6������ u�����)J �DԽl�Z 0(3��� R�5����"5�Dv��Yb@To��
pz
K���mR��^�6Q���K��9�Zk�)cP<y�J��� ���s��)�!����//�*GV�:��A9��+���6��{�Cq���S*���ч���`A����>[@��C����=S�oRKT�#.�lժ$��3�ӲZ�'{�v^�M����}G�7�N�%[�{�4�"Z��EW���V�I��%�wV)7_8IڨJ{�ʵ�|���D3x�Pb���fp�WS�<��C_�$���pE�+���S1�+%7ȣ�T�Qj74�E*<�r������a�!�^�T����}�6:}�l;q�鑐�$|�a#��ԵW�#����W�l�pKߕS--W	�G:g
��F����ϡ���<Lʹ4$�K���ڗ{�"8,R�t�������3����y�9ה���&�ب=���*�2�y �AϷ��P�a8�S�Ü����z��QEQ��a�D*s��e�M��a`ʸ��S*k�YTg�8At��c�Η&N��68�>����;8�L1�s~;v�M'���!�������LEzְSOBIs5Y��B��������,i�I+w��k�`B���e���d��T�}?}������A��Ն�*�#�$j��9Zu��JlǺ�ѷ�ቔ���+N��Y�uk��a���D�'3�>d~@%A'�kp����|~��ۀR:$�N����C:�{�-���͚S���
J��1>:���H|5�.k���	k� O�^s�`\���GH.v�Z�����=�����.��Ya�`!<j誼���Y*BT���.WR=���`G��U Y�{A[���+���J�Z�,�+qp�)��u�QN<���+4�t���������u���٠�����PyY�ַ�oŢ0o���=��1�*b������� ������	gڿ����-�~�@-,�蝇D�
q�* %�hݔ�7�ߥ�뻧�2c����f��+�f9���}c#����Fg��Y�)b��^=��!����u)�C��p����| ��V#E�U��y����Tٮ��*tEI�_���L-�Nj�R�g�͞%~Y��E_�n>�Vr��y��� �R�-�x��q7����o������a�B��а�M�װ^.����zJ�0i+�ii2�l{M�Ya�)�.�|��A�#��U���������^VK����K����i����X��H��C��#�D�tv�9�I7)K�2���7J�����v��94g@yW��UbA�7c��2R�.*�E�*@��/&���8z�K�:3�u�%աȴo3+����|Y��\k�4e@�������� �/P`���>R�8�<_�@0���3T�l%����7���'_wǽ����䲏Fr���A���Y�_3e�����[�]�{}����e0���ےfa��:ƛ^�����#�9Y�m6�^�hu�����T��dࠕ~ء8n+#5�7��>�{��-~J>w-b�d��"gI+��fl��������ӑ�?1�a:q=�������.���i�@MU�8��J15�,�1#��>��w�m���F���^�(�
􊅿2�6�X��.]�ԡ����=�KZn�`�1t�.��4�j��>��q,�K�	�U�ջ^�uR��y�{>1J� ���L��%��~`Bp,{�̻�1�c%���DI���}Q�or�Z�WN�B�*���Ũ�:��Ӟ��(:�Ԯ�?P�+ݓ���"���:c�:�K��u�N_�7�N�t�!jT�ݠ:[��s���Gd� ������zG(���3~n9=I*Bq��(`��0�]�M�"�i,%[�N8�� ��Fm����&�R!OQ#�ߑAF�`�b�?�Zp ]�_���-�������?���d��I����ښ�8ͯ�ggp\e(��B�G#�C���YuW�<�6���]^^qֆ�K�A�}�Ϝ;U��V������������9Qn��ȜI��`DԈ%D�B�~��e����-VH�Zs�O[�B�*F�2m�j��Y����%�W��m�&\j"ZU���}���I�VY)C�5�s�Cï��K���B���c��7�� �A���O�,���]�tѦbt������E�[���va�8�() ��s1��Z(U�%�cd��J�mU�6����@"S��N�d��������sR0�?~��3�j�Oi�h"T� 8:#.Sa��YjBW*a���i�Ud�2&.���ذ�9�f�s	:�Lp�){�H���}��@Q�ңȁ�p+Zf��T�BV�"!��\s4E'��狚B�������g6��)�v,�v깗�����o<sP��Y ���2���An(t���ژ���B�8���M���R�@D�k-�r⾎q ��o��A�x��$� �Mɿ���Λ�V.�fe�Jڥ'i	�dD5�� d��=YT��[$)�U2"���?��d���6���e��8� ���V+}n����x�t'
�\Y��|!�B�n ����c�$�����9Q���$9kc��)��"�tؕ�0���o9J�|�� ��t��Fxd���A�xN0G&MI?K\9"�婔Tfe|�v'\p <`+�6�LTO�;�i%\����x�K�5��n�2��EΪ'{�z���4���|,4%\���@���Cr[����������I��s�<�(r�����q-{un+*�@	���k��y^������+A0!mnZ
��W���,+Gg��<��i62E�5B���C�;���;�{wG?���;KeݷI��85}���_r��s�+��xp���`؏���hq_ޕP�3�\ib�{��zHA$Uk�׺>S-{�9�������N՟��W��*)
��ġ��:�"8���e�����������"F�+����bT
�ɠ����,��&�����1!�K�l,�&*%�I��[�x�J?��[K�K�=j3�E��K���FN���K䄤�G-�N�{�;/W^Ҋ��U����82��6L(<��`͜ZQ�`3�ml���SWO>G�S��0�.��;v��*���iIӲ�=Fԛ\Cr/r��Ƈ��Z���j>��@1�!m��\-f��5�ezMT�X|M
�$�r~^�.�9M
����á���Q�p�%u=�7Q:q��N�K~E}V�@y�.��lo6bg6���N�G(�5�6J�t"��B��%}��a<�N�'����L��}?)5���FA?i<�*}��$�5�Żm���9�qݶ��`�KzY.9r�m��8A��"/9��)�LJ��������^˕)����H���m�&.D���8��.8���I�Q����C�;H��1;����-5�c�s���}��:-A�wssuKW�����5�4���7�׿��>��zZg�,2�^.��8�8�Ie���~KV(jQ��vM���j�B?��gr?�^6t{}M�~��ț�������ۀ�+�s���t��7���(�������gJy���m!=��15ۂ�ym�t�����ʘŨ��xy�:`�i�%��:O��j�`�b��<lM��~�̮��Bӽ�[ XP��Y�C�z.�+h;"j���2g��3����]�����ktP�J����ho��ؼ�TԆG�I�͏9"�1{�|�F�H�ٰ8x��jdBX��m6e�
��]�:�������"vB\3FMx�1i�µ�fx��eW<�z�#��6��*+}�w��#T!�i��K��Y6�B�$�6�d�b����
N0{����9�$g<ׄ�ˈ�x�Fb /6�^7D����Y��K�Hx�1�n�HF�F�/H������2(��<x!80G�%�Fa!�c��7Q���e�&/O�n�}�O%���zM��������u�So�j�i��j"���Q8���e0�T!��`-u���2΍V�:�,��ن�3!��"<BűWBD�ʦ�nC/�M��ț���V#CZ�F�������{#m5��X)[ؔr�6���K��l�e-��#�����cSd��UW��+r��p/[)!G�ʴ�5Yki��=*p��~�RU���dS}g�*���ltM%�UFX�ֺ^��?,J�\~�P�c'�ԑ��<wy����O��~s��ˢ'�����1'L�� 佶���]�����2�<��+>8�mk��u����&�;kW�3� DH�L����VA&ӌ�Ejg����A�����g%L���p�hIꐴ�K��|�r=i#Y|#s<`1�D�^\^Ї��sߡ����{�E��eH*�����X�g���H�>����n�d�Y��N8�g���x\��˖����Y�����/����Ͽ�r07̃ms�H8��Ǐ�v��o���j��w�t��k��g󢱔P���@`i9� �kА�/]nd�>BTu�F���H�g]��EmP��f��,{��Sj(t%�<Zdd�Ⱃ~,��|u�	��u� *�"d;R�-�S�*�y_�Ue#k[�Q�XC�7%�G⩤��G�D��-N$��8����釶��G��ؑ�h����psNX
DR�	�r�""t�6�u{�����7ޯV�6��"B�S�R��i���~z�E��90�#gݸf.=�����͈��:�}m.Xj�m��!�����Te���Ȣh���~���O����Pզ�����mt�{�>|PMoׂd��\���������G���"��UGѱJ� 6���G?��w��GR�S����rE�ņ�����C�WQ����T:�?�����
��R�~����c�EƏb�G�8YS%���a�5tn�L)���@���sn�n��Ġұ���+}����g�,	0d�\-��
�R�澓
Λl'����2���8��8��; �V���T	� ;���� ;?~�#���=.����?���̺Ҷ
��������;����+������a?M�9<qt�V3z8jgzF�W�t}yM�Wtu~)%��n�A���rE��C.'wX�E��2Yd)��]'��z�8F�M�M~������D�ҭv����_���8�N��0e����~����["�����߿�受�~]3?�O��|���~�ǧ�M�:˟����Xf�������������_9e�U ����C0`g�Y+U��ϗ��Q=��;���y��\&2�d^��a�=?�D �R�j���IǍ�:T���<���
��9sX��)�Үׄ�-U��29��8�
����?w�Ռ���԰f��!}uߔ��`�!O ϕ4`Ǆ��'�ߙ�m�l��,R���x%Z�k\�!a��s�%��BȆQ>��gJt`�7l��d2ER�� ŐtC��N�&j�۩n܍��B�,�����4���`e#�+��*ρ[�0���a�]����S:�y|t�x>i?��نd�dDp��
�  ���;�Y�v�?�4^�o6�ԛ6��ʂ��H����ν��GK�
 ��d�Nm�$�l�X�ʸ0e,��㍆�q���s�����d�@�Сj���A׸)�<#U�8�����;!0�&��pu�ZUJ��<+����{�x�<�I� 9���f�/�������� k/S��ɺt���Sa�5�S������ 5�=j\}�W����:P�F����jˇqk*�V�ýT7�Ʀ�5gH֫rш]�pd��%^C�Rļ>�m�2Ъ�t��_~N�t���+uDf��,3�����%o7�k��t(Q\9S=�=G:m��e�5L\S+�D�Rj�M-M����8���q�� ��I��#��@dD؇��r0�!}0^���c�XXo�r���r��B)4T��|AHR-��e��^��ՠ1��#pY��+_�M?4R����[���D�qT0H���2e��#5tJiv٣�y�}Y�^�֯�cU����cU��F"�c*���#�ї\^PWJ�k���n
yx-� M���M����6�hM��cDJ5�8S�8��20I���Tg�2���dN㷑�rj���j�j�m�ø6��hA0���j�L|`�])�+.��s�����Y�!�6�"~�J��g�������������K{���ux��/컊uh�
���r=���}������h���z}��̵q�pL���QO��e�����(D���Iq����񉞞9b�e�0ZKԋ��4�(�"3y	'`C�?�g@`��|ο/�^ |��������2�Ɍ.����|s�V�bi�u�}icôc����� �9��-���ێ�>=0�	y��� sn���ܶȮA�xpr+�..��?��zR��A
ST'x�;��,�f�.��y�D�Y�&q���H���.�㆝c�u��-^ty}I�{�QF�����g���#�s�]�Kg��2�Fi P��)���f=fr6���9ݡ�//9�c�����?o����]�����bޒJ�R%�^#O6�q\�Cɍj��dD\��D!d�NJ�B�e3s��T�&Ol|^�����]�Y0�k���B2����%�K��>S�������T�.��Z7ܭ_�N�^!�R��I0��5:������w��K&�j�=?�n��+�Xz�vP��j�O���f- ���XNvL�i�ӕ���p B�/���1,�D��)���?�"�
���0U�S4���5��VZd咀"��j� ����Q�����I�����v�����rOb�6rb�Ϋ��bhK:S/Q|�Dv0h(��� ;Ҿ�*��=� ��3(��%9�-sRH{$��߼�`hG
�e��7F�߉���<�.�p��+�\.�8����@�
�@T4d0ԕ[�F��b'�������k	���A&�{D/7��ګS���=z�*Ę^=�����F�?���NN��2c%e-ԘqQH�]��>�(M/�Ab;�ׁ�~��~���}b���F�Ü�������{�G����}E��۫�$��pF/~O�
�����6H
�n�ku2�No��`i8_��ZSœ(��@P����
m���J�z�b9�\�mV��gg��
�E���κ[sHs��܄���z �G"6O�TØ��m��o���K�?ਧpT�����>՚	;[��Wx���X��1]8K,�D<�,��5�<-D}R��H�i�q�cJ�;�ξ/Yp '-:Y�N��z�	X�1��0��?� ��d�S5��W,"̣���'��~��,�đ�n�革��Xj�~ڒ]�"Czdx���#8��GRV�7٬0�Fq8%q�U���K�H����9� Og�}LT���v��Q�@!�\��kj_���D�rT��5� �f�[���w��A�H x��+ht"���D���@��eҴ^_6e6���c��މ#���}� ����k6�K�S9����Z�H�j�]T��Poy��*�Sl?Y��*���89;h0B�����߽�M��?������I��e��}<�\�ʛ��m�G���,A0�����3��g ��v; ͶSN�@ST՚��Uޛo.�y���2�(�HR8�f��'pn��lN��}���K�|y����==~��_�O�����k�	׾����M���d]iLW���~����L�[1T�A��=D��[Zm^����������Q����88�s����^1�r�U�>?|����馿a��dp(2@4/�������cZ�9;?�t6D� �Ap�a�f��w-W��"IY2���	��j�ǁ��<//K�
f�پ#H��E�w���d�ț_eC3�n���|��f��wvX@V��I�J�]^]����^ϴZ,h�'7�W�����@���8�ӱ��?E�m��LY{�e��	�������P��/?S�?�X2	ƊL����DT�t/L�� �"7�56Y����)�T�(烆�2B�R�H��P�]�B�Ź�����U)#�Za.{עPd'ХQ�Y<�B&crW����h�ԅ�qc���dK�5�Kp��}�`�J�`��IW�r�۩�3��-�͓G�bk��$����{I�@H%@Ze���0�A<Y|/�w�3�a�psͥO��I#-�*tHʘs���	^��_��+$���e��pvZ�e�ZP�ׁ3S��I_�#�2����jjD��Pv)X�<P_w|�g��ӉO_S��&g	�/��K����+�����c_����"��T�اobryOI.N�"͈��p��J0�V��;�Pua� C���d�m�8&0�y}L5���5�L��V���d(X��Y~�D�oo��O�$r��k������FӂP�9I�Zy#Y�!�Ϥi$����NŘ��Q^RY��$c C�v�TU�?��
{���v|�;v�E��@v�[�(�Q8�Z��@��c��Qt�E�rJ��l��±��aF�9c�(�I�F�0���/�}E�P]`P���l�_�c���g�St/������%"O?s>�J��rԎ��?��%n�`�tCYg�0:����\����2�5UJ��*#>UQ�ھ
��R��!N��߳��]WC�Ϣ�Y53i�E���1��qC��+�oыe.X�k�U~�̪A�Y���u���Ӻ��@�pz���׆\�w�QV�}_�#XD�E����ˆ�<j�տ�o>��7E�H�%�CPP*N�c�T��}�7�MU�(��(i��� 8�U*��W�K�6R��;��6�V/d ��`(�K����4w�v �-�}�^]7����#�,���ț�8_H"m����u�9�;�~���_\��u>ܽ���[q����<�-g�L�������$՝T� *�'A3�z����-V��xO�Ϗ|	o��=��ފJ��_ýZ-��D!o�Ț�f"�7��I��|�$��d�f a� ��" EO����@��gnt�Ne��2,:�:���Rcմ�'�D��gr��L�%r���f�s���Y!;�J�>?���<i�i���ð��/�A� {%{{%����~���0>׈��P��ז/����2&��r�8�F\�=M|��P��/a��)w�K�Tѐnx	1�Ai����A��ʞxl@؄P��2���Z��Z�{���%�)��!�!���}+LA	�İ��8��K�4%O��t�{E��`{I�!M�RpǄd�T�>8��w�g<ʼHF�*�"�*I�nX�Hd�n<��:���Ԫ7%	�M�|}����2-@!!(5be�����@4O� �e|���l>#D��`Uǫ���lJ�2�Ԅ:N�O5���8ܯ�K5.�V��y�ȕT������f�h��)�������Yꝛ'j.?��pṃ-iu�Ns���b�ʺ���L�߲_��
J�oz�#�'?�#P��0e%�t����n={�Ԣ�U(���6@]�M�S���7V�ZT����?U����fR���b�6x���`Ͳ�1���]^��:�I�T�<};1vm]��Q�ӱ�v�����(�ܷ�W	0#�@��|O�� 爷�(�C��q%��o#/N�J�p�de
7>#!���걷9U�N(O�f��9Ǿ�i
�[�n��Q�M�D��go:��P��|��_9'��O�N]Gr�tR�b���d��ɸ�7v
z[,���6� �ī�gU댼݈�m-�}����5�a��5� CVѓ\'	
�XR�7>�$:�EY���'7�_�%Q���@�Z_���Z!Ƒ9�XQI�n�=g��F
.�m��B@���Q�->��ľW&�o�O,��#!R�v1h��o �oI����{I���� ��t!x$��p�$Uv�>��h�#���q�¢�FH�Ѫ��Z�0�}���x�@9��ѽ����".Nm-eA�0������}ز�'y��%�F���?���}�0�K h�AB����領��=v��\.�����Z�Z)S��Ȅ�|Gj4�~�����v�#H$~�{�����/.x}�j[0ip#D�6R���>�v˄�&p�{<˼��V؉��/��f[h������p6�?}�#�i}~|`�<;����;���dD	m;Y��u�I�w.sG��6��3�C��M�~L��
�Ö&O���J��QE]W(��$�@�s!E���9�x�( �앻G��b�:�d�P����լ(I�����K===�=���Z,���h?�����Y��!���|:���hj0�7[�Qd�0���E��+
�A��i��e�-p'L��ė4�I��HAy���;z���/O�,Ɏ�9���D��/�n����5W�]a����r��U@�U7|������1V�Ӯ��@�	���q�m5����H�$xvH0��_M'��U8bB	;i�w8���@B�4q>&�K�Ge%������H��ਙҎZ��"�XE[��S��ց(�P�{�>/��˂�Ո 1�F���D�D.��ժ�p��u�R��W��` U� ,�r7����HR� �)���U� U�l����3n^R�#��%湿�u`�4�)u��d��ٴ����@���Εm��g�!�s�ʁ��qŮ^�'H�Ib�52Na���9Y$����3�ƞ_�s_�v���F	'�,��� �.��Z�۸�t�J>0� /�GX�rh6d^L.��ގ��Ţ}����a��c���hJ.UJT�߷��Zn��~��/�M�qN�h�?$��R������P�
���on�=|�H�8�[��CR�P1�2��+�./k�x���y>o�{Ѐ�|��*xքV�+�N����� ?u6�'���j~��d��; E���7({�}� �*> ~2KiV9�lC���~m�*٪e�<�Zw�7�lW�o������S"v,���o1�H�����P�Ӿ:O�����9X	����>�?s�@~[�Sr�A=U[׌��[�"Dw���i=q�#l{Mц��V�n�X�8�O��]���(d�< 0Pa0�O�tL��N�h$�Zm�R��w饒S5��o
?+X!$��0p���gr@LҪU������qvù�O���E��iqNמ��KZ�W�JQ��B�\���8�TY��R�Y���>&�]�j*�:�%���(����3i$9��kF��T;�dv
�©����%W�����C	e���<]��%��A�:��|:�����^��Gx�ͯ�,�z�tDt��c�챉����U��
4IA�P�	�oʾ{�U�����Ac����N�d��!e�.��Y��"��+szU
�T����R��g\������v@)nτ`u]lb�Z�d�ˠs��N
!S!I�O<���rIO��i���ovt{yM�no����,[`XaPgζS>�ˈ��<�� ,�>��Ʃd�W0�f;h�^2p�_Kmږ�X�h�@+���͖�� x��ۈk޾�c��E�X�<F�}�x|9�n�:vH��j���5&��+Z�������\> v83��;���˟��oH�ҍ�&\���K'蠠q�)�l�W7 �7Y��N��+�
�J�V8s`�1���:y�`r^\����c-���'%$k��:{N�����D�iT����{P�>�n�j@%��DHE�����.dɣ�˙�T��K��o=��;!�� M&��c��PL�:��L��lQL�X��EX�P~H�Y�F��0a��&���&ĸ���0�O\�n[\N�ڿ�\�#�<?�B��J.(m���I�q���4������-R� su:��@���[�C��'�@V[��l5�Ta 2�1�s���\�D�e6��:!��*n�PocM�r? ؙ	y�T^���-C�)oQD�;�D�L�G� ��� �;0�o��(�c�!��_l�e,�G�t�h�T=�����0�s	�^�^��W;~���]^�s߯��zy^T�92��T#RcA��A+(Ax��|J�?�a��6��H� A�E�F2j���_k�����o�*,��g���:�2�^{��uojh���p��x��3{��cm;w�����
n�|�A}�������j�&۝�u������n::��-�dFl�Wku���=�U�ъ�xѰ�˳s&����t�υo�fs�e�9���&�S��bBֆL�M> �[�{Z�y&,$� ����i6���A� 6��i V(z�I�!�|Yr��&?�f`-#�������ʐ6ـ�"�s8�w�����)0R)ҩs�S?d��P"v�b�g�I��V7�U?cFmz����$�?�e͘�_Sf0�ɒ{U�n&�3'�`:�F�H��s�aO��h�NWPP����"5��I�D\I�RA����/�չW>2v�`��,�#��4��gK��Y镥�d5ʡ����4j��0H4�� ��$��Ea�
��2A�	g�L���BY�F;��N_7>>�%����-2*z{ ��#�DM�Wی�A��Q����Y�ǈܱԊ�̬��|���D Y4��S�9�Q�-<d�LZ���rJ3SImGZ^#���T'!)��p+%_���>��g����^?�,�V(�/~z�j6Xo�_��	N.TjT�MW7�d�8��.����7Iǖ�N��i<�쩇���%�N�z$/���C8�%��7w4�{/Ҵ,�@R�5"�,5o�F����i������w��R&9�2��&�'�R5�Wp�W'9�h%Y�@
��j����K��_V�������{�"����%���"����d9��H�-� ��a����MO��|o�&�.�gU
������p�?�g�l!\:��h�ME���u�շq�|/T�|Y�������_.�|o�Ise_�b�0�����mep�n���Gg��U�� v��j�B/��iXI�:K������2��~4bg���&�P!�k�Mn����;�l��\��Y�
���]޹�E� "��kCΠj�$��y6��]�r��)6�$�<<�^:���L7
��t��G�E%ȓ.4#�����)��0���pt��3�2A0�F���){�`f�d���x���p/蠜�(��i�@���%]^]	�_>}����KPQ���^�A��|F�77�Fb�B�4�|*�$��*��<�???�s_�$^��@A? Й3r�F?�K�7X8@5qM��v�\4��#u�z��C�8?t��ܫ,\��=�4tu��ڭ���F�<��D�+�	�:h�b1�%@�,t6더�5b��y+6+���"\�K����:��5�澑�0IC������)�A�$y�x. QS� X//�t�k�sY_bxN�fzt(f<&(o����U�`��}p��-��`qg#,?�w����e0���@��3-��\e*���7��<��H�ч���~��_�����}��=���no��y�̉������~'�g�SG"~�Q�9��l>���ܧW�-`�{:sr�U�y dļBi�^��̫i`e�x"�n`eM�<h�s�E,��޿�w k_���-����ٗ�����hdR߯व�#�X7���FJڋw�£'��*����֖��0C�id��(��g��ȲD���9<Xj������N�ʊ�zևj~�5��2�����G.p%%���b�(�h5�8\�yLg��؝RV\8�G#� �Z4�@��<�E y�ޭN
%�fC[ǈ� �$W%B��'�X�^a�]T�2�ې�)9o{�{��ޑ�B�J�^��Z�<M�L}4�u���O81���>������cm�Ğ�?43#���V%,�'6�����y�X���jT��������-n#���\l/�`��\@A�|vR����� Y?*3�<�sc�ը�jC��H��DT#���
�fŅ��^3�s������Ԁl���AS�-�9x��L�1�ޞ#�7�:,Tؿ'���ÀWz�2sJ9����\qV�Q�y�x�k��ˢ��u��� U�J�!X-EE�"�a��I1�B�귖��:t��v]�_]S�ht�.�R�4�Y@<�X_AD���,�X�����V��ﬔ:��	R�ǣ��X5�N(}��B.�Ua�����7��Yw�`�j\ �g������A.�!�@{�>@���P?@>�SF�%P�R��Gi$�F�>���~}o����s~���g��QG���.��	�o�\��5jU*�]����J�GUff�4By �!�Xt�5��*�%�P��&J�	�
+����=�PM'�mL��Jl��ēVlA
��1���:a���nq��:���TY�XH��^��e�A�'n��b�2R�)ۛ�~�(@���Ӵ`�������I^}�>C�"��N��4�)��<g�1�L�|� ���-G %��i'�ƏO�����跇����S�޳�����,2�@�#p�oz��AdѯZ%@������4ڏ��l;B�`��=Y����QOH�p�\�h����i�p�H��ú�{�)��=�4�U�s�f��KC�H���!N�Fkr���N)m�Y������i�tٞ���%mn�sø2�T؟�0j�����5��E�;6���e���'� �bL�V�I��t��Kt@�H�?J"r]�P��H[��(���B%F^�*�����Jvn����|�r�Ѡ�����f�I%�^Is��؋��<��xp�p����.�IA
�F��ȋ���.//U\��j�DH�D�\8q&�#���"�w1Yx�k(PWـ� &6�y��P��2s}'��XY� �dʑ:>����G�y�>�ٻ~��vLTk�|>�k�"�s�/�ؘ��_g�)<�-X�@?���*��"9�a����
U���������Y�g�z^,����G�(���\a-_g�r��kAh@H���Ղ�ϑV/=�Obb�F�4�I�_�Jwww,�'L��in��iyP(#P
�������m�L��%�I�}x�Q�ֽ����?��\<�s��� en�zw��>�v��-J���tg޽�
/�u��w��Z����\ [M��� K���,��S<X�k8�1������-ؤ��x����ޠQx��oo9^�$���S���|Sqvx��G�9��cJ���3x\;
�|3+Y�w�2��~O��R4�Q�x�ɏ?Ǟ#��,��J�xԀ��l$��(j���xI�Zî"y���X���V��};���T�s8I��AH�Yn�"�,z�/�� �CB�7(�-2VR(��㘹��gd羭	��
?��'�́��)HEȣu�٭� )	"�c}ow�&9�W��q�R5��{�TƳ��dڳ?�Σz=u��o	�=�S��3��{'�A57��K��a|���C$�J�"QF:�_��W-'%T��J����������-�nx�)%-��3��a�s��>Ds
�g��p�����=
rN��|�u��+�;"��D��� ��9�FO�¶R�6���e���C�+%#��w�a �(_�G
�da1���N�b���)8�vG	�R�u��{���>�3���z���zʓ���d�b]6{��r+d�!�}C���_cr�#��5�GR�Ԉ�4��4n��@��}b־S�d%�5Z'J�<�E'��S�:�8��$*(�&ē�@D�7��v��7v<7�Wx��K��ଂC/�lz������n�8GO�O+u�2B�D&�RJ^{`9�8�~�u� e�c���T�GR�S��a 'h����7�T��Y���F��_.������t�S��io�y���>�a�??%�+sn$�M'�Z��{Tt�ڙ_zɢ|Ib$vn����RR�`\e6( d�
 0�e}����t{s+$�Q�N�e��9�%G�d��ڬ8*��I�
�F�g���:��ؘ
n̺8tuDܟ�_�.ài�o�|��?�-�����ؙxz�7��� *f'��lsž�m�- J~�����/t����;��]T�ް���x�����O��G.u�K����Tt8�ʍ,�.1�[QFO��4m$g�h���A�ӯ���W�d��xV��|��^ �lWL��hT�B?sp�r�݊�W��k�k&�g}m�f��!�SenIr�)e�U��f{�S������2o~;j�V+wO�V�e����֨��#~�I��l�p!.�i��B[T��{��ü��U���=��A��/}��vOS��ۡ
�w���JBR����`�	}�
�	�R��qic���Id�,�[��L�5��T���)C�r���.�P@�Чq�iW�R%H1����?�I!�A�#��TK�&e)oy�J���9z�QC�Ɂ��>�t�N7`�2+>}���z��-D�l�h�T�S��@�͒�ohLH�
Dҿ�D�-���x6���͉�
�_q��%{�&�F�P1/Dȉ�=$�B�ً:5���)��e62���wL0.v���U0��7Y�\sڒ0��r� �����GF��N�'���ҌN�B�.W��nD!o���#ϊ>G�[ߝ�3 �T��vDUqj��r�o��Չ�	�(3)��}�1�0`�H ���A�5�7����A�=��Ζ��eԊ:��{�����h�B�!����/��r����?�8����h��
]Y�P��# �D��P��
hb0�#��"eJ�o\fD����Q;vs�R5!YZ�E�X,_�{&�x�-U�j �uG��Ҵ1]\��J���(FR�9�-����9o�y�'I�����-�$�BĜ2��
�@gQ�u��,0�(Y&a�$�N��W\B����_g9��J¬�Q���F5��B��t�79B�'"t��V:υ�>��?�H �A���F��հ�O�b$����j�gr#!�~��$�RE��"����&�^'�F8��g-~����Q��k�!*۸�1�A'�$����w�{������lv�-a�g�uɦDT0w]�O��z�����WK�1W�fer������0���3!��~>�OO�x^p*:@�9Jٞ_r28&_�_���-�β�s1�w�o�����I8��S
���c���g�M�$7�$A3 ~��y�����0�o����0{�y}T1�G\~�1Q5�==��I���_�����8��TEEE�|�:p��k�2$c'a��QF�}��<�P��k�B:���A�r��?��mn�@�70�Qr����YJ���OO����c��v�Ɩ��e�<��_`c�A��:�QCfQ�/�!�鉘IH.x.�dv��n6`O�6��K|�N=��s����-dg���	lE�4 ����_�bT�b$���x�>�1pk���c�?�%�I&7�j)�r-��5}�3��悾�$�w�>�ϟ�xiSo m]4��wmum���3�p~}+�p�ţߎ�����񅓟y���N|�/��]p���i4�� !F/�dϠ�@���59	��}�P@x2iF���y�cX,`�#��97�:*Uo��Y�Xk��@��[�q�cS�7%Tp�Qs�`�o~@pɮ�?��dl�v� �onn�E�K�zp|i�6�)���X�v���4��RQ�*�/��߿�%<�?�*%��kJu����۠�	�<|
��B��1�R?4� ��N*��A���W���,���$�}�����I��D>W��޿�%<����y�Mm$R�l�:r����⒝$���B9hZ��;�p]�7�x�j��k�'!�/���ШnFWY]4�ؾ��( :(�)y��2�{�E+/���`���ӃJIP&�6��i��¼*?�J��3��N ]�9��ѳ��*�)�aT�|�LE���,3�K:�YԆ�}�ڱ�tg!���N�d���)�VrE�b��DL��Fv
@ `a�佺��Y��2f��|m���� �fO}�֤��i��_4U��E�7����pYӆ㾴
�j:M :�xf�T�1��"����0�6*�K�-��e�A�A+�s(���^(�hO��h���0��-�y�d?�Z(<@<��|"�ڪV���2�  cp���][	�5��|i���8S��s�����4�`[�Qw;?�����n�T����3���y��r����p��1�Y���A��۶�Y�L?H ��f����Keg։�㽀�Lu<���gP[��`[���eu���ڲ��9�-�m�*p��ڎ ���F=6�#��������0pǳ�Zaр�#�hwUn�9:�	���U��?�n9��/�l<�L8qL��)ʥ�J�te܌ |�I*8��6g��j/�10�5�M��=�霗��߉B���<G��PaD0m����v�0}�`$;��;5x��a���=��lX�
1lU.a`��� �;�QZX��ac�#�e�'�����A�G�����H_�m(e@U+��ACCs|� ��W��DR���W�?�QB�5''_
�]�c,Y 8Z��1+�qg3�\׫�������3������/�D�K�]�3I�oa/�	��^ڡLf:W������*�(cBy�'��jR�$2yϳß8� ����_�Nl��2gy�`�v����%�`���buβ����GcA]�@����; o!�ɵ'���"ߨ�"�𓮯�'�f�
�4� H#lU��cM$Xk%���k"��M~�s���	���&���y��8z�,�_��|!���m>�uvp,�M�Śe�˧mXō1�b簻�ī�3&�Lv�+_;��A�Ӣ���aI���/.Pv-�և0�{cv��9�����,�����TG�=�ͮ�d�X�^��qP2 	���j�
�)�i�g�gώB�� �S�Jg>���Y�� �d~3��}��|��W�Lp!q�u ���}LLd�	x`��lQ������'�3�/�7^{O���d�N��q���������۷�1�����{=\�=�RĈE��N�Q��Ybؒ�ϱc����K��'��8y�\$o6�8�ک�[��U��	���	�<��`���0`�wL��D�˪J���ӣ�YI������h�� t���Y��p�,��:\��_��\ڨ�4�F�ړ=Twb�p]��p�3 ؆��.`" ��<���Og�����ЕO�G�lo���F�l�d����\DF�������9l��b�uE�Oa���cw�.���Q��1��{H��(�aM_���0����Ǯ�h=���g���F�!N��@�?����r���� 8kp1(kc�4d�Q�	t'�逩Ӣ���3������b��_�g�`�No_vT�xIr�p�U��*���Ͽ�@k��Q�-���/��@p��FA��D/���J<lU&�`h�xx�Ysޯ�8@��ŋ��-�|&�(��H�N��]P:����� E��*[��O�����i�������5u`P�BVԺ�:Ax�{�ʵ����cd�Tz�߮)���HA�����+߇1���vM���aAw������jҹ�Z�>f�X�^��w2`Sf/�d`�֖�y��v��F���}��]�.�h��W��f��l���q���⽬�6��,�p_��	����G>8Z�����v�� >bN.W&�� ��.eGTo�U��!��,�NY�|,��A{H1i�3DG.R��xUr�q>j{��(a�Pw����@*9w��/�y��f���O��y�������̨�'�Ý�� F�KE'�o�|�va�=��h�?��`�)���3p�.T�H�Zt��wm��`�G�0b�x�^r>m���;\�8��%I溚P&t/&)�4�B�<�nC�ʌ�}o�9߇2$�n�^�y���iTr@t{ɺ�]�R�6jN#h�I��+D�uvV_�a���ۙ��W�,��p�vғ��H@��!���N3�n����<�VZ2 ��ŕ��Y�g�3�>v�)����Ͱ��	�mo��__؇3���e���xO�Ő�k~�V������ޏM�9B__ ��f��y�z奯�*u��r�~!;?ΧL.��$��"��Lּ,g�N ��{U�e�8�:m8�G�3c=Ř��������JH̴���f��8�� ���;p 0(�F����M���Q�A��̒k���G�dm�YNA��J�y��t�����/X�����p�Mig�A���:h";�yX?/���s~~IM< fSv1US c]�w�>>�5w�a-�]wɫ���y�mKph�b���9�a�|�L	,\#�
ܷ���7u�ۛ�rb�8^��k8Ur�Y�e��p���a ��O��S�S��S?a7V���l��;_������
ZA(�ۛr�e#���Uب��͘�g9���^�6���2��&��g�Ӻn�W���Sa��m��|a��a>~��h��Y�'xIZYk��k:��6J_����떈�Дw���mtoKw��3U��P|Y7��5z1Y=��<ya�m�.����ן��r�1�R���+�B����\تǭ����/ʳ�6AY#E��~j�_��˚���?���p�8	>=�%�wI%KHJ_��ϟ�����;؊@ׅ�:����̚E�/�]ǿ���6�IL�,B&^~���&l�=��:_߆���CZ���!�9Aæ����Uhs\�~R�-��_q�h��Y<�Qg���6�7j��CT���*L�9�ME�\**��̾:5�0<<�kN%;a~2n}m~&Y��D�Q�#`g�J�磲��G��Q�Z8�� �KT�햿?==���r��R �f]-T�i���1� �@�EZ7e��D_3��g��xo��P���υ��y�r�����U��R�H)>����B����v����H���
w�A][��.z�0;sus�E��g<���Zi#h�V޷���>��!�E�# �j�A�'�����`��ΓJ ޜ�.�g-�='�D��B�`*I$o��sdg�vk����Jݵo���oZ����></���K�]0@ppH������&��}�Q��%a3��?S�p<�D�7~ϏE/>�`6��n��Y�Q��|u��}i����Mq��6�!m@+1a`�(.���{f�9U�&}t|~U��$�l	��j���,fA/���l�5<U�!|�t�gx>˧'�.���c;EjkX��\��Ӊ4
H�n�6���`0��_,.x��#㏮8d�;��3�����Q|�a�Z�%��Vy��Q}Z����o�����!N̷nn�܆|���1~?|il��U�0x��j->- �-�;0^n�m�9y������_0�`|���N�FXtm����I_��2��&ϱ��y�$�L3�umT`;���As�0>G�Xרp�;XRa�R�?��!	`u�=箻���$������-�f��:zp�,Ba��e�S4c(���V��Z��4&�*�yZt��]�]��Es�u,� _�<�Y�{�kykku�0 ��:eܝ�n~G��wb֔g:~�T+�����*�Ff�T�~&�Ƙ�1_(�<)t�DU�����<9�G��rp>\��"Gq؟|����1^�݂��$,��,}��Lj�ys�\x7��[r]v�<#��%��;�i���앛�P�'����R3����'����N�:��i_� E��k(#��Ӛ>��:�F�5*�t�J������*�º�+�a�Q�S��E�	���1��ֹ�fR#f�����*�|���0�zFݠi�ĽidYis=�b@{��h�#����Z��j��y�{���0���tRv@-X�BU����70�k�F�"��8:���ϸ�(���D��}}ր�9�y�*łv����x7'h8�O������b��߄
���8�Ȏ�]�׾�`����{`j5f�W�M��v&���Q�c��.���T��-��ǃ���)z����Q����> �d+ˮ�7�Be�E8��@������{�w,>Ny:1�Ϥr��f^I������5q��b�A�`�+C제���B�=�B���t'D�1�� ��H�e�J`�-O����ڹC�v]�؊7�߄�<'���Z��~M| ��L�9�j&��V������E�G�n�F/փWww�7�}qmن����~�Y>>}
ϟ���}�� y��|�no��7oß^�)���ۭ�a�R�;���9ĩ��� "�01�r�|��'������O�3P'�m]��q�oZ���p�{KР�%`�֚L��r���Y�{�;������Ѹ,���]j��A�l�9��������`'�`�N��h�XCzu#���<\�#N^P`4'n�[��nK
�|f�N]�!v����-E�Nj3�Յ���Hd�H�#T]B�����J&���&��R�Ós7�*�F�����F�SD��A��O?�撂� �/�56���J�,Λ�夃�+�'�:�  H띋m�V�|֫�O����#����N����48��f�|CG7�Z�2ӳ'�D�5�2ѭ�҉��d톷�kN����Z���k6`�/���ͫW��_�_8��'�%����j�����z4z��2_�p��Ťw���$o�Z.��`IV~��so����:P���'h;��y��2�����YC�1�s�������-���m�߰e8>J9�-����%4�W��\L.h	��ٛ0���+8do޾aM짏�3����������v�s���2�9~9�B��]� ������w�*��g�������9�R���������x��е8�ʼ�r��ؾb�,8l�̈-�����(���}�`epc;�6p�[���_�c;e���
�s����) Dӵa��ʣ���.�ʴPp?���~��&�1��Qo�J(xWD���T&T\�"R2;j8�[Eb{P �]�em�W l�v`	�)����v��ǃ˱��v�p�%�na3��7ن�6�� ��\��'�։J?���9���0`bi�Y-����F������i�Xʊ�dκ�u�I&��E30Fϴ�Z
@�f��q�a.h���36q�g-Y� 	�h�?������'�����Q�3��
Xrjs�������pp�%��J��c\\-�뷯����1/ԩ
�-�����}`���>���pP��%�!�1HN��ɛ7��d>�����	y��قr+���`�ԥ���:,��<�4���U�n���m�dA���vt�[�Y�p�_{g�PZ����~��sSZA`��g9?�& �e>�0���J�y������7��bB�>[M�
$�֫g���'��{��u^��[ d�m�l+IG��U^�o��R��뵮�&ʞv���������a<>==��5#����|�&Z����о�s��C�r�~"�$��*��j�.��6H4�l�ac
�*8O�Ma_��v�9�k~�f}�rR�Bs�70����u���k��W���?�G�$�v��l~���c��3��-u�D�L���xޅ��շo/O�/����'�F���B���Q�G��^�i(�0ƛ1�M�~�Ԛ}�Ts�V�\��fHV�]���#��ԅ����<w���8ay��HD#!M=�6̩*)����<�/����!��4�;�-�������I��>:T�dL 2ŧ���������?�~޼z-��F#f�6,��5��>�����?��PP���s��O�v���t���h}~�F:w�B�/!�G�k���k��D���㟋c�p>�8�/~��_�g��S��J1���ac	.ؒ��G�8�ņ�Nmzv�,@̂X߅��<ǹ��� X7W�y����a��.G���z��q����R)zˮ�?����}��C�Z��1��pē��p����i:Ȱ����*�
��cX=���Wg:���]_:ax6��W/uy�;O�������ʳ�֒s�����u��(���rofT��kd���Ǣ1�:3�LS!��R-�ٵ�p�A ������N.�8�v*���l�bvs{�nE�" `0S[{[��1c�J�Ś`�'�P`������Ѻ�V�ZGJ�y�C��6;T?|��c��Ჽ�9�\\s�#5wG��WK3�>5j��O�mjԎ��h����[
+ة�v[�N��©gP'I-͗, ];���&;2���ڞ�Ղ� ����XTGԅ�����������|OV-�����b��u�؁��{�'h}PP�h��+T���m�ǡ�&��(�8W��^%�����cFtuv֐c������tbZ8M�fC���ٌ�c�g
&H�r)P'7�}���g�Gw&�D%J�R���-�!�X7j�(�_A2��9�A��c�>ǧO�D�Q.Ǭ~A������e �s�Ea�+�������6�/��0}����'wd�nq/��/}&����خ���O�:^0��O�|}(_s�gt_���X��c,�/m��gc(�'?��!1��ú#�T��*�C]4����A6K��VN���9�0F�����L�
�(�u�V�֭kEm'FŝJ-�+�3&�C�N���<4۶]vܶy=�U��� ;2���b���>����uk�8��rj"�]�M���U�;8�����I'�Y�/�M��*��V�l�k]�Ȯ����0������0BY�lkA�F֩tK�\C�Ue������߼���/R���C�����b(]��G���$���RU�'@�cV~5p�tx+L��58��)�h�?��v���<�+G�L�uf n� d��[tx��`��b)se�N�d�V`	�U� ��l��e����%�x�,(�$D0�Ԛ �!zٶ[&��w7o�t��T����.7�a�=3�<���IH�BR�=u���Mym��y�����bOS�w�f��Z�f6��Hl���^�^�����qٹ��yY鹒B*�@�3���|�u^��+�/������Hh����c�2�蛁���h���1��;x��XF'vD���q�S�y�<�ٴt�"���ߛNW�%3H)��`� (F0�ky��_�t�21ӆ$��xo7k���&�Y��� d�&�Îa�g"hn�%Zd�P
[	��I��n����O�!e�VL�Wy�"9��0�����X�b�'K�� ��\��k2����f�vdkN�����͡��_�N���m�C|�F�k��!�a��A���`ߍcƎ��žV%�"��J��*�c,ͮ�j;����'�`�^\).
ң�<��5�ڠ��r(f7���� Q�nh�<n���k�U��)�S��zܿ�Hf<��ʖ"�a�ӵⶼ�m����:�P��s����O�D{`�9sF�|5�a�R'�
�;�y�U5��юB��R��O���:L�sLVw���G�X�٨�����t��r�������r�������Z3����$ Oh"������%���A�(���۝3av��)�x�:Ï˰!.���60w?ߚ���v���|��b#��z��o���	_D*����Xp�, WG�^ Pڊ��k��N立��5���h2v�zkR�e6�H��h��UT�V��'�i�D#v�Nu�!���Amn3SG!Q�(���sc�1'��;*
��C�s{\1���������X�) �5�rn��A�2�&�UXL:ES��pAv�B�}��\U9�/��n�
�*�3�.dj2s��\�	[iK���ٵA]a�SQY{�=��/��)({ǎK�++c�oj��P!�7*7'k+�.�w�ŬMg"/�h)�G��J����Y�-8���Z��v{:j*I�d�N嘀�*��:v�%J'�b��%m�8:�����9���|I�cK�n1��gʸu;�ma�]V%s���.%!
6�^]5�TVo��FR�
dB�H��J@U�'���W%��l���P�(�$@�F�]��:e�j�(s����qUW���8��(����ۅϡ3	�ME�pĠ#\9��l����9eӉ����q�c�㏄x�9G-QU<��~���g�Xɀ餣������	�ܟ}�Yc㽕�w���J��t��A���S�J�@]�����Gم���D{�,p� !PFP����M�P� ����& k��B'��*�ٮ�5iRO���SǺ�fCh-g �+`�����v���21��8v(���o�k��(0
 �üh&����ԋ�&d2�"���߳#]�h�`,��2/t��5�18��	$F��b٫Z���d>�JB��	b)"�k�tҦ��`x�[����s�E5�4�T�����so�����wDކ�K_p�W]K�ÖQܕ=�M��;�H��+��侐��1@f�x /+��/�mp
K� �ϵ�U�7�Ȓ�p�Y����b*[�?�7eP������l��J@���x�̼��b�d�Z�@)�%ZN�|�.,l���v�����Ϗ��`���1V�\ �������1	�cg���Ƀ��T:2 >��j�Ewp��d�=肵�kL�-.�%��Q�c��|N�Ue�X�o;���C�e^Q����Q	0u��$1x��� 2����罥~Ѫ��\I��%�z��I2$����'�&%�c�(��7��Ҧ���c�Z]l�}-I8��J��v u�@<6���G��6�c^z��M8p�d���"[͏"���q��( ��t!��PL~$�8<#u����_iu0g}�<�B���?6B�}-��o_4�1�b�V:|��e;��>��>=Bs ������ƶ�� KgA6�mZu����&	�^�L&u�PCuv�8�Z:_`�P�t:3�p[�S�+�<���6�+�O��%�?�*��W(�
��O�g�D��cK[�����yh-�.R�Q:?-D���i��_,r,_^����]x�_+G"& )�����z�x���!<a�ڑ$���!��$v��$�P�V��f�6��!ж������>|Z>��E�wA2�m��A`���_؁���)�X7�&l�\Φs�a!q���6l�y�O�Ǉ�O����>B������Hf��`G7x�V1{����Ʈ��79��oTA<:A�
��m��@t�jSP.lY��1n��p��a�_�{��iȀj��.x�a�t���&Ͼ�	1T�7Z<���b�
p���M�~�� �!x�ⓨ���5!��Ȉ��#8�3>7$D�*k/� ��A/�`|�&��X����89��޹�d�t��8�|L�9Bй�3#������z����y�oC]�/���jK>�&�`1��x�&��B�#(R�[u@��l &4Z��r^\w&Z����ڄ�b@��Y�^9L;�e�Y�T�=`=�0�5�Q�֟����Z���T�_U����u���2ӕ	}�I���פoV����+���
����e�3����-���r-dq>(?�Ш��tEs��	0Q�E�Ǡ�Z�4�����˒�f�sȒ�}m7��:�qt�Z�n�b���^��Y�2 �8�}D�n\K�y�n[&���X�,��̱�(��Nd� :��q�qw{�����Ւ�8?�5LD��42f��� �~i�==�?�9�^*=9,w�vJ��?3�+G������5�5�KF����?u�1 制e�Ƨ`F=?�r���/>Z�9
��.((�߻2�*�4����U���?�]�R)���`�X��+��lA���:f9�Lp_��=����֢��3`>�ɻ�D�;p $�
FL��S~]���x?�����!���,��v�8^O�����8�ч�Y�u��5�����Jl6[��g�7�"�����9/V���߭;Pk�2�[���N[��BϺ_?��!��?�r{�;�`��wl���d�3왪��:�E(O�s�C�[��e-[|�u�Ї��}��u#�?�h\t,+�q��j�+��5�X��(x��
8�;�M:�+P�{@���MM  �wv�0n]�!�߾o� �Ai�y];�f>�/̗��-=g�Ӭܟ$qv 
*I�d�s9�3�V~�����	�w���X�S��,!�0��1�	��\r���;u������{�*KQV������V-η�
 `d1��a��{jp�[k][��hɺ%u���L�-
��YI>n��>Ȯ��+�O�U(v�51���:�r$тٱs��:���g�B(�va�YRM �x&ul~:rej�����Fi<5_Z�^�c�Zy��9��S�_����l��+6����cWf|�N~>�Y��=��l[�G�b����0I��;�W�={�H��?]h$��Mb�����������Q 6Ϝ>m-J���y�-ɰ�V咵i|�a���)?S5�)fzX�^�\��oG���9<�_���c��:�����0;c�f�+Ɨ u@@��$��~���O�aI;��F�C����!��e�߄u�	�����"�4���O��8g0�!ñ�*a�)�=�]>��V�,��<������{�a  ���
o~|C��� X�ϬxX\h�1���pE�����bmY�&2J�P�`v���X�?�G���{0 ��?*q�E-EM��9����2>y)���`���T��� )�w&�;��1@��Ӏg�R1�F#��0$�i}��(�/���O�$˘�d�^/�ú�[��g��ꍆ�����QK�ht7���Q�[�l�;�;�K��1~&�j?�e�� ���,�v����vvʓ�*�{s�Y���m���X���@��rO�F�4,�k�M�:M��[G=�oE'
獲���q��p�$g6E���-�1O�53l�g-9��O
�������ڞ' 8���m�V�E��K��� ��Dd��:w+����$��So��*��l&�{]'+%��m+�p�0�� �'Z�"��?�U0l:�	53x�!�7�Vfs�����B%gD�X�c���CHY,%�Nޜ����ґ�o���v�Q���@�,��2<�Uc̽~�E�b�XEs��ߚ��/�z�[΃����ֱQ׫���p-�7#u	i,2d�ǥtC[�Ϸ/%x�c;��~����e�z�N	�=w�'��n00e����ѩ����3�a�V�����$Fi%��k4́
ՍƔ��H6ΔˠU��dl�%���7h �γ3��ۋڜgi !2(���`�i�fD�I���iǛ��:�l�c8a� ԏ�?|�q�����{��'F�ɦ��S�S'��A��w?��k��,��ڝ����@ܜܑ]g	�z%0�ΰH]���2�8=� �}j��g��]k�~g��������2��6�MpʬFa��K0}7����u@�j]I��q��ڌ�;�������`�4��s+���Mf𖉍�����s���ۈ{�M���(�Dg�Ɉ譫�X�uJG'�~~y&��f`��M�.�J���*6��gh ?̉�6r�F��Y©+L�0
��"ˍ:[�����9<5���'��<�<3+o�H���R�ۜeO������;�#�k�����~��3����ܟ %����,�maq#{�n�dO������o$#x�3���{�0�,���r	x��zyZ�ʾ-�z�e�ɰ=o S�6����v&�W���Ҹ�	�m�.�>&:2	  �ږ�$���y�Ru�'��<�2�6����L-��FnN��_��G��Ϸ<���a�1r_�������|���#�bI�`.Ĩf1-�v�K�k�|����&:@�b��\k���	ɺ�"i���c��1��Ҽ')�5!4�ߡ�S�΢S�ySi� ��D�=L�U�	�Z"1M�}�U;Ap޵_�%����^�L�`cb�Pk��:<�?���=m.$# �y�K3jފ]��=<=��U�����!��O���Xs(��>ͺ[S⁉&�=��l`�	��@	�z�V2�4r1�!	3����;���R��6�V�;�?~�X4� t���@��4D?Q�mkݚ��1��+Ċy}�-d��WҍS��b�$1|�,B��4U�M��ēݑ>2+��t��!`���q8���`~�3C	���c�Ƴ�Y�����5ʰ@��]�4������_9ǗK
�9��>_E-O��#��Vv�d	�`���h�FE&�Yũ��[��O �zaN�g#h-�p��)�2��q� m"��n[�x��|�N�?rʜ��:�� 5!h��
'��$Evb�4M��I��u11�_,�ɄB�"q�F���"\^�2{��l��Z�N-<k�6�௷R��4�(�<giʀ�~�]
��,h(�8�ܽf�>&tG�+Q����W � [
ʉ��C�2hl�(�(�g5��!���k��;8���ЉD}9�ʴ����ҧ�>��58��� ҙU^v0P?+���E�n��ղ-?%@m��@>_��TZ�S��fS� ^ђ0��b�,U3��VQ�RR��b^!(�b<xV�׼Ll��9z��r,t'>Y6�j�J�I��r������e����y9����x�_KŔ4���Ͽ~℆��R�g�-}'���}v�3�V����H��`u��][ɧ-�/��Ɓ����y?���J�ف�k%��"��C�5,�k�*G K2�#as�M߽�Q|�<)L�a���5Ak���� �-x�z=�v��O�u(E�2�vp̙�p�}ꋀ��\���X�3��U#�ͧ4f͎�0Bpܰ�Þ����>G�\q]`f�*���H� i�ǿ�=8��x��������<��SRv���i���������%��𹓁�|,�7�g�E��"�^e?��i]���`��c�NoZc�!��Ru�x�b����YG)&/�2kH��AY�қ.b�X�*?��ɾ J��k�:v>�� �E3�!��(�<��@upBY��5N��o��_�)�(��;�4�:�X�y���d�0Y����5&��qT�(d��|,���0:RQ���:��[+�����EQ������z�	�{�yOV�t^�ɸ����x�r���Aw������n2���A:b=1�n,%��ִm㍁��@�� �C�v���ƞ�؜Jܩ��4|��i�HdkeV�A2u!S��҇ڛ4�:~I�'��Q�2FS~��U�%�������J���I������!�o�J�Wn�(g%��'GI��Y��{#����,�a�=�g��}�.��'�V[�H��S%�0"+��� #�d�>��:�k`����%]8����˶�_uE�J$m�G�ֹ�	�<�� m�3�6��A��çO�S`�=>>�o��A�<��D�� `�q�ݘΟ�`�|��y��]xX=xA/����ک;�j��O����@:�_���`��8�G�h����s:��nKM��~¿���EYş(o�_��Y�G���_B��@Ж��6�K�@h�����ڧ"����G�s}j��P�W�`/,C'���{*�� �9�` ��D� tu~����o�w�af��P5�Z��G��M<-�Q�ίm��u�*j�ζ7 ĵȈ�N��� �X]��dڊ�\��86&t{�1�s�}�϶X���m�1�Bqv<+>����neu&��b����9qJ�+�PV��@ӥ��1m�;Qf���X��MTW��
^�os��21�M��������TͷF�ŗP�yY]�=!NLB,�*�$��N^�6���ZG�h�WY �iS��qoe���R��k<�8#��8�V~$:��(�p�LY�y  h8�i�k�@ji�:w�6�>��J5�DW&�CTQ8|0�ʔM������	D�'��%*42ht�@�X��9� w[�jg+�V�..C9Ga�UR��AUk֮ Բ1���� [�V;x���|���GϬ��؅p�c�����,�ֿ�)�����>�E���>���?�����C@����,�]M���v?�i�� S����籌���l��H#;&Ʃ�qC)
�����z��]%�e�M�y� ��zo�h�t���X�A�����<;�=�wd� ���9;�?gj��I�����=��A�����]& 8g`4#zB[�+"��Jv��Զ�	�ZY0he�1� �J��Sg��C���	| ;�uɞ��Z �*�Ӳ.�;�}�<.��8���P���{n���}y��;�z��Z9h��vN��Y��V�����Ղ߽1��vG�]��k1�����&� M�����s^�"� K*�~7�7NP���T��U�6dRP�4ṁ���C��r���6^�D~��� 3l�D�����7�
�cO���䕘�]K�����C��t�`��WU�bh�{��񡽇�Q������ǃ����[mb��uK�U�����JΙ�����F�b�Z��/�O�J����7��N�<>< l��:z	�Ɵg�q���&�o 6�||3�q��P�s���?`��@сj�mFl�M"�؇�Q�K&���O4��H�����t4ґ��L�v��KW-&ck+��|�=�V�U�P����'u��>�fgI*k��U2�:c#6�=�x��K[���=J�ݖ�y�^���<�9y~�
o�{�bY:���`M�� ���J��q���q	��W��<� X�x�q+p15�0��H�hc�I�;�=�T�L���y���V�U�`�i�+ݑ	RB:e�3ۢ��B��w�^��o߆^�~x��!���J��K:AO������������e>��<nLlX����[�� 6�����	]��XU���'����p�+`�����2�Ke]�3����"�ن?|�m��P�O٦b�8��A�4��g4ɾV�B��m��G��|�-��QN��������}���#;�çl/����y�y�r<�BI�����J������|��Tl/��S�~4}W[o�Ff@��s{{C�y �@�Q󆖉T�nŢq�]_(��_5��`��@U8N�FN��(j�3{��ʐ(�U�����3S��ӃR����e4{xP1z>�T�PH�����;�o-��3�`�
:�u�L�gN�vDǚ��TfL��n�[�. ;��������^\.���C��h�3�壌����3�lˉR<tT*�d�$�Pr�Q�ރ~˲A�o���+��NV ��q����X�l/�\���s�}KlKgF��މts�Z-@gsZ�%c�x�>[�R�-3f��y���t�=���2��q���a�c�#`'x���0�Q�dv��J'
<w��FΔ#|���VB`�Չ3��s��l���Lh|���g �.�v*qC����t����0�i��!c7�ܸym��[70��-n_2i�3^e��rPw�>sѾ�!L_n�K<����k�"��nM^9��>�yL��2ǔ��J)�Z�p�����3�<�U��[�Y��^���g�����f�R"�r�(gdCB�:���Ѿ"���:Yfd��*&S$t;Q�Qw`��_������Q
ec�t6��öA#(����
�z; ��N�����5���4��8?�_�a��2d�۽��)'k��&�!8Kt�����-3�(Q����q}#��f�}}s��x^���LJ{��U�5'��S�p������c�L}�<F�� �����5�i�ތ���VE�B���}pV�A)�ا��`�/j�h�J��>[�G�T	am�s��iR (�b��X����dlL�˯��Yi�f:W��|��t�⡓�V��t!�d�밎���u����XH�-��-Dm�[Ӻ��E
�b�g��@S���93�S��[�k"�U)��r�$u�ݪ�I�/Ůgh��q�HNy��r"A+�?3�u�`�����o�%e����:aH��h��CWs����t����u���`o��S* �ߘ.	~'�C`g��$��v�-�gAƂ�y���٪�l��"�B7�1�NuU0_�&I0Fgr]o�[M�kv<�N+U��M%G�<�	�e�F��������8&��e�/�>��K������fPv�9�^�	��C �Cu��/�7�q`�4,0�D/6;���7qd�c���D��HM2�p-jG	��J�������Y��|J�b��(�_)N�1wԻ�62mb���L|/�7��M���G�(t�h��3�{���uyu�D�S>�E��=q���6�t�����o����`K��3m�I��*/G)j�j��U/<�}��,q��M�0�;��`�lBj���9�����d���L�5�|B��n-�@��;��m���%��QR]j	�<�ϢRc	�T�:�h�#�g�W�ӧ'��(q�5�o�������hXv��ɃY;��q,Pj�͈�Τ�elt������Yo�iE07SgL���*�8�_jt&N�@���V�٭��e�Amj+kC�Ƕb'.x����14�X�p`����(�3��L���������	�-�����Y6ԋ�)���p!�,c���鯬N�ۜCto�	#��#�4�-��JX��^�z����F�v��y	�������0<��h"e|�5c����!��$�6ѵ3�j����O�_���|t~ �D5� :`[�2ي6�l+�m��PC�34r$��AM�ի[ј8���m30M,�莏�Sr���lT]��˕��~�����%fh4�U�����tX�a@F�G�K]�*ֆo6E��7%\�Y<φ_�A��\����Ֆ�R��X/�L2�j��b�2�͍�����/Z!�v��@��}�F�o��m|�5�������OV���z��uV"�r*���j���`͗-�	�H[ lw�m�B�����NB�X�ɐKjS�͟��Ȋy9K�"�������D]r�����άN����5�&:�.;Q̰�D�Tj�H�!�cS@�u+�l��X
7c>�)�sپf͙?t�<������ �-����I׊[����	0�`���k��� ��e��ƍึvxЩ�b/QF�A(8n��)�N?�a^+`k �1�����D��.1p�ݴDИQ�w�}�|s[9@���+�����es�7O:�Ҽ���|>�h�����X�&o^�I̥�G1?��{�{�I{wK3e��y�U��ؾ����n-6��H� A��<��l\Pp��x�&ކ����x���*�B�������|Jm��(��	�~�v\]*Q��N2g����H �R&j��gs�o%��L�1h�p�v��Q(OGR��l�$�rl�9�ɩ�g5��Yɶ�]�m��aY)�l���^R�I����9��u�YW��FC�JW,���}0�q01fXM1i9�Y��'��g�e��BM$6��b�sj�띶j
_�6@M	R�:��	Egڀ��L�E�Iټ��p���<��tSw��}�l������B���l���s�u�ȐGE�4�ԄՄSJd�;�~H�F��X��ܾzR��PE|�۪�6���Y��Y���-���,ϭ3V�nf�H�*�k��[�I���:b֚VuXViXwE�
�ctĢ�s��`D��W�k�N[c �`�����A�6%�H,uƾE���p�Y� ����Bv�*�m�f�5dAV����H�&NɴbYV�����8R��u��Լ����#yoI���9lvbtWS�S�]���/a����������(/_��L2����xP�}�B��f1  a�#4Z��R�s�b��g\s<={(@�S^aX��+[���r}��8#�����K���A� ��=|������ys��5���EC0M_�4'�5u,p�Z�z�z](S߾zm]L�� jt�Ǽ 	/�,^�b a��ű].���;�~|���<�㿇/l��.w�� ���E�4�HT^&#�k�7����0j)�48,�0>�Wٱ�w�����Axd��=%0W��u֪����y���O��c���:H����	� {%��i�C�:�(��9
��-[���ʏ����Q�FQ�]O�t��G��1ﵤtv��Ev����=��S�l���(�!4���ͱ!��<��<��1�<Af�/t;	��Ɂ =S�j9�[`�ՍV�e����q~���p_���xݭ� �Q8���N�f�-])hpZ��:��<;�s=����s�3��@e>�R�_��}�d�����Cc�1�;YJ&�n���Ml�%?�<IY��B����ּ�|Up���P,��}�;���"|�Z���l�N���ˀ�@�L�1��=�8:����������3���6USH��4	�h�+�	��Cf�k�1O�u�(�Y�ZM����%R��]�@���^�[���X��1���������i�[� N�Д��_�)�
�[�=J��h��ӊ� ���jj%���?A~�B`ӡ�*�^�.X����AZdχ]C�
J�Y��JO�g��D��աb6U��b�Uvo��π[�H��g��Ɇ�A�L0ؾ� Ѭ��9�df����ڄZ�����Q	��k�3Ϳ��d'�5��G��k_O/��8.kJ�u��9�3Xg�Q&o8�h��阎ݿQ�ރs&����m���,)g0U��ps�G�Z՚W��ukI>Ub/��i݈����X��L��T��Ȧ��i���p	�������X�#@;�)�<�zƚ|õ���\����B�`��_.��t������u�	�p���B-���'־<a�NlPG��V �~�b�����c��O�������X���*Ln,E�W�]p�Ԅ~���J��(��/��$$��Z�%Ic���Z���kgBj���N��	[�~Q��i��U: i/US�.�/�-`��S��ġ7����|]�e��w�������V֦'�]޾������F�S�b��~��5�0�_k]��7��o>�ѹ}s莜
�2����09�9�y[��,!~��=o����,ΰ���:6�`�m��Uh��5��Y������fs���	��B��iv�<���4�c��̑.��j-��/�m�r�^�d�$x��X�%-ϖ�ֲ��4�+b�l�6�5}	T���H3L�ǫׯx�@8�P���	�������6�)p.SK��/0����ex�,���L�!&���)݃N&�P�?C��!�����K���� j:�����ۻ_�� �c(:F��X��F�s�&}+�{y�a��\7��X����4JF���֌����W2#����a�mA� HѺ6��P�V_��B]���XL���}~@��9@Q;Mu��*�翱�,�"��aa�x;O�
T�µ'bF�"�� �^����lMPϡ������x�Hz*2�w��~��c,�3-�Am����l�\h��q/��Z��g4�v�!{�u,d�GO1�������cl�X��d��.0!��'��n"8&4fh��I�g�5n*�.�(�4fg�"߿W���ל?����ğ>}�q��1B9S���m	��?=��H���RldQع�Z�ezn�n����\���@OD_F}{311�"���̮�1�9@�(�:ׂ@V�C<V�����Rϒ���=�����7׷D��/���h�����]�����P n�@����?���-�/.���Ӱ��t�T���d��h%8�lf3�pA6?�X����[�gǐ �5�ϋ�3�{��x�����kjq�B�,"^@��a�4�9��,<���頟�)�@vC\`ѰY�98�cC�<0�T�9����у�#p������o�ҷ���ƶ�+5�����L�E�m��?����b�L��q�F[?������N�X����[r��M�#�8�M�!����Ku���Zy.+�a���(��=)�Ne�9[������6Et{Ƞ���nniC�V:`�~ ��q��+R�nv,��XC]3��zAy>3�P GP\c@�-��Z�n��<�M��Pե
�( ��@�~`���_ޅw?O��Yy펠=�::-�&0�rQ�)���K�[A� `G-��V���=Έ��XY���]�":�������k��ٶ���,8\ek�x�S_�-�_�EQ����w=���דF�妑�emLh�1
�/�t�����8*��T��	��£�n,s��_e�V�X��b��%�5�{�����Xv�~�� ��Apѵ*�d��Yzz���<�P�b��5?��|�&$���g�����2���`��z��n�:�F[c+���,��� �=���k� �H�@���Y87J��鏱|���wS����*<=-��
Yd����Z�be>�$nLP'ۋ���p���Io�sN�&,��d@���\,Lsqnm��fyT+v�e��G���rзvAcK��A�����X��ĩ����Ya� �������L�x���Kv8��i%!0��L[����"d���1�'O&�X���	��?C�A�k},�d5�^�J�����H�y8u̒'����AM��ھPS`��ݐ����&Pg��|�g?;v��{ �ݲ/`h�U���r�Ev,$�<nns�tw3��^پl�?�3����)�^ˏ�uy�}�����9W�;L��S�8ԏ��'���\h��B=���L�<��T1�*v���Gu�`L���	��g<�rC�>�����"�[n�]mÿ�뿄������Z��{_�s<����=��df�5�ǁ�����~˕i~�u�ml>zGN��>�$�4� )0�Up
K�8���!�] �L'������V�T����6��x�E���J�;oV����d'���L��n"�I�\L�}6(?���;D�x�ć�����S�Ņ5�ɪ���`:`0�m~��X&lgIDL��l�#�q��N!�꾟� ����"���+�)j��@��%����Y8�X�����lE�&bBT����?�Hl��	 w��?��јR����̎o�7F	's][���w��V�r�� ����:9e�(�Q@>�eG��;��FN��l&��Q�	'�>��=L��$���v�� ,�c���bҗ���`�A�c�{qx:��@G���sKa�mxBvm��1����k"v��zKz�?9|��F֦{ו��Ų�l`�./���M �����@�ڟύ���Qth��ϼ��H#��GR���Z����]kmZ	xXiҸ<�(�84��l�n�u� �0�%�,'�g�Je�P�6��w�#g-Es��.Ռ�h��µ���(z(�,� (f�N{�LĒ�(�.��[�9�>�����y��ĳ=.�:,q;�+/N�?zK���َ��o;|:"-��x�K�W,ā}�d$�p���e��w^G�0��"�2ćS����+��A?ڙ��| 
�t�@�Ǻ9X?��Ƣ����=R	����0]js�F���p�*[�ֻ��V�2V#�A��g��� �� ���I�LE[�+�T���;}1�ci5|n ��XY��9%Xv������Z7*��2���h�P)�
��0��x�1p$ńrq��6`�2�UC�س��j�
�`چ�!H16�߳}����㼴�S�{	����q��@�Ѝ�2�?�P��_1B\��K:���#u��?����2mX�����ȋ��J礳0�{���no�]?fp���Ч�t�ͮ'����o�;&x������ľ��1ӛ�!^� ,9���f�r��r�d��~}fG���9�d���>k��J��|�Ϸ&�˚� ���C�n�f�}.Io�*�B u��yNd�TX�%+�����J��7�XuWW,�g����;$���z�����b%at��*�B��$��P�c:bM5��ff�ݛΚtH#f4�+gpM.��2Pɓ��P�5��`�{�"M�R�w�U��5]��PS� ����&d��^c��t#��l���b^��ā5�h��J��>��S@`T<�i��f�y���p�t���'&����~3#�s�1u��4>;�a'vSN����XV��sfŢ� �5�*��d�\�u���2�}��)a�=��y���
�ƒ�$IX��T��:��]�Ls���L���1���R�I
5w���cSk���;K���h���2�_��^�I�F?L���v
U8�~~������
6v6�6V^���� f7�]���)?�;�?VQq �$��u�-̥$ۘP�G�dO1�r΃Oe�-n�M��<M��ܲ�o��t�g��������c�p�f���1����b�3��^���H[S�^(�4̉���_O�	�����ʈ�t� Ct�E�[-����$��B��Y�����&ݼ~Ōe3�,�骸C�s�2c�߻S�߉)�l�#�#+��(��{�:��{^߽���J�R��BV!5�����`����B7�җ{��r��gғ^
����L����,�V-n��Z�%fwM?4y0� �*,BRT�s!��aO�k������Iy�O�=`.���6�ݻ<C=��X��.<*G����^/��$k}me6{	gn	,I|�i�^P��8m��E��Mxzx
��a���.F�Jv��dc�I�쓂�vx��2��- �~��1�����}��ݻ|�6bDM�����Pu#`d��?	~EuxB���Y=8vke�����b��U��� �`�P�"��wi�,3��'�����zu�� ]��E�u�j ��
�� �F '�P#�=�@T�dѼ;+WCk�iq�&V��5�s"��<;�(_����c�k�~�'�<�b�<Xw �?�p�,�#����~�������L��j�ơe�k(�!�P�*_�N��Z����((L�tG��X�v�~�ҕ �V��c�SD�x:n��ei=�yjE ����I`�v*��J��BT��:Xs�4�B��X�x��V-��!"�@`��]�C�=�"گ���2������(���S�:�tv��m��O�eHB�1x?g<H��4=O�z�{�V�lꆡ���GU��#N�΍� ��4�ַ��Ʋ��E)��X���7w4�Ѫ�R��3|Ɏ�k|����80ӡ](�ҵ���*!�|�&��v&,f'�l�bzHȻg��2�Q��L�{���_]���K:��� �Z/�bq&�ԥ`ɓP4U0��==��:ʶ�[�J��$~Rm�%:�ب��ᥑ�vJ�%u%�N�	��m;1v�ymXs�;��Bq�kO1֎���-fl|yk��	:`�(���S��������Eݢ.
�s��4ʒ�x{;�UI�͒SACw<��ԃ%hf�kt�1h��,��XN�ՐxNH�E�f��(6&K=�ْH������
5a����!6vU humM��5���r��/v�L����;�Wo��}�%�0_+�Z�N����/ @��Wo�Q��j3Z�v�p�9 (k���$7�7��g��?�F��u��TL����~��f?�$�������s%��-��mv��<O�B�k�>H������Dx �l/�����֘��8K! �e��ܮ�����/ N�cc\��8����`�>g{�
�;��`s�4�%
Ŝ����X�4�,i{��Fa��f)�ƥ�'6D^p@�mkϡVIc-{����1k!HQ�ΚJ�JZ�땃V���`ê��ئ�s_�i& t����]h��G>X:��0A�N�5�wŒ��bQ�-���U�_��a3�4y����-���X�i�X��Zx�f�ٙT�?(_X( �t��"�򚲤��7%܆D�p��BA�j���m��]��r=��W��A��6�Meh��VE�oŭ�ё3PբA����?��?So���_Y�i�|$c�l�3VuǇ�{���F��Q��yo�{�p,I=DX�r�!n������#�����r��	�?9UyLt�� ���tob��1,�a�b�� \�G��cQ��7:B]\�3(���U'��ޜ��@�h���gn}���b��]�{u�v~��>@�%�l���,S���EP;-��L�R�P�k�žčrڼ�W���Z���2�0����~Ͷ���]X��pO���C��:��r�kҺ�f�k@Ǯg:�Ϭ���b�=C�(*�S������q,�b�k�B� ��~~Z�aY,:u�:G��%����y���Ɯ#��z�����S���g�U�0R!)�8�^����EX�Vt �Vb�]_wG7��
;d
[��R��c���S��1Nm�Fƻ��z�w>�<��;؎}����~G_�d�����o}�i�x��3hs��3��%�b ����-�?jw���ް������B��� ���4��ꦒ�#�}}n�0����V��r ��Kda;�X��oA��Z���Z���ר�F[c�X%�^S��Sh>u����|:j�t����ĕ�¨-L����͡���z�
�vk���YY���h���������r?��[���U�5P8Z���۶G����X�q#���a�-���'�A0��7m�̝�Z�d!�2N8�B���|�����S'=��>����� ��F����G j�ΞD���o+�ڲ�/����Z%CýC�Z���vyr
��x�z:wo^�ujή�Ȯ��OLN\A@"v̒��8sv�2�ՙ2,�n��=����:�]��kX��A6��=*Q���ey^��ϓ�芬f5vHd �q�u�0��U���_���Q�I�֫����j]��k ����r'l �j+�*��Mc�|^���m�w���v����ihPQ���m��g�Y�g��m����;+jk M�쾘73���7�k���y��,�7�f$�X��
`��{��Ob́�@�g�V�b�uo��q-��KLr%�4�Z\�뻻�+�D�vW��=�]o��|ޱ��);6Ke*�{�/}���;���m��ʭl��=��[{��8t��'�J H��_����������Chl�i����6� �������<ۙ�%z��*�S�g�;�!�B�J�>�n��C:L�$���|j u>�dG-�Z�Ѝ}�R vs1�t�dA`�bf�" � Z:�-�9��K��;o��9������J<���"��]�F|Pr��|욊/�J6v{v����J���B݁��}g]�F��8YE`��K�5.�Q�|��d������l�?Ö�y�Q�P�
4�.��dlsP���1v
���Yw%��w�d�#���bv���@��=�+�7s`ق@`'�7	tt��~��2�����|��O��)��)��J�X����m	�p,\yp=|���=�����C}�&Բ�i�>���V��,� ���������@���G�n�0ר5L��\]��+��p6�̎�c.%1�躵a\_l���xfI��S�c�,���v��p+�a��QĘQ ˨ׄƩ ˵8W�dź�]��A�ltQ��pI -� n/�������ʅ�&�����BP�$طP'բ7�fja����y28��5���������w�*�_|�TR�`d,���3 /�������u��P��<(�B��#�)P�f�l����JBaW�D���w�� ��>;(`�M<�߿�%�z����%t&g	�;�˚ ���5��p=�\�bH�k�ʸ:��EE����i�y�9�l@�d�`�#�Yh,m��~͌&	F��y��?������~^�zn�u����/��" d��������]���?��`���T�=��uܾ��y�ùR��3rsk��%n�ք�!��8 ������ '���[�=�:�̿�{ۼq�mpp*����4 �d�����Q���LOY�-��}��Z�nTV�n�E��(�!DP��5�t ��${�Y�۠D�M�<;��z+���s�w;�I��	��T͐iFp�+��]��<g�A��si����=ۛ�˫�K���.��
�bv,v�%$[ˈ� ���)'�f��\e^���@'3�t��2x��*Ɍ+��#�	�G�u%�''Xv�	�`i.��'A<���@�/n�����ow��3��{7w�x���j���שS2F�f,�/���W��'�h.������x�_u-���p P�ff]�76��T��^���A� �ϐ��b��ԙ�4'�# �7W�͏���';u�z��L�0q�y�,7J�V�>������g7�|nl��UbE9*���1u�S#�Jb��'<)��B����OLL��,���b����)QW�HI��b�c��g����;v�X�����>��hy�m��>�}47�,UU�Lj�褶�S�:Lr@�\c��`�ֵ'�f�U�w�{�10Y�&�+����C�!�e�g�Q���V�˖ee�����Kr~Ɣ�W��"FZ�d3��K��\f�"D`L��vN�
` �}��R�!�C�/{���g{�?���*R�5�Z-��{~ZꚒ�Bg�Kvb��9zV�>p��u���v����6�=ҿ9o|�ö ��`�����Mw�m#�_v��/���:+y��k��p_
�O�pq��K�y��]<��)��&��9z�����h�$�����y
��	��˸�b�l�M=�g�ʱ�����V[3��y}�1�_��/���'�#��^�
��+`nMK ��'t���R�.�:���N�������m�q��� W5`��h����!(��k�VU���U������|}�*�c�d������b��f/�ɤ.Z^,}��D2|��Rދ�JJU-�^7����������I9.C��»��C���|�^����W�s4�`�x��Cԍ����I��u2Q({(�_-��	��9�_��������R��zy��_/�^fg����ل��ӏ���&�D0x �����[P�^�������@�ur��|�Ε���pl��-X�(=�͑SW�l��X4�����\j�>7o�.Ki4IJ�Ƴ�,��<�/�&['x��MNR��	�Kf�ҩ%t*��,L����X2Sz�t/[�5�s�<g���&�S��m��Be>W7$��0�cK*�r쭽��΍�^B���EU�8�^-�	��}�i��1�r���C��G��B�=شk�j�]�� �xqND��!���&��va���(Z]&+/�N�h�0���I4��C� P`�X����H��Y�frF(��� ��s�� �aǚ3|>�UZ��+����>;�IP�z8�K:�����8���������ҶS���e�g	���5U^��Y�B�`O�)A�(��6���v7j��1�X��)���Y_RԛТn�8��r�.�JW��\���;_��|�s�����˜NڧQ�ଙ��pJ�lT�hٱ�L_���W�ᐤ�c����:�sޗi`��ロ/ǵ�m�Iu�i[��u�H('F��@��M�lOL�N�*ϋ�f6`��~�Y��@��@��b�/ ��-6�=�ZS�"�hgz:�'d����e���3�n*���ڭ���V>.���!��R�n}r��M�|�߾S�ѵ��G�v���ۗ-� q�_����X�#�B,�����;.I�L9�����E��ښAL��r&x(,�h3�����$`���2�ޚ��* ډ�¾�XK�5;XoT����Tަ�5�l����ʸ./)W)%lZ��u����qR��w򂦎��"K����bi�tT]?�2Ai/C����4����F%KndL����YWuU� ��v�n`,m30g�v��H����:j��o�F@���%Dpg21�E~��_����ɶ�R�}�\�[���4) :���٨2>���Z�Rx�; ��K�}�����7��ȭE�����"i43��������?�w�g<�H�^{f�8@DdUu�I���)��*+32p  �ib <�Tpd1B��jF����j�dj�h�Z��Y  ��7R���z+�������`���y^
����dn���y��Q��]�b,g&�V���N�,F��7�S��֌?O��p�����g!s�k^�Rq�5I���^Hǌs��>�Z%��/i��n���$G(��jz��(2PS�����oY}3�A�L��~� �g�"=���D�r���Q�i�ރ�>�G�Yh㴾�@�LG�%99�
5Ѫ!�[�+�2�5B�\$�`�]��n�j�9�W�Zw3�u�S�b&-j��]�������^0� �s������ڤ���m���!�y��M�VHv�۫72J�=�5�wd�@'F�D��l7��cS:;G����g�J#.������LA�զא���@�I|u�Z�ՠF��3��Fs��;Ʌ`Ч;aC�6L���WDҚ��e�Q�߾���'y�=u��@2%���V+��^S��ygy����à��E��B���745�������8���M]Q��8e���ҹ�e8��`�o�ʇ�<�R%��{�K�%�&B�&N8fe0�!���ke�-<�s��Ƹ��rRoUШ@qC�t��H��.F��S;����ae+�۹a� �go�q<t�?�4��'�K�m6k�Y�m㉑inM�#u�-, �<�|�.6�Ma圇C��T���I;�E�pF�gڂ/j�>ó.4\:0�^�[�H��4x�'�9�utc��0Bg�D�H+�@EY�O�T6�PM��D*]��!��75F#˧� ˚e[*�P$E�xC85���V��M�I�u�fZ���-�>nFl{�V�AB��HR>�TJ�7/Vr{w�ȣ��m��cP��7A_����S���+m �w�NB�n$���N�l��s��}ߪ�,�U�k]�3�;�S����{#c&����'<mt�c���D5�1��f$jW�a��+4^Ca��7�|����\��cE�s~�����Ԧ7C�w�?W@}:3|�W�t�-�E�Ar�x�g�L�|�*A(]���w�}'i����i�]��a<�Qr@pՈ���q�s8��:LT�d�w*3FF4�.}G.4ilmF�hg0L�D�[W6���(  *|�6����G�4��|ޤ�/t�l� ��;I�������c�+��r��V�zy|-� �$��z��n#���\ bg�(<����mWj�|�����i��n��-h�G����H���Rsp���C
,;���`�B��=�	�DK���K�� �� �E;V��%�z�%e��v]!�1�V��SxG:�j4�lbE�\�B������T�q��XV�W�����C�%έ���|�6�ʝcM�Z�r�tj<��������b�w�E9*�G���qk!�l"I��t��+�' L�ۻ[�(��5�/<��b��93��FT3.��$�8���nV�C�)A3��� �0^k<���Ȥ��":\��,�2�p�]˿7��y�,F�_�������6�[�ܼp������;M�)��s;�le�9ds0�� �d灠
ҡ�m�
q��'��Ԍ��N2@�iU�b���U���΢���X�E0<����P0Z�r�m�1���[�QGzR40�`�d��-@bV��&#��N��������c�Y8�A��?����Jv�z�67Vmj�*w�K��5-��V�Bz*u
�(�	�(?���d���ҥk�1��zkd�LɍZA�6d�s��n��p�`�������!�k��y ���P���RP�S�1<F�W��S�SzĽ�E���!�'T0���O��O�9";J$��Q��X[/,jf�Ľ�'6M���E��:����vl��岩�v���|4�Ee1�ȍ�K0Jٌ�B�r�x���<Q��H�i��n��n�>Q���������V~Y��Q�/��/Ţ]�<��wX�>AS�!�P2F���Zγ�R:��Z �X�)Di"k�Ή�/�m�P���4pD�ܴ7��Hh��DR����l��J8�+������-͆Wh�S������tL��g�:�^=U4�S�}>�1�AvX�s���VF^�"�,C�G�:�LNXvw<Z�>]*�b�	Ӥ��AO��!�QA}��kzTO���aD��^F��7Ι�Zn��h�w�����#\6x8w�b��t.v�z=M�á�|i�' � @:���2��~j^��r��TV1�4:nɔ=7c����RNO{�4S%�Ĳ�%<G<��8ԃ�,�Vް�����Q��ȳĽ?^�f��i���c2*��`�
��K*�z�	����i�u��+"���� ?�}0n�6�I�Y��,��G�zo����%��z�P0��A��~� K��v�.2r��mn�b�
�+�����w�ߠ̍��\;V�R� �"��������UR9�idu�����tpq���������߭'K(r6_r/� ��f�ʪ�{�;��Q��\7^�K��<y����e-������+�����3�$�*�LdpN���a��=�l��a����:}�k��:Z5,�P���f�j���{��u�:��`O'Z�AK��V	S#R0%4�6�/g��H�X(���v-������KA�^�T�����곮#9�_�r��Ff��@&TŪ��(�VvpNF�=m,u@�S�{O݊��%�Zr�U�k�� �RoQ�a�p9��p�Y=e���8r��"ga�������x��vw$�~�N�b6Zs���e�/��b\N槚ƴ��2h�� ��)[��f�zV��h�t&.���J:�EhZ���4W�b���L9ڞ!�a&���|$FL�v�=��@xB_��ʝ�+�b,��{��nW��qĚ*Z�Y���7r^vòKW���qa=�ß�@�S�g>2Ht8��^kk�!Jx�k��l%�}�?�Q�<�r����0�9q���;���rŀ ���Ŏ�}�ׂE	G�&�}��OE}L�����5V࠱̕`�݆`��z!�o��r�p�Q�M�T։U����~���t���Q7�����F�i=�\��KsH��ΰ����ј��!��v.3+�2f��8W����3x�4�Gr
�%
00e�� Er���UF���t)�o��,����[0�[iB|�uYOv�"���`�2�*#�C�FF�+ia�j�w���
�����/k��7�N9<�1x�V˞+�����.��go�C�?E��^;:�i`�a]zO����m�泐U�<�n+z�jM1x0NY��bE�F �8`��l5" �/땅t� G��ޛ�\T	H��n�6]V�|�F#J*ě���-�,{}�w��b �ؘQ�o�Qfs�N��4e^�戏��sմ#-7ύ�5�z��of�D��.*(#��}5�Y7�'�S?��ȟ`e&�s��ٮ#C�=R�vz�;%K0���%V��h9<}>�:�l^����C^ A�"�&����j��`�== QtN8�T����E���*q�x|b�n'���a
�߼Q������U��d��$�C �r�(]����H�ďJBF���5yc��m�������i
~��7Z��5��m�� %\�5t�ee;a��5��^�EU�h�-���6`�>W�9�8W�Y�|��1:k�����@=z[�Hi6�(+HL�1/�z�ǧt�X��ϟ�9����_�}$�^{F[u��[����W�&���T�N~EJ�k0�(Z�z����i[�HM�]�+��:伉�Jn�G%�S�R���ʋ�Q��U��jsny�";���k(���sǉ)��oJ�Fd��*�뭌��t��9��\o�� �Ϧ��0֔��)�5X���ƪJ�?�ϞC�x%���ҽ�Ӿ�?k�5G���g��6ر�5��VS���"�
wt}�3}�a>��û}bc�[ַ���ZԴ;mX��UN�Y��1�'�
?��ORt�2%c6<�O)�5��P����U�J���{J�~��F�r4���弁  ��, rD�VQ��`��ъ� �'r�b��ԣ:ϩ�xE�5S�����7G�Ā�A��%X�Q������
���=pk{j�i��
?��R>����eA�4"�
��{0�΍D�{z�Qrc��9f��ﯵ�V's�K�EE���M�>�(wDͯ��	
|0���w�/_�g���z�A2����-�M:h����G5.�C�Sn-���\u蝝�B8��Sh�r�n�D�XCq��:HE�zbID�'})�Q�g��&� �tL��ʉ԰m}�Tg��c�;@�zyy����Y��۝.�LMY��{f����u����T1�J<<�Y�8</b+��ˎ��������X�5�^��r +�|s�����-�&�G�@�0͍:�����m~���)�X��sĵ2Y�1�$�֮�X�~���Q�A���������d���i�2 �L��,{>Q�����|��=�fů��e�4���)�����a� e-\��3A�9I�m�%�����l��V���}�e�M��5ŵ�Y�ɨՂH���U�^���!
0�@�hc���?�.C��͵<��yM%�njģ���"�����%J���j�fT_�+:G��^<{���g��lԚ��pHԠ��0�*3�YKS"r F&K��Q�9�d�;Hm��;ӆQr{�A����F�������,�le��"�F�f�����Ƨ��w}�԰O3w�v���Uw"�/[ʹ�-WYQT�N�"A�2|b\�y� �ʞ6���\Zα����������&ؘ�a�JT�Q��\�ѫ� 4Y���%� ƻ�� �HVaL�3ڄ\MiaO�n��N/��V�l���:�a�{�5�:�Y�gn���`���� 臈V�ح��7*��d^��H����O�j<b������L}p�c��9;��hX.Ov���xh"v&wHA��«�j�&�r��� Nt�="ɍ�>�4X���5;˱�#=�d���R��'Z���ӽVSO���1��d�y��T>���B`��7�l(�ˎ������%A������I��9D���6$�K����G�+n���q`:V�Em!O� +�qO9���� �_�������[�'-TU*�-�sJ�J��	n�����-����~%�U��цe����k �J�l�^�j��3N�.5��h �����[q���Kp)�e��������r�T)�Ty��g�=z�sOY|�Ayȇ ^}��Y��@͗B;�?{eKeN�a�ƺ?�ȪKݹ��
�����ʰ��k�e�9rGǻ����jsD��+��� ����������m,�vD���=pbzt)�%�ɜ/*�="�Q�I�a�ߎ��jVh֎*�E��ʕ��fy$��Ih����&��R�=�3�,*GӧU_��E�Ѷ�«����^>#��:��&�t�bHcv���ƨ���)"ca4%]^v�?5J#�0�z�ʥs�Ƈ����~�ᨰ�X2�y�HcDv���W0��
�"��Dj��r;�;��G�V��F���b@RoΪh�H���̒�S��#���^ѹ�9�%�F��`��Q����S�έ��ʪo�=�۫�o�d}N� �fۙν1
��F��Ut����I�/<_y��gO.�~��Hq��S���'��s\w�+���'����U���P�#�)a�C���i����kE"�����24����5ʰ�m��Uрk'7�4�#w��>pB'����ùX��VA߫��@I���#A�M�e~���,Q�)�MT��#*z4��,x�,��d�!�c�)w���=��$L�\ܱ����=N �QJė��q'g�������م��L�H{J���,�tF����^�sę�4.��1{��)�!o�	����'�˶hx�-���aIS�d�����<�=�3�:(��N�|��X�� � <6]����n
�l��m%�77mB�q \�����^iĀ"j$�@�轤�j��ƩE��N�n���PF���`��E���:'n�j!��ial�> '�6+�N������#�ED���Tk��Q)X0�����q7��	�,
�C;��A���ڮ�2�,�)$�"q/H��K7
JH���-"��Q��i�xM�!1r��5�\�)H���=7c�`>)�
(n�ƻ���?��s�JI]R>�R�H��+���;��2�Z@��Z���[��5�*��� �k��U3z�*ga�P<0&���R�*��	�j��­�Kin��s�(aL��^�RH�������H�uLT�c>�vm��A���7O��Gk�6,Y�et��Lf�����0g�����f��N�p�)��_W��m5���쌞W�0#,e�Y񞟓�̈́���}c:�do���rt����=~L*�0>9��y�h��p��r�a�z�#:��.��3A�luyj��M1��*��j_u�8L�����w)@Q9ar�l`1%���A�2or쵚����!�uPY^��؜�P]C�a���q�E�Ҿ9���d.�0��y����H���*�N��Q���dA}�#����D���ʧ�0��b�a��G| ��,���k�TW2P�墷�*P~
3��ޛq���|��H�IZ�{X]��)�x�&괬"�  Ĕ�K��l��he�I�> v`�w��4KR�������0S���Tx��D��u%5z���+��D�����8oF��zN	��/w�j���F{�
#�,���dI��6EV��O�<���4)mkK�S��z�)T���8��m��p*o>>���Dn@������E��@y�܅間q�7��m�4h�IW�@�����*���2LX��$깧��ﶤ89]�6+�'_�J�NWI���ũ�t��ZZ{ao(�m4�ڋ���?���x���-��q��_��[�1t/D�x��e	��*���\���@� �=u��5�^�	�1*�Q�}�
(�ao�G�"u��L��	�Q���Q��3i5�Qs _����Ǜ�r��MS�	�i��y{�Q�cslM�zB��U�W�l �wI�h���VKm�E5$c��o�sJ�;�w5��6�D�,7]P?9M��;d�\\iF��;B��l���rqA���3��%�,��j�YC��������}z��j]��j?�9��n��WZ+ic���}����k�AFE�+;+%(��f�ĖӺX?h�T����jL�\!g��;�@���`�F_�W�'AQ���q�So�;E�XZ"4�n>�E� pɒVZiԨ"Sʻ�
zrI��3�x�-�#{�bzn�"Z-�����xZ6՛�G)��(�:#A00�w�V����,��f	c@A�]��|+�=��`R�!�:���`�~ް��_���j��C����l�[�Xȕg�>l�z�]�K$���l'af>}���((�T��vr/V=�C�� ߙ�&��ޒ���D� 3�c�92M=����8���Z��9΍ �C���[*Y���F��uٓ�X�@�V��y������P�\%�}ϊZ�U�47�М��f��G�H'�^h~�X��<b���z�ۇ<o���<�9'Q	�a��ѲRזBK#�|Ra�1.�e[��V}bBy %�c�.d��Yd����-�x����TyʿS��X�~s��+�k���h���`jF|j<*P穖�m�����r��RG��!�f\!s�DO������tgB����ԫV�[��5��r[Ѫ:j�z	hW�T�%c'��1�|�h��p]x�_�~##�d�LY~���F\2�j���K�g��A}��/oHG��=0%cmq�8�̱q��%�W���OΪo��t]���u�3�D���}������h0n���X��T�c၀����5��C�+rF>�"i�h�(oD�RIf5qq�:� >����K��A%"6vao��Si:噁c�7������4�)#t�y�n�WI���{�fD�MБ�bc/_����Lv�Q~����閣�R�ꪈJ�
��:�v���l�zB@j�E����^kխ�̤�=�J�;�<�J~�_R�]��iE/�,��苛�;��K/�Ĺe���s��T�3wF7�,�G�@�'����������-u���3����񨐳c+(�g�e��l�@8\W�Ω��}�2���٫��4�KV(���d:�ր���V����jݼh��(����ѫ�ʷ=��>ok՛Z _~<}�Z/�fK�e=6��*2�Hӳ�b%b�&V~Yu{/����h�:"���=X�X�a��ˊ����-R�g��!
=� �^��k���p`��a�,WZw�����Dͨ�ph�]���s�p+��w�m	������N9�]�|� b���J6V��No��N�Y��DNF3Y��^FIv ��>�зw��Z�*��39���|~*�S9I� ~�Hȍ�°��)�4C��	�|������6a�L�v�4{�;�����Z�_���Nzm��I���^�2,�[V�
���Zh7.�q ���Sc�O���� �Ї1�JZ8z��XA�V�����35���C
�fT�Y����A���V-�"��D��G����V��gpǻ����ǜ��p�#Gx�=Ev�,<ʆ_��z%�@�[J�45'����a9Y/kr:���h��r1�*�VҒ���H��8����P�7M78%Rz�=%��%���>���U��M��\�mR�@�ky����^�Y?��o��r/��Ejd������ �4|V�	5x���K;9��)���������;����Ɏ9�@n��s"�`d�;Q0�f������P��G)i��b�^��ڢޯ��Ƌq��p#�gcß�X�j'^����5Ri�.�rNC����:�|���j_�Y{����<�%A.��[�i-Ć�6?�h�r�8`Uq_����/i�����|�=P'��vL���?G�D��(��ٿG��ƽ�_p8�"�~!�%-�!�������gz
�)@N!��) �huTk܁p�{!�^�6ɗ�F����&����xM�A�6/{Xa�����R�<(*�]�
�#��1Yy���p4G����:8c_��x�ǧ��_s-�G��[��r�A��XO4Gg�W� a�*�C�Sw�R�b�#N������7��ںҮ��#�`�G����Q�ʻ�)�L^+�N���Q�F'sng��F� �j�r�؉JL�h�hd\:��㊑'^sG'�#W��[o�ʍ:�B�{��b�h��A#=�v��X��F5�Y���lsڙH�xd�T�#���#Z�ު`"�I+`v�H@G��1��R����YwF��Ϣ뢑�����ʲ��GK��=��V�B�=�,�r�C(� }n��zx�j\;�o��ME�a�L��*���I�s�_;+�����fgU�Z�)�����y�6�*/��A�il)�Z�l�E� @�+^]�+�*t7�ר��Ʌ�ir�iz�����/V,���j�U��@>���|��L���������U��˾�b.�Y�ce*���������G���˶�:��q+���*�i�b��bvi�*v��W�s,+
R�������<�V�o4m-�*f�kG�%5W���b�rF߀?��jR��!��F�+p�ޱ_Q�TpK�5��n	�ؑ�k4�B�؁S`�i���N�(Kȯ��6J�NR�fw�5�� �Sr�$]���Tڨ��"擹����U�W��r>=!?�*�f�� w>����|ڑ��3h��V�Y�PX����X�g![,4��"3�qP���4ۙ7��(���"h��`���t�hdg�SH��%���c��	lH�M��8WB�@�K��=$!}r��N%玡{����W��=6pDFt��4[�m1x�PI4=����^<_"D�8�D�vM�r���yYGK��_�Q'ih8`� �^Z��>6ЇQ>�U��h)�h��Z6��h���pC�JFB���Z���\��겄�v;��U&bte'���)  &m�\E%Yf	��H9X㉅���@7�^���y((�gi��N�fg}j�24�QdV�+vt��˶��z���g��dQ�e	E�W����Q>ƙ_��Q��TT!��Q�-׎����(R����
n�AC�j��WeΡ�J1�5O_�5F��W�9O�G��*�ʈ���5B�j�<�Ⱦ�QYQ@Du���x��O &_,'��տR�S��R��M��c@��])����??�/Scs�}��[5��G�qox-;�38���7�_uM�;�/�*<D��ӓS���O;l\�Қ�J�j�����^^]��w�Ǽ�Ǥ� �FJ��&���h�4	�{Wv���WohK���v�.�:'�w��W�ٜ���?A�;��x�R�!x�� ���ҎzFs���JG����s�Q����!\��)��H[���"[�*Gm��#}{è�.�l�L��Hzk��Ԭ����_:^2�
t�M��F���w��G�^�'a�	#Ju��Ũ8� ��b��>�U���³�cտ d��EP���3c��C���)�Kz��3jS�=j��c�SPGt����ײ�})�k��ݤ��xDU�YH�=�4
��Tt�m�?H�DL��z|����M��̯��L����@P�H��|C���>��J���� �����'��#�����Ľ���R���TV�IӨp��݃L�7�6�9�ej�c�s�hDP�����w�ucі-�>�I��/�H�3:��M��j8�L>���q��>b]��}��C���K�Ƒ�?����D��B�����91�}�9Q$���ZהHu"�1��ɶ��k�/2� ]a���^�\���#���Fq�T��g��Xc���zu�b���Ǩ5�b��F|�r^�NA�� ����y2����x
*�_#}u��H���t�v���h'�6gذ��q��!�: ��(? �a�����4g����&��a{!�/="q��̑�;��$Z�q�b����\N�y;�q��Z�;��͚� �b�֔�cG�o9FO*G�\qz�:y~a��E�����N��|���� �Y���������]KCHx�)9{%�3u9H|�Ye()��t��DT���\m�$%��HL���E9M���٣�mv�jX�h�\l����; ���4����CӪ�~�8	^$!�;��k����U!x���_��$KY�"���$
�h:��l�n�1�'�=C���E�XJV2hf��H�����X��U�P�p5ؙ>FE���z5�1�/�레��faϪ��x��
w���P��ϻ,��6F$�( v�������I~�m��̣����2�Q)o�[�=�N�Ȕ.D$�N#���>jE�`C^IK+-�b(�W~s#Q�&Ms�NB5�J�����l��0b��j;NZF/^��qV��"��*X�*5:����w4J��0��veMwF��?F��{$R(�A��|���p3+�
��d�����`�{�[G�;9*�.GƘ����㠎Ǖ���99��BT�u?�Q���DzUJ�����PߢC�Zf�-A��F��#q����(�9��������i�"(Le p�kD��*:/�̫WW��_rs+�������>��Z�
�hQe}i�:;��=������+���{�T%�o{��\殔)g2!zİ�>�/���ۯ=\t1)�u�ZM�urM�]t��}��;���������
N��q'z���<'��5V Gy��XM��q�����R�Ӽ�W�D�nG�b�U�z-��yJU��VZ!%(�oE�`�#���ۉW�z��thru�b^�;(�1��Ų�3���Z���+����h��#�m��	���қݫ��Jh6"�^F�^aO��"����PPf���"�Mɛ�J\�\�J��)��)�cjN��F	��{���T�z� |�u6[�W� 助{;�#V����KV��N����-TGI/T#�+8���6޴SMW�����M�kSUϦs���|�����n葟Ѷ�C{�E�>���f<�q�~%[�����SU��+/i|�Ǳ�Qq�=� ���C�Z}�@����<eܹf�T�oX�
L �yq�T���'Ѯ�g]����7�����+]��uP����^��A�Ӗg��G��&`zM�8��{�Ȓ1Ѣ�>?��&�Z
^�ņ���꒩[T�澠ߥ�0f�����18#�Rc�a1�]l#�5І���`�Ȍ`j�F�8�	}�L$fi$���2$�N�x>a�,P���(�ҳ/����9?=��$#&�1�Mv�f�\� wX�x� e�(rFe��j���2�D��l��w�b��bO3AU( ���G-)�p�pX
����Q)G�Y���葝�\�4=�ߪ�;�����a(�/�
��wU�!�#�و�AJ���9ӰF}���Ǣ��\NϿ���*K��ui�$L�Q��[]�U��
�9J����J4�d+���e(0L���%%�2c9/.��gB��A"ӅT����V +;�6���XYu3B:'#�Ԑ�\��˜�4��3ł�`���=qh�:r���ܪZ`�e�$����!�7�U�\��+
 JK`j��K�6��Dj�-�yv��MD7-���W�%��2p���6�#��9zZ +c<�t���P��H�w,��k��z!�i��lC1�4#�b(ザ��5���lkʦd����]�ڶ>OZBQ?�:�sX�;��J:�o�������@J�V��C�s���q窄]Ň��� K?�F1���R4�Hb���o�r4�"�\1��OKߪ��r���/�� 6_ZV��JR�)��sǌlnѫd2+�E�ƣ�u#+�i���^URu��+�#�1g�0!�X���J��)V,�<N��d��{�i
�������ɉ�����E���3�^!* �#ۍƻ&Y�dȽ���6��J�7������5���>Z���ZGUnP�Us�sj�'�/ia��+���򫍷���矸��/�G��y��K��t��"�u����\�ľ[�+��b���BM�"C|Z�%-�V��h���yqI]]�����-�(�8k�C����@��*��3t�WN*u�����sEu�m��{9Z8J��"T�����i,�C�Id�v��y��Y���Z�`"A�"���t�H���h��[�1�5��J/�x�2G�9[R��R�dH��Ę��c_�Qh���1;9�If��9U�)�r��ۮ�Ζ}Cd	B'�Zռ�ȕv���n�ӹ�T��Y�^��Z�:h{��^k�F���M�y�W�d	�$���ѮVl�X����0�;���!uգ�	��v9<<=��N���q-�d/ ���`"�ئ�R[�� ��I���%<���i!O������rB���q�f������[�m������J��$���y��"���e_����A�~��P��섫�4�]��k�����kc<�g%|�l��l�J�4��H9Gj���~Cg�M���#�D�m�(;P&L�S9����d�^3H9=lg�,AĊUǆ.B���a|n3�e�v�9=m ���<���C�����d�<F�N�����Ǔ� OL���Nr12��r��X���M96^R�=�S��c�U��.�/�@@qr����z�����,�>������.d���q��3Ƈ8���~!�q�56H6�G��7f4�W��GD����)2��6)��pC�-x@��C�G��B��vG �v�u�h�Ee��3��U���� u�ʪ�i��u��1O�P�f1 �)Fڌ��mG�e�0�Jvvy.��\KC���2�����4iN����\_����&!k�j�ë�L�R����rL��l�e��z�3��9(��}/���B�/E� �%4���_dJ4�[��U8p�@��=%�ҕFl[���6{�?g(�aU:K�R#GA����.����?��J���-J���:� K��<cn��Br�"Ū	����~�ؐ�!m��o��o��h��X��+0��~�^"�=[�RN��D�1	sgc#OU
e�0N����k�����mf~��3x��#_��MNt�B�����v+Q���㜎A�����mͣZ�}�vT�[��~*YhI�ȇ=G�}���Q�0�Ē��q�*$�9x�y�b��� ^ͦ�ٍMA��k�L(s�>�������s�-��>�j��k�??�7!����y�j�[I��=tX
���q���#\�}k{_h򫯼9Nd����VuG�J�E�y�e)�i�v��G&��h�6U��x���c/��ڂ|u
%h��h����s*xN(2��'��y��5�E�%���F�x��a��
KT
B��57O
����F5ʍ�^((�2:�}l�%�ߘ�K��3"���=��ß˶S��v�p�r���/ó>��;jKyϏ�g<qc��G֠�ƟX�9ut���|�߁�|A�h���N��[�,�\���#*k��T �s���"U � X�-���CJ����N���D�:�	��;� �h;��t�ܝ��滼�d=�s�6A��%��<2��七���^
�!XJ�_T��΍�k$�Z�b�;�7��R�/C[g��#�l�<�r��4vۣz��\�=��jZ�"Q������JXmfW�CϵXLƹA��iaSܵ��gC|�^�\u1F�A��X�������ac��n�x����B�J�d�CS.�?TΛX�V=�Z ��.��;���չ�/�x��+���~��� ղ~�����q�*�q
�ߕ��v�z���(�1��6�_�-�XZ��c����#7z֮
��뱨?�|5Y�:r��k~��=[3��b��)zS��?ѠO���K�Ţ��ǚs���4ʎΫhk��e��R��}7xF�T�X�e!�Ff�5�grzv��V�^]��ťQ{t�xx$q���=K���)�<A��dD�z� �(a��{ia��͈l������+r� Z�a��iZ�VL�Sg�H̖BF�s��["zf%�F)�}�k|��|���ެ�7��B6+��n�R�U{�5�q�����:�bO9wvzJ9��x���}�o�fq'+�@��`�Π��j#6>���*����[S�B�ߧ�b�G-Q8Ivvv!���t�Jqg���x�Z���p���K��ܸ��4�79�ڐ	Y�n����^r���四�A�X��w�s����o��:�<)��
�L�o���L�I�A��,uǕA  ��IDAT�j�2�ʣ���m�t���
���Xkz�9�:������<+���ٓ�ڸ��=����2�=¥V��M��,M��s��4b��K�����:����2B�%}i���3Ż��~_�I����P%���Ex��}�)�}Q����R�
pv3E��"p�7��	����r���8W([���h��p���ƙOa4C�����:w;G�⟍a(L�C�]��X�7�A �s�%�R������"@'xt�)a�RW���l���#ꋺ��C}���7=\�Đ�<�b���V� w�ѣݬ���U���t�z2G�`������7ۧ��ט���݃���w�v��V��L�ѣv�"���{wʊq�D\8S��'M�FAH'5�v����Ȯ��"��\Nb�����n��D��:��խl�eD�hD���XA4�xl@�z���7��7
�E/7Ȕ�XA$�rA��O?��{����ʜ�-q��I[���@�ʀ�"�m_CDP0y������jtc��]���0p2��<����8�r����������|�	���
Kf`^XG���_(H�)�Оb�y����v�	��(+����ݫD�V�:��L/�����ƣ����Q�ˆ���8ڨ4.��l�Ÿ�Y��^��9�Z�,�D�.Qr�!�����ҹ���-�����m��l����S:T򂪌������>����/J?u��+�� J%�t*��6Rߥ��ۘ#��_�P�YL���;\��Pݻ~�õTu�^�+�S�H	�(O����\~�3:�q����9��t�:�<��j�j��YYn{kTQ�;��_�d�)ܦ��ܴ�U��qo��@�H�?+���,�O��S�u�ݨ��s���L�W����'02ٲ���/]�����f��XKb���1�^�iU��jN���T޼~'߿�^�^]��@�H���A��R_������[�����1�� f���B�RF��C�?n-�[k��h&��_���#�] �?\`��*��(��H��9��/�uj�w���I�[l�j~.oί�$�����}/.��_��_���([�u�O�'F�l�-i�Ͽ����W�r~v.'I�����u��������{���fEK��>����K�)�NJm��c�e�1�sm���d���덬Ҝ�d6����(��_x���PY��������\���������5�����zw*(D';���FE%V�Y�S��y,۷�٦ie�#��,�:K���,D�게r���p}+���ի�����4�����k�2iF��;��%{Y<�x/u�F�V�����W���V�ˠ <���G�%em���=<�W��o�#�v]&�� 9�T+,�W�eb��P���u��rd�V����Y�q �(�M�M�8�=�x�Ddȯ���-]R�u��'�{KX��Y�upGvj�U\ў�=�h+L囹�`B����"fzE�2!�{I��*�4�	�Q�%B�"~B�l!�Q>�<Ƣ�3��[�r�B�����m�R��͑�@`�v����R��G0�s�� ��iR#��<��=�<���H�Z��;z��K�<��(����w��������L��rz:�����:gA�p� w�w��%�d������$�3�)��7{�CO�'�Z)�7�zIQ\���a���g��h��=���-���t��P��.�t%C���)�Uo����qQ�A��~xg&[pOuH������(eu���z4"\�ij,��D��B[��L���pHs	׸~|Ԓ��<X;��#DY׎��A��<)9q�G`��prS������c�ZT�����A��ߕ�{�1 0'�a���\.��|������g@7��}��:�>g�<s��}�7��ƈ��A�H̉.0�S�8����m��,!ŢwJ���g�a�!��:��y�����������
��F�<|��&���]�3����mq�YU��'Q|vV�s4��Q����4� %�п�'u�q{�Yꐏ�͉��+�ke�������{R?�w������(�
��]���3�9y���R�9�,�I�G��c���� ��t�����rK��$��K~�|��n�Mq J�/�Ǟ�FzM�� �����m���m6�s##�g�j�r.���U��h����ߝ�~���&����h1��#g_�^�;?�}'~�۾�|Cݿ��,)W/��G6���1 ]�Iz��g��ӟ�$��?�oy�浼y�&�@?~�ۛ[�&������ ��x���,Ӥ�|��H��iP�{[1y��	���E����Iyu~!�������t6��ۏ��צ�E�v�c�����E��������2�Ӟ��Ez-�Og�X%]���W��/�������UF��|b��R��_�U�Ͽ��ӏ�?��G���w��F*��\�<������I~��^��X5�`����̽F�-�O�⍜xM+����i�k�c�x	ON���s��r��;$/i�\�]������v�!A�4��l<�~�e������O��.])+�� q���ۻy��gy��Q�Fdr2��5Me�(�����F1}��F��ӫ��Rn�$�XJ��������84�S�p�� I�%%x�&"�z����t�ki�{-�Χ.��0�7�%WDB�'dm�=�-x:�d�h�B�M�o��ƕ�z��v�-�����)֖z*�-�)���)��R�G�M��Yؿ+D��6ؿ�3S_�������Ȟ_,��	����}��߃Ѩ:��kɍ>�H(<L���������i\�Fy�oM��-o�@�7� ��(�!D߄�QÜ[�,M���'�`�Ol�[۔�4���ȑ�09�R"v SRLMO*�]�f+�_�+�y
��]'��axhQ�@:�l~���ryy��'�|V�DzE�
W�(.g�+�=y��+}�F�T
�o��f�-;�f����R�'X�����>y����3��1H�
v�N%b)o��pY�WơI��k~0�*༴�D<���
  #;�|4���̆��$NɵK�R'��rR,�2��/r�q��c�x�\mt?�ڵ9����麻E��ٸ&A�U���G�����f�!�:�L&w��53R�����!ǎ#v��g�ՇǷ2�^ڊ��`;�[��F����`~�3��`��Y'��g����vļ��	w���ΪK�����G�˲��$��E+<`��O#AT񴉧�x:��I���z�����yjn��dZ��O8l<U�i���):{�!�o���ᘅ�(oD��P'��h��Q��c�j��jR0�� �e�#��o�����p�G6��녁�Q��li]-�_u�D��#/k{�Yb����;��<�B�=�I�}����]�������7��ySf��͟��\�4�zO�m�o����g�7�j,^���h�*�ww�����,2�p`�>��c֐�Q�Vlh~z*W����Hc����Y'���������J�W��}�V���H�~��2��r��jG =k�Z���ͽr�%;I1J����.�_��b&w����S�����6?*)N!���ZY�y�@xL�Ӗ�`j�!	0��|��d&���r�,��: �N�sF��7h��ᤗN����pC���ʉM�&/Zç�G?:Fm���SC�3�I��䦇��S���Rtvr�:~$w�;���s��!��|*�����Y(�;�s�L%�Ω���	
�Z�H����
�6=�O����_���Fn��Oiu�!�K��,��@,��Qd�?_1lG� ڷ�X�e������qc e��s�߁ �o���6����O��'Bˑ� /���(Y�P�nq��׫���C����q���9K��RR��?�"H��n�3��������TN���=��5�g��ң (�ƪc�3��}��0>��x�R��b�Ƽy��A��E7�hFL_��[ǬD�c�q,PS��R��x�8��Z٣ϓU%̱�Fs6�n�L��(�]uH,�{:��L�r��0�F�� S�f��yO��	Y@�ZU�\(��}W�(̲��n���8��Jf�*5�]��6}c��l !q\���ȸӓ����%�	`��
�x���8}�UOt��36nTQpk$�;��:��à�U�����o��Oq`tϼQc���R�ܞ�@�Z�z�"�zV�#�K���T�[��1rP_�qpD(�я��@*cٞ����;1�}���g�D�-@�9S��bc�.���������gN�i�Y&�ƯmA�Ζ��Pk���uR&:�P�g�^���](�Ūh� ˑb���(��^��o��Ú#Q�/=\{�/T��#��~�8�m���R���!1����eKV�2RnQ��L\OQ�b��'�\���VG6�Z��F�ȵO�`_˃5]�k��i�jp���bm�i�baQ����C'��:/���g�k*{��W"y}�_y��Y�3'����&�^��Z���6� T�=ȶ~��9Xdu���/Y��l��3�I�����|����. ����ÁEUg=��j�OCoC�rc���?��#�U|y��e���݈G��=���"c��Mۆ,?�¦���N��y~��W*1_�����L.���z��%-�n�ޕ?gO��d���j���s�s��v�dّKz5�,k�H��4龯_����'�so<:��_�?�����ײH�A��yu}���v�����t��2���ѱ�p��樤�)�7�5BP+���>��r�}�Kj�߿��������/2k&2���s*'I?�^g����n�K���N��)DR3,���ɩ�C�Oz���<ggZ�|:���!��I��q-��N�Av�*�[�3�)#5��lȫ3)�k��d4�\�<�@�� |~{/?\�����1�&)��V�jЍ&�@w7�
&��!bg6;մ�i�vgU�@����R����<�^����-��]�1�=]���Q&�O�:T���`\#��a�j50�>̀��*I��>O}ujn��3ϰ�l905�qL0��R��GM|c��#��=ک^�N�[�p�PmPxU�B����&�TU��[NmQ|z#�N�}���p�Δ,��Y�(�Z�~Th.�bp�
�ZhGO�Yq�!���ty�jrM�r� B]��}kRU�Q+�i�N���\�ݮ���^�P'�n�J��_����<�e��V�xU�GS��Ӊ��2�tfp4���^U#�Pp����Q&b��#��C��I��<bs��sW̰h�)���e��'�|��$3g��:���?�@���Eg�
�D�$���5�Lt/����̥���N��ז�.Sc����O��/<�"wjȤ�4�}F9�pC�7P3�[�訵�9��d6S�a�(�M�f�8�Z8_zk�s`���]?���Mz�$����.�FL��}9��CNw��Gj�WS���*��ەe#�"x��G^C���`'2W�E�% �t3s�6Ƒ�	���x�����ZQHaJN�Q�9��{B���b��,�C	҈����]�G�y�k��y�	�����*N�]�c���Ouyԕ�zl.����|���b�~w[�(;��n�*e��K�:D��s��kYf��@#�.��mbk�8�==�"QF�u�ED|\�|?�;��PmjZ����gç�cW�;oةT��̆g���k�L���ֺkH��_��N=�5�#q����)vN�����[
#�Ĩb�h��DMaa�`�}Ws1������=z��p�����G/o��ޗ'�'����p��m}~0K�Za0���~��A���K���!�/����/?�58t��^���Y�6�?� ��}G���x̪հ�u����ziQ�J�������Y��"NmE��5H���9�Q9�$KzK��exz����\�\�ե���(��2}��斑B�+�����}���w*�������>п(P�jʩY������_.����ފ� �B����A���D	�[+����|�WP�H��w�$t3�a�0��ɠ<���ˇ��/�|AY��bE�f�ƏE>����p����yj�f�4��j�F��IL�P:K���O�g'���*�C_q��q�Cu柨'qV:���-� �W��O*r�F�VB��P���Q�d|.��Y�'�U����e�B�mT����tQ*$��= ��:��%cVz�Z�O���e�]y��6�SR��Pd�TW蕣A�F=GI���rt�'GO9(����H�,^�ב��G#f@А��}Y�T5���^2��ލ}�+#9ڳ��XG�8�2{�IRp�jSa��bJ��&��O�rf��_v�R9!�/>���}�U��ϲ���X�J�Y��_1\,�7�p\o�ֆ�6t��iG���H|vE�˽�o��N�P�1E6�';���ho2�҇�c\|Q���~.��
J�o�DՆ�d��.ͫ�U��'39?;e���ى�̧6���|rB�~��\��W��������#ՓB}�����A�|�3�K�x�*<}n��J~`1ܰ^�xWL|�@�-җ�F�UismV �U�%�l=D�xŘ�a�ȏ�HAW J)e��A4[�R��Sq`|+Y�ĢYA�e)�X_$I6`�1`m�J\���}�1>���tB�ȁhx��W��e�8�N�G�X�{�9��ս�����z��P�i�{���l+��.^r�'�s;�;���'�ҏ>n����JNTc�������Y���Y�	���C��J����
�ʎ*F�m5�>('�W���W��g`��������VD�}��k9\�I��N~��T=�k$�{��&j쳏g�68PG��h��x缮e0>{��W���@{/<qʧ@_#��ɲ,h�R��^�����2���6��i㱼\�������#�\���0R۴/��Q!�Gu7::Mq�H���o�_k����lh��`ГGK�s:+�v3������/�%׆VR����~cv^g`����A@����/��,7�7�X>���ӳ �@79����gg�����e>y����W�!��B2��p�i��ӃW��@��g,��f�\�f����3t�]�w��d��{�N'����K�h������o�����z%߉R] "�w�$�b�Ng�<J^�^m�&*�2���I�WK�M��F5ӭ�\���[:Yd�n\��D�Մd�k�����C�7*V�V��4(�A�D8�z��1�NGܬ:��z#w��D�.^��f2J�$�����=C��P�2$ߛ%�g<3� �.__��͇t�i�ٚ��;�p��H�EhYIo���@�9$�{v�J.._��W�d>=���BX���y�('2n��}�&�$�w��n�"�K�([S��:Ŷ�ʓQW���T��>gU��������VO�R�Y	M�+�<M`�N�*��������!$­�"=�I��+���P���p�8�8�Ֆ�u�ev��vY�6!}��u�|L�U�� E�a*��|: ѶR����dri_��� �b��y���3�H�7���F��M=�KəŌؘ��*�$ܩ��c L�,%Zڕ����<�G��X�����BYs^��S��n�L=
]��ν�Z�]�[O��w�qש��;���/>b�|ֆ��ʁ%u� d��$��$����0鸢k&@��|[���h��5X��7� os�[�	�s�=��7O�8�O�O�Lp�-Ao[��X�/��ȼJ�ȧ��~O��R�R�V��y���p�e�M� �3���� �+���{%�FKlƐebo�.�j��l�h��1�ֹ��ӛ��9���(g�J/�X������n�)*�l8w��h�m�Q��yge=7(� N���}�����N�T���t����vg��'��
T��Ze��Gyt')sG�K�Y����)ѝ4%���:����s���;9��f@����Z�k�Zguſ��1�ƣ7L+����J���9@̹7�(nJ1n%��l���2�{��ڈ��f����(�=���Gl��vN����pПa�u
֗�9�z���zW5�S×y����XD������~�3�)���:F�����tо�&ė��`�����%we9>��j���L3��*�J#�i�+r�ؿ����9G��yZ#<{/O��J�x�V]��|��k8�Gɐ��9��O<>,Ԇk��F�;�J!@�A����q�$�����Vk�~���Qc^~UV�2�Ce	Y��=~�v{�Y�T� >�{�������+�E��M��C��`�
���c�S�qy����>?&��P�
���gH}���9fS��n%�d<�R�����{�NfI����ۤmhs�O?��V����
Z�� *�5G ���G[�:ǒ������X<�J�u*ۥ/��N�q�L:���l�u7K�}�#ȉ>zL�UPG2AD4uȖ��|��{w+�Œ�>���|�HtO�n����3Y��u��"���-B$vy�ߟu��a��nc$�uh@�T� H�Z/��z�F�5[C���D������&%���L���@����{V�B���vf'3�3���I,��������vliRjl]������Q�1��
f0z��&�f������圡S��d���Z���J�S{�#7j�I�%cl9JJo��v$w�N��+i�@�ra��c����⦆Q6t�p��"&PT���,�C��[�-7=��|Bƽ�Ih[��r��'z�'�E҈��)�B�w�ޱ�]��,��)x�5���)��QW��)HVo�J�@�Ģ�J�E�P��֌cx���UY�z��:=��EC��u�Xy����-�g���Y)͗��������ѵ�#�����+��w��P&`���ܟ+��U0ƭ�]�/F�� ��ʾ{%-�!�ec��������J�^�r��f�²�-wM�||K�R���QU�Ş{��*G�ų��f1S�O�]O��@K���̦��S��H���&����b=�A�x��K�V����>w�O�l��w)y����YzxY��醦���Y��(_f ;4�{̾�:�J���h4@1���4
g�6�q�`�;c����buR�q:�p	��I���0�q�+��e���h,��W�K��j�����3=.93�؞�v�6<.9��w�k-*�%Y���"�P����ϩ������7���(V��� � |"p`��hocr%ZJ42�hÈ�c� =К��(���;}eLz�y�+܅#o<ip}�(Q������ܴyJf��d�HI���Us�e�1��M�,���m�co��n��Y<�s�ϟܠ�nx귛r'�P��=�=TĀ��k���q�����)뛡�I�����8X��`��2���c?ծ���WN�'U�4�������,���ӱ3=ҝ����� v�!����w�z�O�}�������z88��ub���O��Z����u�����)�1�Q~H���\޾{�����̜3TI�[����m���+�oډ��Hѓ��h��|��O����n{�~�+���Y=�Y�m�ۇ������݁�}B���������e��������M9�<��r�����F#���,��&ȆtM�� �39�(D*���]���ԛp)`B���兜��d.��Y�%�v&�t{��V՘�Eu�#Y&;�O'i�/K��t�ņ�Xqe�t���ײ@�ʮ�9
����=ޓ�ϹH�#p��h{��NY����N�������)Ȁ"���KV+��P�<�����
 �X$\h�#�n��x�y��cT�PL�P��q�;)f�W## �a��*J�;=��ś�d�lb��/?�_���e�}��,RG��5��a�yw&#�MO�pec�Bz���"|}���YMd-㮓�t2�q���~��G����ݻ?$�lNd�D�� ��Z����]/�oY��7���p4hR�iP���:7݁���"��3����/��/���u �ڜE���y��_�G�M*�X-E�|��A����U6��~�z�n��<�}�r��,#�4�(ۜbJS���5�O���9ɕ+�X��?N�\���1n�>�����MX�:Wd�*V���9n��8(�,Əe��q�E^��Ix��̉E����,���r��<����D�"�l���`�z~[��/G�1\��eۺuL�MՀ�|�%��+͖�7J}]d �9���<��ɥ4�'ذ 4
�n�Vh${wq>g��ң���~M&�-8����_�/qߠ�=��}�����q=��1�J�4i4*�I{���}c���*��%�D	X�<.N.��Ɯ��M���������YR�'�Y �5�m�����m�~�3�"D�	*�%y�D�:������i�8Q���˔����
ҦG^�n�3LY�2^�\���n�y��r�p��$Y����Z(�G�V52�|�_6gT� �@��>�h�F��g6{����3�Ͼ��H�#�_���<�QZ����;|���}\��������%*���֟GoU�\�=E��h��與V�BbP�ʳ�Ѧ q�N4Jg6i��l:������Z��ހ����L����Ƣ<T�/:\ϭ􃇪����
 :~�>�`u��Uh՞�\^�ށ=�K����یi�o��jў���9_ �� B&hX��L����Ha����?�۫+r�|��w��'�B���� �]���Z��Q�z����s�P�i5K�vH�z9�v��Aj���욤'���e�+dM��+) #�%�>"wa�UJ{�b��N������ܧ��\_�׍��\�r����Y�/$L���)[ӹ���~Ikö�{��ϖ��!�ڟd�q{5�@����V=z��j�zzh� h���(X1�ěW���=Ð>||/���d~>��ٜ�����[	���Z/���k�*!���aXnDj�M��U�ı�_ي��:�@�K֚���$��}/�����dяK�=�Ȏ��<C��,�4p�|Ǆ�>��:��*Hhc���!Zk����zZ��Ĳ���C�i�AzJVِ�J*'un�K3�{���w�3W�����#���{;o8a��S��y�&o�QØ�B���}$hyo/ӭm�s�A��a��.��{U��DOuK2��ȏCS�#�e�D����M �U�=��y	<'��D�:皾-n��:�}㈮;�մ��������K>����4Ը+��ۮ���r��֞I+mUsĔrm<�� ����;������5�X+��'�,w	���r !	(D��J�#�4Vl��"����y\�pu���!X�XE�����T�:����y�c�_��N�I��
XZ2��71DF�`����qtN�S'䂚b�n9z��N6<m}�<n-B��I�䕐#fp(/��x
D�ى��<�F�K�F�w���鬳vF��c%���%g��!im���]�1-���c����dvN��}Z	2ec�J�����8��P��#��t������*;�*C����=[���@۷ԩW���M��ՆJ���PJ���S��~��k�S�N�M_�Ixu�U%~х]9��Lw;|�
 �>+�(�������k9b�f�����L�A�\��>���+p�LvF�sR�ɗ�SY�����YUI��s����'#u�g�]3����r���u,ͯ�k�H?䈨�
��%�6eM���_�"O)���Ǳv�ޓ;RӦ�B��R�@%)��t�~���l&D�o�+�������@�?��l~*�o�?�t��a|I������ u`�h�U 6`��6j۫-ӷ�U:"G!"�������dBZ�$l�:7@�p�1]���D-��{R;>�\�Ǐ�r{{�^7r}�Q�����5W���\���ř�����k:N6��� ���u�+'P�}>��3��ؘ�&���3����*���n�$���������
=×X�,I�I8�Fm�(dÙci(� �Ԓ�{J|��췵\�9y��M?!��-ѹQ3�W�_˟~������m�8x�z��������i`�ӥ�u��,QV[5�|�=�WB�h-`�P�G<������|��yWtn�h�{�)G7L��ܳ�n��s��������(����>z( �~=����T��W��f��\Q�T�����]��<U1�.���:ܐ���{�Q`��;Y��j��!`���W�^Ʋ�, `�sT�#�9"H�`�ֱ2x���p��n��y���∖���e�)}���r��Q��:��V6��7��=.������Q]��_�8��.�Q�E1�,˖��G�~uz67�&	�h�md��iY*�V������8�4$KǼm���R������1�B6�gT�����h�cr�Å��i�Z����)�hx7�uCE��(����i/�5ơ5N�l����m�m���e�=HI�= ������
 ����7z=���\�;��f)a���3�a�g7����x�@�@�oM'���Ŕ-�G7:7_�����伆�Eb��+�vG�ƽ���1���e@׫�an~T�ZW���?��4�����1�fd�����*z�O�Nc�����k�B���Y�|���^�[ G��#���#�1�E~t���W��1�s4�q�wz����Zo<����u����a����{��{�6бc������N-X�(����i��8�r���Q��j�Λ�=k����lJE?h��Oy��:4>~�(��H��Ժ���QJD��7��vk����ܓO}��6"�������Yl��:��h��pVC�@$
�1(%$h1#�Q26���d������F��EK��c��ﾗW���y��A"����$��9���X�R�)�����r%"ϤQZ�$�Ů<o�}���,�A��-"~p8� ��fߠ�N����/���Ǐr{�@�9���<��R�h���i����by���@�Ӵ�P.8Ȓ�@l�꟢���2
��7h%>�׳�v T(�w��ك3�k�<T�v��5�z��N�� !�8�8�䜎�WG�s̰�o-���Q�gr ��?�	%WT�?h�1S��^_ɟ���ț�7��Ax!rI?��A~��g���{���A�;ms���"�s�^^e�i�ZxF]�ʛ��
����
Z���S������M�G�-As ܴ+"2+���;����_0�a^�W���J����{���AQ�۫�f3$����ٵk��K�aYdo������3����Y$@���xc�(g�=���Ӌ3�&����*��_#V~�J�@E)���Z:���jFn��"�Ƶ��|�l��=G�H�K�ƾ���*3�2�qs+c2#�F}�\��Y�:�����F�K3���B�8Ӏ�l]ǂ��D�|l�v�~ľOK{���fV�Z�c�����^��ng��Mbc��P͌�{�sk� ��Q-r%JW���P~�&?{��^�[6�NPß�(����[�Fո��h�i|�Vܔ���15e&j]��E��v`G;/�Ti �ɣ�{�ÁP1'5�K'0$����;�ĬAvZ��D�"9��I�M�Xu��=�%D��n�ˎ��ֺ{���0�-ˀ��Z�S쓶>&1t�XU����M�I]^^Ȼ���Օ��=3���,�����YVi�������|���6���y+��l`/_A/_�Q����Ϯ..(�g	e�xb_���'Ͱ�%_o����?�E����U������X>]8�+��y����'>J�"���-�+���۞�a���um[���3;��L1�;���Zx�5w,^{������~�#���w}�{�}�;>{����WK��d8�<���~=��R�i>�I2?WZ/N���_�����x���'L,���w�"b9���y��A�|���E��j9#��R1f��E�:�7�u�o��z[�`*8�|r
�ܨ��1�y��b���������g@��:���©M��ɜ 9�w���x��m=���o<DT)�`qe@��>�I���RaHK��a'��X�c�쓏r�����gj���%� ]�.�e�5���$c@�ݹ;��8B�Yh�6��k�ܞ������Rl��_����g����Lh�J�w������<�d1�N�� �@n����{&�6 }vrH~�q/t�L�����`�h�����W�W篗�6�[�e b(XGAIS����q̩���F��pjO}�1��,݂�i�P;h��Ɖ�J�i��8x�8�r�\fu5'���'��Yҁ��Q���CקO���'����/?�"t9l�7 �I5
�NK�ڸ�]v-rG�<�2w򯼾��~푍wt�ɐ�Ck%Fsjzt*��uBF#���M���%c��cn��*[憻2g�Y�y0h�7���������������N�c>�6kJ�hU���>hW"�mg-hbٍ�,�Hƅwz���hT7�r�5�X���5�.\S�@'�Ɂ� �4?���G��*Q���ӱ��@��'4�!�},s3�6ذ��qyue��(���<��	pp����.ק�l�훱V�p1O�wR�W;�'�Q��9���G�R(P!���O����K�s+w��4���*W�v�7�7�����o��Y�?���6�c̛y��Q�Ψ,�1�L�S�r��<2�s~�N^�:aQr'$���w�n'�6�	e� L����1ݧ��H�񟑮;�-�-��b�r@��8��� Ӗ� �8vo��ʼ<+�;�@5����o��N�i�]f⤳�+�vZ=5y� $g�ɽ�����g�����T/�e��.8CQ&�!�u�@3�o،��m$ôu����E:�~�#z�ٿh��o��)e�57��Cų�e��'��F,g�Q�(7���D��W\��sӛ��7���jZp�]��@�~[5����bv�^"}%��'���_O�[9���8	�˿����W�%����G�����"�`ə�����F��00�)&{~���jlJ�ޘ�~����\�����W����cy�1���F׿�[99�s�e����Z�`�������:3��Ľ5�k�Q����*�G�؇T�v8�S��ξ���Ӆ���ux�5�Q��=�e_����3��=	T2�%�|��_��.�g ?��B��	��_��i]�3?^�6j6k�o��;�y;g�O��2c0�|H~W8��Pf��u�\��(i���}2ؗ�~��FhhԦx���� ع�f/��Z�8>�ya�F�`:hd�lP�����������|�C��}z�U��`ܠ�GM��v��}��4��@z�i�,�?S/MR�,�w5��t(����&YNi]Q�6�>�a˪GgzJ9l��Yei�d���Cc�+բ�V��kP�eQkK0u6q� [��A� �r�z���pr�cW�"��A��z����ʥO���P�G0� v���앮k�?��4�����_u~��?Չ��>'{���7��3�� ~/9[V��LA���AM�(N�ѫF�͆љO�Ȥ��)H��
7Dr�D�e����4��4�N��̮�1/^?aB���<�Z*��hjv�� &��q�ϙP���d��0u�it�ic'���]�x"�d)���	!H��L�"yn�&����0�U)��>Kgn�˅Ȳ
�z�1e���T�)�{q�bЉ�B	�l �H�ӥ8Hجq� Y��kK��XT?հ=_������^k��� ������ܲ�M�#��V�x�w���:����	[��
�N̿�����	Pp��6��ٞln>/E2�o���Ys���2ڃ���r� ���:D�U0c�k�H�ۖ6���͵��՘bU�����`@kY{ʓ'f�w8G8�j�q^~��y�<�ܫ`A�ěx�����|ߢU�z�)����5 d��1���;)`^Js��,V #G-��g5!���ѳ�#�����;^T/Z"̜���K�H�o�N`ǇĺI�Qx~~�{@Y.��m�g���S���	�>�^�m�s]��KP5{�/|t��l�hv��&��M�tq,'�\<}�޸�?2���P��9(��G,�w<�qt�G��,~��;�&��$X�FL��b�~�r��N�"�{k��WG���9���k2O���`�+�%��X����).��
���jY�ϿZ#�ֹ��]��(e^��縭��|fy�91�ꨇ������`�=N��� �<��{�3U�챕uF��F���M��5+^~�S<-5�1>����W8���m�L0T������d=�գJh� �u���üU�&�.Oנ�A����ګ`Є\7C�Ւ5 `ga�k�!���VR�d��]3a����+�H$���3:��M7�3Wl=�W�2\���+,���o~��oN�����lNe�	�c�R��%ӓ�ɱ��ɒ9s2�̠q(s��k���[�\_m>��4]�Q̠����%ܭi����Au(q0��`�alv&��<>=0�5P�砭��gn��	�[(d��,;�*� 1*�����f�R+��ĺ����9j\CV�n��3�����b�J�p�`�Rl��߰::~�G[����0WBHߧ5٣4��g0���E�ڌ�š�*6��u9?/;�qZ�Y�#�C�;L�N0�h0lЊT�a�c��V9�B�]5��Lf!yi�g�\�no�����f��>�6�Jd�ʛ5ʯ�X-Y?�e�y�}r,�l0|S{95=��*��B��&��Կ!�<2��2����g����ml����`̍q �Ͷ��)��èm��,��;����S��G�����mL�z��ɨ2��<lh��!�/�xz|J���1�Z"�:-��`@,ܣ��D@��{؃6����[��[��4��>�:j��``����V"V|Q�cO'y�*k��~�;�*H
#�se�l��L
X��I����D�s�ձ{M�=jt�0��a<���fCj� uv�3��l�M���iM ���|�kl�>�]h �!L�����ۻk^*��3��=��
+� @��}Y�}���w�ܾg�q��k hts{)o�\p����%�y��Q5}2�f�M����zd P���"��=� i����޿���� s�4�e�2���_�f]�'p���/���G���	� A�b���2�@��,F�5��,Ӆ�؛+�DBP��ټ1V4V\a�)����g����𔾧1gj�T�%cL�nJ~6������Q=7 �QӃ����oWӄ�=�^>ݢ���u ��j����o]C,l[��6���j��1H���tn���
* �3Ճ��gqƢ��=����0�z��
j���Pg.��%�"w�\��_�	�Ur�U3���P`�M樍��L�!٥�N�w�X��`�A&;QK?���d=+_�G��\�<�����M��F�^ژ[�h�;{犢�¥T虯:p/�^T��_�8��~�#��Ni�����c^����Y&�zv���S��i�;���|B9�~čK8��iM
XY ��)����A(�����':�-�+���دq}�S��2�r�'�A�S�) J0M=���w9�^]]G�e0֮��Y=;�y�h���r��f8>����5>�J_��{(c�����2tS/�W9�p���ğ�f	��c�sF���<�lz���X2:g��Q�nc,���/���]�b~��^����[̮�o����ߗ`�ߟ}��K��VYՁ���T^��Ѓn��=Vm�m�f���|WL�j�l?�p��zߋ>>���_�4��`3x���uٰ�s����ˋ����867�{�#�(׏�mf�{6�N�3�t|buN������(��'��+n�����U�Tm
���zͪ{EA�@���D�#�6���(œ�5*,3crG/��l�5i>踖B�b�}Z8K����K�|m\O�b���	��*���鱭\UK�{��s0$�7�!������E�5���������e'�~:O���N$�%�'=uq�޾eKt 8�� ���"h%~�X�9�4e�0�M�7`Ĉ	d1����@��J�B�o�A�.G|w�k�FP �Ā��FZGC?I��{z-�2��'�i����Hִ�;�����.���Fk^ä���3a��L;�65�<�c+��И�4����G�l���X��d���3K�0�8nz}��;<���3���Y_�e��xd2 ��]���u��;���n_i/��\^ЧE���J�M�k��y��Ϗ����gNL�^z"���"�!oM���I8��n�lk^�Kt:�tq�[��q���7��,-Qt�b/�Y^,ܿ�K���`)>9�	kn�,k(���DG�
��ALv�V�|C)�SP�N�h����g����v�����T��H��h�;C�1r�����i��9���Y]�:_j{i��3A.�n7-;����h���9%�m|T+׏@~���s��D:j�6�	u`g�n�����4v7|^���ml� 1����Or����K�*(w�@�����{��n�-9�`f�{Ϭ&���9 N�4��4��1��!:�2�����y2��t���\Y���uZ���u<��Q�Nvq�dyn�d� ���=�p�%J/5�:���'��1���e��� P���8�
�|ڟ���E�˝��@�9�Q�&�I�+�n���B�p�AT��`�h������o�ln�c�Oc��a�i�K��M8� s�$tu�4ʶ��T��Ű��a:3p'������Ē���o��IFVX��4�kٿ��Z~�k���x��߫�{���nLn.�� ��v�N	v� ��Z��N\���
��&��a�- ����2���c��(}	R���c�����1;�xh�g���n!ƽ��8$���Z�5����D��A��Q��y�5�L�{�m����w�=����i�A�������:wN�`]�*��Y �Z�B>��OΡatf�dp.O>)������ ��I��[^|I����]9@�9����-u�4��(��|.���:u��{C5~n[Δ��NƲhŝ�W��lw�s��Z���� �ܷ��_�=aY�~�g��3P�4�UP\�p�H���� �|?Ғ�FJ;K��E-�{�z�Ύ��z��������r��xe�3+8�=���
�;wP��S0Ʉ���ՠ����q����]lm�c�VL��ʠ�9���~�ͼ���he�#�b0�Fi���b�=Ѕ�� ��
rk��uOD�Jm��s'q�Vc P�'�1��B�h{��@�SN0fJP�t��V:/���,�������'_ė/8k2wʬ5���Ӈ�-e��ԌT{9��!����YL���`��bF��Ab��*�3r0�Y�d�v:Y#0�t>y7Y��� �e�f�2��*�w��g��P��i��	ټg�[-��^�[}v�G��'o��^z�P��l�	��F��*��Mln��Ox����
#O�u='b���zOa�w�W�mϸ�~JS3x�_�w����A[�Wa��^�����D<����S����F�xմE
��'�F^@H�ԍ\_�X*��k��"W�+9�����Q�]�j������Aj�fvc�x:�^��pV�@������n�W�&��K�-ut �$�U>$х6}вE�Z�60��0j�NBrcuT"�v6�ǛiP,�[M5�u֕[d���d���(|9x8kK�Ț��}����gy������0&A78��}/w��)໑���7�@�p�����:^������||�!���6m�X+Z�,@}�_'��+�X0�=7?*g���'��ݤ ,��f/��UKEj�eUN����R1����ُ%���,V�w3x���{q�C쥊�����'�@˸l�NRK$s9_2�~��0P����v��ߝܿyC��QŜ�ss}�2�_>��]X,��\]_�]��W�DN������<��aԘd�=ڿ�^3ji%Pl��Yx�諪�c$U���3x��Nn��^])E
��?�Lb�~��E�<%#s0zw�����o$��5��&wű�{כ4+RT��wO�P��].)��c����~\���X�Zw��<?/Ҹ�Ҙ<���Z-��yU���R����P�!��<��t���|���(���d-�mI�lhT`�'���u�}sw��r
��%���h	��3������J޼���;��2v��7��wo�r�@��Q�{���<p-�}�k|4q5�;-�;�m����9��g�#2R4��|�R T Yf����Bno.	��a�{�������cQ�1����2�*4��b5��t��nכ�Y�lN���c6��N3��#�y�;KU�r��ʺ��?QA�X�Ϯ��#�:�qǧ4˙L�Mw����<˧�4�A��h�h��`*	�x�k��Z���Yx�A|F�������3p2Ӥ )@�f�i�$���|I���`���rLLX�.�a�^��רCbN�(�¤�X:�&ΨU��kc�V4��,��>��% ڑ��^	�3�,�t|c摄q�C5�z��&�����-k�̰Ϡ=�G�YP�-�<�1�=&�,��b�p�Gu������!�:��Å6�4���N~�$���对۝�7�9`�ρ��39M%�[GI��Sa(;,�U�Fc���L{�ݛ{y�V�Q���� ��RV˙�{��fp���{C_������������5��2��B	��F�/A����H<���������HF��r@�'X����'UJO����xp!h��+X3O~���%Y�s�Ե�8J��_�ARj���FA�x{��wgDP�`}���+�ﻆ,^$Q�j���;@���WW+&���{���>n����3��l�H{�����u��B��6o7Gۿ)�*.�����@	��Aك=��J;��v��?h�w�m�|�1�$�����_㐎lg���jE&�1��9�n�?]?����XrGe�W,�Wg�Ŗ���U��g�M�Q^���]�`\��:K�т�	�8δ���b!oҚ���'J�qO��6�ZM�`�g�2* ��g�j����G�4�UϤ�' C�4u�e�!�\�oPm/,�2^�=Њ�E�܈�]������$.2#5(��SjB֮��n���ОE|s
K���E^v',���<q�G�@����Fg�;�.eLp�0���GG���ŝ�:�u=��ih���5���& k�#��6s���^֛�&�)���=��K4��s�g ������2��W����rw���dׯS,��XU˪Do�+�Y�f yP��N������ �ˁr�rus+�w�����X_v�?�����%�߁�ʯ>~���ctɖ G��Bӽ2�`�p�������<m��&��4�(w���
��/U��Kg�?��*r����b\o����"m�7��6��f�f�A�:�yL7a@FF$mNd,\sæ�k�h�o��Ҡ��������Vj�C1��P[�Eٿ�K |�+�G ٸ���^l���9���,�l}�y��%�X�S���D���E5iYq����G4����t{+o޽����^�Դ4��7��]RO� �� æyw{'?���:@[�`$�l�q�Lv��ƞ6o ;t�U+5��wo�ȏ{����<��~���3��(E4�6msްA5(Y11d�MK��AT�1Os�c���n@]r�
�q8\*-�W{5Fb�S���� s�Mn��û�\����HY?.�m!ա�L���ݽ������L�ʫ�zK���<�`�#���:L�
~��'�]n0֬	5��: b]�9~�F�hu�>�8����u�@��A����i����Yr���^cC(�l3W��}Gp�C[�M���r����-�F +�`�5�힁��G��n����4P�mqȪe��=&~��1��]4����ثF�B5���d-��B=��y�+�b�$f;in/Pg��3À7��Z��u��m�B����APV&£��w�?б�m�(h�A�8��b�{
�O��g�`�o�/^p�=k�6̡�3�(�ء� 6�n��F�;X2�:�RvY�`b߽u�#s�e������hm78k���_�3e6�/z|�h�V���g�0:(K��Р6����x�-�U�{4�:���j�J�_+)ml�Q5��B��ò��q΍%3�����:��J������ s�9d{:3��Q��/E�r긿&��s�i��_���˱__��i,�^��Lc���(|��I�A�T�[�'`��6N�QE~��q{�Z� S��?�f����M�����c�H<a]='_ ��>tZ�i���w?���៘������Y���1kb"C�N��߷��0��6Lڟ~��%�س��yH�9� �`U�9�l�u٤��p�Z�?�p�斌P$��"s���d3e �3�)�syZ􀒭m�bt�A�m�����/����*�1��I��ɗ��  �R��7��9�}�6�4z�9m ���
e�8'd�7�4�jU�*���_@��0iv��.��T踿��W@K�vJc?5- ��Y X2@����`4
T#a�r��&~�8�8�`��n�}e��ɚV`~�XǶ���������x�x�����&r��e�Pl��t���@͌��`��y{{E���.���@�"��i����NEhq�Sؚ��U
j{yHk)X�:�/*!�
�����S<_$ջ�>���D�u?՞e���y̟U��uj�[��'F���5)�I�F��{<Gh��n�Ǔ{����B�<`qtI	O,MY�5A��%8�gF�0�aء=��b�N�(��3��Z_��n��ű�|y��ѦO~��b��#?�w�p��Ψ�Tc2(���|��/�/y$2���]���^q\�� �L?&h���&� ���1*��M��ݼc@�C�	Qi�5 ���ϒM��pl�k���?����0|?Ə�������M�(��٥�����<Ѧ�Cr���R���x���g&m�v���������vy\?����w?� ����� ��M.����[��G9S�(��A��-A��d��`�m:�5[�*B��,n(��!xߏ?�M��/�0���̒u��Jh��P�VY�m���`'D��@��i�i}$��ޅ��
1���Z4�������|����U����g��1�P�t��v�A���nL���2M�9�ptE�&�2i�QA �MO��j�6d|�!𸽾e6�~`)͆:1�jX�Y�[��pgcmm�EKW4y�Y) ����p)|�h��n����E(8�9����1Qw8~�1�./��?9
^S.1�4�v��i|0�q�o2:M�%�$R49�~͂ �-�2��b�GC(Ҡ���|�0���U�7TwG�	VPddh��8�.�Yt���T�urB�rE�eIt}`x3����X�*�B�H:�wi"�S���,�Κ"�*�5��723C��� R������Hy<�QՌ�����4g��Pn�[���13���5?Y/���Jk��a�d*l=�����m0���=f�V�p�Pf��y�����N���,�IA�fO�H��,mr���`�oQ���%{��S�q0��{�h �e�����.�?�)ʿ��ZF�ͻF���Lm��A�{��÷�U �i����=��05)�j[����X)�p��{�NC�6�r�رR��v�ۮ!3�uv|�k�Ę���43�ca�`Om��R���N�;�D��S�:f�M�{�o>~� fW��*Ǫ�싹X|>;�;bd�q�q4VkO�O7j@c��5�#u�\o �P�g��tŊ��-v5(�0@��Z�S���	�g�:|��Q�d�s������ �t���CN�����L������K=�8gs�S�u��J��郬x�Go��L^ ���,�a�I:�*�>�iO��6[��}�kr2��q��}��&s�׮���e�1��˅���)[�q	`��P�T���F�l�'A����wvsm�p��`Ì,YR����G2$Z	8h҆e ui�������%����`�!h-9&c��.��߮o/���H{>�\�l�j�"���lP�[�~N�i�k����&z��-�9�X T5�i���LA/��͍2��,��e��?Z�ߚM�I��\�S�=���*� ��V�ոGH� ��Z5@1_v[��-Bg����o�o��-M���i�io	�G�9�5f到������_;�
�7b�U8����Ӹ�b�Nn��j��cv�5�0�Ta�|���
���?|������1~��7��p9�ٮ�N!y¿����L�^��Q��9�)��=�Ǐ�G���laL�cEd�*+)��K%�\i^z��QɆ.k�1ג�v�R-���V�H׎��i]�A�G�����?ɬ�L�� �.���N$��_�|,�I*���%��`��*-}���?f����t�oo�Ȓ��˦�8������YL��o@]2�2�!��;n�1ݓ�����;��V!*���6� 0�z���adQQiި�L�]y�Zy�]NSL���2tV�v���ؘ�T���A,B/�|1iC�)��vl`�)��!���wo��K�>ʇ�O����lv�Dˎi"R@	ukdZ��J@� _�QOO,����^�޽���I��O��sg�L�/��&�#��8d�W�
�+��>��腍�*]E�:�!�ۏ�l�W@f���m��*�= ��i���*QEk��9, 8�슄LW����+�4��?������=]��n�P�G��c� o��B-#��" �n7i?p;s0��-+�C˅Q0��*�]��DSDv5P� '��c�.�K����M��%�r��b��ɒY.y���A9P�)s-��f��\\�3��l�e�TQ��5�3�l6G��t��!pD�)I�qq 5p~pO ��@�i�L'�:4��D]s+�ٳ�� U����3��5A�@zl��T���� �T$~�R�.gb�;-}
���+-�Q0*X9n
�6��U�,��1 �8^�.X����3�9֦�iٰ��������S��(��Ƨg�u�
��k)�� �_�|��ԟ���=��H�n4jYId��cL�؂��{qn��F�[b[+޴�v{l�{ch ���R�֤��X��L6h%�tl������� lӛh��/64�/y䌗ފ1�jw&J�?�"Yđ���s��旟;�r*͂LO�I빋.b��i
l ˯�s ^�,p�.lK�6ߒ]� ���ϲcG�G��኎�T[ !�38��w��]X�L8��'�}f�!kG꼬	�Ѳ�����v�Q��Z�s.������C��:.�Y�9����c���f����э�mu�l"�����	�4 �c9J>gq�L<P�qjB�ￔ��'?JaO���{d({�d�-��v�Lmm��Upv��3rcZ�a>H���-���Jio��D�7X `�����lă��vsŠaG�<e܆F���y�VK��n��h
��r.����E�a�ϲ@�q[4��:�@?2}?���5J�P�y�f��@_G,�Yl�rE/w`m�L>2��[/V�N�C���E�2�}��kK��� K)�$�C���� �?a�����\���t�O�\v,վ�Ap���bA0  �~U�eP���K��=�y�g.���rأl��F�%rZ뮓ޛ�u��+�X��JOPv��t8w 0Z2�e��u})O	ng�ɼ嘀��P�D�������%\#�2�Ax������Gk�\�rhjhɔ�����D�C���>j"R��ݓ�R��d�@�RGIK͠��q�oJ`n,.uS��)��Q�M���<��|E1�և��91y��P־� x���qb�&����L��]'���ĤN��c�%�C��FL ��w���yAjSL� ���q�Yu�(�ѩ����e���/���V2X�<��7-c�2��DiB��uW SN�6
�g���{Ơ�-������^K� Oq�?��G4::p(�]|�˦��rr03Q�2ZeRL��?�ݧ>�=��I��q�k���Z.X����d�GB
�hÈ]��/�/��ǟInyڮ�k{=�V�Z���Q����\�ï3ҩ�9�&��o�)����%t�5t��8��g]��z���ے�[��,?.�c`�������v�I�$�����7�1�P{n�����;���책�-���M��q�M�L��������G��.���l��
ebK=�K*�(yF��$�5ہ�꾽�ҡ�C{G��ϫ/�N���!����,�M�M?�Ϧ���OA�pllȻ2��fؿ]v=�CK2J�r{�&9�|��O��_U�#�����;�����f742>Vd� x����c�q:06��W�٦���	:E;ꅌ6�p��@pB@���Hl���
!���g&�=XW����K�̐�%}�72�3e��@�����e$]�9����H������W\�a���S����邳�l?�Aս�����F]?��$dĞ�7�[@����e�����(�*�ȎpX��ޥ���eI��������0�*��:=��ɸ�B�����B�3wA�{��j&MtӉ�g��F����B��?Os���&a�?~�D�dU�fF�38��oԩ���gv���/i����m�;�%�F�c�	�?�呝lqP!TC&��EtP;���j���J�=s�jd@=��� ��24PWۏ�a���J3��oY�g�A?�� �^j����*N�g�/a��=�|�{��Zq@2�B�W`ǅ@G�4�]i{�����ڱ3��m�T�&;���ɜ��lE�Y�kL$�A�1��N!;�)ݻv��z��9#g0���&~����Gsx���wY� �_��X_�l(����A$6+`�nf�� W�Qq&�Cf毩���������]ϰWqq�M+{c��d�a`K��c����=�����h�����}UU�U�ч���J��N��pϿ�Q��ו;.�_�Ó�M!'��c>G_K����}��1��%�e�9��^� _�I�([+'��><���VY1H\_�ٞ�����G�o�����C����@re=��]�	��9�أY҅��wʔ��Q�&m�;�O�j�(5������t`���*譽�`I�0B���l��	��ٰ�+���5���5q׬Bn!t�7s�h{����H�+��5��gs�Kd��%�e�+G) � ู�`2K�1z�q�Y����SG
�48@�0�ϊ�"�{��3�=��Aɚ�����J�%f������MΔͥI��l|~L�T�H�X��Qo��M�VP~):7Wd
᚝�������/9������K���bᅼ�^�����ܴ�������iMZ�o���{L3'�pĚ���"������ր��C��Tw@�� �o�5z%h�1�^ӆ"��V��a�
'��^p̝��M���T3�aq�/�>��}�*���G���r8c��%�{c�=�Y�Ie��wܓ��C{�M�g�w�V�#:��f���ߊEH�Z�RGK���ـfh3�Dݩ�ےk�oj�ZYj0��7y>W�S���� Q��-˘�޽�W�k�&�q2�%i�>�+�.���,�s�k w�ޥc��ۻ�pL��<�����yEq�dR�8΍��#¶�3y����\�(-[o���t�5�Z��r,*�F'\w����t��GK�'���ك��S܉����L��>�a���]�j�6�y�miUڤq�&�K�%�xz*K'�)0�O�)(@M�م�]J�eR��d�d Q�5�.C�W�wm�\y�Ę�\Y�S�.8����b�K��3[�o4/S������/��F>qb�9���`Q"�L ������������EY_5U�����EШp�|y����+�3X��~��I��� �d�ulʤ׏��Jl.Hs�1���O�?~ ݖ�sM�x��nI1�?GJ2�����4P���X(V�;��;)��l��n�3��2{���{*�gm>��3[����4??��1���o�4z;��Z���2�a��稭2[�Us�L׌`�v�	*�ERcY�����B�?�+��-j�%��	���t�-:}�� Cj���i�ҡ�01������=����u��Q����P�����#���Z#S�.ʤ��8K��"cʬ\:��WQ?��ь$ꯑ1���� l����u`ٟwܙ�
�W=����}�{@��B���?����5����'=xP~lC���u�i��5^��^3�1�j#KW��9|<"�{���^��;��vNf�a����-�/�}�]&���Kd?�s��i}&�P�I���C��"��q�nx'ߟ��89t܂L��o����۱���,�P�.n1�u]~�@ h�i4�mb��B=ۯ]o�<���6��E�KK��\�6-if�<���<C�-9C�.Q�[�Dƌ���̎��E˴"���(k��K��&�����E��lM`�)޾�ꎫcJʸe�[s���5��h�B��or�s���QJ+�XVg�N�>�m���g��N]�o
��$��V_��l���c�n�|-�QU�Ce�%���V^��� 5%(�7E�؝*�T݈|^.���(��1���
�{ 'ѱ:x�oW׷fp� f�hyrԖ�؃��M�m}~~br��N��(��i\]wd�P+�Yh>��{�h>w5������5,�l	?���2������lxc.[�N`���#Kw���(� 7�\��5 �6�h�@�_+C �!;z����uc��1�a�@?�ּ`6i���y Q$�cs�cX�_�����蘔:��Wt�w�~%�Ǡ�zEzθ޹�D#�qhC�p?TT�Hsa��YeVq�{V2ΟO���\r-2���ȔM��� �)[�ǀ����*�] ��C�����d �}́G%�+R����1������% /�~j��9���� ���� �o/3�5g{g�U�U�:�Z0�>�b��Mp@ǆ�MM��8��c<������{m�(d�+qj3NF+?���߳�0Ū�X�O|}�W��+>g}Z�)'��Yn�a��%^����hܤq�L`�6,����A���7xL�_mc����T���hBv�	\�qT���;5I�>�&�����uk��Ꞻ3d��\���ۿ� 7͝\,���f>X�[K�Nf F}_�N�5n7O�u�$�pŲ�4��5p��Cs�zi��6j����6����=���$3���yl�D�����5b��g�=V����7k�x��=m��ȗwְ�y�f�S��6���羦�ي��F��*��V���d��aS�'!�*�>q���E7��At7�}�_?�"�)pEK2��*K�k�az\?��=�gH�d���w7"� �t���l�n2�G�<�XTc�b��$�*��v���k�n����,������J~�������{B�L翔v~���N��B9 �:ໂ�`Q�y�B8�z����8`��.h/�L���#E	�H��?'�&�I��m8?���r���A��C6�$l�Λ`��	OcSnLշ1 �:7�'2F��4W-��r���j�����i,�6��b�m}��-H�.8o�0f ����'�[2Hp�-�W�*C��a�N������� �Y%m!g8f���� �-�Bblg�`C�9a��
!����%���@�ƅ�N:ϙ���G��a}�����yo��1k� ����t�h��^�6Ӛq8Q�gb(�0&�`m�Yc�u�uћ��:�}@�Y>:c���8j`��1pnnny��1 ��p/"��A�?�D��}����+P����^Y(�N�>%�w궕�uZֆ7�F~y���;����03���&[3d`e}����3���D��>�go⼼*w؂j2�f)7�;�7�5��,��fZ�����6F��fN����I�ծ��V�Rt�l�Y���o��=�T����s�.@�|���z/���� ���K%�#�Z{�2�Nڅ��1X󌘱��M*2;��$\\��ԠeTީ嬳N�b��_dl�jm;�1D�И�aDe׹���>Ap��ݣ�~F�jE�ۭ����p������v�t`�i�D�a�x�vd�e�/�����x��0vJ�ـ��{L0�(�l@1�ٝJoa�{v�&W����z��NH67��S_���5���
��0��_Ù7U��#O��f5i�꾁N�>��D;�;���g���L@�X����d�k�'c}���J��!�� �m/�mk��uI6������1'�����z���r/��W d��2#�	��|���t�a��g�����o`�I�?X�H#veC6z8��:e�1��~�^��=���`9���nr�����HL�{̺k�>�D��>�p8� t���' -�;���@ͼV��<�`WG��7ô�)D���9��!Z6L]79FȌ�=fuqM}"t{d��L�l�֍&����Sv l�2mm�a�.���5�T��#�^}�����߯Og(���IU��8��вz>�sc�j���Ҿ���3���Օ���-j���R�~p�9�D|��G�QQ{k{ ��®Q�ey��%�$�}�,�`�*Y4��xW���\�BRJe��� ����	��`)�V�F��X㱆�=9��~A���!kp�K�79H}�<��8����r��?F�o��8P@9�FPA=Rnη|��wy�#���4��hԿ�lB��4{��	ZT�JeU�%�3r<~U��h>'K�*�%��ƽ���3!6��l-K�F;��Y�]�q7żtp\�}Y�s��C��ig�:�������������7r��1����IN�yb>g��8����9�%���R/[AH
p��?/�Ko�=h���k��	ԈT�����h+nG<Y����Ӹ~��/?H�oT0�Zc�W�y�Z�A�FFRQ��q��x�i�MU���r}����2�>�j����HR&vZ��7_�#Kg���ry)('����9m>�i��:����t�R�ɓ`Dx�.���J��V�,yx~�vې����V��]��tdcV���m�YhTy7o��Ď?=Rj�o޽M��]
ږ����,��`$,Ҥ�NǼLF�2:�4��P({V6";1��L��p�w<<��޶-����z��#<Q�ȒsI�?�9)q����
�as�$��b�09���� �|���Qk�V� �	�9h��KnҨ�G�;*X(�% ����� ��N��쯟?�@	L׈�(�C�J�w|o<f�:��pWL��H7�n[a��^ˌӞ�;6u #l'�(���Ԯ����-7K��o2��L缝�Ӣ7����܁O��`��Y�����Y6�dd � ��F���ۘ�u��y��x�w8O@�Y�4t��9�d15;'vQFSC���2
���yBS��6��vK�i���B0�l
�`�J���x�k ���m:���˞2P���gl�X��ZH���\ ��h�����M`��h��n�i?=n��s8XyR:�Y��z�;�aԳI�m���e0��� �(�d	�`�x�z"S��j\&�N�}^�A���W+��1���)^�d���������rH�<�(��r�:}��*(;��[R�jY�k{^+WN��-N/�:�g`G�6b�%�b�49��b�"��f�y6���o�epF�5��r��S�ju������23fk��ʕW��l��V�=> ����ۦ�!<�	#Og,�1jG:�]�����-��q�$'�8�vX��F��{)� c��S�$������|��{�S6��8��5 J@�\�8�l��$� u;Yu��՘�jɰ�P�p_[�|Bu��5�4+K��&.���tO��/�QO{9�%��ߗ�?�a�~��L�Y�3�Z���޻~|� �{`g��I�N��Ē~,	
���8�O��F��s����겑��Ρ�FS`G˻��e:�C�\L�חϟӹ>[Qֱ��<����@P��wQ�\��,[.��������ލ�K�ԼhP�C2Q�y:�u���9w�����k���G�,!��Xv<����vM.���	�\u�ViPD�:h�3�(�erà���^�sf�yk�e%R����鴬.���:�y���sI�b۽x�#h�x�vd����/����f�=8�,N>]E9�a���;[#������W��E<�ae͢�ے'��:`��}��}�s 7Z���"�I��q�V�@��n `�Z�$i����O&ՎK��Aa�f���g��?5/�O����*ڜ*�=ēM����"���ꗧQ�n~o�[=p��NɃL�D��!��5�u�����}�ʨ2��t����χ����9��~�3Ì�;e�^,e#�G١1�o�����>��9�&6Or�tK�]�Wޞ]d^��K�����1G��r)���b�V�����
���A8����`�ުo��K��
�����/�g�l��u�;2�Y�I�Y7�����K�H�h�X��$s�����ڑ��tg��\���.��1�bqxQl�ړ����$��h���fqamOc�,4�S�-m�bp��^�`e2zG��|�0�7]4�#���h7S�a��5��k9�UP���@DϩQZ?�~|�V�w�o�����Kޔ���t]�EyN6�� �������T�A߂��H�uJ�Y�ꢛ������}�<F��Di��dN �Pg�6Y�谼fN�A�`������f�R�p���� ���nh@� �Nc���ܨ��h�� ��K`�rlؾ�]	�4��[�4���b��Ghb��8Fxh�r�hf2tl��j��� .��*Wz8�<tԅ�
�
�,Qz�Z�'
l
2�,��΅w�N.A���I���UѝJ�c�a���-�۞�-�/�a���8g�?��J�� ��g�x��1�׍g�ʬY�zϹ�A��i��y��ީ�}ޛq���[���#p^�Za�P`��%�kI�d'>~���E��Hd��@��4ĵR�	�1;�����[�P۶�~p&!�l&/=v�.g�l�DT-��SD~Ԛ}�E�i��o a�i3��#՜���%m��>c�q�o>W��a0�t=�tn�.� $����VA恵�-m���� �_�p&�Ө`��	E�d�5m�]>��ߟ�&�Mʳu�c��]�]j�I�ZoѮY��e�k'�|_��S�
j+8$&:��n�;4��X��p,@�N��� ��.��N���f��6V~03qҘ[�����A��{�S�Q3He�\i4�Fw4�/q\�cg5u���qvO�o��S~���v"pE�t������X*�6Y;���N�X;������ �ߒoK��uo�;B	:�@U��L�����H�O����p��{c%d`�x#�>����}�)X��DS���V3٬��'�[
_��&ص{�+^��90���x�2 <�vs�����p~�MW��׆{����??|�uk���\]\��(X�z��s��G��ր<�� ԹX�e�V�N�@F�`���:$a,H�F���{�u`{����1�U�]�� ;Gem�M��_�Z�P���N�殮_	�6|,0?��aPE�vnh�����n�9����>��h�F1�͖�!:j�(k��}���K� `!�ֲ9�2]��RgIyh{��"D�����>��bI�_�b��#���c�S��^wNj�h@�v���X����Njm��Ie�L�)�H��!�9�o���t��0�mm�'h)�C{��\e�1�1x`[
�����DG��OM)�.ِ�߉׌��Ѽ��6�r�
����v�ó��SdB�+�R;��!?U:�Ε�hEА�!Q"�Z�1H�0���*b씭2�$2V�	�X�� �k�oQ_��P��\
� | ��~�_~��|~�,��Ky��9�=9�����v NĀ�R��W�l-�R�A>}��v����"nEE�v�V�N�=c��S\�:��֨��24�� �SMĉ�Ŭ�q?�g]�`dD���ϙQ�\=�1p����c;��w����9`�.�'�	A��NoY������h=wA����Y	3���������Ai��e�s
Gp���f�~�'�I��)� 5��h���+Х�!a2,Q�����[��I{2�o������A7��AY#�[L��x��(��͸�n��R=j;��@��[=:���U��y�c�N�L!FHA�Յ;3r
��N��KZy6V ����Vu��Vo��&N�-)�L��l蠴60\@ ���&� sd!�Ŋ�<1���ٸԨ��Cx1*J2�f���E[	�z7WP��]T�]h��3[E7H�3APg�N�D��%�d����X7֤�U�J�ƭ�V�L:�8��r-��A�.�M
�"�ڂ�e�Th)����~7k�I����ރ�sВF�S��f4�
w��s���t����Y,͓��>B&�j�]:�#�A(��.N 9�����#y�m���x7��ksQ�m���K���C �*6D郊�&'�"��:d�h2�� �����kF���<�mtA���8�.89��gv ����{yl�DF�5fT����5D��o�lL��Hz������8�1�� j�`a�߈1m���oBq��$��`k��R��f�YV�,�������ӕ�C4��b�d�."��v��?b�{xL��[�Y�ٽ*@�|ںQ�!eF��j,�}y.����L��[�eW��i�|��Uv�
v��b��q4[�N�:�:H^V�}̡�(Z�".j�G�A ��QYJG��֍���?�D�{�����ۍP�:�2�_�8�Z�����i���~���*|�G�
 �#�Ҩ��r:R|,�i�^�3��sb� ��Q�3O_�ç@7,v(m��OA�S�-����M/��{�H�[�9�"��`��v��S�c�7��^ l��DЈsVm�F$)#�-F;����+Y�<L�c/ڦ}y�~fr
�ą�W[�%C �eB��gy\�2�5Q[����M�����+���u�����4��W�@}��t.��v�aq�����t*���;������Z��Lz� Fإ�Ɩ�D�Q���>�Y�S-$�F�4�jr��)��c�I)�#<����p�=Y�;���<���Z\-aML]_ߚ����L<X�9�1��[qZ&칵��dNh�5T������ɂ~4�h�D#v�bٙ
X����>Z����q$���%�Vn7' Եi��{�i���k�o�<0Y�����փ]���vڨo������Ŀ��i�g�$n�%�=�������7�oC�Xse0}S���6����V���`;�˛�ƛd�����Bi#��Ŧ�����]�"	z,+�#�ke�l������k��4��JL,B@�˧��<u��UA�"r���ʿ��d���3�U�����A5�z#@���'Xbe^��Sm��ҕ�h�+lFKh�>C2q�|^{Sl�_P�{\C���]�Һ��$LB.��������rnu9�&��5����� UH� hм{�S
8n������h�2 ���o:=H>l�&��3�?��T;d�Y辵ۘ�t���G��5�/'���n�CFĨ};(�c8�:
P���_�|f����Gy��y��G���c�o��(�#[�/� |��k�KAv��$����_yy�m�ڥ	j�>�sfD�Am:�*i��3��=�^�^WoPy����h����C1=�.Mu	)^a4�hY�-�!��a~��2�@�@��69qa#δ��)T�ҡ���ܹ�MDǑYh�h��7�]H����	���P�LXD���M�Ss�D焛k
��[X�M�8�Ն%�@�%&t���V;wE��l��R�~P�\�zCb�r2��^?~��r��Y9�u�|�]##��6�p�R�X�X��c�r��l�����ӎ�"o�J���=�W!��YF:Y�94�!ɺ�����h�*@fh��Ϗ� B����#���D|�Z���^S�l����z���:���N넹Q�N�;��r��O�c��m������� g��fCt��VK$�-nw�Xk�áKuPFg�Hi��A�gk%��e
pb����H�O���t:�h14���U ��Ō�:6TA�~&�)�*;�'_��:x�I��hYi-�����]gx�
�Rc|SPǀ�&_�tD�g�Q��9���aP5��'����v�0ji3r� ��u�<���iiD)���7�R���뎆~���O��!�C��9��Ы �����4�X�НЦb��;{�@;�Ʊ/�fvfPay���.w�3��b��j7}cK��U-���G�����G(��u�L���~��;���d-��=Ш3���
�[2��Fո�@"�&�(��9��
��0�ڱ3���t@_o+_T�W�I9�ޥ��MDlK�t�W)`4��X	�`/V�c)�j��lv���o@����ܾ2�ԉ���QL�eG�V[�Gm�A}Zj׎����Z�G�;@�n�S �D�!re���o�k�3�@�Q�s#��V�'�T�O5�v�����i���E����T�^Ǳ9��Y���9@^hzc��oY.��;XC`�tcp6�v!���5'3���G]�ވ��~���(���I4x#�k�k3���:,}���=K����T`�v��;�_�X_\���#y�v��ԉ߯ό
P��T����/�<�4!Wvh���d�7�{���5!%���y���󎺈��^Ũ����*SjN�X�|�y��9	 |�#�4D�D�꺉1�ra�g���G��:C�X _�G�<��o���/[��TSn��V̕����Պ�pڶ>��Y�����B����y�hI�7@���u�jL����M&���4�C���X����«�i��|鳇C����ҭ@}	v��qk]ogZ�W@�(�QD��$��Z�,3&oԵKێ5yY��LNT��j���X��ƛov�x�Va���˨�$rr�?|�z��������ϛ> �
o��B�������3{��9��I��+�Gf�/�"����Or}�n6)����sq%ϫY_\J��<o�a�h����y���7q^���Auܫ��b�� C�QQ���m��d���^��_@���e;1Y`��Gy����K���?�!�t�׫k:��,�ѳ���좜�JjǠ,��}��/����m��`�'�V)ʨǾ(w}M`�5�P|HQy}f�&���:��� u�Z��b-E��$�)CA�VU�Q�s�o��	l�x��3ۄ��˥��Zp¿�9��1�[�����q�3y���-:4�Vl��2"���V������ǜ�n�3m��W�p�yӄ���7��#���!�Eֽ<���y�ɩm�P��x#�y�8�-y�J{�V��а( ��C6��ҁ���+��*`�N��D����V�8��zǱh�v[50r��)؜~F=��>Ճ������s�w�ZQ���Q�I�9Dl}G����+��d5��[��Õ�90�N���D��;	H��OA����M0sG�,�h�끔ہ�%\'uS���~`�R���i=�\�wO]7�\+M|�/�l�)[�t���0�T\�(�߀��n�Q�I,;T+)aX~A�I��9�4�gca���z0P'��s<�0�1Z��P���$��<��W����	��$��f�����_/���1k�T�P��q�&��5�ǁ1$�#Bx�b}[Ǿ������pa�&�|Y�ka�cG8��L'CE^�{�VnnoYƪvo���v��T`���]+S�9��n��P��!�?P�MY�ޞ^�muO����c��5���k�c�O����w�.k�ꑳ�#>��&By�8:;N�DO�����ybO�o'�Q�x*�E����� �Q�4&�ee0�o��l��v{kB���]������?�v\d[����Dm3Y��N�K��Gu�y���9cf�3���B�_���A�Z-CUb��ӵ��^�l`�In���3>]85g|���nf���?w�jM�X�kU/��qm!=T�Z��M�g�����a4 �7&�`�~��G�>Q������.��
��X
��8&l<�k�MW�<y6�3�\�6/U[�{�,.f��s�r6���d��A��+�)��2���S��k�����f�%���'���������W�P�o[�2=B֓��=�u�U�<Sˎl��K-��״ԫ�1z�L��H�1ʩv���<��l�=�س�N����A3���ngK���:�l8`��}�A���z��җ��93��9=��Ϯ��3EV{y<./mi���L`��\�P�A��P;.�y�g�e�1hŘ��<&ː`���mJ3����E��
E��~��=g��l�є�Q��㈾�:E�C[�$�U�h�K��A������]3v�o0�Zg,y2�jJ��woɀZ�n�2�<��-�P���mS�ߝ=��ߙ�@qvi�*�Ǟ�Db̙�®�X5���ǵh��3x%!��+_�8BƎұ
V&Y��i���+��{'?������M-�9jvG�r�&�M��v�@���qC�	�k��vɰ�Ќ :���e�������]8� �J��]E��Q���3�z�΁%lFgb9��Q�~L�����:
�_����]����]�lP���f�'��#p3��bV���`���u������/�������ېi�F������|0��9�
 �T���x�( �pkp�&�
��cN�e+e�ssq5|�=:tA�
��e6�il3Vc�`�Ό"�W/�(A�$Qh^�/�����j�[k`mP/�cAtG{^kV��*����lyI
3-�k�[�c^-l1 �leE�ꅐK���7`倽Ѡ���sCk�m���	UD\�
�Gү)�|�GP�Z-���4= up]��"�Tfhf �x{}Mp������A�88ZL�d�����c�ekG��9���5�E7��ׂ�;��2��t�:o�y�jv-��]/�2Y�8׬��D�4;�1����`
 �D]]��{`kz�A�c����CG0P�7-Yi��Uj���J�Z���8[@�Ώ�-�,��
 ���F��A�\��A��r�/MH�OEM��FW�D���r8��QW�l�~Ut��@b?���}@F۸[��%;h��騸�	[w]E�=H�Lϥ�X���t��-����v[37��xe�N^�5���f�jf��ܱ�3��������Mo�Lg����;��ۘ��e�\����}�'8uL]շ4L�W��,��'��^��(��&����L6L]�%o��ȿ�ۿ��woU�,k�����B���;�3:�$���'�v�D�udAഁ�-5/ֲM��.ٔǇyHOtj�]�l�!8�S?�<x�{��%���WX��IZy��d<�9L/���_\Iub��`>=hun���ua�a�v����Q-�����'{���[�����̀::8�dx�G�Ƅ$Ȁ$�q�1�V;�Vڙ�`~h��\��������sU���*�?�&�EI�k/��v�9Xq���p���"ځ6�Β�\�G7r�|0'��3A��I��lu�R�u��9hS	�������-��.��L����+g��ϛغ�Q4Z�94hywV@L�5d
/�HV�2�Rws��&b�-����6��`,׀�8��*陮O泪˂K��Y����e"��b�<l@(j�5d��e��Wd�#4�'=׽����1���f�N�V|E�[�5Z~ϟ;Y�Y��ߣe��<����Y�@�|��E>�7��:��(�[�&&)[2� q���C��^V�=Y����{M]+v�j�7-����`���%��܋௉���W��;�.ʙ�Oԉ��T��y�q�s�A�_�?g�x�������hv�L2��6?���:/�˟�����7��HC2Ĳ�	��X�.�X:�V\,	��o����Ǝ���w�^AW
"�Д=Zb��9ZS�<h�1��s:B�QZ��s�ZTY�J����`��+^�:��wo(!v<u�b��$9KxF��ְ �/�����4�C�dBR���1�?Ʊ"X�΢��lKÒĴ��.?g?oz���_�~�&���Fg�4�?�^��+h��L�&����z�l�*��޽K�5���<&Gb��d�oVW�&m4����NS�5���a��(����Ӊ.X/�F�<P��\_�ؤY7�-����S�|'� �:,�Dp��jG�k��]�T����gy8~T��ĢB��������c����|�}dǡ�62J]�(��$���~�f�~Kd��׽E^�nt4���F���J#
��Օf�PK�� �(�m��:�-���H� Z��ś/p���@����2��5�UtN�Gz�F�UZ.�K�"m0
4YP��X�穯��)�wn29�� �s�N����lF �Ѣ��5�ޞ3����r�d��#ރlǪ����i���P�M�\{&��a�l&�³��,=�\�ma��4��{����wX-H��.\-�'��?�	 `L��V��V�Ǩ�0B � ���M�EV8H`-����;��դ�jÀ���Q)=��4�!ן�}r���!́���~l]��Y�d?8]�)d��h��nzH����4��b������_���e
  �A�Ȭ ���ñ����/��6N����1�s��+��z���\�T�� �-������u�okyzڰ�Mg�6K.|�����>��=�c|��N_;q�Ħ�g\�^v���L���㔃�|)�d�-Q(s˅Cv�Nb�3WV�����Vr�⠍;p��-,�xr�)�P������2J��l�6�dG�R��ލV®�!�P�6�8Kf�@&��[=����%��к�&mI�"���D���ltZ� ���Vnon9O���#��lz��@G� 7:L�u��ڹ���h�\�����jq�p^W�� ��3�qG��(����15�,�(�<��G��Z^{�N��֊:-�z�x�H��}�>7=����9��Wc���S���N���|xh=�:s)�#Nl��Q�ɿ�g`n�9��{�A!��,k��yLi7/{�%4"�H�l��G4M���u.��CNJ(�;P�N�3�=ʸL�[�V�W� #Pb`�$Ȝ��zv�t����MP}I�z��taЮ]����Y�Kd���v}}�q�5��	ߙ�s�hl��>��ͥ�:�̷#;���0��p��ș�.,����q��M�Y�� ���df���c�g����be?�Ȭ��t��tw��d^q�	��T�=��#3Ydu��S���f�ޡOU�0��F�����]UR��6O��*PD�;!pv��a��$�϶a�P�<FA�
FB����ګq*�.Dݫ刭����}B`bN?���9�(b:j�w��&!�����kWX߫�v�D�V�lܙ�mC�p<գ��Kr!���9�0��䒯�H{\�S�����gg�&_�wA9xvX4m��-��y�������q���'�up=�ǘN9w�]�<���*{5M�l�ygD;	>��}�"o~�j)�֊Tha����[&�}m<�{�ydO�h�b8�sǱ���cx�}O��q��G [�>gA�[1��Z��)��d�<YQt=����Z��/&���+4�Bb�@���Z���A����~~Ⴒx�E1��߽n���t�cy�������P1����T�A����`�&���<$Dt�pN�Z彣B�l���)-�{����)�v2$sd�*�|4TP2�K����p� �:�{��w.�4�S)�<
�m�1�g>i�&�q����}�JbY�!b��>~4�Z��]&���el�������k"o���S�ts�CB��9������Û��<$�<�>�ކ?���/���w����ޖ�g�t�H�jr�8Ef���Y���?�@���k��E�D���-dG{L��/\+Pμ�&K�|G��,;��}�}����:�����?�C�����u���n���v���yz��i��cVZ&`�R��	�������n�C��R9�!�y����F��~Gg�2]�����.��.���1���g�x�l$5���6r|[n�@`-��M��+'��:I�+���$OQ��W�\�䈷e���	d���s�
�jOT��Wep�<��>�y�X�Bk�����:�~�: �$�㆞���O�&��O>���Vp88�^ `�`�#u����y��u2�׎��H�C
�Bh܇F�0�]鸒a��#Ď�Sr&%kڶ5oT
gܰ�Y�_���p�7�/�����-�l�;^G;��y~^^p���ӈcp.����`(����(bu��'t&��w�e��trz�s&q�DU7�aҐS�}��^lRy����6�����U�p��F������I�#���N���j���	G�<b��Kɻ7o_��߼"Q�|�yG�K��z�'J���;�c���Mx�ӧ���h�2�#n�Q%��,�_�!Ϲ?��C����W��NYeQ�Ί41����{�"|̶w>����'���M��H�çK���1q���#�it.��9 ҳ��q���١K�*aC��'�i�����;�B�j�pb���l)G�3��<CF��7I��C���b�|-�(N��Z����7�)�v�j��0�%��C����JR�v��������­�	&�*U�jk1p�"�r��Fh��-&��J]��6�$2IM��fɀ1Z�������ӓ��ͫWy��.���u٣| �w�Ni�O?2I��N��H��X�kCR��A�m�Ye_><p�ù��sqQ��|-��D��a�bpg�`��}��M���Jm3 �o�4������]>�O���χ��@o]��o��T#��꣎��C�:��� �Ajh�=�r��G��IͿ��`���+5���~ߊ��Ak� ��]�?7��/�Oid��~LS���b���9�����b��4|���U���(c�SU)أ��fqp���|6ϯUw���|����o�Yq$���o�C�1PvX	f��"
D�觪��e~���LZ���ݠ��j��BZ�>����U�%��k�G`�xUJX ��6��$$i��s�B)�
�ٗ�����p��Y8�!�s^e�������_�_ M�Xl�M��f�[��m���D�7en�ro�($���IY��> }^J����%&s�޳ea~
K�y�B�"�8�<��Zj�7��^��i񴙉�������@�ïǼ�=�I��&ۣ{w��{�_B�_�w���\�!r,0
���5�c��
�-���Gfس|ޗ����F@�F��}�l5�Ae��J"!�w{5�`z����o�6�2�������w�������m.H���Z�nf� �
�yLR�������췤�[6Ӧ�����f�'��H�߭�,Rk$�8���V7F��}��^"e?�r�Sj�%3-%Fo�qx�q�Б7�=���=vtE#�N	�-�q+�Wj��1E�f�X4y��w����oy�p�P��<�@�'�cF{�&��΄'��lZQ���U��"�K��;���$��Ĺ�B5�z�>��D���c����PF�&���}
T�	��j��Qeo����*��]�eB�ϳ���F�A�"�����Z,#�����(e]v�X�i�*�J��FT\�}}�����D�}~97"_��o�XŸz�6������:/�؂hn��2-1H�$K6�����t�(v�����-�ҳ�ts�);N�E�|{�|��z6�P��Z��7�ߕ$w�}���<_�/;���po�J�Fd�����8�C 7��q��;3����h��̬���e��w�s!�D�*%��!��F;�%vNO+f���A��,X-�M�~�Ѡ�}���9{����;��{�}��_u�ȳ��ҴȜ��b%�rި���syuN�,pxL45�����X�o�$л������o]�f,K��3UW!F��MB$�mp�28tS�����g��Q<6t4�n����}��������������p~v�y�*��St+�.Oj֦�7�pr@!����#�`E�l������,�'�����c^����,�n�A(�N*�U��NJu.�\ͣ623<�VI��� ��L����ovޡ*Z�e�ߪ�X�
1Gp/q}��z�SmxV�xް�]�N���B�$��=���t�Qw2fNi'K����`K@q���I����a�iC2������<�^^�U�f�a�Ǵ*���mv�VBGe��W8��4�Bt�BNlN�|/ooD�(Bs���=�j*A���e��<<މ@3i���*����T���ٳ��7�#���1�Lq�=Oʒ>�_t�}�d�~���؎�)ޟ9U{��A��M�Hk\i�B����Ŷ������S=v��$�FG�=1�rJb+���h.a&��}x�����F.�h��G0�J�%#����B�( !�:�s��-Z<�߿��m���wy��C*��jW@���ȨV�j}A�I��hm#`b;J�;�Nqyλ���aI�
%�����*Z%*:-6�v�۠뢐�Ӯ X��v�o|��7?����3?�I���
��ܪ48a�G��xB�aWb5^bG�09G-�5�c�oUP�"�Mі_�
s�G�\3|��91A�8�
C�sXs����GV{1˿"�x�By�B_U�d�γ�Wu���.��J�҇���`1%�������Eo՜(�B�m�o�.2�iʠxN�\�p�眨�xӬifӅP�.̶Sr_��i[���v9&1�͗�� �,#(�4�9�ءp�ٹ�P%��a���O�$��7��Z��%��Ö��!�Y|�o��F�:�㨽������d����:�V,ٙTޟw�<F[�
 �B�;@=!1�$�lZ���"��خ!BV���p��ulWn
���MIO�'O�H��:&�����?�%)��`�*�n�뱶��N
G](�%����s����>������t�'k��T">��/v��2����,���.P;h'���}f6UXõ M��T"�����Ђ���#�[�8�+A��v7S[��:U����I�C� vh��6��}�� _2<�'�A:b���|Ԯ~��������sb�_��>+���芨>�Q�hǊ�pg�pC8�k"��r^�x^]�`��]0�î�gg*V������c�(�$cs�5��?�*�Q��ʒy;H*�w|��ˋe���
//����m�x�)<���ֻ���{<�>��Oq�g~�~�{��(���~�q�������>-ʜ�q�߬�w̀8��o�+���kC�HO�˾�� ���TRJ�-��ƪ��O�����r�iӾ2����CP�憐�l͉�`�R���_^��{��p{w��wy<�֓<�Բ���_d�/�_R�j���Ȧ���'���/�k6F�,l�OdA�<p���߼zKR�ӳ��	�����wW�n�Z����Us�����&�O�k<�_�6�h��J:�(ڍ���u&kI�[��F$t`����QI��Jf��Nu��*�4��	b#k�b�6dHq�`����٪InՖ��$6�h�d�Mo�Mʾ8��J�ә���!��x����p��2\]_1y���y��s�`���Z���i�(����#�@cҐ�n�Jac��Hx�����>}� �)Ae��s�N��7!bPr�B�2���:��aШPQf}��H�ׅ��T��LE�+K�B�}�J��\sP����d���ڌ8ꪜ��|Sk�r'
�#�o�C�Ӊ	 I��7"=D;���)�ċ�|���<�n[C\m�S�կ�Y��%���h2�u��5K�{�uN��QM���0� �$ȞI�mG����Ԣ]\[��E��L*cr=��9�cHz�t.��T�dv��tý),�a@�����m�/_^�a��{���)�9Hf^I�1pղY��gd�a���=��5���ߣ�:l�P=�ҳ�D�����x�ώ�x�� ��(�k�g�%��y��]ϟ��UI�O�6�8��u�T:U�GD�C�d8Q�ƞ����Y��	�9:��������7,��F�Vs��Cŗ�ƻ�\��;XgXsh)A2�v7�$��Ґ���/�g�-�f�V�L����NU�� d���}���N$P
W������E�-�N��=������ӧ��O�cx�c͖ �����d�w%yRg��Һte��c�y$�c	��_IZ��6�7�̍�3�ǐW|�(�s��8 ��]|���QU�A>e���ݮ�@˖��S�e��P�a������|'N�����;#!7"LC�N�,�4I�Z�1��~0��0�}��zK�:�f-�v��%%�[_(
\��c�T~�w��8Z�5Z�E����o6�"����T�*k��1i����Co%'�W�vL����Ğ$�%jĹ���>�v�6��`m��'5=ܢ���
�<1�	#$��]き8;E%��y�ש�9���)��LP��ⁱkq��Y�߂�dW�6_�����lEc���do�5��b�w�g����gJ.�x����k�%�k��YOT�;YH�����2���#N9F�U�\#�t�1�6�I�1j*�5q1��d��"
v�$#��"��VL�Lj��}g��фn�x��mi������_��0��=�%�������_xUI�v��O���$�%!�^�q��B�,���s��ET���Q�`>��2/�(��E\��KG	+��X� =�� �Đ<*{�{����o��u"5e�s�|��f|6�&����?��������n�����寈_���y�N;��wڲs٘jl�[F�qRe��k��9vK�l�a����*��s|οz��s�����ܡIE�lx�M��E4���2T��W5�a+&	�w�\��y��Z�3&^C��+"h��z�8�at��
�3X��}<#�w�+��j�U����l���ѽ��	B�������Ϗ��<Q7������fԒs'�6��+L��ϓ�!k���a��i��>���\m<Q�$��Vɝ6���̈́�H3Sђ4z�ĥ�$8 VUd������]cR��Z��;ɴO�T7Ur�	�8��mb��l�7ѪgƇb�����^�`�����[�����W���*���Kp�܆�O7T&ZQ������DV6L3�pgr�
�k�A�:\ )�el�f��1��X�5��`c�6v,������gsI�N�f�������;S13�m��\mU���E�;�g�<�M��+��f�yV;g2kNH.�XMJ^�b����|�ު`ɲ��Őd#�$����+B��4EF�I������Ϭ+��<34�C˱��|�$�D���N�ּ�ΒT�M�r	'��i��|����<����2�Z���'�N;�F�-I������T�FL���< �����-�=͛��8�W˕��ҭ���Ag���� ��Q�s����g�7��������g6�Ã�~x*�����ʖ��D��\� ��<��ѹu��Y�=���,�����9q�����c)�˾��ʈ
����Jmn�
��o��l�<۸�˫l/�������W$H��y<�;��uE)���[����l�
5߮su��8�{��@�Y�֐���,.UVD0LrR����� �f.��8�O~"!t�m��m��{�����m��w����դݻ_�����z�`w_s��O�}8����;>������	z���ƙ�_���']�=ǯ=������"e�Q4ج�:��N�CCP�����!�-��&U� ��ϴ)J$����4{�B���ÔJ��T&	�(�,xj�#::I��n$�����G�";�^�:�99JD�hH���S=���m��7�dۮ��Gk��^-����a�4����YI�'���L����3���������ֵ��k��?"�����ko�׹T(�h��)�q��8y�En�e�����Pz��hn�s�ѭr&j?1a���	^�OWIKF�Z[a��Iz��DJf�����)���g��%=ܞ�=�o18G�8�Ri���������J�D�;Q�%�ΤRq��g�v₂+��ϵުȋVs�ƦH�>��1���[N@/��P�݆y�'#��!��ܙ'[~��2@�%%+��:�o��m�W��7�+������c��2��4c�}=KR��$9�h�\R](����Kq�'d]��Z�z�-j�2\fu
z�v�v���u���x=i�Y��(j��!6�$rDU(L�Y��Sq��~�r��^^����	17N�k�id[���h{�r��p�&�m�\�㑵5?�v~Y�%}�k��������-~�O���7y���_x4�>|6��`�^��hI�d`ۖ�U��d��ߩ���C���x*ڍ�Q�|�ͫpq�d��笚�\�����r�CrG�~*Y�.�=רv�8lxon�qx��f@${zA5�&o�,�$�t�K1�'K�D��������z��C"c>;��ix�?�Ǽaߤ��h�������Ϡ�X�.*���M�"zĒ8]gr��B�����@8F�oh���ܬy�9!�ڤ��۞������Iض��Fn�?t�j%>x��a�)bn�7�P9RCr�g98���
��	��?�{����QQs����{�m�����X�m��SPA�Qj�wo�?$���儃4�o��ݮyNtVՑ��z�(�
�1wL���cvv����!E�����!V�U���#Zf.^+�ɉ��{:s[�Z���X�s=7�9�A�t�nZ�K���۵�T�����B,�'g�pq��ǋtTE<,�:ht\�R�*9|�m}��{5QJ1>�|%	M��T��3�������=`� �	9�:w7�!�D�9hX�Jގ��9�AV���疪�A5Z&�u���S�'�;ݗ>�w���|/��3UZ�B*u�������!��&:�xζ���X���[��<���oK�`����}f�<���1��t�eO�'7�����>v<�3B>��&T��FҠd5�C��|*"�������v���*\]^�o���ϫ�K�e0����O7y���~JqH�|xN��9��NT�l�C��n��r�7������c������9,�P�W��	>�q������G�F?��t!�Q���t�_�����O?�no?�5����qp{�ʍO���h<	i�Bw0�,aXn���Ë��=�s�
���z,�ɯ��!��~�u���}���[�cO��~�V��e�G����۞�ٹP��ڂ{ʙo雀�H�i]xep	�!7_�܂�N���K���>���|���{�qﬨɢ��fj�&�ή���VtƅF:9���}tbd��6�jy�|e��6r(�u�c��C�IZ��1�
����W۹��з��X	�f:��w(�镉_4j%���Y/���H��7)���}q���ڱ�{%d/�%U��n�dں:i�[�������#%-��0]���Zļ}���;Γ�u6TX,m�
���^�2KH[<B$e^����`b �m��4��?�ڰ���p6����/z�!�'@bGbCS�W(`!Q@�5�&U�����x�U0eAi��8p�ܺ?�9[#��D��b*H
q��-M��j����sM�V�F�÷\@�E�(��$:���T
�6{&�73=��aV��'7���)|�;=�$�#�ܜ���	��|�3Ѓh�0N`�ՖŃ��6���K�-uXw��`�L@��f��~�B��/�^͌;���o�T��y�~�\^�C��u�ww��k��)�V_]���?���������w���m�{�#�J]r�x��t1��*A�<H����zi��9�b�7��+ڨ�C�;G�V�L���ʳ��̔�ɉ�n 5�t�09 S� Ne�P=��9n�4�&k�ٴ��8	�o%9:�?FI��Y?&�x��� �ZkP��KU��nE���[ Fv�7�Wo�`5$������E^����$���vRE�g��*�,S<;�H���~L��8����9�OS��N��Y-��$��/P���oc��X���؆9�:�Yg��h(�	��L%*DH&��� 7��8_�|P�ό��3:? �����?[
���YP�+; un�1��0*H�Y�H$g�) ݀~tr�@&��k^%��	6H��șpdn�-3��P0�ր��\l,I!n����aJ��71>sf����y�+��r�e�I�}%���PP��A]'9�C�noH���*�}g����`M������(��n�c�9�Pb���T��/�4� �s��N�6��y=/�ж��H�� v������̔F{F�*��O�/��m3����#��Y��U3��!�4�T�Z�΍�:#��pAA�q��\��k*�r�d��� ��Nz��A*CF����q�T�)
0�Q{9(q�qo�QK���{���H
�)�	��*�
>�Dq�Az�`��*ab�oL���g�gϘ½���Ļ9fO�o����g�%¾���D��G�9XHj��͐�.�O�^�VZV�k�Uo��g����7��o�%�ΛׯM�rˤ
�U��ߑ<!yf?�];�m��L9:J�� ��V�e��Tk孬�D>��Fޙ��Z���یH� E��%��z��;S�ل�/��pyIT�7�:�1 һ�O���I
��Ҋ5���>r�[H%C~���]���s��W=F�O|�����/��#|�#Y&�E�	أ��^�;\�㴦�^��}{�,z'�h���D���b�2� ��H��9d�J�*P�vs��g۶�<�(tP�H�xK9��-��j�0�<�T��(
�ړ�Ż��@���`�d���a��y.*a='������ԉ�(Q�������лj��8�m��'zBt��oe#J,Y��Q�kʄ�=n�x]U�KZ�L�I�C�_!���N	C�b���vu�m:?"�}�M6=�Z��-���Dt�c���l�%<�2/�����-�Xl:������I���R���J ���'n��+�K�_'6}_Ҹ'��V{@�;��ӄNG���_��F��ە{�d��c(��ڔ�+����Yբb�BkR��bE�=���:к��-�t�cK��yb!ɢ�~t�5m�K2�Yb�U�d� n��]��t���\v)�H��m�Bb�2ڎ�(����'2�
�#�s�/��H%u�XW�!�^�1G2�����ʨ %[е��Hm��z��Ă���
(U�꾊ŉ�[;���5���W���^]]����~z�S���vg�k\��J����z�ݔ�����g����B����Hq��@V����٘]u������##�3i4�^�#Ƕ+����]�"�FB^�٠���U��Y_���>���A��;	���'�`� ��T~��4���a^2y�V�ņ�ɛ��x�\p��s���NЂ�8�]X��a�z�/��m9�`P=?�����v�(H�A���\]^�dr6m���.��M�a������6f�T���ALْ5��":�N=���6���N���|��@Pٛ�O���=	��
:Z��� BT�wR�o�Ά��q�7�b�9VY�7� �E����ܨ�9*��FD���Ƀ�jFK2���`㫣�dl�ܸ<���;���ូE��eB��/0���Aq
�� �&�)�1��,%�lu-�N���"���:������"�1�	0�G�Ūe~�ʄ,��?�gb���1_�8�ض9�L�M���/pP!9��Ž޲w~mR�r��s ��&��F���H�po�y��0I{;��q%�9���1�����{[]��W/�|B �P���%��̻��NI(<<�/��RHV�*�{��D��/圧����{�����'�<��/�ӥ�5���5��F�2�kp�������)� �ֺ"'��;fcg���Ql��������F^a�衲�o�pZe��T�3�����ީq�i�F�6��c�1�̖��<�_\�*���߇���")+��>~�>~�޿{��i�-w����Sq=��pv�ue��qg�&|����e��}��j�4�;s�I�Z�#T��z+dybJ>ڦ�a�Q�� ��X<R1pE'��h�z��Uxy}MQ��}����f�m�������{ګ[J�m��`��G_Zɬ%��F��}��I���ü[�ù��:_~İ?��YٯO	}����-���A�������u��*��|�e�/�v��4�@���F�:"[V��sq_J�����(���U�t�w��p.�?O慓�D�[�B��Y%h$җE�3#����pi�PR�Ss��yJ2��˟�_�}O����pWBeR���ی@�5��h��ɪ$��>;1D�P�D�XWI2CZ;	^���ެ���NL@�*��1qe	7\c�Hf��Vm�K�m��hIn�������=��c��
,j��.��iY�Ǌgl���g<���\
�`B_�E���ϔ4�Ϲ</�]��/C�����I����}O��RD�_�Λ5&���ǐ���ɔJh�f��I�Z��[��@�O&��j�"'Rߛ�H]���m�v4�]����\V�3�pu}.�{⑕���n4��d�:|��lCĳ��j����p��fN������a��	�Q<f������P-N��c�Z���$��WW��s%WSZ�\�A�L*릷�Ѷ��U�R�u��i��M�[�H��m 챯�&8��9���(���i�}����n�>�~�y�M��￧8�Cgh�F2�����{�䍟72����+bHl��>)�}��5���=����
��T� J�F->Xl�+�r���:��du˂��6�H�<aD�����ce6�7i��F�Sl�mK8��;����ھ��26�`5H )2Q��H��A9�C2��:|�����o�|��'�*��"��#�o�@BƵ�e흐��%Q������|��Mȯ+���@a@]��Ș�U./�m&�z/s �I�ӒO$��q+��'<Fc������7�5<7G �c�5WU�'r��"YD��6o�n)��!��)�"D.L\�IY��J����}��7cAg�5�~g�	�ml�L@��h-X"�\�{bF�om�!ٖ���~a�p]}P����=K:Z"2���)T PA����A��@b�*sU���\J1��1�
c�*��I�Z�O�
�?[U��:y���=��z%^�G�^�!� �.��/V�<��������8�0��7���a�����7/�c���J����@b){� �����v��5E29ߖ��Y������v<����M�T�֓AR݀MSj'�ymH�Bk�в�ѴH���?,Y)���tF���3[{��n۫PU�8r��s�vPn�y�Υ��GeJi���!4�{#���ÑC�|_��%�ޒQd�2'�y8�(��w���R>�%G?��mA�?�[6���Ǧ���s)��ك[2�3�}�=;ꨟ}?��F�0F'�d�==�{w�m}9�QH���d�Mkߋm���A�Y9�εUT�Xɡ뜤�m�#U�[�@�����iJ^��߼o�����5�Ψ�C����L� ͂�95~
�q��\U=$s`#1��-s�/W�)6k}��}��..ŦW��Pژ������&G��B�NaO�n�,A���_ ������o�?����I��{�X�4�	�K�ѝO��U��ű�I>���W�z���6���VЏ���$qs���{����޿��ds�J{�h��}T��;vҚ!?N7p� �����Q��9�V#$7)�{����ݖ�]�	!p϶`>)�����~ƽ�y?4@Cb���)C��?~�@^	W��Ə9�-��WU�����Ӝ�f�����p�5���Q�S��h{!rnc��^Uy��q��5�����(�5���%��Ǿ�h��V:!m��>S�4��ƈЉ�5e�`�],�V�%���UL.U*m}?����U��?b�u�渢�H&��t�"�$�g<�[�VL�_'_ז"��R���`h
?oS��u>��'�*�r��m�"g��rⳓ�˜g����vM���H���I��B?L���O��d��p5/��O�ŧ����|jhh&��q��;�to	!��������<�&��=D��H���Ȫm�i�lRT>yK��������a�ŀS��.�p�l@4�yuҾe8܆��їB���=��q��<�����;��SW����Q/��qRyÃd7�B6�w�U���4I��WS���*d�D��+�|�b;k[���|�_����ylc ���1rN��j�n�N���g��o���B�r�]��mb��i^�?~|�*��U��������R�
|o��f��QF|���b٠�|r�K��ɾ~춏|Ee͊7��� �rǎW�+�e�'C<����c�Ѱ�}����$�$�n�h�>�h�9L�FO�>*��?K�V�@�	�}��P!�?P�g�̶f 7?BW�� �!�٘�H��3i�&N�ǳ+΋'m��J6��UM���J��#��7�M6R�[U���fX)1yy�Gd+V����*��-U}7a1Df(���K! �A��	���ޠ1zfW�P:Y-�.���W/�x�Z{��N��>yBX������H�������1H��Y^��U[X�%gA�V�aB��dIe(�^�����]ov�`�vN�V/�W�`~�H8�(X�L���.Zꍮ�7c�>��JЀ����$7���Jr��Վ\)�7wt6��9as#!X%�vk�����8՘���m*n�3�S��N ӳىd(�8@vㇾT8���*�إ�˚+!X��JG�����)�ı�Z��tip�%���|6���F���ɷ +f`�V��>�`�i�����:��m��_	4IF��������zO���y��7�v]m�Ϡ̓R󏏆��9���V�#S��x�F:ý��	������m�4ۧ�&H����"��N0�J�!py �s��*��G5� �/����ݻ���h�B/5Z&��L�իU�q#�LT}jIn܏���X�A�u^GM���$\_]0�!����{�	�Vl�|Ϛ�#�g�1��-*�5���q���k�n��ouC>�[��۰ᅑ�O�����3�� g�x�i|���������WA�Q{p��C�\Z���.���
m�P�{�Ai��/34i�^�u�n��oބ��ۿ���wT�������!���C�h��9�Z����&�Z\)OU=C L�~W�i[%q�rN��$�\i�
� j]�x[�Fo~�;_h5���LH	��{��Aؙ��.|�m�%d�A�j<jLj忣��w�$� �c�����G$ɝ4������Pۄ��NR���9<�8�5��s�6������tX��ԻK�C�֣ ��2���Bܙ��vcsE�Ô^�T#Pؓa[1!�k��}�5Qh3�*_o^���L�@���7%�J1����>�/@����q�<t�,�|x�!|�����Ka޼��k���|v��}���7E��� �ѿCQ�����B��D�
�P�[^���	�=��֮��D�����1�ة��ڒ���{���Q�O$]Uڵ���KP0km6�}ƿkk����؋Dc�=l&e�^�PʫZӍ��I��G���D½FƎ�=Cbd��w�g@.ݢ�|� %�|M�-��,�]���_�W+`��֍''=�<v�R�Js������i*�U�ȬQ��5���VV�	���k���G{��;�q��~�H(��`��w��,���s�2~"
����ċ�2"|$�������y~�J�9�fS�JQT*[��y$�G�%#�rD� -��<��Ŏq���1�Q����aQ�F������2��9����wţ�0���ҁ]�JbT�QJ�~�?�3*�k|�-������	]u2�N�o�qoX\z���i��sE���wA�+ :�������*}���H��,��d&��TG���D�O$=��:��߇닫���0����n����Z�I���QD�7�L�"��G�˅�n��S�����8v�d��{.�S��E�*v�XN|��y��TOo	�+%��S�PB� T�c��f��JC��(���?�����V�N����׌8~�&�	syu�*&H�lP�K��䞑<�MD���;�����h����CH��,�������z���}~>���ۮ�ﻻ.<os�&9��ݰ�[C��hN�W�dЇ�\O6�����=�X�=���T�<�WT>�����	�����(@������f�Eɤ���z��{�@u.�3���ϧ>���Ւ��c$ė˚�i]���;��Ě��$� �B9��I�|���n�m�⎢�
�Db
����rOK �@z:Q5����}�Y����M��]�wK��S�Y��ȁ{��e�'a�m9fF<��Vv��@U��}8=�2��<��/�	s�c=�y���Z1!�3�`��lx���IC��Tq�Ʊs�Kͱ����bq�V�I3�����X8��8�T��Ul�b|��b��hJw�o"��r\���>�5���	Gj�j8z8&��Hd�;��=���$�Z Z�ǂZqH�~v�D���š��˞�ӆ��_]_]�'�8N��/�1����Fr���bnoO�p�+�� ���:}��gI^���8����Q�N�)�e� ��T��Zc���;mN��ivv�u^��OC��'j�����`���HV&�q�Ϛ���~��u�]��v�a�����	q�[�W�߆�������B1�v=�d��R|�j�a$�cV�k�疵`)I��aU\Kڇ(M�e�*��|���/^�O�իW�?�shA���?���+R���4z�=�q���Z2\V=ZP���M�.�!��d��X�jT�)AG�'l[�u�s�֥��mV�W�Hg��3���r���k�S�6��l��D?bL�����>~���m� �,�9��sU�j�%3Ws4i�<�y_e�>�(E�`�0�^���{�]�;�_��=�E�M�T��+���.�86���34nUw�hR"����l��=�>���K�@j���
L�C�#!�,��D� �Gym�O��'�1���w�4'���V�i�m-�3��4e�[	|��ڱ�8�^��mH!vl!bb�F��+��
 ����F,rT�=W K,�`/幡P޷컱�}R1��₵�ȇ�����~0~@��@��J6a���uB��y!
F=��߷1ޖ�c�9ܻ���j�]o|.Jj�`E��B�֐CjU��j|�|�ށ�����";TP;[5^�&�13U3GV�,�J�I��H�(��ڙ"}��s�b�TWS�\�	�,J
������3>���8��:�Uؘ��i�V(�R9���%�x[�Sh�P��@�0��}�e�{�Ww�p��p����{1?�r��ص���m~�Ԓ~���Q��4(�f�k�"��lW�\+���WJ��LG����?������g�ś{GM�Û��X�u�/��㴷�|�1ϩ����9���B,��a��.�gW�J,]9nt�.8I�֠�z[̇9-ګT
Oxh�W�,����)?";`{�8�:ƖX;l�܊��U��Ӽ�f��� ���oއ*?��a�������]{��C�D�d��q��ٻ�>���}�g'�g��6���������𼆹�~?�|�Am�[�%��=x�A+�V���C�,у�np2#I"�<1�[!Gpc��Xq�n����CpN��tZ��'���.;�$#ۺ|b,���p���>���v'���'R��w�J���!2�vۅۼq|��1|�x>|��n�7�i� EDV:��ו�#� 5ؼڟ=qt�cy�_�%Ar[$
�Ȋ���TT'��"�PG��W��O����+��I������bjd��8��]�!�'���-����t���Z�W�{���Q!�2����]F|1�Fu��~��` �<&�3���jŖ����C5�@u��9�����G�5�}��?��D��uV	��`��IO6rb��7cuI���	��z� ��ٹ����)�7L сd������C�B��r&���*+"D�����eb���$Nbr��-U-C�T�%�Y�/	��&�٭xoٲg�@�D����A�\�R�
8����gB	xr��]wgo�����b��k��Qan�sbֻ{���g��������F��Â��� )��U������·SV$�'����hS�֠ ��1_�Nb�dfD��ih�����r�B���vI'�k��`�]�Fwm�u�X���Ƅ$�3�:�����Q:[��K[e�;���Hg1z�"}Ԏ�D1<m��=�xR����=~��)�����[�B�R�1э�ql4��Q��5ނ���߼��>x�m$o������չ%Z��
�s�۰�cR�jW0㼶��X�-1��u�*���σ%w`�P��T�kgj�|9�3��hm�tH{a��:ܪڈDk۪߹/��lj	U�^��~��{��U���l���]^h_D�⒴Ly�1B�X�'�U�	)��_tF΃�Iz�O}r�=�,��Q��}|I�7�Rv��C�,�s;�)OV�L���k!���0����u;*+� ����v����D'��
�1�'[�.j&	NO��e�S���!<a�62��:�5�Љ������$���	�X�9�B��r@O������ϥނy�a��kA��Zl����HC������8ڙ��V��W��lH��z~��$d�Z�PlY���s���pD��V'��rvv%dL��iŖ�_o*����hwޚ��+OR�Ta
y&� n��*�����p'rw)�&����]�cd*��Y%n'QFa��"�
�����?�^p߅M�F���"�}~q�Ď�kS<b��� ��&��SuǇ�$�3F����yW�T�8:��]��5�}{��"̈�Qa�9���iI��f]
��� �o	G%���
sf�$�(J�:��D�\����Z�JA"zr�(;B,-Y(x��tre-![+��y�J=��7|ĒЭu>$G��7O� �g�����&\�U�2?sh �� i��d~�Ea���i��|��<����_�|�?��
�.ע	�x�Vn��	��'��4����κf<	>��!�1�X�GE^;6���t5�^��g�����;��YhW�}�]4�Eb�������������w�0X��R�
�MBd@S�������a2�P��fՆd�7+�_n�oC�~�'�y~�*��8`��H<�j�/��݃%u8yS�.�i�w�b���W7�o�D1h:z�w��m�+z�w����)d!��]x��.o��w7a���`/?����9F���c�5����ת7<b���k9��'��۵�Xz�TJ@�1~��`��'V��ߡ�s7Q����#��ŗ�$�c~��=�#T{����۱����Y+��س��|	��xrI "�;硍[��Q^28�'w�M�+���!�[c�͘��)��>zՔ���D���X,����U��$Ԇ�Q�7����p^e烄�Me��}�����ps��|H�����|�@[dHl�D�}]C1�#�
OI�G��g�	���Mq^�!��]�W����y}�����-�-IOg��s�n� I�`�)X��TD�ǿ[���0(9�m��4
Z��Q���_aȣ�3�:�-�/r�Ȅ5�pX���qD��Ў6AYKg�I��X!azqv*�r��z���#QrCW6(;-$�v�<n{�j
�'ԕ�j��T	��0���R�p�h牡�N��m�/�5g0��>C;J/�d�8?�9_5��PQ�+�1��=Ȫ�h�f�wGu�������8r8��u8pʅ_0,��<�a((�c ��m�ҹZ+�3.A��u4O$��_L÷��.�����lm�I�>~b��5U� C^+gf-&l�6���tH�;��9K��ҫ�Rj̞$C������rE� ��f�TI���yw��ػl�½�'������#ص˫+K@���N��\If��6
M8_�e$�oo'��^��ш{I�]���_����8�G,�+-=�1v��[����
Lު�����{�_?���{���������H�I߻�!+�Gm��E6&�B���L�I?g��������X�k�*{#�H<�`�|��'N��u�������\�֖����#[;q;�?JIG"�qΑ���&$�UB�<'�U#���{�I�j�"+�4�)+V��s%�糓�vNy���wK>��#;\z�$=�����m�-�c&�gX�v,Ha���	S �N</�����g1?#;)R�ӏ���
J|����V�ނ};��0���N�vOO41lEd��/p�ޖT>�ٔ���X�Ga�D����;�I#��9B�A�E���
�s����>-�7�s�~d�X�����oC<0`4��i�BL�|�<�%��L-X@�\v�$ؖ��Oz���}-�V�F�B�4S�:��e("9S�~L�_E4�T}��n����(�P�Lt��Bk�|��@Ԗ��~ۉ��3'�� �a	v˯�s���R㝞��k�CŖ�K�Z������*f��b����9�l��HV��={�fr�V�?M�dq~g���S|�5����ڎ�}b$�m���x��I�az�f��O$���U�YvK�֡@��J���Ba�t���������9�:�7ڽ��K���F�ګ=���H��đ�x�*�[<�)<q�ܗ;L����&�������IE�zD�9e0��<�t9��|�)��9@<ɛ
�C��LĉG	U���#���#��6Ȕ'����W����9:��y6�C(=<�j��'�h��9��|mU�,cz���*FB
0���a�6���F�2$��,�a�Y�]�6��M�7���)]d��h��..cVn�9b1�ԟ�8�,%�P�/�zo�o�艐b�75����#о�dR�6@kx���cv�ԏ��ip��T�`�UC�	�X ~�n�"ϬTA��9{�����d��8���+E��$0�������㪀�ｷ��al~=��PG�/T��D��N*8�ʔXl\-A�@_��ΓOP�(	9J|`~̙�2�a%��fc�Q�;����ϬϽ�%2�0��Qd�hA�Ch`�\zpE�%AŃ���9!�j��r�����V�|�7��[T9�+9�w7Bi&^I�F�r�4��'�X���6}���N��擼�������xb�.U%Z���|{XY/���{�T��n쟻J��w�X�*�H�ft�.ɫs��0;%V���|�o��6�����O8����`̽EE�ÞmQ�h'@�l�۬{"���Sa] 7/��@�Qꕼ+�|g�M�d�n�"�+��8�6mq�qΘs�Dmcx�+v��d��mH�%�Y�Je�ǿ�c��N���+v �1����IC���LO$+�v<����k�g�(�[�J�)���e[�T��������������/��/��C���ϦZ��`�Y@;�*�35��ƪ{lä�e;�s���D� �����s��B"8��E>�-���5s�%P�G�dW�`r	d�v:�����x21εH��>X�*�q��2�ib77�l�F��E0��Q������$������9x89����%?�X���K�s������J����hvʏ��t<i��W�/����;F����P��vI%�k�(R�P�%�vJߣ�l��{���]��D�a/�ب=�I�]�7k�QI7%�ek�~��;ð�R1�{��v|������P$����ޮ�-���;o߱�mR[;��|Q}�Ч䷚��Ӌp~qUZo��'F�G�	H�V��ճ�a����}.�VN���Ub��tLi�68^3H�;�C3�s���]�[�|������w�]\�Sm�=��7<φ��R�r�
UNr�W��O�iK�5�d]��W&�!����nʀ{:�m�LΈ>�N���ݝ$���!��D3�R�\/�me�7'u�n�N���߼UY MNU�V[�6�ꜞRyvf�N�[k���n?��I���te<<n�-�{��3��Q�F�S����(&�����#E�ule�˷%�w�&� ծ+ƀI�~l+�N�C��{�E|>�6��k��z���*����-$�ĉC�8��c�M��-������	ݜ�'��R D$/�!�IFy�yD=)#%�$�����WH@c�iFEc�ލxwLQ���>7Ϊ��/�ϗ���ûw�&����/c�~�"ۈ���y�*��ix��u���*|�e>'tȼ��N����X�����q�g�-�[#,���G��a��3o�˱�|�LE��|�3���a�����6c��0� ��N���G��iQ��ٹ-2���"��m�]v�Vd���w@#�u<�~@�
��8��Y���zzUѶRbo0@�I��N�m�>F8X~1� q��T�8d1a���L�$��}#�*�d��R�U{m@���n��JR�܅񏃊��D��ތ#+s����~�h��l�J[S�~8!�I
���+����(jTA[n�{�����58M��
��	�՜�19m@�TJv������R�y�$�{�y$&"h�b�*��D�� � ��J?[*U(�RZ�W0�|y�}�DG-.�`��N��@k�􄄙�7��uZ�u�����Bno����IAUg�[�zﳱC;C�j]۩�<��6�݇5z��D��:_�� ,}���a�T��iTI�V��c��j���L����yc�R*n��ԜDrN/�Tq����d�s��RgA���p�E��Z���}p��I8|jû���T ��|q���J=�8Wʳ.��
�3�4{U�W�Lň�\����̥��Cћ�m�������K6I
T��Fr�:�*��O^k���TA�۠j���zk��	�$�^}΄s�r�cm���a��o�����x�����]��^���=�m�j��!�ӌk.�I���ʰ�q'&���~�]�y��li��`7�i/�~b&�=b<xV����ئ>���o�QG��R���*%KdT�J��(h�Sm�	������y����!���9u(��U�P�V)G����ɞ�F.ܚ*__��+S�1���|"�rQ�?l,�����N~����~�ƐG���yFtܫ/�b�Y{0�4x�}����|M�,��}訮��$�5���kql�u���"��.x1���������sF�li���B����9���������9d9L���Mi��b��)h�`~ᾆ�{!jwBb��)`�]$-�Bu��X-�6T-��>��E��'�R$�ىT6�;(la?�����ҧ�(Qr��`:(�Sn�`_�PJP�V�];�Q˴G,`�uQ��S{-K|ژ�2&��j��ٕ'��ж�$�ԊF���&�9d���I�3��_#�?�m�\|/1�'g#MV���~bx��_;Ǫp�n
՜��gO�R E�j[���wP�7�ɜI$q1����5]�#
��1��Ƶ��\��Iev��5�g$�P�$9�tN#TX�6�9!�%�u�G���n��B�Q�Y�I:�g<5�B~D�Ƀ-[i.[^p��w�|G2�%UH����"�y*D07Ώ#40���yF�;t#���MO�z,K2OjKj�7d=����S�U ��C�c۾r�fi��h]����-������
X�Ԙ��*�� �unHnSp�#���ڴ���9��p~�`W����j�������<�U,��OԊ7� 9��n��Ue�fU�d%V�y~����fe�s�v�<����ds]1đQ0�J6��(�`-n�r�p$�fgD鞅Y�7����|� ]i�V+k�b�AȝҖ5ξ�����_��=�a͍/wx���O�|�]m������ʒ�0�E���Nh�ؙ���Ԥ����h)���_?� ob�lHVjAp�j�����܌\Y�XKiǝDT���@��H�@�_��!S�(�.V?bIZ5�[�q�FU���G�I���`�����"�`!�;(c��A���;9���bۻ�I��I;�
Yua�$�LDAM�{d:L������2yJ�؊�Ax�9x���B�Ley�O��ᑼѣf��f�  ��IDAT�;�@{��Q��)�����!���*%y�S�1���������+�Zgw۸�,/�	�ά��PI�\��d�j�ArD-I�xc*ĻR%��v�#�*a�P(wLqz�d�H��R	CZ�yr�%r�ݏ���g"j�r��f���0�<���y�9�	���k�{�:����ڧ�v�=*o��GOޣ�Z+�v
$��5Ib��f�c�{*Oe�m�[���z���Et�[�1G!9��8H2�I��'��Ёz�wv�G��[J7Z�Ȅ3�`����������V�;�t�hpERk�O�|mԺ��3+' Q�<I�2孵���6���u5�(%5rH�S�n�R'I�DT%Uj&���R˞=yNMKk��F;��Ax+��W<���oε��c�M��Ȧ�0�qx߀�a�Ҍ?<:�'���9�?��㟇gz��y���`O�l��H�a��C)����<&��Tȳ�������1��?�c�����S�&1��˧rO̯�suu�*k�*�̘�B5���V�`m��,�K�:�E*���0ٰG_����w�~�����P�hC�_�����o���>|�޿����\ϫׯÏ?�޿G��}�����W�l� Fm��N���L�p=.�L�o�+�:�9���+���ڸ���Äj0�p��y 7�����T~�1S}߱c��ٞ���|l�=S�`�Lj��l\��:�a$惀�������G��#t�6�%Q<3r���n[�lT�v(����(p���U-B`p�Z��GÄdEr�f"�@\��g�+m)��ȸ�.<̝*��R���Lx��)�=TL�,����oǢh�s:��gG�
����'�G�5{&���U�'j1oU�g��'D�B�4�1�|��ߗ$���� ��NE�d%xR�u3���<L�M�c�L��(�L-iV3�q�'W=�S�0U[�Z�F%>CC43��H��W�m�i�G�u\\�@a$D���&��ij�t��Lit���x�@��;��~�◶���ɉ�]���)p�P�!�-��Tg�!�����&���D�zWs�B�N��ľ
X@��H0�.��A��d���$Ǚ�ԶU�i�E���$�p�p���>F%�a"G�=����~h(��l'S�k��LI�PYWA���&��]�d�q��.\���<����7�v���J��2�/���lͯ�m͗��,�sb��q@�iynm�@$�E�s�D��ۻM�����w�����vh�/^p-�����}Z �.�!��1d;�2��l� [��ٔ�D�P4�́{l� 0��ox�y|.�ʚ��=���X�}G=���r����C�����$oȲQ�f1�S� :e��/?�!�������&�v+fh���&���aن~���;E��ts4/��D��:�t�<���m!+7����!��(d���$���M5�@n�6؉��Z��7:��<6v�(i�'����Sm� w��M4��}6+zX���T^?���UC����v;]�?y�2t�C�����c}\j��J}ڒ�ru��6�H4ũ�ڢT�a�'�j+#/r����f�1�B%B5�v�l���	����lJI���m�|ܲ�Jh����#�Q����zKpy�M��ޫC!>%��[EQP�9O�N*E]+�:$k�8�����KS��8!bmdžah{�{\��	��o��6���JJ�QF{'(/�_��*jp�ھ�ߥ��l���1P]��h��l::MꥏA��5d�>���ޠ�� �����4L�A�o��Ϭ�����}�L�����
�Ne^�wʽn�W���E�nno�&�H':�����yBӧLqN˫妶��1V��6`�E�H�
�ꋷ� I���9]�@S�8�&҃C�èᬣ�z��f[%�v��1�rum�&]�=b�����>�%��yB⋏�}+ߒ��I˯*���ގ��`�������Qx�k�8'U%]h���VN�;�}p�_��N}8�>�ɸ8z�ND��
�U���c��'�;f��z��:��nIv9iJ2	l�_������KV`����?�)��|�u-KΉ���\I�J��a���,3�j[k��!��v.�|���ƚmYF`̟Q'�
�2�f/;�y��{8���Y��L���}��/Y�CѨ*�pcTy��J��H@=5�/�s�e݇��t��~���z/Ŧw�;:�}R�jcI��c.�R�1e��{;��<��y����a�(y�{���=�6i[l*��T�B�Q�$o{24��:HvΟR��?�Q�����W����L2�w"�L�/x'�)�S%`�]Ūm�@+|�A�=�m�(�L�����J"R-X�B��$G���pYXD
���N��ow>���A"�bb�w����Q��>�O#���@�}����ne{@��k�v(G�j�@-T�s�ɖT��s�0l[+�׭�X�6��xn�̨���pw���m^�~V�����[ ����ji�v/�T\�����'q* ��\�:!"�%���H��5I��H��C��^��J�@�h#ޤZ*�a��M�'R�̧�����-i�"��UiL����a�ַU=w����۾ꒄ�����e�Q{���̐i���I~������'�|w�1Z�9���vS��5�*(��Dl����8N��Q*x��N+C�|t2��}2��y�}����Zq�i1����j�2*���>�+E�G��V��}�PsO���vg��mş�G���/�Rp��-5�UR��;m��-�4�.'y_��U�ex����|c��5����Hџ�Z����(��X��G�꧒<� �ue*���/��P;R�����-�K�ז�e�佶Y	�w:h<����C���p�����E������_�����'r�xj��� j	����ˣ�t��i��w�[hy���{ұx�>dy�A����W��>��2)\��m��錜�ğЯo���}�Z�����>��?���puqM	��R�-O��އ����+��݄�/hW����-)ؐ���e��x�˖� Nɋ�2;W/%;|rB$P��P~��4cX�h=���n��q��͛ ����
��}"r4&uh�f���@`�j���;��1��H��P�l����'��TU��I��#��G+AŐ�)�,�Enޱ�7&�ȃ��;������L38�vE����iA%a8Z;��8�BȡĽ�d��B�4��f�{kD_�@;3�M��:R������l��;W
8q�P�q�@���� �ْX��#�'a�JU�Ƚ
Qbb�f;;�`���C���z��Sp��ƴY�\(�5䗒q����M#1���?�����j.��'DW,��J8������8�as��Ո�oK��e����ߕH7+T��)Z��8����h
�22t���]�ދ�����}�C�_��5~��66ѓ��:�ل��B��[K6�����������cqrNg��tβs9Z8@�|PVYY�ʻ*Ck�g@dATۙ�#���p�M=��MW
)�=$v��c7�`!'���y�'����:9��ه�Lʨ:�ѓ*���5V.�iz�s�������Q�'jMV�݋�f��y��f���6��n�r�������'7�\!����!�ӛJԸ7�Q�c��^~G�l?0o$��6l��q��-��ܷ��wyq��o�&lW�����>���9� �ڱZ_�+���,�	�VWF|ٗ���+$"���tX1Jr�!2�|N�s4��nI�VN�� N�tΟ��#CH���H$njs\��!�/������Ě>�A�?�˿���1�IC^��<��>��}�so;�9�^��o�R�R�����e��B$QIj;�]J�`Nr(��|bw@l�$�۰��B<}d��у�q���A)��v�G���O���dO��>���A�q����9�WKCq�?����8y,T.�ή�k��VP��(�	v`��Jpj-���)9D�X���{�1�w��� �����V�*�����
�U��]���n���û��S��z����a�GW$��q��J�`�.��gŏ,��*S��3.@Yy��b
�n�GE&_n>�k���;1j�4� KV�+��+�P�R5^�^��.�d�f#*�>��6�;��j�
��(��'b2s��q���e���� Q��/5<���&�Yq��Y�`|���!�쓈cK��`�O���h}R�×�����*ʧL�I���?�>>�s��[��O�&Rbw��5��cQ���X�?�"�^6�r��ǕMUP�f� {ڔ�W@ϳ=<˶��x1�Kh3��,���k�&qW���g@*[+UA�v�%���B�����(��a���:��"8��[S�M/���Սg Ԟ^\_�����#�ck-r��:+DS��r����ؓ��i4�~x,ŉa)�����z��u���{�d�X�ALHB0�ɸn�X�����$�w����W��߽�߼���9���)�?,�^;�6<��*�Ι"���i��i)�t���*+�gũK�F	aYw�W��|�nwUI� �DlGP�]�cW��8�b͎�G&d��2ۈ�ׯׯ���1��?�5���U��A
56$�'�qߎ��#.��?z��ὣr���Ņ�/��G��p0�4'ځ��ޤ����~��N��]�����IFP�7���W�����j��^�m
���������E�_a�ڗ�z��+�����I�����d�sbls���ce��qv5Yg	@|�rR��*#��/�I,è-���Yv 	��`�*f:
�uׇ�����|����:K��$� 1�Ҽ�����i�#14�ŝ����E�u�=�	p4��NM�`->�#V�g�b?�!��Y�rRL�{_XkS���9T峩�[]>��/�p�{�r��ƧR~����%���������K$ă!���L*(2�7ƅ��U���pJ���{M0�2)���������X��n�?�6
jǖˮ+���E�Ag��,V�~2��OOO^���K��1�䉥|���q � dA��s%��xC�Cf*�~
����	�7#{'�C���)|�H���5�ɩD�VReÖϝ�V���QITw��Cd��V�&(�f�ITGq*-"���T21RʎD������
���g��4NL��q'ɐ>G�?�f���`ɎW���w�sď%j���7�a��G��aq��}��-�i}�(�=s�DGcvB�8�b�Fv%�������[�'����HȖ��s"`�ߡ}
o�
�q�s����Z���&��(�w�����[%gz�ƨ�RA9
&�J�V�|������1�����l�B[U}�K�y�%�̳F��D	�WѰ?�8�w``�L�tD��IF����J�i<�x��e�:;=/^�/�����c�=�I�lA� �d2eɞy�3{ξ��Cv�~�O�g��Kf&������{��E  �̪�7^���paڮ�H�N^y���Yi��z�]�Խ��`Qbd�㧗���j�<�R�����0N�����n#Z!7T�H��!�13��P�*|��(&�������(^��X0@p��ٕ�/�ܦ��UiWÎϲD�p��nk��n�7���K�i���IE�~p�P�z�Rs'$��u�{ƛDR�n3��rz�hj��w���Y<�7Yŧ|8�:���L���2f8�^��zx�v$�����k��|����݋�B�"Q,5+e��t���<~.�Cg�[@(��c��a%�k��Ԩ#dP*cR�N)�6�=WN��aFm@�1R��UtOg�w�S��2bX�IxD���E�z��rj�h5m�6�K��Gq'�%0�N"5-�Z��GeO1�G�D@�WġBT���7��-�R�����1Y��+�e_}����N2	I�lk�Ez$��_�xR��7^�;���JU� ��4+bs����ŋ#��ׯ��_�q�޽�|��Dѡ�0��եaQyj���UH�3�qw�Q�Rx!)nK�\�!G�� ��1��#p}��1�EtuJ�$�+;C��(�)����q$�|:�y�R��qo�1����TI��t�;0Z*;瀉b����}ߕp&Oo��gkƝ����x��N�?�mp��bm7�)%�lp,0�Ɂ�h$QK��=R����c� ����z�,%~M�4�����ģla�w�т�w�k~'�Txt����V����`��	��	F �����{�ͷ)G��ꣻ��#C^��Ը���������w�ξ;;_��OsV� -Ri<���x�&�z��ӆ�ʃ��!����|�Vϥ�^O��Hi>[t�l	_�N�kcFj��$�X���1OaN�*�K読�PrL�1 ac~YQlhӄJEJĭ���@�,�z�P\���R��ܝrp���QB�������M��k�#�a?Bm�ڤ���Z1p[T%m?�M�̨S���'I� ޏ��DOԸ�
e�+J ^S[8F�JFGY��@\T2-�_<+bX0����W:5ұ�IO���"Ԑ#��+���o�8�|x]B��+�Ч��D��^s�D��s��l�lR�\#Ξg�y��b��I��Zᕭ�k3�$���&r?87y:�i}6�!�4���xĒS�*�}ޅ�&��`k'E<�31��z�tA}ԁq硾�X�Cv�~��L$�Q��ϝf�zԁ�����
'mc�L�+�"��a�9��\�$<3[;B�{�����I��D˭�8H
�2�d�d����TaD�����nog����NO^�f�u��4ы��WЧW��Àz`�K�� ���[�4J�2��;J������!xD_���WX.�ǎx�x�Bv*qea�"K�Ȑ�e��iޙD��R���l��+�Ѩ�w���/+?>��^���\iS�ɲ�T8u.;����ܕm��`�
�M.�g��<Ӿ�̕������$]����ϩ<ţǙ$���5���D0��O�����^��)]��f0����Z����X���A�i0a�G��q �l�%c�7Ǿw�r�kS/�S��߷d� ����b�X
�ɄF�i�!�5�������:dZ~g��0�H5�,���)T�`��(��Lӈ����7I2�W��5R�$��U���T�B��,5?%�	1�,Y�D&^"�!�ٖ�`����,����v�j��i~��h�<G�*Ҳ��b��wQQ}����/^�6�oԈ*�YwY	Q��sbFvK)-��FpO-����mS=��=CO�VY	�0h��3MK"Ʊg:�NЪ�0�!��X5�=�2�o���}��{����)*�"P�ꚅ.��c!˂oq-Ԙcwè�qd�aH���5Պ�š��h{��"�W#�i��!�jk:t��j}jd)w� ���������Q�G����S�^�x�_]K��8�g����!HҝKx��>���A_�P�䖜nd��l���u��Ն��l���#ĥg�+��$�y��:c$�	TWŴ�a�� �����{�IF����Q���"AB>o�=T]�����UV�#�k��r���]��U��ÕgQx{��}����9���f�YJe������;��w�˙;�����;���.?2�gy7w�Q��g�zmT���h��-�4+;���{)BBԠ�B ӽ�%L�v�ך���#�+e1��I�A�"]B1��׼uZR8oX�s��Mףb�O��s��?⛱_��w����Z��l�	)B��ҟ�5��6�1Uj�{�wO�`��:+;�\rt|�N^��G��3�h#��ûѩ����s"��� �
U|��I@�����:�>\���d��r7�r�׷LA�;=& ���dB ��a����L�b �R�z����kE����M4A�ק|Q� �z�Յ�q��1X2�U8��=Q���E�C.W�<}�XN���Iq�:3�ۻ��.﵂Q��޸�_��
U:�IA�)+A��6���RŲ0h�m��T��h��H3'ƞ��V?N��I}�tc�r�����74���b�)=�q}�x�6�Qc����ѳ��-�3Y}e&73��7�����R����6��C�[*�"S�����:�ǟ��f<B����=�(�7�p1w���%���m|n�rǾ���o�&��~e�U�"��� i�MU&��`�_�}%P�)���]&�T�dX�
0y�Ut~�V�S2�Z�}Ec�ۉ�nj�Hl2���sdg_l�G75F�҄�<�{�>'ZmPs�>[c�J�4��3~M�H�nӠ<r����d��t�	���I�Ѻ/-".U�q����YIqF,����[�h�g3�8oё�-�	��fĦ�S�2��ĵ�iD��F���o�:�t�Tn�gP��ok����i���zuB�_JڑD#�����b����i5A��#R%��72ƕ*����ݰ��I�K�������gL����4!=��U��!ډ8�Z��}DQLgb���d�Ob�J��%jj��b�X*L��%r#���B�K�9�yMMQ�TLZ,�!&�-�o祲�9��ްQH��,#���z��?��d-5�Rf�%�j�����Z���(D��d�}������w�O�I�M��Az��3:i��}��Gw-e�t�t�(^�45�a�V&�c�Ҡ&��R4�!X3�b�9���
����x.2Rz����h��{gA\K��;��1���'(�J[0��E����W�x���#Bv>GB})��|Sn�3�p��V��ǅb��	΢0�WҲ�-��[���>M섬��C�c�
D-`��{'�覨�!�UD�@� �j�%�����Q�<��`us�xˢ�0y���9C$i���f�!DԠ"�kE�mB�Ӹ���2B�xT:Ϗ�����	����sg�nȬ�� ʲ!����+w���ґ'����칋�a}b4Bݽߡ%4��"�%�[�:�=٪��0Ԩ��R���g�ݦ� ���Rw~���w٨3�0��cp��#Dd� 5�Z	�O_v�a���3�cr�n���+��>�_��ŧ�Q��e��$2�����.T(A��B�ė
T�ޣ��K��#?��N��Vm|�Žݸ���F�`��}'�$0� 4ʤD�A�!��˔�����5��vea �B�>�l.��O�a�}284,]�CL'` @��������[���y*<E�wTC�Ov��i&�����RC�;����s�=���|~�jqZEfh�QA$�[+% �@�!��=�r<��*X��<Y�G�"�	׍F�&ߧ�ʞ���"�I#�GXK��n=�Z��SqD���a�`�R�^z<�ERe�g({�HE��T-e�g�V=��88�3G�	ƃ󒚵ԊA��	��#��#P�m����n �CcA�F!k�4��4��#un��*�,W�/h�B5O��m-�pggg�J	�=w�ܓ�R�=ҐF%����� ����+���ruLK}(�o¦}�R��s/F�	"w�~��,�jI`#'�^m������Z��PJ{T#��>��ɘ����`�����h�e��~�x����R�U�KE!/�S�n�!̾��SI��K;r4�t�Q��)�2+d�\��ɺ<D��|�'#�uǢ_Ű�İӛ�I�e��tK�s׸d��P6q^��J��:\��������y�H�f�P�h=F?�V&���Jo*�xF��>���kXgp� G���;��pZ)ՌRu	�󎕻�4�q��I����|��YO���˄X����H��I5�e1��-���3+�0�@����v�~�=���H���Wb��"�k
w���o���@�Nz�gX�@(�e��=2�@`�L'�xKN��֛7o�7�|���;w�yj//?�Q8���Q�yBZ5���N�9p2\]����h�ה�@�Rψ�)����¡�U
}�O8g$}OR�Vʫu)h,�����h�	�=�B����jt^X{�ZM�}H��#޼z-���a�CM'�W�O���V�r<`{&��m��T�<.ɑf�Z7�غ}��@��3pL��戯"v�ò�m�	Lx@�sl>�߆xm����(��3��_���F�k?U������8����p1\�^���wu~�Z��y4���5���󅐞��T(1�g#��P�,�t
�_{QhD��񷇮��On���4*�/�@��+HJ�jy�.�Q"s.Lm�y�3�v���:�U1q�Ѣ4�I?ʦ�=��j������_���͗1řXbʋ]7�k���;c����4MUJ��G�t�&#�Ɇ��*̈́�2r�wj�Z�Y�תKd����!JT̄"]��B���Tfs��()z���I'�w�Y\уg���RbEvwO*r���'a���p3B������RP�~9g���leÕв�z5�b��.x=0`�$�ѡF`8�>��7�{�z�=��F9�oJ�TG5�m�\���_��k%CSb�*Y&�%U��Jq��ϙ�㡅g�{��
"E��2�"�ƙ�ƍAݝBa0>A@hQ� ���0�ƢN�����-g�?�:IK��~�uw��A���b�9�;K���r�t@sGK�f��>�	��}Ȋ�~��=Zze��Q3Y�T���4��k4* ƕ_߿gx�90��q}�O7��ǒ��{x�E����:^��jx��x���?s�H���)�Dg�g���"
җ	�"{˩>q��P�����/KB�ujrXi\0~kUy�r�'�����ҟ��J�����<�j�p%L{3Z�Ubrg��8�*q43��тܝ�җ�a��.�}lqyI+3Iu/5��0>�!�'1�4L1a*�]}�Ҡ`���e��ߌ��t�/�+?I(N����Ѥ��X �W�Lj�O;iS��4ƽD0F��_�lDJ�J.�u(��c�5����:�*�ͤ��x[�����4F��B{64]_^����I+Jq�]�C<A�;�Ayh�34��0"����` ��*E���h��KT�8%:�Y�P�i|_-y=V�Z,�B`'�?���ԤH�����0���j�X[�t��cj��0To����L->æ#�'^�u�Q�h��X�V"c����l��G8TP�iW(]l! �_^��� ~�(��R�a�Q��� P��9(p��\*��/@�Q�Q{{,HdFI)��_{�X&����Ա�]#��BZ��e�OJ��K<X[H�ۡAgW�v��g�����< o�X#�����Ҵ�{�4�d	�^eȄ�ik:�E'~���_���|���o��	���ԅ�B���VJ�D�Aތ�ܽ���a�	q������O���^�x�U��R��ƅptp�.@���t�ɝ��.�>JI�6�L3��r{ά$��1~��'���g]D�V���xߝF(
s/ON���7(�9w�bXE�=i]\��q���y����$�m+���i����kB&�ڧ��DA�~�����#��2��C}��n��~�,�Ǻ4B%��T���'��TU��Ӓ��,�ĸ�Q-To��t�˶�MSۓ���F���oFE��Q	3*��OG��oL����J��*�R���"����I�VКk%� � ��F��9O�,�.����;����4pSF�R��-=1H	�(�Px#�Q���O�������5[�~.#�\������|x���Ph�[;0g ,wV��Y��a���]���������?+�-��]P�
߉�ش����`����=�;v�9?4�ͻ�}.#tr����,ӓ�g%6�)!J�8�XKxذ�㚻��q�����B��`i�(8��������h3�� �P��e��޲��aUL�m��J���A@R'����g!i��d2�����`Uu�q/��I��{�}�<Iz'/cgSI%c���S���L������(
�o�k ���c� �JIS�~��/?�L:���[���K<�q���V��=�K��r.�J�т{�Y^�F�/��NX|ci�M��uo4["�TS�,��^��ןC�F/�FiB)��
.G���2c/)������޸�RDG��l�����`.;N@���f��Hg;Wpa��2��eCK�:@�[}6��=��VU�����N����M&9}|X�Ό�#%,=������J���)gƗϒ���V-m0
��'K§�,}��-45)�b�Rh3�*��d(���sۑ�԰�2]���������������B
��T�1�pB5VD%�uw_���z;8�@�q?8ؑ!Z�4���b��;F��Ѩ㎕��5�t�UÜ�`�����פjw2���1�S7Sb.Zvz��{ɸ5�4�Ps�����@�T2������ѩqT��#x)��v��ח���8b.��_�R*D�y?��>��<�=�;�F�+O�b4��:sq&�D��>::��S� ��uE¨�񾹻f4M����M%v ���4�x &��9�us�	R�p������S��r��_��z��["��EGPAP7����T�[:S�]��T��q��t�j�~���-g��&J2)�5��AK�u\x�*L��w!��3��91$;*)�]��������{��{��ۉ�b��R�̳�ٴi��`�F���^��_�z�n�"��b�P�6p̢�@E(y�@;5�p��ߴ��<�T���S���O��_~qw�Q���0�s�ǫ;w��I�D�RQ�Ę)Ye������:epM�a=���7ƤmP�,Ǧ����za�^��>�?[U�P]2]o`A/m�P�-o���K˒0P��m��q�B�9��֞������6�[6"׷S�	.����8Ι@��u���Вk_^T/��.�xz�#�[<�R���[%��dȿ��3���g�Q�w���W���̍���J����bLl4
a!���A�/	�gU4r����ކ����%����/��n6ï�1��SRWo
�<�C~Ul���(#�8�_
���R��%=��e��90-�%u乌���y-n�$���JQv�8X����]���)�t��ϳ��r��VD�X��������>�CaƩ�gP�%=��SN�>�
k��E꽵����[u��aI?��MR�t'
����*B��.��E\o��^��!iW�a�wtZ�ŘC�Μ�ދ� K��8u�}��{��-S�p.��MG���i��mo�N�EX�����y���Q� ���)�6~�|��T�Js4
�ĸ�; �
B*�x%�́}�U!�Xx��㹸���X�U+�1��x(3��>�~�A�F+����ݻ(p�� z{s���g��$�2�ֻys��2�Cm O�ۅ��B����T��׽�^�r-?��k���^��eC]	�K,]�u����J`6���D�ՠo����B�'�"E�IG�B���Җ)rc}yTKF4U{�n�������l��>�;d9�ʩ;1�x�O����L�I�leG��w���E�M�I����BKAc�V�����,A�O���ޮ"y��������	+%<��
/F|���$�D���|3 �Nrb��J��R�ҵBm�R�"D� }��D:-S`�,hE�Tݯ�R�~)������2�DDvIf�ÈՉ�sFG��¡��;-M-Q�+��
嗉Ѭ��mf;	�^��U�V�*�� i�%�Lu.�Jz<���q��K+Z�����ެ��ݰ�\�4O���[*
r�����
*�{o�N��[�Xs8��0��O�?�y�չ;��++�}π�F��X��Q'���#�w`�I)m0V�.El�g��v�9�:��z�4���?�ƽ�V��`D��bI�{e�v���uq�,��\aU ��qF�v�F�a���L:�<�DE{�]wz��]��u��\��̅������L�dB����K7	ty�Ҧ��$���5���_�\��^E�`�y�П���&[��61��징�p%h��0a�qc���J A������'_�w_}�ph�g7����<E��ƍ��D��F���l#�D��Q(�����4*��W&��-���XV,�	��5҆�a �� *3l2v�6.������ˏ�����ٸ�Q9{��������P�6
�{������c���e$�
����l}u��"��ld	d3?��B| �f��&.���R���fH�c�&4���$�L��s���Lme�[1i��� X1���R��W��;HƣN��/��0G2�[�r0un\�!<�y֔�g��>�����|��d���u���oG����"R���[�"f^�~iҞ �E��4�@AŚt��U�iK�(��!�g*�a�d\���h�����J�t��B��3����-K�iT#	4����$����r�p�4	���r!�#�q���ށc�,�UOቑ��F=�ݹ&�$A�_�|#r�Ff��Bb��=v#];����:}vM�p��_^NCb2���p#"DR��!�{�����UL�*4��tb��0�ĭ���[fi1`��	A�����Q��%����>�D*5L�v5��`��v���G��5K���2M��He���o�w�}�z�N��R�ʀL�k���=�T�Y�>��v�� �:]��9f*"<�]䫍v�J��O�P$��Wx��sI@�7"q14�{��萩Y�|��{�l(D"]^^����:<���́�+L��Ź�������� 
¯_�&�;H�8��P�(K�~��W#��ُ�@{1����@^I��7Xv|���c����W��;�BZ9���'�hAٍ�xkH]��r��+�9�J�W(]��c{x�mz�N�y�H�
�1�$�K�X��o50<�eZ8���o:?�C3���,�0�9��>�D|��+S�Wb�D��23��d)X�A%��M�c$��<�۪#yF�����~��b/��xS����?�ҚJ9��'�J9�U��YIv��0
7((�t�"�P��*���㵦31���*y�@�����iUM5���cV�Z�G���9#m�td�?�s&��S�5�h���-u%���G�K�N5��QYg�h�yG�36?��"p(�mZZr��#,{~/x>\/�grƩ��<N#���V�����
ߩ� �*/��i]�5���{ф�#�����<G�'�Yԍ�ŵ�ߜ���3�o��/���I_�2�g�
@��d��|>w��F��7A�ͽ;}qJݻ[	x���CAǆ�pX#p��y�f�eѻ��뾈p�9�<��U^�쪱k����D�~��ʘ�G��F��wÈB��]|�ӣ7?�|;ʨ��]wz��c���z����=Q~�gK(�RW���ƌ��R�I�O^3%�+�~:���=3~�50�$OM�{�jyZO��k%�=5�4LV����/� 5�B�w�O�={��ᇿ����C���E�����W߸/_ƅz�~��g%b'Q�l�ֽ~�F<��e ��Q�)Υ,@l&b`�<�{�MJ�ݹ��ן~��JB�A�.(^E"��x��	�1f�By�x��'!D�z��a!t4z ܣO}ȫ�4�/��?���� d}��c�ճ�~�/Ңy����5�2*����Y����f�^q��~��T�:�C�;��nK�V���@�;7�zip���W�S�(0bO�*=9n#͚���vԩ�ѫ�Ò�3^V2A�����Um#��V�4`�=HDZ�N���:M�,�BD57���e2t�`��H!�ĥ�w�2����v	�<��T�f����C�r��F��@df�(~�u�UX�h*Cv��mk&(�.���4��ƭeJ�P��ޒG�e�`H/I�T ťW�	�,��Ɣ)����>X�A64�q~�B.M���Æ��(��D<�4,F�����#o]�(�0��� @oq�tZ´q�_�r���$�����J��#o��_��\�f�����PE�-˚�
!R�j�J�N�R����љ��K����B�l���DI����ۿ8p���///���2�8���'w~y�n�"�@����0]}`%������?h�曯�@z�^F�����S��Ogg�pV3�Md+(l��p�/�|۾���ݑ&.�
�g��ĬI6E�VGA����`�u��y�^e��d�t��>*�,I������×�E��C\�<s.;�
	���#e<Bx��릫�D���э(�Mʚ{�H���n0?CZQX_c���йc�킩c��9�M��F_���@}�-E�iD~�C��p����C����QH!G�7���wg�Q�P��D��1��ר%:"���D��R�,��(>d�m0��H��4Q�I���$"ĜUM��!�w�3��Y��u� j��'QV�;��uw�n��7���3_�SM�"EF0�KJl\'�;W�~φqF�S3�ʐ��±������`���'L�?;�D����>�}��K�eKg��8���0B|Gs�*s5��OA�.�"�_���)P1p"��bK�W9��
'Y�X���/�!r��1���>7���ק/����Xd���.���~d�,�P��Ľ<y��ǟ��p?����z�����vw��I`�T���֑���������T�p�&��i���"k�V鬃_7`�'v
�՘)iL�OfSI3Zt�:��w�~�������tWq�6��O?������l�Q�:�������?��O���)�����}:�DA�������W/���6^�_HcΫ+i����T(���[�D��JhzGR���_�������;�x���P����ӛ�wܱ�j�Q��S�2s�����5��ɥ��W�z'�.	4�t��|���L�?��(CN��ܲi�\ff�ϩ/=P��Iՠ&�2R.Ѫd��Z�R����V(T�ʸc�����?Z{||�f�9�6seD͌;J��/#�}dL$g�D Iu)*b�aI��R��zX�0^��C������Q���ėb��'�����O���/����>2�;2H1nÛ��FE���.$��k��3�����b䙢
��f!��'u$�9��*�{#nLq
؞HޏM���/���Z	��s�M2F�]#�6ө�@��*{	�V�Q��X�����I��$I;A�j|W*�MĨ����O�-�X:�3"�@k��8˞�H�ҫW/ݫ����_}�z��.���@n?�0̘�zz�lxU�5#�@�'/���CМ��M��#�K��j5*��F+`��*~����l:�A�Ĺ�,���L�B����y�� ȧ/^P�i5u����^V�;�
NĔ��{-���7����7v����`�0z�"���k ������������>�֡���͐��|��Z��$�Ey��7,��m!��c�4�!"��{��N�p[.��F:�������l��{���Γ�g)L!��d��q�uZn��Ҏ�5�P��e������e���036�>��=�>=ft*������.X�1Ui}�T�C�,�u�O�V�l]�|�3k����G%�Ľ8A�k�_�Vs��N��T�wAj��4�aA��N	�k��+�'D(;����P+�(!�>>�t[8�;����P��Ϋ����A}�shA]2Ff\
�����؄�0�!����}w}��v�Y ������0��Ӏ���$���:�2����ʚ�$�K�3�.Dj�����z}�ޜ��߾r��;�1�������/V�^���[��a�`�����Q��_f�D��@b�
���ݓO�R�J+x���FR�{�VY���&�9b���RK�c*��O�<�2dU�T�Bivv�(�"=�统�y�M�A��!����Ʀe'�a]�X?y��Ki��L��C��~�}Jyw�H�.�A��n��d�)��U��}.y��鼀��ЁP�E��#!z)!X  ����O?��(\�� ��2fWwQ��u��[w�������ŭ��5{S�v�+������nv	os\̫¨c�w����{44�9��L+M)��#.����_�_}	Ǎ�<����x�&�	�m��7'`� 2��?%���@ܻ����|5l�>.�z��WOCH|�|J7��CB�\�,�D!��z�Ͽ���cPZa�U��?��%Y��l��IQI��H�N��x�������y��D�]y��D�~�&R�Eф��J���~�t��#Q9�`vڡTu�*�n��Č�^"1:�S�yp+g鑩���&��a���@�eX�F't�"Y����|>�͆΢#��$����V�[.���� Ѓ��_�v���1n��+�~�=cvRP�b�y�ĉq�Ѵ�ZQ�4�'�MJ�sZ��dCd*��T�_׃�9sD~ӴI��R�
���uF�	�5Y�d�[���IF�� �sw���=1�0�ȴ:�ӵN���h��Rʿ���3A�P�R�M����@0fT^�{�qa�vF���[F�`?�,�����7܅F=�V ١f��#8 ���J-@ű+F��i|�w�K�Ż�9E���%�6p��m|���3!�K����7o���������ĩz��M쯤X³�O`\^�'�����A��t�/�����ل�Y>��:f�Q��w���Ǣ�@$|ܮ�8���s�l�1^�T���HTBwqK���G�qK7딞�����'\;Ohq�w�xW���yD�M�'C���T��|�<�3���2j\�yI+��ݥ��c�-�>OLw&[�����"Gl�,J��s�~�Ʀd0ӾRaF�(�e��[��r�4o1QN���s6/iP0���w�:�X@���j�������X����EF�Ag��4Zd"�h���!Xڙ<�}g�޵X�8�rԌ@�������h� P�r^VQ1-9o��v����5�tIw������0�Z�r��æ����8r߼9u���x�������Gs�/>E^����}$_G ��^8�&������ ~	�
~g�H��{{R��5 �ލ�<��p��g����1��R�5r��x���h\<ee�h�b(r�b�ny���c������0ٝ���>�#���mD�s 9EBv�؜����_}A��V�k�;�v��MC�����G~{
��.G;�^����mO�i���q!���I!���PpD�͇(���Eʝ��z5_��v�Ǜ���^ܹ��|,]��]\p��n�؉��;��i�����]NR�|���?"��o,�-�a�\iu���ᱻ�u?��#��]jmn�@aĹa(�]T��՜�2���lM`	:ק��y��(A��S9�����,�Z;���_�R�
�����mN㐖���l�I�V��������C�e�	�Hy�l���������M������:rC̝�~o���9ù�8���>�~�.7`��hF�}suiϽ�
F��X  � ��f%D

 R�L��`ր��+�79�B�"�/\/����X�Ge�o77�4�R��
�bc��0=���1ت��s���G��	;�e�� ������1��έ-F�g�m�:�15��l���w�=����C�=��n�༂-��VEDeԬy�ڊaGS��V=\�d$�>ăU�+���*M&�K� ��7I ��-�����:�Q�N� �ר�ɷ_����3+V@ �Z��/���*�8^V����QD��5���4�C@E��|�)ؚG�V�޿/�D/�|��\���Cxo�������Pqy�P�*-���Y8Oc��߱^�y�޾}�~��g��r�^�\�zȌ`�;����n�j�<�q�<�x�N"�^�yK�Q@�g����_���;G�(>yA�!D�����[�U�[4����G�7�~�$W���H6S�u�Z�:�}S���<egB��v����B%��{0�K�aJ5zXG�.��:���d�Ŗ=���.^y��5l�r���T,dܤ�1	5�y�K�#{�P�ba��?��|^?}��1ps7]�ӆ;S�!�LE�F���^�w���E|�	Ղ-(����h���͠$k�EƐB�T�ݙ: �:�VjX�����3�U�!�D�؀�F��9�h\	jͨ�^严��?���]ԧ�~)��hL�r�t`�A5'�O�eOA�Y��B8�Q��Uw�qF�>��ƾ�k�$}e�y���F�x����S��4�$�����˿D~�/����=�o��/X!��_~R�XO0��=)�A�9�ѣH��_a,����G�t�@����#����~�<#j79����k�z!iY�}�g��j���s�3��7i]�Pg���-#ﾽ\$����{�w��gP��}��=�t�'�n�p߽|q�����do�L;T�T���|nSޥo�@���/�)ez��Xs�o>SH�*E��㏧b�I<~�P�E�ǒr��	����0y�к�(H��`��H��`0���0� �
��$ �΁pm 1�B�H)�b��5�/!�Ol����!2�W~蔇����W���1
��'�N�g�D*/�!�ɐc��5�*m�6�GEQLp����Ř�$�lܑT,e��n�L	U#{*CN�ik����~�mn3����t�}��keN�i�嶒?(L,�Fx�_:ǭ�m�ܲ4��mdzQ!���cJ�'<�EԦw�j�H�� 8> v���'�F0NXO�q�OZ�'�V���jNVC�:J2ݻR��C#�Ya|nMsZ�˧�d(��\~�gu�׭/����V��§)\o���E�h�t�e�V�6���� �2�k'$S��+��Z����f������:D�X�LN�<w.�d!��YӤ��i���e���N"�}C�	R�.M3�<!�H�B?yp_��ì�g���Z���;�R�5,��YSd��� ڄ@*�Tf��_�)�#Bh�B��v���I�h -�`�BJ">�#<�������5S�O������kF�|8;#(�Ҁ�������ޱ��ws������4�T<�Xxc���*U1�������ma˫�����c��F���m��|��hZ�ϕۍF�(�U�:7GX�Q����qǻ�;9�jf���Ψ:�}��P�hc����9���=ژ!�W�,`�G�mt�D���Z�+�&k^��5�G���Q}�FI�К�(?��2U(Z�J1`��4#���;Ű�SD�a�wی�)պZ��X4Q�c��j,��╳hõ1�ek�B�*k-V˄�f)Z�Ö0�:�`.��7^�H)yu��E��R�,:�w�X��������7л��kDb-����{d�Lt����k����U'E��jq�#�"uP�ii\o,�1c:=#�u^p-���i;M�����Z:\�w���ȇ�2� {�|A�{��T0�DJZi����HrZA��z_���Xg�%����X2x�R�+��)S�8|0&bM �b������Bw�b	�j��l$�U��j���F��T�N��V5���h�fq�a'�Z<Ou���Ě
x����;yq��������a~&,|��O'���������Z����)<�p,xk[�.	~0�fQ��+�������~�IF�N	pP���5���*��
eZ`�[��MV�N.מ�]%�7k����:���u���Z2�P���tź�n�A��v}��
 �b�إ+�a�^7X�W�����?l��q:*�����v��oe�$��o���!�V{zC��i��zV�)+I����j������%qRnn�Qa�cJ֌��Gn?2��hs�v���[�
GH߸���﷼��-�g�I�A��?�j")�ju)_.dZ����_�3�d-�}iP �_�4j��q(��v-y(�{E75�[�Db�
�4}����[i�/�O0 �B������y��[j
N�$Ú�9*�o�MD�zWxA}ѽ���}��j��հC�%��9��n��� x�,��S~)�z�T��`6LY��g�CH3�֞Wo5�/y�I�3[V�<��b!%K Q
Pzy���#Y��kJ"C˵��s�(\��Y�j�@�أXa��?<p�'���˗�ʸ�������ǎ�xoov��P�ư'/XYF` FA��$��h��\����4����}���|p��͜�P��*�Mq��=`ΡQ�x왒#dC/E���%�w��G�!������a)gm~��>}1�r�E6���_J�X֤,������rfz�j��׺�
L�hb5��U{(�n�)bI#v�5Zn��9gMN�%�OU���4[ �,������)����)��j��V�A�	�^u���D��:l%��Ug�24s��4� r�E_1�H+=� }VٲjZ�D�����[w���9]g�����g��I���"Q�k�X�jZ<ƹ낦|�ŵ]r��>�hpa��1�h�;й����a2O	��G�|	}��+�0���G��ܝ_\�O�>Ѹ��d+��k���ȦF�if S٣m�O���z���	"dҰ�}�;0c��}w�.��A����<�İ�ߌx����ŀ����c��<�(�pə���do,�H���D�b�V+(��������k�Q�To�JSLWS��YS�V�)d��Ɨ҆�˷�5�u	�M�>���/���U��0b;(��|��J���� .L��n�:��=%�D������\X��_Ɖ����n��孛��k����������K~�>�'FDkF*B�&1�B9���Y����U�nԈSZ��J�[����y�h��l�5���Y�&���ư�6T�����..�BH)���8WO[��2Uk��Uu�إ�la0t�Տ��"It4xvuX^!?JV{D�E��5}���o�V
�������Z}�耺��c���.���=[ʀh��dL���1����{[Q5`�M���h�.�����f2a,	�	;}�Lz#a��6�c$��k��2��(E��[��5RGCN(&�E��T��c��»Ty�G��Q��':��$&m/����ܣ<��S󮚒T�1!�%��f��)2�ˬÙ`'��H�|o)o&�o �'y��x�r�N��B���D�t)%�k�Dw�!u_�٫ǗUJ&�bQYr�/�K�k�2�b�G�}�(�R�o%p"��!BD�6
h,e}�TU@��9�吮�Z�
TM���Vj�D�(�]�F(�g'�p���b����P^�����L)@:��E|<�
�Ϯۙ��y�/(ҼN�8���;:8r�f��)��I�W��EU�y���C5�Og��`�;����\���N�R��93�^W��ID���Ct1��$I����D94ާH�z٫����[��\u'	��|b�si�>.�n@
���w������K�}�}n{ic���鐁�~�H�vi�o=f�����7�g�j�\�D��ݹ��W]�o}�YV�dx����*�n�����Cm���w�b^�Zpq}��Á��*}���R�:����bԬ�#�Y���E�ES�wv�nog�i����%ٔ�<�l�=�����T}���qp���E��|ăH��KI_f�x̰#x)���L��*U���H]�Ư�{�ү�ϭ�g����ԗdGL���k�hMUN�P��L�T:�I��kP�9���jd��ʆ#�-���RSҖ��A4ͧ�s���".$�f�D�*K�)��0������y�C�kI�F2i`�Az�W�
�utx���8}P�����ܷU�'�X�d)�[|2��owY�r7^o��);5�H#���"����(\����u�ȿ��E. |��8I�s��Q֟�=3Ej�9�|/�PM�Kz���b����,4��h]���֕�`ulV���*l<9���7CzNo<ϥ�f�]d�?;�..�6*Tѓ%`<�o���� ;<N ��O���v��g{�hq�w������x��.���vN,(4!"˿���kgD !�0J"�wi&��Bk�>��N�`@oM
;��B+
�X�W.�_�6�%�%d�{������\U,��	�vqJ��ҊO�����5�C��$2;vȤ�yl��q����yJ��5�����	YA���\2��T���y�%e�ko���㔫blcz�s�����a]H�'����}J��.K��n�ؔ`F���[`��-1�j�Mַ�c0r�=Ԉ�Z{FJ`�m��4�ݚ�[<�H4r�7�Wҕ����Cp_zI���$�Y +n��]��L�����#
�45�i F��c^ha��ҰB.k$YM�� �r�m!�k:����m���Og�O��`DJ��Z=��We$�1�A9@�	H�d���nMRp�.>��v)0�g�Q��^��g!�,*0�9
t�D��x�2�t/�UY�L��)�4	�*���$�@k�,iYw�p-WJ1'H;[.w������"6����E|��0��UA�sIɄ���
��(x:;�н�T�	��!=�g����0�*Ar��>%�U�0���@N�k�d~],+C��c���.G�(��K�oS��0҄�������X��\>Q�2r��e�������$�4y��XN(ߪn&cѦ�'�uC��(~�S�{��|~�w�#�y���zM��ZyH��8VIu5�����g�2��ba-������TN&[�g̠ϾW�f�.T[%aP��@T��<���Y�IDzKg�������H���;�)kŀ�E��G�?E��,=�S�E7��C9�TxyM���F��w��k��a`PJ��%}|�`��g�.M�9�8RLך���!E��p/%!�؃�fK��7��t�zgm]�:���_=�vC�'"bʇN�!+:S�[���;בG]]���"����R�����}��۬V�h��oP�Q�8�Pˡ#KQ�8�YᔁQgN�Β/���x�}$r�U0�^�4��)N���OI�P�̍���(r������h�)_S6�F�pݣ5˯/�!��!ۉ�Lw��t�>S|��?�R�z�Sia��c8�C���wC�N��%'���<^g9��~������1��S��k��t����*�ċ� �H���t���������G(��~n�=oqq��v�����õ!D��_��eVo��D�q�h5YH����jc�7+>	(�M�W�[a�|��6d�L��F���=��nF�����l�X#�u�7oc�	?
�'m��=��a��eX�]W,�FM��W`�٦D5�Г-��.E &��X�GBL����`*3�s��Z�S?S�4l�Z�Zc�T��SI(�*������_�le#E���ؐ�9�-}F[�Uuˌ�ite��*���<�.+<A�h��KG���w������b�J�yI��¨xKx��0{�Ʉ���&Z�B �;�����D���OB��I�n��1�)�"xr��vC��*p�9p��y�B�'(�l�Ɣ������^�p��"���nV�K}�{�\�� �"n�s8�c��3N�$�D��� s >����G�ݻwf����?��(H������)���a��Ǐ���c��WREl�#�w��u?���Ʀׯ_��/ܿ��R.���e�S�<�-|DK�%�P��K��{JI$ʻ30���1��2Hx!l�Gm�0��;1��X��[k����B��ZOo#47��Oƽ�!=�UջCaa^�i:Z+���!He��.�P�ap�'�΄�:x��M\��b��t�u%�W�c)� �MݪS@3��4,3���:�V��-�\z-���n�1��$�T�oA��^e���jhxT��t��T�r�˴��4|cy�K*���o2�{|���-}�1��b�:��O�w}��}|���@[�hL��p��d���a��D��2}N�s��sM���oo�$�6�Ҿ�oon��3�x:OV�ң
����1��On��Q�l�����=#�	��j�%= ����3 �n?�������aT����Խ���ypt�.���{/V0�x� N�7��K��o��,����C}u�oJ�2�S�$f_�삅�U�J�Tl�NA:�97WW����i�9�?����2�:^{*T��9��!|��7W�4���󇿺������������I?>xR(���dlz������v�'�02_�>~�cu�Z����-�J�K��R����:��l����(�~v�� `���?�崃�[B�Exj�`��d��nE��9A��B��R��0��*�8��K���mKaM�~'��&q�Zy�My���c�1|����jܥO�v�t������v\*����w��P�`��{ov�a�5*��JZ��ahi�����K�l���\1ƈ���hzo��K,�**�����̨�����+eőRt}u)Q0��V?�(V��=��ک������*��3B�vF���g��׿���u���膐@�-d�F��0�d����'5��J;�r�0��BW|v�o��|�!�°s��x����>�}t���u�^���|��?��>��H!π
bf�b%��;w��<
���jpHM���]������w������B�[�7�����^i:D�S�"m�!��|��.���s��m���o�3�)�c�C�w�8����iߍ���ߍO�OA��-�/~�I�{�����+�9���fu�Rˎ/�,U��d b5�H+w��ne�/z!��Z%k�Ҕ\i�T�k�/�ƣ_Eu���T1]��_��b@�lf����;��܋��4b�!����i(����*���t>}���HP�U������^-խk�T}��p:FqVH*֍��t�����0�|6�[����<I�|��0ªXwr@�"d��Ɵ'��z�p���q_sk�}L��V��e��*Eܲ8�V��4Rƌ)M ��<0��i��Jk���n�f����/<�i��;�b��g�X;<>t?��i���ʕ�55ݩc�1^��ݍ�������Mc��nN�cڐ�����e�j`H2� <v�Fis�z!=�[J�>����v!N�<N���u�$�:Ww7���HXv;m�r-��QG��K=2���ϝ�}�!��*&�tY1Щ�����M�\IF��	���~�H�0��:HC+�IL)����Z�Qމ?b���ˏ�~z[�>��+"t]��W�Nv��HT6�t�R
��i��nİg�~o�����ǯ+L�B�� �dĩo/���_�;�X|�&6�z��H�2���@~��+������`&�"�$����=^��I>���F0q�0f����D�v�xG4;��4����1�o�9:I�>~��ڨhi:w�����%�]UAA��Z���']�����S�ԙ�LZ�p-�"��P�0Y�c���˨Q;�E�b���֝(�P����I�S�%�.��bbH���d*^O� ����*F�������0ҽ�
B9s�g@/�35�G�����g㷕G����?��C����_<�c�����c��s���G���=Z���#�a[J|o%8���ꙭ�UjA,
ʹ���c�CCznEŲ�N v[)^CŜ��R�q��Q�U�jD0�}Mq�P�ҚddY�@B���S�/-����m��>A����6���3I�k���Y��?�E�l���Fx[O�����]MVZ��c$�T9�/æi�"`���J�V4D[�ݠ��5+C"���A������#<����e��E0��d	\�F�sUP�V�T���|�)ܸ��%�5�iԻ��0�QtD��CZ�l��X8�v��-��,<a^������$>[|~�2@{�|�x�V�g�SYӵy�lK^�G[�}�o�/]N�^o�M��͚�Z�P>�5�m�Gpe�[݊�z�z�ç�uO����[tK
�(w��3 w��nqg��\D�P�q.橎���9��ʧ�qz��1�)���3������,<�38�xov��\�ֶ[�үI	���¨S�
��<�	8_pc����k���?��F3��2�\�B�m��yt_J��j���o0bz!6#w���� T��5�7��/��s��>�Sy��r��%{�B�~`��؏�Ε�W:��S0��i6�$�
�W��j�~�j��MQN��Hv50dc��L遤}YD�'aL�Mf�
�R�m�4v�����~ �{�{��7�	@���N�@�Ȍ�p�[A���Щ�8Gش]ϝ HM˃O�+Ty݅A0�ISx�� ?J�P�<<�L�m�"�$@���o�D(ԉL�r�S�sv�3�h0y �"�}����Vv��@�}ñ�L$4F�08M���h�+��R��%U��BS򞵛�ۛO,�7�Q������;y��bz�*gM�|ho��-m�/y���н�v�w��7^j˷|�q�Z�[E�4�����R)S��$�T���D74f<P!�4P���{Å�C#s$K�<H�"�$3�侓2� s���b��4�ʹ�]�+��מ�	U��Њf|���191d�H���F�a�z�l���+֋���1�^UC��Uh�]��73�e})?��&��
b�ʃ`X��{w۬h�XY$��o��;����	��P� �9D�^JUH|���������uR`��iJ�����~���O{��Z��i�e�&�a_}E䍕�����9�
k8�8�b��gn�bF��VΆ��iъ����P�bW#�oY1l��:�c��/F�T��W���p�l�B��ǧ4��ַ�߇7�[��jk�;�����y:k戴��
�*c���V@����J�b�̦���x}���WB,�W x����	c���7'b�&�3.��v	S`�P�e~;2��55A��kH?���ǽ`���L��:'^zb��}�;=�\4%Z��U��)`M��j�\6	��!���o��!��j�c��zRDߘ�j%\S�(�^V6�9f�7!�('�x�ȣ�*e,Z��w���Ҍ漭m��5G�a�؍�d[۪t�U��l�d�r���m�QHA��!X�c8q���M"��[*�sEģ��B��g!G$=<�O�����	��P)j�ըƶX0ȬE�|�� ��Q>��7.��IO��-x��F���d��p7SO�F��y�t�F��Y9��X�R�k�:�*l��R��QK��t�V�0|�)�� z��>����9p/ ��ʚg������8e��c,����B�������i/D��KQ�pﮓj=� {�>�U�xE�.�C�S��#���g�ZQ��{(��d����ۿG���hƏ�n�nf�G#]oK�\d�{�4zH��	V�� ���R�~�DK�8�=�a�~�,��FKpk�H�;��.9�̓H֦j[+�9��|$�s/�>k�KZ��,x�)��p�8�T�T\&(t9b�j������#��)[�����u�߂+��8Ů�L᪕ �6|�O����q*��h�{ ]Kg��f���
o��F�9+��K��F�11��d��7[$D�"h2�)����y��EQ���!��0f/s�����ux}{#cA��Q���e,��Rek`��@�8�?�Qk�CV>+���Tm������\V<lÌ����F��|�\���h��\�6┄fh,��u��l��x�0�Z��'���m����PW���sz�Z���u�@{V���v�v]8��PgSB"|�8�	T_je�Pa��P�*ǳ�=]���BI,���{�M�C3�72\/����W���v#���/���y�&�Uzp��t���l���;��-���>�F�ilC�V9ʏ�ۍw�\1��h�������A�*7�3�_���N�Z��S~k�vtS�ئ!C��`�rPa�Y�á�7��Zw�OC�L!��bx�.��3&��j:U���$�ܺص����ږȆ�L���ằ�'�/���h�9f!�j�ϾU��r�9uK濼�w��'��Ҩ������K�G�
V&���d�"g�ggF�%v��c�$h�ʄ9����/P&���!���1TZ5�t�L�y1���J�j�P��97̀��y`�1� �J, ��W,�JL�N@��_��,�����yav>�}d�םݙ�<K�~�ag/
��ؖ��^���ƾH�w�*ߕ�CJ�.S��յ��L=t�뮔��o��0ð�1��ݰu6���T�b�z�R�"Y�>�s��Z��chL�!
Z��lr�/ȁ���{���Sr5�?U���K�u��J��;�0�8"��[���	~d�Ы�=����O�-�QB^B>�ߔ@ގVV��L�}�HVe<��m_�]_�O�7�w!��7�q��V�R�h�>]�^�,�o@���ᵨf��vp���`!j�.ҸT�5G�O{�*�`�r]�/z=�-=�Pۼ#��:W) iCı[�qgZ:Kg�����# v�j%|�x3�;��#��is����4>E�[�+�1+�R�r�Q~��@��i:)lA�owG�
#F��:M$�SÚD�J�1ү(Dyy~�R!D� ��A
�����"��-�u��x�»����ý}XF��~���kPR�m���&�HZyƄ��_M}-�'�(!�׾�E�4 ���IJЙ�!6�>Ya@��K޻��wP���!/,��	�5X�,��7|OA�a�==fqz����Zܻ� $��WYdӢ+�sk���i������RH���b����PEޣ����g��L��^�p��T��'h@����L���T(����/_�80�}-���G�\��Fƶ�mdfR�^(1��~~��s�f�_EY8��_�z~W*��4��\�m����܆{����*$Eg�t'K���<�g:�R�o�V�������2%Ǯ
&�r�����R�B�y4}y7j�3��0�M�_)j�iH�8$�=:��618s���K�(lJ6�'�����O��O�i�y(6�y�4��3fF�]>Ƨ*?zi�]V~>r�Z6�J��p��Q��V4�0��<_|���6Z=����X�F�B��gt<�L6{���:"���E�~���1?#ʥ�Ls� aѯ�yO��TA�v�1X*_�!x6{�|uu�*Q������9V˯4<_R����|2�� �NJ1ެ� "��/����<=����(
����z��-���j;�`�(���b��9^��_��V��Ao�D�`L 6y�ehR���68wg�&�C�~�3�cɌ=����7䙎a�:�(犭1X�ٌ���&j�K�)�:��5�!�A�.WiO(q=:��R��ɔ�P?�O�7
^_���!�L���Z���y�_�o�`�z���a�WM�B��Pzr��?k�6KJ~M��>v��uZͶc�^k�S��ƐF���駶mc�x��F�i�����l�'^Q��%���+����4�[��K�]N+q:��oc��k��@|�"j6���"VJò>U� �>^�[����M]Jɔ������3&ErxY��[�7FUHd
��0��I3!��%ҕ��W���a�����3UhĈ5�{���9��V1���<4�"Y�8�g
�٠3/�O/���%��;0u�˘��(ܨG_�߱H��_�m��F^�BD,`0_$C�W�ȧ@�E>� �0��pv@�����P�F�c���$mۉ�j�Nh�]d�Ѭ�j24�[��f��� �����a)�̙nƈ_�qM��*Y�ƈZ�!fsX0@d	���5k/��]9;�z��\�ך�zBƜ+���{I)�@�t͂�W�)X�s�$YS���g���Q�f��;q"^��b�&���孤�Ul�����m Px�2f�X�OK�A�C,�X��gg��a�N��'�ڲ'�q�F$3���`�,,����Z�+��WE�*�UQ@�P�T�� �>�i�y�D߈�]�0��鱩p���hc����Y�])�؅֘vy�[�h���??uΊ��_�Ԅ�,�T�I.�����o�@I}�'�iO�<<����5�/m���%!y�>��{��]a�.�<��wV��,Li���m:�XB�si���$LB�GM	*1��jҐ�ׂN"��1�a}T��V���B%�ziThJ�0\�r<�X�y����vo_6��L���X��*^v�狽��/n��Q�c��YQ�#A���)�&sE�s�Z�V�Os��^[�( �fM�}>�?o:�~�y�271n��������#3�ٓ��B�9��`��3`��A9��;�r׉3�Gx�P�"�egZCpcp�9==��x�K����M!��=S�
<��ԁ`�[�O	XlkC�Ԍ-b��{������Ȝ�+q$�i�샀<C�8��Je���x P�j���+<�S0j�QF�tZ��k�><˲�k0R�9�R$Lu/��ҹV%�#����Su(���w�y��F�X�Iv��BֻEb�����'��8�ܗ�l����4֒�f*����"�F�f���=t�a^�M~�t"Tcfi����P�F��5RR����l#�����n�t�q��#݃�1�o�Q��L߇����-�D���m_��Wf�u\�-��CT��پ�V�Z��u��U�5oL���q����b�����\6��e�z!w��U�[�hP'�ۛ��=�吊��]�W�;��ʏբ.�B�+��%_��i��<ﳬdO�KdN#�3�(2t��i�YR�Dt�`�0R��`��&��~|�x:�����܁#NTv\(��ᓠ��z�_�նXYj��b8f"�4��a'�m
?K��r뗚�mix�SzM���������:����4�{������*n�������c�fD�,��4X�`R�P�QA��	:�����}Ȝu�p���V��N�畧Wkp�>B�r�۬<DV��M,B´��&]���P��8����JSn ��ɧEru��7_ݻe���;���%���e��DǬ^�!�#Bͱ��o���n.����O��g�Y�j��i�p��q���C+'>	,y���%`�W�+gz�1�GL�)�74�l���B�\[����O�ئ�|���:�����"��i��>���n<c`���ߛo5V���K��|������u����>>�R���Tr���U��rx3hH��������}�����*�Rt~(ܕ_��wn�����N<k�q.) �nY�*Wn>.GwJ4�E���8W�|6�UtA�g�ۼy]�g8�Z_@Y�>H�$�
!�����x:���i����0s������M�"�v%
�^:川��R�M�.��Z&]�\���t�@Z�c��2 �4�??to߼u;4`��f�t�	�s�挂�H������i�,��7o޸�������/L[B/vvE��!kG�<B��� I#��`�q3�����L�Lr���x�5��~����uI������x���WQ����so߾�W� ���W/y���E��+�^KTԚ�LS�;�G`��yXƹ��eXH�B�K����n� �~�V�	����	�蛠��>KGZ�Uׂ�y7k��&��"�+�>�=�.���FǓ��.�9����o��Os�����.�)3 ?�2��-��C;[~7
��C㳡�	��+l�*�ə��yb����a��S�ϙ�m80�������m,&�������8:��P�b��6�@泡7�6? LI��~��	�����vpX�k'��w�e�Ӧ
z���9{� ���x-V��f�Yc ��ޢX�3,:>^T���V�sw��w�1��������K�(�㧳O����]^]�?�y�:����4��O���J�z|�+�� ]f��bB'"c��"�$��d�����_��[�r���� ˉ���^�CzR��>�
վv�3�	� ��j.����K,��8��7ۛG���H�u��Gʠw�[W������0�.5F����{Y�϶�׋��:���,͉Q�m�B��E�Mt�4&`�F��P;ۥ��n�r�{�s��q��aP�<1<NR�G�3G�z�'��sA�:��תU����-j\V���r�������7�s��XWp���H����*U�N�?<��<�0?|�.��`�1¡W(���s��#�뙂�ȵ�{m�6�`u��\W�֕�Ǟ��=��F�$�^��}��dтC�F���v�ѩZ��C/�Z���ۤ���U���C0�?W�����4=�x�����0�<��q<�$�R��c�\£ax�,]~�|�a�q�Lg�:��#'�mIPY��~O���`i6���Np[ĸ���뎎�M"L"#M;����^��0�1���ޢ>t`|���*�2wbtb�s�.BЁq���*���Y�sd����{���^Q0�_^\����C�H���T��F��7�ƨ6�*H��\��e��	�k��H?�~��b4�8�FsIb�EA��ҷ�ܸ�y�H6��U4�z)O�R17�|q �؟˫Kg�XFmU�&S�E�$�>xQ>1#���2�R�S��4t�$� �����J�����*�����=����LB��!Er���#pu��_�8S�-ij�_y��2��g����z��&Mj[�iaf!%�
kJ����7�������mI~�i�"���z����kϕ�����Εks�1�������x2�4�ެ���V�g�7|��<G�H;ɗg���+��G�����Ҹ$�/Pur�O��n���䋈��x���u��~��k=.����&�)�c��Oܛo9�[� ))��̬��v��_���_e��t���Zr�]1�����V)"A���pW�˃h����z!��G\ ��ݿ�8<�t�,\\��ξ`�y�91{>}z	_%z4�;?�!�
�eм/_>�Y��;c��`ڱ�̘�M����>�Y�@	~���D�N��Cfs�&�L ��Jߋ�eo��$(BHu��5�=_�^ �s7���'����1wp�G�����q���\���ۮ��>z˞�I.Ǿ�3�痗p5b�PG;�,�H�N���?�:�\��~J���α��Й0�fT޵���ޱ]��aW�FԖD.�"�*�(L���>���b$v�Ї��c�� Δ)��8� �� ����7=�?߽�������*|��Ͷఔ����:V7P�2�b8q&��ݭ��tR� �îZA�mM���
��TI�^����A�|�&��H�l3���R��M���|Rr��F٪���yS��zN˰b=�@�D�:8p�X,�&��./s�v�J��z���cu̖�׊v�M(�r�'�>�vR�.7��L��f��T�fs�������oLt81僉�/���5��zu��15�D7���=�R*�i�Dal8mJtC?�0.o���w�` 0 ����6��{;�I��.d��pi��M�A���Y.���G�������<��m�΁YT�	@!z�hh�{����C����Ǽ��\�d��o��;���C���q0d 6���N+���d��IfI��}hAE`��Bכ�� OROH!"����KX��R;�]�YHW``˾# 
�}�N��NG�ι޽ R����F�(R�¼���������R;�����>w�ю?�t�Dw�,��N~���ϿumE��UxG/��� �>���%��Pb{�L�:�z�}�'�zw���2c88����W���)�R�=��НS�C�c�z8w�i�7-���~N{%yR�$�t�eZ�髫�����x!�)cx������m���8�K򒽇���[F�k���8�i�=sG�߫Ԙ�U�$��~wQ΍�Mt��8G����i���N�aF|{{nF���j���
��Mݞ���I��.�|^Fި��l%]&���<�L�^�pz�(�0�� '�;�;�B	��C`��?�"߁���]S
d�E�������E8�;�a� ��]߄3h �Cg^��u�F�@>��/�^0��w�C�w.`�vvAXfY�a����M��eS� ��G���cg�CWlߋs�(pF4��kI
��]�I�E�ŐXz8�v�~q���F俊�p���pz=M0h�`2 \�Wn�D�m!9���n���8(�q�����3u"L�r�[]�d��*�'�D�ܾ�_��`���R�6ۈ����;AS͎l{��5�X�_o5�8�#|5$	�YM"�W�$���Zc���ӽ89اpJ��W<����� �g�y��jϧ�擁���9�.�48ܟ��/۫�&�D:���ݗ��v���=�ٹ��m�/�+������V��"\s�m�����h�9�z�:���o��e�i�4��'��}���I#�����l��D�=�;�7�[���R���K�pM8�%r��E��E�Jp�K�טrX�30s.�!�����}xϑ�6�������#���|"gx`Ӿl�,v�(��RYv��C��lր�����exw��4nH�e``��[f �}@k�G�ڇ��������_/i� �����5�|pF�	3[2Ga�G$M���k��
�ދ�Т_�y�5�j}�����hז��99FpH�l��#`דdqI&i��FFY�j��m� �9#�P��jk#
�
м�лjb�%\>E����08hzu���C��u�}��$�4���v��>�O�AK�6*�b���T�'+���
&�H�c����0k�y������u+�|����yO��Sppʖ56g[p�Y����f��^�~�N���eu��!�cg����KE�f�\��I�S�����>(�ZwH�,�1C�9&V�j�zղ��F��4l�IƇ�#?��"�D����U��Ό���U������k��,S�o���ܔ��F3;�h8�,��Ɯ
�̔	4q�.�T���|F���7��ڷ��ѦŹ�Zɠ �5*`I��J'Z���!:�%��I�@��A�s61��N4q6D4�9!hՊ��A	�HL�H "��4b��D�4vb'B���@`Ġ�wc�ρ�����.(���l9�����Y������s.�����)t{��o�}Ha:���P�]�A�Gmi��b=N����X(��v�,}��<��[;\cv#8z~|�w�q�b�*��Ѐ���&;\ZH�Qf�`�ߏ �6�/O�����߈�nqh���C�Ie�J��n�'��̄�V�����-{٠95M���Q��ֈ#Iޒߛ.������T�;��J��J���Z��|#b9~�lg���dM��$���CH��{u���^f���������o�(KCݿs�	��j� >��<A���<��\��i��W
���u�ɜ�|�3sMW`_��>�X���
'Z��O<c�� �9x|�_���6������֤x�<Q�$���/�3�x�c]�|����a�<}N��߿��>�WWgD�n�n)�'9�{~
�m/_�yqOZ;gH�0��N��P �.�����=���͚`���ݑ_����̏���گA��E��4u�G���FT�W���?�����?���R�L+���P��(�}���?�`�@��33���K��~���1���A��� ��J�u�'��Ȃ�(��h/�?�N¼B�U˪��~v0& ��`��z`L٤���YXZ�5�E1IS'ؼ64d�� MC�����K�]|���)�iP�9��	;�r��|F[H�K����6��X��LAY(���5w���3�s�v�@��l��d-�FQ�u�x.����?��\�L�T���:���ǏN�t8QS�C�#��Z�.:�`3!G�:W�ټ�T �?PZU&S!u�d�"0O�����δ�LJ<.2@pB޵T�*���*U�/�#erc�}&8\�ɬ	�6+�SX�U:���q��	z���Y��1��S�i�4Iz��\ǎ���A}��f���<?�VPd)�Q>����H�����v� �)���H�)V�rs-���\Q �gt?��4�$
)N�?�)�H3ю�(2���;sdҸ!�eq�� \4�/��3C�ԛ�?k��0�k�AM���՘?��v3�-�S�Vg�,�!6��t#hɼ�I��y�<���d��x�����DGä���!K�2�����sǺcU[pFY�'I`P�m�@&r٨cg��I#.��Ɲ$\=;J�D cML����8�r[�ǧq?�>��e��ۈh���ק�{�}�w=�O:n����1�1�:%7�u_r���erD٘��4�ҥs���.��'���x�b��"ZbN��tL��)j��N���܉��Mj&3�5e������Ƙ(�(?R1͛��s���&�;�H���z%�~+S��%�X=�&v�sfs.A����L�Qfm��W��^�������6�ց��;��<�87"��X��f�2X�R���dx��k�퉾�=�J����
gm�&l��2���>S$Mu���hI��-�<����$I�jo%R�����Ux���H��� �AO����=�˗:4�;P�@��A?]wڸ�t�"Y�y��˘��j�w#��%����i������gDw9��CR/�ٽi<�y���g�_��5\�\]��@�<Ʋ����1�>ɏ��?��3i��13P�)0��|Ez�F!�
w�c ZRWF�~�u�}Ϫ�K�_��h�������OL�2�c���~!?�V���y����6�!H2����A{/`X犮�A#��嚙L�z/:�纃��葩�xl��p�;aV�$�h�F1��"Ԑ����A�w�R;�וF���ϴ�a�ޞ������������:�3�2�,4��_'�]��	%�F����XA�2��ɚ`�.��e�I���0��h���)_5;g�4�ê����BE43��ټ���M}K�9���g��gpL�y �ؾWj���CU������S��f���t��Hk��3��PI9�X�)X�G�O�k���P���s,�{>�9��B��'��j�*3X#=�Q$�Ҹ���3t��-y!ZE�,��ht�1q�p�2�J�}��#��l�<+&�����&��\�V�������!���*�1��k_�pt:��Ō�NH=G�Ll>N�9b�M����C�[fB��I`�fD�ڟ����g��,��̠Kb�]��_h���ͻ�5���c��6�@M6 \ūw3Vv�LR���[���n�9�$�ɵ��˙�]�9�
f����u�`� ��j�1�wJ�Β79�`n��d�|?}��~A����2��N",���e�D�Y�U��謩��
N�ؖ$=�F���&��	������9�����TV���R��~�+�����9��R#��m���)��ô��>>*�k̓��er��_�Z�~w $�����N6�N�p�&�1��<���eP���j,y�jo��&9hp6�������^�v�V]��0&�w�Jo��Rf�rz%b��1�����7���c0Y�
~�U,w탙>�]��֫�}��f�cx|*��
[١��8i�����lD�a2���Ţ-F�u������e���Wܾ��\4Z��M� .��	�k���÷�Rz�F��
��_�oݞL~.�F�qwv0zeӬ��k��A���}�Y/�C�'�!q4e�u�dJG���0F �^�/�fo&F=I�����q���f���,X�Rp(��Q3�2�u������o�s8�x^��iq�S=��ghh�������b �Lm/� 
��^�;]*1�ӿ{����|�Ë̩"K�d&��{I�4��A�c��HfI"h��6�휢kt��_{�څ9 �X�es��c�6��P���! )�/���`�&�`��:fN�Ś�޽�er�hk�3@��Ň���!���p�Q�[iU?!k��2�E��$ �A���~��pU�)W��>?N���5;R��8���á�6+=�z[k�?s������6ٳO8M��)L&yȽq4���M�SV���I2V�C��[Ge�ᨮ-8��S�������X�~�)#S������Y�)b��۟jm���i���\fF�w'���%��JZ���z��Q#i-c>(�����Q��<?֒�y�HxBe�>�&�l��l��	4�_�-`�|s}=��0G��#�\���I5;�ځ�X�@St��wu3拰� Ј娚AA|ѩ�5��`C/�SO4"Fh尖+�BD;J&P9ЌI�14ؘ9�����-�0�4�ĩ�FoD0a�
3�WҤ݈d0��X9HTK�@����~�#�_C��;��u����~�4��"�v���ĳ����o�ѥ)����A��y�j�_���Bf(�<�2U)W�BKu�3��*i���E�c�.�	�����B��;	�����8!n�o(�yZ�Ǝf�& ���{�����F�ORjZn���D��M�0���^t D��N6���S�HE�N��lQYz�PVh&�6*+6aW��!�#�s[uC�m�do����M�Ʊ�z5�����Ǡ�V��M&y�=��}����t�s�ܠxo�G�:Nxo�,�D�=����ij�T<L��c�;)� �\&O��P�'m�ɖ�8\�O+~�5���s=#�����,]�R��h;�����������U�D��&D1U�Я�/���Wt^�}��L�_JdJ2�re�����EYvUϠT(�k��;��]���g�򞩒X6����̪�H	̞���O͡'M����$��b���.<���_�ԗK��dQ��I�Âì��P"�m��+��<>=��۠�>��`&R�7C�eu�3����� �?~$������ӿ_໼� ��"�1#�.?|�@e�=�6պ%)�N��ۘ}�Q�nH�̙O�>I(��;�M՚"�/����Ζ��	h���>;?[�}sA��<�<��k'j����Y���*1G�4Y�e��w�{fi��3�g��R��%<&�Us�%�V�V�m�ʴ���;�`�m!��M���LP~,n��۝u��߹
��69��<�7��������T�ה�z�꽓��ߐ��m:^�B�	щ9R�&���kB:��ә�i���ST*��O��K�S,�Q�4^�G{��\��S��Z����I�Ԫ�<�R�������o;�	tg��oO�P�,1A׶.�@�h�%n�f���uӾ⺱֎�9�t|�LS�,@S�8!��#���}�$l�Utl^+��l
Eڷ=k�l���~��8���6$���{h�F�6"AV�$�0�6 �+�.�sL���ܣ�u㾠z�L�pc*KO1-��-	�8�L�t.tp}:>fsmhC0XH�(Y�+����y	�0��oEc��T���N�$$%M������[�ܑ�f�������fIZ����%�q�܁H�K%/ɫ�z��>�STLD
�e/�
6����;�A���`� �<Η�/d��3p��u0B:��w_��%��<O�(��I,R*��C`֞���5>�g�N^����j��:�e���txJ��:���~�?��W�N�(�ْ��!�����e��\�z�O"��� I׵�{fͨ�V>�{D�ss秌����\UuNGA�?�=�uҖ��!"8�B�;xld��<^����5��X��'���}�P��
�`���`�^�����]�Qn�й���Y�����i���Կ-�2�k�,�Wm�f�n�V�e�:���>u���M�!'V�"Q4'���������q��^V�+���t�����`�V��$�&�A+$Q�S3�N�V�j؞���@ ;pX�B�§ϗ�~��d��!�\X4'e>�Y�#�ל?2�8�������FΒ��g��ߊ_�KD�:[�?!b����O?�LZ:��������C5{����.���O���H�����L��FL�s�l�w�]`g��|��5�;�P�)�_~l������$9�:��Մ�`�]�S��M�޾d�q�(��'�ë��AT�9�����Ki[��P>x꾒d�Pf-db	��@�do�a��۶��(�F(d.ܽL�c�]�Qs{�O�lo �']G��磃�FC��Iݾ��'��3�k�W��R*�~��1|� 2S'�!�Fi眄�l����1P�|��[�it�+�]|���U��Q��ڇ�h�1�/&�9C/?��̗T����oe��ʴ!㨌��?zKx��������3}���L�gL�z�a1r3��7
��D�&�27(P������31��'�4�}b�@����'`�!���腦�F:�F�3�J�4�"V��r���I��(���^��'X[��A��T�ʔA�7�#%�PJtK��̝��}V���-�g���K��ѭ g6+#9n�P�2^�ڴ�YrYc�<�G�j��;�g�~V��[�+L�������_�l���;[�؁T������*�*����J+�i��`�·��S������ϋ��ý�F!�J�2`6iG��	�!�r�u"5��b_z�*s�ӑ�O3Pŝ,}�S=���z7g-NO�d��F�+@`+���A��<��{���8�a�C5����w���Vm:�2��6���h���fL��皩�k5��� �/�6�;�3ud��=сτ��j��5s6�<�Z��T��nS�mr���8�Q{M�}_s2�g %M��i�XY:<~��B��<* �{�Q��[�h��P!��yI�p�,� .�tx|چ�8�����yg`
."9�[l8*0��13T%`��ܰV����j���H�`���6İ�`���ގ4>d�4BDI\�|���͇ ��*��~����yp�-fv �����c8�?7m�~}}MH�:�$�#���;�ֹ��#�>0�3�"S	�|L��O�O>�Z�i�~�L� �3����^��f'Q6 l�`��Q�n\츲�p�3�v�}�ïK���|�b���/�.�,���>����������t���!қN�Y/���L >
6����%h�Y�kzպ�0R��,7�G�Y̷~B˜��ʽ0*���踕W�����������T͎�9q�T�i@ ��k��I!�ǲ��E9��.�|���G�Z�j�e���kpӧYd(�x����-���\h�63?�C�a��9w9��|�X�-FWr�����|�Q��F?O���8�ze�Iu�\D��#�9�sC��h�z֊��*�[/��%q��F�"�ˊ�'���H^FZ�*fI����q7l)p;�-�{��� ���I�v��f�!�sկ.D�>�����^����ś�ag��s:�M�RF
朙0D��{3M���0{:�$�%�W#��4�/�i����}�~C� U=�'3�P�^�j1�C�tX]�/����N�#������'-y>��eS�Wfl;q
B/���k�(����گ��o.<Я��,�����{��㯤��Yo-�E�0��-��G`���u���tu�#����Y��p�i|7�8h���N�?�8�x�q��kʠq�B�H78�t*�Ҫ�2p��ҏ�ڈ�߳��?6�.�1�x�\G�s�x-�t 񁦥�qG��z>`̩֜�@�|�ӵu��o��^�6	DR�>�Mv��\=cG���.��}9��c]_y�Z|�p֫J��`L]��K���C�m䍍�M!�Ɣ��T�9*{cfY���9�Fg.���}`������m�<�a���dz��\H���if�MsZlIs�1���휿�m���"-QqI�tKO)2���J����@�b��MV
�=0�ȗ�$�L�}F� h�HxuV�f�T �nRg����@t{{C�b6����%�f-Y�0W`Ҥ�kh����b'��q�a4����jb���2Y��6-.��J���!��Щ�׋�\0i���|� t+�9�(o����&��F^�yϦg��ŦO
�{�y�Y��^����̟���-�礑��L�N&�v�!�9���Q�f"����Zÿa�5��x������Wx�<���3$&�V"El#q�d�f-1̷NqC��f�Y����)9�
/d��.}֔4S�&iU���G
�S�ձ�Y�^�^��f�$b���̞Xf����Y:�+�Su��%N�c�9�X�綄�o�6�)�ч�}祬ٓ+�J��Ly<K��#����j�7Q4��,U��f�}EaBL��>k-����.S[;ӂ��$�`+������sJAq�l��|��_(��cGZ�-���ӯ�xp�]\|�#APg�Ah2 K�����B���~�:�Pf�nC-����4t{}|�#mڐ?[`�� B��t�d�������ӾAe5H�Q�)�X7-�A�t��e��ח����IHdp:f�y�60�	�"�9-�p�rws˾v�y�W ���LQ�+0cg!;��,4>|]�X�pu�	Ogd��\?����N�{�4�5�Rp�sav�qs����/�p��ѝk��6��k3���/\��~�~z~�����@ �3�qҽ�@����G���pq�7����8 /��{ݚ-bnoE�N��346?W�2}�4ʖ�g������fʛ성c�lh����f���L�c]��b^>�餻ˤ�˯#4
m7�s0�t���1D�\e�[�y:w��=�Zr %���9 ��k��Y�6�' �>]\���:&����C�ơQV&����S�Ne:�F��������^�T,��.U�����Y�Yku�zV�7$(::��1{j�]�_m�nɥE����L)�fGƈ��&�:Y�����]�
 �-�p�S�D!?)����XW9�>���9��"0KR�&_0�TA��KRi��5-/7��خC���^�S#?�\Ab'Y��f�v{)f\$	͍Q3��L����J��_l�O��شM�i�$�(DZ0D�4kG���N|!��aG�K
�0лu*1sH��_��v?|�^�_�iك�/�n��HM��M�FO�?��V�,�؄
��~?&F%L#�9(C�������ҟ �`D����İ��>�z�|6���.���,|�����{,>�p( �\������2��7�\���$չ�H�5���%��d�uH��bk��o��9�݉s\|vR�\�5*���m�ؕM�s��(�����e�Г�:�9��/�����g,�I�ڦy_�!������[i[��Et���Ho5��w��2��m��ٮR���F��w��y[ԡ�� @�<��@�䙷©�!y�=-��+��n1���ف+kmV��5v��p��H���:�W2�ƞ�����^���)�aK��a�IV$l�ٲt���f6b��,p�Z7v���� V��c�a.�� �3� [G�y-sL����1-'�8fj-Ek�~xv�E���]d� �����4��x~���$��9>0�F>!��X�;*����[;�z^n��4ǮCi�}��uc�ע����@��O�s�鞞9�9��/�~�ɳ'�Ï�a�\��QB�p��@*"|�[���eH��Fڮ���d�O���%ך;k���%l�i ;|��`�Z�:�@Ҝt�lcSΧuۧS���|N�u����&��+���0��i��t3���F�y������Q6��"Kpy�uZ۫7������Nɉu�%{WR�F�&����of^pwS5��!��Z?i����pK���e������Xs�,������lYʈ�D��ECȡΐ�Y9{]��u��uY��NJ� �g N�ՙSM���'��n^W�C����$�	���a5(H���M7:�uҗB�3
  �L�S�}��6��c�2۰\-��z��	1V����.@K�<�UF�^����a��)c���'�0���"X
a.��1^�����Ⴄ~������܂��ݞ��J�^�b��3���7���������Bi��A�w�b��3'2��yKZ@�;d���H!��4�M�pX"���|M�vg�1�`�:�3̥�#�K8x��/Ί����^#��5u�F��1��K*�UӉ��1�NӢn�|���"��8�읲w;�8���A�Di�H9�p?*��K]Υ$óm�l���y#D������Ⱦn\ m��I��Z=��<�C}�O��w���ϕ^Z�(�2�c�!3/���}���̄��YU� };)��|�I�9����`���.��j2I�<Ws"Eq?-�(�׵�RI��_��XcK�2�R�ߜ�l�*X��f��9\k�@�k;D����oT���v']?^�G_�������=�aא{�L���d�k*ٓDB���թ&^�e��YzE,K�"Q��	�|��I���7�L�����2������_G���L&Lx`ѳY �`�7Q�*j�	�^�_v���\]\^���(�g\��O�9���[.#�_@0s�yF��#�M<�H�:��e�S�g�
ژR�)L��d<e�Q&,�+��ՅN��N�A0V�����ے�P1x(�%���{`���N딓�/�H�da�~	�_�����d��X�(&Z�|���\�q�g��*�7#���� ǐ�$�A����gW�d�g�Ɣ׸AgT|^�I`��� 
���~���1p{�!5�:~)�TkD���`L�z�o�� ��D�$M^��*�E�O�M,�Q��1k]��%�W��T��ЄTºna�:��L�;sS��,����M���j)U��䲑hf��5� ?Ll�����s�Eۋ��CW���9���7'��%4�D�s�JrUΙB)�գ�;=���\�>�9&�������EE�ϧI������塩�QJ�~�Ҳ�.�8������V�P�]%ξ�&�7�^4��h�Hn��QCP����#�(��@uP�{��� P1�H�ĉ��ӹ(?��o�����6d��0��+v��Hä��V���|2�9M`M�.8�S��M�G��;�w��FZzC����3�j��s��T���S���w�1P�=9&�c���fG�<<<�o�70�no�(ʇ� f9!>s�!<><��~�-���G��0vs{CeA����L�
;����G�5��fL�����RW���F�I$L���k�� ޅ�����!�D_��m���K����(�����k!�yB�Ii�^u�D5fT���_�QGı;��z�̠�tC�ĥ+a�BKv��(���=9�*�w�,������=Kޔ0'2c��}G�Q����NM?�/��s�n���`9����)�7r���J�8W�4?!��P �8mP�eG�� {T������Y\��g&(ơ��f\i��~��ppB�&Ĉ!�H����~�_�Co1KB���j�L��n�B�f����Z�/�]ڹK�lCh<!�U_�?*���nYo��Fs�,h�\)/!�ry�սҞ��.��� �Y�a��.֘����D�k��J�J�c� `�ڄs$	'@[_^����A{'H[��O���b�x~&�;D9>F�X�V���.�qp�@7��%_]j�	���X��
�H��!l��o<�c�D=�l��PXtY{���	�M�/eXS��N�?����2"�=�[
z�t�(���qܬ�V?ӫcsjJ�uX��~
��$h�`�.��	�;
�i�e�Ք˯�dα�'��1�$�����[#��2���u1���2��!s��-��_����8�x���a��
�N�d[�G�����&��܆���᯿���
��
R�Nlݱ��D�s������w��eA̲��@�:�`�G��g�a���ɶ��C\��}���@���/:x��g���!D�pAŇ�=IA�A�
f���e�A��������#�_�u�}��8+��ǳ���>b�M�T�}�;L�����q���$i�\F���o��兆���!� �5���f��	���*_�O�B���A�|*�͒���ՆsTh�(�~�WI�<o_��Ơ&D�WN��.�bڐ�5�o��0UV0w==8�Ԏ�_o����103�=��L 'K��m�5��+��]�Gr����պ��!M�!`����vi�u�~�:qA�I:�� l� 6���&��|ȰO�h{�[s>���(JԆ��@�v��9XuK�_����}'*�}kɄjh+�gWg�<����q������7ZA1V�< ��ݽ#��0z��>ח������$��;��Ұ��}q�UF m ,�cP�=�9�GDgF&�31s��:H~AĮ�ۻ;6������-��������~�-���g����x���c�6)���V��2�d^�V,`z�~Gz���X��2 O�^�Q�*9;103�P7���f=�L���}��������Tu3���3�����b�$k� �B����]%t+kMijt�s
$���;���S��A �˞�3$�'����� ��I��D#��Iu3�A��Њ@�XnZ�����ose�а+�IS���Yq����C*�lk�5ZU�b�J�3��F�X���%\�J`��[�pN��	��4�6�����v���YL��u����p=3�
U��1j�Y�[e2�\�7C���9���x��|�r�CW�y�}3�ٽcf:��)�'3��_�\��k[�|c�z4�U���������=�7�ZB��-Xks�E��?�����&���AL��SXpq�ߋp;3���Xd��P0�VS���a��A����}�W4�^_G�s��GZ�@��6�Yx���mث��Q�c�������sr�'�������N�Z�S@���
и���������zG�8�է�'b� {lԤ����-1��@������BSDNQ>��/���p�+	��+��O 1�K���MO���r�����D=-;��!���q��>=���͘/�#C�����lh������Z^"+�ê�9�=ט�����[�t�p�>X�j&�q�D��0n��`���oZkCP)(΃e���K��p�4l�h����
/�.�$&�v����W(�-�$Դ�U5�H�(�4Ӯ��f/�dYG��2:�\�	<�Jܽ����]��� �N�.��Ç���ƍ�}�:<�A!I��6�x* �4�c���v��E�ua�d���ŖD��Rϕ��35��-w6_�fs���%/%KV��_���o<��`x�1i��$��	��e�*QԬ���|��~��+�gS���̔��.K�Ƥ�E��ğ�SdB�wOBr�X(5���\	B��e9�R��~�y����9�+��	��B��-(����IՎs�T��&dsđjN6j;y�'6ځ#_�o���wN��CA�'�0���
�C=��j<UN����"����Q��8`�\���3��`��l���\0V�$a>S���P?0)``Gѝ�i�ښd���P x�E�3#�͚�]�c,p�V쥭{�.��w���$b����1�*uA=��PK҂�6�1��̛͚�B�oD*}�����wY
8HNVG�p}w4�PG��ߝ0�nD�G'��1�������H��j�`:A��:t#��T�_^�/�l�F)��,���L�H���+C���H�\�������[�1i���N�kA¬���N?�vw[�ժ�C&��J
ݞ������K���;�|��Ҁ������K��*�mLh�{[ײd_Dq��68�����ê���4�B#yO���.M�_Dg�E3qv�B��:��8Γ�"����||Y����z�B!$��u���-T�������h��\(�2>+�3���!k��6�\*�"���J}����}ϐ��T�+.���L�=W�Ce��9�b��q�f[�?���h���g`�BkO��j���kL�-�YL��	(�
�L���~��.�$�ʝ\���x$M�W�4��5�^f��ZE���l�����N�.�y���:gg�puuF4�'�	�H��D�wP o��6ǉ�1H ��l�w����2F�L0Z(�&"n�>��)x E!I���E�
����윂8P ����F����CP��f��(�$ڬ�+���R�c���i2ݍDC��W�8t�����ߑe�c�ӫ�6�
���o�b#aB���
�:F٪��'�|�u��3!�y�)p�%V�P5Z�T���H`V�C�no�bAN���jS��au�"�p:1J����Ք�sʆ�3?���|
�Ǜ)��A3tQt�2��9������Ͽ�%<�`���^����`��$~#��=��<�9r8�V8�Do���F�S%�F!��8C��/%T��%�OY䤪��tM_3�Z,9=�MW�]����+��TiO8^�����uZa�,H���.}�{�����
�5*���b6����9�L�5,�y�[l%��S̏x��~l�+�C�4��J�;9O��ퟬ�Ǚ�&9|%�Ke@���T0�0e���K��Dx�:�$kݰ��\1�fPdi���:�ٓ���:jΥ����	&� �~wrd.Z4��Hh��t�l��YL@pϚ-� �sd.�@�ŽH~�6���5��/���)���ca�AӋ/�6Ayd���F:P��Y������(��0�0F�,��G�[��!�į���{r�(��m��I��E�P�s*�Sƀ2�(2�ꌄI� �ec4�W0p p��{�����Wg#�m%��!e�ϣ̗�0�:�4�/��Ak����=i%vd�	�W�1�؎���O����shX ���#�𘢭�ô`�t�����qG����Nc���9�5xB��r�h�,�=�~IA%���'�8��4*]���D���b�u.�/�cGo�_zȿ�b�@����kzX���1EsϜ_,�9�w�@��*x�/K�Izt��a���=�s����j��e�����9[R�vk>��Q)�9^���j���e���NB?���{cB����)+���)�C���zy��eƪ����/ʟ�6R����7���|Q��Ə�8�
rz	ŝͯq�����ΚM���?y �oT�^��|X੯J)���v��FA�7D�Uu�1՛p�l{�,Fz��(Q�+`
m6��7����L'�E�Y##���m��_��xOJ+r����	���d�i/;a����ԧ�^�͈�i�K���?$(�1Sg;�/���� 1����7&���#�!~�H�2D���@nS��@iW1mJ=�����M��6֛��	ʰsi[�I���/c��B�5�0zf�N�;Q��(L�8b���䛼X/��.mGвϯ�� �j8{��)}2���D�p���.z!c�������+ .j��E�Hz(���ȗ�E� ���GH/ ��M� 䂵{���^��7���Eu�����4���\�J@4�����S+5��5�9����H�-lװ
�4�t�j��C/|�e�������[r�U����[J�F�Os+�����!ҿ�ak��F�n]$�lRfN_�~S�����1j���M"����l[��
��Xך(e�Х�Vh�=�ɝ�����V�r�R���y�P'�
����b28�:3�'l����]��Y�#Z917�tI��/@�}y���lO�.��lC4P(O.����!��!|x��,4!�+N+-�<�x+C�#~�@_�8�yl�օ2�.��)�cA��a0�B/�H@��Ά�3���%���59�Q��A�Y�I�����m���B��̠��8�{�I&&��M%�lj(tv<�:�9��xUM"b�!��J�Os���:�����Jf]�c+�0:��Cz��˗�p�H4�H��]�\���;V�H`�<>�fϫD#S�q\ x��Au�B���L�*Z����W�uO�/�k��<o���7h]�E���-��I޿�b��}fȘ�%I�F�i��ɥ�SiJ>�ۛ��fiM{��q晫X�I�:4t�n���EYy�/J�N��5��YG��ͯ��=%"aJ���~Vl��M26s%;A��fZ
nRs
�g�X�w�qE��IU[��q��ώ�3)^LI�$�Cn[���/�i�ƭ|����/ed8zl>]� ��W�G�G�7֌��RA5I���FC�k��t$MT�b�iH�1�&C���F�<`x��`�S53�|����y�a&�.����D#rD�%��.�D����td�'����A^�\�i(	�o'�7�^�uCOk���:��_�O����CZ��5	2�T���뀞�y�vc�:��e�c���&���V+!�ƞ�r �Y��4h%�(���q35��G����}%���6��؋߹ּs3褽�q%���������_�5v�MR�{>YW)NĞ�i���QuQQA`��7�e��H����}���c���u�P/4	�����������ˍ�0+bS�>�d��
nz6�f
���o/`������9��a�X��Jf��94��K7+4�Ynz�D�=�OJ^��c(�B���4�C�
~=���%��M���s�����yt�+o����9R�P�� �p����λ�=�(]�Y���]��zH+$)J�����/_�b�n�]N�|v�1	J�0�V]'�k��dZ�:[��ꦲ�ƟsoB�b�%KW�]h ����vb���:�%�A�c��K���wf���٩s8rf
x�K�lq��&{�]T�ǌ�q�%Ud������*H��	f0P=KʁԬw�
�v���d_h�]��O� ��d�WIJ��2c��e��"�Y���� PM�p�V�&D��QF:;�Ė�5�v�^hǞ��@UȌ�a�5�Q0* ��zO@� ɟ��,�A�C(�*̢.����%iW�ܝ�A�M�K�t`n�$�De��ag���&5�"P*m;''��  ��������%�	�:�~���|��	�×�?������=����F偑�!.)|<�� �3�#͞�}j�Ȏ���Ђ�Ah���;�>�� M���T�ɬk��h��S��UX�s�3b줰�g�]�'����R��Z;Et�zCi��r���Z�J[���6���.��T%�`�ꠐR)�:�i��!}ɋ���kOIr8|����a�~na�8�H�pw�x7������"T���n�q*�<%��1��_��S��	�4��Tm� .�r���փ��4[��^����z�d�S��u���I�\QACU�^/sJ�'�����E�B'�`a�����e����e,j$u\�g-�O��^�üuL�.Jസ$�h�η�X�%�1LT�X���H�H��0vF,s�=���؁�C�:�+H@2�8���B��L���_����.��H�^�8j���H��fX�n��T@�ߌXd|OC��92܀�d�#ܷ��8�%�ހ~�����:*c��_�j�.9��v :HZ˄����L2�}�L���tq�w+}y��M*����L������.:�kn����p���mO���~������}���5|��,�7�s��p���B(z��4���эO�8ꆳwu����4��0r�IJXJ��0��Q�!���@����"TM�,\זĲ*)�4�K�l��!�i<�^t3�mEB:t��q�Jj.��M=�㜟ϔI_ �2��wY���5�=�r̀C�n֘��3W*���C�n´J>��u��i��2�Zej��@�շ)\���c�#��+�<i�M䦏b��>`�Ǳ+�q�3@T�s�8�Ǳ@�b!(&9-}��٤JHu���L�*K�l� ���d4g���~�hOj��I�<������j�;K�M��U�3x��rTf���.��R/N-��X�Z�[��R ��?�D�I�4�m�"T�s�,2��m�뉑�#�$A�#&0�^��oE����"���0A2����B0�"s9��
�;(�?`-�x� (�|8���Hwֳ0��K�D�ڊ6�JN�Ƌ"zt=�k���~�z"����H���ِC�'�&��GbP�Y4� ��L���~���"J��	f�?�0�4���!f�Ã-�!I�y�'��d�<oԌ�lّw'��غf�bI��<�U͖���i�x���,S��
��%��2���ސm[xT҃CL(π��5ꗁ�ϳ��0�ܷ1���N��$�۪kf�Z07�v�J�*�'Ek�l�6u��	�P�4��!�4�\�e�b�D�j�2���� a,R��K���Hkh���g�@t@�q��(}�±�5Tj�k��>T���z���~W���������^sA�R�:�ϸ�'P�/1��m~�NpL�<hԿFgl߷Q��嵈�M����P~p�GՄ�sL��`�_�F(�:`����l���EBl�4k̷��t.A���Izs�����}T���O�/����噝��Ξ_<�I�� ��<��)���{l���Q:}�A����0v4B$�!	Y�J�B�w3�H3h�F�ǌ�e'A����|�ξq�9x�i6[��^c'j9��M#\p]7}���p�x��V6YHd#>v������◇���8���GR5'��� l�s��~x���p�:o��<�p�nb[u/��y	I�Ij�Lv8t�����6�13b�ZP�ze3)W7_פ���qȇ7#E3���wi�uɤ�W:��;��	 @��F��ѨK,��I�ÙN�?�j�}�F(Y��uM�{����C�ibk����ܩۭ���xY>.<ax{�e8��W<�,��>5�zs�GS��]Y�u(U����>�I��tfD��+���&�*E�ɗU���3�A�|��r�N�5(|(�S%ij���;����$cd��Q-̹A�I�@��d0f�������=EǢ�t~q�$
H� |vb���Vl�$�7E����:Ѿ��	G@��YB���;?}�H�#W��p~���2c�0���f�<����*�W�	�e5n�/W�8��"~0#m!?�Ss�̦%�����`�]P�*t��4l.�`&�{�|�i9�32O�م{gb>�_�#�E}��ݻw$ż���>���#BЎ�u#���j�R���|������s�̝��k���8b��������Y���N�)���Ǿ�.0�З�"s+�Cuى9�9�N`|u�!�V$�(��[�h���iWt�ֳ����L�0_r���L�C��<��[����>vQW8��H�'�����>c�C�/�v�������b���e���{�z��jZ/9c�|���R%�{F�)�:�}>+����!����3�$״�̑�80C���D��&G�ۿ*4&���BSS>{���![�Iv��"&ue-w7�;����ok���1��T5x���g�m3w5!�j�f�������zݧ�L���k4ZQy�ێ�#=ɡ�����`�������P[.Ȅ�M�W��G�&���ߒ;�͎�O����܇�h�9�_�ێˋ3\ ����W҄}|~�_��ׯDA���#�/ԧ�1�(��2b�(2f���o�^4e1�H�L��X��LN�ӂ �鎘8��ْ��m�#Kb��S(�����ꚃ�z�ѳ���BP�oe�)!�}�tj��>�~������oUŖ>���װ�����#�t�u�v�r��_����=ݕʶ�!sT�^0������p�N�*�V)#걚h�Y+	H���n5C�z�c�$�ɸ8�E�=$����W�kJ�rZD��03P'�*�8��1r�e�2 �RU�'����0��QZ�NHcU��_�DJ��n�̊NT-)�ݡl��-�C]��G�q��P�z)f�J��T��Z�{�F'���y����
,,�P֣�7���;[����XP�3���_�a��]�i~�f�Fy��ƥ9Efb������I���Ś��"a ɼ&E=ۨC��j�D�KT��L�H����H�cTKB��o��;!e��]$�f �;-)�CzD�8;	��!�4�3�6�rM-�DM[�_8�C�񔉱��{��.�ڍjn�ڑ�>�&��ZO�T��l��w�[�4ݘI�p�ܧH&�V|�%��vQrj3 U���o	����:��Q��������	$ H`���r��f�X#	��z{�EGcv��+G�Bw���=1K0�~��G���3�L��}��>|x�A�`>~����IK
�>�!��uA�m0�[���0㧓�F��$��y���ͦff�&&h�cgg�0����@^l9���2��p�yЅ=�B�c��b%�t�����[�F'{�b�#��c�`���pC�)�B����?ܖ6�P�~��?v�x�|��|m�-�����a6�iiy9Y����xr�����ץ�Jf^���(�ﰺ�A���A�|J�s�r]����e-��:�aC�:��o;|Rպğ'4q�V�Y��)QGvj@���#�:�RKKs-�C[��E;,f3�r?��t�G����_9�e[����`�yӤ�uO�r��mK��b�LCv)��2A�51��ܮ�ơ�W.�t�ޚ��4��*�^n�`0J���H0��}|�!�ES��K�:2�j)&�+2�%i�j4/��Շ�s�� MV8QÈʆ���>����^B��)<�܇�Ӟ� ���Bc����� Spqh��Q��f�BB�wv���"���J�l�$bm%��ŚE[��h����I��$2����!ݙ���� 
%��E�?;�ST-o7�Q\�$7�ew�}1c��U�8�#�����Sf�ጓ4��IkE��; ,��<�,���~��k�j�('S�h�B�������A�%D��M�N*g�b��]v< ^ҡE��k�}�����yLE�MV���Rƃ/�F�����K{(Yxy��Q��rZ�Lj<�8�=���2��uC VH}�]Z|*�W,���fM@4��'o,��d�Ԉ��G(HTFb�9�}�J��՘���2���be#BI���l*�VW`K�ZiC0���r�J�������Q���W��o�Ml���\��� �����w-�:SMd�*�k����p�]�q�r��*����	�V((-Z���3뻖?������}b����A��Ĕ�``�o!���}!nU���Y�~ Ǆ2+4�s���?K;b�P���L�����;�4���7i��{'�)��XO�_^�a�JaI��XnZ��9h��}r����y/hR�_����P$\ ��$�f�$H�����T؊�\���E�$"M�X酱��]#-6M���+h�Sg�xֶa�1s��C�Ͼ	Ј�84V�r�|��A��9,)k����0������h��$}<�Oh�b�񇹒D#CZ��ձ�6~���� �����믿�T���m�駟»������ᑞ}���ѿvT�����{Q	_��ٳ)4�^��I�vM(_��)Ei�f�1S�.0G���Ǘ'�c_l(�� ���t/k al��<O�@����p�or���G۬���ļ�Otn=��C�X��܌�c�f_�Ǣ���lWE�t��=�5�R���fLwW�V�
f��E+����?�Ut�EqF���lQS�y�(k��o���E�	�:�1��)�}�6齖��,�h�%E��m��pe��B&��}��TK��$��İS3�?ZA������C!�1r3���G�)�����>��E!�g�и���������AKX�����/.HBdF�h���Yۍ���M)���_���G����ZJ:�B�,碔�u�Z7����a"M���2���|�p�nv�o&�笙K�� P.;��"G��׳۰@�t�|�90��G�B�u�^��������+B�����_6�V��&�I�1�f�����
�Q�6�4p�j�@���u��τ;i�0����`����]�G��Az�}h1�a�M�	c�d�1��a�<��<�.�Z�dr�[o��.![24�G�|�Sp0M�S.;���waK�i�OPkN]���Ƕ����c�G^��Yw#IF��8��n��qŢ]�]nsMq���|*t�1�T��v�7G�g��)�>i�g��΃˜�H�y��^��s��%�Tb�0���/���Yx,��U�:�f����J|��L��� -�$��/)m��@�V�L���EV�x�ө�[�H�A��ɒ���J�?��{.�țu����|�ı�Tԧ]ʜG���O�t�d�Lޱ"�����ԕum�]_��{~"����2C��G��ڍi����Ő�)�V1*�@'_ߊ��}���sH�al��V>����U��!I�D��[�+Mx/sBzzꆙ�U���DG>�q���:;݂�MTl�Q�4@�{�r��9�S!�8:K���/��t��iBΟ�縷>[��%�-��t��Q���	C50�G3�{P�F8T0S����Gg"=;r� v�A���@G�s�X~D��$;�ޚ� 0�h�w��;C���fmQA����j��/�0��4�݆P#_����~��1knnn� ސ`~���̩qZLΤ�}3e�����Q.4r �aF�����&����T��G�c����8�ܒ(j ��3�e�s������)6i�`Fq�~��D�n���9\{��j��ޯ���A���b���hn&eY���t����R�0G7���s�`����+��s_��	���!ۯ���L��(���nfϳD?�-�WYPӋ�Μ���N�A��>+ty�h'Wx��*5���lWv��}/c���묦b:����ؘ�-<�[��_)L�v�q��Y��s8G�R5S�����:Z��-�9�g���^���xJk
�/ ����s6��S��O�u���_�y\���$��̩h��U��\�Q�o{sK�=�w�V�t:6���Q�k��`�spT�� D��
q�d��/��*v� A ���eX����[R��d�u6{��=Sdj8I~ݾ�4͑1�?��#Ί����6��s0kʂ���n\�M�S��X C�65*����� �(�Ήǲ�v@�-iX���gט:�,�+���ɯ�2ttt"����O~����)dM���Z�2��|V@��飤���oP�st�_����U��6o"�<P&�1lr��0�dp�s]����^iޏR�4U�dF  �u����Bq�	֬/�	�ie�i荋e�p~ER
N���R�uzR��C�G���~v$��Y}�})�/mo��Q5�3�2�<q�yKiZ�v�R���i��3a����*�TN����,^��t�b�͕������󕊶M��!���V]3�}Y���"��ǚ���.c�1a˞�w��'�)4���_s�)b&}
�q�]�J��9N�0�\-�zhT e���w
��m�m6]�~η"�I$����,R�l�#��-��XII*��{��n�o`-��<�	�A�8�j��`���.{b��u���������H�zb�q!F3�";~�=c�S������Tq�-�}��Q���:p�<#i?!?����)l���q�&�hꩌ��{
A,0>c�փ��4���ӎ4��i?���I�'{1K,e33Ў��˫���ÇpssMfS��}�8���31`H%��db�@=�1��%���A@m��������a�~?�������#�!�����31���%GF#�ȾsV�ؚ�73��mE��ȇ�@����X��	��R�0�NƟ'@Tl���h�q���+{\N�8��ϙ�{&����y�od�Xm�Lbk�����C4é�4)��H�Eʝ죿�t���xB�%!d=��f6G�|�0�E��<��mr���l��lBY�BF�p��}���5��2;G'L{=�+%�amS��YN�����أ�7��|ݫ<b6G�L<J=���N�l~�¤�Ƭ`�T�9�C��vo:�e��j�1r�R�Tz�d��}L[-M�sPq���d7��)h~��]�����[���=�����:�t�T�S�4މ�Z0�̈Ʉ#�E�Z��@/��h���b�M77������2�8�!,�#g���v<C��$(P&��Q{u����0�"�w��A��HB���C0������v�#�<�@c:�%�:c�g����f�*ik ��H��cs� e�~�/+��cm�A��Z	]��tXl��i�!���[Io��%�r-�j%�j����(fr*�u�Smz���v]��R%���[;��Y8�洫�Z�;X��ӝߵ-5���e����6�+p�8�������	Xvj�kl�U]L�x�3����)�msW�]�j���!���HVR��fF�{�� �]N9�����N��W
��:��|�奫�b�O�w��&k�;��Ȝ=�2�x���pt%�������C?�U��L�Ϳ����q��N��c6���I%Y�_�2ˏ��T�/4�;��O	���H4W��䁭�A�c����r�į�(���E�@��J��z��?r�c	?�s�h	̓����CL�A%x,A��!͝���0�?88�p�0��n	�qD���:�FA}���0�0��2\���1̆=�����R�����̡���A���A��eڤ�5~�	7��͒$yC�r�d�_`Qu/���#쇽a�!�myP�w�e��� �H��]����̓�ۛp{{Gm���u�?��#���o���{�n�1FL�����(BV�~�V93+�|�Dm�8�����M��1���Z?��a:i������uK�|�U4�.�CM���1C5JM��d&7�t��1�PJ���<q-;Vw�T1��ٸZ�8���F�,���O}35����\E=�g>�4��b���r�g<��VW�A�g�U��'\���&qyBzr�s�Cʰh^Q��aq�6�*�3�0I�d�d��i��zåQ�k{��,�J�Lƞ�1�RFC1� �lR(�;��� ��~g�E$�S|ܺ�T7۵-ӈw<�JF폎��=O�nx#<�e��F�����Ժ�N��G�\�:r2;e��j�=�W��֞�Qد��/�^��(A�s��3��WV�`김������l5��E�k;�x�j���*5J�
'��5E�}$:�Tc�5�w��4w��C�D��9��gVlM��&�Ġ�C���/�W@��mː�0�e�"V!�F�2g�2�������m��s�$a�55e޺O�:�<dzT�{홙Jie�؎��>@��c��9��f�&�nS�V�#�q��J��^�=KֵE���i#����`��*�ŇC��x��i@�%v{�f�V��h�>*&e��Oyb�LR7�!;��Yg��feb�~��9�b�?H�*j�] �~���ظ|O�w��kj:�͖�网�& i^��CR��գ�v�ڝ�ı/������*˹�+6�EU?L�)'%z�'��i}��J+���ծs6�����|%���)HRg��������N���QC��CD�B���ʱV���'0�1 ��S���́h{�:��E� 5�^�����R��KC;#��N|��̝k����=����ȉ�$n��;��L-��&��oϑ���ݻw��{���	///���4\Hf,���:�W�Tv���z0㉵P4��űS������� g���HM{�4�-��/ ����m�ɰ�u}vKa��.����BL��~��خ{jk�@����o�8�Wc����P�`p�Q�32E��~;����-�L�G0�����c�I�	�Y��`�簰�0w���Ű��2�~ds�"^B��o��Im� Tlg\�w�ó�Jo�'�G�"���?�8�٬|�ciz��_�M+k��85���gg�O��J3䟦FG�5O	?��s�r�="g��<�l��\Ӥ�3�V���	 	!;p����홏�eL�i�[uDț�\7o��k��H�f�g�����ji�T�M�ّ>�z8�ʚt���2���q]Tx4L�q�5�j��̰bP\�GS����ћ��z4s*�L�+��`�ґ�
��t��gL��x��$�	���6/XC���]��aq����0U�qz��,��o��nC�����(��l��7��{%��y��q�:�oh�cl�O��֮�������D{w�&�V�H���vX��e������-����@�-��`z�Ly��o]�0��N3�|Ϥ�q~�LV_^�-�	oy�-�P���G
6��I�#9�7�t8�������:�[�Mz�e���(#3���cH�'�>��r���^�C��tmGR�^T�)��'ٗ�yf@�C���7ҋ�֖�D�?�T��K�ܩ��}<'P��<�R��)�x���ՠGy@L	��y�s��\�������T�T�$�&u�1z;h���rC����!�Ku��q�-�Lo6���k��6b���F�d�6K;{M sV��R�tza!gY3q����|��ס�v[�݇Kf�>T1j��W����)HØ���@�� (`"'���\����P�rߑU�0�=5���X����G�k���� ���U��>š��8�_bw��ri�z�n��H0�D���#���3`����`����	�Ƌ�G�b&�.����:q)��:yzz
��?�V�!�B����LL%H��t)s���i�dN��*fQ��R�.Ω_��M�k2F�D{���z8Ć3�gn/@�|0,��C�����FX���Թ���c�}}�'��/��Z40�B�h_[j+�U��A�����#�������ٻۻp{s����b�u"tٳ�td0Z���L����m�>�H2l�c&ݖ�P`��Cѱ��"����V�����9cu�tl��e��J�����׽;��j��4)��Q��;�4�w�M����j����	r�M~��\����h�/��ry��)5H<�n�`ʨ�{(K�����Or���y�?y�T3�t��7{>Q<h��Ֆ��jƦo��,��U.��֛�McFq�[TS�Vq?����ْ�$h�8���äS8�}`5��k�a��7�P��^��3��g������w\MC4�#fF�'��XM�YuGZ'�>�Ijخ�t�~�l���y0b,�Xc���$��݂͚)��v�]���	pڬ�v��F�>d��
��_:��g�D3ooo�7��H� � wc�#���9�|V<`�MQ�Ʋ�m���h��@#Q�P������>��u�����̫A�������5�w#��m��}PLHc4|�W�8�T_q�Q�H&Qq~+��,z�<��e��$L3[UH7�Fq�i�mp�m<Q�̋��a����z��|�|ǫ�~4�_�k'm�����c��Q���E}&��8w����,�-1w�H};qJ�y�cD�Pt��<�>�?QJa�s���)�J�V
��Z>�k�,�JeC�\��U�kbz�?�o���4��y�&����S��$ ǈT�F���F����`ʧ��9a<��8��JʸiW�z�ʕ2m���6�9�*J��I�ܯۃ���՞s��g��i,�	^
��)dM�r80���1I�t���>���Z��!�¦����H���,A�ۡΒyD���o2b� �`�K�*R)�/W�3R�FF�hQ4��aB��^���C{��� gKa�y�u��������:4gp��M��CR��o!b�Eg�j��d	̡^�A��ϴ�>�����'�����5H��g�rA�����!\^^�����!U�/�޽#�.��8�ڑ� {D��{�`�t��8�>d�i���UՄi#T�'��+Q�fӿ����_~�i���v�~����#}��I|!�
T�����*�\]ӳ�c_����O4��V0}����;�#�)c'B-~Kt��h���N}��u��^=�}�&f���T �ƶ�B
0b4�����uI:,����
l��a�HRG�ǘ��&���/۵�:��>�=X�G^2t\JM�D��N����GSwO�E�����̛�M3�Bq B#T|r�
h���Ij$�!k�(	�SW
^�X��������5��e������ �.8ԛ��:�J��+H���5َ�wp��·^�P!�Lv��[ج��ѻ��N�E@��.�������1�Ǥ�b	�E�t9�L�����F����NϘ�`�l��?y��g���(��I�W�K8��>�^���51��_X�A��5�rl!P�0���EgT�	�ԈR�1E�E��6����/�v���/����h!E�|~_?}_>�d3pb2	�Q?���C!�;x�^�Jcdf�V3=9Yf�m5�B� ���4�g��-��m%�o�%S4
�u�d^&��y�B��瓛7
��G�l��r��Ib�S�oV�/�<� A�0W,������Խi��ȑ-��R�]���r$ӛgzf2��"�$3jH�t�]k�@(�q�� YU�Iμ��U�������q3Ŋ��Xx�`�����8���a�u��QCw�Z�,��l��F���+�k�7����:y���qG�e��<��9%:lJ��30�ڹ���>��1��  ��IDATSc�����HI^���q��s��k	>�>
��Gsg��Fi��a(�Y��9��%����BӮY��i�jn�������p�C�sLO/���Q��s
�����,���O�z�e�Ny���~t/�uV�u �/��������s�]����A1�Fk|:�M�9���x���i�P]߫�1�C�̵���r�|:";C�tV����I�':��~�ˈA�W=���J�=e�*K��ֶٽ60��,�9��aC�h���2FXcD6�쮈���6��C�����y�zp���<���!8��m��گ����|�*?|"��7oI��&c�:���k�HUb�� �}�� Zώ�T6����HF1��_��t{ 	����H���$�%��޽�g$�`k��`TU2��KF�X������7X7�c�?�A�:Xzxz�d�dВ�?�r���`��+s�����[���k�h�
�G��ݖ�]'�5t��v�6�9K��X�6���E0�@�Zמ���(�=���3 ������N�i2�;���IrPE���v�4�mg��Ez�}L�@�5�FK#����ڧ#��h�U�~d�U�f%�l�!�f�De�ȇ��Ql��������,1�qJ���"�xIƅ�?��A<9h�V�sqT]j�9|��μ�7#b�����`&�'�v+�Y��ؐ9q������p��=Ӛ,:ۆ���;?g5��x4f��9�z#��p��]�|�7s[��4��3.�rT�$\'֏�x���h�K�G�#�Jǰ�ڿ'�`|��*�-o�m̥��?���CȔv��|&�M��9�p9y�V��lU���Im����p����Jҝ���%�A"�>l{�~tQ&H�,�WL�����o�0�fwt��cWѿ����5�����j%N�O;ko/�;,�:��FKD%pf�WѮ��S�D� Y��p\a�l7�����A/jS���؏�x/�M�ɝǚ,��.�݅����(��d�v�BR��N��wwD��:��sR��u<��9i�DE�S��z���hH�,H������q�m��)����ς;s�*s ����"����ML��Q��ޗ��C׾�²�s}|�"9a�����g�X)��}���'�d@�N	��t�L��0�U���Z��R��#�tl�}����os1v�IP]�m�9FG����dHꘗĳ^��}�~��pz.`�
Ց ��zF�� G���WJj4��k���3V��J�#�2?�^�U�uj�&�Ƿ��+�'#��Ma���v���0/(�Xˮg.F�3�6��Z˒��0�{����:��b&��O�~�,���̧P �u���R'R���:�3{�w1}��ߛ\s6uG��x�YsslC>�UA����ȉ�7�PbF{{o'Fvd|mF
�0УU���͑�bYoN38�נּ�H�9˔�H����]��k ��E��HB��t�-� �u�0���1���Y��P+A�֟;b����3�3$P薮Ă86�-���z�����o�r��1�?"f�`Χ�_���P�wo���w:�γ���]�ᅿ�qA��k0&�lL�^)�!��,�j����E�����$rDg,v�X��c�{E�A����_�|� 6�8��i���5� m�<�K[�?�pt�K�y��{w/�x=� 0V��y�+�gD4��
3�K����W�$#���t��mLc�Q����H�C`$��y�mF2���VB�F�h]��� ������'dP�A���!�
���+�e72}NF���g����<��2}g��� ��|��m\(�H�} ]��;tۃ9������0�:mg��h&zcn�8y���q��lq��Z�����X�sɘ�[�3����k2�ن2���G�n���ٳ���f�����ջ'tǩ-��v�g8�<L�y������8�%���*'��:��I��X�<G��d��-=���~�sL�Զk����k-5^�qf��T,n��9���m3^a
UB��
r$������������^��w�q�[�u<��AM�6�@�
yrv0�a��V��+5E�B�B<�?t��$%�I]__0������k��\��=�R��AO �ܸ=������p��d��Q��P�ݲJ:w��BQ�M�j5�Qm3���c�k�ɇ�{�� �^-��yJ��c�E����E��.�C��c�_�'茇H�L�Z.�D\�]L:���ͣ|��%����j��Py?�K՚S�d6 �K�R{��7y>�.u�.��V50�n��g�nM��-�5�U�-��XCQ|�;q����2S�[w��y���P��M��[q\'Q���cE���p�֓{`Q]s~�"��!l�2n`��;���)0��+g�UA9<N��On�Ӊl?�Ȩ?��&;u�>�����N��<3�;����YB=�e4�J0�X�Y6!]+�lXٵ�L�jއ��R�oF�����g:����]���p�3�ы�;���q��7�U[	����˟���)���ܪ7��b���&>C�E��ZO��ajE���u�/�=E�����h���|�q&Nۑ�f�_��U0�>�D�18�uΒ�^��w��B�Zn�C'��{!,�[;��b���sA������nOg�$�=*��~�!�QK{��#��h%�������)gˡі�o�ݘ�h��h��EKmA\|v�s��/��޿�w7o����zK������gK�p���L���7~�^�8�+G�(A����{f���ɀނa�F+��� w�.neMl����d{��5#���O��A7*A��^9pt����.J)16Eʪ��b�:��}��J��x�g�Ga�7��z�9p��.X@�t��X=�VPS|���m{	��~������sVK%C�O���~y~� �ř�0?<����!��f��xG4ρA���K��0~�6
 �Z��
���v�yU�b�Һ��E�K�Հ��X,K�Z�2MvTr+��Oʁ�;u���~.�*}/Rdj�k�^u/�~?f�����1z�la��\.b^������C[s���ө����4rav��8�,R�@�=�8�%�|>�}�磝;����w� �����%L���;�2#�wt����e޻]^|�l��RƷp�b���M��u��;f.�sd��k�{�J���\L�h�/�`Cc��`�2��L�ֵ�y��	Ġ��eV�y
�D�(3f	n�ɲ=��!��U��2t��͍\߼Izm��� 4E��=������WIW^�L r֐��Ʊ�D%��R~�y��f�z�v�2(J��?���ߔ��C�����GXv�Z�~@�ʏ���قA-˨�zF=�^i�V(ׂ�½t�u�u�@[�,p��Vf�� ZG	��9΃N�6A�d�4�4i�7�~�6m�E'�}����|s�z�c�����}"�l�d^<�'k2��¤��E�UB6��8�J�����w}Z1g;�:�-<X�����&Gz�D�xp>L2���)�bHd~OL�т����Tϗ�x�Î7Du,���O�z�:�"�F�_s#�2�vr�]��H!���B�:�T��$et��<6����٬�]x��G�<���m��*�,��V�E0_i��m_��<��b}��n8�=��
�Wu��=y���^��iTrK��zt�9&���ߓ,ďl�́*Pp�q�@(]5"%�S���v�o�W���ز��Qt����sT*�1����h.�z���q�����r�Ҋ��l�_b	�B���X�:�����"�%V�wt�Qރ�@� Q��%l-S��P�/�Q���nC2z�É������q��+V��ب�����:��qe4���~Ԁ��.W0���׿�A��?�1C��r����`�k�Y@� @���;�Ug��=ˎ�OK���E2�&کJK�P���������}/���	E�(y#nk&�1��6큣��#	c�����g��K�^�#	;�f"K�`�nn�|��d\n���E��r�L�w?��c�{G0�ӧO�����.��L0�{o�ޚ�C��he얱f{x��B΍9��	m^z��k(�Z.�T��=#}�pG(;�%l$��*���W�7�9�����g �6�.�S�X�b&0غ���9���=�D�*�,�|%ٛm�oB�L��-��T�����JbM��;���-��*M����Q,O�(�=^�3b�>S{G�q)~m�9kjz���!M��T��t�� nM��ȷ9
J�;�,��[7���Q"ܙ�|�j�=�w&��Mǭ8�������U`��_ʭu�ʁ�a"k
:xԄ��xF�4:
׍� 9��>�j��-����g�|A�]����Ŋ�$��U�ޓ$�;"J�a�����s��L��n��u� k��,/��<�n���[�!��A�!�&���
����:m6l� t,�R��� ϐJ�8P�u1t�&��,zd�f����H���@$�6]�8^s�l�kd�~^$���$ضg����k���I��Vr�-�Ð��3X��`Aȫ�n�����A��"���,�#~���kR��?�	�۷ň���� 8�������8���Y��-�_�L�J�v/j
�+��ړJ�K���7���XƊǵ�c�T���!mow2�=�qa_'z���B�y�E�Ϲ`�4���b��=�z��������Ȉ���jWs��p��`|0���N� L��"���mK��i��붩Q�g��Jb��5���_�:�I^C<3�j����U+ό�������\�=�W�1߇�˽_�ѽ���':��0�i��0c��~^��t�"�G���g�����(�yj�֘�]N��s1p�Ϫ���ﱬ���?����U��B�3b� 
E��u����ˡD?7�s�pް�ٜܴ�j�o�Yڂ�&\�~��{m
b'�˵Tl/�Ph��&?�ڀ@�%E`����؅`	 �p���Q)�����
�5�{���=���~��Ncq�����@���+9��f���h#�FtO���Y��D���x���D�FBK��m��!�=р��pM�E� ���V��gH�\5�	#�r㌲a|��Z}T�2v���F�| ��-�'���>m��"Jga�J0�?}��_����|���ƹ5��m�8$�cdh�xٸ ��f��e*1"��#{	�=����N��l����4됌{����IX����%���i\���?�?h��jMg����Y��M㭜]�q_�c�vK`��h��*R7[�2����i@�vf��{a�s�꛳"p�f�9"��j�Q���߲�;q]'�%���_�V�d�o��.��?d;6%��#,�z�m��`�k�{�E�˧O%��]�3�Λ)_n,GwG��1e��0�,|�X 6�����̓�s�P�#_"����r����?�<o�?�8��콻�V��9#���y�C>sQ�vz���M������=�_5p�`i�"��<��P����qI�2��V�8#WL4e���p�]3ɴ�Y�'��"��Õ\'}�-�N�I�W<��27Vj�X�7�=@'��M�]�(M��c�8U0������v�R�/��u*�	��I�C��AVR�}+9���6+�q���O�gv�\4��}��{�>����|�+|}/�������\;��iw�E�.v]QL�0>�3'���E������|��������T���]�R�-�u0�XU��5.���2t�PvF��i�?�<��)���5ݝ0'��߲҅q��x{�_8<�*�3��_��i_4��NfU����~j2!�}�� (�1'93��[���#���C�ǆ�|j��s�����E��X���Z��4�#�rT��D���R�h����H���un9s�1��5���-я�Í��<���Cu�u韣C�'M� U�,�)�rU$�G	����	��If�����\}f��֘T���k��i�͛ܢu�,�7kD��MU6L�NK�|<)Rg�(����[��8����E�FZ#W�W���{fڞ��'�OS�R2�s�Mt[��X�X �5k��"������Q�hH����%R� H��l$��t̻���19�x�m����T���흴�d Z�J�4���ᅛֶ�9 k���$�E�E�� ����O�;ZF�$ʾ�r�`���[	 ���v��Ҭ@�=��.d&AsT��@̹hV��;�y4�g��r�x<�X<?E'���q���3f�i�<����?�"���3	����5؈"�=v$���q4�	�ߑ��	c����>������}�*�w��xw'ח���ȷ���r ��{ ��t����4N7ϕ�I��@�	B�]z�[]+�d�A;�FB�~T��V��h0��t��md��r�u��u�T���P�[�k���#�ǙʫX�g�v�Q$�њ���2��<_��W8/�������?���8��G>"��~}�gs�:ҡv$��Rgҏ|���Îl�������7ǉ��</��mM��MQGF�X�*�5�M��%�ܧn�����AF�ABm��ϧ����SN����%�.��i-A��G�ݨ9���A�#&W�TՓ���3�B���%R�N�������H�e҉��1C����bۮ�S�)ʜ����ᆜ6,���S�Л�A��|~H�?������`h�t<�>x7K�k�Dow^�b���KuȠY.�,Y����u��1Y�ݖƱO����wPn{���T`�brÃ�ĝ��=!;���Z0�}�R���B��Zv�۱Y�>�o�qsW"�����~/z$��3����Qei���m�8#�g��0��IuT��y��Ԝ<9ڢ]*�%��G}��IB�XV%�r�r��՘ss{;��.Y9�!Ɛ�UԉYX��q�[}o0�]���⤅��y��l�L!��F��k�\�ϳ@,m����nF�ƣ;���|.C	2�X��)���~|9�Jqbty��~/_�~O�_^�"1�ܸ��v��<��#ʆ��=T�32����/���;���<�����p�8ѹe;ʎ�|�
�h��ξ��PL��P�wdX:$���r�|*����gĎԕi���
Y��b)���b���F�h�0�G��1��������E��4N� Y/����N��z�`�~��#�|������:��� -��d]]]�۷�������]��v���x'�i0�~�z�s֔gg6C�4���<�^i}�h���ȕ���+�������[��(|3��w<.�($�=;'9.�eL~���,��<^>�ׯr� ��X	���n��0.�`��Jdh��'�����ٸVa�<2�wwrs}��k%ΎZ�tт�!�C��Ьg�f�i�m�ײ��>�c����B#�D�1�4�z$|�T������Ʋ��(B���4F?������i�x,\��Ƹ�r<o��u�.]� 5��T�~(c ����N���i��۵�H�vBAF��`Z��dR�A+z�xf(SC'��4�B9�4�=T(a�!�p�5��jM������sJό�}�Sf�2Y����;k��y9W�=�-0���v���Ҏ�֦��5�M�ׯ�:�H����81����(�8�*A���h3�N�L|���@�,�v*�:?��cM�����y�#�0n��z+��RRT��<��z5J��'J��Q�U�����Q�r�Ҩ�����9z\'��#�K/u:�Uˠ$�w�ӗ.r���a���m���߸m��$�EBQt���x��19�E�RB�s-�Eb ���c��B��Wp��|*��'D���i+�J;���Z�]]ȪM�W:LԬh (��d�|j{48����v4��J�wuq�~��nd�f8�O��,9���Ѯ^2�HT����1�1,(6�A9������L�2�c(H��{Y0+j�|���Ymv�o��KA��J��~�s��i���"G��I�==�$�%5��,�̝̻��7ouΠKߴe���󁝩>;������>������w͜���c͍�k.�u;E:	0��-r݀݋x�Wt�6!JSE~��0D���p0��Y�����Fx����"�?{��d�E�^���S}�8������p������f�d�21�	-)R�f�?�4}��?˸� �H����y,�P<��f��q#�*"���d��*�[��9�fz�|>��b���i�@Fb��ɜ<=��1g������!)��r$�}���W��3�����Q�J̀����{�C���7<���S�Wש�5��{@��y}=_om�V?�JQZZ�Ȕ��"mb&�E�!�N4hc%Y�3�p0T��@��,�Qd�g�s�h�v�����{�a�d0��ii%1xAB���L���gu��T������,ژyP�5�`\�vҶ:c����K�>�����(�o���vs����wyqN'�G`ݼ�y/,�"c M``���kz���B��Y<��@8Q8�����yqlv`�]��,�A�Q�3!�FEi����d�g��d��64��m��M��l9[�D��0���A`(�� 
PL�bPǺu�$��h�jD@�Qb6#oFg�_}���H��?ҰF�3�@j���	�E�X��d~o�q��a���y��K`a��D:�t����-�N���{�"�C--�wɧpP��8���z��}h�R��g=�	� J�8���4��m�f�ap�uo)�\Ҳ����|;��4�FD���P��������O�8�����EX��������5���т�&GNu���_�x�~����W���[����kͳ�9Bujl4tu�"L>0���!?�������a�9��^��N�(�}l3�@M���gL�L���4�ќ~*��6��w�2����ʢ�+{�H���`l�m��b���u�xl'FG^�RO_��@PX�iL>*A��J��!s�@.#��v����l�hii�e���5K���ה��w����f�юT�*|��|����o%�i7���F���,�AB��9��ϓ�[�$;���I����Gc�=��v�\����Ѿ��s塇���%�^=�~����5m>ڟ��<J)�r>�"���6p����g��#6�dQ��4�ӛ}@tm�����"W� I���C���%iZ�H����q�Dn"��퀝�n�쎪�!�R��6� �"F'���g�W#v�kv(~�o:�G��Ԫ4oVteaoc���mv�^9��>O>��A���1��W� z��gux~�	��&	��`1�\9��Z���̘�`Jk��ٓKg�6��������������\Ѕ�-_�ű�>�R́�(�����΃����_l�1=6�L+m��[TA�Pu�
2
��uٜ,��g���3Bu���Z6~�)�K}�#;�[��Q\��p+�1bcΨ}y!�=�w?9��`��s��S��ϳ�T�zǚ��e��Y��;��6������K�;/����*S:�V��D����kF_-%�WJ�,喹�줹k�}?�9�j�q��G�.�E�u��$�d��=C�F�"��.c�!���ݕv���NST���h*�z�v.��~{����^��*R�e�
�]p
����Ȥ}:5�0� �<���>4�|�L<?��?���p��a�|T��ZE򸰍sTco��������پ�i�4+j��U2��72\͂h�IA����@�N�c����F�eh���������g��%	�b]p��(���<m�l�A�Ԋď+� ���sbN��f�Va�g���2A&���W�Ʒ�3��Q��&�)��GC��E��K�j�M���B訐�bY�~�.��q�R*-M��`h;����Ȭ	g_-�l�eY�u)�5^�\�h�/�~��O���Y�� ��r���m�kY����M�F*�MeX�1��.4���"�1��9�R1�����FP���<`��Hp�.f�Y@�������B�������-J���-��}L��@d�u="$��=C��m�-���8rH�t��xF�)�+˶�9Sn��dǋ���l]g�R첐��ˊz�9��9b��|U��P��Jf���IA؜:���9�M��P���dd]�+��|'�H�՗S���9^U��_�+���e@�1k;J���|Ʈ�8N�G��F:��4�����G�'M�X0!Vz�>�U��W)��'�f��s�A�h��H�ɑ�0�f�Zbg���_B����|&C}���v?Ղ��J���c|��>���N�ns�����\1�}���*�Pl �c�~ϟ�ؖ����d��Z*4&C��K�G�$s(]���i���@�]�w��b�>Aߤ�I��v"H� �.�\֘��"UQ��w��;������C��pβ%�F�n�^X����{�|���V>�����Lή/���I�K�z��ƘD��N�p�K����m�C�����%{�k4���{IX�ShF|�+!W�9M^���]KZɰ4}���ȓ�pO;�t������$?^�����#*F�[g�ן�^�K�l0�O��&=�Q���xM�\��	�N�)���k��ȱ��+/�a/�ߺ=���Y�k�e�|�0��ѱ�w&Λ9�9b~40�4\������xs�[	J�ƹ}��pw8 �X���NM;��T�O"3�ކ5F����FQjd��0�@((���sc�3W*�,ap�ì�#Xf�Z&epΟ�<�,�B�ѻ��mv���I	�(K��]	p�2U��<,?��O�5#zP��ǩ��E�(x�V���*Z$� \�ǜ�A#��c���AƝDD��\̡��ޘ�de��|�����AF�O�p�+R>��~v���܈�s��j9���<��L@L��1�}�`0 ߻�~>y��7�-���ʨx���|L��cvع6�J�$hW ^�x=ȡ�\�ř�HS��VJ,MI2�g@[-����y�W �nh+��"B�敮C��,+�|`����F}+Tj��,	�.
��vz�:����LOy����k�7���yq:�ı��3��Oˡ��&�ū�
$��fN%Lƅ{[���nT ��� D���㏄2��X�<J�6���܆,=��8� bfa�6������<��J�G�_AЅA#p�����ƃƮ����J����<,gW�rw{'��=@� �r��h���=��B�1p�t�^YW�k�p{�����{k������F�gg�,�I��k�u�R����f�Q7򸁄�~$���h��r���!K�А�c�[��˔p��^�k%��K���n��ׂ3@-�c�?@����Mz���l���Ͽ�"����_��|vz	��b�OsY����h�"���8d�$AP��=�.Ƞ�3 ��Z����*�$�D�Yه�G���gl�繑��=��7����{b h���q\���٪4<��4T���hZ�}�׏ַ���!�8�[ɝ>�FY�+���l�i�,�w����;�e��Ev�ˇ��T���j��[k3�QՅ�N^�{_�(����m<���9�����<@��0�d����%Ww6�lãk�3X|u���8�V4^K��`�B�ʜ%�����Z/�6�s0V��2X��&�_�n���2�f������P&է�Ԃ(����wp�����|9n(TϦ��R(�D�$V1��E���ABA���,Q�lo7�󘮣)c�:y��T?��#��������L�!��H�a۴�
���<-*���.��Q�4i3�/�S(��v�i �O�Ѕp� ���n��@��%/nJ�q�
A���>�u�C����aY-y���;;�S���E�������\�;yO}��=��Q��{f�����vL4P��AQ��[P������f~U�9.>������;�C�х��`���B�}����4k:4 �:ni���YX91�#�9^Ά�9;[ʪI~f��P�ҵ`���E	��������	e휒��x����EGy�E]�M��o�Nv����R��B���^g1�e��7n��o��
�� ��ʂҝԎ���lYۧ�F3�j��>_˵���Y��W��W94@d�9�F�^�e-�ÊE^zf��\3Cn�n��A��͢8еm��0���l��5ӟm㿻 ��8��	�6�54��A/��&L��܊�gE!�Έ�{�F_�]�cT"3��-h�\^������E��T+�!"��(�?	��P�i@sk$N�t�B=_^��}�(sH� �^[�g��7�%~�l��9��V%<7������FK"���3J��R3,��1:j�}��e0t�vh�L�F��]�� ���ڬfme�4���,K���F�>�hnFC�.�:m��O<
j�s5�!�q��8˕Š���Z�A���M޶��)*�h=�$fĄ�fe�����,�
��|PdI�0"��J^��^	�
ڂ��|�	�;��l�9�])��`ݥ�A'D��%�ź]�nȔ��C s��{,]�o)��`]�4�ϥ�@��Ԍ�A�3�c�[b_��o��7H�i\�֖�Kk���
H�>Ȼwچ����O�Q�e^g��:#��Z8�M�g�����o;�{-���r��$��A��?Cnk|V����%�h�qDˌ�& J�K���� h�V����Z0!3	�k��؝v��U�\3�� ���"�98j�9����,��\-9s爠V9�|�\� گ:�VҪ���N �Vޭ*UYA2?a0�����^�u������T��v�lv�u��~�s��d؟u\#�u�����)2�R�"��q�KH��2�����մQK��G�Ŭ�N.��� �[A��fx٨���r��i�k���UaQt����2b��Đ	T�Q"��}���ӿ�v�+�$��NZ��3�0r��UrW� :I�������Tc9L˱���v��we���J�+��2��IV�ѩ4���B�=��z�P�!O��gxd�T���D��LK�A�$}ӵ49��#SCE�R�ި��ιy����0�=Y<s���0�ј���.>�k�A݌
Y��IG�}�w�(;}�@4g�^�k��*�
�<4��M�s����j�����(2�j�Q�͎����Jc�y�ZM��������P�s~A�d:�;�S/T~	��`��q��k��!顖�9_�|��U�{���G@c�l�4G���2[�ja��jy�ܿ����?r�.�l��`��5�w����ߣ�{C��R�ۯ�r�d ;Z�s5I��͚p���q=j>�U!D�ɉ���B���'E�*��V�r0ݯ<�� 3� D5���ބ��@�*�m�D:�&]�r5�I�9��c156��20&�"�2~��\���������wUgN}zJ�MEM(o�g�S/�����}�O}fv����r;D"v��Fpgi���q頡�2\��T8T���v$U�0�8���Ap9&�A�|�&���2����pӂi|��[�X[ݜY����c?;�v�h�g^�9"ؑ⸚�:9��1�P5s�1W���4��E]�+G��8X"���D2����,�.�A,0��Τ63y��ĨG�J"f��E��y��R���'m!\1�g�U�z�/\G/�;<�s��AU�56 y�q����N=k='CQ4��j�� �/�I-aj3"��0�zsحgp�����7�M�CܙӋ`����}@j��kl����PJ"R8Y��J�u��iP�mm��������m��n�b�(*���l3�p��Jچ���Z&ӻ�������w9{��5��p�c���u�˽ �m¢ۘ��p�t]\���6�F��J3R�x4`�-��<BFj+�����qe (h�op�_k�M���d�!�y �I:%8l����A��S|���R�+�MFSr��%��@�!c����ӂ���
��y�b�ö,��%thsz}������m�m��IG�n�� !�� A�L ���֜꘱�@λH�vYV����3��/Znx���!G�Ϝ�Q΃��\3��"�Dă�_�&@� +I�t�r���V�Y��[i�F�V�A���M�~���V�0f�(�{��lL����b-ޱ��޽7���E�[ߪ\ix]}��uj�������ޟ��`]]�h����B9
����.���	d�9߽/o޾�{�/�h��=ܧ�I.��MF=�v�T�	��-�V�����8H� c��/�4�!UѨ %����9�o�:�ʺN�K��r�9ԏ>��8�Sma��C$Gk8��:QԎ��*���v��vɬX_V��Jk���o�Rm�W�u��8v�Tc!���}�Ү��6�"�|���G����+-�h�>�z���B�BCNv��1O��3t�&�
�M~��I����o߰���"e�^�u�ra|��N�3��1��_��:��A���NGccϨ*}<5t�JF>E�LU�Ã C�$��SOFcO:��q�����h�A8dY��2�˭u��,H�H�R���"�o�5��Xr,���.�n�G�+n�����M{C�Ub�l%nhT;�����8�	���:j�H6��;��@���]�)Γ-s�&��h�l�i���PO@�����hT��s?\盫�/n����s�3ɖ�>�����̷i��Ч�r��Y�h����R&���`2�6E�X�To�}!�gi4�~�F�9g���TGi>,��=BZ��'�/�:���*$q6h	�����\����$����]����([A�T�}~�]`B�¯�Ӕ�l̗����0V|Ek���.�/�1\�y:3Zos�EUw���"?���{���5�Ck�a�z�x����,-u���<]�c���0�����S@��:�b!����W�K���f�a�D����J����x�,����d��䚢t��5:�%�����QL!�3�d8�Jt��i�yU�rkrZ7�[�E3�-7�������u4q,�ql.�~܃Ζ�<�</��S9R2R�����v��!羢��`��A��ʗ�-�l���	����;�'+7&sn<�*S��hj؄��CP�[CD���}b���k��-ZUX@�4!�(g��cF��i�b~_���M�R�X< �����;kk�MtJ2d���,0l�I�!��)�l�K��ʤrKj��o4+����"do�繡n�d�?����^/%s���NA�u�\=��<0'[�� �xm�����F`H6�`�M��m2z�����ip��y��H6l2�{���Ó|���ݦ�hAi�%�hq��dւe��8��`��:L�֫���g!���4k��)��5�t��|jA�C�xr�(���k�.����X8q��}���m���� N{�tXa�$���ɝ�z�^��:?'�%M�!q�;s��Z�3����8Sd�`V��h{R܇UpK��鳓y0ع�e���
d����Z�򾱀�;�In��ȓ���fdP.�"��VVw�>ڢ�,y�ۈ�Y9/W���hD�'/�Xۘ2�,@4���ʣekk�"ș����e��q���N�"(���H����L�3B��#��=������Uz?R���Kt�1��Y:�6�G�=����Z-]$�&��E%�Vq�V>�V"�7��dR;5B�R�:e/������sV��0s�Oj<_�G(�?iл<������	��FJ��w�^q^Ñ���g��5[e��n�/tQ}��^߱_w��x���S��`±P������ƞ?TG��O9גA�ֹ&_yNr�X�n(x`�4��5�:L��rBƺG���]!�};栶��u1��*e���#O
�=�7!�}�Cȼ<~��|�/�9'������NU��	�G6�̨�װir�*�~���Am=JOd������7y-��(6���&�i�/'��qPV;5��&������)�F4}9ׁ�-�������r�YୌK�M�Ms4��7�{��r �����zb�|2HhΙ xx:�T�;Q�� ��"}ޮ�[��x�y��!*��`���(-�^�pO��HV�Z`��li��ۮ'u������t�v��$|��ݿ�l�KS��A	����е� �k��P��_��Ll�͹6H`J�x��eXOߒ���ٲh��RM�Q���Fx���>Y(d��N�h��CNF�ZML4Q:�vʻϼ�;��Ɨޯ�m5��1��X;�B��kX�%�4[�XH��Νc�&c� ��s*'`}a`��h=C�$8e�a/���l��I�0}nh���$���fƍyG��w�*ZZ�V+�<�|�D���!oY�^�"Mu�m<-�����EɈw5�h����Zi���~S��@!����9�X���t+�̳�"�-�%�U�0��q�L�r=�����&ω1Ͽj��6Z&h�D�^��'��t<�q*{ߵ�2eG�rGJk�*��+�����T���Nד�e4M1$*�b�����?�ٜ�:ɬmf�[����s�:�8��ɓ96}E���X���R�)�z,���]�8Aw�ߌ�$�{�<����*���Y������d�B��DEXM��?g��N�^��e���Ī^o_��!h��%����u�_�^�hs�p+����?l�9�"�Ԙ44c� �#�3� Q�������;7o�ǲF�
ʂM���p�1N(���U��<���5o�M�f<H�	l�������;�r@� �-^8�U�	y�,�ׯ_�t/8���
���ΘY�p�dh�#i���N?�(;k���r��}��@��������h �Aoe=��:J�f�P/+]�NQV��Rj,"��2�%���9�<W���!3�r����{"X�����:[OE����ie���ܥ}���ip�QO�8�����dt��83L�N�5�|N��M>�Y.�cc��˾S�g /���c?�0������3Ǆl^!p�}1/W���Œ��lE� <?��kY��"X��2ݧ=uv&[�c%��W? �K��a��r��y�e��D��?�V�.�Ѿs�W�}��\���l�(�y��m�b\�����6�á�%����+8�����k�;���QJl��ge��ӤV}?֜"�����|,O\��u�48���g�s�y�"0��*�Rm╒�e�H��V���t���ю�$!�T�ܚr�i=(ҭ�ZcH?���`�טm�Ѣ�;�6]�(vr���tyTJ��
��Ό+d�7��q�ď���;>�������֫�m�����{��j��e0��vd�)jG��sB����;�"��#ꤳɊ=T�}���i�F�,���v|�&}T%���2W����u�f�������Oh��$�HT�֩�
�������t�C�J��Bp�%�i���8]���)�ޒ�t@I-w{��$��� ڧ�����:ExfڀX٩>�R>���ݞm��h6u��sm%�N��M/2ϑ�8����H�4Z����.���Ǥ��M�ц&���j%ò_rJ��6���"u2'�;�)�����]�^���穭H���`��Ǽo�ut��龟����)����EfvQۍ�R��cy���~L�:V�q��������� <��\(�BHYXI����~��k�k���H��9c�@�=��Ш���{�rH���v�,�8EFk�H���l0��*�GK���l ����5�%�[���0�e�����L�݃l���B7��p���Fόh��J�]���H���[�&�'2�$iI�R;��wd�[ur�
�9lr;�Q@L5Xv�C	vi��Ɏ8���淃|�tr�e?T0ǻT��=w�C=/��"�k��@{F���;-kj�M�3��Z�0��q4I�\H&�}�%�<>��e�����
��68�� ��?�O|�@Q@~��-��@�GRU
�k�mW�L/�9��%�Xל3P�1��J?�1:C(Xg������3_[h�%�T��S�ʐ����h.�픛�b�����
���[����q$L���2e�;T�R���M��2C!������$�(%pf<���M��}r������Ϲ����o3����P8����/�K��?���߳>A�"%"�t�W�Ւ3>�</��h��5�K�,�g%��G�-%�ch�~P' ������c����q�с)ͅO�?Q��˿�����-��<���}zݲ��#�J�e���%ɻ[5��BP$�=�J���B��d����9����ai�w��-�;���А�7h���sl���%!�1 ����ȗ�Q���{~����Ge�~�c�Z��姿����39Ư3؜�� �n�ݪ@.��s�����R<:�7�u=�	)}VK펆R���_�Vq]h�
�=i<�����<`����YF��i\\}���Fw� 桓�}z��Mz�y!n���'�!�nΝ��M�H�::��سN9������L3�]Gy�'Y������5�r��-��s+]���4)RD(h���yZ�J
�F����k�y(*n�6�	��S�ý����ĘL��f%�*�����M�yO�/�FI�$�ne�Yc�S����xN���dhT��ɺ�>�d$h|ƙ���?�3w�>�2���9[�ھ��=�N���(�6+Е�J����ai���+���0�q�X�+��0�H��J����1"�= �\6,��Hv8h�X��]����K�{��\��,��6~"��{��W�ю�{��7����4�D��ǋh�T\O�cy�U��Q��@�9���w��2D�j���N���a���g��|��1��E��E�8�>;B�/���zECz���+�|^$xfy5���|�=m�E�e+����V0��'6,[Gbȝh�J���#���͉�	���	;k�!";e�y��7���{Y���1}�OI_�[z=$���}rG�N�=�&U����s�L�h�E���H�xB�}>"��W�}�\;���:�v�[czg+��-W-	@�®yH:zz���Vr�J���L��4�o�,ᨢ1�˳�.R���m���Vy�������Vub�����!��8�����;�xLxD?�ܩ�X�pe7,�Fh�?�J�2�y񗘎x�9��+������sΌ�����%H��r�;��Vgi�#B����Ez��	�_8�y�:�O���~�d�*9n�%�%y���6v�9�^�f�zC��V!����D��ؠ�5��nYG0�E_z�jF/���{�Z�����t/���(���ꌮ�|}��	� ԙ�x%!i�j� |޸%鞶�=АV�B�I��Jʙ��5n)�-��'*k� =Q�N�^�$;T��C�S��oSQ��}"fǧ^K�Y��+r�ܢ��k��j��G:m�7e�,�g��$g�ᑥ�<�9������Ɖf8٨,6��l�*��8	��]WJ�6d�}�D�4XV��v �U�%/�)9��i�~����|�����]z=��<#�A�$kVޚϷG7�M�g�@��Y';39l;��PTFo�&4�F���Yj���~��&CS�g� ��xk[�%9n�m$�aw�m�ӵ�{{.�ߝsp�%�{����-�@!4hr��x`M�zp'T��`�Dz��ǹ9�!	�;Д��g����s�3�
�Gg��ɩ����Zֵ/�}�!!2������(�d��%�=f����>y]Xh��l�.U��~0����|7F{+�B�e�� P;���������(ׁ� _d��^l�s��E��X�K+'�}��!�AZC��K��7�O46�l@���J&���h�yK8�̹sh.�\2h`p��G�o���o߽�9������B���ᗤ�j!��ן�j�3C�D�21`�x��8nў�W���ݎ|Ӏ`k\E�(;8٦!f��Ÿ�'#�`�ׅ`����������ۯD�<�8��{�6��������Ը�����F�f���S���]܁���*�T�v�O��ƍ� U�H�[��@� �/�W}�t!8��텼}s�`&�k��Y>$��I84���3�#���g|�s��T"v���H��n�N��\cSn�Ukp|��30P]ֱC�A��*3O2��N~T�?���/P�� b�ݙ O���Ǩ��oQZ��r؊^DY�8T>m��V�S٬�ޯ�
�A�K�<n5��~@�)Z�ĴHP�;`��]�ۋ���H��a۬><���]h�����ĈWrdƨ��ڭ��ГD�Zp6%�:,.��Kzuex]��IW-�Ɉr_xF�hA��jU7"vVfそb�kl6Ț��c!��4����ʱ#&���u���yN�xK�[����,kF���l�,_LuY '����=\d��=�]٬vN����0
%Z d�����k��>�ҚA2sMΙ�e����K�Yƕlρ���.�H�A����A�.�̓���3rŵl��?(g� H. ���
@��6����/b|�޾�p���}Iv79�bf�7V�5xi�x�f��h��=�7��KB�<W���Q��4�H@���'�c�+Y��9�6�I�k2�q��9J���џ��`��C%3��6������qr:+��%�`[L���Y��ܳ��9�Μ�i�sf��^����9��-�s�{����g'>°��+Qᅌ{�n��N1�)��Z���je]шXɮ�-h-��~����;�o����!t{�p�wo��۴�e��������+,��O���/�F�+e�f��)�;�$�p�2"\_�/N��E&��Ό+���/�<U*�*������c��b�Yvtv�<������ ��N��eǀ�6-꧇�����=��77����&)�sF�.�{�Μ?�uG�����(/K���1��grt�m(Y��Q�(�}rv�;-i����G���OQ��q]�d·�͔[�_��я�	�|J�J���~����>g�:�
V�2dC��%�q٤��/i���)��i�v�˦����Y*��;Sz]�Q�-ߊ�	ft��$D
1����LO��9��<�,�K��ЊR���f���>���r���H�Q7�wϟ��!h�]Z�!VC�f39���Z.9�˄H�Td�Ҹ-�hQ�.�v�+U
:wG�͠�mTrCm���Eoe5�9�Or�q���u�Ȑ:��o�A��@@����>9�_�$!������P�|R�k������$ۜѝAe�����Q���r�lzƜ�3�;?_����
m�/.�86?}�_~�Y���?3+vw�5���@N����u����$���Cy8���I�Cc����c#P���Go#D��>�6[���������%?�����ؽ
-�Њ$��lX;Z5D�p���`2׵�`C90��,�d���F^��DDΖ��u�χ�x]ۄ�����]e�f.�n���~{b��@���x��h�w�6��!�� ���(���½����v9�'�����>�SzI�#w��<����4�^||?�Dfヲ�?�2r�^@�I)�R��u�c׎ˆ���W�A��6�� �:m�� !t2��<Y�]&��%*�;ġ,���X!p{��a�2���/� @�� ���A`W�-���a������]��´�a/�$j���/���?��,�b/�[�v�m�T�*��2�*��Iq�]�V�����a	�xtx�'��\�9�xF�̘ı�:�����2���۫t�N�P�g��-��mCq���/�jI޻�2Ð��}��J,�M]U%"iK1:d�]׿u�����<M��]�����?�ֻ��A��㯿&��(���%���g�K�/�ɛ�쁕�"9e�~��hO�����f���>Z4%q�@���g녠�g�$���(jr��VE���jE�Gd#�X�Յʁ"*�T8�^N�Zwh=w<������n�	�j�i���"�N^�.���3��J�<1F���$��~[,��d����5�Ku3Ɓ�fԨ'w|�iW�2��X�cu���^�/�2�V�-��!�͠"���@f��A��q����R�oӵl������gy��-�1�₉o��XhB���@hj{���@7Q]k�s!���� _-V��tmon�$��k�2$�'c$  �0&П�?=telɏT�_���ʞLo�?�5_�z�Ş�w]Z�E�g ��A2���F 6�lgJ]_�������w꠫%ַ&O�L/�g�e�����/��@V�*�T����G�g2��U��C��s�o�۶E�B�1-��}�z�)���H-��j�5�=���;��Z�:��GIєW'�H74B���QR9��:m'�M�@�5y�����_�����#����o������!���Cr>>��������."�:�c2��b�Cp��@;Yr�)WG�ok�a
���T��
���ri��A��:��������1�!h�p����@�ɫ���������ɏ?�>9Z�$'���&9��>��UL�"9h�v�� !��H�69����C+xr(����C)Sn��֯r xc���t0�� ƞ���q�0#P-�z&�R??_�1��g!�05�^�{�GA�����ر|�<+b[)d1��U��y7f\Th]�gX떯�Q��J-;��9�*TR6س�|��*�fY Cx'.9�1XiN8yԱ����2?sp�b4�	�+̿�J�~n��yz��Y�����X��9�r�Gӹ�9� �!-���X7���A3����{�v�9 1$�q�2~O�� /�k����{x���v�-����'����ָW�_����h��>��*bh���񮅢��	�e���'zk/�d�*�I����Y��Ą��+���wɰz���D�� L�駟�O����1�'o�P��G��
oĜu��݃3���3����h���zc���Y�}2��|����4�`��@|h Aġ/p���~����� 7��M��&��.�{�<|��:~�GX�ˎ�^ αc���Mm���N�Y�`:������L����sM��%
(�B����5><��Y|��[�������}���O�>������8f�z`��h{x��������I y\*'i�o����~����g�:0��z<# ��~�d���j@����j�]�:�y4��>���D�$U|�{�/Ә<1��Y�gg����z�;��G�9�D�v[�a8�.�	�٦w��@T+�x� �$���8���n!��k�g=�Q�a�{jx�S� /���0V��	K+խeyA�fvpr� �,O�J�ޯ�C���##}�և�Gr��� ����=�c��Q�T��|��~�K̾��0����؀�t7m�ؗ��D�,/�@�u���6R�*�/(ˢ�r�%5�;�}�h3�z�?ƕ�����\���`�Z&��;��T����3�q�ݓ%�PFy�Z��fZ�6&'3��R�v�>�n:yD,����v�uxYb�@��FK�٪�џ1>�sl9>@T�]���\6�ʝq�2��*282�E��0�^��~^�{��^XN��"��+�Ʒכ3=h�Ѷj�ʘ��q.�i�!V������A/�o�cx`Gy'"���b���͉:��n���t�7
]c�/].u�ښkH)t\zC7z�˅�� �3�EI��~�˟^r5/�b)P�ҵ?�����7D�$�h~��Ly咽��E�}���l4`����l��V��w���"����噜�4N�e�#��Rr���.��
I��.��C�A������Mz�2	͵���m�έZևn]����1�4g��5�+{�F`精�|��uI�l:vp���zE���J�D�_��o�ZtC#�����}��!��/��z���#�֝u������?����^���	φ�]����dz%��= ���{l?��߰�P��h�����[��'�2"���Z���#��g.�c�E����	�����}�h: ���~
=?����<ʗ�?'����� ��r!������  w������xJ��egנ�l�r��B�VϺ���#)@E�-h�w8	X�OOkmї�'Q�v��}�]*��C)e��w�(jxl� d5]G2,�m;:��eA$ ]��������NP��|�p��.p�ŝso�\��WӁ�|h�H����1d���K4� CE�<Es*���&��P�a`��vOOg|������-3hj���^s�Nc���2��� �A1`����i��S�<L;�?C�I߁�պ!����[�6r�4A��2�+\7XV������	�'��M�9G���t���qr~��ۛ~���L6�!9�;-���PSt���d�49��1�ig$�D�yFʸ����J�����>ؚ�4�u}PCmխx<WI�n�(�vA��R4kԳlD�8��t��	��dK����M�A�)ÎA��a�4�cc�N(c�{��0��� �X�/�Ɉ!�H���ϋX}Ϗ����w�ry���<"� R�{�?���<8gXO4H�^
��і�:��[���#�$׽]<ə��+�<n�vqK�
CD E6ۭ��6`>��Ap>!�ruyE�D�?�e�o `���a5��6�ey珏�h%T��A ���R���L�-q�Yp�9��k�z��M@B�.ҵ�];�O�'�p���#�:����K����O���'��^_�|Uc<V���=׹������o��;����3G�Y�Ac�ȯ��)�.�*GP>�v��#���8l��>���Y��Q�a l��k�_�?Ngݴ�#�YG�=K���������M�����7t�IT-�yM��#�����A����|�:�,c�%p\
����3������y�%"r�
�σoFKb��UY�:��N�g�,�"�]w����P-0.A�#2�ѽ�ULڝ���� 1��w�ݟއ�c9����3��K�� fû)I��~�~�ޘ�_zKD��Ca"h���"ˇ�Uw`��ѽ5!ס�y���-5E	W[� Ro�"��6ٕ������xj.��]Ѧ���J�n�$��6(��a��S��c�k�*ue-�{}�,Q�D�kf���i;#iy��r���;��;�Pf
}�m�Q�T�#`�t:j�+��i��b:/ֶvc��B�{�2U vE�H�wO�y�7PaY$�Eޔ0��Vs-Lk�N�ڱ����2���J�hh@��ykQ޿{#���Wy���������v&6�5��6�9(.2*t�_�� |�]��Yp��^DJ�|�Uχ�;~���X�}�R'm�6��ܳ��)�bNՑd�j��e$��;$ғ�^��l�JE��(-�<Df~��!=�3�t �w$�X��)fK����Z?��3ѫ���w�Ǡ�@gO�һd�4Q_k�j�����n�k��\�sm#88�����>�߫��������Q�Q�x��Ye���{
O�s�wٱ�㦼DKv�y�:w@�<�S�A��JhC-��"�+�嘋�9=���l��+���j5��&���Τ+~6�x��g�c<��m����)[Q��T�u�fK��U�:
���w}f#���
]V����P#��m	�4mǈ0j���@.�Y>}�w���������U���4�;&-��ӣ�@C9 �رx�"��8��]A�#PW,��Z���v�Hž�-����9�I#�W�z���ց�?�̓Ƹ�u�+��V82�R��trr�;#�� ���U�9}���;�9d��@�=D�����͎�y����oBQxyV��ɂ���F��'v�0:։�L�3��)1��&����w�󏷰t#�+�w�P�"�K,	�l�t�
��O�V�jرEc4'ӌ/�!�x��GԱ)�[f�GVH2�e3�3��ugN��h��q@B�\�_CA9Y����.��� ��yQ\~�zgɒA��Fh�vò�9V� J#�!i��N�z�2������Y�A'<�]�A  ���"��%ב�ޓ�1Z�7�A8�پ<q���'�gˠ=�q~H�y��\�氆ƽ�J��ӒK
�w�)�W�I��	���H�M�I���f�V��x���&ۀ'#H�:ak��(
E[��^�SP^��g-�V:�,��ZyB��v�d=%9�k���0���r?�%b�I�n���9�a�/�#k��$�@�d@���m9G�Ye�k�)��,ͣ��5ruy��w���;V���vv�8�s/f�Yp%�U4�HvD� d~��ۯw��������K}vJV����(�e�p�3V�������#{B���!����=�&��k�O���H���޶d�uw���/$Pr��8tD$7 p���|�lf�����s���	{��s�\ǜ8j��8 ���@�@:d��	�@���I�C�+聺�ip��O�YH���'ޗ��4%��V�8\.V6W-{���iԹ[�\
$?�27����.���w�g�s��#���A� -�{��y����
�TS4�x�
4G?Q��ρ����� �lPǕD�Z������C� ���&���>��Ir!��N�O��"-�V�;�6��Re������<����$����D��wDX��7L ��K�9�tlc��>[w@��H$2���F��FE������u�)9hR��h���L�䘄I�3�b��W���� i��Ѥ����ς<|�Fg`
zp���ظ����JS0~@%݋�(�"��I����;���<��M;�"�^"���+�mi��zG]���I�]].�_��?�?��?�a��ׯ���R>|�l	�	v�@�s�F�\ls�)�#0ƹmL��}�y�P�0�����5��5�H�3y�v-��W�����]��x  ���� �g�8��O�z��M:������.V���XvTYz=�9���,gƍ
�9��p��\]^�s��x#����Y�^9��d)ht��%� ���h�N��X��X�Y�Ҏ��CKt+�[�bכ#�K����r}��8s~y2�:;�R�$C�r���Hl2�"��Ҽ�hs�?�1�d�`j��ܖ��i�6���)>d�G6�����'�;l�1��;Ӳ{SA"���ڔ���}��:�xU��1�a���;�ݼr�[犭��P>�J<��� �ߦ���8�<B��[��t�=_��H���(�� ����)|�tD���������޺�HP�	%ҍ�<S;��n����O!9����w�,��Nh����� ��
���Y�����NjF �OLާ��li�h9jY�,�I8֛�epZ+y��Т@�ql����nhT3��-ڤ�L4��~c�vу����Y��Z
�H��pr�y���e.�l�����oL�k<���$���y;�ϭp�郴һ�"먎"��w7Akǵ=�"v�R~�Y6�#I�F7�x�@�ao� ^��P^i�I�9s��l���);SX��x�$+,G�M��C����6�7^_y=ww_��M��ϼnt�u7��Z�HEN`�Z�e�'��匲�;��;:'��g�KB �0���A��o=�Rc�d��C71�N�u�p�=�3�����"��.�?�!��"��`���G1����@����Z�r�����B9�^�;����~��+�D�����˿�"�@8v=� 8�n���Noz�d���T�7�=��d�5��0�`������e��E�b��v1l�!MG��d,�I߃�����YK���c`����]D�=Q�����t��e�����݂��������{3��T�yH2z��F��> 2�_�;����i0�Ç_�׏��^K�`x�kh��`��õ� suG\$�8�޽����N�?2ι2��M�:�u財�D�4��\"����]r���y�����$�XC�����TC�$\V��;���=�ER�u���,�L���N5��[����C��ȶJpHe�&���)��٭���<mX���S��Mz��c��E�_��9dd����%)A������U��)t���Z,SY;��ّQ�-���ɶ�a��2@�S��Z}�=�9ذ����}<(�$_y}In�V���0��F���Pގ&�<�c(;>����M�:�/Ð�M�T:������ĉn��F�-��h,��|*~��*�e@jdG��/�~&WU'8� �����}.?��2�!�C��ρ���ö �MZ�K�)z�G)M���]d[���^���-�<z�p�	QE"�Hf�A!D���!���n�ڒ��Ӄ��+;"i���>�8!�����A |��_�S��v�eL���\���L�x4��'U�q���f�D�+To{��|\�#92�����7mrɲ�����rQfeu���c6���Ę�|y�m�]�i�P�$��9wqH�Bʬz�TD� ��]�=7l�f���x�o?�ۛ����C��tɠy&;��`X	.5 �͠�+KV�G&^�fC[	b�%9/yH��]����@�w7���Թ�5�^fJ:1A���.h�=�(��PF�e}�[�٬�I� �2�J��c��7�G������x�DR�I�s�5@p�s�!�$����97������?���l���9���[x��C�������S�_�i�H�M��/ZG�'m͎f/k�a,�V���V�jc�f,�/�2Z��t�RlAd�!N(��e����< g�5ʯAw�I�V:Q��ݣ��_m�<�):����
�?��[�W{�8��[���	[��'�?�Dy����J���̋�v���	�]���?�c'H��fn��eK�Ν@U��'i�ǎ�J���K�4�/�18������5^�$�$֎�X-��"��=���@X� v�o�P�hI�ؔ�U�:<�h��Ln��hx�EvrV��T�7�ZW����$��s4(U
�QJ�!J���Rɓb\Z�=��P@%�$���Br�S�Z�#�g3�`�垓��eّYj�Q.���Z��â�� ��ͨ��m	�SOƤ�&�\F��߽M���5�j~'��ם@�p�K���f��ք&�+&-KS�Ă��m��<wE��N��Fԩ���'B i�Q݃���:в#�ri��xn��d�|�2N�{�u,*���b8c�0�Ϳ���Y��Z�(�܁����v<GFcs]��p�;-{#I^� bl�C�%3�f����A�,dkJ��~�5R=p�,�5[DG�9��l'r�����u(JP���q}�%��k'�o�N���z>�P�Wb5�
�!wL�ٗGZE�('V(�/ӣRz��S=g�Q�nN(�A)���!�-�ӯ�yS�T��LהN{}�:�42�B��\<u�Xg�s�|�k`K��a8=?#4��qL8��H�7�bp��@
rM0�����=�ు����N5B���$�޳�!h�?J��^	y74�N�
���5Q9��8s�3A�	rr����!4Y敍x�q~�����/�d��S��3H�����h[v�[�f�8���~��� |��W>c�����r$�"����/���1�mȟ�2�F\�<\�Z�����2���R· x�j$uO�F>�>p�C߂�z��^	�.4m�6��L�6%�]|7�$u�Xr���J�${����*;&7��9{�����PJ��b�X��
D[��M�P-�j���{4=��b��oG���ǬNI0X��F�ľ�0M�&�Z�ج�T�o~s�k������������TbW�i$p���`��_UI�vD��`��`R���NK;M�-�Z�<�%j���8��K��1h�'����{{^��#�-P��q]��]2fG�,;�7Y&�X�B]��K$�~�=8f)h��IP4�I�ǲ�_��;SB�!X���ƸN�Utr.�Ć��#A�u,��7١�;�A�L�7i�U��@���·k6G9>��l	��@� ��r�j]�gh�i0k:��ߛ�.O@��o�8TL.''�w���!Sqh�?�[����᷀��������߽�z�]����'W�PA�ۂ��/��1���Z�s$ؕ�yD�3m��<���#��"{O�*Ll�\܄�]~�5h��H��Y���37��4��*_s�g��(��C��f�P�Sv(-�Q���;�؁�e���м��T��r�Dv��|	,-\�g�_���g�'<�ӡ�����X�PD쌝[e�XL2$ԲI�i�0T���I����|��rr�}�(�۬�O�N�m��%��fH��[���F�IQ:Ɨ�ү
X�T6y�5�k�i�?����T�o>��+��ۖh����-ܷ�S8v�$����<������w���9l�ow}]2��BX���ڵ��#q���ٌ�(Ս�W�"{�X]�-�5$����-�E�H��( Z�#�E��[�gF�]��,a���i8��+ٚ;�[�]�؁�r�uCm�-�D�k$f��޲c&ǥ2��{���s�A��[��%4?���B��/^<˂ꌄZ$�� |������mL�7@�*�:|Q!���~2�&U�� �JJ��M#u���6��_۪$�ܒ߽���,�6��Z*e�D=�^�x��k�9[���$�ա������N:��VT���NG���:�N�_�A��/詡)<&ՍZtPp3�$�\d��4A�G��a���&m4��k%Y���)W���zsf��S����K�W(�<�/.�e������0�F7
1e���N䪐��k=��n�^2{����:���r^E$�=�N�s�Bf���q���p8�pT�@vEZ<����p�Xc	Z7�1n=�Ϡ�eܫ N2�oσ;�ƛcH%�U�g9�vg��miи<�'��?�+;ן�������A:����uE��WH�WZ`oZ0q`B-�i�3����Y�?�B.h�x (����8�駿��g��0Bv�9�|B��%�.�e~�Ҝ�24{��a|#���Q���߲��?�@'	�s}{�`H��V��طk��5��ߛ�I���9K�B��Z�i��g�m���~��>�_~�%������lxޓ�ڏON�i�N�K��w�_'��@/�(���k���k��	7�C	0�N�,��M#d�I���*�9;�DY2�=;ο{%|�z�3º9���qA�픤��/W#�����p�R���|�7!�SH>5�*��ܟ����-��o��9�D�YIB2��M�A�X5��|���|x��U��oE��U�G�d���U��d�19j��$��β�[��F҂;;�D	�iШ�ڗ)�S�o�`ɤ�C�mC��g:ܗ��1��4��� �ۯ�>,IvϾT9W;N<(��E�l�ؗ����WC({��}��#k�3�E�X�L��o�o-K���N��+�,)�6�ٹ��)�b�Z��C�� �޷���`��Ȁ��"2�7ʁ��J�e�P��[P'#p�脵v�J!0�CkW��d�����LzEIv�v#�]5ˁ��n� %G}����c�.���-����W���"?a�����8��`5��o&w�?�	���*��׮���
v+���XP5��T���߆�����Q�����;Ad䟐[�]�H�Å�YE��䛫7�L #��v�ҠAm��Pf=�l�8��nFA�@���Y�����<<���A�.q?�; �����ˀj���nÏ�G����z�\9Ϟ�Q��1n@_���R�1V��d26&S��ٚ\Q�DR��-���9��: =���7D!��\p�wy�B��aL��; L7�S�:�؉�����(J��A]��Uޏ���W4�m�blސ�Ȥã�� Q�d�p :� @�Ю��b�F!��U��까��/3*A�K�=�\N�^yD�M�~O�D�gpg5FZ����/^3��ve_r��h�=�?��;">[���]�T�7����/�T?�rٮ��,�h��f��ʢ�2�*���
=�<���N�y�"��%yfVlkeS7�rv
襴��i��Ƀ��ad�Ǐ��eH�f�
�$m���"�N�xfc�mo� -�{}��A�[lV��Δ0�'w���|����сP�.�4hɖ�W�6�482:O���2c>�:���7��31E9�⓬&�@`-�#vU)Ϫ�β�(Ք�u�s'��ئ��	i�0R��m��:ۢ���T���vl�6�nh���W�*C��
'�<͂���n�04���� T��t9I�橒�Aɔ#�┴���l�۲�g�9���Q�,�����0�A�G�3� �b�� M�B6_�(����˼�v��Z�|��yhº٨�Yuv0ơ@�>��I�w@�@� �Ivƾ'�\C6K����ֳl�D�z�L�d��ʹ<|�lI����i�6�[����i��k��4��R�������*�D��ޢ�[�4�	�Ux>(�dv���L�����Lff�"шHE�'u�m�5,oH�B��'��Q:=I�+"l`ᄐ۷����,\^Jf�82V$�	?><a���[����7߼b0��H��"K`؂?�J�1�j��{�C�E~�V2���I �WgE��dI�c��R�z�����9o~����~�����4��ٙt�������A�����m9��
\r�y_�@ ��v�ׇ8~j�meH͙^��/sb2U�(�T�F��=��5(/���\/�4`�/��㎓y�j`[�CH��=�{���B���깍�w�/"J��;�訢ez8���,�#�%sJ�u�E	
�Z��a^��y<�I��J�Z!�%�Lƥ��)v�NӅ����R�s����V�^CL�3��gpղM�iK<���8`*i��%�Ko��WW.��t�P%󪽋]0�s�F���8�~c�RnI
*S�t�#D/�kK�Â
�egr��O&ίٜ&��k���Ǒ�Oc�hA�X�q�ˇ]>n��L��&��������GJ>�	�M�ŎN�)���򒘝i\YY��3�(Ϥ ��B��",S�<�n�X0�#�-�%i������1�'��D�4F(oz,(W!�Cr��vw���<9WĦ �"&a+EE!�ַy#��ʾ�؏��kV�~f?�K��σ۱MFE!jSa�m��\�uv$�Q�$�(�k�/$n$H�`�ke������B�,w8vzi��HA�k�s����nL(�1��}���$<G�$��'+�C@�%��x�q����"ܠݶ�;@�$�F�����hǎ�\dPp�dP*ς4w	�݇�Y�K��S��eΧ<?�y0��n�%�4%$C�/\#�2I�߲NE�﷯�a)��'�!a^�c�$t$���ں����dr���J�P�&_��AyG>�r���h�Ft^�	�O��lg~swM[���ϰ�+̯B��؏��%*,��s�}2s绛|��{M�G�N��;���\^����3t�sL�O^�pa���vs��]���2b�]'�����1���O�H�;i�='���2��v�Q����?'�j+cH�$�����rI]@F��a�����?�(�/j`QFx-k��֍+v�r�22ˋ���_~�9�=z.?|$��ʛ��.��γ��x^�|��,z�H��re$��^�)���B����CF�`���n�3h���i/B=��(�.��GW��8\P��T,"MϠiSIlz�7��8�LZ�#)'�[�����Xϖ�	?Z��g�f="���@V����R�TQ�&�nT�S�j���j'�$��ј��'$W�'�PBF��]�����ؠXM���ZgQ�R,C�$��l��� ӑ������@\5��2�}�XA9��E�@�P��\�5̇��pr���o���<�PA;�X�:���t�	u��=(?�u��JG�2���z^~�mx��פ^�s#�3�G�سf���!����5�C��~�>^������m7�Y��5��%X.��	��ԗw/۲����:�b>ǳٺ7�,jV������F����=�Խ9 �!����4��I1C�Uf���*c^����[�U����9��`ԡ�SbN����Z.Ο�W/ç�lq��͛l�-�"�lp��t���Rn�Pr��X�Z��:6r�Z�ф��>ϓc`�����ݷ߅��.���0H !8o�����uܰ�@HAQ��!����{��_ï��&������,�`�dcO�a���U�&�a��Pq�hw��^B�?	|^�
�6˖څ�}h���(�Ν"��޻�̄ALΟ|��38^y̠�h#���k��鲣w�u��~�����[rݑ��=kEHW,��jq����8\�x� 5q}Ȃ�Xi�وc!��g��pߝ�B>�\87��@d�B˨;��Ij��x����$��֮ׯ����#z̜�T	�����P$��Ѷy�%#
�=8{�k3ռV^n߷�G��X���y�[�6]��9N|�
�|�r�zC'wn���b�?#AY8g=�HD��h�`�$�������bZ�a���:�����H�S(��8�����t�����.b� �):88ʲ�5����En�������J��V��\��K����uI�ù��~�>9�@P�������D�Y�dʑt'�c�+'*�	Q�֘�պfP�4��=϶�R��!Z�A\��*rZ�Ԣ�ޢ�[Kž��5��9�Q��<�Q)x̨M/�� ��DA��w�`��������V��q����,��]�QQ��BoK@�V����vO�k��?˲�����ݫ�«o��M�@���)h@d+;9���!���{~���p��
Ċ��d���Q�� _^�g������ɩ�e�kyN�{6�Y�U�ʺ�W��GZ��`��/��Q���:o4`�K6j�ASn�T6��@t��7�^e�,��_��y��//����4Z��	�gqv3
2��a�b�uL~���Td��q�z��.�ZRO�(YH�[�O���W��A����X�v=�z�TF��od�v�.}:���t=L�/I�v��:~T��q���Й�I�=ŷ�i��̶�����y�~?ξ��x�1S��V�F��o�w���}�v��p�P���v|a��2M�Re@���1D��!�q����� �`�
�e`���8j7�R,(Ԛ�u�a�3洍Zrv�$]V'��$u��x� ��D���B	]XbӔ �)#��"��#���E� �%a��ϒe�1�*ba��@C�N�rJ�1�:jP�'ߘ���yFC�g�/<�|���T��3%�Z`_����ʔ�)��S1�ms�f�N����V�v���c�vY��jY�+u=^��i�#���&�$�>�cԠ��~"lR�M�,�I��?E^�gS�j�ޞgp��%A`�AI�Yx���L&;Gw2d`�b�Zm���C�.硰�B(�]k�3�!��7�R~9��Cgk#ق�f�M�q*G���Ѡ�zo��1�$cp�I����a�*�h7��·��q����J
�:|�wS���9C��ʸ�6���]�����}�F���L��Ǭ���xҕh��} ��ų���A���B��M/�O:G<�����=�,�([�.8Dsd�ސ<�w�H9�Q~���4������=�7W��Ex��g�@�dY���K`P�qG�t
o�>���o«��@i�{q��";�c��}y��C��c�u4˼&�Z��gcA�>�����~����'r <���C������5�ʷ�}G�g8I����
��*0�K�+�\�4m#]���#�Nݵ�5�D5ZQ ލe���׫p����N���s>���n��-x��z��IۑS�"8i��(Ϗ(� (9NPM��o��[�KJ��JX�ٞ���Z�+��л@bn �/r�� ���A�$��%3
.��}M)�w�X�u���$�+f���F	M,��ۤ�ufѳu�gk�lfm�k�d2g[	m�T�뽦��3�?��K�A�`�D�q���X�3� B�7 �(��9��4d8��8�7Bd�r>	�a)�n4�∠d�r�*�T�omIvIC�7\�ѭXg�׷ٹ]с�3G��V%pOʃ��dؘ(il�CdI�= /k��>��zqq8wdO�NÏ��#P�6��t R���Nd0dU��&v����]�>�M�4 �40��4�ܩu�7�̓)�Y�䶄�K�Jb�oyY 9hw�u��^��F��v+�#w�<]��ēnc�[�h��uD�-1:X�)E6�me���}vdd�d��q�����7�-ˁ���(��p��A�! A.4��dt<��Oj�;G�g��L����s25����X��&m�(�㵝f?
I�S$��d�Q���#A�KSh
�M7BR�}n��=�;
K d��x$|6(�e��}>�����u�D�!)�c;$��w��Դ���L6�!K���ǂ\Ú�_I��
��$�5��2s���h�2�g�XP=T�W�*ojYh�o��fG>��g?�v|��?�J;�Y��z}�4��1��±�s�#T��[%t��Ӕ�&��fOi�T6����ˬ��?t�8I^U�ߏj�E�����3<;{F���NJ
́BY	<��F�%�r'/Y���M9`�o~{C��O?�k�]�?�,dqn
��;�%P�A�3c%B4�!h}g��G�����������C��x�0�1�����|����3P�l0��&h��2G��)%^�⤍���v���E��s[q��=k���}��3�f�����Iy3}~&�w�[���ry�@�����3a���5V�g}�S�~몊 ���?��K�����4\t?o�)v]u0�6���UW=s����X��8���-Y�dKqtW��A�6]���6fS($�I��I$��(<8l�L���臕���N�i��w*Ї��Ͽ��o�3����	�l�h-��y���ƈ�G��)�nk�u��ҝH���*��6FZ=�d�HY�tȥ���a
��������Oe���#<?����$���r�~5�/F�k���>X���U�w�2�?d��&w��F��%�����h,"H#�9`b�t���%�o�['_��V�}�NW���x��S���䵱sG�g 0��.h4ݰ�lO� ��d��}�x���	�W�^q����J���������C��<Aj2��f�a��F�u �.�ۛk)%|�����[���q��[G�,��CY��q~ d�ﯿ��@J�-���'f�Wk!O�'���5;6[��-�,��x�ۓ��?�����Y�������g���\lU�.d\cy�=�)#Lb=a>�ly����p���*�Z8�	�:���+�OWYG���@<ڳSO���8)�ZT�0�{V���Z��M����@�I�U�Q�N;�̠��i��!B�dvp;h�?�&��$	�� �t^��b�x�����~w�?���N}[�����;�r��gIe�9��B��J��Q�\4�.�N���aLQI���cx�MVRi�|t&%��%�铷7+Ȯʬ����+K����h�פX(�'�29[�^��2����o�L$�R�C��� MEÀ
�|�-��54��J:�J �Q����?�/*����p�= �J$�ta%bP;�.7�sl��b�(UN��;��N[Y�����(	�,\k��%r��������ijT�^��a������v6Y@��5T()�4�6Q� F�;���Ygl�+��Qj�%-%�uJ�&ll֭��F--�=`�@�*RJ��zo���z6�x6�l���Χ���_d���[�2��j�$
Of?�ק�6�^ ��E�������[�g�
H[<K�K\t~��x�F�F��|��p�}|��5����u$���=���ۯ��g�%���鄫h�m �S��
�;D�Ӌ$Ʀ�7�����6�_j%A�R_E�cLO��!�zvȧ[蹻�~��گ����t�0�w�5ɌQ(�e�L�"��|��J��~�;=�ħq!'�����^��=[�_���G��W�ڦB9V�S�������y&�r-�x�p�`=i�]h��82�ߑZ��~�F�fA	8!��A���d�dz}>8�B��0���f2~=� )��:��~�dD��!����E�C!"�ae�K���e+�������ex��g�aX�Շ�4ܱ,P���y' r��£�$a�q�P���Xji{]3����VJ���4T�My��1�=s�&ĝ�Vπ�=�n���-�7�㗶��c�bA�o~ݓ��\�G�ՠp�B.64E��-c�n)���1���?�]\}^�N�;��6�XH`z'��M,ı�"̊�m�2D�fjx6Z�U�{ްV�M�K妲5�HT���]=��1#x '�Us��!Sz�00�e+\/�Z��������s��ᠯ6��\��n���c�����e����R*��P��I�^�q���^dʞ����a�2�ec����u6J��iޗ]�;M�g��u>�x�d���#�� ��6N&��j��YHI����i<�g��E����٩�	�8l5�S�"��9&��QA� ��C� |7�`�.I>z@4�y6̤���`�]C�鍶J罠cW>'��0�lN��7�Hွy�;;v�ȆяkCV�=��]�0@���!��2*��&�EdSy��Gp<�/_2�od����=�L�NS5i�F��c�Ao���km��&Vrtd�1g�� ܱ.�}��-� ��c Z'g��ǂNr��s�Y�=�����:�}0��ְ@d�v`��l'�I�K>G�Ϣ�$(7�讎��! �����r��<�sV��١����1��N(ɛ�{N�g�w��)ȓ��~�fo��7eVL�*,c�����q~�+�K�9 �X�ҠcO��0�\i-�HF�"�IRq*�[CF��T��xɇź$�e`���v���>����^��3h�1�9�{vZ��H�8��h����-�������xa�V�k-�B@ƨ�y@`@le�E�`&���r@�觛�������Z��G�IPw���|Q���k�L&;�T�]�?l���>��P��3n�>H!T�٣s/ڽ�-�3���y�����q�RE}�IP��)Z2���+AtOD�\��:���dҎ�� ����J�@Ωd���1��U���w0��\�Al0$�Q� �E�N��8��@�QI�9���eD�X��۲OzK����������D�{��\B�h�wo�Va�Bh�6T����.�sH���1�I@� �YW�?��ͧG���gY� ��r��I*�q�p)�yR�ׄ
��3��?*xFZA!�V@D�Q��^S.� p������^�H�l���p��� �����p��9!؉�5�9z	tI�J�@|?��5��P��"Eg�����}�X=�n,�~"��陻)�L7[H>�CI�K�o���Iի����:k������8G�?{��uv�s
�O����gN[�FRE�e��M^ ����tN"J�녁��!)#�8��(xE�A !��R�ù�a\�����c<ޭ�6~�	�50Pc]�իNj����Y�E�
�������0�q��h�&���bזA��8���K�7&︓l��0x�9�ɍ�vVR�*N�l���DZ�/�
��r>{t��k�}=/�&���:��0qn�� �D|�62#�7��2�l�?�5MG�k�C10�����,x��������Pa��Q.(�W� ��������	g�m��4�hCX���t�(�=#h�+8�wY	.;Q����>5��O
0lD��xE�>;d4�묘:s�:�d���T~��֛�,ao�0�H�7�_Cm0���3$N�q��D%�窑kO�w�MוfL�2|�[���6Ui�ڨ�F�Xg٘�%׷wB�����H��>���������}�W������nG���2u��~�Q)�A;,�0&���yx�LH1O�̄�o����0��HbKps+�Qʸh0�5(�E�܂���w:%�L�`�@�Bb\'�'	s�����`��ĵ�c"�0�0A�������'�5�� <Ƽ�R869qb�:��xX�s�Q�.�Z$2^�:�Ϭ�޿{���SORt$���@(C�h)�S��S��&.�z�_1z;z#P�Уj�N�J;�4�.0HKs$Qp����n�)����h"����bq�|\<�ߨrL���}B�N^U��:)�}%l���u��N�t����S���_c	e$�G#�b�=p5�m$гφ�4@�W����.�f6�!�BA��I�M��1����Tm�]�a��k��\�Ϝ�8�&fa�S]�C?������~���Q��B�rN����fd�H �Wu~Z�L�aX7���<'V�K 2;�K!^��F��n
��j[u,�W��.*��I�OIp��� m��x]ﳓ|}��hl�2�����������N�
���^�7\�]�&�_��@�[;����j�,�޳�b����:��q�5Q<��ꅖ��i�d'#`�: ���� ��k�hw.JF��i-c���P*�P���*���&�d:ë�q�\������$h��cfY)�'����ŧ/v�D29J"���`�DA�TP�bC�f���Dur#D���YQ�X3�FK���D	�����	I�TD`*J�d����	}2�C�x�\��S�������޼�-����"m�v�G*�+[B	���H�@�!oo��E��K�p���=mT6���X#��r��xA�{x|Ƞ"�Ju�718UB~+��z��S���l�����(��^�m�R�; u�����p�HB�-�ɥ������e��ϣIx���.�����!�E�[���.l��i�R	d�����;s�|Ŗ�A�sxzX/��y���437(W���c[�������S�]��a���	��b�l+���� q"j�7B�u�9���(���pc��FH����c����(h�FB�W�GFR��'L��zu,G#�;Ʊc�!C*��R�������T3���sĞ��]9�Q)Χ�֌+'��� �r���vf��5J�ւAU������w��y��a��U"�p=U�MM���ȫԦJڃ.�mA�'���&v?�Ւ2{;�l���w��v|��q�c�!�n@GG�XM53�
����gn��8i������լ��ܱE&���N�3�ِ�3� B�u�4Q�� ���K���%ɕ}�kB=B|�N%��L�;i��p7P��em�fD�;�X��hY�j-���Y�V憭�1U�N��}����pz|�y�M���Wf�`�a�`@���֡�ۗ"\IU��A�>����ϟS�aI�b�N<��A7���%+�� P�Tq��������*��Q��*;-�&�� P0躅����yC���������W��)y 0��2r_�[]]���ka�d�����=�x��"�?΅�z`V�^��VDŸ!p���[�K���(�:qt��1)a6^7	�������JʄQ�%�*]%�CԢS�b#�Ü-�Njt���'�0ñ[:�Vu\�q����Ed�^�H�2�Bh;e8ƣ�QjB�sF-U5(�0,��6z<#o�@�$ ��U��Lu���5�C����B*N������Zrk�?%�B�e�f��D�m���L�?��ٖ�w��|�2��!�� v^@=ߠ�~T�D�N�_��$�#��BXj�va
Kk���r�J�6�S߱e���63�cыelΧ�bFu\T���r(�Y�a�߭m�%2��QU��������.D�����z	vBnQ1א�vZy�����y+;m����WR��d�h]��|�F��{Iʰ���k2W���=ʰ�4jJᵠ�ʼ嘅�3��H��f�<��>�qK�ٯr�G���>YV�֨,0;DI�Yr�G��%��6D `d�y��o�B����/D�5z5�ǳؠĿ�~��A���U5��e���i���J���|M�Hf��(��# WՈ �$�r8B{�=I�D��_[�d��S�%$ #>M_���5���A����'Hw�n�-��%<H��k$>���><���c�|��W�ZK�26隸���^��E��J�E�b�UY|{�u��T�҅��<�H��Q��t��MBp��V�C����jO�6-�:��EOu�w������#_�Tv�Ӄ˽���u����:���FV:Sd�񛪔YA:��������f�)��4��:9f�s�g�m�ؤ�b�E���_������)KFo�L �l�h��Pt�(P�u/D��Yܨ��d��=kE�F�f�xH555�ƀ��� �O5a$���Qʘbi����v*�!�;��΍�^	�s��'��h�������F�lw���23%h�n�s�Y�:(��P9SF,6��Pϫ<)���/�$��Z%_�yِ!�Bq����V ���܄��m~��#(;f7a桄��L��b��ޯ���+���9*ג����:�]ۖ̓�XY��fJz�R/� ��
���Rm�p�kdӂ�'q̏�a���5�\KMf��ÂS0Ġ5xzϬ!�Ch\~�$���7o��o�HF�]�ϧ�Ny������y^�:;^�k���ہ�֜А��3�C�`��_~�)����?�۷oH\~��.�`>_�B�6���aD��e� ��cㅱC�����	��&�(�"*M���hϪ� Ĉ��@<��נ	 �Q jeN�ZtE����s/�!i���gn��C���	
-�Y���h���u���o~ci�J�>^JW��D��ɫ!%�A(�����������)����/�H3H�6j�J���6+���g>��;%衖�u
.�����Kٯk����R����(�[M~� T8��r�YR����2�9y�^#mL�Ӯ�:�H*,dI�Cpn�ƻ�)R�i��Gu0׽���(d�@V�Y�@fA�`���p�X�W=���j/_?hi�MҸ%�'��Z�W��l�h�N�u0�i$���-�~��R9���G���q�{��'�$�몛��%2��y]�ڶkt���-sO�)ߢ�~S����KG@<Stp��6�K��t�����%{wjo��d�o�ɤԧ�}�S)WD��>/��:eWVob$�V'��V�E��!��D]OUp��qT�fd���6[�(��(��?d;�-�R�i�k�ڇ}Ib˲X�ѮM(�)���$�q�Q�A��~�����ݗx(�8�ӏA@N�bO���l���0:rp�|A�\P{/��������γ.9gb��OWW1��]*���Tv'�0}�+��ʾ�tk�.fkG�-NHB9/�"i/��Ř����t,|����1��rΌ��6��m��߸��N��T(��(��K�;�$10~��D�/��/�Y�'�[�=p	g�-�C��_^�D;I sP�݂Nm�
^ī�
P�����{��-��cW>'����FI�\�����;��另3,��i��9f��� ~���Û��W:w;w6]�|>;�I�p^P�(�W�^���3���O��s埾�m�un\P�y���<����d:�b-|툚���R�c2�	=4���;��W�+�aQ���m'�߉�_v	8�����K�~�O��V��eg7�v�F�5ݵ�P��ȮQ
Y��ߌ]Թ0�\jX{7��!n��,I"��Uȡ���B��S�,KF<�D�Kz|.Ų��5d�c���zr2S`n��BQC�E�`�b���4Hw�NQz�ڈ��Q��ݏ�:�J�G��Y�%�#��ֶ�$v�ij����TڵM�-�v���UU9����e�i
b�F�48��/�q���G�Ltp�|�*��\��T�4���&]ON_�'@U��=�0� B4
J�-ECQH@��8�d�����.��� h�M���;��/�'���O���t�X��~�]Z��*��Pu^�Q�Z���Z��F�F�>G��
�Ƃ?`!�0�Ȳַ��@m�ӴwYP�����c�ɖ��*S��Iu���<t?C�����e�K1�����lP����X���|�wR�)���JҒ�2�(�����l؂3Y�Ţ��	�d��ǘJ97�IDd�7��T(ߍ���Lx���72�
]���Ї��.ܵ�D���6�����z}��ݫ!'�(- BA dP��@$Q�i��Bk�6_�q�H ��AI|Ij,�)�X�o�(�R�kD����Xe�RyF�\�/��Y����J m:�`]T��0CA�ٺw���:БCl=����{�9���DPW�aib��Ak���d(Aם��]��lIE[%�(����H��y~�Ԁ��l�YQ.�&T��PZ�Γ��a�n��g��,����GgcC�P�GYɉ�gK�����"��t�]�>�0�Pq�3N����|��z��2��N����^�L�Q�+����sY��K�')��M��s�Y	��rjg�:�$�.���k�NA����]/�a�;�`��Mԇ�Dqd����8�x�"|��>GY�ҭ�����~Ar���'X�JI��2o�])��r/#I�����n�����_��~/�g��c�H������'H�G-@�@j���#~D��7�ف�u"�r{w#�$�1Y�/ӽ�ܜL��cäC�~�}E����T�F�b��<A/Y 9:���v��X����,�������L~�,y��]����)s5��1D">��y�u����2вZ�f�����Ko����T���.&��e*�+�[�R� s.*ɴ!����A=�ФF�\�P�:v�B���3��AP�	�u�P\�]�0�����6� W7�H]]]rN��H����m��3��F=	��ֻ�<�$�TZ�<E��x���w���HT9�gI��S��9� ����2�.�XUE��p��]�B��m�D�g�6�5j���a0�m�a�>�������j]a+�tepD��˻�ή'�6˘|q"^�H�:��,�m%Y}��c��Щ�k�zG.߭��_'�4�I������T}o�S���{�!ΎE�'�������D�t�nW��U��f�r*��F�ӬL?N�!�9ʽ�b��bHy��٭��bJ�o�J*��?��tq�e�٫�h��/�$�K�Q���ڻ�19��0�:\�z͸e=<��a"5���:ѹu�v�[g׊hϸ��Y���+�S����,)c��F�q��T�vMVX75k��ٴ� ��-�۱����=ݜ�Z�s3
aw�T�zYU����s�V
`�[��$D���ŋ���2��m�_�R!E�r߱���j�UaY�2*P�t���	����H���H @v!#İ_x��)�E�CC��_��Q�	o�x@��+f�4xE8�F�V�CK�Pڙ6��Q�|�������%[e��;�U��tp���TG5Q]�0S:�.��	�;�:6>n,��v����e����ɴX�Z]V�T٬�)ꒆ��յ;?|�Yf�H�aݓ����3�Z��i�N����ֺjZ����n�c��ؿS�N���ѡ��LBI/�"�Q|�WY���Z��M�uDD}�����e�:��D��I� ��$��Sd
Y��ρ1^Ҹ��h3��U�ɉ�K�Ni���H]A�b���\sF�;5DN�e~Me�괘\��qqnGG���ɟє�c,�=�^u'k`�>�$0=N޳e��ɟ�ݫ���2�����jY&*��P���ޭ·#:��ϐ��Iv��XY�`N`�V�Bu���[�z� c#7�ʪQ����6�ܜ;��s�%u�k��%�q6��!Z��D������h}^�C-�G���xQǶ&돊���(9r��KZ����d��]!��Oi�n���a4y[����5 �2���O4��X=9��K2.8:��_�j�^\r���÷�}~��/�cq=�[.��|Y���<�6(AF��B&�9��woߑ���s#JDq,��[ 4��?|����������Z.KrfEU�p�!�ة���>'@�k�%/Z�J��?�+�o:����|� nG�;oIS�o�+��ceM��ZV�-Z���$B-!t0�C�@���"���z�bg�5KoQ7h�A-�����O+�딯�|4�X.�z�d-7@�@�b^�*\��Xj���3~A��;��ʄ�A0�k��<s>�JG�m�aO,J�#�Ɋs㚥ˢ Y����d�͑�A���+:�Ӯvza�k��J���Kx���؍��x(��,/O�W�x1��bYq>���ixyq�m���xA���p����3�f�X�1��!��އy�^�����lC����(���I�K��h"1��N۪#�K�~���"j�Ԩ}0�J,6�g#M��S.�Qڽ�b,j��&2PPƁɞ�	�}�� vꈖ!B��U�O<��]ԯ�nU�B��CMbi�Z�b�O���&�U	���w�j�Yw+�b��ޡ��o�L�iA�z�V-�E4٘��x���ޏt%`�[�X��x��j[wU=��Ǳ�ɇ��w�ʹ��-D�>�:���%وZP̾�X��5ɕ�A5��Z�,���F�7�G-<��:r3.�P�'����3�ω8���ݞYS�����'Ҋ1]e�Ä��Zl�sp>]�����O���M�Z�[�ڄ{e�O2V���_�����f&b=�J��Pv�Q�nV�T�p��;� �����cD����̡����#��@h�"x0�vs�r�\��Rzdphi���uP�ؘ�]Jy�{[�^��b��;�NI�4�c&��W�r2E%&�F��P�u������d�� �g�c#�D[ +��}�5R���04�"b�f�`h������qm�0�>��='.�g�K 5��^}���XKq<S@�I,y�$2d'(�j�4O����8Щџ�#;ǻkKV����`h�^��_)_Z�3]ŀ�vd�m�1��1ONN���r/���{ІA$�a����;c� �&��$�j���"ܒ_s�/�k&��u�ڄ�0hK��k\�kr�1Aa����Tg���I_C�4�-E�*MvH�I&P\�$�鷢�*lN��۽��R����rzG���4Vv��Z�T�NK-m+��[s����@G�.�p���:�Ԅ�ub�~��9o���a����&�y`g�����l��i�Ln���]�ߜ��<Q���&�@�U.�a���S\�@a��IA��)�F�>4����	v+&�d��ͬ�9�$��k5J�;�p��d�2��"��X�$<tƍ��ы��e��i�Au&�#:���@��6����� m�E�ݝv����0Q��z`��m�5��rTۮe�wC�d%I���fɃ��
e2缮���+oJ��q��ǂf����]�W.���2Rb;��ͩk�x��Ґ|\�T�s�d�ʨ	�F(J�+��c�?�$j�P�q��AQ@�h�0�'�|7�z�LJ�B��6�#
�����s�M ���by?<���#�;-�b��M?�.�G��H5B����+0ܦ�b,��&�$2JIZ���]<�v�n�s��H�l���v�0��G���D
!�޽��2o��s��b���ێ��|�s�{����j���]$w������y�wu�銼:}��(��J�RA��krEfjo^-0q���1D��k�/�l�T��s<��n�D^�]Ρi�X�^��S��w�2�\D��=��v��i[qdk��ԯ���I���'���V�94M2�5��no�v��,��"b���m��ݒ��;2>�|���������磊�k@3���/�El���.X��3[���J����S����強;7�/������עbD�6{�{������f���#i���u^?`���O�R������7�.)��H�H�Bd
�<�4�����:�}_Jzbu#�}�d(Mc�"~�v�U�#��wh#M�?�KKQm�ީ�Me�L���Љ+ȨY�3Lh�%���ef��A��lp�U����Pi���ކ�we*�ɤ*cS;��K�!�V�kߌY�%�a��*�n�_c��X,IP,�3��,o޼���mQ7�u�|D�FN/�l9S�Ύ7P��$k�A۸����lC	������aw59V��W%a��[���=9k��^zC�a]xq0���t}�#I�[�N��-*ϫA;A��t�Pb�r,�K�{]Iv��9�𹵗I��L0aHsM��Q�O�G�FFs�\!�FGd�כ������W�	\��VA�������9sR�ո"\��$Ư�r� ��'�/�4s��_o5�L���4���J��M��ڸ���W�uvG�+lC�g��.vƃg���\^V�3����z�ϖl��mG@H���g��+��ē��uz�<q��ʗ]���0I	چ
��I��-�{�9x��X�}Lmw'�N���*�rWY��тcXg.ȧ��r��($#)_����B��ul?�H6ۇ�,+Q
�vӝ�CJ8�9�R�DS���P�I��P,U�^:S�%�;CkZ��S��_��3�5�]g�������[�=t,�:o8⾝�����Q�D�6,� ��+A �)|�D�2`�'��+	�s��US����xe�#�b��WA��Pб�0?$H��`8
�|�A�.���U��Q��λ����<�[������(��-�k#�:��yà	��H�Z���X��Ey�M2y��TU�.���g�n�9?\��4�.-���^��Ҩ�lGr�,?"�9�w7ԛ�ߘ�+���v;��w���-;jW6& ��fW��=�3���<����	:�?��?��k���<?(���7���o_	B)?�_��%�(�J"$�68Ǟ�/Ӵ�F��+C;�]h�d�Ϊ�;U�+U��(F��x��=�_� �vvL�6C���"��6W�c=��P��:iu���M�^_��w����X[NzH�#�3	A��ф���H�r�i�	�n���~M���c쌺��X�z��q��h0��1���%��6njз��
lݜ �T�D�B�\!}�U����&�zp�n
�M~�OB�zl�ֱ�Y�籘�����&��}/�£%�x�`��8�.�M˪��S�@�z��D��d�������~U��w�A�M!��B'�'f��rA]���g��2`FBkF3�V[��A�]"yN=$D�����,JI��P�44�`a�����B*���yR�e��τ��:��A�����˘��K�2�לM3�i;u"��^m�U6lZ%�q��w��C�A;	zd��cT��*�3W��!@� �F�]��3��d����v�rH�-��ڔ���jGh�)�K�{4���Ϗ-y{_����H�2�A�'�]����	�s�$XG��6��`�<hKv�6��l�����h�sj�Ts؀�^��1�aȲ���߇X�n�p�<���X毡]��0h�m#�&�q*ݓ��#T��;V�[f�N	����g�j��!��+�q��T�� z�ϙK��g��.�ڒ�t�˻"C��oI�l��cuQw�� i��R_.���"��;�0�ʔMJԓ$N?+_/:uz�}�:3���|�Vl�Ɠts�Ԗ��gȣ��P2�r�E��7��VS+�7eX��>�q w��j!N�LK���܃�!|���,��"X����>��DY�Q.\��kCi	�Qd#@��P�	��RFEt!�QZ4f��P�,�Y(��S���9����Y���KY#H��e��m����]эd^1�X�g����<�u]E�(5B����D�3���xH}F��`��T|/U�UM�B�P���I�m2 �u�+2􃎳�oxN@��Dm�Rٹ)�>Di�n�3��҅��a��I�{��Dt������1�$�1M�:��!--��+9M��Ji�u���/2�|rE������WA\�5��XP�M�&�tZ���a����9(/�0M���XX$��u�NPΤQ���!�s��<<q~����)�����^�u�������{1d�ڈ䊲R��n�C�+��׉�ڒ��N[��蟷���n,���a�Z?����li_��
��^��'��?,9}U��'oiǽ}���c�Qb���(�)u�:-b�
������bh>܉O�]��1��e'�x�&צ�f疤~��&��~��A� >t|�y�$��(�&�w�����z�btR7Q������9`�xͱC���|�ī����c����S���i2g���0Q�r>� "T�}_�YV�� �NZXZi	�uNR�7�[d�k��FI�,{��Ғ�(��,���;nH�&�2KM��\[R�XE��fٺԺ�Ag?.H�k|�+Re�%8P�v�c��b���D�ip23Wqd Ǹ7�pnc�M�Ӏ��;�[�e`�J����Y�<_G%V��<N'@�A��8�F�u�@��e�����Nz���t�]��g���&��x	.Z����A\��ѐffR�m���`� ���xM�	ɹt{G�A;�,#赖l�x�+�_����
Ad���"��Kv�����ݷ߱���|N��:�G�5�y����:����� �EE�\�s����>����f�u��:<<	���ㆀ����m�S'�gҕI	�J�����k����6/Ryx�/6v�Q/E�-�����?B-?/E��\���T������f���x��k�)�r+���f�U6�i�����P�6} �	�����`� �eJ��y\&~��w�v,��X��~��Ow�ɯq����8{�O�v���{��w��>� 2Y���0�� X(H�d7�;֞�Jd�g�<H"�[EZ�gP�����5]]P��h�̏�~��<a�!D�`�fY��&<ܭ��ev&?~$�� :S�M����f��7�V�1�=� ���I���\7wl���W�ο�^���4��fu$J��l+d}��(�H��!��5�������ڬ���[����ߞ�c	���堉���3���NuP�8�d���H�n�T�@@�2X>A���Nc���u��D(����=��k��yU/Ą���mR^6R����b��DK ��7�f9��4-�/C��ϩ�еeED_rIy|��6�"���Y��F��r����T����<�"F�6���>�����캊�
����&��;7�co�H$��G�KXX�"�zh��N��5a��f�fE�����{��(�Y�o^�G�/:���ۯ���N���^�w�W�����/**�^~��ܚ,E��÷]*~�n��fݪv��붴�/M7>4�����u�?y�'�9�%"^י�n(���]Q��:�O��q�ۓ ��R}ȝFf��Կn��~�*�e�Z�ׄ���P�s�ag�Xښb�d y���&��Q:�m߮uvu���p�e�� 4�����r��i%L:ӓ��#�~��2_�{UF<���q,��]%Fƨ��F��k��!�6�^O¶+��Qʞ�26W�y&��8�� ��0��`D� �,���1��f�,�tU� �h�up(�\[�d'�	��ع3�8c�G��O�*x�ׅ!����ut�h�쒴�ГI���([ +#S���?[����@��a��3E�\r$�C˳Rv��"��C�!�r�����l���aPR�>�Q�7��2��m��=�r��t=��uG1E��^m,�������C~��{��ۀ�hђ����ć��OU�Ϡ�Q���P_�B�Òh8
y��C����)2I=5�]�_�����i��GZ�o�N�$s\?���x��
"�E�A{N�ӆ�E�̣���'�p�^^C:m6�C���ƛ;�O�����C;?��6j�;n��Ǿfrhߞ{"3{ޮ?�����(�s��d�7����R�N���e�A�?c56���g�eu�*?����9d��iA�'a�F�2�����d�ӨBG��"���*�m��p��9�� L	�e�kcz�Dc	�T��SjH�d�.Q�J�حG߭�kԎ��G��Ƀ�d1d,Jy��$v5^�KAˏ[�Y9�mS�ȍ&Z��x�#�I���3ؑ d)�44,�K�We���#+A��妡�4`-��e%6�|]�
�w���Hyi��Մ�d)��=9^��[�J��w2O�Q<)�7�'5��</J;�����Sb�I�F,��c�qQ�AJ��_t/�D���DX��|�l�D�/�=K��!��$�V%:�Ն����Ԅ�	��\@��ن�.N�7(
6H�TZ`�u(��Q�?�4-b�U[$��P���o1�ynT�C���l����^���k�*GP��>�B��t��,�;;=��,e���69+���5��B�HI�����Q�񇿰�z}��Z<�����v��2���!|�� ���qC/'�U��~���F�gS݊م�M�j�
�L>�tj��~����}���^����}���ʾ�������m�V��;�>�HS�ϸ�/z���l1x<gب;\�j1Ԓ?���
�V�����2O$�*cb��cB��q�8TF���5�Q/T�6��\�ŉ�%Y���*��^-���}��rwn�S��!X�*(ܳ�9����~ͬH��B}��k۞:nX�!�N�(��i_��o>��ܱ,e���(�:ȅ����xN��{�P�����!(n��т���Ĺ�h��hmU�l��o��؆�i�K;C<;c�!Ƴb��9�xB=5��`P����Z�eG�CC�l>l0�VQ24�U��80#�H�[�m:����'B�K���C�
猷�V��s7&E����������U��ɘ�l�b���iw�c=X���O�������2�� �Fy�p]�j�!�s~=��(]�g#)_G_ X�Xi]1.ۡ�`�ɪ��
3���6K7���[�0gb��3�v�"
g#m^�	0�N�bD�������e��Ƒs/@����=�����&����E��Et.A;\t�A��>�?���	7��\3�O�w�Y�V����nA��kٺf��>xT��:Tm��߅숟3<�u��6;��p�*�����(��o[!!_t\��0	Jה^g�t��yJ��lñ1�ױѠ�Ӈ߃_|�6WfZ)��\��u�x������0*�LJ$w*M�I[f��:x�q��Z<�?F�*��́o� �;)ٲ�0�bP=b�;��G[�]}۱j�!ǲ8��阆�mh��H8i%c�p��	z�_�;���dC�.���#��eA�����βf�C"�df����9o�K,��`W$���0�����D3����w�G����|�`�ʫ��x0,�b�j"�@ؼRG|.�� qt'�C�$��r��&3*%˅�޿�V���j-�3�9J`]�#�p�d@$�F�X�;00��k"� ׶���l(�^l�AeQ8��7���7�?N#�<���~����@{N�;���C,Z�`��ƥ�Z�F:�9�Ϫ�g�$��q��'�w����>�>�z|>@	g}h�Q�������o�= �p���x��ŷ���	��k��sӀ���	?�H�P�qM6�������_�c#�t����m�͟.Û<߽y#A' �0W�)tjQ��%m�,�Dh��
��ws��x��/h��g�V�j�T/�C�յT>��J�\P闬�8��ke�o$L���u[[����g��s�x�
�qǹ��Y����wv]P���:��Ug���ԙ��Kp���oU*l��~���~�ύ�n���N8��[���!�%���'�y�)���1�D�e��2�V���ٞ	[Hf���7�]
��nX���2V�"H�B��=Nr_p��OeJ5r!��3��k>�}��s�� }z찡�Me,v]wy~Z�ϊ��L�4eyD!� R+�}��,�<��q��89gҹ�9m��6�c��ܦ*�Sd�@Ĺ��/|���|��b,wf7��I`������\X�I�)w���0Gj���(����Fy�n-���!�t��	6��PX�F	iT���:�A�"��a�s^Sv�����ׯ�|Ѷ���^+�EI:���8��-t.ID�����yT�s�i�U�L��9���a����1�gV�M�4W;�B�k��$���|?��c ���j�Ǽ�ϯ����M�`G#���֌���Z�3��s�$�������P���.�F/b4n�ٹ�U�=�p����>���O�;8;��3��tC#c��zX��$� ��l�5p��*d��H{vz�k��q|v��A�~�t)�R8�Ţ�?�}y ��Ad���=!T���2�ꐜ9-9�r���߇ш��ŋ���;� ���R�?�dl�״�Z�_�{\�I6BW�V;�(:)ENDgQ�E��dt ���<�z����P�r�����i�߱R��p�R�>��6�7>�����8�B
��<h����G�3e���d�t�4 x���2�֐��p�1H`����Y#s�����3�0y��ލe�Z̛4L��n���m7M���w�y�a<b��(m7bp��]S��d
�l:��&�L%�>f9=^�*�cC�I�A'wP�TRW��u������F�~��~_V:.ey�൰�*�(�L�k����PЕc�R8v9:]��4X���vRA!��xW'-3�nW�g��!XAr�|�8���	�R��?�ί������.C�?����J9�准�%�-��N��ۮ$H��#W�f�:�i�Dk��b�ƞ��c�e�:$�4�פ�_�Q��)�1j�����a�����oNl��I/�Yk`G�_tiA��%���@[R��tm;В�LR<�1��}tz��ć'�׆ 	����n���D�
d�,i��"i�|�F����*����U�N�+c�?;��Ckqg72�2o�{�N���<�x�ݿ�C���>���R곬�VJaY�=&��e~�_j��ܯ����8>:�OI���+2v*��ˁ�A����U�E���;����1:�6�V3��l"�A����JER&���-$��������t����ReW��w��]�c�[��]�&Y���A�c�F~�Ќ��K�O�s	P�t�&B&�p)V��n�&eM��K���]���W�b�9Ru5%R�̱���3X��5��[+�9�àDh�6��O}3h,j�yqP��6k�\�K��w�s���#����\�{r��o�#qqq��γ`��ʠ�V!���Oc��쌠�|Y�@���/�)H����a�~m�\�#zB�jR.��3>��$6��L�8	�LS��5�$��4�'����#�Զ+v����ƙO���M1����9G�La��~2����ݙ�g��]Ԇz]�m�fo�L_���]�d��!A��F�z��o�̵�H�#���T��؃��A�dD�G��pJ�E�@|���Ӭ��?{.�wktH����,���1 ��Jf�j�)ڶ@�{f����A�
��ǀ$�(�YKg���2\d#�~$��w��vW]+	�H'��<�4:�ݮ����PQH��!Q9�E�.XXKk��(���R#�|:I`��,��:�w���uҁ:���^�s��c'A��po�옶ҙ�
�� 8�w2?���9+�3�C�`�ځ�S��Z;���9ò9�Ûi�%j� �.[�,�ͽV��5�b���������'b����=�G�!˗?��oW�+�%�l ���l�-A֙_����X<�Ɲ��=�����Rj�#]8��_I�/�8#+'N�،�pyĀ��@~�0�3�:8^ӑ:ȿoz2s>��ρ��ԁLG)J>]��T�~�������v3ۉ�'�SrG���M�_J�p|��m�J�$I���b:���&^hm�D��?,hP�S7F��	�!�Z��N]��Z�}X8�&��Z���mF���á�4��m�%�/_fg$;$�Gٱ=8��B�B�
�����P��)p�Fv�k	��W���k�-�ܣ�kI[AI';k˾Ϩ�v?���ԉ�Z��:�<�=���yw�_锳�����&�ӋyTl=^h􆲖H8q����F�x�؋֍F.ʻ�j/J[�F���I,�\����wԆ8��(@ʍ�C�]�.���8[�o�Q�-�c�x�rEDQ� E���y��,c��O�D����kᤁ<���|9:>��hEAN��]�Z�R�*rV�V{���hMGX��x��i�A�~�`����_���������oD������ԝƓ�sW�54@q,�^���[��gϒ:>N{g2{A� ���qӔ���tX��Bk���r���V��#�ZR����q�oCBs��oqgH�,�a�������+|�CB�Pn�27�U������dh᎝�:_�k���9bΩ�|�Y�!����!�T ��~}��r�g�7Bo���aw˵����a6���>���m����I���������_�k~����FZ��Vʬ�x�q�D�B����o�[�Iػ��p��|�\P;X�@(s=G�й���쏉�<^G��p-Fs�����v�1��㇏D�d݌Գ-y 1~g����_$s^��TT�[�k��u�	��S��<f�OSe�+X_��X�^׉�\��
7z�PwL�a�*~|}��ˏ�+�8�g��=��%}.��gl鑿�?O�R8ɊA4�m��d+A��@_x�'�>�-#�I��5�vm�Fh�zҕ}�q�oBw�-6���LU����i�{����⓻�eM�3� AY"���7�Js�d5���j
�'yAԘÙ�.w'��fW�N:�JVa����]���SqB�#�c�0��;�#��i
��(#��:%�6���[��>��ZFU�;�\�ͺKP#���nk��Z~�(���*G�b��|yf4��,���D�Ǐ_���k���6����U�t��N~�R��ƾ�ty��Q[0�I���d��1�/�p D��*D�0TRp�`��^f1̤�	�e�La��~v�ٷlQ�d�z����yiΑ�p�|�QG预�ڛSgc2����8��O���SE=1 �>�;�H����YR.���Y�Y���<㶹i�р)qs(�ݢ�6�l���³i-��(����˜YP�3� ��1�|y#��m#ϰ��7�x�<\�t	C�Q�e-h['��\W�B��"�t��O�2��8�1F�+uJر#��r#(��?��fF��;Fi���WqN�i�b ����.����2���(脓�E <�� ��]�@�ȀJ�������Z�1 צc���/I���˗���s87�ِ����ɩ }`<�;������n]���d���H׉�8/�	u@�9��y~��N�����,jP�ei�W�X�k��[��{إc	�l��T�H���(��~��!+T�/<;�^�
?����ͫo�������͛���[�����ub�!:A�ب�Su*Sv��c�+�힙t��4��,�����ޯ>�nz���dn��E�ﻇǟn�"d��1T�:�D�9?��ׯ���|���?G��?{o��8�$	� �~ŝGMu�������������k��2+�?y ���f I?"<#�{�w'A;TEEE�n��><	�G�MN�����f}@�������k��M��n`�TU���Q�6Ӳ��?(2@]��ki��wO��
�%Z�+7,��ʘ�z(6 	��IVQ�R/�Jc[JaT��4ݵ��-8?b^õ�k�\�L ����?��T׍��5���a~)U�}�
IQj�}GZ����x)>s�
 �F� �@yk�ض)e4���5��Q �+M��
�H��;-6�h�髕uL[�
xʫ�m%K�5�ń�{�tۘ2���IH�?�C�s*��<�K?c��p�a�5R����N��]30F��Y�6�O?</>������#Kw� @k6�1w�\e�ԫ���"fD����1�f?|��\����� F�V�M�����۵�l�c7ñ���`��>c�5!��W,c��FR�a2�Us�������������b��!��r}3�sA��A�V^�7?�k�	��š��t.��FƐ�YR��5�/�g_8LݐG��й�m�c[��?m����߲^7F2�b�=�6���_1��5Z���B�*��5�c�w��Đ���߷��RV��T�ؿ��'{�����c����n鷘���,��OR��|��D�A	��,�r��:�q� #�W+j=�Q�:qȨB�:�./e�.��pP��:]kD"�b�F�hPp�õ*Xӱg��t<~��ήc�oN�3�e� ��q���ay�{�kD���9-D�������Ie��!��tbp��^�ij�Id{��W���y�X5���@�Ք��T�0i���T��-G]�*�B�֌����R�5ҹ&���IU�` �ٵ�6���k��Gnj7�:R��lE ���#�6e��`��N�`d>=}Bv�8�����q0p,��h
�T�hٶ'����seЈq޳�w��NLCT��#@[��Q�BJ����r䳙w�T^n�R�ӊs��v�D5;[��Ƴ�&�V���ѹ�l�~=�>��1O^��;3�F�i�T7T� �T�5����
����w��*J�F���3Hh��Xo��w����<kê�
S�V9�-��3ҡQ���3ip6����28?` ����%wa�YT���!�QT�j�vd�z��{8��f;��CFՂ�#D��x}8�����=����3�ݹ�r�Y3�T;���<��	�s�j0&����{�ǅAܩÅc �aJ�v6��kb����q��m��s΃����,�mz��99�,�8� ����y*A~KN�O«W���O������?��OR=o��~������9�~���J`tQg�Z�� vzc�����+r����&�f,`N���T9��@�C��%��݇;�N�0#�����;�z�uv�ō-�*���� D�o<��k�s��YL�L����kI�J}�SSgO���=̋q�/f�O�i%�-�l�_�t�/e�S�D.�����?�B�A�i��qt=��L%vRV��������0������ҶK����5�T��JAl���)��'���V�2����*f�V��q=�$��^s+��� ]�i� �4��p��ˏ�р���iC!U�鋪cGv-l&��A��fN��B�[3���4����~�c/��g��n�+�*W�D_8��p��v'+����X^��T-��V���nGj��f�c���}����Ӳ�!A����s�}]�3jHZiͅبm�뢁�궵��f�&�A�����*�?���5 A/�,����۰l�7��r��-�9�#�!��&kY?��d�X����k�������2u�&\\_z�>�����b k�>1e��O�I�B]��z���L2��}&��X�-�jFF�	�z��5�����������d����`,��"�H�<?�����\��n\#N�F���bÛg�'�;5��Ac��`>�'�p�ɶ,�þ��5�;�b�m_��ze�E��<���QMT5G;�z�f+/-M0��(���WYF�}<z'޺�}>��;��cV�m�R>�4y/x�;�������h��t֡�6�F��m3���x�'���}�Ue>�S,��1j���pf��B��7��Nγ��ӧO�u�?u�׬#�@̩�Ot}��6�n��r�Y3����M��R�ؼ��!�N�o�D��S�}��{\G��Gbܤ�@�(����%�d��L�,tkh@�.��iZ�Оe!�3�����seV0�d!�v��� ��A�Jd�n���y�)h�:��8sd-��ٳگI��U>�2��_x�ȟ��}��b_�Q�/F䒖����V�cts�y��LATF#�7*Dk�X|	,�)�ch3.�)h�Μ�^�|��Ï����p�yݠ���Xj@q�����Z��q7���Ҡ P�Γ�Sn@%>
�4\��^���:���)$��Zkn~�~��Y�w�U'D�8f�+9o�_�������o�dqL���Y8��qx��sP��A�~��?W�^\[ce����J}��!Ʃi��T��ce@�L{1c�4i �<=|:�a�����P��ncL�z0�E$�``�2򽔌[������?����ó���j>����� F��5�)���7�n�-ho��4�JI��8Q�8q����[�M��/�F\���������u�<u�_B[g��p�DP��0/�S�A�fW��R�j�,5
M��>�3�3����52[YQ{"�ͫI���i��s��Y��ϩ��m�� �� �G��0 ����.�.Rn��������_�1�� ��lL{ĘhK
�^�:l}`C��:���A����e�մ���[ �:%�O$i��6Hlձ9�~J��ȶ�rpG*2* �AR�:Z��y8V=�{���ը����	 r*��<�V���� -%6º;� �p��cvp\� ��jZ�a�0[��EJ=3�T�%e�n�:W�3�9���(kU �� �H)E���o�?{F�Z �4�QI%D�t��!#��H+	.5JX� ��)rvv���dM�%Ϟ=/�u�]Ѐ�2�W�?���,0� �m�`���(��d�5^i.P�j�y�z8�U��1U�y�A%�V��ެ��c���1m�+t΃}	�\<���\�wg�L[n��8<��b�uwM����(¹`m:���[����P�:,�9��DWR�<Z��H�v�"�}Y��W���;�Fm{�C1'�P`X7��܅v��_G�Ӌ.��+�Wg��d/���*��X޸fLM�X$�,�*��އ�_g,�E��Ƃ=Պ_`E���Ϭb�q����ܬ��0e��ӿ{5-��=P+o��j�>>E�cA� 0d^�{>}�>~��T��#I�~����r���,�<}¾>�IХ�7�����������/����Q�|q&A�͊���h���ZN?�>h<D0}`��&����������Rv��N�i�c�{�����o�=|6x�](����/~��X�[�K`�6݂��h�'P2�l�vk�ꡆ̯�L��Ӯ�ݮ��Mf��E��h��E�_�����ab�j�Ǩ���X�U���{����r�E��(���j,��%5���O���S��"@�?&n�{L�����N��/�;�V����\��(�QǾ���V`~?
��$u�E�ޗRw-{hs�H���w�9�l��ڗ����q�Ug���*
�S��À��+aH]q^5*���Z��M,�0w �,/�h�`�f�~��9@�F*� �v����!Q�@���Kq��l�J�J<�sZ�V�R�Է.�+2np��Eb2��nTxn��u�m��ü�S�pd,RM���C�
m#Qj1dp�^}��y̟�ā�g`a BjiB�'���R�/h?��[1��rE-��^u���3��?����`�m��ɨ��l�E�3ϷY�|ޓ�� %���h�Fd��`�-�1d��?:��u 8.4MҀ��[Z��A��Hp��R��9P��R���DX)H7j��O�X��_��'�����1�x����/��/��`hc�X��0t�X��&�7�տ��/�ZF��V�zԲ�"2�1ݙ��^��b?N��!����ZMD�Ԡ��v����`;������O?�5%-���=T���^(�(=*�g�>X��F��ߦO`�}���YDwh���fazљP�� ���M��G�W2�3�Y0E�0l�hv���AсR[]O��u�^B�6�Lt�OZ�>���J�r��|K1n�Wm���)�}�l�n��]��-��1�n�yq#H@6!��!���`�#@���[2�`ē�5V������Z�v�]8� ����y�f��?0�c�MD�=�%V�Z0�����2 Ɯۭ����� ���ޭ�c�%�d'�?��۫��0KD0] �F�2�ƹ�dD�]:aYb���4[|s>tg ���6d�JP�:�p����X��iB �a�J@m�ᚇ1�f���5N+e%c���o9�!�(`B�Ό���a�����)���{� �0���գ�c}_������_�v����ß���a��d_�@�H��ۿ��C��,��k��`�a��=�F ���-Mh�<}&��ķ��ҙ^y�ITUjhk '�S����>�(lF ����Q���ᙜ<=	/~x^~�׈�˹k�pg"hC��)�X_��wu��g��?�c�����^|�4��Oy=7WRe1*����;v�>l��>?}�
U�a����s����pn��g� �DÅl���T�Yu9U��M�R�c�"������uys�ʒHSHm�҉ �!͗)tm7�U�~/����V1V�R��J�J5�je���eX�>|� �����P�}~y�]�_^��:��F�a�>l*�i��?�T����`�.��\��o"N�
��������q��N3����sRD�2���[�>x9x����*����7���y v�t^|'�}ó@`��N�촸���cƬ���&X�,m�v��y�:�;�p��gس�ܔQ�" T ��S��2ak����P꼶�NdkRQ��w�E����_�=>������;����u�m?��+�8�z������d�˛���Aϲ�S��~0=�|@��F��#��ةEs��!���6uF`$B���)�c:F��!Qn���5L\�j8�}�r�Iu�ϵ*�3�dbȺ��hZCGD���(TV�v[�ksplR�j��Ӣ���iy��'�{����������3\3<)��T��	��	��#�S+�t_T������V�S>�1�Q#2F#�~X�a���(D=�j��S��gq���(B��H�	�Qgl�Z�I(��R��cM��Ο&o�˕2vD��ʉ�*"lt�����:	�ؽ��Қ���J��,�'�����������|���F+���p}t�5e�W]D�`mmȾXI޸�ʔ�Ψo_<K��,X�\�����K��f-U`į�D�gէ�w�:-Qk):��՚��4�� a�70�$*�� =~��1��4��F�Ѫ8��B�>/�ԣ�����r��qc�F�DT�e�� �mp�h������%#ME�0?�}�܂6�VV�^[`D��ZEx֪SD�'m�>�gR�/.t��V�JLZ��"�-�=��d[�zL��g�1k�����e
5 @�*��ƉEꄅ1��K�x:�e$���i���k��Ӊ~	�P����@Z���~��Ȯ������X�%�՟��5,<8��n6�8h`%����J�\Dk�('L�� ��V�1`s�e�Y�(�Ye�З2��WL%�%z��N���54��|����k��O��������y����*�B@LR Y%n&��]g��*��DG����P�������å�0�UQ_��#0�޾cz1�Z@p)�=��C��@��E(6R��
`W,(a�L��O�RYB�ag����`����N��y��ka�&��}/"���e&�o@��7T�������E]9/�+���6ۯ�4�Ņ����V!P�[��C��=ognWQ�oX� 	p3�	�ڽ�t�$�����Zm���A���M�9Ř��Xe������zIk5������B���c����]�!'밆�mh��	�C����*f��\� %tp�H($���W�8S��֏�ٚ^�
�����N��{ٟW\s���F
n�L1�B�ϕ�g�{�H��Ԩx��7������ZamE���.N�O���`�UI�C)�^)�#}�r���I���u�s����8�C��iIlݞv�F��zK;�`�o�I@�Z˘���w�H�f��ꒊ.mF5_*��]1HS%��mu]���}@�@�^�<�6�#3~�����RɈ�	�˧}�g�Վ;�\<9k������d�z4>��y��P(����+�"�x�����X�h��h�_!XIҰ�4:�Z���{JʖQ���UU�ONV�͒^�Z�` �������9��t@k��]��#��jyN�d�j#F��Z'�VK��w��Q���Q!<ɋ������c0v�mf�N����ߵ��S|�#��>N��{QA�(����yҩ�Ue�9��aqDeI���O�J.�  ��IDAT�h���|��I�\f���!��3�� ���48�0�tAOUa8�}���q�95v��9�P,��p�10"�
#�3*�5����K�b-�6G�F���њ)	����Y��5��e���kN}.!O#��z�!��l4{D�P��ܓ��"[m%5�#���S� V*�7j�EF�R���֫�TVF�����Q�!�l 3��c������P�w������d}g%j[)��p�7���:Y<�����+ɨq��P�I-AT�"ϕ��,�yB�s��1�k��l���:�hh{���|��8Mp�OO���e`�6Ѽ
���6N�S_%�:-ul��-���l&K���$9������u\�
��U�s��{e�$m��@�HƸ��ԕ�	��A7fj"ݙ;` ��0�kOy�����dq_���`<�Xe���H��evm�4,1�M�.8�g�	�!���p���6���Y�h��=��=����V���g2v>/����L�5�;H)���L��> �в#�S����pN�1�F�u�)
X�{�k�Fj/�� �a7i��n��}+����R��I����ԓ�\�'�!
����������JE����韨����Բ¸�&#����EG�L��b�����3e�R�x����� x�#.cZo�r��1��-��v5pf��kZm���5���:W��́�zej�ϲϰ��U:m7�`�� �J*>�u.9�k5AEj������=g�a_����Se���B��U��j�m<�*Q��t�5��]�����~���^Y�חH�9�m���,Bå[��P�΂�L�ms�Vzl���.\[%8A{xp�^�\"k�3"��%)h�y/`bPVX����1�����6G� �	���;��k�����A�ZvvP'�z��IYC����?���7Le����'{�׿����}���Q0I@3eQɜ�q���l�I �c���5u.�zM2c�Ύ���P衬�F�s[��Kۣa*��Y��\��"Kz��J+�Z�Q�Ba3C�
c�fu�Ǯ�H�Ko�D�=���s4z}�;�c߱]�n�X��:%ڄ�٬+�G�,��N�" f��'�nӾ���FN���d��~E�<ٯ[�1�j���f�EƇ5�"d#�ь��Q-A�/<�5�GMw�>��6jk=�������o�f;����QS=�f�(���~�"�b¤��c�Ă���ϲ�q���w�އ7o�0��*�LcѾ�׹N>�dp!k��q���+2+ �fƚ�((pc�&�L@[���c]Ewۋ��q��x7@w�y�1�vڷ��Ĝ�J�X�g��R����P�`����!����8��dutD���i��9P����95�k��x0D��W�R��:�,=VJ�]��S v���w� }T��E!F�}WG����\�Po���Iڍ��P�O�J��vIDz�Fٌ� ��\��DCJ��/k� �	���C"KVI��Pt��҇ h�}�(UE�G�2W�ZfD����#Iԁ��ʚ�ύD� t�T+y�ȷOaMF�'Ƭ�Ʈi�Y��Fۭ��������D�r�p��D�M��^���L���c�ٰj�
���6����g	�1�u���$:�[OLS���醓g�Үh8��k@n	��hژQ�=R�F�U� (I��}3�*�l|RQ�o�)[_�Mh �����V l1e �l�J����έ���|!Xn�q�y�Y�)�D�0�v�R6�t*Fm�Fey�ު����Hr��W
�l:)��ɴ}�{��X΂ʾ���&�����{l����؉� �Cd��pN��m���"=�W6�@�6�0r:�F:��Ǐ�Q굤5�T�X�����,�������9�皎cx:e8�8���c�N�;,c�?�{V�>�����l�,lk�5���j3��qM��K;���`��d�6i�G��?}J0UkV���k�Հ����麰��p`b.��L;>Q|��	�6�=�-{M���t�m���}���C�� ���"Ml��O~na���
6H�0J�Â�!�&��j��hշJ�� q�RYK��z��,�r�߬�w�5��$������8��؀֗jM�#'i*ŕk9Ŏ�z�s� ��G��0��b^W��ylM�����
H3�;�"V�w�����y�FU�D��<�L%��q�6i�7R%�XL�cƘB����^��#��fk���o��k�g�� �#S&�{�϶3���a|h�n���7W!����<�����>�Ai_u��:���S-�����6Y�g��[�/�/T� G����]�X�)N�Ơ�!�}+i� �dh<�I6u�D�96��x�5���ͤz�QǨh��"��g	d��1�m�6�C�}��`fay]��_.�Ѿ���8�V��TWI�~����S^��k��NH��Z>�N�Rx9��b��!����
�a1�l'm�]�/_�Yǉ����F���Q��w�(�g�-[1�k�ݸ�'�}�#���Hx����������nMk�^SK�,�T��2�5�8 u郈ٛ7o	�`�:9@ �-������?3�����d�ܬ�C�K��ӓ��4����:/�sC(HmIIݲ��6�B���ѬSpgWd��b�䋰�7l���c$c��"�݈
�`@U�Z#I�b����0*!r��?����yX�6���Ӱ>%��.��C�N����p�Ѿ(��*�A�p���;|9Yg�N�%J���
^��_����#�e�@Wc)��`C�t�h�{�U�W��뤕�Pu��6Ju6�7���2�L ʨ��Z42�31����ڬ�p���h A�FXi��v�8�T��F��VB��>Q`/+}U��q�^*�	�g-�^e%9��R�
��LD�+�Sb>8*G�ߏUPv�85�8AJ����ｺJ�^/�d�ǚ3�_��	�� ~ 
_�_�np�pmk;}V#?df\�j/8�V_����6�HU1�7��������qjj�9�K�zlq�3�K@�*�)Z� º�K���hʴE���G1.},�Ah|�9B4<J#���cm ����,iv'�a����h�1w�*�&��A8&�JZ���8�g��{�-F�*�����(��/��m�N�=�g���T'A���^;*�u`��錮�G�xC����tƵ����B��M�P�`� 4%�2Ҷ~�����S��Ç�ç�q�Y��W���)�dU�Ȱ��zc`��#�;�����f�?m��x�1��:a�vvc�b'q�-]N>cj������m5xR4�@�3Պ��I@l��vR�~�t��C�d�h{a�F��J�-d��iXC>|B��k���YG�0��m&�.gF�F��k{�D'a�Y�m*��Y
PD�)�[(cv-�����`�3J6�W��2���dx'�v�����:�
�4�kH��Kqk�y�Xo����W�
�u��=�Qs}5���2p�������4ع�F@��{��F�Y�I��ܗ�T6��*C�Ie�a��5�")�5��
(o����3����7��(ʿ��`M�P�<5�TTٺ��� �R�댥�3J�1L��bQJX�ꔉ-@`�(�nO�����SV�-�G��}z��o7�נ� h䚊T��g�����v`�:���\�}���n/���q}t�>X�k*�*�,��o�g{�M�6+��땦�7��d:t��/�`�<�Ɔ�u�\F����OE��l7��nc��GǓ�x�ط�*�T����];y��"��d�}� >�`Q�8ve�M�Dc��-��q띻�=���?6`�����1��m�3R�~!C�íg�� U������t����!��L:���%Ƥ�2�V���u�V��0���A����]@��F��g��~�D�وR��L���97�ĪIn��rnu�04�F�e�1y�qNsd
Ǎ{sܰU"�*ʤ/�8��2�L+P\SʒbU	��A�(أW�wj8�Y��e:;���CF烕:����H ��f,|��#M�ۂU�T@N�8ʢ5�>�{�������j}��,�Hm���p���?�U'ۣ`Bi�I+�tJ�f�Z���
F�F���5#�'F�S�����j-��$Vz��tk��#�B���%K#�T{�����Z�
Fo�"�FU7+���uZm)��NҏC(*��J�ke�Z�TU@vZ�y�� p�/��g�@��6�\�saA�*��1��U�f4��`BE�gdQ	%|���s�%R�g��`y���~E)�d1���tp�����0��`���ap��Q���n������}�ee��D�P9Xf�0��� ��>&����G�����rE y/>���=��_w�1Uu,m4�a>���t�C�ߥ"�@}�`Z��F��c����`�t�yy��n��!Ô��P��WFC_��T�{�r���)�e���=�]�N�}��ޱ�\����3�XY
��3LłC���#e�ɆU�n���YJF1�2/K���u,+�Q�8UTK��J�3����UX\*h���
�ʢ8o��;�c�l,�4jX�g����������(i�eMd����C���6GhǺ��8c�]�|m��U�,�ak��a�?�uM1r�v-�G�SD&4V���)�UV���g�s�s֮�[�롔4���b���c��"�� �h�Y�t��Z�E�^�R��̣�-�ZU�v�6��<�((���z%�����32oU?�v��%mg9����n'��������W�`o:�Q綑G�z=�J+�(Ҿ�b	�v*�0��u�s\��#l�����C9���j5f��Eo4�=x_�dN�DC�4��|���%�*ӜӗRw�W�9_�z�/<#c��i�fO�v��=�9�S��@�֙��6孝RȬ�}�)����}�;:�}���$���x����;L�^}cK�?	��[m��}��ߤ;:��t�������q�{(3��3�Mtvsz��N�M�3<4P����#�3\�Z�8�t�5��/_��B��I�N���sa�u2�p�:i_F2��N �N:�- ��C��IlQ7a�1����ܶ@���ؽNg���K���`�y�U6d�١½Ry��&�}����� �m0���idQ�����5
�d>��ϡh8?���Z)i���Q�	�y�oy��s�6o�]��Wȹg;��Ћ��UB��~L�x�/����XU�PH` �j2!
"��K��`��ϥ�6x��U8X�7"�gBuj�ر佋�o�̬P�D-I��Y�0d��T��,E��\�J=���NJ4ad������5���N�0��Z9j����h�I�X�Y�U���C�>P㡈*�'ӆP3������H�gT;� �����l�MK�:mN<%
&Z���iwA�5%7�����TL�I�T�%�;<-�4���0�1
G�T�C)m�9gE]iCc0�ѪzO��/�w3���o���^��$׳\+Z�1k�X��(�[d����6E����F�а}QI�R�= +E�B�9el|�z��{
������o�M�K��6bǜR�Js(g���sa0��������Uۆ9��$����5=#��>���(���	^Ϥ��F|�	�h�^����A�i "��amH��0�n��zg����S�L�i��|Y.�����*�k��ؘV�>�Ac͆h���K߃��L��@�fh_T���ܷ�������������8X���� ����\�i�L��;��C6c�ٚ��Td6��I���3u$uYJ]{ E���]�����3���Z-��6@i�j��s�c����&�;�H��4�`��jF��B2ÕE���!���T�oބwo�]uM{�l*k��`�U���L��ʮ��4��j�d�$UIg�m{tz��֬�t��22x&�֊kx�u��=�C��p���	(�zN��������ӑ����0�Y��j���u�ob��q2pq�TjG
&���8��}����z?�x]���آ���ds�ϥ��v�7IK�G�Z��(=��
��vO�$(js� ��`�MIP,�5d�P���9�G��^��:g�T���y@K���}>��r�P���V�Df,���[�^I��[-�m9�~���Al�v~_[�����|�Yg�F���nc�8��˃>x�����h�{��:Ct�^�M�ZU��P���''F�� y����EĨ�L&٣#)����3gUj8���[���eY�����r�����tG3�D�m���p�X��;�����**CE�|DeT5|oF��V�x6�k�jJtug��������~qq> ������^(�Ɉ�==�ی�d�	�2��6��4ң�p���Ձˡ�G��F���"�o�Gڨ���B��\E���8 ��Ӫ�7,޸W\�U�2]'0E�,cEm�5U)� �?V�b|�9�l2X���T���&K���X�6�w���E��Y"Ctԕ��Y�����|�
۱�Em��ձi��F5�84���aN��jĵJ�7���e��8�oBT;j$�!dl�2���F��jFHZ�a�D�xm�$˟H�aIlԑ�=�#�l��_kJ�>G߁qO
�pm�_(���.�{�uO�Ty^�q|/VZL$�5�^ D�<�惦,�R&��'Q��iI�FP����i5�x�'a�_���J�q�]Lh���8W,���ꉓ�����q�9a��
��1n�y�F5[��U�V�z������Fҵ0_��٫�8@ ��rA��`�"]�`�F*մ:�3���S���ԇ���J�S3EA���@��/L>�3��T0��W>����2�$�=��R���Źm��L��
�_��2�Z�P�Ki�(�aE&h������򡮚8�p�_����r1����U8c}C���M�'�����[��Y9W�k�c�\;e0�O���sh�|*s���/..�O?�M�������*�H\{�b���Z�J���a.6���p�1_/�Y����^>PЛ����,5؍��<���� $�_���热{|8��wX%� �LJ���s�c�J�i3|�sI�������Ë:O��	�/�5l�ĺ�dF��<Ɇv��������Ra	��X��Y�Q��`P�g�hZ.L�	 ��V�b�2��SX*��yw�ؚ�
��x/�>�X���5��a����	�hH
+2u^u�C��V05
�\���+)pZ���\w���Q�v4e�:Y	�\Q�"��u�4��b�Y�$��P�K�Ùuc �e��6��1�q��m`�Xx�m�o�km������X�P���)��p����������^63����O�nC\�
xw8�m���Ú��S���!�n��L�/Z:�9H�5Z�h�l��ݧ�gdClZ���K����=�4T�A$�����׳�h� ;,[�v[�>+]V��fM��L���Hj\����	ٌ���w�!��N%@�g5#���a��Uϟ?%��*�o��K�m��Z�g>_|�r#Q��zI�24�1�H6n�тN�h��qd5�.�4ɂS�nȮ���F~̑6QZ�v ����_�x�tv\L9�����Yz�u��6���y��iU���k��R6k�R��s��98"�%�)�^����ӪC� J�|�} ,��v�ЍW8�`�o�	�uCȚ���4J���Q�u7�`�D1J7��S"h1�`%:�n��E�:o�vi�&V��h�#a,�
V+�SK���yeƼ��`ЂU#,/ N-_^���)�wj)3
�D���lA�M^��L�)~��OfZ6�H٨�8W��
�?	�����V�W(�]�%�>�DL��U5ڸ�r9�}ZSKgu��`W�ib�Eת�v� Z��k���i�ܴ�<r�8�A��6~��&r�����5��J]�~J+L�J��aLa����5�^�Ӷj��M�y�~H���t�ZJR3�2��4j�P��ru}���Sf��Zu��	!G�ߘ�U�>/��or�p��|%�3=�;���i��M
ԮWf���$�Uν��4�O(<���.�n��8X�>�}b[SSm&�1e��j�ds�D[������:��g�	���a���y �,(u�F�2���c^(0<GJF[��2�xA٪}�7�Pl6q�M��>þ��u^�`�XE��%:RK�_`�u(X[�X������AWøA5O� J	�N�\��2�Mb�&{���B��9Ю����`�
�5R6{�4���Z4�`g8�s0w�2jg�^"4t�h2@�L0_��Z��j¡-0ޫ��ڵ'a{�%0���e�!x��k�N��{X�d�բM���0��t� X��}�m���D��iJ&젢Єm�F��a/���L����Թ�2��U��KX��R��U<������\n�׏���ܪ{�X��_
�&�
.�M��1�/J;�>~,u3��(��PjF;��UA�9���>���Ӹ������� �����z`��+�C�������"ƀ�m�`�[1~���p���D���lZh���4��F{p����I%`=Ŕ
�3� Y (q�4�!�؈3�I�/+�o+н/e�^�V�`�o�j��T| �瀰&@I�JB���KH�.����c)7���tT>��b I�?�6J���3���~`'�v+^�ڀU��&���J=$�joF/.��� �R�N�L�w���H�-\X!����L*.uQ����c��p�������C�e'��Wtds��*9�("}��B�����~��wtT�j́�.�*އ�����~���!���Ø�nU9�S#is��a������ߧ��J��a�*U7��c����`����`�}�|FF��O�]����֣�w�r�54{�e�rê]�%�;�5bFMB��[ڙt[�o��s��6��	=���)#��$�(J�u�f�0�떆5x��0?�>�>r�^�]ɳ�f�Y�n�=�>�H�F�CP�� �L��iq@��xƹ���hQҝDT9Wڸ�dv*����;�;�����H.��K���,pMn�AFi�q��&�LB٦�m%JC>o�}�.�(�Q9*�÷3��m���c~��Ư�fg�^���$]��W+je���m; 6 �5�Թ�m�w�AFڐ��ZU?�HpF�a)�&�W����i��]ֺ+�
�V:��l��z]n��1Z�&ۨ��j�d�Yv����g�7�$�����O�B�دS2�W��# r#�痬R�����U,e�v�Z*���u8=9�~�V\�_Xߐ�ÔK�w�nk)2��T����:��6�s+ƽ7\PGS�d�{9��=A� ��H�������?�>���C���xd�֪-�^+����t���1O  d�ʼU�M�q�L"������&�>�!EƇu��[y~y�:���߇H�i53�cc���p�1pp�v�S�;j� ���3M�$�)!�N�!��+�1�֤���3��!ؼ���1/o��5�L��s�R�$5Z��kW]�O�a�E?D��Z}C;�����~��M(�p�>ꚑ7<�!p�R����X�5/f�X���5x,p��[�#�� ���U,�f֏�%y�<r�*k��6'��]���P�C�o����2��Xf�P���D�T0��V�GU��{��M����VXc�|��m�mL��ͫ��W홖m�s��U���u ��큛.�[����y ���������w�Yd$ݽ��1���v��Tv��@��!�ܛs���c���$R���a��;k$Ku[� �"�`�����ZAT0��0�"zǛF�:�("(�3�kr1��Ӆ��a�kta�-%�#�9Bh�ot�g4�|����+e����z�L��҉ID��J4��j͒�I;��@(��mḮ��uZ���R�8' Kq��Dؠs<I�ڃeb�0h0R�MR[VZea�H%��CGТS� Uɇ�C�쏨�,eG��P-8� �Nz��)֌©4�)QF1� F�>�(7�ަId���!��Չ���V'1�J�t|D�Я�hb��&�U`"0�U@��p܋�:�#��
4�
����V��R-��*��k�BM��r=�뫰N06������9Z!X4�"G�8Aӫ"��u�Άհ�:n�R��3�șqF��礞���4��`?���zp\/��@'G��a�M�&�I�d�H*��"<)b������'��w��9�\�ތϙjaXY_ {���։(7ل덏W����;�޽l�����H* �1[K�]�����Rig���٣��&Bm�V-"��Jė�������n�o��V�5f�ܲ�/��{�:���������}���y���eI�Ե�*���1�/`.���q���	��*�`�5���EԔ��J_KO��4�
IS3ԑ��ܷJ�n~�`�[j/����[vb�Y���T~�3�B� wvڂ���(Wt�o�> tF�X����i�f�c�������v���d:�"R&�1t�i�Pe�NSFﻥQ;埮Y�b)���LD�FY%+����%ȡհ�0�u����ڥ�R�U�87"��g����\ I��@� X�x��lX �҆�5 ����w�͛7�훷�Ç"�|p���:FO���?X=���� ���IoKF+�%`�A\ٜzj�G!Kn�w�Q+r��  ��em�@�b�.����VV͓vP���LٌK�;у�I=����^�aV��dmE���RS��o��O�=�`m���J�~ ����)Ŧ�O����P�ϙ�2�  s�8�R%,8 ;���1��5:GX,}��5�mTt���j�\��RҼ��AA$�K��`,�I@�pLK�v`G�s�@�O�%+�J��^J���Y]�~o�h�"��{T�\��$^�{ĩ�}�o)
ʕ���L�}H��6�D��vM�����`�5�-����7�qc�Ŏ�ZR��qww��ǵD�����?��ŴM��Ř���Mv��>?8m�r�-��plM��=�d�zm�d�_1�i�̉/d$Է��~��b��>�[��ϭX:�����m�w` eP���c�T#�1�ŝ)$�4^`lbr>@��ᘛ���j�C��/���vE:
JI���T����K�EʬnH��&�N���D3e�T�yRi�R�ܷ4��9'�L�0B=ZX�}���v�Ҏ.+�F���i#ʾh�M�|0��:̯f4TI³��Nq�b�F���`�UW�0'fLi9dY\?"�8�(a�X�Q����@� ��}�zU���c~d��u%�R-���(5:�`�4�p M
׎�tx������ZJ]�g�F.ʨZ��`q�¿b`��C `��ҜК�+Z�t3L�Q�
%���Yn<12 D��DP}���oy���`�V�G��38Z�̨TD�S]�j��V�}0:H�l"˪�dU�	���V\��q/�Eѳ��ɭedn�s���C�A�P<P}�QYe �Ю�g7�Z���o�/����[QQ톹���^S����btl���ce.C�p���aP{�&j��jc��p��V�X�(�~I�mDP�N�g����z9���vHy>��l{�:L�<���.f�r�eۈ7�}4[Q59B�g��gS�x}9A&�wk!m��w�+�����][t�����[����u_����'�d��2Nظ{��.'���;V�/Z<��U�"V�
�P��Vwh�N�9��*/����z��Q��7�.��3g�Ř�P�T�d>m�C�*�r`k�cKu�����g'��
�unf�Q�{)���9�RKJ_�S�`��[>1]���p+�#���y,��l%�q4����E#���;��w%%V :Օ�׷Iӱ0��y<:���x�`�·�;DJ���N�<eUQ��v"suM�돟?���އO���BA�P�B10��059G[�v��o�{�X	�a�\��K*B�s�fsH���d������@�x�]\�3ힶǦUQd�(�S1�JSV�UX9}z�a��Z�����kT��Ze�Q��q<�>�@S���Ǜ+�h��A��ze��dAR*Ci�'e$��2Z#�c`|�jd�Tgs5s�;���u
�V�J�y!h*|�GR��W`HQ?�W�V-⽰ ꚁ%`aCAf����Ss������m�����Wl�:���[���A4��`�X�T]0P�G�?{N�:� �F��\�),�MS3üt�䄏��Z��D��=�*��)�Q�y�W S���@��-���n��֭�7���^��ʲ�&3��g�q*���t#FM:�vo_>��k���hv��l��:��k(��׸�}g�C���v؅���1?m�4Z��������\�����'IpB��a��L��U���Z�-
�<zt�1~�_�����S鍊�>J�,��M�����(}��N��ƚ\��:����8E��	�J3.�X�)�������u	����<�=|뒋�j3�M x�
��l���=���������l �� �ݐ�6tE�w��z)��T �	)3e�V�,4���2�2��2 G*CE70����{�`�V��)N��:=����Xq��ķ�(�$�-u�(�g[��6ad��~"��G��DtL?���sf����1Z��e̗�3#�,����Z1`(�9|cg�j��.kl�C�b������ȱh���΅�aH�1��7C�;����>�
A&n�<L����T��ȷ=8��D��E�uJ+�R��;_27TU��2	��<"��>�P�E(�-���(>E����Q*R\�`D?q�*~'9�:�F���o�	�-m��i��Xm]�`12
D����_��T���s�n����mY[� QK-%�z� Ü�~�����^�\�M�p0��f�O��ꐺ	�u�R����X�su��1�hp�5���C])�)`C���F��D�@�0�?�~���v�##�l+r���o��#�T(}/�}' Rul]���L̬������?�3Lj�N����H���lr(�����>����]6H��Sa$�y���͊;�c�N/qz/{�R��B��hhUX�_鯕A~g���*$��:x��~��*XkNWR�����y<?���h�lh`�aT��|���[n6+�qpm|�BC�S�Ql��h�kÌf�ɀ�{e��|�:1uFXlN���j�rm4�?-�އ��2?�)걸����w���Og���:rx O �k8�ʤ�b5�T��٬�V�	��	@���`S �����s�Z���svv�߿�/�ç�O����jE�L�v�"َ1F�:�:�Ķ�T��:M�U`��5j ��C��=�3��H�]vP���A8Z��'�d���z�i4v��I�yyCP�vX3"�\И[k��T���a�N�E!0�y^4v��L��H�����a��	lk!���Asߌ��d�,�68c�o�i��<Q�t����PƩ��i�0����:�ÚzҨm��R�+��@3��Q��p*1��k,mW���5��Q�����d-��	�b�@2��˗��uxt�����IkR���p��{���Y��m�g�|�*-�.�c1��E�=��'5>�Χr�~��ɖ��ɇ:�$[��t��:��]�!�0G[�����A���l�����m��Ŗ�_,���g�3#��q��n[���{xܦ�!����7�gl��v\�����8�=�i��okD4*RԵ.��Eu:Gșw��w�O���e�a���}�|��[~�_����r������%��5 �Ԧػ9�S�]˺�.< �.1�>qN���Y"�`��&dTw����?�ɿ�S���XP-]���eh���Ғ��+�ݚA(w3�OF�
`
�����b���tZ�IT��漳2�����m
����d��8����������x\ɣ�[[���۶�H�*��u���!iD�����`��8/mIÅ1Ӌ�� �:��tE�t����V˵���\2/�F*1�Ȳ��}�{����T�Q�V�� :=�ډeK{����?���!�i��`��0c���u���(*�J� �A��fqL8t�����)�\�P�=��JJM'Q'�#��Ǧև��d�(�`�K�l)�U&�Jm�.֪��}�k` ��BI�u�u�A�m�4z�����&�5G��ʲ�t>����
���AS�:Ӱ��Ε����y~�3��"%x�Z�v�B�@�@�����(4t�����%Eo�rk~G�S�9zk���ڡ�d2A�`T�|�<�c��r�ۍ�o�e��L�U�,�ΐ>���}���̡���Vx�8؝ǡk詆���_3M*I` ����췖ys;����
�)>�|���,G�#>B�Ok2a�G�	$�����9�Wg{FKSLi�q#g��� ��g��25VZ���i1c�e���bM�}�1{�~��GC��iN�9�&�,k��g�ώ�8&g*ǫ�蘛g*�����8��W7����u2:�!�y�2O#��5��9���kS���m��������|��4�״�`/�}�	ZK7dYm�\�-�>��:{:k\�Z#��^�n�������,���M�mrqu���B;̥�*�zr>���`�	�
HXie.cvRp�ߛa||>�����`�c�f@)I@���O᧟"�l!����1�	�� ���#�R�2�u��&����8^��/L�p�_	h�uB:�� +�i���"Ŧ�Y����ąU��ֻ�I+��&�ۭ:�ת^
p�I%2T�2VZP{��"��&0֙��bN�=�T���k{��6F���g��V���*�I�X2����dޑ��U=/kwa�j�X8��.��7�"ju���5�g���[�
T'_����DLw\���1n�̯�	�3A����~������Wm�(5(����f=����"d���ܽ��&��]kӫ2�9pL��#7��i�a IٓoGh|��w{�V�:��:2 C6(�~aN�h�Q�7V�����>��,����*cO�S�Qt4��,�Ǵ�Ɲ��o߄��g�~�Q��j4�(B�S����JJ���.=�1���ܒ�Β(?Jt��h���VZBY�(���"��K�Ҷ<�{nI����eN��J��H�q?�s�s���Y�Q3#��+M�k[�#f�J`��//������W���H%��UļR�N"qI�����,�:�Jb��ȭ. �F"fK
MJ�͞TlY޽�q`�ͯ	��a�4��h �������f�{�6���ϼ��{q(J�I*�H+[��I�C8������̓V��u6������	��JԅJZnN;�ZI���T�X�ќ-�*MI�X��Dx�Ю��e%hq�U��{�~�#Ut��k��S��;�/�˾�hky�b2
�����P�<%ն�Y*uN!(�WS��/��A�*v-�ra^Zj�bK�m˔�8�m�Uã���ؼ�o
^�L��}w,9{��M�8���)�V��vg�d6�ʶ�� ?�[�g���>�{��4-�bu2<T���W����sc�G0�hW���4��D���.����+뼱�x�I��h��\mD�U�?��#s�h�TL��r��)ޛ8h�t��[��2T�^�2�������6AS�'�u 5��� m��y���1�l# �	�Zias4�$%��'xS�bݑJ@��.e��\� t@:��`:�΢������Z}6���B�Z�����@�֧b����:l�������SۓӧRU�7�m�� �ReA0����U�Fo�\���:̪`s�
�?\߈�0�;x�R�pl�|U��s/X��9���3���'�UH���rPFǃk�s8�jǤ��:[�>�+� �?��vD�UEs��7Aw�f�Z�7Ik�aj���T+󧤴'�3����.Xd�*�B�(��T�`�� ��L����u��b�x֊��&.�\h�(+l��넌�cʜ�xܚd��upI�ٹ����>�߶X��p3�H�͐ɱƠ�t�o�h��;�%�L��`O���nm�T���#pG������gY܏��=��{l�9}61�Q�T5�}�4�GP~�[~¿*��s�uo~�K1�s��yG�r�K41��;r�U�]:k��}��Z�o��m��m��;�#�*(�+!y�<P�\,!����;��6���#�����5#8W�7PH>�*��cq"�P��m2���}30,�3�"Ewa�$]dqaY�Nt>����R�1����f�u[�E�� ��JŠ#Y�
[� �і�uGRL[g�e���G�t%@����Ѵ�Jˈ��h�>�%�F4�8����B�h�`���$���P�%+F��HBWFiJ0������|�-����M������+�M�n��Š2-��,ڇ�K����o��%s�͡�H����4�X/�6��9��w΃Fݠ�PI����O1�F�Q��Uo�J�-�`ݥ0���m)�(%Hg<�=?;����D�߫p��	�%_Xr�ю�oȜW������]������7�G�(l,��A�0�~
�h�ʪ^�jrj,Wb
�U���2��,�X\d�y����[kr9E�J��P^�85;�gӿ\	B�
��w|�_�md�?�oe���?��wv~�"y��#E1��Yz��;�ج��i�dN�X�V�mAAf�`�x �R)F�g�A`����8�M�7{J�K
9��F�4�+�Y�i kY(`�cf�ib��"`ء,�	���S���>��R������*[������cz_!�g���ɕ�ݰ{�t8���F�"�kL�J��l��\����Mo����jf����Pȁ���C����:��dT��2�=8�8�'d�F�PA�W�)�c
{A�Q;T��*$��1�JY�Vs�y����T��oF���Y�����i~���������2�cZ79Fp@	zy� ��k�@T����ܴ�,�EP�g�@�	�� _�~�J9K���+֗T ;�}�A��Y;���T�l�~��E��Qӗ�����������9)K��J��Ǿ[�~���*��PӶ�p���]�?�.�]è!�6���p����/�ç��ݿvwih*��Mb�u۶���ir�=�d�v����FȆ�. d�1������5�
يutd_���&�;��W�
�5���E[�lʟ���O�IZ�M��ةm�a�u����L��]F��b�����>���7e�R~�x/�7��'�4��l��σE%~�{�Ie|���.�ZEC�01�Dܯ��$MQD_�}x/����$UTuw�7Ra�K AX�H ��^���<�y-���W�� v������ 1v�d'�.7Z�#���c�y̶ ��ۍ���v?nf  ?.~�wJ4��yҩ�$�h�s���w���E�=��V魍Qg����A�͡��墖�����)-Uu6*�x�t��?~6ط��u#CP�ݨ"|c��ۡ��{M��i��:	0��e^ot`щ�&���Ϭ�QDy5�Ϫ��f����e��,6>�v��bb�rGf\TU.9�+��4b�x@A���`si��J���X��&xMj���e�e̓caeU��h�c�],�����Ɇ߽�\����;f{zu��оu=�#i�0s�-Rx�s��%�'0���<�וƯ�yf@��/�� ��{q�5_�����|7ۀ@	��!�$�A��'ϟ>�R�����,��k��.pܮ�4h��X����ˇ���r�j`K���B�.w�1ѮW�^X�"U̕y�Z�f�F�M������إ��mf�%H�W��$\X���F�4:�p�+)%]��Q��	M� ��)�Cc����CfV��}r?4m*�.z�����K�h�̯]�r���Ӥ�ܞ9��������֫ ��:�Vhꅍ�MY�YY#xd�J��1S�B������y��y��lׅ{�Tx���\�Kow��Md�`Q���N�3h2uU�j���L-8c�df��N�ϬB��reZy��Z��6�� XB��pys��2U]�G�6бV]��? �i�(�r�g�zyE��DT���e�YR�T;J� H���l�9e���yI�����@�X�e�T��Yu�^�����ӵM*�ɹ�����ɲ"����KZ���ѡ�)�2�0�n_���Ѷ
C���z�dK�V���$Af�Ze)�nK�(1��H�c�.uy��y�X��Ѷ�j�Ύ��]�ܬ�#a�{�Ǒ�7��n]G��ݰz����}�f؅m�F�;E�;�R~��������!&p���e��0/����xr�K��g�$���;ٮ~�o���l~���5}��x�Ɍw������6�s�Ki(��#q�)�$N�:��N�ŤUcO<`�|>;c[@q�3R7�#�� BS��X���=W�>^`�ԁ�]�j�]�!�H:��,%���J���Q��'���a��'��C<gt�`O>�#:�(%#i;��{�d�yU0,�8����O����gv12L�,δ58=�"��Q��꧈m׹q��Wّ�R.)r��(���L���ua�G�W�N�%��-�0b��4�4A�p�٧q��M��gϵV��ג�R�m�7�ɮ�@�1E�P�������*6q�����G��'L���$*ur�.�!А}[����ūW�勗�O�&vZ�*��tX�ik*.H��7̨�l|;�#�9n���8F��v�u2I����(���:ec	����L��"�<&�ԃ�p%X��G8��w�n�԰��Ic��3i7�W�sZ�rw�h~0����-���r�}�?���W :X���W1�����1 U�~��S�&��˶���~U��d녲?�3ΛZ����-:���hkR h�-/����n56��T�Ђ�TD�Lӯd
�ۂ*:�E8ZfFI+�LC]��j��!M�Jb; U�Z}	��H��{Wl��AM���J[���G�����r��,��m�óQlL�ye,K�$�y�V�VB�4�D��$VT2��)���ۧ�>`��D�*e�����smS�9ffV2��������0ujP�{x�x� S�pM�ά��P% J}}�*��t�{r]f
�HX`�5]FV�i#���N�s�ff&ZxZLm@���E�����(.�Fz
A����%4��!���+�CO�	j��z��d V�h,քJ����I�-dݑ���5J�����\~m����
��j:Qx)� Licz!(5�U�g��� 7?�3��݇�y�����]j%���sI�R��0�3��4���������J� l���^�H�-N~�۾��(�]_~��qM���xD�G�ۋ�H"��W�k������q�/�����i?^���ap�yqM���u��_����<�]�Q�k���m���?��
'��$Q�JƮ�F�%*]��ȯ�cVE1�k9b�lQ��320[����`B%ݝ�<����I��/4����t��KQY�͌����#c�e�J�����P��ch��>��3�"��.f�J<�[umE����i��09yrʣ@��˲�x����F�L�Q�@��
�Y�@Z����jM�atP+d���C���Չ��j �ǌբ=dҤa��%z9�Q�[��Z)�L=�k�b��+?�v�~�,���l�+�/cc�ց�q��܁Q�(�R�p���A�k�F����w߇��^�gj�[?Hߜ0[�$z�f��*c�HI�U:S �`�rD�B���Z5Q��ҝd�yz��0�'`��m���?OnP�7y�Ԑ)���8���s��S`���K9Vv�^��UH��S��ZN�^T@ �i���<�-�R�_vY��)���Pس�O��g|l�w?��,��`�����|[�ٿٸ��X�;�5���9���
��l���zP�K�!���t���倴F��$�>��FƓ��ټB`̎o�,�����mD���B� �:���N<���+SN��V����ؽ�˧o�d��{*�b?Ԑ�>���蘉~K��1c�}��l3����m	$���u�,�F��Y�)$-�GDL��y�RQ����b�3�d/��4�)A��*���}��m\h@�J��g�}�`��
E���`��ت�2Z{��'�sY�ԃe�F�y�D�s��4	��ټ!����M-�x���/��������4M̪�����0�j�o�L(�������^��U'[�QP����Z����X��h1��B���M �fZ�|웃j N�dvO�q�;����~3�/S��
���qak��ɼL<�Ӗv���FtaS�C�x��� �`�W`W�o�7.Yyx�k��jyþ%=�G��u��>�Z+C��O}�}��l�9L2�F�)��͡=vĭ�x��x�V4�؊�q��M?=����)�\ˇ�t���|���s5�F�ӹ��)�h�lo�A��b�u���h�ʤ�t�<`o7�R�s�2��'��[_��1(ʁiN�}�����o��{x���b��ݟ=�`N�;$��t�.�\@�2�	�VdX�Ek�u-�H�E�lb7��X^c1��%Q��a5���6�+kܒBk�8�{5<�E���d��*3X,�c߰Y";
|�"̘����h�M�"#'z��[}h
��IH�9�`�po��53����:"0�j�;���fɶ�Z��H��,E=N� ���C��=��U�2��F�PLu=�{�M��o���~k�z=6�ץ��i��GJ���\���������-/~Ğ�IEH�O"D,y����Y �ؖ-����j�C54�����V)v���`�]�XX=xV0�[�HfO�F��@	��o��N�h�H�dR�M��Ζ�_��TF𽗅]��nq�}��֫�JQ-�Y^V*wN)��ht0ѣ�)�q)J�^e:*yM���|-;����r}�Z�������]=��N��e[���m����2�mJ�!4��i�s])���l��6����I���{;���i�e��d���y��C�O�����b|�4�ӓ>��}��8P��ܣ�E�A��(�t� �]X����gy~��;Fr��$����A:����|�Z�L����X�'����/��sͭZ,�⺪�i�}3�z��P.���Rum��)�����d��n�<���I����AK�pq�4�Ra���s~�,
�k���Jo���rK���d�Dm��L��W^��s%)�2b�-#��d$�|9Gfo�E}�LC�Tc+p�k����!�t,]�?�N��2]�N�͒�cV4�L�N�E/]���6��y	MF )ԽIɁ������������Q-"�^�gs��6�>#e;�9}+�R-�՝��.U��$ih���
QL��9q��^|�s��{cw_ҿu|��jM�yG��Nc^���B��J����Px�&�T=΁u�gG�w�ꩽqMJl�J5k��-��~�x7	�Y��g��)����'��8a��4[4٘,���E��@�ʙ�7,�+����v���x�C�_�9־7�Wn������id�|�ey�9z2����󙮙F���Dl֘����tkJ�i�4�+���<X펫Z5����O�yG�װ;�ά��p������;�����[q�=� ����m�W9q�b'?�������ph����u�y��~�<WGعz�Dݩ/���I��ϛ���F$z5�h��Y0:uЪ�\T�"��
�Nд˽�Nsև���7_lJ:k6&m��?5�DDX��������Ij0���w���q����FޗGo��Y�ؘͫ0�/�=E��b������a��,�E�zd�qY�j���C61��I��%�`d�s	ZY�`O����CMv/[N�՟�P1%|m/"Y�VB%�
�痟���R�DF)k1D�YԳ���3'ôu��j��%�c�	)�b!0�j�t�Z�RC]�$�:�yDP��#�}�?U����W�W�������M+5��9�4�[oEbI�z%�H�Ŷ({`�ee��`H��^<I3|C56`w�%�7���Sd�ɩ�!�G�=�����ro&p_;9�T8��~]e���m<��1I�X��s�]�8�F��?�l_������s��?͝�=�]���g�`���p�� ��#�8h��뚔�����~Ȏ��e3U
wԀ�)Íf&�Rudܱ������,�;@f��C}��$�5���BK̎����F؈�1#u<t�� iܐ9�Wj{��Z�[�e�Yգ�/�PѢ}����w`h�9�m�����ձ�;�]�����1:���H&�* .���Iݱ�`tB��Ț3��V�0��f�J5b�"j������˳K)k+/մX�>��[.om��<��:��[� ;�Z[��[���X.@� ��}Y�3�*�;����!�־ϟ?�O?��G��U��6ڿ`���U����
�^�\Yc`����벭���T�U�b�V��j���|3�[�{��g�0�ǖ�b��
ϝ�C�t����W��?nc��l�ɸ�1.�Q�CRݠl�{]*����m��mU���o�1Pm�}M�Z���r�"V���@�t͌;��8�e���!<��8���'y��>�-�������֑�t�q�b�T{ ��g9}~E��ƹ��Ƙ��u1��J��ٔ�ge���s�A���t�?��6��x����潱�\�]�+M~�+i����)}�m�W��.�(�s�z�Hzzl�X��W��D���*P#�	�&W�5Xl�{tB�VF�<6a�YȖlL����g"l�E�Z�pݑ���h�����"���;��Uj����13DJ�@� AJ���Ѳ�V�ߔ(���������u���}�{����kK=d���J�Ţ���"e'T)zϓ����i/��a*Ԛ�a�y޼~���>D0����)N�gG�|f���^��k������&��ϟ?q���<4)P��������j0��)�^��캔;VY�Z4��-�Dk��	v�7�4���F��Ϸ���?{���8��	�d�̬,��rgg����{����i�Z�"?�x����%�{v��$�KsSn"W�$	� �����H=�U�|ͫY�S�b�"�M��y{���.��x�����'���������㓖p	��/jq<��	Bّb0��}`��{���+�*?NT��b�P���\��
�B�[��-����lġ��>V�xoo�aɴsN�2�t���ynQ2 L
eW��un��Je����}�G�v�%���l1��|�r���>,�`�ђ���݃Ċ����޴�y-v�aM|Go�yE�&m��W�p�x���:҅�s�c��%�
�LQ�t�8e5�Ls���;U�M�gk
)�f���@�>9dõk�K�`�%F�����_���\l�:Eד���~����@\��%L�����@�J��Z���va!BՅ��f7�w�ީ�3����_YLPv~Ԃcp�nm,]���ZF�U��(����ih�xJ��堌N���>�n��p5�;��'�t����p[��6-v`F����a�ྚ��$4�u�t�2�gQ/��H���~�}E)�o�����X|/+v1s�_����F��x�@��̛Nt��w�MT��?Ȣ��:��n�|�|.��K���Ri�'� C-2��C��՜'���;���HB< Ɛ�j9��b����;A���R����l܂�֤<*&�s ȡ��E�Dgʺ�3�0�ŉUC��P�Hr�T����%�}���-�O����8q� �O�_��������!��fe�-�I�*X����
�xl��T��$�CH�)�Gqf	��LwE]�Xy,I�1�.��ZC{>g��j�Z����>U�6!�����Ba����V����׺Y��`t��WHf����|_�DlN�M��j�@'fr����[��� �|r	&���4k����A��p)�{/L&��z���

Ȇ�0f�B&�k�&m�.�Q�'��X?�#�}�{@m5ma_�g�A�k�ﱁ�c��R�^�*�6���%��_�<�x6�6�"�[J�4��11}�@�p��w(�1�Q�ؐ�&H; �cpĠ����閵Q�XG�]N�Y���N�L��5�	Ƌ�J=����9dp�hf�fK17X� zIpz��e��jV��q���LR씤<,�[���������f�Muٵl��"V$�]�����	�}�Y�*�bϕVI��J�2w�J��j4��83��\,��U��`^����ts�E-<�O�?K�B�����e�S�u3�P��$�?��aZǱ�6��p?�����Z<�N������L���MC�����c#(5+�F������>�i6'�`�!=��`�B�D���YpP��^��y
��a\բ�5I?,�俴m #�Sg}�C=p1:H��
�sP6}I�nX^�c�E�g�{��	X�Q�T�(��T��u�(�CX�4w�p�p��Wڿ�-/9>s~-��#�RӴ,�;}�l�	�U�����Q�(.��m/�O�P����g�?,3�7S�kC�����L����! �$pS�"�쫺��AOH�e���_���w��h�?<S�10.�<{���^�@���LC�{`�����Ħl0So=y!� �h��9�{A��O楟{X���������-��ڼ!M� ���_�l^M]Z���d�aR7�MHLI7?�A�5�hJ(hT�#J{N�F��&�Q�~"����2é��:�N���������k��2�I�r�Y��)L���;��5�Q�wh��㏆F3�������,H���S`�����j���C�7��N���`t�P��@0�8O��>��U.����%���@�?����|W�ؔ�r'���sC����.'��TBT��v}��:'U��5;a]�zq�z�(gV*.�T.��w�΍�tY��������Ӌ�=���R�d�Y����\@&��[(����qn?���v� iwKEJ*�h0#s"�I�;Uvs�Bv�*� �����!��
�ZQTg+�j��a�:Y��B �9�ÏZ���1��0��t�\�dm��DC�F^~����.�j1��(U���2�Rō�Xg�뚊,ch���u<�����]�e���r�1���������1b�y����.5����oU�K\����o���@���%�0�{��nn����^wߒ\�:�c�x+04p�^��'Dw�|?��o0]������w~��v�N	��!��yX���sP��ֽk<�Nx�1\5%Φݗ�B1)������J��� ����{��]g�V���������~���>������ˑ�i-�S��txf���%�Sf}X�9������i>[�R��mٿOR��;��rI��k�U�8	�|���5�~�f�%�/R��9�QW6���V�H�z�c��j���Y��9Л�&Lz��jc���"p����^�.?�n�x.p���]�gc��	��jI�̢��XX�M�v�V���Z/(qcf�c�H���>�Xr7#�pej���!3D��nR|��B��I���������`mS5��h���HE]�n-E�X-��WH�f0e��c{Hܱ�zz[%����ԅ���"�͡;����X2�j���"�Dl�V�8�%���A3a&�f@4k�f�b+�軟�U���lby�X�
s�i|�%dF�.D� �'����e:a��v�iX՚��a�Oc	������ک��Sicq7Po�,�j�y2,�	+�[����cPli������z��E���~r$�O�K�9���X�Q�3T� �؈%WP��]��X�S�l(wU���ngp��lV�&�q�L��4����rIJ��y�Y��F��J�/�ʜ�8#��g� c����յ�����C�+����R����[Y�L+Lu~?pv����З�q}|~gm�F�� ~�ٺB$�Տ����e�N��t�:��m��H!�VS�W��4�g/;���8�<LB/�M�R�k!٘� ������`R��z�r���ctέ�H�dD��;[w�S:�����;»��������s{�8�%A�\�,YJ��w�I�hsE�������c��7���Y�Ҵ�Ȱ��Ż�\<�;_��Ǐ�o?<����H��>���,g�[̱��%��s@S����H�?]�ڄbĺQ$&�Κ�D���Z��3���^�Q�`|.�$w��}m�j�t�m��̅o4�Y�p�7���'���h;���+������Ak�dY���i�l]�^xHs��\��4B��:�ݏu�!�|t'(-��KZĚ>��Q���ͧ+v~t�:���OP�W	D�O$[(����3|d��@2�Hݭ�f�9<�橝�7�����D� #���W.(�$Á1\n��)-Me��H�V�S�(�6�y&�qݽ�U5��d�Z��
�La=��̃���LeW�&ӂ�"�ۑ2#U�R�3j���6F�=��w���L���s��A����s�per��D]�0wU,�4�U@�X#��6n�@u�~g����Ü�<��	��0��}�,#j��j'�SM��Q�{�/�KPd����}������]�_x�Ef.Y���
q�*��d#)�7����β:(#�`��D��g���n~.��%1-������ə���H��=��K�����m��v�fW�{�Ԏ����R43I�hse`�{�@#�-tڤ�;��Eӝ1�B��t��Ei9Uz����5a���JTZV�cT��\ 4�j�-����Rg� K�Ϋ���r`M���-I�0����M({#]y�$���"���Զ� �沒�(�����a��П��N�#��3v]۷�~DAP�Y�(nϐ.Stx+?�7�'|7X������\�\x_��m����1�X��rPtX�{�e�H�/��N����2�מ-V�'����=ˮ9�����No���IP�+^��`�e��nyfk�Aj�G�U�<2+}�(Ǫ�[K(}"+�V#�BB{v�����:C�M�{Ʉ����?f�ݷ�}��z1�B�C�y��ȩ���K��9��(Vdә���\)�nŚ��-�,k$���\�$�U��W`=�9��Ă*[@h2�i����x�e��a�!+s�F.QuM�*������xrIn��U���:]�p��,���A����R,�C|A��0��ګ�3Y⠜���N~h�V�ău>���<nԙl^��:�|�_xb�:�=����Ǿ��a���?I�`��A`j6��,���1���� ``�O����[���T�6Ls��EO�~����LE�j5?�1s��9ɚޙ?��/8)V,�\9�8+v�B��S��)?9��0!h�\�1F6�R5	�ww���g%�S9���Ll�̦�77���#���h=��O�u;���4�r�%�Ů�y"�S;%�W$�IR����KnC\c�F�J�KgA�{?�E֤0G%;�P}�()̚�+��K&x5���g)��k�荚�j_9KԵB�1����M��DP�S���Е���{<wk�b׊Z�*�T���Έ�	�E��S���(Ҡ��F2ZYV+�2,.[6!3�0w�E����DR-�NN���lr��qg�#����o�������-݊�KPSg���Uc���	3pNOn�D������H�$]/'b��q�LT�>���I�8[?���2{�O_�	k����'�5�1-�L��(J�LX�R{Ya!U�*K��i�9u��q�@�Ֆ3�MI�s]�?+���o�N|�K��z?��v�qA�gֹ���s()+S�?;�GFk�Y��<��U�z��Y����褉IkUMX��+l�'�?ƍ������>ê�z�ӌ�YAD�g��F�Î�Q�k��g����Ʌ1�|!Mg,-Y {~0�ρ�cf��z�+֤,��B#�
bP�Ê�[K�=�VڡI�'�'S~�W,|�����Z<��c�*/ֵs��G�C��ۊ7V��;H��C��*s�����~Oew��¬}ɪ��.�Z[��fP"���b`�Wd�jJF��yQ���`�`�\O;j�iM��[h�,gF��2�����E�(���C�������`a5�d��\�}n�[VX��E-p]A��y8����	d$��*�,aݣ�Y��O�c�,e���������"e�6�k2_��ռ��7�|�s��;SR���YiKMo{-�^̅T��o�}�@+�Z��v>9�%��R���-Zy��ad����`��c<F}�
���������GZ��n>����%ه�]�����ͼo�d^�(g��BI	��T�E��o���~w�1�j'&H�o�r4|��4��W��wp��0_�D��PVJF���v�'�;���g)���&�*?!�[�L��8�/O$Ӆb��� �G��Kg�0�'O��wr����K��W��_M��gW���	`ǂ0�l�sg�g��ۗ�����K�mΞ����o�����C_>��?�@���B�������������^���+�`N�.[��}zv.�����ﯫ�K�p&��M�k�`�ѻb���ވ0�Qa��7����i,L�Y���9]\\x&-��F��'�aEԧO��$���FL�9x0q�8/2�$d��	�"��(����bF.iɫ�o�"wGN���T��Ɗ3����ͦ�J�K�8���w��v��.r+-gYp�9�n���r<�A����Sn�61ڄt�,�LB�e��@���l7�1��Bf'Yۦy�S���@P�~�Y��L�~�)tqrJ���AO���A�ORa(2rE;[J���z�Q@�tQ���m�2�Ř��� �a���f�P1�XX�eVΤBd�[�Rd�"��Bx�	�N�͊�	'b4$�0���-��\d�g����t]���|Z��]�	�:+N)[��U���ث~��7�)�,�7���'�{%���莥��M0{3���" �(<P�����Y�}�(::2�� �������p��v��?x�|�|&dn��a�.��U,#9��(�)qdk5����i�p{{��n58츗�;��9ݞ��8��Z(i3A��L�Cbi���N��!H;�=�(�����t���+>7љ@B�-F�����՛�"�9�d2e��j��	+�����:�[�`�"�8�Y�(���="������ן���ð>�-|7�,,'����n�ok�ZP'�&�;v�\^O�}�β�@`$��d8���O��vG�gW��F(�v�-E-�/�'�.�8����r@a��?�)�_[��7��WNq9a��t�������P�I��v�{�kXJ��$b�L5tO#9��H�F~�`k��!�d/�F_�:��Ͷ�Ѓ �^bީPWa ����KF�u�)HA����!y*�Ӡ��( ��&pj��0��a
�S��*��{����w[�p�Ӭ�9���� +����c>Dl�&��|@L�h�X
�<�w9|��E�����w4����x�eS�o����� s�~(�?}mx��P��K�A����,�Pf4e�>ct�Z�j�d�`���P�t�2���r���� �x�Urx�a�Wv��M�t�,�L�@�`���1A8����Vߌs�xp���W��T`��|�/�?�9[-��q����l�u��/]^ Y�� �O�g�Q�%]�iNP`n�2JvUhl��pyqA?|�����e̿�7�MŬ1kz������_ӿ�˿���%����������������W��_�������~�;Q��S����_� ;�Qb��J���'��Z�N9ʊ$���o���.&���n'V8b�S�Y�h�
f�Xi�1Ǡ�`��mO��O�~���J��$�X@��*@���N�r�����V|�%CȠ
��f p �e��G��,�DU����M�;�h��ӂy��ľ���{�%چx��_�}�,:�8o],x��ו�?h<]���6��"`b��QM�����b�=�Z��m�d�d�v:ݻ�`�cNH@��������p^���le�>�:uř؁���^��l�s}b�ș%e6W�;C�V�W��*>d�T3���`��z�ⴻ3�����O!��:sZ�P�8ɪk�����:jc c���%�p-O!P�`��)n�w�b�\9���1wH�-(�.3S�7�~���b���>}��͐v�?%�ad:c�9��6lj0�9~E�Lx��)�,Z;!��~�D[5�Z,H��b��^�ܑ�����i�q�|oY���Nvڳ5����&�"u�Xe�A������. i����،�������\��֦K�q�;��V̻�p�5��	q��g�N��=u�I����2(��z,��
qFo_�Dae/[���C).�^Dqb8B���� ��D�`���na�%�%:�JD	v��5Ш)[27���]�c�kz>FW��\���g�KDasW'����]I�u���O`y��i;v$�{���t��N�I.i���\�`0�D,�{(�R����zG"�=>Pf��ep�zI�QQ���e���S�F�VU��.X��V.�+�K��S��iy�U֧��W��u�|%ټ��Rmp<�X���š��G5��*�ƚ��Az|�9ܕ��#֝(�-2o��^W��l^0�U� ��0D�<�
\�\��\��P��a.�j��ɿl�;�v�ᛢ���7<�3Ly��gW�{�ᠯX�U1 +���.����(�wx�R��9l�FC٫֦ecFW��f����3����}�ǘ���O+� ,pj�~D9Kս)0��Sw��]�6tzrF����������?���G!�@^��`�+z��9�\_��o^|#׾��[�Χ�\[���Z��apW�bU0��i����ǚ]��/�%�&[�|����|�"١Tx�%�53J�B��9߼|Aϟ?ײ�齋�a����]����իW���g��ܺ�zF�S}�'r�"�� <L����B�i��[Y�캲�}h�DS�1AsF�I���)W9�gT�G3QY)󽂓�ն��ͮ�>��o�����[]������;AAx�������|׉?�u��t����3�;�@V-�+g������"�����VQ��So�օX<c��Q���:ܱ0���	�E�&d��Nlr���)e��;�+
+���f��1���,��	b�5c���X��`�o����g�݂��R4�R�:NL��©�~���v�����;ӽ�1�Z��Z^g���F�P~�`��a�g�:���d#Q�8�[]�����.����_P�$�q��nX|a�;�{Uh�#"d���[g�Mq@Z���
V����4SO�xj*l�z��ԍ��߭f��`��|/s�i
���4� ƥ���촂-��bem^�,4BH��p?	�ǊIsՠ�Rl>��D�U�%}�nw'���f���8v�-��Yqĉ�����*X��Z�Y(]PdAy0e�u�pg�AB�s������a�Lr=M�:mBi2G�B����R���~:D���
\�� ��c��ʁ�ˁ�k�(Ð��\�y��ė��x��2*�z�#u+W>$b�=��t���8oMYh�ܰ���&��y��6Q	w�G�]�f��ZŮ��u�.Xs�)fQ�q8a��@+�F�]�.7����wJ�6Gf�X|��@eL �x��uh�[��5R���\�o��A_�����NT���\2�"���r<7���8�m,��5eph��~šC�y^��пٕ����P2b�(5��y4��2�xSj����R�Y,�� {�-J�K;�Q�����QZ�������5Ɋ�oV�ף��T��:�N�)W�PɌc�S��m�E�ߤ�_怲 s�2��U \͸�IST�p�}V��6[?�"6� ��9ee����eD�J�>Лׯ�,���ӳ�7��XY��['����d�X��܈k����P�cU0P�	�>�i�dd�߅��ܳ���Ŋ���;�������ǩ��kK���#����������tz�c��"��g����8�
�A�޽�A�ع��������������./.E)&�a6_b*\B�\L}�ѼX���,'����̀wt���D��w�Cq�6�u�f)*��m1nW��.�σ�9�>~7�I�B��J9z�	zЮ���6�ˉ�(F�5��	����`�;|��Օ	R[3��]��s��L�-�jo�ޟ�fʌtM`ۈ�CL��r ��/�����~�E��_(u��U�����[�i�`��5���I��ad�m:�=R�y�������{�3Ti�l�)LL �=���/�[gزBv��QIr3��%��9��1��g��:��ٖ��m�-q�Y�죟F�8����%e������.g�I�d��d5�A1f5��|N��!X3��+����}�qIJ��3��9�So���ն&�L�ҝq��?����1w�E/�W|�v4�.�%���-cE�3h
 aѓ$7ٟܸ�2P5{�J%�n6��;e�#A���}.b������H'��Dhe)C���U�SM�L֜'{���z8O��|�}}�+��O���ZU��'iV��-��Z����~�����b�t�1��r�����`����-q�łX�V�m�~�t�EY�E���.P ��F����n9>�ݟ��C�}��~�p���1��ndk��蠔k9N�.�>��q'KA�JZ�Ҍ���LS���1�f����+�f��<��!J�Dsu-�\lo<N<J �����;�&<����ag�<7k��Y�k��F4��`�f�a?̧��kX�v˦���ٖ�xPJ�3N�~�������<�����'+v���g/��<Y��CA[��29�X@52�~][މ������h�54�u���k/�${v*J�����7�7�ޠ>�bB|r-L+v�MVz�����o߼�8&�S}����wֶT9�1vد_L�u��Dj����r?�gs�����-���ҧϟ���w*8t������ufp��]��>�H��ݞNNO���݊5�<al�Ì���0U��ň��{..�����d��SQ~��5��<ud��T�|�Ȣ�y\��R%��+��!�`f��������ػ�AK�lΈ(�|��`D���ﳉPRsl��[� ;�3�p��j��9��n����J�t�t���ņ�;�`EC��cfzGe�+:�\� m�pF�b���&u��m0]I8���BVc��s�-8�&�}���X A	i�KR4�"�+it�b��Z����$�Q�U�#�D�z��Y�� ��\2̡���f�;9{v^���n��-��l�-�X�/�wԵo�X�t��c\��Ū8o����'��=9�p۩��`��ޅP�����\7`N�
�v�X�r�Q2�k�-\Z�YX i�7�֑LD��r+T��[��-�e�����<v�����D�0�����̥r�Lֆ�S�cc�sF�+�d���_�BRi�5^�]���ǻQz�A}òG3k�u%X�b�j�4���+�r��2!VZ莧g���S���,�������VK`2�[�A,�%�zz|�<�2��_��G�ȸO5�j0�E�\�8���Bnc'�Wτ���=\��=�#+����om5d�*��3YY���<V���\��u㺅�7�jW�iui_ �F�vk�ZJ��Gin������a"YI�)K#�<�Wγ(�B6���pSήKK癠�[Tv����|O��S8�L�D�(��@�-�{�;�h;܉k<��-�?[�}���_�;�9 KG�Ӱ����e��}���(���x-�of-ec�b^p�^��{���V�5�ҵS�� v��O�<�NB�ڑr�ꌝ.�^���p���
�A(x_
�����@9��;K�z:!zl�Ç�ai����ĉ��-8͙SC0u��
D��掗����RW�h��0�M�Q�Rb1C��z@h�[��Ȉ�c8���-;��f�L�Y���G���pb�9�����&!�/����M�2�7�#�2h㺯՝`�l��E� ,v	3����2��3�	 r�:hJ�ݮ%�?3Hwww�@�#끹}�f:��a���(`� &J*��5����z�gBjU%���
	�ಗ��L��
p�1V�--���%o����U��B���Pӭ2�^�lV�#)K����A!vTP�+�`�sV��S�97�Z�M0w�U����x�=�[�kR%ǈ�$[���hd�M̕2w�)�pO����oiy�C��|�櫽���f�����y̢��s�㙕U	�#-g���[9�mj���U,V]
$�ǌyg���ʣ��#
f{m���C%�6Xlŝ��fI��"�6�{��M��~����E;�ױe�F܏����VH�����4",��G3��N��~tw@X�_�Zk*�(�X�
-�l��Hՠ�(v������kAHRQ�M���[?��ٴ
AC0��W찢���*9���8���i�)��&����2�,|)�u�#����׬~�E]�����Ć  �����E�Uɔ=��ڛՒ+_:�?��96w��H ���]R4�V�\�ͬn��]M�3��r:rΰ%'�T-��	�s�4�^ƙ���ŭ�WWP\��hEq^f)ֈ�p��T�@�r���'��t�n'������G���v��̻��>�C�f+�&�#��*��_4l���X�i�^xv��]�p�LGg5���Ú���F��B��湒)���g֘�m�=��{XtK|Y	���\6D[�i�(D��R|I�+�q�~��w͔:QO�}m׺���^M�����	U`�b9J;�ج���%_�*β�5��q>��%3�pK�j��ݹ�͜/@�3����ܰ,�����c��#k�=�+zj_�8$h*x߰��/���JM�����1v����0c�3.� \[ր�-�I��r��l�J�N3}�}M��
����'z��.�.���?�2������$�|��Jqך��lQ��ݟ����d��������$����8-���`" <CHH��[�����F� ��g:���v�vw���(��98ɸ�����ߋR���
*�+.U3��9#����P��Ƙ~Ĭ<&3���^����$�:E�8m.�+h��#8׊ō�A�;	�8�:'���� lZ����9���eAp�ࠖOf&��L���b,GP�3QJ�9���df���n���j�M�`y�ʝ�i�L�lx	�;���2��%��3�:�ư��9��>�ŕ1],�$��fE�C`�<�rB��Y}]w��؅%��mX%���[��P㺖�+�{�5���� �Y��oQ�TM��Џb�%��8��Ǧj�����V���=�T�D������Wt/Z�S���p``��Szu����@�.YN߱5����Ս�����Ǡ�)=/K� �0�b'Y� RUk.?Q�)S��b��l��Ic�3��,<T����l�i�XJ���D�R�c����B�%�YfD��M�A�3D$!��Y�x�s>�G�6�fgq�`Q�G�� �|k A&/{�GULJW�b�����O��'J+��6v�v�F&/d%�ˁ��20uN�\A��yh��mw�����ǖ>������u��O�c��A�!lW�<�v��|�i7׷r4N���Z�6�C5_�:�<$���Q�O��'w����[U����*F������X�F!9/.\'�InF�J�\�G�"��������KM;~�����-3+���ӫv0�
�aP&J�K�ay���?�C��ĭz����X�d8��ͼ�!nk�����}�/"(�s�~�����51f2�H������C�k��X�"j�������_5�Rg�sv�ov�?�%[&�N�ݚ,��\3o8�qZ�C��x>�n&$����� J���7y��#��Z�B��)+늝��y"YB}�3ym����]�'�������8g؀�*e��#�]��;~���Ъb�h,���3��y��5]\^�	��?|/1i8����kAt�l�sww�R����򹽹��I��"̿�!�������y"����"�ݬnnn'&~�XA���ޚ�+wpz��LW{%~�_�L����
J�wzJ�i�9���ܰ҈]�.�/�ŋ��+�xL���Vg`Dqkm=f'��U]����At�/T�&8v|�����-G� ��o)���CMS��J���zgL���ց���Z밥�pCl/�)�/8��	]N��9�JH,%�_�LD��)�D(=q�Cs���Uɂ5ةmW4ͭ�E���pY��ToQW#�?�s��Ԇt?�1N�B��i΍�Fzl:J�8�i��2����Κ	nV�>�p���8�sZ��(V��p�[vA#p.ղ��0]���!��C.M&,(bG�9Yf;�xuNs���^�x�	fwCU����ո[g i�GS����J�y�X�f>)vL:%��S�.y1��^����e���*
�έHe9͍���Џ�\�F�Jq�5�h�G��U��ag�u��Pa+�I��Ji�Zl���!�vb��<��;��-��ܘ�Of0m�Y���,$�Р�^��&lj�7c��]�k����Tجu58�C�!����BR��Ϥ��d�W��e�1�����û6�D࣒�,Y_䷊��	]���]q�g�͢�k�sUx�;���/� �f]��.%ܿ��K;�ҳ���Ff5���~f1��
FЁ��]�A�Ngf^U�.a"Lq��gJ+O��㰴#�LsZ��d�������U��"׳�� %�ޭ#�'��:�J�����漋�H}\QR�����s	E(*�9�龷[ʌ���ѹ�~����+����6�}͸��ژ�K3Ay���T"�w�� RY��4<	k�l�d$��]��E��n��ղU��)I��sP�Wn�Z��#���8^�"-�P�������ΏeE`R��r������Ǐ,v������PW��@��&���/#��z�����s�p8euf!����[�!���j��Z���b�5F�1�-���܇Y96�.�&a���7�t��і^~�R҂�|��(O�Qd�W�_��7o%��珟D9r{s#�p �+Ζ���X��ɱ�#�����F�`����b�<1>w�0z���?�@Ϟ����s:;=��[���7��1%[����Gv���^ݩ�ib"f�vbut+ʢ�k��gϞ�B�ﾓ�ɧ�Sa�xll���s���ӓS�� gir!���1g��-�,h��`��$<�:&�Un�Ê�������S��c��'�ʱG+��C"ܙ�SY��N��(�iL;u��lv��O[lb���i/�uO�\��������wΨ����mQ��!FF>w7���)�0����'��@�,dK�-�ł��^����KS��ț�.itjw+�9��׫�V���Z\ڶ�Ş�K5��CXI]�F's4�B�fvzY�����T��`�Ä����hr-�$�7�J�2�II�Z)N�Ȳ�tFY�7ht�>�;X:�A�Tz ���}�;=s��ю��׌m$n|d�J�mV^�{��v�\LH���N�D�H��'�P�d�I�kK%�F�g��f�ra���:��0�n��k��
)�$]	�S�8�Ւ��)�d�Y�ɸ8�?����SW��t� T4rX����ĭ��tX_3�������x��߈���K���'�(�Y����]f�1n��}�w�N�|7n4|7�w�Vv<z��s��B����w�K9�XgQ87Z���) �٤�=�/���,������c� ��@A\��eZ���_gYG��wI�XmuZ��cS%�R?r&��p��}�a>�j�j����js�$)͉�:��V#�gjK; �}�F��	]�<@�^k�����ms����v�jd��/pM��΂��U����&ƦE�WҦ ���I
B�G6g�l�ݼ wq?�O�RЅ�[�w�M�D��#�]������~m�չ��0V��)�5����2�����] �\�9L�Ao�)P�L4/We�B�n,2Os����/G��KY��a���?�5�p)�>����1���J@0���C������g�:d���t��/���;3��P,����iV�O��z��')?v���pS�M��V�E�)!����r��W#ƽi�����t���>�H���W	�'��'s��ۜ�����$X�xU�(vД����s�~P�h:���smp,ƨ��{e������Ǐ���:ٜг�����3!D���1_�v�%��;i�ӧ�b�Sʵ(s��h'�f�w��/��U���7��vj�߹��E�W��-�8��vI��	F8���1�w�|s��pB���I�}�E&k6e�ۼd���ڃ'p�-�Gˑ{|�9�3B�5����.��h���{QO-�� Lx����2e���|9��Eϩ��L�n8+���)C��(L�u��,���!�O���P�:��D�����]����\L��TX0����D�O��Q<F���i�B�:���������]x����YiԚ+��ԣ4s�x����� ^��x(.�2Y�]��P�{'��q�i���x�GVH����s��Yӻ{�3�f��~bbX^��ԩ*�@����X�K�qk�b]�.��YM#�oc�|]}.(-hm�`�@�f���b�eQ�0��b�ٹ�NRݚe�c�ᦦ¶>�D������%xr��k�������o�`98�h�} ��X�?2%2+��潄���T�u_�B�S=�P�]�М�#� �/陱��G4��%���@��|��0p�3�K�N�f� ��+�\:�/��@� ��k
_]��ק�3��B�^���-��L�Z4@6U������zif�$�5�$����,oL0u��bG]�l�sjs�w��$h�ܵo�GJS�rmJ�3�������
�̽��]�O����U��T	
U[�<^�ҹ<	܄g:K4R��2ݛ+vJ�W�\u�/*	f�u��X	�����ơ]�Oߏ��3�J����V�V�����:Rʁ�1�P��t����
r��،��8֧���J �-n�騳*�y���?g�o�_��O�����a��g����P�̕a�0Tb�jp)? ���a����/Z�@���<����W)��3��3Z�7�Q�����L���K��(��컟�5-1̒���_������/7��+U��$잜���3Q�\�_�3N~vF�6�X������h�zZ��Ʉ��6/�I�}�XU�^߈���~��R��tzz&8�ykk�,��?{&��O}|���˟�Do߾���|�+�X�t1���o�����^���m���\�����͛7ӻo%P�`>�r��Ef�͘��U���̜e[�Ϙ�9@��
���[�v�|5
<̞��O�UX��W\�U��77��D����;�*3�;ږ�N�u>�`��O��{�I�F�J,�x �0g�@�6������o���6�\�}G�^�=��.F<�T^��[A�� ˗�yi��ݼ����S�b��?@6)l7�	p0>�1ޯ	�-�3��7&]�F��I����vD�7~
�l�j� ]��s��}�@���ߥ�V�$�5�����N�V����;Q�rBx�s�G8�V�w{��XG(t2S'ܰ ��D��!�6g6�}����MY��gB��D0���5��h�2(M ����|�u�	Y�J���p>D��r�vDmW�ъ��7q�e�*��:;?�h�eryK�G��1"Ô�ɝ�]Į��x�m��݅�j0�zŲ$�� c+ŭY�9M��{�j{*"�T8�����3�-�d�A,��ieS��Ɲ�^Q_��(!��˰{uw�#�.7�=�ٵbu�.�/���%p��Ų��!�a���#�476`'B���m� f���c��9�:�]�1�_Tck��zG�i�xgGD�Z�kƥ�:�ג���<�b�X���(E���aeV�����R )U�F&}���m��%dLm(��,Pz�Oȼ��6q�H3%N)i�m^�3�O�̺�ٶB�� �vC�k�:�`�;�Ҕh�d��q��s$|�C�>\�~(�vK�a��(�0δO����N���4�e7��R���S�>X�D��n��4����U�|�b��a��kc,yಸ��R3�^N���V9��E��9�z�%��+!��nE'8���{��5\kMD����J�Ob��O��������sw�=-h���^k�^����/�ߣf�zYz["g��tb+���qr\��>�_��g	�Ɍ+QX��1h�JfCϟ?�t�l��ʢ���Iztv[:?���Eu�t� �`P�l0[6וb�U5E����O�ǉ鹡�>I�dt̩�����}v�8���@l��qs,|)��O�x<wҧ�gW���/_ҋ:�|�$c��5}x�~b�>�"H׍���y
B�9S�0�x�`�V���A\T�4 �^�#�St��D�g&|�!'�_Q�n~;�1J�ׅ)0�#?�7u?�l	a��T	y7��k�nb�8�4[�Op~�و��v�f�D�'=ŗX���p�9̺$�\gA��i�>��60�C׺�ue�1v�,ښ���a�,1�z#�rGM�(�>o����y�2�\��AM)mv3y"�f���#��Oڵ�WlR�51�6�n�`���e�[�cʝf�b�ލ3��C]�=J�V[�� �l�#�l�3�r(��օ��:D�������B h2��51��e����`��|x&���ގ:��=S���E����r#�c�{[i�"qDp��p<�T�Bi�����x�x=�ڕlw�S�aa��s����	�G�uK�X�>PYmw��wtw'u��e�S�Z�5��p��P��@�j���pE�Fwu$��"�d�Cqf��ȳdО���~j�:�s�u�]�^Ӛv^���%��\�����h�������+�V�ΕN1#@���c�gs��\g�ԔQ�R@/�����\�����m��H4��T��p~�u�lv]k1�4�$�MZ��μ��7K�`А�%���Fa�b��=XBi�(Q��Y�r���quHmv6��&f������
���!�Q6��`b�}�^�d�g���Ĥ��ʟ���8w��7�ܒsg �>�D��hd�?wٗ%ޅ�f/���ZY���Ȼ����8^���{��Ϫ�����ڮ�a~T��"�r�V�x� чl����$<�����wd<|TV,����Yj���ʌ��{+�<ן�{u��dęJs)!�c�'-�"0])8}���e�o���	ǌ9=w�+?X����k���XĜlO�D���.��߼|I������ﾥ��SQ������ǌ�0|��n�L{t9�_y_`ͣN���K��S���l�<~v&��w�B�cQ��_�@�>{���߽�9�X&�������?� V=��e���7o�Y͖:�pI�w;-��A�;�y<cS�0�>/Q~n���rEQ�ז�0��C�G~4+
2mD_���,ǹ�k% ��G+�bӻ�e��%p�Mcb���/���8���IG�3��ݫ	��r��g���#|=є��\Y��C����h~�{	Ժ�SN�@V����%)@*S��g��(*��
���:���Y����VcCP]�ZRU�r�h�,Oz2SUH�����6?�J79��biJ�OsA�C #'�>/�`�%����6��2{�T�b�(��>�3��t�Ni0�EO7���g���Lغ�	>�;����*��_$ 5[��bD��2ap��Bjy�dr�'�U-�8�jW	�5����\�嘣� ���+2���E�`�%�-z�J=��`XC�F��([�X�Zdsr���_��;���<^�OB�jI�9P8�MD<X�F��,���P|}"]�(v6[aN�aonև1!+�������s��a�@+��{Ґ*����Fܦ$d����l�g6O�v��rh|�藅h�R�)p\����-u"O�
�L��
{s�$�z߳�����|�6�`t�gX`�u�5 Ҳ#+}�sȧ�=+t&����b���'�w��t�Ǯ`�b
&2��??�4swG��5�� �����R�3���{8�.5�+#�F�s�}�Į$*�>�q�R��dΒ�KJ�/����YW��|�a5麎p�
<�����t���n^��l��0�z(�bޑA}�A���AC{�ʏa���q��U�b9}8P�:s3�V�Jw%�[N;��+=1���<T��!6Y,@Ko�O���h1�<�"�
�S��h�ށB�
t���d�Y��u���D����˱.g:>w�w9��kR�|nߓ�s����Q��������6�jz���oS��Z��ǂ��q�k	��_W��w֩Z6��KP���Ǘ����ś��I�=9;��$��=R�j	�w:	����ffY�#��[Q��;�9�L+z�|�"�2�}��	9f�R͈5��7���� b)��f���A��k�Xm%(��Ds'��0CHa.ʧ�[����Z��ӯ~��a+��a�-�v�������/�q���R������Z�>J̠0M�T�� ��icm�kN+�fĘNj��V`�ր��)O�E"��`�b�1�.K�o��4�&\e&�ʾ� �5�ѵ�l�\ ��(�%�L�y��P�^�؜ѳ�3���݈R�ŠZDyGl�)�H<�x`����Dӑ�f�Rw,dQ�Æ����qaμ �ΰ�CM۵LZ�́{���o~�-��������}�l�h˻�9#���ln�ڏl\�ۃ%ǵF��P�8�_0������&G;x���%�v�3�~��I�3z<r&�遛ir���t�+��"�-_@J��$_���p�����h�p��<=)���x��f�4��p�53wl) !ǋ�Fk��߱~�� =�^���&����|����p5�1K'�Ŕ�}�g;�Rj�E�|o3h܂3���sl�Kro��aAH�Eԣ�zǴ���a9^��fY��:��n��v	�����co1�evY6>�hS.�E	��P�V����$��+)L����+=�
L��$ ��X����M���ꖻ���)v��4��>�csdcB���:�p~.	$.�/��"D\}_a/��Nf��hE�f������ķ�\ ӬXf�hn/P@�5b1\��
M�>�����b2��ʤB��A+��
?څB%[�B�cB�"K��d㱩w�L�K�X�ܔhwѶU촆<�|�����[N�?��(@�SA@�m�U�t`�� <�&+vJ�`�M�Y׊�3��h>�,¼UCy� ��Vz���싼�����Opȇ�,?�\r���,�U���T[�V��^+h�6^=Ƭ=�������C�3�G9*��B�?�68����L���@V�
=��	�mE��+Dט�������%��׍o�yhJ�^��
4���p)���D����{_?��
���ߋ��(vz�u3H���Om�uIbל��Ӎ,����vsJC$@2��}��E�H�lT�È�ӊ���=����I��ӭ7�V��0ӝ5i�,N1�^G�/��J���.�.$K[�|��Y��}bk��4����~�J��Թ�������u�|y�ʨo���� ���?���?�C2 �[g:' Z�mX!�0�9�@Z��%��j�rg~Rw��"v����dSRs�O.ˢ�9!I �|ݏ 4���)]��	Z�:�c���b��$�Ն�H�t�.�]M0���L�u.��*�q�ʡ�`���NXJ"����	�	\��%eu'i�O6��!�+9��K<�Tg�^��cX�����)+8le�3D��W�rA���l
+v�\� ��읚��T�T电wU���o�`d�:����T�S�L�S��4��=?�d�L��ו�g=�~�	5y&�oI��Y����z�>��|V|�%��z!�<lˆ*�g��β��ZV,����Dƀc�5Po8�d=�4WG���m�3�e>Ӏ��Nؕ9V��l2�(�P�kQ�q0���Gw��uhD���E(N���γ����m>���q�
^xJ����
̃B�Z�ˢ^�z[�۬$�Y�/�I-֥��\�+�8�1�F0&X���X�@�5,�4�M�R�$����V4|{h�E)�'+��s�\�4�p����7����-n+y��r-��*�6���bTi�4Ӎ��\S�]ĸ���d�N|�}ݫ5��Km�ן���[l<�~�57�_/tO��g>�X��_ʁ��"́2%�jem��Q#J~g(��'���;��kC8�/�j�xBb���g�1����<�Q�&�+by�7%Y�E?
��vh��1�^�]� Sy�g�d@K�of]�yz3�e�:���l������TC�nR�;k��
��}K�{�2�j2��'��%�%�v"f�.A;�/��z��^}���^{}�F�z���Ŷ87��0�Q��aE�����E����"w��1�v&;����`Ѻ���9�?���8:ܯ�Y�+�>���SxVos^�ǨO�Nq��&�A��je.��G���+��
_���_2�w�]�	�i���S����4�樖�7"�������\ ���1+ee.2.n�JmHUܚ���Ŋ�ėO����~�G�����@��ʕ/����$��|<�an5�9���.`[����N���7�o����X�7߼�F��{�N���>��GܴH�>��no5��ׯ�O�����3+�g���;\9����[����zz#�F/$[���y����y���� h�+d
�֤�kk�#lMˑ`JSj�n��gq���hI���kq��B�b.����ħ�#c�ӳ�XӾ�)����O=���F���v%x�H=��2��O�=9��Ջ+��ꌾ9������bk'�����w�,u�]�o��C�f�$��J'S��vCg��m�Q�0�uzb�)��ॵq�~27���`��f�Ŝ������ +uX�C&�$L[W%�'��̛*�4�P03�b���4�a�B(�:��l^�:�SbM���m����0�к��iO^�g ��TX��9/���q���ǝZ)N��; �v�e��m5�~:ku��I��-Y��ZA�iE� �K�i��</��m��:�R,�OW�Wa��� ��ڹ@���O��R�q���I�N�+�Ȅp�\dFi�x��2o�G�z�ZK�w����T�EXp���-M!S��pڹ�?0���5p�W$�jqT"вtI��2)�pl^{���d\����I'��CqU0*Qg{���Tw��O>[��J��?Sr���O�� ��������,�?��Ze�D)�JJ�1_;�Oh;nE��]�����Ջ{4�����Q0�� N�O$~���]^��ٳ��8�ʣ��U^��<����;�6R|��;%�%����b隀���T��d̬'�-Q��T���:���j��Ԫ����>,�T��#��b-�
sǁ�}3�x��g����6Y4��waBy� 1��JZ�G�F���f<��1���xE��#���Ȩ;O#�q>�]��I�b-������\�er������aP����
��ݻg Y�3���������[�p���~��Nh�,2�jI���{z��}��>�,�G��ņ.�>*>))��OX2i��|�9����r�<@i�~t7�_,8r�K
Н�*�n�g�����J^�Z���Kul���/ن��)u�y����x�X=q4����W��ǔ�N8��!�8_���3=p���b�;�:Mt�
�8%n��73���ʵ<1�9*�@89��X'��Xnon�p�:&6�ܟ�xN�����~8�@��]�3U𻆟4����-��ވ��qvq>}?���aDF��N�/;>�,�VS���3ɾ���=+���ܲ2P���'ל	�O�~�ߊu��w�D���9i��J�OH������~��^<A�g���saZ���;!D����+�\_�������pJ�[VfM��6��ߋ҉3V����7�%x)g��7�G�Q�0�P�������ŇEG9ͭf!�\�0ȹ6��a�-�*2y��cVCc]�xn혱Nl�#6���'W8���g�W����ijS�[��r����̂[�7L�)���kB�w�>�w������o雳�.&p�Mp9Nk}*���0]�b��涒�G:�ĥ��M �R&��S����]�D��u��_c�QtM\�J8�!Lb<�Y3$ax��uJ�©b� ����H��4/��3\�p	)�$w�2&�M�%Å����z��Kӟ%����*���\Jܼ?1�2/}3$�+�(qj��!��Y1��D'U�?1�'�|���	���f��b.7%Bl��3djmh���J\d�����ę.��E	�0�y���gm�����{X�mg���9�M�Ժjn2߆�Uw4�vk<�9۔�ܤz2�B3i�T L��t�dZ�� ��GDvp�z���Xi�&$�wQlP��PD�=�7F�b�'%���¯��>#]�ט7}�,�����)1�
'w�ہ��G�r�P̂@�F�y �����)vN�|F>�ʢ���o��b�aQ�i�mpN�ZL�ޭ��o�J+�&: ��YP��_�n����N\|��A��4����Φ��k������r�(.�(�-�C�+��3_Ö�z0�2̇�6�X ?��Y�����`��t˘�výg�`⅃<o��S�-e�����e�g�6we�Yx�rED��5J�|V�K�pd9P���5S�
Q�L���|4���,C���k���ձ�W]�-�k�";u�	�8�&���@�c�6K��M@љ��מj��cj�jVFq��5ccߩ�J��uA���.�N]Ѥ$�7dV�ɻ�*�*gt���b�����^�<�,� �@!6&�b���Yǂ4�A�����b�Z�$���3��3���奬[����������!�7��o]�]M���iLM���u���Q�W��%!9�)�ȏ|O���G�����X�Bo����#���+V��Y�W.�	ں`$f(3yjv���?�����~��<��CH%8�c������r�k�+�@�a�K�gI�կ���45S���ҙ�Jh�8�=I�iȒ��ń��}�� �I�e˖��N�4d'9�+Z^~����r�bQ��
��b��FPw�� {zr&���q"��vJ���tj�r��O�?Nu~%�E��p
w���K\�q"�liî[�tuu)�٪g��U�3*�E����W���>^�a�L��>���bbř�6����S�yL��^��c���ز+]B^�,32Ae�t��+��mzO��@�'�|�0��A�׫
!=[��.EKan:#2����z���v���nOr��
�#8�h���{��If,֨qƫ�i�S����\�:딠s�;v1b�ɠ���R�+6AF��jNB&ri�%�5�?]5w%�xZuk�0~Z�W?l��<EeyWT�cJ��N��9��U�-֤��5K��$f
ϪA`M�I5aX3Yqmy��q
�#���a�2�<Z�ww�!U$��P�I��G��d�Gd0����s\�rkPA��qN�:�۝��NV���͍q������:��ҿ�o��b������pKw�H��iTW��K�\�UH�73��>�E��5L�>���V�8 ؙ�%g c,aF��6rl�p��{l��X�u�5;DT����4�1�,��邛(�H���J�U<����}l�[Z���f=��J╚
b�H��
���~l�~i��ݪs�� (��Ѵe�_0�$��c�����q���`���y�~	�[\�����W;��)��K@���-DH>�x�pfΡ�C�^��/z�H�f��-\q\��S�\U�#���G$�W'��������m�a7x*�R����:,��JR��r_8��h�C�S���9�r*�c��W��Q����% D\7kM���L�j�P&^�ܻRJ-�- ��U�!��L��Q���l?���q݊K�~�)up�gg��_:*����m\q�q��1D�Ar_񍌯*JCm�  �=ߙ"T]Q���d��3~u�P��!R������+9��Z�\$��)+�
��eT'b�w?
�
̳���t�q��f��͍�609��n��y�b�iEeV=,�l:=�=;�8��nCW���T�+q���V�����u�u�ң��c^�I����S�T�W�ч�k�?~DO��x0xrެ�N�X\ �ec?�b+?!��c�v2lek��դ�pH�d��k����]��v�A��Uҗs<�	qܜ��s:�=[�����j���bǧ���=��w�������law&�H�֚-pJ��h�vu}}#�z�rp��K�}fI%.BHٌ�ӗ��v���Ϧg���ʻ������o�H=�	��_K��ruq%A�����?�J�pvvF?}���N4HyB��$bf��v��=� h� �����JuaS�@\�8��>���ժ�&<�Dd�O�� ���~�-ɔ��\'�A��b��8���;6��r�6�e���2�x:N�)P�'*�qo�Z?�8OOΟ
j�%ɇ��Y�5��v��϶Eb윰�C��\��V�T�@��ߪ%�R���ʳBn�/�Y�@�Uc�N�?ML!���&(/�ipZeI{1��~�`K0�.�Ǩ�X;�9怨ś�<�<n�U�7��/ƉPLh�F�>QTab翪 L�ZtώC����΃dt� ��YR��)8ǅ�I� Yrn�c�ǂ9���"s�"p;d�t�4(��@�5q��ת'�f��
�\���v}m�a�%�ϑ�1��`4*
��X%Z?9���t�>L���Aa�ܥ�ܫ5�߄0Y����yLn.��ʏz~׶`V����J��j��Y���$@�m�rײ���f�S@�l0��ԯbb�
�&U�H�d^��\?pL�V:M�V3{����*k|�̌�bcp˴���w�nc�
�w? f`�%��B�i8���B.Il+^;�"�X�2�Y�jn�$U��Ca͢�"�2iX���ž���7�(�
c�,��.[���-�)'��n�����K�u^�+dE���ωYh�>�� (��/5h
�2�R>�pfS�Ro�
�v�%Xq�a���F\��vx����x�d{;D,��bs�`c�oo�*�Yl-¼�jwC'�QdM۔^������y�:x�dd��q ]�?�h�2%��D'��ggm����>�h1b)���z�����h���H��q3�As��.[i�7��,@�<b�$�2ي��0X�o��K���iμ��K����[�L�뙇>��ׂ�a���a"FK�����V�s E�M�'��_�RUM�����(vN��?Q���x?�����gz����d.ԏ��*S�:�F����B��0+�����2G��:�NS���f�d�Q���m:�6NAW�:�
�Xԟ��}�^��+�Z^з�J�Z=<����T[#M��z0���#�csL�.�e��膳`mOĚ�8���d�i�A@�X����p1R{��}��Aܒ�t���������Ӊ��F�2_�xf*6KeǦ���)� wyB܌��X��\�Ԉ�.[뼜������޹�̸�	4[�������?�i��FLh�a��oK���b��s!�)��/�/�1����dSk'v�ؙ)rgi����o��5>���qF0"7��2�yg4~9M��A���c�>y���9�F�����b�I�>h���|C�8��t��#���a�`h�S"��߉&g3�=3|2TE`fw6&{R���2��O��$5	C`̢���P��H����f�z�|�:��v0k��\�q��/2�Md�Y�FI$2�e*	��]�c_�kI�G�����VDӽ�8w�,�rNn���)v��Cx����R6)��~e�-A�u���j(��څA�+���Op:�)iQ�Nw�n{���QRx"�{�]g.�&Wi��A���L����ŷC���YSkJ�	��~:�YC���V7dm	{g�xj�]($B)��\�F,��+�R��A'҅�t��
5]��Y/W����^�Յ������H����P���d�I����,L��HJ�Csp�ԙ�Ǹ�̚UKgB�3���s��%r��ě5]D�%�B����;���GY�.�⊢�_0w��"D�|�U�k��p����q�x�,�´Oo�;�oV1�r�V��*�)����@���>~�$�B����!�Ѝr@�1��ot�x���X�dQ��ŉ���w�����B^\\H�E9Ԙ��^�Зk�a�}���f�<֕��	,�`��[|��2�"�+	������~(X�1��G�]^	ߊ��&+�޽O�?~��C= D0|V�1�fU*<���VbrY}�}ouc�d�/��E����M$J^s��߉5:x���F�Y���w$V6���~�2��]}�����@�(?̇��S�:=We���u;�)_n����V�\o�j&;HT�&���r��r/A�G�����4_��;���鉌}�̼��'g�;۩[�Ѯ���J��
��e��R�t��s>̮�no�VQl��<��qX��Ӈ�+�Η>^�CF�ř!���3������b���14k��_��2?�q��k�/R֘�<�ܚ�"��=$L���K��ϟ��Dx�t�OJ~�t�@�6 &���]k+���O����`��[��������g�D��JQ��g���OU��F�t���i�Qb��Z���Sr��+[�̊����i����DO�Z��83�g�������%Q!A�|�ӵ3���׿���y����Ql����%��^L�5P��Z��	��w�;M�V_,g:=��c���덑fB+��f^~��U��'�3x;ݜNsr.�`�i�q�f.k�΅��ĸq�Z��W��ӈ�Ed�7�K��|���o,�� '���^,��Nz������ȱ��A�WD���X��N���l�A�jE���XaeQ1�	$�Q�3�Ŭ�%V>@P殇5F� }�sdF=pr"��<�91}�g�Z��)�P�R�O�?�����g�^�H:�$Z(L�k� 3��h�#O@N	�c��Nª1��X�C��T���Z �!�s�>�2v0��i ���'|ͮgݰwX#���Q�D���r�Z�b����k����x|] ��c�s`��`'�<PK���W�<�a�)E��(�~,��2gn*ֆ+E�B�:�5�t�?�]�-��%�6�ʈ`��)�F3��^����-���*x�?��P�$�!�9 �ݴ����b���b����P�l���J���P�����D�xw�"�����߶>�����~7�^L��� �ⰹ�\�<��ti]��������K`� ߫�j��0�;�o��̼ݧϟ�*��G�NP7�:�>�c��>	ʇ�xV�;������*:����������,�8+ ޾K}��޾{+�E�!����ꊦj���e�
E�*y�+��-_�X�c�>Õk�K7����5��T!p�=��}~��#���+z5}�B�c0��d8���פ�I����V�c1�dm�]
��q7�5����Tu��@����L<��/�Di�
��f8�~�V2���*,	?kW4�(��84O;��
5�_)P3+KX����������Lx��3��v=��	.�}� t��5O����,A�/Rq�	�����#w,����^쀤�<�b�~���8O��g%[j��$L���^�7���d��q���Z~)��x�q8�Y����P��U�@`��V��1�S���;?T|�b�?��*�42��=Bs�w����䌡	#z�j���yw��3Cļ���,5����c�	-#ӏ�?���GɈ�Z�Oag�v~q!�9L����QN ؊��y��W��X�ӭ�hf�@҄O���۷T����n���r P�� f��T��āݧ޾}7!�?�����:L��η�7��Q�|"���˾|�L�I�=Oąj#
�{���W�� �󵛩V�~�޽{O�S?"��N8��Ǫ�%���m����8�B�llbM 
�V�8ى����m<@\5��`X��K��KbQ2�U[���^M�Gu4��SUR{��
��|��O۳��oe���A����~Z��yo$����7�XL�dy_j��~F$�J��	h��~��\�媾�`$�����e±{5݃1�1���f$,�ZVc�,=ꦇPb�'QĆ�u�{k�mi�Y
�+/��'��K�d�ɬ1�X�"l0Rj�?�i���?{o�%9�[�H�Ǿ�Y-�խ~��;f�Û3��F��Zs����I^ f��GFfU�J��,��p��fF3p\l ;������
�����Fk�H�+���W��#����KV*�i�q0�Q~1���� �F��	,����Uߌc'{�N�D��+��F�HI��y�c�_<ʍ�㛡�U'�����#@����s�OrS��Eg� 9�JU(ͨ�a�7�ߎ~M�cDrԒL�q��՘�S]�ʔOe�Ft���+��)_4��_��9�m�\�a��0��hz�I$V��ؑr��s�OK4Ύ��pC^s�U����"�=�F �wk���)�x�TGͷ�jn+K��й�w[�-Ѧz�����A�@�Fk����sX� �	�XY������Us'�u��j�+MoGz=}5��,-Q^�bH8{|{���Nἐ�������8�1
g[�:�C��8
�M(h�~��L���17�F究E�/���\/%��E����\t�AQT{�z��a�'u��mD�	tbD��Y+���@0v�P�O􈲎'R>_�o2H׋:�:KQ�#k���ϟ�~>�Ȣ�w�Ju\D����8$GY�Pc�Y���vZ��)Q�+��I<�8�N�ؖ:ݫS}FQ���Z��x�G���ؾ7��ʛ�������=]��f�L��?c:��;s�U���kHM�c%�Kz��k����j�E$����Mc�;����eef%�㋌�_�H����ƪ�˹SI�wɦ��d{����=�į:��N�����E�>�|��X�]�~�>�����8S��'ՆR�_[7b������Z�ص��[>N�b��_(���|7I�����!���E�jW7׃zo~����t�I7~��jYq�O�:d�]�iQ�M��{e�gZ��jE��6ڌL�v|/CP�m������QW>���t�<�ԯ��#�B_n�nFam����띞���;PEވ�I7Dޜ~��nT�57z��*,�9� �޾}+o߼�
`�a;Q�n"
И2�jo���o�M�~���f�u�Ua Pf:��/�;Yv�"�m7��)�9h�{�Z��A�� �|�y��N�j�� �J���jy�V��dצ1�����c��q��O��A52�B#��k4J|	M6`G�I)�Nj�Zr�DT*Ud
�0=�Tpa��+�bi_5�3xyQF��2n�D�$�J
��m�3 &j�u\a�'q@q��'�JX�����<���jm%�9]Z<���(�;����uI�L^��ǹ��t���X2ݣ�xd�js�� N����m(;��F[�j�B�E�)@PG��\��s	��x�[��r�
��<E��r�h�	!�5�e�ō7N�[Gr��ң�v���2)��3�?��GV�
�8z�����7;_�9RR��w�����+��P�Ѥ+i���/����<uct02�2A�]+���b��a��".��l����uZ[1(f�XV`Vo$�*�f� 3���SA�@?dv��o���s."Ȅ��II�u��]p�_6�8��1\d�Vs!2Z#��6P狴����k�놅+������	�pos�ut::���>E4�O��c8�k��De�y�/�)R�aHC_Bd�U3-�^��^U���g�NJ���)"gMF������k��0x�T��-a~yqQ��m/�z��0jHI� �nŀR� a�Pҹ�㩤ֽE�@��9DrawPع�������jH�J�N�n_)�NS�������7Hq$�|��/�ժ�
������T��q=A;[�������g&����s/X;��)�c7�^��M̫��	-�l^�dxٯmN� 
�����5�l�Y��ۿ���F����7r��Ry���R�U�`��~�Z�P{$lD��.�("��/##�U�yhŴ�NA�]y�5��\�C�)s��a��Tj�T����ܴe�Բ8O֎M��;۶�-M�q����_���Uǃl��I����N��H䞋{�AW�*;J�D���0of.�䙥1Q�\����%}��<��TB㞹�1���O���DWC�>�y<$I���%�q4�V�����q�Y�
$\ )YW��
� ����^놺���J\֙�@绿�U���R���ADϻ7o�}��Q����1d��4Bqc��h�^����^�w/}�a�,'	���� ��|x�Q��Aެ�&�@�l�-�����%M��SP����P('Ne���}"r�������ͩwR�,�Ƣ��a�<�[/�h�U���@����gX��bm��i�^�/+�3�	6MM���1����Yx�MO�j��=7N}��T��htՌ�<}���	�̮]�Ź�^������rm��ǵW�& ;�_��r���e���AS�:�x%�D����ȻY�m��D�R�z���|W��{?�!�����\G�Li:n�� s*߉�9h��c���h��&d�A�]S�Dc��W"'���� f�T�m偪� �`.$!��5�K��������3E,K[�li8����+�D˚��#����3dX�sg����v��{�K#uT�h�-V��w�� (������e*�\�ذ��O/�Ը�M �J�Ķ8eF*w��,J��L:�tJfeG4G3&��2�]ջ:2a��Ji]@����ܻ"�gPGP4� 3.��@d��̵�M-�k��`+��Ҧ����gW)T�}��d��W(T�Q;1~��c��%�Y����}`�_�RZ;�P�A�
ZD��s��aJ�s��$d��ֵ��c�Y�_zZ��X����ETμ��c�l����(1
Mi��g�r�D3��UuL*�4"�����zzJڥ�w�d��U�t�?3u;O��/�lM����(�G�UL%�b|Z^�I��:�F
0f)�Dޓ��ɍ�J�N�=�g3r���vc���)��ޝ։��:�v]Dob�d��b�(��g>3�	d�`/M�s,������GD�7%R;�����UR-e?sR'�EY��H@\wa#R�8����Uv��_�-�"R���[J+\�y��߻sR` ,�/��������h�u�0��e��<J���$S����J7㸁m�ET?�K���tM(�Ӹ�^�ݘn�����!����6x��Z�i��3�i���Ԯ;�`�k�Rq#�&��m�0�,�PG�4�Xh�n�u2w�#�"�b����"7�g&�K��]nS�o��.�|!E;��*�6}:��TY�_s���N�y}���Fy�w��}����4|�XB���F@����*7�j\��*��g����:��g��\��N�p��C��:�hH���-\1� �ZU�b�[�b_�j2死������
c
2(N�޾WP����U�aÅ�a� "N�ٛ�~R���������kC��ZSa26��7��1�7~ɔ��񺨬U�r��F�
��8sp-������ ��=�fx����\kD߀�	-d��*�!:	�����m0�XˈrX+��]EX�o�zHZ��H,h!�٢b:3Y]��C;�d��cj�އ�QU���
�����!ʟ;����^����Q�nǼ�3���ߨ�Kf���[,d�x�a2n�5\�ޭ��%�Fm[l��Dn����G� )pPǋ�"���Ӱ����q%�O= �s��4U��=_�&��ˍ\ɪ�� ��5ξ���u�)��}cV���R���^�Jr�PNi,���RiC���<�oQ�MV�9��ͩR\%G�kx)��y�ig+�R���,d�m�4`$Z�i�O1І�İ}P�_�8 ��=�b������+A��+�ᾋ�i��n��Ԋm�L"����=����PǢ��Q�8g�Q���!�d�Q��\<�js;��ܺ<8���{	S�X�u�ơ��Zj����s'�g����|l4ұg)�Q��T��9U��[d�΃II�@�E]dMA��u��	�e|_�Oߴ4���2/
?� [eI����1��8����>f^�� J_�����]��o6���~��kg�9��ZeS��ڏH��S-Ԙ�3�Y����d]�
pݑ
L�?9�,Z����(�UEU�5���9�Aߩ&`��k0m��M�>�gS�7�aaU��7%�X��C&������T�5yqc`N�QVeπ�������	�a|WR��о9A���;J �"Z�
J6�ފ�螈�F�U蘚��0@ǸxʻF�i�N\'���H9�����T�d�q�07���7H=�eS
 �N�E[���Z9n�,if������f�)�$�kJ�& ze�?u$E�O#^���i
�E��Z[�ۮ<B�Y6�7�B*C�FZ$o�� V��M4!XJ�{S�e�s�`Y�� ���>A{$�X)��V�������X���#�o���N1�����hw�3T�j��)+ß6ͼ��T���}��m�Snϥ�D<�ϢU71�oo�-ܳ	t�ר�������d��Ї��Y��W=(���ײ,H������{��ᢜH�W���	1G&�A����G���0#�9
�>����4]��� � �d�������\2���\cᵪ/L��M�ܢ�K-R6�])Y\�U��.2�rMz�c���%O^�&t��=1.|��)6Tz.�wJmMY�ܸ+9̱UΚ�"o4�[l�#����@̖���o� �Y�����
�z�O��ԸaT�t)( q����)�+=����Pr���K-K�0D�#�L	�R��)gzէ�$�� 	�yc��Z�e�hH�0����xzp,�ǧr���4i���g�iшvm�L�L�PT|�/1������<P2�^#\���&��d�o9R��!2���{3�zk��osl�!�R�9�He�9>8��#M��=��5�M�S��oר=��&� �Q*�"
��ߜ���=��]5i���;��PX��Cֈ�6	�)�6	����2!�sj�rs�^w��s5 �6�B�$M?�;;�T^�	�j�PR�"�9�gib,S��b��Dр�vԢ6WCUzUꌎ�(�����x�x19'̆�k�;��D�V�բ��џ���X�͍��a���*ټ�2��Ȓ�j��b\L���wA��u�ܧ�k<��WI���p�O�췩98#�4M�Gh�#�+ГJ�kC0a[��{����`�u�%�q��J �wS�lzNs�x�C��S��!�"ʄh,�X�k��s��v���Ύ�"9�߭]4���pB|OD��8���W�������5�[ ;�@�Dt׿E�HHptz�T�(�8�#[���j[��i-�$���WﭘrC�p��[W��M%T��TW��h� �d5�;�(��j�#*zRczd�H.�������V���5U"��w��$��4�U�r��
Ф�s����s�%���l`u�coL��R�V5��$�24�ƪ���ug�W�6֙��q��zmzm�7
8H���s��ʪ�Vtö��l���j����t�Zc�#����[s��/���b��='��d�r���:�x.q5�����5�{`�q�m?"§����}�K�N�I� VĨc^�
�����r�wb�Y�qV^�r ��(jjXy�L:Ҍ�h�(�譯qߛ(x�9A-�U����WT������<r}��&�3Gxl�>�Kp���G�6��)3]��:&�������C=M�e�܀H�<f.*F��Ĩ�c6lEW*'�P���R����ǴRR�����3��%B$K�C�t�k9��m2y��s�����a��n��5�}�徱���x���R��������z[�Q�� ��B�H�=�y��S���k0���R�.n��X��:�����i����R�4���A�0��'ڂ~��R�C�8������
.%�r���/�(�oEd�z���Cg�N�0/Qc�M �YQ}�p�r������h�/�q��徦�QބR^ɟ���"�Y��UC�{ܰ�n���>�wߺ"�'?r��pjY;:k勏������\$��ɣ�c�K��9�ށ�q��*ָɷ�JFN��ִу�F�:��nH�%~��~��9�9e͏��A]�ص,ů�F����%jd�(�4�f�|K5X���=s�U}/;�Z+E��H�U%�ʃ���0����ȸ���|6��o��f1��1��g���Iūi��g5I]y��ךp��H�#m�����^��6@cq����s��!k�*/H\W�؆���f�4�d�Y	����ӿ�Øؘ<;����q��J�� ���`~��lr��syZ�)ˬ�A����dœ��7�^AC��oY��zqse����ܛ����U���O��2���ؙ�q=�R'FrS���Q|ϩa"�eK��#��=�l}�A�A�`�9��.�P|��U�Q7�[���d���שz�[��C@�uCӃ�r�р٢�m���)eo)c^��_Cī& �������[��Q��gz���}g�$���@�v2�\��bz�3����t��^%Ձ$WQ�"� 7�l�z&t:���C� M �h��D���*�Q�����'=OT����+�L�'%�@�h��	��������{ED+{�2=x�S����YwyD�sVp�?�l�T�c�9�O����]�ß�^Su��M���;�������e=-��C$�������ͨ�~��JЛC1Q�и������O��ۅ�V�x�cvIc}\#��K�h<��W��Xk�����K�!"�\�Q�u�K<'T�E�ܣ�c�7��ӧ���0'��[;/_F��K��ɢ0Z��uB:+~�ǖȝ��%>�w������U=��_� ;)�ϾM�t�gx���a��
�����7iM�'�H7�m���N��+�_w�Y�`jוׇ��Ӛ2��B�#a厒����,����_���� �H�!�j2$H`�X*	�!�rT��Exe �4�[7 �m݃R¹�@gu� ��-�x ����m�	�W�bjy��G�G����ڶ�w 4����>J���ø7ڂ�ʠ�=��ņ��o��l<rS��R�3e����j�/�P��3F�o�D��!��������P�<y,�=V�
ii{
f-@R�����K=��Ge�0ʕbQ�V�|��i5�X\^I�q�co��gJ$����:Ӵ�mǦbkz�)� u��,ZM�::ܗvu3k�}4��ԥ(�m��P�X�2MzA�U���K�_F�L_&;�@h�ɦ�g�����K*�b���K��ৡ��d��T�����0��=.),�-9C(J��Z�S�{�����6���;�˶��]ᨔC��	�JOr.)Uue�D.*�RaUr5�4${OU2O �-K�����M݁��\�.�bQ����5���@�8����w/u�K����2�6ǫ���F4/��BI�A�g�zM=�DrE�O�=Ln5�D6�xK�
P�J���d������5��3e�9044�Aӥ��xư����NV�#���)�P���π�V�����y��^wUS6}���[6��|��LAT˚4�®[aTG��"h{����}?�_���������ECWd��<���պN���QWb5��H+��9�kU�N9�~�5�}D&K�x��[{$J�ҝ�+���[���*M�T�!W$����<�u���t#{�+�?�6�C���4��Y�Z5T���C�*]ޮ�z]�}}N��+~4�22Um`�:!����FE�>�c����u[�Jb�
׏��Rq�e�� �2�槎��堌�m���d^�"�z��M)99�4�b�tѾ$���u��TesTa�rF�kZ���<*�neo���"��c �99T��g|FJp�S8�i�轑)�vr�7DD���$J+�����h;8�(�/nW�����r���:�p���v*�a�q3���Ob �����iz�|R��y�T�&F����_��T)�-Ơ���z \�rN�:UDV�]}f������=��:��:�����LAf9�es��#C g	G�d0������l�4a�I�ᲙJ�T���l�&G���ZH{�"�Q�xre����2l"MCL�0�<���{VO����;��葜����D.)xu�;�V�,���c��]U���(,A@���k˫F���Z�'��c\H��n�Kл`J}g���߀
T�_�H`�G�C�0�R�$k*��s�Gʭ�
��38�!|zz� ��5�5G�G�n_�����X �{o��A�衕���J����Ct9J}ݰE���ue�8Ni����c��g���Sy���V�B��ba���w1�`�wB�L�Jo�ttc�˅o]����p�����|:�g���H�����Q+�3�󋮱��wb홋Z�F�ǲkƹ�����;ç���Ƹ�+��͍W\���6�\�Tv�@��yA�o�C���[Ԗ9�J�o��S��,'����e���<s��sC�IS�,y�ϳ{�=��(�����g*m1]ݫ6�(��\�P��&X\.ME�R�I�+a�Xۜ�&�6Sy��'���A��T
�9��b�m��ت�����c��\#ݓ�������FSm:���ǀЃej��f�[E6�5"ahF%�-U�t�4��bR� v�d�>���D�{����� �àR��#N~SQ���8��V��uϑ���}�/��*��5���d���B��(\p(���.#�ϋTx[j`���Pw�!�U����T��L���2m�������!!�㖦��?K/6����?EX@�%�-=��^91���l�E�z���ą��d^�t=+
	��j�*y/�5��yT��~���4�Ć�W��b=�x)��(��X�n�:�C���w՚��,���#�52ߵ��s4u��M���Yv�F�"Jp۲S��&��6^�,��H`�c��{O��U�>�q������W�(x�,�`���w6mC���� Խān�O��4��k��t*�Uid�����c (�G��P:���[���w�<��ʱ��P�猣�q�k�K\G���� h�0���:O�r���{>[#�^{DT?y�Z��l��د�.�)�� �Rۅ����b�:j�v^ͫQٷv���S9>��jD�?9bip�w�ݘ�F���s�N�`����d��G�s���|m�.fEh��s�{c-���p�v��͓p��Q�~��S����?�ӱ��%��±�Bu����c�u�I�_�������Tw1��3'�m&�i�Ty������_0�����sa�o��2/�H-D��Z���Ry�C�J�К��'%�81�՗X1 Q8��x�ꕼ|��F���pB<crwR`'_Sa�W +�8�X�&#�����x�V�T4�JZ�Dl� [�ٹ.|a�^�9�(Y~vz:� �/ 1�{\Z	A��������P����Ty���%�E�hDO騥����i	��^U�7�GR�(O=��H��*���߼}y� �n���T׌uΡ�r���������ݻw����^�>}"o^������Vv�=-kϧ&G�6��� G�ϧ���^�Ѽz�������J���lv6�P�-�I4�#5�ޜ����)q��Jq�{�����ͳs�������_Y$�(W�^��\<mlj	�mj����j̠!VB�ū��4�X�Jt]���Íg��%:��>C1�Y��E���BTn����	���'��]��-#���O7���h���k9���҂���zƈ=y(t��ѕҢ����h�Yg|��}�b<*�Fx�sS�Değ9װ)%�ܵ�g��� ������V����7Ɨ4D*o6�a��H	$���$҈�Jc7+����������N.�j��#ϕ~�Ig��aX���/d�h_�O\W��N��� ��g�$���z~}��Թ�R��y6n��d��}��
�W	e)����m嵧� �" \��rC�S�\��i�c�1g0��j_I�IB������C�9�?}��d[��szɸך���F�"�����"~����H��su���g�^��T���#��*�q%��I�)��h�ZF�$� �>�&Pz��՝�IGh�Fs����sǐ0~����S]s:�V@��P�������K��3Л�>.����=ǝs��P9onU�sI	��Н��`��,d�Q�(|mͮ�3RV�<w�V8C��Q�C���3�e����F��ӡ��>p4�}-:��a�������8 ���#�oF���h�u���׏c��'��v �@f!�Ye�X���rgp=��}Ur��L%"�H��*[3�B�PȨ��Wҹ�j|����.<e�������C+a�}=�y(��GY�}0�S�)Qu�"�Q�v/ӗ��Zc�g��޶o�٦�����M�y��]�����ȹ�6������-��Sb|�����˗��ic���`�8a�>�m��M����7�J��g���w�~W�_�A[��ڦ�1����QX��*\6��e���(z�͕-#9�t[ �TE���u� v&
[]v���AY�y�7Q�_��"��Ӭ
��+���O��5�i[<Z1H���&����hFu^�������
�BޥT�.��&�9xC���,?5}�D�P�[�$��h4���{t�<8�M���O�/��/��a8�n�+[T�H-��H�V�ICK?9J_6�.��|S	��A��pLs�S��_�c��$��G>�f�����Z7څ���X�@F�U�a�����c�5���2؈QU���P݁^���) �����{zm��+6�ƿ,��:��5n&I,J;�q�99=Q`�ʴ������ՋWc߯5z	�<�߽�y�|8w7V9Oж�=���&��Ovxp������0n�^�
堞���Cm�B�\��MKU����Xl v\� �9>��5*�㹷��7��H���>�AU
�s��K�b'-� DeG�Z��-"���77$��1�$L/�>��%!'1#$[�ԛ��r	C�ۖ�����@U�9���ڦ�GP+�;O�M;����B�\<�i��R�"5Wf#�E$��8���0�'���g��|=�g�ʵ��¯+�B��jm����I��걊������Q��"@�;�(K
(�G6��Dܪ��XO�% z��X�}�eo�� C�����X9�'�[`�ﱍ��/*q�������U@9;� z�Ư |�������,�o�p}�cr�~߫��q��[p4ܮ�\쏿�hT �y,-M���9�$?/Uk�c<\k���l��d|�{�Ҫ	�`�VE�e��C�l�����)K6�XJĂ�7���ށq���QnF=�V$'XF%hB���q�N�ꅋ<rj`c̻Ų�=l-:�R�$�1Mn��/E���P9�,��^�w �l��Ǿw����4����GS"��C?L�~] �@����q��Qך}f�C�������/_x!�CE�������țҴ����`��z��;�[���F�)�!��hfA�w�@5�U����E��������= v��x./^��o^}����ߏ��Հ,TK��������#y����A>|��A���ӽW�*[+g�� �a'� �{��_�L�����}��;	=��i�2GcN�9�"O���2W'n��3�m���ʲ+��
]gB��' �?
� �| �:׹;�x�B��7���tΌ�|կ��ʸ�=�@P�+I��DT�����ڱ�0~�~�@�����%�y ��;t���y���'�^��o�p�����|���ъ�Z5�� �nn#C@Ӱ��/R��?��~��Bm+��*� g*m����)�HWW��Q=�W8��*WI*up	u���U8t�荿°�(w�]B*`g0A*�&�Bu�Ơ�@e$W?��v�/q��W뾯�:�9��}��[O���&�3�gߐI��E�,<l,%\s�,6+��d��=5����R�)���i}��5,����ʶ�°Z����";���v�^��s�E�g �+eA�J�O*�����Ƌ  ��IDATP�,�2�q-?|��o���n(Z��ӕ\}������kE�����^��$�yЕB�!�"�	�e�5�n��z�e�FH���"�

�����Fl��;s�#DaIk(��*3������:I\k~Z�Уr�3>��k\$]��dF�QM� ���wZ���p-�*�	粂C�y	��wz�1�������/����?�Iۏ������z� �����VA�䀚�s����Ѹ!aĳ��:�q�g\�h$6�}��6@-�L���@�F��0�m�{J$��X���#�dbNEO���][�P~��7�Y�D�A�~\�͸�e9�����؏g��JۗF�
���q���No�����H���փ���V�N��z��%���g�Ā ��Ri,�|�y��#�����"��&��T����Topϋ[ZY����h��NӈDO4IV-�D�8�|�ȱ��՞?S�j����=�մ��l� ��%��/@Ym	p����q��shp�1���1V%��v�B4��;���`V6n��e����)�)�SaP@4�����C���#'�U��~/�f�
h�
:�m5c&��)C/��݃U�{jiJL=�\ɗ �-)�TC���=�-�L���8�_.Ch��aww�83�z3�}��82��u��{v�#��-��˯!�y����r�-Ć��x��0,��g�K����aˀT�+�x˴��&����XZjGlRoX�{�VJnS���T�#�(�E�l�����s��U�ϸ[G�_�L�4f]΄���2�1������#�#�o<��]�Fܿl��T�Zy�]��,Ĵ����e)l���7�9���F���c�(]���1����X���Doib(bq�:�r���uo�8�Sn���߃�p�:ؓgO4���ﾓ�����ahʚ���6�؇���0�"�����L��z!���������^����	��O� �;h���39�~��﷢�Σm T���	=�r���s.4�^�[#M��)+C�ubZ��/�ʾL9F�QC�DRe/L�y�<���F�ݔ���!#�p��QQ w�v�z��q�0�}�(r��xO��,���=���'(Ǧ���Z����z\s�J͖������y�Z{�q��6~?���_���)G��=���D� ��s6O��m���j�ұ.���y�9=��ӧ
�]�^˛�o��Ǐz�w�����8��jt]�W�\
�-G��7;>�W}ёʏ$,�����>�6Aٗ}'㠣�g��/j�l�q��^pg����.uMN�n�`G�g(������j@���z��)�7bGf��-����y�]_���ɳ��G}���t���aQ�-����޸1�����<>$�0ra�w㢻��f\����L�E�v�i���� ��
o]��-(��=v��o�m9H٬L���6�����U��Z�SB1�?T"���b�H��!�Ӷ��C��p��>7��R����⓼�F79��4D~56���B[-���r�]!H%}�i��Me<+�;;�?�O]�Qqvv��xT�M@(���3t��8�z!h� �=m��q<9Ξ֐P���Y��%h���R�zl�bs@�<غa�o�4�0�ja{�j}#�����1��(9Rа�|������������O�Rrs}#�߾�?���fc�J�ҫ�i5��+�.,���c��<QϘ�(�J6c�)]��� ��ց)_	a�Zy�See��J�髷�q�x�i��
���bTiK ��Z/���o����K��~g@�)5w"�y�P�L�5r4v�������ɣrl�ٕ��ZQ�� RgX[�J*�3b�����'Bp'qp����Kb*�4�����C�*-&Y*V�4^!Ng����eǛ<�������*��sO��<߯=�OO�x J�@O�?�(�6������^;�ຜ�X�R@��UidPPT�Ƶ�>�G@��7�����T?��k�254c���m��J��Z"�+�^��Z����
_�)��B_�~�&��=1RZ�	鋀�����3Y���) ۧ�:V�U����!�:@9Ѻ��͎�lyʓR� �����1���Ib�g���6�C����ԅ�d|$�;Z�c5��ӱ�|i	P��ΈA���=�A��+Y!E�=*��9;��X�bݗ��*(;�B�s��s���H�٠Mƞ㐶�X�l��u\��ؑ�`��dejh�xbI��e�0}�~� XL[_*�k�uֹ�reGJ�c�gv/��լR���T#���/�tf��0�-%��{z��y�+�M��� ����R���-Mw��%xi�sj�i+Л͵�TD���z�����}��F=����%h�\�\��3t���39u=u�AWu�����ئ��BR��Q������pS=����H�����T#u���?ȋQ�B����}/����o��y����{�L'��,�������8�r<�m26�~��G���~�[�,�M-�}k �A�^�28�jXL��}�j����aӹLn^n��A:��x�:K/B�So��Jx��֢��yi:R3v�Ei�ݰԩٚ�
�"�XUٮ�3����:+��x����Q�\4����W�8�k͢m:��>w���YwFuж�����}��|Ex>7W:7��~����z��X<W��Q����XJh>�}���������&�����G�4�`��c�6�Lq�QS��q�u�^�F�/u��v_��q��_�ӏ"�VT 7��J��2q����{[F�<�j	���cJ�-�\�R`*c��:�s�����AH@W�oB�Q2�=�[��<}�TN�Ŋ	�׾6��Q�c���iJ�d��\`�)C(��gy�Q�7����`|i�z;ͱ�b��W���5K����8r+nF�瓹ԍ3ї�Q�������'��wEK~�b��.ح���;�عx�A>"=��U\��-!�VȫkI����oC�f�(�^����n׉�ĠD e�I"d��O�����~�{�Z���&eA�L&+��3t# S��y��O�v���
u��b����qX��:�v��M�6	��2�

���b񹥇5��2��7l�:�c��F-���dDyʭ���/��po��K�*h$67�Ř H���A�1&�Σ���S��'��x���?�fh�XՁ��sD/�$��\ќ����񔃼V��.�h��v��m�QL�G���e��o?�=�@�����O�5����"%��?��Xז��Zӕ�4�l�P�T=1	�Cf��������Yʺ*Bo>oʚֵ���# �(NaR^�
T�}��[@�����.�j�B��m�%ZM{5�<w)���Az�Im[�����5�u\_*�V������p�ĥ1DM^�� �7�ݣ"˖Ͽ���To�Ns�)͢��T!�Vfz��B��ڴ�uI�! D3�����Oe��h�ة+3�2�� $��z�\�a��#����?��$��o{��ϼ�i穓G1��k[.��S%��k&�Hl�Ě�kƐ������#�H�j[��B���A��;�/�����/뚎'n �.v�^��� ���8̀H�F_&�=�k�3��)F&R�+������+�.���N�|��΢���R�Q��~�w�O-�qwk���&|�p4�������s2��'�Jppp��9��F����֪R,{�S�4Mni�:G����?����|��w�����f���������G������VZ %/_���ϞZUׅ��w�f������NNvN�6����-	��BBc]�Q�������Bݕ��!��H����@�"^é �kI%
=��	׃h ���5�)U�,�
SS�7+>�"�NFM�u��E��ܕ
�-���f����	�NÜS�(�T��,u��k��f�:���p�z3"��>h��,��8R����=(҂h=8�WN�ix���� �J�U����w�$5���o�.Б��pL���P���q��o �:��ٙ����K���/?&;_��~����`�@��Uv�a��)�A6r8� ���@X��{r�XC�4��Ή�F�qus�װɣ�x�;�(�����ٷ����ft�hIkj�F�@�׏yOh@q��P��%E�88ߌ��rِ�.�7|����R�˔�Z�ئ7��g
�*h*��'��p!�>��Ꭵtâc����(�[�������Ub�*�gK����6 q�6}P ȅ5ƈ%[A6#��P8��Tb(�(UA�Ӕ,�����(J�]7���kn��o݈=�.R�&1�id�����4bf���ʁ�@�|��^��m��
�\E4�G8������z��y����OgJ�ro��t|^����1Ŏ�{�-�Y��  �D��X����{����{s���ژ���BL�(G޿ ���c�m����B�܍!��. �㵟;ك�}u�3�'�q[ ��sQ�|V���61&x9wUN�P�7L�������?=�����KܐӅ6�) �������XX�������__&�6N��-��BI���V��v�j�4��ޜ�Ǵ��HzQ׆�<-����(�����w�y6������z����J�$M9l=]Υ0eo|�	x��-���v�m��x��zn��#���;2�4�g~�ς��=!�WR-��qD��!{��U/�1�+[�b��f��P��z���S�ߍ�#P`�f˹ۺ[�ŝc�k�*�1����E'��k*`'^������xH�lM�C�)>�K�	���L�/�W�S����}r��)��vw�i�Z�d$��� �-{���\.�?�bImEBǔ�sͨ����,��|.��0:��A.���k����5��֘���(���t�����h�4�������A�v��R�$@�"��q�˅�g�8~��O4b�(����x���Nލm�
�t�����b4x�ݗ/���"o��B+���絺[I��2��&���q]��lɣC�9:ȃ�'���J2��s�J��Wm}�|�lLG�걝=CMrY��8HF��"�G=O�ϫk. �ZY�/s^[��zu��ׂQa>�'&�T�팻	vҋ�͢��5���u�Ո��*�Z�N��Z*- dV�V��jl��8_/�h88[���i�`�i�7��ٹ\���V�ʋ����g�[��]}�i�ϰZ�ڷG�筴]�M���aO.[������<�����/4�݃4��?���upS�D��P�@���Y�o��eyB�˵7���  @h$Kk���T 	\��Uzn�"��揮Ef�����s��L��A&�3�Gx��Wq�MJإ1��b�����sӍl�b��VRXkIo�(������I޼y#�?��Kx\ƱʕrOS�*���wYZ}��*�<��BZӰ�7bG[LN*DIO���{g���~1[�)R�"R\(T
\�E	'E�ZcBEC��)2�7�X��{�b��t&b:'�.���T�(���V^1M�I*��r}�I../4�}���5������ݨ(������˼kk�r/;�ԡU���b��e��cSԪwα�
"��D)�K'�.e>u�R>���pb�!�	�TPB].9s"�ZBT�v�W�@�놰?G�i��8f{c��Ư�!��c�N�R��H�"0r̓#2!-Ne��{����Y�t?��W-aC\�]�M�E���������yC&m�eCie|}v�ٔQ�LO�����o�9ʻ�25?�� u�@��O���KDc�S�4(��_;Im���ݔ�AI���z�w��ƍ�"��H�c��񚽓�G8U����C��>/��VS�*�_ٖ9�R޺N4�_Cs2Ih�om�l�J}�l�=�%u���������U�R��f{�:RSTN!�z���8w��x�����K��44�ӗ�-�sW�T��s�õ�K�gȽJn�:9OL���?�泽����!��x���߱h���D�8qr�'��T��bp�T�<�FG^8����y9����)�Qz��$l��c<��G�^r*�W�Q��.�Ğɔ���R��:�DbDW�~R���&�u�*�˾������[u�6�(-�2�R�L�e�P^��L��\�-�P ~P�IE�)W���mV���O��R��b�G)�m9�垎'��&�L<��nb�Or�*vJ��i����9�8)|������Z���)Z�ѫCU�URCE��3�h�tX��/��0���q�N#A�J��s�#P/H�F�i�3��{��]hɥ�T��?:�T�x~ƽ��W�.�����,����9iq�� �<!υ.�˱qu�"��l��T+����h#M�R��+�4���h-~�t�ȹļ����c9?;W 	�P�|󍜌��F0w0�>]_�8�eq�yaq �������K f����U��o��;O
�<��F�g����'�u%g�7��G7��\m�;~���� lu��X��"�^������4O�)z%��=�ƿ��3�< E�6eBK}����Vpg=
������%##T�A
Q�1�E�	��|�����Ҁ�t *�f�1�M��1��r�Vr����}��� ;�Mh�hA��1���<�_ys�[;Ed���@����͌��B���v�!�ܨ,�-�8��]VE`�Ts�X(�����|����]so�I����o�S�)E`�M4�&�7X�(��#_�x�.�@�<���o��u���
��C���.F�[��^����T�q��k
s����&GiQd]I�b?q(����e�u,J���;�T�M�J	�\����w	q��m2��L����~�h�x��,��JF��бH�
T�̯I������v�m����N�"���Y�H����ᑫ�d�Rp}�=��m4���DJ��TN������H����|wQ�����O,D�S���m��z�g���Fy�p���Hy�*�ո��
D0�Mb�\N4�k���;)*(�l�}�Pd#�~\��c��J5g�G �P�D�3M�S)9���-ь[���D����|f���r���+S�ř�س�D�V����{Վ[��¿\���3����1x��R�u�����cm�# Q� �������n�rkS�"�h,G�R���v��c�ܪ�K/U�j�1i�5&c�K��)O>�4���7�_I�Y�.V:V}��<�?!U�����ik�<�!��a��!�:B��\Q�EC�rx
g���G�ز�5V�ש�?O�n"��X��%4�c1G	c�C��^��K�"]G���T��F��S ����1Ѕ@}�u�^�`Ӹ^���lܭJj�=w���[�i@D�+�6��R��q���}�{�Q}	����]���J�q<�Q��H���CD���H��,`�v�IKEj�S��Vv����[�W�6ǒ�/C�!�.!yg���TK�Ɂ�_ ;��A�P.}����P���w_?y"/^����cY"kʏ�N��è�^z�Z������ɣG��n����jh7�S׫w�G6��$R��/9��E�h�:��@���<����ѡِ��e&���9N�����)P�����ߊ܁[ȝ����3�1;ַ��������?��mp�g�1u��l��~��؛�N��o}t�<�f�e�W9*����|H~Ӈ
&'�2�`�NhD�Y��#���Q������cEү>]ˇ�����R.6��P><0�'Q@&�����z���y�� �W*�"Հ���F����\��G�N�������L��6Z#9Uc;pA�#29ꀔ�~���S���6@�~����e���ym?LȚ5���ܸ@U8
7�Me���s�T��=������~[�ic��JB	5��!R��c���ƞ�?��Bw���Q) V"1��)*�+�x���/.���8ό�5k$��,ݸk0_��N���/N0��hγGl%�FB:���}&HD�:���ɔD��ZyM�s�m<�RrD�ȍ���n4�2�������}]���q�?��O٪0�5�G��]U���-����5NVJ��_�;�P ��y���bA
�����/F� /^�W�4��b{Ō?��gd醝�5��h�E��O1�Jh}�����;@*.kӶ�Wآp��/�/����*Äk3�f|�R�"J�'5N�J��8Q���V�4|�S�"�PR"�(��)ś^������2�Mɓ�@�ү��0���grч��xz�LP(����P�&�4U>b����+��o����Ӗ)|����������ַ	�er�Y?M�A��B�<.`;��9�.~22�O������+M+�EaN��r�݁s�8v�|J�W)�� �wf�/sc&���k�����o:u����l�m5�
��M�����p�3>��&A&��\_�L��Q�M�-��@M��[�F���'T���0�fԏn��FO�f�Q�\���^�9$�6P ��juF�B,}|�)�p !�Q�j�+w�qa���ꙹp�4N�O��z���84��tS/�Eר;�p �]��iB��k��}?�k��� ��鸚�$�l%�=��� @�� ���ܰ7 ���У����p0��9�q"rv���IL�c$G�n�K��������7����`Ng'O��)�E�ʻ$�竽�8��-�x�����y�䙼x�B�=&G��Zv������y��������������3y���O�����	*��9ڬՓ�=��֫�,�V��i�B�Ѭc�/_k�����#��AZ�YQ-���H�ӟ�����.%?8�O�.����\|��
X���*��uT�7M�^����f��~N����I����D�Ѡ<T�g�*��!���@}��RvjV�)�����yϽ6���4G ;�@%�1���º��Sw1.��ryzi�nn4��1x��nF�P6�v���^�]��mH���h���ً�w��N��m��;Uڐ��:A��� �3�[�ꮇu���f0���h�)I�0���7@���z՚�lڼh��[���r�Z��Ql*�م��.K ��(
�7�
�y�������TmOUW�h�z/%y[_���Yq����1BYü/�r�!���IA���l��/�w�x[F��x�b��S��V��������w�X���"�˸����%Gw�pۆ%���^9`	o6Bx���j	T �P�Ka�s�JY�~��g���9[jb�̚yÙ���e�W,c(��ḿ�z"�񦝶��kc������ӏ��ͨ��ƅ����Q�/��&1pG����}���_j*�u:�%�|]6���̄Į���Z���qM8�g���ck߷�Cû 8�[�[��E�_�U �d��G��U����U��H�w1rv���kn���GqN�;�=oS}n������*`O��;plĒFci�u}���QE�A��B�6p���<�D�Ld�8*cV�%. M^����ָ�л⫷�"n�[�$�~�q��tYɹ~+nD�<�R���r� �fk���B�҇�ss��Y���$>�<y2�%�s��V��	��� �oֹw)X�x�7�Jf�SVx\{�N;�vtr�'�\��^+��f_O[�7�������0P�J���UO��?����[8	��[f$�c#uŻјx�J^+��T��X}ҕ,UĎ�;�b��D6�Z�>���-u�5��<ٗ�ő0�]#]���鄓s O�/�I=���c�W��dF�>&�ˌ��VSj<�f|o�4��\i��*"��VW$*�����x��n���S5=�5v�N�s7'd����8qVie�0�̘�f4����+�����xq!'�DuR EH{��QP(��
��g�x�e�$J0�\F�x9�iN��[)Ӻ���V��X���Ȝ��D�Vya�'龕�>%Y�����L�	�X.ݞ9����x�R�����k�?�(���}�#�5���Q��Fg"����H�Q�X����s��H/pk&K��s\Eiz�O0�p6U��|qÑPP����� Α9GZI�W(P������\T����~�#*k��i4x.���"Yu�6�lA���(����a�\N��\��g_��c�(�Apf����K��6��Z6��;M���4g�χn�����������K�ٯ�b=|M����w�]�+I�@0��|8��(��j8g��0�T9)ע%���Ȓ�𶫁���`]ߗ��39{tf��H�r�K�:G�L[��6��g�`;>9�45���AU Dŀ��Zh���J���*�p�C�	����^���
GSV��t��O>q�]11�� }B��[���"n������Q�d�Ad�kVm���!�m�LY(l�s�9���u�y12�E#�i�����T�%۳va�fy�F�d�E����y����x�.|GP�X�|�,�K�\����Bզ�jf=œ��8)f��ZN
P�x�C_t�n�m��Y�s#��H'��u��W�6lN8k�?��AX�¼l$����q�Y��.cϱ�w޲ƫYy���I�P����;Ջ����4�WH��3� ʘ�z���<��騄���'�!��� ��K{٨b��[j\{�������:W�	��k(�21�^�t�kq�җ\S_I��{�%��a;*0�^��BZ�Py�h6���zps�o�!����}زo4n����>w(�T	�=��t�
&k��
\)%S	��ҡ\�'�<�pjQ|*Ɖ�_�Xڛ�ʥ�k�ؚr3�4���[��_���YT�/iH^=��&�[�<�N����N̸��UTS�WD�"�z���Զ�yyh~�znGd���t�>�{�� ����ʇ��g�~ԍ�S�0�]>	�{�3m
$V7����
pbE1g�h��7���}��>��F�r4O��UQ~T�Ξ����������U�4�?~?��y�,��i˨�@����]B�K!��f��\���I��Ӕ��C���x��(ZK�e������M���G�58�0�H�M�z�"��B��&����B�g�3�/���%qӨ�V�E��Ր���
��q��:�>t�	�����ڹo�8��D�6�W��>����Sv�� vg���� kֽ0(�Ջ���EW�m���kL<s�ݳ�xp��O���D=~,ϟ���U�G��H��u�U�:"�{�	��Rgr��tQ�,"����<�BǏ��F��UPc������8i�ʹ�h�D��~����)�����/:RC�4s�i���-����U��K�,��
]�D��+�m�A�xl��EoQJW������u��Ӭ����]�w�8tKj��#�:��9;?��5��GP:��gU�0w��3�s����-�:��������('�s�1� "�n�o"2��5m��*�=dq2�������h�������A��ף��K�[��E��
'����b���:5�m��s�g�t0��s=���z���:���MY0�fv�\}�����3dx�-+�h�[OM�5��7m;�u���*rkS���hl��;��}���%az�<�'G�Ko�q�]���}GS��;��!�G�ʑ�A���JeHtk�y^N�ldG�� �m�i"V1�4,��|������e���)h��� ���{�N77T����}lJ�^~#G��_��r��~����^�1��
R\ 7_�} ����q��x;��VQ"�?%��N]��O7;&��Bh➭W��Rݕ�dnx :a0�gP4����Q�'J��I2��OܘOh�B��ݬM�s/��՗H������y����!Q~�F�Q_���y%J��)�])��k�~Vh�&t@������k��Zy���1��6A�֦�c�C'��Ҷ�nN���>~���@_��̀�PP�������1Ͱ)�Mq�<ŋ���!�yT�d�q����� vj����W����.
9�k���K��1Fs+G�z>�_��a�C��k�H;�҇�5�=��x�6)0 ��]>��q[D9�#֮��f4kĈ���UT���)�K�_�_��ގsN�|�����T�ivl>�-V{��<U��iQy�o�JAMR�����ĵ�����#+��I,\5�"�*"~�����;�;=�Bb�G���WnJۓ+�Q?Y[��$S�?g�_B	.��H�)�!A���n�����]����4�d=Y�vm���|�3�t����9���%��*�T릾�?ּ���GmXo��5�m
�lo�N�|�\��Җ�ֈ��J2�q1ί}5��B�^��\vG��3�]����l{��L޸��%�N�>[3�;�m�����ñ��RZ|�L���\/�V"* ����i�Y-Kw��A�Y�7�Y3�,J$�Qdm�E08���XQ�K���NB��2�՞�e 6Y,�ͤQ��zU��{�p�w(��c�ֹx{9��w���%���]��3UzO�.��xR �R��:��$��8�jupp��T�\�`��p:�L�wpJ���:��g��C�����7�*��SvG�&eP��j�
pB~8��x��F� �䅦��'�EP{�o{xZ���,J�/=����@����՛���Rǿs瘎���[��&tƐ-�C�[f�j���@~�@b!���"��ۃ�; �N����1����� V�1�"��F�+���:��_���q�%��Қ��Y�Vc@{1�΄1P�*�  ~��>d�}�V޽~�c����rpv�� ̂ܐ��2��4Gk�:]5.����x. b�<�����{��9�ߗӓSt���k���켨!'*�=�����O?�|��z�������ԲJ]m8Vu����
��&@�}.ɴH�F�}bcϖ�>�ڸ&��~���Ф�d��-�ޟ���-��Mͳ���;)N�
͡��&��4~�����$n ��R�@o)��	ֶ%qXR>���:�J�����]��@����I?7��O���/�ū��R{� �f���M|����v`��t~.�����p�pGa��R�۵�lb�GD��G��r��H���?h[�?{6
�3������>��E#I�al4(�ث�Wd�#�@�C��Z�Bc�պ�5�܈(�6�R���C���I\��,�D%Wz��X4���kj$�=4���h� _cdO�V$�b@� ��^���!��pP��r3�{r�t����	�p2�;�(q���L�2���*��J\�v�7�G�fڵ�`�B}I{��E�D9#7�z����M7J�c�v����Y��,Mj���Gͻ1�|�˱Go�1q�wwD&$%Ex��_&ߐ[�>��5�U�6x�}FT�6i�^C;
`��\)Z"v")��}���g�i�u`�V֨��%Y�})'��Wy��5����.3un �ם��v�c�pg�������Ú�5�H:S�U�6�[��Vs.����$'�$ 1ov�9y���"�Z�%ٽ��p�s�ij�d�Y��1���ٹ��:����ϸ��(�� �8û��V�.$�(�����J9�4�@l5(���R��M`���w�s�%vj�\�@q�k��69/�� �Ko�7�*�c@`�����r��nv��v�Ք
OA�=�j_z̯Q���;�����{Je5�~�Ȕ�V �C�-2�ƬV8��1��Dga҂���eB�5d7+��P)::�M�#�����Sr��Np G{'^�i_�D��$��"j�> 7#Md��<���C����]�����	Pi9�ÏN���FK���ƹu��\z 0rgctx|"���������7��ul{��45�=
>�����S�"¤7�]�$/��R@���c���+�Ta��Q���{{���{T���c;�V���[��p}N��W��=���:�5�z�\-�� b�G $A��V	�)��y%�.�Ls�ͨ!V��l�1�<y�2���f��w��#/�pp�Y�]������~�k���[!�Dyh.>�/��X��w��ǣ]�t'�>�+������5z��Z�GO�m+%3I�Up:�E�9>_�A�Jm/�y%������;p`v^���s2�Z5��{�:������0EЗ��\m5��C�\����~�{�@�Nb���X�t<G�������#�,l~R�o��l�ZD(ŋG�9����ǽcT�^��K��/U�����7���1k�߲��}s�ͅ�p�W��S�X��F�����*Ӑt]�#�����z�J�y�w*=}��2�8��x�=�QQj�� �# �@�����ȧ�RҨ�_|Rp��gϞ�g$� ��/���>?>�pAD�`\ޘ��>�QHh'�g���s.泃4$�S0(%O�q�����K���0SD���o�x�J��nDM�e�f
ȡB���L$�ŘJ�H�TUbVx�O
$<H��h�a�8)��d@O4��&f.|�Uɲ�,�$�6T�axq��A�}I��KT��s�4Nz������0��A�\f�!�KD��z8px)�u�餲��ok��^��}����镆M�i�&2o8�HUJ��+4�}\ޛ��le$f�)�]�6��i���nj���#�rIA�V��!�����%k�s�5�Z��^Z28o��:f3oO'e�9^�3� i�г�ikY_l��fp\l9��'f�a��w#��px�K�j�ot#��;�W
�J���ǌ�ƌ�r�D�_Ѩ�H�i�;"��PZV�I�K𷊚c��#�F[]�����nG_j����\>�
L�% lo��'��D��4]��t��2.U_�f���$�MA���h\�і������V���9��>��@���n������9 ��gP�>�e$���[�Gn{G>�Oe�7�����i v\x�9i�M�<8�A�Ȇ�7>G����ԧ�u���D�����D�D�+�;�'s�=��$���<Y���Jt��F~8W��,����`,u�6&���V&u��2��� �uq ��!��|�yo��~+���S�'�G�������ޫ"q�s�Y*�[0���|!/^��ӳ�p��=�u������u^L��u��t������) ��gV��9"jL���=�=�|�ż�b���9��9#'i߱za��'���Z#�V�\����"xw8f"yr/������0��S�?U�O��Q�CJ!�R*r[��`Nb>R��J��B!P�TΚC�'9M߿}+�����z��y���/����c@T|zx"�K�d���6���Yɛ$� @�<U�nc M㜩����Er`g���{��Zc�����3�@�qyq�QY������G�p��ү ^�����Ow�N�E|��3�:"�K�F8y+YA�,ۆ/_!Ip�\���c�1���j���(2�ס�r)�GwxR��q��Y6��p�T_��>���@���u��9��&�a�Ռz�T7bL�bƳG`4Սj��7ۜ���F�58�h~woo_?z"�������?��������/��U3����y���,ֹ��_X��/>��͝\����f9*X��^]˧�O�X�A&w��x���3�FA�`��>������y��_��*W)4�}WD���zR�L)� ������9KW�.L8.x-َ�@O��α��w���1K�W�S�O��h�?_8?�6=/����00�?6���v�id��u����Oݰ\��<�	`�N�a��+�EV�6�0�����[O�G��\���G��`�yoV�y 9"@>��P`�����@���Dr��� �'bl�{�p0BGS o�ܵV�K#ͲϞdi 8O� � ���C)�l����T���[dq��	#f,R �%_]S�g��S�<h4�S3iز�yYz��*g+k�7n�KD� +i�<��4�5��t���"	�)�"\鹖.n�~</'�K�w.�؀�:;uV�D���X�i#���ڗ�	*��0������������<m�5O����T����Ġ@����f�<U�}?xjG9~��#�~���j �l�����؏��Ajh���=�q��F<֟���4��&/�s2�K�/(�Z���=�a )7��P�.#g-��H1�5ݨ!�/�~b�=�#���0ҵI�8��=צ�;)��S�*F����k�f��铥��h(���ǎ9�'}���.�{�I���Ֆ��.�1khF5.�{nU�~�,���3'�Q'm�Nm��09�����P #¶�17����)Y����$��q�J�F����*�+�]�<�8:C]�M-����*A_��S͘^�]W���H�M[�=0*Շ�b�MegQ#Q�˅��0�l��H������
��������M�AԆV_u_��rKzTx�|(�''�����1��GAŭV!��a�V�T�N'�0b�~�8z����o�J ?F<���5t��A �:V��V����h���_�
�:p�a���ng��\YZӥ�8�2x4�2�+o�lMV~��g��8�X sZ�R;��9���c���@�J�_���j�G�G���� �R�:�Gt����<�1���d|< ;�&KD�0�c��`���'�8;�L6�sF�x��̈́�[OKk��&٦�>aژ�����+��"�?"E�h�?���+�:'�E��W:���=�8���SM��[Y���g8(��/�r5Λne\B�r%���%RG�&w8�z�L� O���\ ��w���25��{o0���*�0���O��t�7WϜJmڨ`J� ݣ5�g_��o�B����}�~�_�Pw��~�xF���A	/[���wk��9�"�96�T���e�.a��5�j޾�e����T^�|%�^���_��q#��ǟ��o���?���@��2C�BP����T��k�s�h��(��Q���13ôR��ݽ���"�9ܳH���,c�����=	|�L�D�d�������1�߇�lK�THr���[�3�^19ԩ��Q���d�D�dơ<����������f�jh�����=Ӡm�b@pq�9���p2p���7^� J��G�{��q$Y�������hrfz���w�����ݙ�&	
�(]��׏)�PY�3�&+E��f�͎��6+�yU1s8�ը����'�j[]����3�()KM�im7Seߖ����fB����3	�p���T���Q⹄��
찂�@+�b�j�]��vߖ���2�l�q+n�=Ρ,� �!�œ2���r)�k�wJ+$�-B���R��$`�pUQ.AG��N���8��M$��(�Q3��%��F�U[�3�|��<N�	3�V��b�m*����Ʒ�a�#e�ʕ�Π�uz���ھ��l��ͣ�I�u�X'fJ�j�oe
r����J� ������ a!���6�4�Y9�s�n�=���Q�V)��*�uhš55�b701e1��R���9�f��ʀHrN
�\q�-g�3����t�M]�Cw�s���E`}��a����͉֯-��
���wH�=8b~�as�|�Uu�ks�!�K�sqEw�Bf<���J�|�RqۨzZ���pG��]���S^�x��k���;��E�Y���A�{f���QbU3a�K �u����y~G|L�*�m�s �04�B�����?/(!w�:��4��M�k�n1d��d��tKԉ�m��Y�@a�g�N�<�F����!�ܔ:W�m��<O�@��~fo�~��7>��ID67�{���-��-ޔ��¾�+�P���?5����$�<@���R� ��e�&�*�?y�0(�c�F^�/$}��G������[n��]��[��7�6��>e�C�Ȅz}��J��^#`5d��k{��l��t���A`���?��7�B�n�?�z���[�ܣ��8<:d0�ǐ�˻o���"&6���x����%F��jR
	뗹��d�n��d#� 9�����̮g�tvrJ��_��|;O8֎��$���Д�� O�q�dkN��X���MY��
�Y��Ӛ��c�n�TZ�םpf)����`0R<ܗ���l4�*�k�쩩]��٠ް�:�	(��V��t��+��h�cp0yp<z�������F�vC�#��g�&��%�v��@�>�L���@�Cw>��V��x�<�\�8 ��. Ѩ��+Ss�m����w��5f��u}o�"�Z�b�KaX�0�n�@o��i�;�"ª�6������׿� ?y��~��5�����o����OBđ��pB����e��(	|x��"p�����% o���:�w,�N�gߤ��Bh  ��	�E��V�n]%�����خ�-9�< T�u��v�ZO��6��&י��Ņ�|)�&w��9�!F?�ۛ�w|7��d4J��а�W8w��V2׳˺׿��ʧ4b�9�`%l���\V�ZI�E�k6G.�8��\��wd�tr�&-@��|�\ j��0���k��� 7�%V�J�@����U��e�����cϹ��KjR���8kT�n�Ǐ�#� WY]��!��� ����~SE��w�w� OB�Z)y�j��v��ƒ��e�0XzwC�dB뚎�[g�*�����*A+-��z��%��ؐ��/vp_�T�ǟ��%Ɍ���<]�ߎ��9���;^ˀQ�l��Mjk���X$b��WQ����j�Ĕ�{��
Ղv{��6��6��9'�y�N��ų���%]�.2#�»pǻ�^����Tgk�dK�\d1�Q��EwS׆�H�t�u��$nض9{!s�2�|�y۶��U�=���r��]I�ҷ+������dX�V|���A���UȚ��᫕x����w�w9Z^31x&U^d�D�����|�j,sL)���_��#ڰLK��A�n���}\�'7Y���+%��1�<�0p�_#����,�0��#�7y��)�g�`#�{i����< Ӗf��GT�u'~�#����U�Gk+N^+�9���Ol�Y�q�J���5��Afll	5Y��]��~��mk�5�ü-��Ѫ0���f
�� r��f<���)����
@��.�ͅx�1��(�,8Z�>ܱ��' .���	��h������[�*��8���j����/�� d@��m��>���BK\�����Z3㚧8��A�(\LhT ��*��K$S��T��$�@]�Sh>c�z@'d�z��7����E/1w�$��� �p����M;�H��g�=:sV����D���:⽦�f0���c�ϜA�u{�ܶt����3�����<7�+�����{$�j� c�d�ѳ3�_��N�ɻ>>%���;I�^��Ѭl(S���Im�����Y�����VJ�\k;���9�a��)l3x�̻]�IfA�?I���~��G:~~LK���u�;���I$ �7����d#O+� �|�u��c���_b�?�X�h����`_#�Y�(�9�Y�G�����Ƶv�Ah�ft�����tV�	c�~�Q�1��k��\�i��!��1�#{[d�����h�Z��,S��� �X�٧ ��8~A?|�'yz��-�����32��wB��p��v�������A�u�����.� f��[;��3�� PB�<Β.�t��9(���v�x��肠��Iy9,�%�b�!���p{4�׈�����lG#�q�q���Z��]�n�y&M�z��=�<��y޸w��®�Y��7(���J��L����r�uݑ+��E�rݛ����"�aP ?�4���1�1RM��qS��j�&	%���K�(2�ԯ�4I�czq��l1j�rb�ժ�,r�ۛk^8�p���S	�Ty���X-D�����o��y��	������;�t\C%LKˣ-�|��^;�^�P/���[ާ��gفk+)�����,r�0x�lo�~�Xbc�a���F@d�Ɇ�yosd�V����ɦbk��P����_��G�֗��� �F�h<0f�ٻ�e���l.wN�ʘ�*l�+�6�fݝ:�A�!sw�i���r�sc9fzk�C��O��<̓�;����A+�Z�<��W��D5� (�eæJ�ƊCufi]Aܿ��1{�Kcn[w�#Kp�X��5�J<���ܛR߾a�&b�y�D~֮W@��R�.��x�z�F׭�w�
�ⱚ�X�r��P���ת��DSo����V��e(6[5�g��\}��|�,��k>Ǝ.�����:�z�X��`s *��z�i��}?�Ř92�����K9a�uŐ��_I<v��j|e��(oTyH�>#{�ɭe����R3����s��dc)*�V��u-l��:�aX'�˒�0Xدn�aCh��!�{�ڴ�-n�I&�~Ir�^yՋʣ;���rJ�{���e�_2b�y�!��l���`�_I���$��|�X�n��`�����5���tp�R�C���x�K׋����w��S��� urrB޾c� �o{g˽t�s�68�oy�봼q{#�Nn�
�qإ{����BL-�m�ؼ�d�L��4�i��\��=�V w�lo���ХY�El��,  ��;�`�Ƹ�^��\;�`m+�ۋ�l��EX;�`O$�Z'ա��k�mv����2o�`o���-'�9T�66�L��}P�2�V��X�6:���%�
���x��G_�7�~�����O<f`�1Șd�ݝd�2����=�uq��� j�{ɢN���c�;����v*�PN�hdZ:y��a9܄�zJ �ץ��k�I�����w��>�|��nL���R�\[�-L�x
�ℚ2��0���{ǎ��}�ʪX��k$���`�)c�x�Fh��j���ЇL,���و(����G�1�ؽ����ګ]�^�BbT��M����ʮܺ����A���$^qb��1w�m�m�NR��� �/��(WQL���#�|@��3��ds{�6��M���eF|�s�#����{�"��	!3���mj|/<��`�c�&=�6��*c�;@�g����8xx'd���0I����Fw2���!F��R��-x�o��0����:�,�ǋB���џ�6�p����켙Rb��ε�A�2��\�1��WlRA4�
��7Ea���0+�=�r˥���EF�teǲ|U������/,��Du�����q�s�!����=�C A������`ޕ��x�TE�8!��0� Dq���")�Pswŭ��=~���m��]�:��vk�"ۥn=�|�6���K�#�Ju�ޚ��fE[sp�z���u*3�X���j@��r�
���qW"�d&�\�sI\�E0��v.��:����b����/ʎ׬V＠�tNa���(�S۸�6~�Z�_�7�	�P�<���X4B�(�u�Ag	�c�
��=��%Ozh���=LAJ_)����q����ON�U��<�L�j��u��b^/�b`�L3�ilTNc;ˢt�.{-`A�s\Y2���%)�X�eŎ97�`2��J�b�JZe荗Ae�X����]u��O�2�r�]��U��5�U�E8V���K9F�f�'�"�?�>��:�}�G7B��ch���[�9}���w�yM��v-_% c���F�Qj�8��e���L��h���"2��4���Z�&��K����L���*��G>vxϢxq���i�1��j.@�����(�kX6zp��q�Q�ܙxX��^-�:�árAe���q�F��6�I��l����fcئ��vĩ��A#�9��Y-K���.�4�1�!�X#���=�b#��Iu�1� �\��<��;̳3go�H/.������ú��}�G+¯����`<9�h�t�M����n/���P�Pl�|e6�A�[��Y{��*�ƙ���iߥ� t\�2p����/4|�V��(q׬g�ݖ�{��6x�0K-�6(�	�i�謜)u���5�v^Ã��>�|�˫��u�9����<U�����@B�,�{�>�dk0]'�ᴎ�� o��C��C�W
$�4��D��J���ӓ3z~|LO�>���t��������t{#ˍ%G2 @�������' ��Ì7�S���u�9]I�/���=|��1�4spK�;�->��ή a��������O:�����m�{?�|s�WO6g?�P�"��sl�r��Q
����\�6�7@%��cGf�p����Ҷ�ԭx07]�;��oN @��W���쩱#�@D��w�̏�����:��^��z��ޚa'�/Zѿ�y���+��F�*����M �EaMt�g뽆��Қ�5�K�{��a���h�y�:S�H�3��ޑ��*z�Y$z�7Ү`��� /�"GZq�H!�\���T5��� ��4�M�@f\�u����ƪ,�=
�3�Q�iLf�t���쪊�b1��ߗ�tˆ������wx��q:��n����xqvNW�twy�g	o#CvYV��9Ь3�*��$*C�,�x�x$�Rtra�g�}������U #3���:e�02�i�
�
�&tAT;Ǟ����P��X0�Sv7�xND�$c�3㩢�S�����2[5�x���6d�VA ����C_�9�+��0�l��=2W]&��I+���(c!�l�)8�< E��/l����|����B�1hb���sGf涵��b��d6i��Isr;)��s��ۿ�P,��+}B��B�˶\Y�B�	�g+���J�(��:.�����Ɛ<w���C�C�fl�2�g	)��C��ʤͦ�L<9�ڒu�������׎C��2v���8�g�B

&�,	~��e�(�֯�M���`�	�t�):8N�����$����H[%��pGŰ��:��#;�0W�%��t�Jە�}�����P�w�
0ϋ���m'�d�x�3
��\;$�8��n�ٙ�36H ��Z;Sޞ:P�?E�/���ϡ�)�=|�~�VyR�@�w�L�i� a�Jh�3(�o㞵�Ŋ�V�_�+/I>�b�a��*N*D{ω�f�� �P�G��l���e���s_�hy,��3v���ʥ*�x�-
er�0X��>���;+�|���u~Qt̀��;�b��&�\/�)�3�F=�q�]=i8�@á�1 ER��:�$�U.@ �g2=D $�tg��F�H�%��� w��ó���嫗����$�%�C'�I�(�N�ï�d���{���I7����,�6���zT�QA<�T赁��-��ن����c��ysk��~Cy����sDCz+�m��9Z(P�Y�f
f��A��J�`p8��-T
(e�A(N� � ϙ��K:;;co}D|8y��t2�")�p_(�4 ����/�����]�TtoC�
עԎ1�+�ժ�Tݖ��un�;B�[p(����)�TG�o��N��68y��q¡d�W >'ۜ3�6�� mP�'��$",}�)?s$�8��̢�@��y)�Y�<J�R�b��7?w�tpx������y����(�ڂ�W��-%�c��ϸm��t ��fU8�����<�2UE���é{Z�-g�znk�����QFD�@���0�E�X~��Ywtʭ+7�)��B~��٪ �'r�x|�
v'-��8T4�������C��ŭ��,t������䤟��ƫ�� �0���m�x�¤>~v�:-�
�I�E��f�#$��C�b�I^��OvL�d��yM�u�B��5���(7�f/��YHµr{w�� %�Hϻ�I�<v�A@����KI��$� ����޼yK�U���6-�t�;!�� ��!t���ڛL�H��%#���B���4�,KY���'����p�,�v���s#�_�<?��ޠ�H_�i���l�w�w��vRv�#����F,z.d6�N�e�E[����A;|)��S6*^��N��r��]�kÄ�=�n�2dB�B�x�i����+�b<�ȗz2wE�b��47��k7)���X�}2��*v[�3�xz,��
��/\3�q���k	��]G!gWzU���;��l�/�)$ �L{1�k�"��J1c�<�Y<��n)�0��؂�#��Nt�Z���zAÓ��&�[y[SNb���u���"�:����O����w���Uc����*�l��M}^�a!~�=�_牅}�cc)��3�g	�oa��)/,�]�y,W�O6�P�v�H�X�
0���!�i>����Բ�f�����K4����l�4_A�� U��:�Y�5٣�U�m�J��"�BY�o0@6�)P& YG� ��\��7�����,���ν��+�G�R�:"�m�@g ɽ#C*_�%���:���\Q����A�jD�\��ly}�\�:����B:"_ 1��T�˴�������2\=��hs�l�5�R�����J����k2�T9|rȩ�b.��J�I� ��8m�A%��� ���^ �yz=y�Š0�Z�N��/�[�g�^���}N� R[�L4�\i��YU��(�(x?c�f��*�Yy�ܚ�4�L49�HcÌ	��$M6gRB����@<2�ɳUY��<������ry��r�9WI'��6{N!l��{�x��t��`��M���L�R�f��0D�Q_���Mƒ4�U]�yJ�.��\^^��
;�������f[c��׿ү��B���'�8�H�?�o���TȊ�s�8j�Q��ȞXQhxА���J���b���7�K� ����v����˗t� )���9;(0�=d:�/���ԯS�N�N���΃M ����=����lV^7W�tx�qH��[�[cS�p��;�d�#���؆���]�?���J� ����*��v��%�N��t�fd���kC8�f�&G>��
R��ȩ4_�oV.ƭ)J�C�U�P�L&�س���8�"�����猶^}�d0���JH)�����f���,����K��9&c��vQ�����B`���w�E����Ъsv��ӂ���C��0-d@��)ނm(`.PO����[z��("�}B�_�'��}s��S �T�j�v��N�S�p��Nɯc�}��~+�]=��d��[i��+����aAC��gP߈V��}a̓���a�c?���2��Px��Q#61/���[8b�*�b��H�u*����GT�?���NRİ�A����0����45�97ބ�]\=���)��q��Hs�b�,���i��%<����hg�kI)b2����>����$D�'���ٸ0~�f���-����c瞝��))��r��	a�G1Wt>W
�Tn/H�0���}�8��������t�vp�NACŔD���SF�Wװ�`6N�8x��F�1 h�:��|Y1p;U�>�zy!H��;�S�B)�e��D���V K�B�(V�ѣWF%+���!�H�T`��N����_�l��|�l�&�u�̍g�d�����m
�c��(��_
��i8q<v]�����Y$���B��[v2G<��������w?vg�nD�ԩ-�{��n:7\[]����1���s?�0���Xi�9;�9	�8c�������/O�s��div@��x+��n7��i�F�y�����i،ΝV1HX�J��F��:�=7z�GN6�sYx�����ˍ6KZ��5�=����n4" 6��I�$촍�ذ��|s���8e�y
|��H�ײZU���4Fh|w+?Q�4�S�fF��PA�Q>Я��ka����7V�xK�F���Lh� ��ACpi��|��a�sv��2o8,�S��?�Ca���D��J@o� �`K����.�pz&Q����tG���Q�#�o�-=���ڹ�=�5ߛ=ãn�R�Q�����R�Q 0!�F��A:u���������i+ҽEp}	��z���F�>l�ݍ=����BR�om3�S_��6���cmP.��eI��u3���1�z���&{�ɓ#�ڀ�6����'�ln�r���-�X��eo���}�c[�^2-�Ni�l6u6�{v��.�pq^���٪��>7��¸�B��<�'g�w��������z��T�C��GB��_��y)�����_�}��#�1⋹)�D�7b�(�,��6)���(��G5����$A������(I@w�wq��]�d����H=�=�O�_���AR wv��8	���ү�_g�V]��d�K��3�zw�񆮒1|}u��O�-��uI7�0����V�:	��$Q��孱�0�n2�����Z�u�X��@�7������>��DL3�=�9�,ֺ�gBN 5x�hF^&�9T�� ú���@�;�=�!��o�{w_4�0�Nw�CQXcʀN�\^���E3�c��R��0F*����ȏ��&�I^�3�1)Bx�*iI�),�PdP�V�8����������o�vG,\��l�כ2��Ç��I�}�rZQ^g�y�>��]�m�P����]U�X��i!\S���;�i��ڠ��m��٤��9m4Kр����ϵ`$��/�b�fP'���v�Li�d��2/��\ ]���'�]q� O5�?�g	��(V���~[���r��nы����g4	־�<����˗�͔>��Ez��lh���f��:�;r�zy���,�X��C
쥅C�n���}�
S��e&
�dˑ���3:�2��{���5UU���0�Ī�5�&Z?�s�Æ:�A7f�Y"��X���2/�[w�O���b���ݷ����2��A���ͥ�b.�@����JC����k>�,��u��!9��R`���
�D���<��0rMG,���s�� ^�B��u��� ��)��ԡ6ɻ� �<����'m�eq7S����<n9L�b^�ܲ1߫���Ne�
`�ɔA��潄��S���h� E[I�g6���6j݊M��0�$��֦p�D��?�E��MP�)x���~�ӓӤ����l[~Dy>�����u _��rtx�	LĘo��a��<�����<ݴ���#\<9�t��l�����3b�h$�Z�Z=JfE�"�o�����j9���D�9�d�z�Q�w�3ۡ�٦���9[- �H�Y������/�vqŤ���� @��h��C���U�0��{ިF��6�/�~�����itP�(a-�}�z�Tts�S�V����w��&1)�WH����M�Z�؛�o�I����/���)s��^[�ۼ��޵��ު�����|}a���,���6����}�ß��o��o���AC�b�������3�)���~��7t|��N�NY/�I68�0��r���C2��Wj8^��`�7�M�,�~��\r�P	�>� 9s!�\nhY��e�)�����+_� �ӿh���V�;T���Ş"_.�=����slq�,�"��W[۴{��^{찾�Vx�`r$�w�(}wttD���������`� �R�G��ޥ���Nk����W/��ӧL���cč^�k��O�%SP\��׷����#�^�%C�yR����g't��96N��X�m��Bh��E����cl�xRYt���3`�<aN��iA�л����p�+H�pخ�er�6��(��yB�����}	��NϺ��5\wN�cǕ]���Q
᳸�6�� 5/	j=p��l����#���B���9�S�:sG�]�e�T'�!�L\{Kk3�2$�F���)�8'�d.�4~qM�怸��2ȡ��Z2|P�?x	����BX���>����C\�k͛��l���-]�Q���?�7TaZR��m���U��Μ�v�	vb��b!��k��#y�:ԑ=B�?d�����Iv���VHusWJ ͬ�v�$����VɻC3ΈQF�=�[x����TG= �Ǽ����{>r���k�Ȃp��e��J�}"�P����V\�F��_���RoL&M�?N���e�~M��������j��)Hg�We��@�x���P��n�ca�&����1]�$�� ��L9v$�B$
}Eye��*�\_���6�VOc	�_�LȮ��j�����f�9akv��f6��3<���bv$;����W�X)?����n���c)+{���^!�J����8m��Q���5k��e�����R>T����6.ôy�2ؖ�J�g�F�	U�yޚA�7�T�S�f_�b��%�Ⱥni�����z�at)c��+5*C�`�o���ق�E�3KuKIۼb� �W�V��o��3I2ʌ����p����f)�O��|�������#��C��5T^�.���[�2Gx;��	%4��^Ⱥh�(8�x���n���3!�6.\#��x� ,�Y�WX����Ӊ=�S=7VR�"����S�/d��fsϖ��t=��6�-pҌ]��p��lG[r"��o�aL�g��ﯘ�1{�T�e��!�N6�A�4�;;�a�X�\G��ܻ��1�2�����il"Bbkg��/*u���y�$��e���_J� ��V�m� �6!��&[ �B��-n��>]5�{�IlR� £�6��������[Ћ�-��J<~�l;�q�/m*]�Y�+�_�}p\4LY	��BGY�N]V>������j�1� �Î�A6R}>�c��'
���*���~ߔ�����k��N��4�;1�v,O�3`���E�4�vw����_����Á��0M�����1@�?���VVp��1鋗/��7��K^7@�o�R0՟��1Hsvq���֘�c�����������k�Z��?�ϯ�[�؃��{%��Ͽ�B���cW��Ix�b��f����K��ߘ+����ȿ얀�Ub�u��*;,�Ko�0�\*5����N~�X�����^��N��_����
��綐�2$ρr���^Uu�w�^A��'����e����!s���v��!c�[U�(f`n���n#f0Y�ͤ�-Vn��Š�=/��Ȏ�6�
Y>���Ӎ�m��e�M׽�kH˵��u��Gd����a�PԴ�2�+��Z$�pA�IJ$�������ӳý�]d��Z�[Qbj�0��n]x���R �@/�C1�*����Eh��x�6�I)c��Jv�,�&+Ǳ����󎻍�@k���)�L�ȣޜO����㙇JpG];��md��q��+�ִY?�v�H澒�K
l��.Q~���e���nGݱaB#@��e�M4D +9	k5Z1�,k�C���Ʋ	r_o�b	i*�.G�oFphj8��(��A���q]9�UN��c�[��*���󺇂]lU��*x�;3�����!���=�B�e��P���I�6�z�^�@`-����n��7ɟ�v�+�fYv����;xm
B���XD�a�zk���
��)H�W��aӦ�R�D�[E�ڦ��q�@�ԋ�M���Z&.�����G���F9޽{Ko�����t�R8p"}��]i�&��H��&,����w���￧���,۞%����=뭭M�2��{��FcC6�j�}�'�<�? H�~�ٌ�Y'7�8��d��������9�d������ W��B��no���{�"4c�x;�m��ٽ��Z�d��m =��m�t���/^��$�yS�R�i%�0F@<�T�	,W U@'���S���ѽ��x�P�KVE�B���Z��W9p�k|���J(�� �޼}��E�q˅9N���I���O?1����¸`���+�\ 4N:,��.���J�Я$Y2aqyS{ ���l2�@sx=}�����/����o�����-�Ԙ�5ޱ �6��Y�@����:xr$^=�v�m�+��a�Y�Y'�.���t����N�AϮh��-���2=[�r0�4���U��|�̽�>p`�{Ҕ�1�g��������c[�GN�[�5f쿙p��i�+�����ƌS��0�~�' ��ޔ�)N�HbP-5���.Y�A@�a_	Y��d<a�,>��r 7�Btq�Qxx���M�,��|ws-Y��}xϬ�+��>��c�1�P�ꜥE�^ÿ�f¢�]�fuɱ�Pjb�X1洁Ku?W��E�q:���|_}2�۱(w^�/�� v��P�f>�cS^?�Q)�=��Y���U$rv+y+9U�)�`��dF�ǷF�ͿX��t@2��U�r��(�.&#�k�J�w�IBmVX8���[�"/)�y������/ԼH�9��� �U\�2��	��wYp���q�A@�X,2e3��Aܭ�V��k�/�Wy�����_-t-H8L�h���}��O������n�F���2?Y�פ'���,�ɼ�A��s�y8ˎ\���b�I�JKm,���c�L޴�y#ת���'�6�E���o��n\sd���������9�����������Qvl�܋�AW����Sr��Ŗ�<\	���	�Tʡ`��{Y�N�YY�l���oR��Kk���T���ᴖ����3��K;(T�Hf$�}�X�Ĥ<���rv��{3Fm���Tl�8����bn���*6� >����k��&�+����]Ƈ�ԉk����FN1C�AE�xUy�,5�K�yа_����+�:��Z�r���."�� 9�'�p̯3+�u�}����C�I9����D��ѽr�#[���R��e�_�BC+I���+�lG=r���N�y�9�l���Y��ԩ__t��1^�o�O�S�m�,�cc��Dҧ��u�̝��n��g�L�=+��S������@ �12�,�!K���M��.�d�
u�A��dp��|�����L���뙶<z�aYm�YB
x7�T�>f���.8_�m���� p�3g)�!d.��߾}��C�޽��gg�m�$��.`Ǭ6�7I����LI��_�@1��V7��>V��t���Me������|N����mU��e\(7���g*[�l\-W9����tI��čZ�(mu�A����\� !H�t�}�\<:���6�mﱧ�ֆ�\__1�1?���Ͳ��ʴ�����^ qf�T���F�7���d�j��<�/��~����9[{�,�d�Vw���P�%��6�?6p����<&�!o���)g�B�a�p�y5��ۚ��0ә��G��/˥5�ot����L���؈�P?���M��Un���W?f�v���B�y�h��a��U�{F��S_Um��w���s�|o���gXĨj��4�ɖ�X�7���}x�@n�ID�n7Mč�+�W����K���?��`�Dd���F���>>�'Ϟ���.��p��bp�I#�C�H�D9�wZ�Av���t�h&jN�Dl4����5������g7
�p�)�h�&:����	j+�3n�X�4�Ir,.�Y1��v��qJP�]2����I�^=��ﱈX�I�ή�mY�����*%�����w@ݫ�Ua��Ks�<���V�{&��,}y�mb.�N�L�ɘ&;����J�/�`o��[��\�-Ӣ����yÙ�X��x�᪤�j���L�H�Y����B)�ԝJ�T1���/�5��4n�Z���{��?�G�P�Ts94��)��#t�Y(�c�VR�6��lW���4���7��h�v7i3}Y�yV�i�����g����>W*�h�ԅ��d�V���7��{+=?��R���>u��VZ9~%��\Whװ1�����>�߮��8�P��x�f1��L����Ӝ���ڕ]0,j]-�*�WY����ǭ�k�*ʝ���yLG��A��1����Av��ht�TN%2��z��|$k@����K[�)�m;���cKKK^!=0�|�S��?t�����s�b(�w�ͥ� �غ�)í��<�o=�t�$N���%�K�u��ۛQ��s��
R_�Z@,	�U�C��k�ū�v�ji�2d�m&����%1����\�/�r��12_��0�t�.�ѻS,̧��>��^�=��+�>Fӏ��O�H��`z��T�u�QŊy���ASZ+^Ԟ԰�$ːf�z�R�fp�2�3���&� �O�����m�x��6�z�w�������U��|,���K�ˬz�	�!Řu� !���ʞ�H�_���L�kT�b�dK���ybׁ?P@֜��d@=���Jxvv�sD/_��W����gϘH������-}x��~���d����WB\����Y	iu��˅�kF�:W����l�pV���z��5K��-��w�;�7�g�3~�l��3�N�<��:��0�33��Z�{�����g'�Ɖ`8�g�b���vmU_@?#�
z�kMOк�
�=}B��ϙ���g�I��.=�6�#��u\.�h�C���JϺcO������__�7�_-�/�o���%&ֈ�0���UZ�V�-�z��;y��=�~{��=���cٸ�%{���A�ޒ�3 �������3����@+  �l��4@D� 8���޶4Δ��ѐ-�s9`�a�D�	���M���Þ0�gY��:��:!oMJz[\�+�Ӈ�#1�R����B�)7�?��뎙��l}���+k�����RdD��\��o�ᆩ+�ߗ���@^��s<�(
(/~��e��5�p�26N�<p`��W�0 ^�T�R��KvW����ΠŽ,�뺹��J�$�+<+Q$Y��=����gES�2)i��J�����0�EjKP��cKoZ5BN{��>�bP��xH�MQ 5\�_-?��C�ksg���;�u�]J��-Rc����^;U�lyF�B)��Y��D��-6��߿W�������чX�g��b^� S�*�L6-(��9݊�,/��JUP46\�(���)���L�=g��'���V3pH�K�hň�X�ٽ�I�ٸ!
�"��Ѳ~�NV�Ap�T��U2��`/��Л�����{�4�\��o4<p���f%�#�3ˆ=���s��IϏ�h�Y���Ʉ�7��ib���o]��P�Ck�|ǁ���M ��`��}�W�I`'�t����9�˹��F�~=$��z�P����X<�S���i��r���q�E[ѷ�<��H�{ѣ��>�/��0+~�HI1k\�c�^b%���6��lK�b�kz8���݇ȁ����ש�c���͗�4���$�Q�0���������ڟ�xq�'yF�_K������d��{�wx_��^E�1QN��ŏ��>�~,ך��V�ֶ��K�O��폆�4����}�=�.k�o�6��C�~er��d#�����&yWw+�����e��ac�bL/�>������p�@N֋M��tѩ*Oߞ9o$��ڨ�d�:�������Sŷ�)��.�w�+#���q)*�!dO�*���"������w�7A���\�^�H�V���M��\9}��xA�� ����ՃrB��@K�]z��ma��ΉGv�y����r��p������1���9�}�������D=�������!��^���7�7����G�5n���s����%��hlҁr�x�_��A�8���	�@�l �@�<ʳ�f@���3�x&ְ�B���rC6��|����T��ϪɞZ��㨊�=���+I₰+qJv�a� '��o�?@ x�`��ͻw����p�^�=�+�T�4�c��V��܎+1Ød.�@Η�M}�� M(��S��L��ic��kX];��x���#��ζ�y�4�5���@]��5DN�X�{K�^��PMĽ���*� D�SQ��g�~�<<�n����0��'v(%L�xHV�l~�5��MF���2i�Dc�CV迬#���?"ߩ���?�Q�J�jȿY�0с�#�R�����p#B�q�i�.�Q=õno�\)���&�$y3�E��w���d����U����f2.�c@(�@���G}�3�J�����s^8 bĴ��b^*����ǡY����s�Y-����0߫%�"Sl�wB����̪�ͰUL�ݐ%W����{씞?%`4���'o��MV&ew��v����aS�:�\���wb5ef�UF�KP6i\���	��K��#$�3�"�]:�7(.Xtx�+�+^HT��ԣX��e|A�R�����xqu���6�l�q}P:��/w���v9��#n2��3�m���~x�]&�MvO�i���f�%����_�.���N[t��E�OR��n���2��\{�c٘��������G���.�0aԍ�m1����	�GRG��>�~L�>Y���=0�c������eʉ�� G��-y���c��:����N�s;/6Q��슉�d`�5��;P��2{L��6"�t�ãkP4w��k�'i/cWѳ����4 �;����F^���Ǉ�Y5̢�bُ�⯩tx��Gc�d�,h:�:� \/�;�5m�^<j�5s		x�a���$�d�J��;����:�/�:S�<z"!����G(d���[��崡P�V����x�(��7eCѥ������MUp��s�u��j5��rB�[Y�j��w��A���fY�NB3�$hĐ���m�i�[$����	P��"tAe�ͰI�ǁ��r!�J�-����w�я?��z5±�����'t{�r6'���t��gϟӷ�}˴��`����_���_��}����M`�/��flܫ-���落r�>{�܂0��Y�y����A9�%�dj����� �!�'����K�A�ʏ��K��f�yDW���c�.Kեx�E=��FAϲ�G��l��s� ����z�W/^���1=�6Ħ32��R��ש,/>r62<�H�nD �����\S�G�/$��(��8�K"z ����^7ё� ޚ��+z���+E�D g ���s� C��G��}�����駟��P�>�0*o��Âf��2�9p�5L���6�~�r�h<W�8><|B��zrpH����޿c/"��Š2Y���k}^�&*B����˿�������_����<�����d3���Ļ_7�-3�y˭䫕+
��m�F��m_
LR���K�����v��c���z����u�㏙)��f�L���h��:G_U��!� �<��&P�p�뿗��|s�� Vp86Ԋ>x ���j�.g�v̈"����"�x��L�č��**_�z%a���Z�
�]��#�|0�JB�8�f����(��%�_K^n�b����/3ZBt�OSd+��5 ���nV��A i�"ԩ up����Gk ���;��7뀝���=c�����"�ۢ\r���TZ���G�E{[0�x�����zg������sU�Z���5�[N�?�
���5�`��y_��0�V+�XısSiL9����!ʇ]��f��ϳz�������B���27_��ϣvR�_��\q�B��ZŤm�~R.���ݚS�,xL*%�R��j��IL�� �`a����t@���_���J�7��R�h���F�\U�2��_�pC�1'��g���9Y,�2�c0E�&	�7�c���=}�Ҩ�tW�m����͙�Qe��<0:�k���c1Tl�����m�)�5���p���ĥ)D�>nc���eBY����m�嫝����{ꌓ  9���[KCm�v|-9
#}�`�=]������{ng��ǌ�����F;'�R`���� ˉ
�1mC�����F�̉�ud���YF��:R?UƉ�}�@�X�:�<�1e��9Zdz��Z�гK�;����� �7��B��o6�mn1�b+!��5�5��yS���p����N��7.)�f���"��S�^h�c:v�SB�#t���w�?<}�������?` `�j%�s������3���o���6� V���MA%��4Ll%���g&!@Fk�TI�"��Ï?Ы��$[�z�@�aO���3�@śe[���zh<��~��&Zƹ�4/6�������̽5�S[zx<���z��s��D���\�w����ɓC:~�L��C	�bʉ�d�=99a�����ɇ܇�G���^���H!(�K<@��yӐt�H�ӷ�j�� X�_
���g�x]
( +#�������4.�g�}��	�_�~ͩ�LA߄'Q�d�v�?�Iu�����T�M����ڒ���00�����D;I�>J�������.���/�i���t��%�q�����F�����d�!�@&��`��o�"�<b[��~�]�F�9.,�䔉�����c�m?}���{�P�����}D�^����ߕ��ĵ�s�lW�R��;f�/K�:�����������eO�)����BR�RM/�O%���Pv#�Ӿ�T0X���ʛ��^,�Jt�`�	ɔh3N�9Q���dp��f!��ݠ9²�k�$��@�8�"H��}X�f�U��00%1��p{P@2�̕[�Y�NZͼb D<�k��ң��}o\;U�S e��=vm�sy�)`Ǿ/��������l�B�1凌���"�>��1&cԳX�lpr&�UuV�T���sBA1�M�2�ݦ��vw�nB��]:�]�$�=(2(��M�Y1(��F�=\ny�����N��"� P����a!]�;I�	� ���su�������I�\w}�^�t4����2��xA�d,Ї��<)0A��x�j�Ӻkl����]�����������u^���b߄)[Q����
��Ǻ�x97\���1�N���&řA3��4)�b���W� ���S˚��`eٽ�-c1N�:b#�g��/�,�>�WJ��nܕ;�t�"�� {z�B�O�E�ԙ���[R4f���ډ1W����S�z�9t蟓���t���Y����,� ��>�\�����1��.��Ƶ0��/A8d� zn�  �mօ�y�`�y,�S��R	�ެ��8�������y`Y�u�kx~ßF5@kb{v����Ə9��zk�X5Ǻ��?=���醞�dq�dBE���\�V��I����=1j	�F��'��Yq4��iK�3��H�i�{
R��H��V`�_^'���ɓ��ӟ�s&��|�!7��㏢�PI�۰\�̈́��	�/�8�9�f�&��g�S��mī F��9�� 0b�77��W�������Ke�������k>y�7��'�%}JcB�A/��u{w�ab?�ˏ\&�mm��rx�5N��<H��'J�,6���F�^]n@]g�L! ��������W�"�@�jRy�>''����� ������TP �����>����k��xV:nf止0�9؀@��X�r������kN���Y��b��gϞы�/���s�*�0����9���������8%�ح7%������n�K���2
�i�X�9�e���h���N��_	��`�)���������?~���ч����xS���ԯ�{��u8:b ������/��J����~8��]�E ���,W���m3��Lk٠����W�����+�zL��_�~��5�X`�m���+rf�@1g���Iξ�!ө(��R���K��nh�X�;Dy7�ڂ��ĕ�.���9�ճ0:tVN��@֭���M�	��n�<��Ŝ]�W|y7}V�����+8��~� 2��*�b�p�����b�\ql%.UkS����pC��p@���V�� M	��}�LC�:�ӻ����r'ʮ�z�f]V�)������Ǝ��Cd�j�3���R���9�Ԇm�fTF�{`���B���.�{�;��]���C:IϹ����l�0r´�sv����Vw(@.
�d���d��LC�(���8��V+q������W߼b�	����Ш)�;r.�P�t̀�tz��W�J���5��cΓ�Y%`���7�O�c'M0΄�-�����xVY��Q�dR�_��{����S�ɧ�ke��Ycb�1�zj��ào�ls�-�ugPi-�r�C*�NE=��4c\��9��ڿ�w4��5���=u0�Q�;R1y�`U�\��T�	bsHdH̡XZ�~�[oF�Q�c��������z{�嗄�v�����+�����266'��ţ�[qy�����!}��E��OE��d��7p�Ot��s��e�-z�vP@�:Σ��e�mo��5Kn���
�\>{t]�̓�k������_��~#�z�4�ח����/���^���Z>s�,�b�ǐ=}��CDjd��2fϞ���ٴ��z��:zw�����S_C�C�Uo0oo����)���KQ����o��f�@%���z��&�a��'�q�q����l^�rI�%;g7Z)P�F�x7	p�������!�3KI�}'�0��j��9u���%٤��j1�L���Jh����I���z>IV+	�(ƠT�aO�W���������z/��}�kt@!xԹ��e��Dx.g�R��Z�BC������G�k���4�aU��%:Ay�˛7�MV�r�7�I7����e�?�gP:���G:�k>!M��w���__3�R�1K�g��#�-l&��Æ5s@E��8��6�2@�;�Ж���q�!��^D N�����Md(���g��)BY�F�om
�A-e@�ַ��S*�/�J�߽c��=ɘs���U[����[��nk�y�dY��SGx������,������YE��O�[���>6�S��t+�^�+ڧzf��9���������t���A��M�Ӻx�ʣt��U���!^���l��2LǕ���IZZ�L�$���u@�3"�R6"�͒dO�����퍜�)C!L��lk�ǀ�7q(3��x5RZ`��+*Q��~�^I�߭�YL�ȳy��ѱS�݁6���gn��a�,L ^�nb���Ho�n�ٓ�Z![m$��h�N���Q��}�;�3g�Dd�N���S���GP��}O�1`g�|{�����*�Fy��C�3���d'��!r5V�������U�xv#���g���S��zrtċR��xl�~�7Q 0h��J,���V�\�K.��V�[PO�Ca��]��<}�~���#RY�>�g�$��Ǆ�4պ��X�m�a8��0w��`o�J8@����K��=�,X���'��߿��y��]j�gdػ���Txc��K�c�F��x�yq���4b<v�L}���BN|��M���?���~��ܪ3 ��s�6	Nh��t�c�	C#0k3��8Q��\j9y���'Yt�)�8J���PV�1��鷕��e�6���O�����/�"3 ���t���K��P�4�����qL������yS�&����'���� �eQ C�$U}�c@�\�� {f<$zB�P9��¸�l�AO��b^����'"��/�2G7����ؗ)cu K=Cep��Szx�Q�㲿����57�m�]� �+����o>.���e��#��?2��G�ଛm��H�^Z�Z�����~é�K�1g�Lfۺ�2{�Wt�t���?3����������]8-y�_�gS��N���I:3<L.�?:�0�z�Yz���.l�$6B�.`�> 2F$6���I�k�����/���"�O"@a�<Y�4<��A�Y��?x���ʇ��<k#��h�F�.)�_��m��Z�MU�d �+!�F9 ,|�������/�ޚ�v���[�"��6=8<L}p$��
���H�#����#�l���c�g%���	g[�����Y��6%)�����2@�)�e�.	�x���$@�� B{2ǒ����������0����m��s{K���k*����)�Q3IzÜr��G�j�6��q�Uos;ö����_����F�Y*B����a]͊�˙�53,{�����t��&����:�8��TN��[�.����R��~����L�m�j[l���ޯS{`C�/?��,"H��˻�(�,#E�u~T�Ǟ��a�n�������Rl��2m�ͷ-*��c��6R��5����M��Z�S��'����@�{X�����GoU��t��,E���vk���#\�,b�I��j�9���_�dw���I�pY�x��ո�	튴w��O��p)0q-��f�
a]Kk����/��n%�����ƣB��N��q�@�בz�u��Y���Uc��uX��1 {���phj�6=��e�*ߗ�\������M,�W�;U⻶��F$����3ި����r迭�/X�����<s�5O+,��v��R����N}:ox���F�q�i�u�)X
����5 ��\���EZȠĔ��L��.��&ݑq��y���V��Th쥟<{>e�jN�~����&l���͛;"(b"��OM�9�e�F'�ׂĢ�#�N.Ѹ��� �t�s��D����Œ�;�kSw��֞u���Ͼ�<y��o�x#����(&��v�R9���>�05dw��[N1�ϧs�PϢ�0�%�o�xW��f-����10��^�|�[��H�㎐��Xԭ;�ƮY�ɲ��^�J�=�:V�g,��G  ��a���v�����b��{(>w?�KS�R�;քu�O寣�hCa�M����#�<��T��9)s�/��75�����)�<���(҈�o�5�+�P��c�NS���_�ͤ[/p �蕪jZ
�����*�rP�M�4�V�CDǨ�,�������+�|�$���=��C���MT�{�&� 3Q�0-���Ɖg� �B�ή�!TB��8 aeB^���+M�O�"ey06�Y�Z��o����tvz���x�l*�0�) �6j\c��ͽ�|�Mg���ܨ;x�p��S��nz6�{�R;ާ�6������i��:���A�i� v�_��:�w�o�to5�}Ʂx�UZ3�˟�������l\�(�r�Bƞ��P7d�� s�^�s���D�_]r��J[���{t������sz��-ݴ�VnE�}�m��p�]�h��6���P�p���x���	��ݵx�/f���� C������Bs���k�;l\�3Y�m�2���l���t�G3�{�O�~�pI_�12�xF��I0~l�K��zK?u��5,H��Om��>~��>g֪����I�9cI7r2�*�,�#d)>q�����s�s�����~���S���G:^��R���#���)��%�2����َg�zW�4gB�<�R�"bh�����@�NjA�5R�����a� !=�����9	b���<3�µj�uA�+1ۊ�3� sF��I`Am8+�� �)�p�0h��{o�['{��3���ߔ^7vN��'� ����T�|6��)�%|�$wJ�kKp�vUp�wMɭ�Yx���Y��7���)V"���XVA�����^Nu�\ML�<��y�����n�7)h�+�L�1*	���H�cҹ:���>��;�hd��[�}[q��X�y��vu�䕄�؃��t�U�ܟ�R�S�*��o;ą69>�z��un�G3�j��G*��	.��o�� ���L-��O&��8Z�kWQx��\&��L^>��+�-�� ���?�c����`d�p�[�M=��C��t�X�.�8��~
���Ϗ�Or����~,���u}D�a,>�m5,�)��A3aЈ�ݯ��Oc�)�Ԡ�����p�X�]H'd���
�,�.�� ��}�E�l�����Cd#}���|�cc�S�n�9^U�hv�w��S�l���bgn�N�ɶ��7]�sZTO���E�s&
h���X��8�B-�X(��Asц��gy��y'u�Η�n��#��r+ތ?"�L�up�����q/ߠ�U[Cښؗ�qm���Z���=��i���5�vu���H��3L����yU@#���2�2�c�V&��� �+�7�P�,T�U ��\)�/?^0�.�C�`�/����� a�Nk�V���FI�8l��of�252�|6M����L�!\�>��.^LP(�#�lM�I����zB�pMҨ�����W\��^��:5C`��p�e}vv�i�ц��o8J�<*�a]I��g6簡Z���xH�L��s͌��8�,H4ʽ��_˂k\7;�;����[�k�#�����]�Qp�C
���k(
''�D���R�4� (��A�����c���7�e~���@���u�ڍ	�� �p+i�>�
��O?���i��y�m�7����a��r�p���!#:� z�Q�.�jӘ|B�����}��ڑ����Tϋ4�����y�MN��7���٦W�^�7/_�MN��퍴���풽����AUm������5�*c�@϶�f&r^��#rbp<L`RJ�`�ӵ���P-��JpOHv��E��C���I6gq�;kf�e��V!�UlB\��E�ؿ����n�)s����~h�\w[������Ӱ#��a}j$~9�`�_��ϼ>�$(�) d�����JX�
���A�|5c:�E�#��; ;�й��=�o�X�l�8㧚ρ �p�b%r��8�U�l�4T�ٱ��C��B�٠����Z.$����%P�ٰb��f���-�wL� �1��2|ː~�k���X`�<x�8vp�oV���Y~?�>)/��z��Z ��eeQp��t�E�0�t:_r�p)G����+̺L/�C�����A[ȝ-l}͛A9����.�7+�F���N�«jku��n(Z&X+GŃ=a��jL@t�=�3i�Mz�x[5쑳QG�I,<v���xc�Q|*ͪî�m6�CY�}w��n,咮v�FMtn�6�c�'�{�V��D=�ldk|6<B��;*
�%�^D}�A��=�,��q���]�Y���S�[�r=s�T;1\��da0�-��I�+��^,���t�.yo�4���r�0�c���M�\k��#�m�+��"��y#=p�hk���A�~=�
,��ظ�VM��/�C��c7|���t�5�`�(�$�w��P�h�8�������Џ�\��s�D%�x��b��'ك�I����w7���g��v\�,dt�Q۠ӆ�A�-����W�'_�u�k�Lq%�#oHvh��@�p���axǼvz�v8 � ́>�ټ��'%����C:;=�͓-���fP�<�)Z�x����W�����䑙��0!�����6	�G���O��ș���,e�^9I?}��9�Ȁ�C� �Э F u�f��A��Az���t�9o��M霍�Q�2�����_3�'d53R���-%���T�.��4� ^;;��{/�TJ�lL��I�����o^�1{̳�Roq�#�����@(]n�� �F��-�}��t[p��$���7���lc��J�G4Ahk�����db�4�P~<�߸�>�'x��w�^�����p�Y�l��ŉm�L�]6簴�dJ_	�B�d�Ёc�Qf��q����S��&~j@�zA�Q{F���=y���B=���NF�=Җ�lmU�W�����Y�T�ֳcf�|5��hjk$I���?����U��'�zD��-1��W}�c��� (~���W	�"8E3�Ů+��5�we[v��~�ԩٓD2I�L0P��R[xp�"`��Բ$H5 �FS��k��o�{᳧�8�gw@0�Z���q�mZ|n��?�+%9����Y��DF���&/ �&���84�r��b��%;���c�!%���kK�ff����8P�|̈�o^x�m��!�X�s�2�m��)@� !X� ���~��1W�wwܙ�y��̇���~�.����ΔP����W��1Ѳz�)�?;J�?�!|Y �[��am��ho�S��Ҁ^�0^��m��煖�d��U� }m�)gL6����Ƕ[�h���=����ݚ��_��	e~�||]�ݟ�^IZ���3p��3��x����?�c{�9òV�}�.$R��e�j�ހ$<��W�.r�m��Wz���C�J�W���ϜԝJ� -%tN}�c�;�L	���q�y���Pȃ^Q�u)���G��EU���!c�!���w&�p����cG��i��@*���Ӌ�u��h�O�g�;���2�d=}���$=`Ħ��v��#_�&�>W�F���/n�g_8�O�@Y�2p�,��Ɠyb,�����&�e�7=Y��qvrJ�gg�J{���ؓf�a�b��j�:4s��f����ʵ� 4a���+�!��zt�f;<~f3/;�n�eCⴍ���c�铧��]��'�DOh#����p3����C�@B����Tj�zmNJ���0w��K'����o�ߦ�!����J2}̓]�R{˳�!���S� s��]��dO�=���9����y␠@�۷I����lc v�������î���%����>m���3s~P���Lfi��g�~��Bd�$�E��n�$x�'�R��X��Lm3�~bJ�Ν�Tgx����&����K��]\0y���	�G���'ח_��7���%��N�����%��2��"<n��v�:��'#8�ʉj��������ؕ�rt��#¯�Ȑ����U"���c�]c�h/�}�cMI;���Z��$?��\��]�w~>�0K��X���ֿ6��sU-tc�3GB���u�׆���K`�e����l$��	V�ų�Ab���ϻ$�(�o���"�d�bab�{o�� �ι�U2Z[v��<A.�`Âts{�1ȍe�j,8?��J	�;�����b�N�����q�_�CL���T߄=B�P���S��@؍���}�=^x��snz�
k��!�E?����nP � <A�,Ȃ�=S#��,?�<C�_
�e�C�更���X�*!I�J��	��Tv�֝!|�]+��P�~����;gG����#�y�)���5���>}�_�Ǯrjʷ�E������A��=c���4���u�R��X�U�8 7(����Z��F�ןxh%�l�~��g>��I`Z����ϗ���1i�S��G,ײ��3n��o�������R�^�>,v?�u�h��������@�,�[��n
��.��)o���[�4�����y�9�?���2����eb�m�������ﱔ�)PH��_���6ͺ��U����|(���5����e�y_2�����oe�G�އ����C�	ЩSi�z#>�S���[(���d}z˧��1�D���p���Ƽ]������ma�N��D%� � �E��ON�3�3�\�{��!	:+�c�u~~�d��y���$=O�v���6C�0��'���׆yk��R�-R��W ����{p��>ѦחW̏�>@���WH6ٶ���t������(�I��<g����.59�� �e�.#��$��9�l��w5M١��H@���قH2�p�B�g����x��{���М�}q��M��C���`�=�$��WvT(#N��-��=��:�������s%!�=�e f5�𺕁kjW���f;  `�mXK��f�͙����J�!�s��h�LI`k�y�0(��»���	�9'''��syI�f��u�"lmq��� `���Gz��%'[��p���	X��.x�����Ǉ MB�@藧��{���ԝ��y��p£ױ��]ݳ_��2��<ě1�x�6|���'����N�����	��y�&n�������������P(Bqh��l��ۅ�����C���Oȩ�;�(��>=@-�8N��J�{�${伕�T��$J:��C����� 	K?�=���	��ӳ�L��ܾH�fgc���s�����n	Py=I-��V�6<��������.HR��55F�\�;}�&~��{�Ĥn�k&�<\;����{˲#�Wd*�휱C�`B�)\��� �*Q�S��Q�B�ݨ5���t���y��u�X`XnK�i�?�5w�� ��%$z���+���g�]�����h��%v��4��E�^=��cKw�B��Y���!oBOD!~���Cd8�Y����1��c�yaK��:54�Z���u�����h10�h���j����e^�y.O^�����fo��E���'n׽�gR�[&���a�p�>l��j_�4�Y����M��u(Ճ.�k�!�)�xY2Iiw��3VZ���5x|���0c���!���A�xl�h�0�������߷1���a�a|D����Dg=��t�㌅��<�j}}�ב!S�˰��2�����?P���<)�D�lb��������O�i�p(~yH���'��AU{�cDL�����T�7q��uHh�&(�t�5{�5��dEYSW�y�ú�.��y�t�U�������	������� �B���s��^!�S2��Ի@����^0�V�2�w������F=��`�Cwg��t�:�<��Խ���Fr-h �ܳ�V�I6[�~s�̙����ZzT7YkV����w��UlI �23 8���]7��^˵W����6�?���G��?1�Y���{&FFF��o��}0�W�#t��y���x�)���ˏ�9����B~�� ��y�T2bA���p�}�Ǧil�ሞV���
}�ܬ�'�9(���!���v�� ̹�_������[��������� o�"�$�fX���&Y�E�/pXH���?0_{b}����;����nS�6��_�@2>ړ�c����gz��w4;<����N��pq~��珿��ZS�s+���7ɫ_x��������}������;�/�&W(W�̝Uh?d<�T�޿�_gt��'��?�����~���ޅ�)J�84}|��eS�e��cԒ��rk�	x�%{^7|���O:dSTL�d}�O/�b�?g�p�h�� ��0@1X��-4&�۝<��Q�q16{�����0|LX�(9��{l�GW!��1��ld.����a� �-��3�+o�]ഁ!φhM"��P�J[v/�_RtSW�F�Lru L��qƛU-�00gL
`g��p?v��0HpP�,�w���b"�K���'ҹ����M���%*��,˾�A"�V ܙL��v�de����z��5��$�zZ�y16�S���!�;�_�N��"�$%"8_�:8}��|���ɲd�R�=o|FM�q����	�������a1�����y�� �x_,<��n�^1�L��5�Lv��2�l���l]�-w��]�ͽA/�|w<7���ti�MA�Xz�O�m��	�Ϛ�>�hCZO(.k�U�q
�Qg�l��݀�<�;�m9:�h�T�oQ��X �����󲞸�n푅�g�я�nU�g��<�O���k,���Uv��+�+�w���U%��)��1ka��$wӼw���q
�v�{��:zD�������,�R�N���|=$��l2t&�c�$����u��i�=��U~���~�(G���=w��@��kWZZ�w*���0����*ݕﲩ��KJ���7XU��cJד���1��qs{�!V��}|��=w@6w����� .u�a����g�	��p�rɟ���i�a!��&�s-%;3�5B�k��k�>� h&�!��`6�Cx��ϱ.Kl���ku R!��CRl627���FV�X.�0���%�Y7>��-4�]Bs8�����&뵢�i2l4�Y���*؄{Д�NRU)ߐ�b�$�+}�g��׉�=��:�d)<;��-�q��<�@ic�"�Rg��y#�$�e_�^q������oFC��+	�c�g�ĆĠ�O|�|qH_��~|?q3}ߊ�56(,�J&`��d 	m��H/4	��>�{�u���9un����[L�	7���'<�,#m�@ԊA��+�j4� �� �1�cC��zJ���g�E1d���龇����[��՛ݻ��|}�}��u�q�-��뎪�N�p��p�"* ;[�!����3����ž>x�׭|7Tv<[,Ǟ�V@���X�c�~�1����N�	�"��Ejk��q�^G��˽��4�Q8��W%ի��;*N�9%�FvEv���A�5xp }���	����TNb]��u�tq 1�t~���=|�����F+2P���Rwzs��y���C����g�3�N���4&~��%����w�0����`de�h��p,�c�9(��0��qࡽ+W�ȍ�a[�� 3����h=A�dAݸ�.]\~�R5��kV,�"�ݨc/؛/�:��.��Z������9�<��.�Z�kD��B���Ȳ�bg^G;Mخ���fG���N��
���D@�)܅qMvd��q�Z�}as�Mpi��i���H�{��v	v���q���i�.�Ǯ�|��ѯ8�/�����t���B�gz��f�������0𳭽�����)����Ґ��^��&�Q��[w�0�?����uq����O���>M6$*�}����s�-z���;����<%�,_'�?�����V���|��'��?/��P\�9PE3�xΐ�_�±��I:�I*o�@�y���<;�I�����w��e�������-��0����_�S$�tD6���gt��=?���8t<(�� ���0�O>HR�L��,\��İL����쩫�fF�#��p$���� ��~wuÙ�8c�������ˑ��������݌ya�]ßdO�Q�b�:X�� u`���2���>;a�"3E]���Kd6].ycw2+D�T⥭����jV�U#</u��'�6>q�%�l˨����rH�f�5�����3��K�zX&3� n�7�Ǣ\
@��I �֫u$�F{NVS���3Zq��咮��0��,�nC�{%}h���Ck�Ž��a�E�ɲ�����s� $�>�5M�P�l�i��@�E�4�3��!���b� " "<�Ļ������f͌۱b�&�p0�ee�}�U-�Vp�#�"/��7�w���OY{Lҵ�����ʈ��ہcA$#��-M
ѐ�i��H����|=�,śӴ�� �.��(F�]��T������2��y3���-�g���,|��)n@��B�6*E:���@�m�~ftqh��0�4Ŕf�RԚ\J�Š�M�}ʌ�j���<�TL�@���<�%����]V�V @Cĝ���Ө��2?J�S`�\b�Z!�7>
�Zɹ!`�*`�ۄ��&^k݇r��n`��?��r	L�����mǸ��c���^9pa����7oް��c���Ǐ̱suuŻy(�=�~ƅ�i"ؑ�-?"���3�GW��_X��P8'@�T����A'�@���2��"����>`�������v�1�8_�c����**��B��#g��Y��zmb6/nG����={,�I���.D�T������=����I�s���6IԖ#�M��wf�rm�Ur�$�&�Q!`nx�ɤ���9�̧4s���d�񄷎�
x���q&����u���:�l�\�|��r����t����on��}��I{�A�fOX��������R��ݴ0Q��+��Zὗ�n�ψ_f�Z$�O��R�{�d鑕,z�b��5��{�	r��a�O���<y�%�v�IeW�mvZl���1N�\��o��cض�L����;�^|���y7z��%�S~�	߿�u�4�����L�U�r��c��@�u��{���ٮ�<uU�ˊ�m���2{��{~I�@�Tv[.���_�./�G��r�V�e�H����%M�쪉oF@��ATt��U�j�Iߓ��:�m�a4��P_їϗ�O������iͼ~���X�E:0+	u� gJ=<�Óc:]�ї��{�N2Oqx��ɨ64AP�d"�B٫)��ynj�*p���С>�}�?������㾹e��3�`��$����~��߃.�fzx�����\_�n�����Ib���1��0�q�pX�`%�R����) 5�Zyk�Ay̞�ЗW�);a`I�X�KI�;�k�L8U�l򝞜0�B�$
���-�:�>X����&���5���7ڇ���Z�ս�l^q�J�p-�b�W�ڙ�g�=��׵xX�����aQ�a�� ��ݬ��its6tcos�L@V��6l����:�61`ɩ�׼Ygf���5���mT������8-<<{4��B׎O��O+M���ȴUʺַ�Md�J[�t�r[7�u��CQ��LǑZ�{��5n��'����޲�~�QE�h"u��8?W���%�N��6�o:���U���}��qqn�q��|����[Y�2PǷnsf���o�׬�\Ɲf�aX3���:m7�1�S'80�K�h�zU��p�:�z��3W�[�S��nZ��������}��Ex����I AjX  ^x-���0�C��b&���)�Ä�3�ZL,4̻�{�G	�h ~,�a!e�߈���Y�n��z�G�,1�KVN��W���ЭZ�{�� �@�3ȟ~�����W?a p� ���d^�)9ؓ{�q3�|�@7��@��D�)Yy(9��s }�ݐ�FI�U!¢�Ew:�)j�s$��T�}�F �z�Wx�5��q�J.�k��	��s���E�:H m�� �i%��P��r��gg�)�e�EO1,L1�Z��,� ܖ���@���><�zr6;bPҩ��b� JG�J�����d>��E$���Om;se���2�E��T�:	w�3�
w�;�'���cs��4��lx����:
v��ϰ���w^�#s��������=潒���dO;d����пr�J-%ǩLv��.<|�$�*�?�6�U+���p<�4�F�QW&Y��O��+ٻϯaA�õ>��0�'��U�e��n*���H�>�*#o�2��a:�r��k�\�=ڷ���Sw�7�hQ�a�C(�߈�y���w���	5~�:V��~[�[�����
��$�zvX?��Y綽����ۼޣGi:|�ޮ�#u�mG��|Aj*�����1�2ٝ�tR~�J9oX�k��8�w��v`��*H�Afу�8H�q�V�A{��/gl���<��s{��a㉧T#/̞=� A-��lF96lٛDC�p?��<�	o�c'�H/?����7��6���uG���!��u�ę3'�qL���K~�q�����~���_�=�VW�� 脚O�tvB�����oi��#��/��z(�A�����'�3&�f�B�<>9=�/�Rw �^�s�������Z�/��zXC�␢���sM>��ϟ+���m !�-�M�{d)B���$ ����޼zM'g�\?���~�U�|B�0�Ӯ��}WJs�~a�V��C�i���p*�$j�uv�ܧ���)�y�dH�����Bg�0��L���x#C����j����P�y/�G'4�<��M�ca~��2�����������E�Q���Kɐ�$��h̲QOo�ݤ c����k:hT?{g*��Bǝ�����n��r�����֛ކt[Xw�����>��y7�%QWp���|��M�u���m_��G�W��AO]�����Қ�ҿ]�j)A�p�Q(h�����y����!���1���.�6�|E/�;�)ԧ���"�{�H�lw�yh46\4���$��P��X�ۛz���a4�"�ʋ�pXziE$�+�u�<H��|�iD�l������U��ᴈ�$.zZ�bN6���s��Tq<�WV{jǿsln!��F]
�%�P�U�b�A�RS1"-�*DX��Mj*�so�}�.�3�aA�F�kX����o Q��B�x��ɋ%uر���~nD�%�1�H�v�$���3� �e��#��G�c�xd�Qt-䮉��,��#Ϙ�˩��r�F��b���L�i�@i���3&cc��s�3����z��� 5�I�v���3~n��y��yX��:>��_`"2/�o�&��\�|��b�v� B��bzr8�C����׌X���TzVh���ڱwx=ײ�u��[m����c}���o��׶��V��{�#�O�)��#���3��4���i�&{����ّ;�Y�zKV��CΡX�!d�.�J�j/��kyI`�f/ڝX��c�{����W���ElZwk?�}}��:��:�
L�bF�1��h?t��>"�Za�6NG��u���}��z^tA+����Jlv����կ����EZߎl�n���;j5K�{���q�����so=�����"}! �#��J����c�G�cv�յvOI���7}���^o����u�<v�8�𙹄�=�	�ON8S¯�Os��l�ͬj��5�~?����V[r�R($���y�ِXЬM0�+�j��b!�� X��Fk�s��r䃿���J�S>���?%{������S�7
R0��J@�H�Q��wѵ��Զ�wz��9��ǟ�=�HH�%<��Mە������8/�7߿���؈,T��m ��PX�Bp������{ܼ�S��x��9m�����t������F�ۍy�ؘj4�:����w���1B{��=�^Z��b���O]��Xg� s�����Jt\yǲs�.���t+Rf-xq���\Ǔ�:<�D&F���0�w�d��ּNؼi"]��B7�!:A��8��<r��F�S�(�Z�m���ز;�{�����d�j[�H�IY�R�j=�{��m�a�Ę�$zfe�u�I8��O�������Ւ�:�4��AWdPG�LP�j&\�Y��o�Q ��<&`O6���*����=׫Bc0����-�,7��r���n�(1P���]Km#/v����$ɖ�ω�=�G��P ��̤�#�$גJ@����\vM��p)�+|�e e��#�������s!�� ���\Y\�3`�K.��ξ�."c�;v?���p+Ki`G8f�V���z���d�GM�>\9��h���͓��������Ъ�x�4�x�iˡ�8�����B���\-�� �P���d�����:]�dA�'xqߋ���`Eo%�wE0/;�Bk���wC1;<>�R3*�+ލI��e��" k>O���AY�5�'�M�c� ̉���yv�_��a�'�ȓB��Z�[7f�)��{;������`+jXIk�����m5Fǌ��(��b����~���c[�v���G��w�k�� ��3ťK��[d��+?j�EMɋ���m�O��%� ;^�B]F��}F	�3�ր�>��_�|���M��'~a���Xy����G}��9�Od��}�{٬����H�K�1�CwY�C�)��t������V!������;T�a�k�]�p���#��DC�&�D�3��o�\VL~�˿����� &��
M��QU'�%t���u�9M��Қk�Qc[�������?�{,#�4������w6>ς�~�ϳgA���]g�;�%sB�!�w���������)��r�h�p�a���k��K��@Е�L���K�Ѽ�MB���T����h�"Uy�[�����%���N�$m:@���s�_k��Y�w/�R�}&�I�:2��9̛uAx=p[n����$�)��yƈ�#���: 9tDd�Xu��٦�:�'8�R��$��'�lt�O���12ᬻ�����q�<���C��z�:��	%�l��F,�1 ;�/.x|��`�&�/]�j�ll����Ʈ��؊��<6���GG��ӪQ���Zɫ�9�e����52������4�����'�I�B��|����g��Ħ�� �[�&7 z(J'��-.�aG��� �ē����|z�m^���cS���2�ӝ;Q����
W~ٴ���8����_1�D�*�-+�UA	�]l@Oԩ����Pw0iZﳭW���W�t�h0��K�6@v��� ]�����L�uX(n��Xx�)��~�劾��5��xyH���,�9!n�H*�uc B#�-�s`^=�8Rt��	o~P�X;W�%ﲰ��y')�e�B��p��!:lYs�̧ϗt����y���g2e�'#!���N�(��C*��?�z�t	��r@���Ǐ��/��⃿���E�H���c�߭��=x��xL��X@�O y!8s�; -P���uݎ,i�7��n�֣�LM f9����A�1~�J��R=h�ҋ�,x��bB�� u⹳f���àpq�tx.���ݰ�4^'�����܁pne\O:venQ|%!!���+Zo=��;�>Rev��GBn�쉃���p���|�`�'vg���i�;Ѝz�܂�T�m�r�?�L����=��#�BVԶ��@�x�p��n�ٽ���pcg�����ٵ9�w�˹-/7�z��6�v~6��XO6�@m[���^�]�l\$Y���f��-��seԱJwK�c��r����y;�5��رU�{�X���ԔN�T��X.=�gv�������C��W2�������ۛb��+��}��!��~���@���m�u�<��:�tT��p�0qC��㷗9����6�1v:|JÛ�Qʥ����uʈ߹v2�r�fp���#�$5=/=�
�,DFr�q���AA��c���<���S!�Er���$�ys��@����{6��6`����n����'�����Eғ�bI8���6PGt�:5t �H��)�_r&'�E�{q���0��B/b �'�k�(���qK�Q1��%���)��tx�}e�q�e>-�ݑ��YT��rl��f�ͽ����d�LC�Gjq�R���\2>q����uY��/cm��KZ�"c,�{ ������}Gǡ���
����쑵2���X*8����qy�?�M7�4��j���x�s�������em�M�)o�W�_s���h�JLN�@7w�@w<��668�N��q������+xP'��b!c�"�"�
Q\#{�Ÿ�؞��Wc*��N�+��m��A뗃:�� g�S���t���E�f��.Ui�r�⽏��V`���N(�����ۦdɑ�Kܫ�8	�#�<�w�r�z�[���?����u�B0F*ڭ�s�s��W�6,�1�f�93�|���=�����gvcs�����[681��@�����-�u�&&%�ea١ĳU�B0�b6��Ɗ�<�m�5IN ��O)�PP���g�$k�>"����I��D�����Z��x�ؕ0�*Zݯ�z��C��}���x���],�pE|���Ǿ
�S1�o� �e/J����?詓+�Owr`�����d��n!V �â� �y�|��TOq.��JwVJ%���u����5�k�I\�w��yə�l����M`b���8��B�Z��*������*,2��y+��Nc���=�&S	�z�K(�j�U��hLbFjH,�P"P�(:f���1(5��u#;`��J�V�6�*p�*���e�ʔ\�u��Lftrt@g ����D汳a`;L���Q��
�����)Y0}��IՉ#`��]&�{d^@=��<��v��J�Ɠa[�ǟ�O)�MC���i���#�Nnd��K�u�|v�P��4�}�]��xSyl�FKn��� �51�
��g55r~��J�Ց(�7�6I2@��fV�td������{_{�u5�mN�	K*��2y����Cm �)�[��g"�Nc�/�q�U�{��;����֘��m��~mխ���uӌj]��x�xiy����#m��u:&[�8�}�ͻ|���՝>��E�wR�ԉ�_ �xj�<UV�Æ�l贽}�U+�"nj��� A�3W�$h`�`-aRg�g���AV�#�9<0�]H<V�l��PK�y�=gZ}��غ���P��d|�	�)��aT�zCɝ�' ^L��GȽ�5���e��)B}�I���8p-�i�P@_�(�B{�v��,�c�Y��?�yl(���b��'����(�����>~�T�����[��̋�o���lN���p���,�	Q
3�U�J��WP�C�W$wEhJ 9\r}`�=��?��'�c���s����]t� �ft�C�P4������$���֬�l95Bx��YR`�3NyHe����￧ӳ3z��wt쏏?��_�N�=�0�U���g²���ﾧ7o^�����)�kDg�[
�<�`��VD�4o�VB�POo����ls4(�wɾ�^������tM1�oc,��ic�Y���m^���$-bւic�Ր��Z�K���~P܍ K/�y�D`�{�ѩ��bn�����w\�G.S��|���~T��k�%���� ׺x��~���]�����0L�/�a�7"��(LT�����Q���%���)�-n���uÈ����0���$���Y�E�4�'S�7�(n��0���(8�"!Y��E��t^]HyAzX�-�|��2�U������_����ir5,�w
����a	/Fm7땑S�O�^x=ܩ5��Wo߾�� dXx\3��`v6Y\�wO^�m�^c���L�;I�v�S����n���5v�
���LY�s3�!N�P��x"#�6��Fu��ظ�� 5<�@�v8vX�A^�6�"�ψ���Ob�`���F
������Pۂm�.�I��`�����wC������[�<���p��»�������:F7 ���+`�i��V�~��u��]��O5jd����}�y�5੕o���}��Х�U�5m�h֮_�>�k�x���i�FK��LI�%�J*�C��O2fZ��<��6ɵ���xI����߷y���[��Z{��aw�#EIA##k�6_R��ޙT�|]���׮ܖsC��0��::��A�.�q@-~�X{±E���g���[��}ߥ�>p�_���Z��K��Ո�jE�؁�Z�$��bY"�,\�ʊ-�_u��R+g����B�y�d��u�1p#:�Yrw{Ϻ>�ԃc�yn��9,��Pkh�|��Y($������ĺ$ݯP�Z�)���}zr*ٱ�+�4��M��� J�d͠]@�<B�^�zɶ�l>e�d�RѳY�0xyMаYob�'�:'u�.�}�dӖ����%�!ԟ=ITWsD���8�+#�"VxP-CtXr��R��'4;��t�ܓ>�sؐz�rJn#"�2h甊�7�Ύ<�z�K�p"���ݤv��9蚜uV�go����h�>Nþ���3D� ̃�d�ynY�.��]~������Ʀ(�`������t���˗t� ��������y��9���J2��#���;dK{�݅��ګ�86��`���:�\��	�J�\�����uB<a~��lu������6o���I=�\��}��X���~\Ɉ�°|
��c�;�v]���R�@�Ǜ�Qk`ӎ���0Y���d�ҝx�,�$��q������D?����۰`�Cë+
��9��x��Gp�TtA8\]_�@��K/�MyK\A:Gx�0:�����z}�Q��PFT���m�F�VV�r��
r6��W����t�By}���{Z֞�ۛkrMA�7w�,n�b����SW��.� w@�{�9�1���յWA(q���C�������B� �X�,�n����� Y��Z9]d7c?O�ǂ;6.-D���=���[��9�)a���n��ZH�1�1�[�8"d��8``�����M��:'�+%S����໖,��=ev������}�g�4pI��/;㋒��(2��,�Y��f3����s^��ȕ��qL�
#��a�M+:>mV!�X��8�9��Ӆux�h&�0'U�,3^�fl$h��Xh`�1�L{	���n�!Ï�֑����S�"9�d�&��-w���c�W���S{0��?A��F|��iZt��,g��]��B)u,D�[�M�*�<�� ���Mw�]����n���yRr��7��	2&}�X2Ӊa��U�~~��B(�;�2���-��=w?�=x��m��Te�)0�=��־�O�O�n�b� �j�;���E`�?��r8g)�cؕyKe2$F8Q$�Cš+>�'X`�Cpvև�H[���wxFltc�7Y6uܼ#�y�&�p�h���%�"U@�(��+#�5I�\H��������)�;�ѬK��^��d��	z(�m� �y����@g�|����h�0�X�G��8��j-���/x�Fk��Ĝ8�>)Xr����F-��\�/o��no�0^�xEX5���xX	W��F7,㰅bq8��tEp��*��1��l����L��`�s�Ք�C;�����%"x�\�W�EL6�>�(��p��(���8yݳ}@���<��y�>}���a0������]\\P�B���޼�xI7_������8?=��*��wB�����{���������F������Q ����D:�%[�d����?��|h}�?3��ˌ�{�v�*9�dz�7I�r�E>�3M	h��F��_:���lD���+ہV��`�C�)*�X�	��*�܍��+[
�Og�d?��-|99�7���Ç즗�JB�^�yC߽����=�Y5㰝�o��_��W� ��<T����R�*�7�"i�!�wj֒�Q2H�:�*%Q��ͽ�\!SW�h3� !��(��f�UIk/k8�����0�N@�5�EސnA�� $] v��@F]�� ��2<��B��������,��M"zϬ
Q��(	�!�����nr��]��ТmW��d�&�-[�ˉ�M�zVo�hYqȾ���MA�"s=�&�?:<`� ���E�O��4����9�1"]�y|L�3��)�[j�쵭h-�����xe(
�f�0B�S�}uWe�drX*_�J��V[�lX�7�.��R��Jq�f�Q��E����1�A�$��,Z_�D�����B�{��ֶ�p�z�� x%s:���d>��ʅ��Ty�"�-�ƻ/#��>�0�(��U��͘��e��%_��A9�uVu��qA������uJ��&�$?��w�2���;Oo���oC����V\��|=5n-4��p����F(�֩}�+O<?kr��������C)+�^���;�]/7쉖@!?��ّ�G�{��������|�����o���LY��+����̮�eB�!t�uM�d/�l3E 1S�����F*:t�:=�V���B+_�/���O]�קy�"zɸv��L����fS
: D���Y�}����Λ��[��˛H^�f2�AdE���W�g�|&����n�F���i !!�B$|}u-!W�Q���b�Sp�lֲIS&�i~��)�>�ab�"�ރ��أ��i��B���n���V����!��t0��e�׃z�ߑ�y^��y�������K���U��C��������;8y&�z�O�:b-�^%�2�Pڇ����:��x�M�c�I��c��N���p�$�$n�󏂿G����5�7�|u���h�ڵi"���K.�;�
�,4 �*��<��p�����/l���as1� l!���2��
W��ۂyl�}A���b�Z(ߐ�հ�X�C��Y���=a��ָ��;��3����[Z,���;�C������89<���M�[�\��6���7z�y��=}����Ѡ�@�!��/	�ꍌ=d5[�NAl�e[,��y���(���Z�`X$�h���+����Ң�t�vW����ݭ�]���/#�����E���L��EΚ��б�<9�j���H��g.������\��0u�7l����'��v߀�eB���z�.�0'?z���s]e1��(^�oxC����v�jqI��g�ݛ���ﾣ��gl����ӻ���_������w��Xɇ�����|���,f�©��6�E��rC�p��!Nw*$l��I�lU�aC*8��b��E!`N�4uzcn�v<8�Ʊ ��p�=��a�)ћJ	v��P׀,�cx�c���($k�&<w���*�{^L�,gKz(��Z3ћ@Pi�I�,L������S!a.��~�ИmF�S�x�w]p���B�K'q��@�yKyne��;C�Z9����C���"�

��@�WNxy����n�^y;��Fa�o�;	�+���DM~	`��;Kkyww�^7����HF(	S%H�>F�//NKx� ���Y��4Ԩ7�6'��H�8;�f�io�;2��5x��ףNL�][�������NRhcW�b#Vtf�f����?Fm>�p��pF��a���a��&���_���˶S) ��O�θ�o�	�lA��f2��~��w,j�;��oz��1��/�\��|��|\�� E�}��Aŧ�\�>.���H�}Z����ԻB�.)\qg���q�.� v*�7�`�US�����UK��[�z����Q��[a��x�J�W}��{��N?ؐ��j�$ѧ�B�0��z�x����g�)�8F�F�e�DS�)����䁣�:�u�]��d�cV�a��G��csy�#7������y�d%�!Q��L.}i�_�s�7�`@{��aU��#�N6.�^ �,Q=��*��	K:�DF���R�n���S��_��܉�qp�@���y�X��QkÒtܖ}�ykj�\$96`gS3���1�8B۩���M���o�#��rqvN��i�M:�����{a�i����p.��������`o��/\�4 +x�/»Acc�ɉ���u�Z<�I�7�hnl>��T�q���h(�$���ڰ�haT�����(�V �*�)�`q1�F���b�m9J'�Sik��J&2远*]9Q��W_�Ii.?�����_�4�� �-�R:b�)ُ���_L���
lF�K'n�"� |�~nj�p�B�SvV��<�.��0�g� j�[�_���5}>8d �O%�q�x��^\<�0B�	��lm��@�]�Ɵ_����gT
��%��x�Wy�%�\����֖\�T�(s�`��!jCr&w�Cm��{��)��5O��g�c4��M������b���lՃ�����·��@ٕ��S�q�$��*�#%K�ܮ(�
b
Z�g�{�E��0�Ae8�K�k�uΥ�+�F���߷m|� X������W�����]����hjBp�|������|�񣈩��F��0��͆w@��L?�eh>���3&ׂ<YV˅,~
 1���{uk-hB����ZN��t�@��ud�R�:fت�(�:2z���p�	���e��A��U�v*��|A�bʡ%�A�9E!�����B,�"0�e��O�N���Ȥ�g)�����=v�[�r\�3��r�[caWr_╁`�2bɢ=��1D��{�� ��w��(,N�P�=ct��T�E���K�!s� +7�������eSr�s�6L�'���� ��8�6�
�S�]���xޢ��"y��#$� ��F��1#'� ��N���	c���D�"��	 ����Z�6q�I��h&�v��݅`�=iQ�����|?s;� �JL-��j!/�f�H(%q��|���d��:�z�4p���ad��o��瓊�7v�B2x�I�n�m"�6v�� S:�������!	�/�\v#^��
�]�G�`UVT�p0)�<E�o��Q�c��0�7o��#B�����ĥ��a���6~ܶ�[�P�ј�&�ڤ�Iwi�����������*�)m�C�yl�Í�Y��]�1�:U�oU���8���o����w�s��>�m��;�4\�l��ѭm�v}R�{��*+����)�Y�Q���p6�?!3�&�3���k�{�I�vb��~�����5a�$��Ç������_�{���%'����� �B7��k�7�&1�'�9p�����fƲx��H��^<
ʐ�p�0W�������Նù���Odo��?\2�x+Q_�rBv�ٜyV������<����m����@�5�߬d3�7�4ǢP6�᧜}* V���Hʢ��p*P4�&z�3��S�%�ͷ�K�3����\l<���G�Z�o�R���観x�8X�^ښ5U�{&\~�]�g��J腡X>�/�Ͳ��JXR����Ar��P���x�ς����w�F�z�p�7�B*EA�X�X�Hۗy!5CdQX���� ����T޽���_9�0��Rq�2{�#/������ZI��,����	�:�)O��g��+n�S#!y�kx���I@��cV�or�\i��9~�Z8�����iԡ:�ҘZL�K��GV:l���|5� eB�:Hݿ�T]-EM4"?�Х�v��or#!{4�?u��s_������rC?̂�}Eo^����09���ӥ�O��³f>��0�/�U��W��Z�P�ĄጺCXӳ������2��/�o</
p�pt��E۪�Ó`H�������'��PA�	`g��]�!��t֋��srvJg����✎��Y8W�C=on�Yy��Άu�v���d�^��� XV5ֳ �$��L�	A��tV-��t'��~*��a<9x��2�[h,�U^�C26MX��05 (�����=r���c��ȫ����2i{�B�w�qX�׼�,��[��{�y�=,Mdv��,ة���uܡ�l��`W�.k{�\�yj.��a�a��S�.�P�MX���Ġ�8���ٖ4-���"t�2T���;A�B��n��F����N�v]���h��H �8C��	��:��ǐש?H\�h��j*͊�6��ؒ	k��K���vx�4bk�C��5azF�>��X�Է[����K]ݿ׫?V��b�;i�=�&W��>.�}jT�:E3�J�V�r1��
 {��%���I�!Zh��12U���pkԨt�H�Ѫ��2�
nW��{��n�y��ۡ����^3|��}���'�  ����-On�ԛLn̓f�c��;��ۢs�����a]�d�W��w��A�g�"�售�_~�'���KG�%٘��7�ݝ�!�����Cv.�.j�D�`�ץ��%Ӵ�l)5���Ʋ'�c���2�-�B�=��a v�q���g����.?|�p��R�G�x� �(g� L�� ��V,��6��CuC'���?���)�@���_���o�W��?p�#l�8Y��5�;�P��|��Ȅt~~�@	<7޿G�������./?�'4�d���Mvp7$��`6WAxc�`'%C�LN̹��d���Kϛ�ļ��1��bpk��핋��Q
�i�
W�PG��r�J��d�e<���{��0~�u�|�00N��ύQ���c�<�,6l[!\�7ֱ!�p7�yB�!��� HQI�w�p��b�8��*����C�k/y̔1����=ؚ���IU�d�����,��_*σ��Lq�#4۹���L&�>���)�Lٔ�t�D`��x�(s��5��a=�.�爑4��F��ȵ��Î�X�g�3K����Q��`���ݬŽ-6i���Ʈ=*�d8�h��%�
K��{Kut��\�ҥ�4��^ t�	di��	
���O���G��]=Hq�h=@Ȅ��01!D�B�A��Sz��5�x����!ޒ�F))�WB5�F����@B��a��G�ttr� ��W��0�;s�Q ۈgP� � �"�t�!}�����#v͔bCgG'tv|JǇ�t��3��ᝠpHV��$/��Z��`����eRD��F�d����k�e텽�-ى�<p�aR��pjnu)5��G�b�O�1�g��y��^;��E���`R���q�JUH<Lt.�6�;i]71e���¢�q\
HtPj���������d2i[�^�]P:�+�1�=�ik���ZvNx��HRfV����mY�e��u� iZMD;<8
�h�{[2J���{�\��Y�R��+�~���|J��RZ"�y�����-gp�&�X�T��Nn ����Φ���n�}p�cَ?�=��}�^�ӊ���3�c`n��o��Gzkn{�2XB>N{�) h���WA�#��UaNbw��y�'/�a>�r�H#}ڽԝ�������qa 	[�Y���o��	�!�{48���ݛM�3bO�'�q\��@�V�e���`|1�>���1D,��[��^�^��EDu�{x���G�h�k��绣�v�ݎ��tA�?店f ����姳a���g��Nn�ݥW�s�dR�Wk����p���s����=��c����4�p������BBr�rY��\�Έ�T�uW<�CK8�����˂�I����X� �X2̈́��{�" ���dOD��3��6��G�yV���pp�U����a$n,LL�e���P�e���C�����G䰱M)�����r������۷�������M�Xw7=��xsf�5#Ե  ��IDAT��!-aH���y�Sڕ3���w�M�*n�&��2�5t��e���VA��-k�l�I�/´���N҇C�Gl��ũɧ��n��:�ܞH����Rލ��dC��t�����I�@(d�Z�w�ٰlˊ5�Ŷ! �k�u�z�z����e\;�i�t	hq�E�&�۲f���J�=c�0BK��Y�d��\��x��N(!#�7Xm����S�@<戩W��uҍ�PlT�@@=�{XE��#�E�m����ȵ|�����K{.��k�6/�dgoȵ*G�wU_�����@�{�,����9R+���<�U���c(O��#[�]�����i�v�{��!m�B\M�xw",� v8�2���[�t��.//9$+,q��U�f�����cw-d�x�g/���`�L�b,��s�p,r�h?\JA��(��/W�����?��fS?
0l������$,��\v!��26�C�F��L��[������/���Yp���s��]���Y/7��MV(�}ɠS��E����Ӯ�/G��vě��Ɵ�e^6�o{�h�n^V����1n��xs=Pg(|�7Su�ǩTh�P �m����r�3����S`��kF�م�)��Y�G\J�r�;b�� �?��x��j)� ���<X�8n[|\�PP���r���"���s�1����a�v6��+B�����Ӏ�?4�����:�v^�LĞa����n�"^������G����d�Se��JI���y���Yǐ�h?�ױ���{�s��W�h-���y�"�} K�i��"�����3�.��m\�C��U�u؁��0�0 ��@(���\�/$��o���E����ٲ������>��R�j���|�-G���)���J-g}�D���7ޫ~����J�"��\v.�[�~�x�Ԯ����؇�(�5�`Ǫ�p_��փ�4p��*d64�voո�V����Ҥ#��#��~�D�u���f����H*��Wd��^9=�s��5��@A��%�a��dCC�g���oVS�uU���P����Fu֢WJ�ˡ4�da�����G��
¢x�
`�C-������7�2֋�b��I&&�(��hD7��W������9$}ZV�Ǒi��+��1/k<�5C���$��?��>����@�tO�5�ӊS[� ؀� �����gPɫ��g@,D#�7>�Х3�B����4�T��{�6�J
�^��zP7"�Ri^�����F6$��J��4d[����$z����Ijv$�w�k��\�e�}���B�6�-ocx�F+?U!�HB�2�ȟ_J"�F�$��/��:ũ�9�l��M�c�u�4Y��:�X��e�22�]h��bS�B�8��aU�`����q���xI�O��B$�.)�{\��r���m}]X�x*d`x�� ��U~'�x�����}��ǂ:�Jt�ׁkM_kE��ddw�_.w�U#�J�p��U~S������x���:\����y<�w�R-�=sZV�.z�%�<O���w�/�ǐ�cN�|ȃ_�e8��o��36Z��D&s)���ͭ�aB]<A?��#�t!�H������d����b!韃 ��?>>bω�^qʻw��чw���~ef����ó�����;��?���&�B�0ܿ���=�^��.��~���]:��c�����������^\���P���_߱�:�Y��z^ ��k�������E9p�%�K��ɍ�=wv�K"���bjyRN��1`�;�b�'���$">�����B��Jyw�d�S׃�7�.��d�(�C�*Q��"ʑo��J�r٥'{l5>&�Bb�!��I������Zql1�_�_8�v.�ᅅ��y�%��kP0l7I�S�$;]��!*��T��ЬP5^������=/ n8[�KxO ����ty�����R���SƁ8+z��Rt~��@Ol�j�V��24�Ua���qP��U!�@�ZȓK'��x?�ԥ[��y���-�	@Hn�_{�]���.�cp�_��~��m�����#��崔׾�u�f4�Y��R?���=�������<1�$�o�5��i�T7�
FB�J/%p2	mq0��S G��I²#�#;�b����m������6tz��ə1���ܵ;����,�� `U%��!*��O߂N���HE��(=���?ƭ^�k�x�[N���ӗ�ߵ�֬ӛ�K��	�\���\���%�R���d���΀N�cb����>�5����8͎	���)o�yL*O˛^�},�B%5o���gc����.�MK袐9��1�6J�5��d��W���R&+o!�Vw�Y�i�'�r�q����]���x��u,�R���ЯA~>��A���*B{Ĩ��2���(������>��o�o�7�y���IR?�>��������pvڔ͊9����߈���h7��<v���>;=㈁52�柆/��S@� #k��� ����ě��l%�h���h���N�G�7�r��9
6 �w~r���#�̩��(�T!c6���O,Tqc#���8ha^�R]`�Q8[k���ÃC{H��LV��<�5����)}�ds�S8����F-q�5�|���X�D�����0r�m�\?pm���@�J�$Raʙl˴q��9mB�<s�)�d�{4n��#��a���?M�~ݡ@]�NT���	{� 矮�W��6�DQy�!�K�GU�b@cGBnڠN�~�lp���	�1��҅]��9��������!s��X�d�,%����y�� H���4@�E0�1��A(��ҟ����ׯx���?~���3G\.�^d�4��w��@�/�����'���.��O>0�tzrJ�^��Z�����D�.X�!0�B����9��l�	�^^~���;/_�����>����M��2?	\)ُ������|���A�tG�n�9J-^dj	b/�aV14I���*1vR���;1�b�\j�km�Qc�cy,������X�p���o]gG������IU��sQ�Le�3"W�}��p�.���QH��R)|B��3�L����I�6B��E�S1��B̍��<�	�$�汓;x�Q/�b��Jл0.?\~`�Q >V���N¸
eC��826Χ;h�P4�ɭ�=�0�Մ��/Xo	�)8vN�?J��j#ٯ��r�QO����^qˢQ�&�<2
�7;k��};߸o��n#�Q��;���c�~͟���?�ި���{S��d��Q�F=�m���$�K��i#�U��rF���j��@e���Yy0��c:89�E�	J�,�*ri�GI���7Q%��j�e���b��VP���N9��u�ܣ��'%Y�Y��&]�ɦo��� e���.fe$��qE�g��=�B�o��h�n��)���y/!��]�v���L���d!Ӟ��M�����w�i8�h�豇���vjZ�g;g�����#z��YC���2΀���V&R�4 �^�GA?��z�hxv��8��W��E�=�Ɔ���0�7=����9g���YB�>�,�3��	��c��<8fВ��W���m�5�ǐ!���#� [L/4`���9o�]�:O�܍3�Y MBЏ�a.���U v��P�,D3#�֍�B�����t~6�]�ݍz��Ʀds����W�}	��3�8H��[�}O�n��
'LA�dk��g��;�z&�0��oj���$!�g*�R�-Dv���!�^���rt����^��Ō��E�a�i�ג�Q��jRŴ�&�s��"Qؓ@�D��2�R��8����[����NP�`M����� |��n���4狹/U�?��~�L�B�b��2�N5�� '�E�fɡ] ���iM��:�'a,>c[�+_�Lm��c�l�+�ʛ3��`��{�
7\E���:]��Ew�b{��=ᴽ��C��z&��c*p~�g�mG�S�Zd�[*�:����شYe��/탗[U�&-۷:�YGQ���6_��cv���`�6�ZotP�i�Sܦ�p���)�FL0P��Sif�:�M�ŀ2#w®��
���� �����	������t��}F�9���[6����[a1AC��9]2n=��F�D��vt�]����e.�c͂��I��*/;��!�7n1�>?���_��~�冚U�DɌ�tH<�H�}Є�A�Y��(�ia�u#�1材{��aPyxU7�V���fJ�ԍwD2�ZՎ�N`�y�X�ۏ���+\�Yf<�F@6�M���Rc�+]��3�P��5ߕ��B�(�L��k���&�M���"��VҺ:.��`���/�����d��k���J�M*
�8�9PLTG�DV�!��t�p��F2x5�
Gjt�*�)�-M�t���/.��)Tj��\96\�hz5�X����g��L�'�����x����wK�uyGւ;�O�vV�ǠW��E��==Vt����Rm%$�a��x���{�m��[�䋩���;G�N��Lx"#5Wn�n�$3�g'83j�8����x��f˰��Q��nk97v��]f_qܤ��`a[���x���|N)�@��`�����]���N�ç�`���}f�ĝ�L):��ҩ�<��t���K�p�6qZ�G
��޷�:����}���4TF>^�Ƈ�]��(n|.�i���ϋ�)��e올�����FN�)��Y��2d��&���@.Y'�HX�qtp|H˓%'�X�-�͠C[|��/�rk�98�x!<��Y�OӒ3�ֺO'�I���<���:�Sʯ"��S��2{)|$��w���=a#jƃ�A��wyz.�D�Z3v��=x9����3=���
����QU5YC*I��6/�F��We�(���pф�]���G���[�3���W ��x���(z'�,�-�q�H�g�/nb��yy�=������D1k�{x~�y=��pr%gI=?:�Ⅷ����|v��,���oi#W��D���on�:J�řbө�����2Mf������bE7�+�x�zy~A���iOd�U�+�_^�&d�i(�ek����<u\V�kK�������9%}�Ƴ�h38{�=�`�4�v?�G[ۘQ���s��\@��lK�����eUg�vY��	�u���q�z~�U�d|vb�r��r1)�L����P$�� X߫L:�ǎ	��	��Vn��[�z&��D����W�2���:��߈
�؎�}�(�L��v�w��u�Nv|"��0�^�� `np��Ŋ�i��Vx�h�{�(.�;@{!�8idA���F ��uM�y��wtw����i�;L^ ;���E����6S�C��/�:��$3/>���q��F/����I��I	�����p����7���5�;Uj6K�.1Q��$�.�p>��Ǽ\��I��c/���s�X��HL�v��7�d�f��m��e)�3r���b���|8��YY���|a�9��E��w;2#@��Խ4z}�'R�Y��{�y�a�d� ɤ���t�j3��(���%Y0L�M�JR��m�*�c��E^q������E�Q΅}��)��;�������Qp)��V7Z�h�*���pI vȑe�b!aw^���1'$�>n���p��x�16��{<�ط;�c���-��|�`�u�wl�u������Z^m!u�0t��m���?6΃!�W�Wnڈq��T�K�{V|iGS����l��N�՘4rS�lt�[��&��������W.��Kmߟ�٥�Yp�-��5p���\��-��N��܎M~5~��������F�q'�5-Y���v�c���
�Ń:#cG�{��އn�l�S��6%����*���D�vdZ��kO��k�͐R�	g�Y��܀��-�^e����?2c�U�.E�%Q���0�csix>��.��K��'A0hYP8����dI7�d^{&sX֨��4iC�(�Ӏ�B����a&&�]jNQ-�da9N��ٻ��!Yb%�8����$��k�LX9�Q�~��Z�n�A7F2���Wd�"&�x�V�W�|"�����=�ⲣ�>n���%_7)q�����)�f������������$��It�gϞѪٰ��/�e�>�gJjGݠ7%_����x�����ú�=M<�h�6���&�^���8�pqz&�U�WR���Z����yl�K߫�)��2�,ӣ�[�o��!�M��{<ag�� }l�yX���\����O����Q�o�c������%u��$��Σ4^�v)��B��ϫ}"�>MǁDx��R�K޴��,����j�c�7ˌ��)��t�?�do�KzoL����D��"ʤب8��@�QW���:�=���ի��$�U����=��M9����k�?�Gv>*���8z�#.b�28b���Z.����å>�J�'�j�5��8E�*x�4A����R�)������t���g�,<�0�-���*��Wtw{ˠ�g�Z	#?���s���̶ a�r�.�����SiL�x�2>a�BB��H�/�%��	�$���	���O���<l8�JK9�}������xͪ撠�C�,͟�݈�*� ����rf�	�!O�vL���+�2�f�a�r�M6'[P�L�ww\�O�
���h��z1Ӌ� �~��`�rNb�_��t��(�f���N x��Sv,$�S��<.� ��$�]��!/�'b�A�4�����o��/���;���������m��a�nmR��g���X	��CSr�k��vG��VMź��l�A4���ڵ��*G)��*بn�>�e �GV��ќ紁1U+���}����׏l������kAb��(3�g�}�U��u�Z��J�I�^f�Epf���!_o�wQ��3���$�����Ì�\Y�S�g��?~>�w�H�*uQˀ5X��2"��G;�&�d�݆���m J��m��H��;|��c���b�����Q���W��[��U��8�8q��^#�-���p������!��n�>�d��	pYD�TB@kZV�����d�A�F�jٰ��t�� eN<��p%K}������ԑ7kA<�\E�����ˌ�8KG��>V���g}3|[��7F�Ux��B��=�=>�d�`$jY#�=��T0��Z=4'xF�h�σ�?<������q��pY�;���_&C���`9'	�sX�ʙ��u��᥍��`-�${R	Qq���5͸z�����vC�5�D���82е��C�h��q�A��;��
�/v��-7k����`ױM5��^��="8�|󸷤"��x#ܛgw��jQ���M�Bm���*�t0.&$�1��!'�'܆xB7`u�j�\�fj�1��z�Aa���Јl���e���|)��j��C3	��q#�w[�.x�#+����0�rd���9d��=��.?�X~�+2���� ˃����+����S�;:�qtx�Y��Y�gRa���t�gg��x~���u$M�x�,��\&,@+��/��1�C������Z���Eu:e�1��V���%+J��Hȯ�{j ^`P��V=xֆz���׋6)����W�Ǯ��-2��P��o������I�&��Jond�z,�;;/&�2��,�R�g%ϛ��mE�.��J��Bĳ)�6WP�^�q�V��K�B����uU
p�b-\Q/�%.������?����4����4#Lp��#�#;H�+D���x�a�WC$}� K�X�crdp���Ҭ\���_HX���~��ն�O�����ح��7��w����Jaw|�,�6�}�o��O�;w���OY1��HΖcH��c�ִ����'���HZ�[�������٦�� ��ak;�x�@�y�4�N!NBl��	��z�,7a.Oj��������"�<�F5�IA�-�Υ
�Km��[nT��o��p%���I�v1�\��7;�@F�*|Zi�E��p#HO������&��1�ڎ#[�j�,T.�M�-�~a׾8���(���>���%�n5�ե�����*J5���0���8iF�}�pYx�>�=<��PZ�aAf���)|љU�Wu̘E>��UDs9{R;$Q�뗪�"Tԉ���������P�s]�<Oln�[NJ֭ �p�#/F4�j��k�-ېl�Z�&�I�2\�|(� �)�U��U*�I�;c,o<��G�S~�J�Up��p3��6VjmS�������~U�/�����У��lX��_��\�hl]��h�v�R;'���vv�s��	{,�FCߦѓȲomԣ��^� a V8�K9�̣�1��hأ�l�8��J�NjkW����n�!��a:
񸪊���e7b�1�6�+�3fs�@��dr��a~O%z�ճ�PBeo�����=R�F��7��@9l�YA��g4����$�sD�r��#�k=I�E�.>QωB��L�T�_}ıc6W��垠�n��UmɊmKb�hwzJ�-a��_u��v�����ʬ���=�\3E��c�c�BO���F/����Cڗן9���4L������+_:������U�Gt����g���K�HUn�� ؼ�xN��'L�~Xrj�/�>�͗kz�b�D���F�
٘<��h�,�l[���݂wi���;��ֵ��P��p���{!�o8��'�^�@��,�If&�J�״�����#s-���3.Ɵőڽ9P{��\[��������:�P-�����³�'�~�4*BzKo$vw�m���1�^)��k,Ԧ�����R�v-+<�NNN9�:�oSK��R3XX��23��*KM�8 �Ɣ��0WGi��ңm�Y�<>:����d���O����r�W�>)�Q�l��c'�.�T�;f4�|�����o���%~���k� �1$̐�d��-FTﲝ@���=+�u*����M�$7��M鞓d���8ʴ,�>��[є��l�8z�kU܆�d��f'��2�_��&(�̽ݖ7�f�f�[�N{~�k�J_>���A�yn��]I����J�����鉇m^�1"#g݊!�j��յ�{�ߴ�	��9Ha����8�y��j-3n]����A8����}����v�]�"`j+�G����h:]~o�z[;5u�q����:���-�������"�=���5Z��)��-ۊ����F�ș�Y�7�"��zMA5��[p���L����)+?�E6ɜx�0o��dY�\��+pQr���!Ȓ��4���#���e%�!�+/!��C*Wei.E��^�>hҠ������ĎƸ��.��V ޫ��ȝ�.b.���V��bpj���f��.��e=�K�'�2i��ށ7c*n��6%M�1�	y��C��ߡ���(x�#@������4���6�i���>����d'�蓼#�}h���� �c��e�uD��/_�p�����.�ba�\U1����'����ǗF譍�d@3��U�-���/��ƴ!�����OL�њ�	��.0�\������ѕ٤���f�B���m㮳J���ߐ�&��la�%eam�Y���nU��!5q��v�ݫ؁�/���x߽��3��x"�~�GT������k&^�b~�I«�����>~���s�a���_��������i2^�3+�txv@ϞћWo<���aA���dʤ�0�q�u��'����%�^]�Y�j!��ų!����\x���NG�9ntSn�wqY-����t6q�4��z��T�XW+���Kx������J�]0�=��Fw=�,n���<\�Y��^][��@���%�3]u�`uS����y�U�ݓs�ݷ���)C��E{�)��!�p2`G2��Q�����0g�&��N�m�����kx�̓B���www��b�C���a�:�VC9���b�uZ
�������`T#����d�|&^;�U[�|�1rc_V�Y\��Y���J�R��Ӗ�䇕���I���0�]Rg=m����}ˎ5x�5�C���k�{�ӈ7SK�n����_~>4�h?'�%/1��)^J��I!��@9i�u��:W3i�'�(g��)M0�+�%��+$��\jB��ث���	>��x[����vE�x����Ks�Z-�3b��[�	�4���v���X���C�\��.��;��-��(kȑ�n��;<�ƟK�P�j���{>�z_��d��!?Ǽk3��c�3��^`öpJV��{��+�n���q>�|���k�]�ޡc��P��<%�&�w��4�ր��lZ��i"��9��N^7�|^���	T��3�Ch�T������={�B�FݧJL���K��Sx5 [�4x0����y#�=m2�nˀ�φ�|�t��g��?�Ȅ�]~�D_����e���3�Q�#3�iؓg^l�l��z����9QT���P�(��v����"��56�gF5��D���o���.#$�Y����V:���zq6���+޼rI���N�ez��v
�M�CF�f���נPO�Dw���(�8ai��WH�hK���&Q�������H�rM+����%{)h��\�N�����}�#2�Kƴ`�1�l���z��#ˉ	2�a`c���@9x�Gj�Bӭ[�4 ��Ё'�A�3��:���.B�5�Y�õ�awB��bV┽R�J��}�ڋ�MЧ@�<\��֩!�6��i����:��'���2)�Ĭoa�q��I��<��*ry�� ����#>I�m��?�ȅlZ�em�`AxM�$�t���AL�3��,�t��W_�����O��a-�����~{��q(��W�^s��O?����Y����g�����|�?��:������:�w<��\�q�SaQ����b�.� G;:>���:	?a��hq����:;���j��OBY��
�D�Bو�<=9��*�`�o^�8E%���&dx�
�O�����4 rT�YLj��r��c�@9�(���=��b�q��z�������������.��)�`q|�;Mq�䅰��o��>��j&�^o�ݻ���6��.�hrJj�4� ���( ����]4��U1���l�B|��zE�]��|�߃w:��>Y6��@�<Y���̽�$Yr&�/"3KW���0���	όώ �;�3-K��x|���YU�30f�+E�']|���!�ΣW�1UhH��WV��DO��o�==�4�f�����PH���D��t�9��_O|g_�/��M�f�PNzz����Bc�L�Iu�W��X������Cp�Ü?���
��+�0Y�\�Yp����=����9v$/G���t7}�b���ff>X?R��RUf����O�85v��Z߳���XL�#�{ ��
V�����{�FʩO���#J�>��m׃TDh�i�U5x���g��j@�I�N��H�x;��2hel���m��|Uz)�;�ʗ��(�C�A�{�s�d����L���܈s�O˜_�������A-��L�Yàم�I���n=�iy�j^�T+A�bk�� ��~���	r�P�Q���"�y������r�H6�k8�2睔|/35`��	�Հ��r���ye���j�	Kl.tz��λ7�Z׻wo�����'s��?}�H7�o��Ǐ�^B*ym=���t�&?���k�H́2�+��enŃG�.�@��sƠ�[�~��˳/�9�������_�S���ןi�kr�,y�?$y6Ldo� �Ы豃��
���r"%U����3Ԗ��~�:�H4}|vPh;�g��|}M�?~��!�$v�|�^=VƋ�C38�S�,˼3��$���iqrd�0܌r�����K�_���-(�K��O�U�t��T�:ݾ���ѡ	��W.�DYD�^mG��Y�Q��I,���2ef�3����=R�c'�A�e�'���D��Q�<ԸG�?�R���=5 R�N�j]�u��U�%��x_6��+�����/���M��+A���!T�9$�����{��,20���ӟ�;�￧����c`�rU����3[�$㻫��\�6@���@$*���9~ qxM9�D�1���r���/���2�{���}W��1�G'� ��殴CB��[N9H��ySv�Z�j�bl�&�``s<)%B��,�ڼQb����T��x�X!Ύ����bm�:�)WwK mV=g�Ap6�ur$�i�ZF�۪P�e��p,��:.�.|��Ɖ�\s��������_>0�PG�)��b��2dI�q-��M��?�ïRb���ma��p�/{��1�4�㲦_�z��f/��\�/��3��4���!Qx�)�+��sK��!5������1V�-'��}��б�ÿ����E)~��wx��,O��|���#��1�M�k&Z��=��wx��)�_5=U����F��Sm���C~紆�EM�Z�Ov�66T�$?@?Ӑ~�Q?� _�[]4��ju"�H&�oV1���3��D�Pn!�"�%Ձ�.P75��W�bW��3p4�cΛ;zcM}�ҍ7Z����Z�tՐ���9|�h�x�f|4ޓ����0���Y���?���+�AG���|����xL�w�6�#㍞�}���)���[����z�q3{��i\��u�� O�wMd�N��2-o:�5x�5<���(�#��k�z"�?I��ك^�?~�|�����D��B�}���X�sr]����2[���H(����rqqΠ~�"��!T@ć�������2�s����	+�H
�aO�yg̴��u{�W@�~�tH�}�T�E6�^t=��l{q�$Յ���h�_�����r�0�<v��������-m�����#<���>U/#\b�;H����>� ��X4l�rsM��O�?�I�tH�_Xj�I���s��&��Q�6�n��P3����JEǮ�f�9Y���9W<�._Ο3�� ޗ�"+���"�n�mػ(뚳��9y�J�0I��)��@� ׍:�b%��˹3���sXj:�U9��/��ؠ�P�;�7r'E�����%��=��)�(e�*��b�˧��g�1��N
�J�7t��#c���O<�1O����G����I�3��. �̠���~�!�=��<��`�����Ǟ�GG���q<o�Ѿ��w�OG&/aL � >6i��;M*	�(���)��z��N/�������a~���C����-��=6�O���.���UـG�Y !?��`����Kz��������0���\�{|���5ǫW������˗WL�@}��w�Y� > q^� t�`�3���7���v���Ï���߾c�&q�f�,N��d�q: $*C�$k����͠0�
�ض�S��8`�4#'��5��̃�1�Lyz>���b��������*bU�F�N���L<��P�Z\a�"�lT�3%��lkS�����	�Ґ\���38�֮�\i�T�z���G�FN�u�������+X`�~�*�i����v�k#7rC}��;���'v�?�����?��>��b [�)?��򬫲�wb����$́�;���hR����8��g��r
��T�V���"�GT�$R�![��)�:�����a��g�}� �g�1�rx�(;&���C׺�g�O�7����8�����m��"x���^K{���'
����3j
W``6o��A�ƾ
΍or��"Svͅ3}~�=�'�y�z@aI������͎���;���w�R�l]N���<�Uぬ�Eжu"Ģ��L�����@�(7����ȡ	2u� 2�,�l/�_#x�D��%���b���>q�X2R�u��T���������g�Y8�`�$�u�r(���G�%�L���N�U���*N�<���l�l�r�.	>&�v�V����E�o�
�J��A�����#Z1Z�@E&�����������f_C�3�7��e�G�}�n�9�O���}���I��9h���	=sr�$7��'(o�Og���,/u���o� ^���e:��~4�4a���)�W���bmӰ�F��Sǉ�A�$��*�
� r.Z�xa ���2i���Qux�u{�}Ԓ'x��:�\���n��I�{R��r���͒Å8io�0�9'aF���UJ��y� F�����p0U�$ �u�6i�$�����*�>ХPY��X��0�]`| � �RRO(����%�	r�5��В'�47�ν^DV��f��![ivգ��W���䌚Ҿ�=��ʮ����{x���>��зޮٸ��"8�!�I��گ�h�ve����$Y2{�#���60�`mk�Iz�� �F����$�\Ջ�br��ZyM���҄0ɬω��s]e��x5�|DO|�d��q]΁~}�+���@�þ<�n�m��d9]�ˁ�E]�u�@��\�f����>fv��]t�^*v5шP&�!hr�/��1��8?����ҍz��.�E���&eqI�q�$���1+�/�tr~�I�N�N�8"y՗��������ϟ�CL	nz>}�����wz��%/�'�6uy�@6%\8~Y�O?�D�������^�]�Ӌ7��>&��)�X:���Boi���[G�I��q�9.i�f�M�I�P��<���A���jJ��j
�X^.���ɑ�Z��c쫒îIͧ%畔��Ē��5�¹b�#�ڌ�Lg������c�s�w���ށ�8��Uĕe:r%$�����J��-�W�t!g�S����q�V��³��@ε�<�.�yh�Y��Ev��pE��A\�bq��:�^�����~��{�@$���[� �(��?����������>���t���LQܳE80���(3,�� !}�Xf����/"ѧ���(�|�!(3���MR��.I�
�ri��>nSz�i���N:tn���"��{??�!m������ʫ�D�����z��v��:&�H�_w�D���E0��0��O^���Ja�g�T��=#=�{��$��U��~U0��n�`5r�q���s~Qج���Fտc� �3����.Z$�{��!^���j��Q$��f��Z�G��)Q�Kf2R��{�6J��M/��侮�<�r�xB�������OA|}`1�TiK��+�E���>i�Y) �w�/&��������͍59J�Y*>%	ݳjFNE��b}\,���v����#���e��c�;� ����.)K�2&!	x�x�z�F|c�3��Ɔ�I�G|u�մ��}��1�CA�H�>�z�]�r�No^��2��ˇY�=@�qٳ?����+qU+�/����c#b����32wi��I���@.6���E;�����G���y��i�Bx��s�k�M�v���a�t<ֻ5-7��H�V�<�qS�}�^��j� D��؀���;������� �{����CM�8�5 `˩e���W�[+T�fU��4
�:�g��N0��Ҡ�;�/r伟�L������^���+:C'z��9�J"��q�Jޡ��%m5L����Z�v �Y�qd`�|�d��5{�5�ϧ*��>�Þ��� PA�<�<����9�G��P
cɺ���:��`�]q.X�25}@5n����!�d |���H�v�k�u�Q��YB��!���F�܇p���tiϛ��G����f��8�SY�2n���T��G7:��b�o���1�~J4Of���qPg�A��|̎Ȳ�'�bb�]����=��"~�0(������ٷHv��'HM󰺧���g���{� |�իW\��H6�ӟ~�?�ǟ�?��g�x� ��k�:������L\(�������#gg�J���+��Ҍ�,g��%�����|d�߬V�
1�^F�&����U�t�>�m���Ԙ�Z]�<g�V9f����
US��?��pXR��ƽ�p�� ��r��7����!��g�Z��%]/z��Ha2�1�_�չ�Wc
�P	�%�ïp9�c�m}��Z-��f���H�삢>��Ƚ�^��.�}'I�n��$�<y޾{K�}�=������?�G�/ ��wo���ׯi]�����|�����MYO�t{sC =uO���p�:��vp����=�g<uDA�	�!z3%����F;�uެ8�0���k����Ƒ��T�;�y����y_Re�æ����{����S�c�����8�g����i��=u!蹏z�ᳪ��ѥ;q<z���0� K�N�x��Dÿ�]JnLf�TppG�/��k�{���K1�oLcg�/p! �	�E���s!��V�1Q�օ[�{Qj=�μN'�U�=� ~<���[�����ѿ���F��6\���<u�֝b�Z�٨��c��z��ZI2n�}W۠ ��s�!��r�7v{PU2�g��{��Y\���:չ��Ys�C}��J;M	IR�U��>��)�&��Q��C�?p��%�,Q���[�-Ԋ�%���t,���=6<�j���`�t��͇�T����!.�u����n1zI�ιp�N��h�������-q�D=#�K��CAY5/��m@�&ލM�E���d�y�R��`T�����\݈q�c��<��c���=&��e��Bb��l��&;�0GxdL�a\}2t�� H��0�]oV�v3N�Am����~� �wb�� ԣ�x�q$QF��w�Fp�.T���z��*gI�"�5��Ҧ�&��'�x!wj���Qʆ��ל�������'|X>W�/en���)�K�����ӏ�&��+<RXX|Ѿ��-da荓�!�I颎���i�@;(�?ڨ��8 gk�� (��y�3�o^��+�����KP�6&���0��v�w��#�@���V#�!Ne��E�򏿼gͶf�u#hi��H�n>� �^����+T�Z�?�/�����J0*n�j o���[.���]>�U#Pc@�I�@4����J�c��C����n�+FwqާO�����vk.?7D���,[TrM<� B*Ia�Բ�kB�<v��a�L�_7�(\*;ы&�z��N��9�N<g�\_�Y��xV���m�[�Y��
���Ӧ����g��X{�#�s!ǘ���02�	T�V͒۞[�#���-|��65��1Ђ��咭!p�o/�^���G��������=�}���-����^ n�m������c�����? Pᙜׇ�>���3`�.p�\�oI�P���ё!��
g|^��<m��r�G������F>��r��ψU�M�?�;�<w����zb��Ӓ���ߔ:��(]�f�׸b�,Nv�I�kMa�uo�?)<�W6�,�kR�������S������uk��1�d>'S�SX��*x�[r�\wHԤ��x=��i�y�ڞ�9$K�y�sO[
��8xPPl�)���;�塯��ۧ�+^`�W�n�lC �ɐ�%�C�w�$�T^�c/�|�"�	[fu���~N?����b_�+�sN6��I�/�j���9���G�a��ڱғmb���`��f$z؊����6Tz��5q��?�� 6��[�=|0 _Z�u�,�Hl�Ml=zX`<��W��^@ܙ����'�/�r^���¸�B��h��cC����*���Xj>I��~z������R�0 [�>�^���U!g��˾�"����R_e'M��۹��6+�Ƹ��W[Z��L8��#Me `�z�d�E�ٲ�ֱ�� ��G9!m}��|߀k�5b��e@t~�����w"k�Lm�~#�͖C�,�l��H�LXJU���T����l�w�m��~យ�=�������m �:N���;�y����l�ԧ����g̩�j�u�H�ʣ�'�ϣ�^*M�`��ţ`��PZ~v;���lG��fT��#U�}H�~F3�q2�t[��9�58�
F�۲�R��%�=
E���N6�b!I��, Y�XI�&�r�y'J*p�&B�9$	��z���N��n��m��'��ᖸ���k����'h�R%W�;�b���x�o�z�f���YA8N���	�ן�l�������peH�,3���c�Au틕�(�ʌ�� ��:ݩ��^�K;��p�5���y�g�?kl�0&d���s�0�������%���@�ʝ�7��b��d�F��X_�y��k�l�*U���(@ͧ���^��\c���k����%)�h�%�ʐ��Ջ����[Nz�l<�	�����k	�������J����`���R�I�vb��-wk���aÁ�;l%�j �7:rv7��W���'��L |��iz�8��3���4���3д(_��8C�"��;�9)�s�@���t����o1�����w{��ęÑ�ё���'W��.��k⺈�xVűT�:�ڍ�O�e�������Y���v�
���S�B��?z���UkēP���6J���\�3�V�Sx�Uy�ව
���z��.4����F�{M��'2���ßё'���5�G_z��ʕ�0|��^�>(s�*�����&�QɎ=`Lꘋ�"�����쉨�J}��*����4��d�������dL�Mu8(�1� H�ַ)��߮��n��Uů&��_3:��y��9�&O����Gw��>Jİ��Ts;Q��J]ll�����p�t^�Zf��*BR׹�:�p�P'�L�F��EZx���={�y���[#�Q�}�9G��{6�>�֭9Y��%�Ұ��0Y������/_1=���q����I�۝&�����c���C�jb���) ��CC���
�͟��q9x~�z��8��1�_���K�7�u���Z���Wn��i�*��h����/�!O����7�����x�������e �ۆHx�h���h�ο�ou���x��^�-@�3���x~D�e��Od���G�7b���1�tT<���Z�K�%r#�x-���d�E��P���������VA>z&�`�@��v��ƿ�����z���H�x�<٘��7S�����$r�T>z%�4�>�����A����9��$ƒ�g;��@�X֝�B�v����a��5��7��Z��{!L� ��|�1X,g"��^L��[uzE���
B� ���[��\�y�PM�U�:Fӱ�����m�\@� î��w�g� �TϨ։�uc�����q�=s�	~�d�<oAظ�0��{;�2�%�5]W�!*#i�0b�,��+!��x�
�r�0�-ǜo=k�Pڭ�����yU���IU�0p��P���_�+�T���q�4B4z�����<9���5X{ Go�����5�\@�P�y�;��-�V��&���8"-�PX嫡 $�%<pH�o+�n�$S���K�_Ǎ�y���N=+�ɑ�tH)Ww=w�)��K�g����2�횲��4|����G��*>Ѐ�8l{9��������S��nV+
Z���@ש�2�a��+cI������2H���7Z��,��|9M��$�=�YB�p�f����B
^܋�O*�J�	Sf��Ϣ�n<.[��RN?�Q�6�m��+�1OPI�x��h�������^���['U��1O�I4O�g	��r�bH�(�
�v��ԣ*xK?��k�7�;����M�X�^Ri�pz������IUnvr蓯�^��A5NrU>&A���+���Y�vwDߟ�Oz�ϚS���{���}�2\�j�j\s%vd�3���1�f��T22��e��$ᑿ���
˽챮�?�,9�1<,�k�Ś�r�b9W��+�Y�ro i���W���H�	�`'F�r0��q���,n6�g��6��xl��"M]�����فr��*G*���)g���R�� �O���8vrz�UY����"ߺ��f�����f EA�Ɠ.����U?�u�L�wox��<"�6�}/9��Þ]e��^�@||*9K;�bȵ"`�ɚ���Y�ܯo;��@>˫���ȶ�Qw�6�[���E�H>�.�{�G���ǯE3LG������T�$�Y�HӁ��S���g {�W���7����a�υ�2���ő*A�zS��-_��W�M&�}�$O٭S�a��b�T/9h�v������gIKYK���� ���0J��f.�W�IE%��W��4�Bɲ��Q�A!7Ma.�b���Z*zv���d�;�����Q��F�2;ZmG�5]��N�[`����5�ʳ�l|x�`/�Y fٓ��׸���(�������#�c�A���5x0��7gf���qg��;W,$��$�ˡX*��4Ok���ڹ����t�Z!p,���?��AN��0�ׯ�p�7�8��=�|�D7��\��_�s�R�յPCgY�۬$����h>�X��y�4�e(���A�p���ԧ
������݇O�����
��Daؗη\*M��+������ĪD��[��uD���玕�g�;tqxUP��t��c|����Il��a��CJ�`���R��sGH���ޟ��S�,c�b[D;�X;�����г�=�O�I�T��s�DG���
��
]�%�cA_��nU�<A[N2��
�*����H���U�Ԣ�%�Ѐ�']v�����y�u�G���p���4�p�x�\�$c�/SDfi�z���=�^fR&W@�����=��b��b�^8&
H�^�*��Y[��R�c���a~����wu�O�y���⢇�@�k�i���d�K�
��a�D���.�q�Qt=V_�����Te�|š��ik�؎xH�tisJSm��:�L9Ջ؁���������h�|��������k����<,��kk�S���n���2'�-�>��C9�è�OR����{�i�	`����{���/�p*x2[~�j45u�t�E[�_���~�^�|A�?b�yb:�ZE�,m�0�Vi��m_���#y���{��wiD���"D	@~��8>>�*����������|�4���1��8�?h>��o��H�"s�f�- ���e- ܺ��##J�kn6&cLgHJ�g�J��Q.vst�z����� 4��-^�3���^\�wo��~��fk�*G�<#�<�J���{R�w�7o��✓H��ٿ�G���k(K�g"C��> ���A?�;�l)4\�6��F��Å�'�TE�o8�i!��%[Y�O帨��E����j�2���ѵgN���``g��;�X��ʽi�}�A޳�}-�ו���!/��$Y����&�S�t���F��q]�xua��[$��^<�y�$�>2���c�-i�;٘GD�$Qd�I���y��ik(�;����e��Z��G�*����YÄ���r�G;��$]���fh����Ҫ%C,ڬ\Ì���a�n ��ZH~�x�4�m
�y%��X[,�y�4��a�tWu���T�H�+*��W�/�(���K'oYX��_f�=��2Qw%��[e�֒�]��f���D��o�cy�7��֞̉��l�������� 朕���9�����;��cy�S���{��LyY����
A		�����B6�������#�ȑ���۸�����`s�����ޛJ���Ƀ�j\��������,kSe�7P����Yy�ZH�L�_Y?���3�=7�A��x�&�ȼ�w��KN�\%;���F7�r�����w�'�.W��DLR�����c?=O�4�ؼۑMs;�Ø�Rbk��� Sdќ��>)�)c=S�P�Z��`>�J��nWs��cp�)�!�����+�0]����eg8��V�wR�m|}���O���{}I���H��E׺'�מ��<�G��8e{lF$�H�=�H�y�r�p"��4�Q�Ka,�>T�ڷ�f#���~�`{[�������5�4�<qkڥi��(8��aH�H�9R�bR�`!{�,�A��4���1Z�ז�Ь��-���8쑠���K��O�Ť�O���[�d�y-ʼ�0Oϳ��a��#��Y���������0$.!���ͧ/�2��E��EYS���gtVe�7�~n���-�T2d���h[�6�작������)���{�9���'�����g�٘�#�&�����������6[�c}�	Oq���@�T�����p?d˅V�g�vFqͰ��b�������G��z���/��߫�]n�xGq"�ű o
���}Ϟ��W/����Y#9 Q�@S־XT��^�N-q��=�5��V�m+ ^��/���m�,�n��J64��9��\�C� �̀�Kùz N�J��r�:<�Q��|훇�D5T��*������1a�i4MN9�!>M]��!��./�����$�I��9���3�x���2���`�o�-�j��1���������8vX�1�%�����j���V/�zIu#uP!q��1�00Cc��MI��!��ɦ9+��w�����˅J�[�����m}Lt��uxa�����-OƜ�ޘҤ�4[<r�G���9lrc��'%���R
�v��u�|�k/����IQ��:�XҹW�K��C���4��N�-W�/w�^��Pe��/�%�Z����� 8GM���bW,����pKQ�wS���4�Zu����xU<\��n:�J��Bժ�s��q�v6����g���c���c;��8+K��o�s���S�l���^��s�m\f<�$�X#+�=u��� �VK�* ��3(������V
R�.s7s/ -G\��J��?\���Ao�\b<bNY�Y�"�O/́��=u ���5���/>��f}� ����Y�cv(lŃ��.mY�clTtҰ�� �G�|���3�4^�����db�a�r)	硁�Q�O}d�\9�/Nʩ����-��q�a�r���#%>��� ���~�n���!K)4{��J.Q�0�n��e�	���l}�=��N+�@ �H��v���F���9r	%ɃQKs�x͏��Rrq!
�f�+Z?,����Șe����K�Ya+tm�|`Z�piR%,�ǒ�B���^A�p�xZ�X��X��aH6V�V�F����Y��)�+]�F'��Bs���Ǫ5Y=ul��0��B�&-2ѩ�`iϢ�Q�z��D~�Zm�Dٱ&���-+�M�^m���X{�2�	C������3�/��{4n|m"�4�p}1�H���&]�&vJ�A�x�g�xM���C���:(r��M������p1���u��tFǇ�f��_�StU��!ϒwQ���#��.��<\�EU�$�>�r^gk7K�t਌��<9]`�b�HC�9mR$�����No���@��,؛yѐ+�2Ǫې�/����-��{�(� �^/_�� ��K\��jA�l!�S,��m��*�t5w
0ll X�zB�OY>�3�9Dc���!�ZCæq��,%A���*�JI�mi�y�X2a�N�5�^&�e
4���Ї,j s�9D�����
�;^����K�>AE�/����g���������W��o�O�?�����ט�{*�}k��a�3��h�^��zJi
���?����8�j�S=e�4a�Ϛ�Nu�pA�q�;�P�=9;�1G� [G0F d�R��MOw 3� t�,�̒R�r�)�vR@mৎ,^JR�+̖�Q�Cu5z5Q f���B��^m��9���;�Bʭic�o	�}��Fe2G���x�D(�5�|�(nL�}����Ifg���M53��BJ�:_���e2�;������x�`��0�3n�c�qK��"���6����~���pBO~�����2�GMfWF"
<õ`}�m���
4�p��+�����K�Z��-�X����" p�JQ` Y-5�(l�����N���X��2)����PU���@�T����R�����6�r�xݸG	������
�@�!	˫��L�FR�N��!'S�?��>Gy�6S�1�l�א,Έ��!ga�bK^��sq�M�p!8���b�k�kY�"0K�5�-��Ĩ�E��b��@
�j��M���8�e�7��ʖ��Dx���1-��Z	/�in��IyS�R���n�u��g�O�~�獻`|%^|���$v +�Y�o,��^��W�6�zo���#)k��.,����pp��t��@!�q��8�f�oQ�&B�S�P-}ʒY�=&��zF૗��W�su�ƴ$tl�76�T���d� *Y{+-� _����v����N�:k
�b�#��� H�CB�v�����yupWNh�� �d-{���I��n]�U��?���@mLE3oP�P���E��l\q��A�����N�lB�Y�e����h�[���'rpu�:��Mx�������0r��Ve�O����l�[:�4TC��cP�\����e��
�OI��<7D���itV�d��J%��N|�)8�T��*�!̩��FQVΝ�E�{�%��Zo)�J��e8���vG!׺�E)8�c��Vpm��#�0�������z���W������3�ٓ��vik��v-����v/4�Ϝ�*R�ʵu��3ZxC!#���	r�ٯI�oCP���t0U`GA��k۽%���Pߛ�Pi*�Z �ώ���B�tI��z̈؛��&|v��|V=�C{䴚�RJx�a-�00�%�����,xT�>Kf���({�T�!�v��#�>��2~���{I�!y�<�8�_��7���[�޾��h'tx����ϒ_�Ñּe��u?|����+���}���O���3����W��SI������9�ѣ����ٍ�l���aT��G�2}%��;+�r�[ <��Id	#�H�'i7�֧��~0O2urZ&ʓ��+�Ӂ,�Xg���G� �	�9�Ok��O�}8\9؞���T�k���8�z����`#��������c'�I?��(H��!��Y������� ����0V��1	A�]]�=�\��.���kj���4���Ss�l]-'A���g`�V���x�S����zј'�M�J�{�j!�v���������.���|98E�� 1M�������R���P��Y6�y�(�7V{Z8�ƌ����	��B��uU��\r^����k�����^�	e\�e�t�V@�Q�Mt��w���"����%��������k���]�a{(έ��#�'��ȱ�M�Rm;�ad))jK�\vm�V�|�+� �'�q���~�ale�[k��	)p��hJfe���֬�Na���č��{�]��{C=wп1͚f���x���e!8W���	��¯2w��n��
�Ivsk�5(I�7��M�&�9�Nz��?g_�������7;F�o�1"��(�VjXt���yrE�nٕMrcm��
�{��!�# �ܹ�]�$��b���Wʺܮvt��V��ټ��ɒs ��Eni����N��*�.�T%�T����xu5L��~#	A�r�sᖝǏ� iO8��_!:Ei �B��[e�L�5���@jx=`���R�'iRjl��[$:�H>ʺ|�po�<Q��N�]�{'pY=jm��g�`��+DQ�λ����[[5��%5n�Ӵ�"7�P?��5-^��Η����<<�+וs�M��)����������*�Gb�@(��:5.�����=�*RkD���$ގ}��e�s���ܖW��۔q���"o�}�N\���o�V�|X�>?geyT$��F��A"�b������UV	�l�x4˻:���yQ��*��oQd���3�ؐ0<�q�"3Lk����ݻ	�N��	�*�i�9` �w��5��rDҐ���M9�V�Sں�͕5W�W��T�ᒁ��#9/�TwPp
��
mga9�}�������./.�y��U�M_pN&��勗�����섁��P��%}����|��ٕuu}C�~ˠ����&r0�h��ZY��?��qX���>|�@3x�=�\9*.�;�X˙�eY^���c�*�<����{[�aPcO}����HA3t�3����4hOo�~� ƸQ%���#�N.�a����"*���:�`�oyD�����'���_�<&_���{.4M��1�<ՂG������͊�Q�����1�=��&�iԮ��*w�fJ0zᎄ��n��5���'4����������^B TDP���j"J)�-��jrI���;B�h��_���>Ԏ0�a:�B��y�)C����1�B�30G�[3�ı�<Ҟ�w_�T�s�$O��mE�j���ս��hX^��A'�u�&=[;���v_����)D�O�2�j���A6~ L�>�%ɭ����>�l�p�ղ0�{	ź��k�k��W�rW�:��&�4��1W�Y�Mpr������\���k��{�v
S�㯟qGo�^��j.f��H��C		^	#u�����f�yQ�ڄ�F���޺�s3MW��p�+�NU�}�Zf\F.�//qAW�6��Xzr�����0�򾆰@1a!9��q'����J*�M��&o԰�S��ڐ�L�9�^��y��<��i��Pd�������y�a���ꌖ8������u�9�'q�1*px�-$�(pT��E����k�$�/�XoV�?�`�nؠŜs(�����x����4^�C����-��LO��ȱ'�$��ޑP���"��Y��;�°:9^T��"��^Ih�����^ ���y0��J�K�[?L'3��ݔ�&e���!��Q�N���x&n����w[ԑ��ι�E�5ߘ�B�:	��i)eU�	�#����Y�d��e%~��[@>����Qg���c�{�o�g(�:\�r��,�'������ʧ��	h�2��y�!���l-1���(�8��M�,/���x��w*��eaD�/���@G��N�{o�ӈ�^��To��r���T1���o�Sr��]��Fib=�t�bmkra�z�7ٽI����������`@�0V/�x]�y�����?��
��f��D_؋����i��� X�c&�z ����)}`���n�w�=���n��k���x��*`<v3�@8��O�_��������|A;�N�?H��m�|X��;df7R[�(�ʗ}|zqN�"�o{	��hsE沾%���z�ث��s��/�A�=tr?ڭ�"x��kz����O�N�m��̈́��N6��Y��1t&�"_��������W���'�a����ۄ�z��qr�oH�W�#0s�������O��N�z�1��5a�[��Ñށ|���j/�9ӓ���a�z���=!����z�vR��Pd>=$�n�����oG�(c�� �b����k�`�s�y�[���lԢe�ð>�1�3�i戹�S����)8вf�%�mܾM<��SX�Y�Q�2���a��tY.��Z?�5�;���2�3j雏���$%���w��˗/�9����Ã$m�����)J�Ly)`�z��+�=p> |6�(e#C,�
��u䉮[Wm`���
=��#�G 	(͞3F?�*�6��N)��"�fQ3b�D�+����2����^L��u���.��	ɑ\՝���B[ԓ*T��ǁ^��s�)M���$?S�����#��B"��P�f�S%�`7��*��C]]��,X�l�Y6��$�E(q9����X�V�gȟ2����,<��ݓ���A8�"�ڐJ���n�P2o�_r�����*�6�P�X��[?Κ�N�\�e7!�[~}B�QXB�|�t�C�5��]�cAx>[0}B�2̕	sl�D�Ι �Hri^T���٨���$�}�rB�g��<�+��0%FL����ݜ�%���o}�k�ܒ��2<�_ � <��(�������8���L ���?�,�zj�:���T��\��(���3��8E�=-S����;��l��&��7+�I ��홹�1%A[��z��9ƺ�u�5@��G�,�6�i�7Jwsko�Y "�?'}AF�:]̏��%��"�MQ%��N������7�V���}�㞳�Z��+�͕�ī�.���s틆���+(�P�$$F�1j�7h�p�lc9nL�C%�A�=�q��)?IF�U��mnI����N�\���V�P懽-��@ � ������v�p����S�������=i�ɡ�e�C�z�Wr{^�Xj=���^*K%�P�4 ѓ��yek����=��{�����˜�d-XeFT�:��`�7o����k��rM_>}ao���S������;�z��޼{W�U���"�Y��/�0���#�p���isW>�>��e,�^g����oǹ�:��O���=]�_�ey�{�{���_�_�(t`�^r�8��fCV}���Ots{��
/�����W�0�*z�n�	�f��e<�Q�Kg1�1���K��j��m}aO���S���=�H���̸i��A�n���w*W�~9r�G���P�2��̉�d�o9��ʝ��LALN���?��F����<��2�����
bȏSko�yۄF>�=	9�;�lj��z�}��O��8�J�E����
7kM�����+CA��O�C��e�WJ��@�]5��G/dfGE���.�v���+&��wROK�3�S�6syP,�8WϜh1�/�y�yw�lk�*sOJ�#�ڿ��'�N~�?,���^��L!3������R�4��y[%��%���0��EG�_�`&��$'��6�����tR˪0L 9޿�*X x��g�bFZE��F��a�����7�ZüͺN¾�����0G�۶C�:g�����7�᜴���?���e��j`儷��r�d�����Ώ�@HE��{�8�L� ��a~�O��ԃ_�`��)�_����K�N[_Ɲ���L|7�q�6���Mu���\��K7��Ѝ9�d�+|�V@�fQ�x�߫w�'�d��`-;`bDwE�[�7,���Զ%��f5N��&�͵��O��W�8��tϞ��f�`ot���Y
G�؉y}m����8�=�i=?������l&,Ie[8�B�D����P3[P{r�Vy3F�N��������P�7P9���Y���)�;񤜙�f����Κ��G�y5�8ڣ�{b�<!�>|լg�;�\�-���$�K��ۼO%���
 `�f8�/6O#`e;���Q�hֈ�Eև<@p��ƀ��#�ݒ��h�m�N�ѻ �򦬇=p�e�L�n& �n�������
jSI.-�s{��ŞOe�6}y�Z[�ؖ1�2���7��t��]��ʬ�@ iǪ*��0^*ɵ�ɼ�;rPB�߷�������W��eќ�*��y3�
^��'�D-��,$\���|��� $�s�!�@#Jy��r�����" ��j;�< rm��ՃF���:={`�ɮLF��t��6�"�����gԤ��(ˡX���T��n��)��~@�
����F��R�ɟ�����/����%�B7d�1��PW7�Ѽ�&{��(	�r���ށ�����駟��/̻z��s�� )�  8?~��>���k���>@nx���}0F7m��k��k-U�|}���w������n�o���V�58//�8l��[d	��^D�fx�uG<fHc��$�;�"�b��=<����=ldG=M�>�W܂��x�>�P�h��휿�f~���W�1��O��<yR�{jÐ�ĹL�1s�ʓ{����ء0�u2���j��E���[L4�IC�"��Qz�������{��!���O4�f���9aX'Zz���9��|��`B>�f�����E�V7v�W�^;��Tv,nv��_�VöϚ�1�c�u�@��W�d1�j-�Z�y�ɒ9�h�s:u�=֗�v�Ms�$�F���u1#�x����e^g푊�~)��z��g��~�s0�x�n5��{�����7��5�R�1F��sqvB��:^5�%�ر���/�L�ҾUa`��',���>~xO����� E�)[T(�+b�(g\-A��]ϪX�
p52��(�
���69t$ђt`�Eb]�+4���z:x�W��>��u���1��󧉑aKpqn�:�i[���M�����$7�t�$�t�X������+�}~��\�l�L�$9V:�d,�!ڠ@O�}�{��:�&�$���840U�s���!�VUҽ������%qq�ě&3
+:@���5/@r�l�"�k�?\ox܎Y�hh^X6���5���L7'�~L��{���k�A ns�<�:��r���HD���g2Uea긐�dQ�fe�S�ZQ�('�߇�sA�S`}'�tn6_�'C�� 5M�$i��E@)����6͖�O�ʸ��șoy�� �׫��^{>"\e�,�CG���Qaə3f	�j�B
hYs5Xg��%��܏������C��o,�fJ�������NÄ�w�sț�.Qv��-�����^>�6հ	 �����`��Z�I���$7�Usy��{���6��?�m�×(_"������;ƈ�S mw���f�����>��M�]3?�Zp9C^����]O(�V�nˉW��x_�ƕ�iA�,�/��Ph��1�\�2H���|i,Ϟ$���{  ��U��TC�*����o9�d�63�'��4� {�J�]�g�C��}��P4/�~�a�3͉�\�9�՚;9?�q8��
@<��
(�?���8q�����N�Kcy+�!�Z3��kت������U׳T���A��F�z�>�Y@<��	�����k���N���\�T������#�ŮW��Ɍ���߅� h��� X�כ�k��x�`����#���j�������%+ �� i^�z��`^��~@(ӧ闟�|47w��Z�-�~���䝞��k/e/�vRe��h���p	�Xf��xyJt@�j=�N�70��k1 �u�Z�9X7w�M�O鼼f���3�m�8?���5+�?-{����c�����y����0����o�h�M�dl�΄u+��eޓ�=��ճi�~T�[���<v�ok�c�L_�� ��Z��_CG��ω*��֢˪)/A��8�1��q�~V�X:qL�����\�oL�����F�Q���Y&��ʉ�'�%�����o)�Κ4�~����=�z� �
o���WEq�Й��ɬ��-b7}.��@Mv�7�XR��+9|QER�Z7��(�c0E�K���0fv�1�.�c�� � �(�lLխ�r|�j[%���b��p&cP�n3-�im�}�\C�Lh�mL�S+o�f�"� ̡�h��f�B[a4�< \
!QH�֨?�X>�[F�Ԁ�dB�$���pׅ��e�˳O��3˛�"4͋"?+�ES1W�����>���;f�X3�l�o8l�,cI�_�^��o�RD���.�ou6��1�O2���?�I���禮Ū��aM��їZ�{Q���s�������sF辸&[>�
&�m�>���,!,�rf]� �� �����_���*_��r��t�mw��y	g�����s:.k��dGg'���^���1ҐGt�I��n�
U�F�+�r�9
�>:����H�x�10�!�5�72���k��X���u��R_�K��G��D��W�-ݕ�Ek]�s�.����˲W�iN'E�zX�������"�e��g7vݨfbJXfwk2��@�8 &��^�Ck�ߣ.E��U�/��tXXEr�q�o�HBʵ���*�wz��)���5|��K��[0�b�{Y�w���V�[��خ�<֛JH��l�aYg�g|�R2���0�&��B����
�|&��V����;h���kB2#���s8+�fUu(���I��O��i�)D�U�!
GQ�r��3�z2.4]rq���Ii6lA�3+&�*���N��4�����2����d�(�`���0Ӳ��F��[��a�c9��u.U0�[CId����g�@���8�����.FcLA��X_͉k�AY�g��I��kh���p�9�1�)k,!�x�Y(��fI�7��̂�s�FY���5��+�S�"�77�)�We'-��;::]
�@hҜfG��5�'-�����1XDqaM���@/,����יÏ��d2��D�l���q9��ƽ���G�N�k���!te��N��VB�/�x^,����C���3����O����K菶�d^m�$���=R;yB]��&O+ɵv�A����n�s�4�z>���m'>��l�(?���� �����*��9y���,�՛�zG�9ɛ(y�������+z�����t�o������'��B��Y�!���$ǜ�����U���D¨8�vCV��~@a�P"�/��çt�0���8��qUx1<�T����L�S�n7��ZR笡�uZr�yV�/��ٰ~�п�V���h[��>uy~�<��������	'|~��-�A��W�zS��nCfd�T��=ZI����*�0�5��U��dj��ĞG�c f��8q�>��{F��'��6��1�v�/�� ?a�3U�����7�J�f�ϸ��x�c'�W��\��P['�<$ٍ�Y&�XL`w>鷮u���4*^kGt/�9 �\ҷ���y��Ȧ"�{�-��J�M>
�v�W�n��긥��C�zMI�9��{��Z>��J_&k�Jԁ�'�eD��a�۳��z��5���)�1W��5*���W�IIAO�TJ�.o����;16�DJn5Q�y�#��e<�rNeF�����pX�K���
1��������J�,I[a4�;�M��$ɜy���'Q��������%�!��\���	,��]A�;*��9�������6n��k�h?��̄���iƌ�@�㳼����`� uʺm�5���|�C�/�sE��nsaX��(1oEkE�/W��I���R�
0�.b��
b����,i�e�c_%�"�e"���7�Sc����)�L��&1Y� 9�d�S@���A`G/d�bJM�Y��3�s���m[�;]5X~� lVo��$�����A|(J�m�/wt��1��� ���<v�ȝ�?ly���yj�C&gGK:;^��WW���K�����­����r:�6�2�(dP�V,��t��Z�(�\�n�8re���9����:�ce+�C�m��K��v�\Z{��V|w	���W����/wts��O��ep^R\���|U�<�~��iO�ܧ�N��b l���1�"�4�W��Gm��� *�1�`�e�u���j�y0f�(iN��&#�z̺X�G��ꍜ)9U��<:ee*#$�#��ΰ�ڋr��ьZ� l�Tx�+4=���ɧ�;e}�sau_^wEh�xhr������~�������-����Gtw{S�Y�M�Td�q�{�9�,�ϐ���ؓ�� C _P�B�K��Fh�X�!g�m�����[J�U�`��e�ʪ-������/L1t����H&�<�7j���D>�rƴ��Y�YXJ(! FYto�����u�W��-��k�2�2˿�%Vt���˺oN[��8j��jɩWj+^rLk�|c�qa��+-L�4Z5��yn5�i���ʓ���}-�ϩ*H�7>��q˞7e���"��������$��-�e�!�	/+j�&�F_ �oEQ^��rO���f
Q�< �p=��9M�QR�^f�_��|�a@�����
�9�:��@�ۅT?c���n�r�Q���4�^�'��iTY���"�|���%�U�L��w�2�J��n>�:/^��/_�U��./�X.:99 l����zU�������a,��uc���tww�yM����e#Vͩ�xu)����B#ǚ��a�Vs���HuJ��|�ә�Z���(!{Yă��Hz�
��X����aٽsأ�/:���|�|J��(���(����+�<;��e��[e���w�圔6��V_IX|�����~`��e��?
X��d��-�|�7��7���C�SYL�of`�1{�c�O[�Ae�����]��|[~�,�������u�	�w��Ȋ��T0���ʱ�uP�};�?׶j$00��4
�m-�2�Iy�ϗ��k]��A�������yK䷼��-��rM�nKǷu�yKH��'��6��\�zu�ތ3�[�=���}��P���y��6����	��LZwfFÜ���[��z���w�@����o� ��F<��9�kJ��O�(���d\�&��"��}VTߑ0��+(ᓉ7i g2a�&�.&��vh��S�Tr�&Wu�-QM�;���̂�A�R�F����TDQ�V>qKu��h�^���M�QaCb\�
,����Ǝ�'�%$��^����t?�6��J&W����Yv� ;y!�,+��Yx�z�y�8�,q��G�OO���bS��\��mg��%�` ��S�g�U$��V��U����ڠ��U;��M
��U��� :N�O$��b!n�x��<�>�k�v�dA�=����cÓU[���W�m�E�N�[�%��*��<G�Rz���൵��ل�,��� mv�!��qiF�'�Hx��J�2��gG��Y����H���*�y�a���(#�L���X�,7MVpTT�$ �ݲ���:�%I���*Vd�|�=E}ǊV�My@��Ֆ����͊n���Yo`Aϴ.��Jz�1���x�7p��N��v��[:?*���h~B��u��f�ҙ� ��Ҏ��VP6�ƹ�0;���5m���d��p���-L�78O��G�O_7|��m�z|��v��m���,y����e}���z�Mt]H��UG�7�l���sv���*ӢC��#����(�]��\�B�fe<ge� �-Z:>����Y7��=y@�Y�jf��p\��{��c�D�kUy!WZ�<�x�]I6L9T]�-��s,�)�H��JY�/�pĉ_Y�[��{(<�Ї���W�:%�R�9�H��vŰ���=�mC�����>�qh+����Szy��Х�_#_A�m)� �͋p�_�t|V��I��Z[h2/�晝 ��G[I<c}�<��Ƶ�}�6�c�R�X0�k|�{6h����4���{g����,���6˞�(^\�8���<ɫ��ns8K"'�9��r� ��D	x�\G�Q���q��!�b�t�Ktj%痌k���R��`�^��ԣ���p����)p �Jze|�Ɗ)<j�[V��cbNf���v\A�W=A�jk���3����i����36�@�mOZ-99=���9 69LV��v�z�����Qy�V���}p�(/�k3x� �ā
������c�����3{Vh����%kQ!���0�[H��C�?ʻ����yJ: ���F�r�WWh�f+^�Y��kU^�H��������
¿a=e��QnW���r�y�q~+�:C�0L�W��SM���91#�揔�٢A�� �aY���}G���G�ʥTH^͚t�r����������@ ��p>����Ks��� ?��2�̽L�*��$��qR��"3b�C�$�30��ww���'�����o�<	%C��%-����VCF1Vl�mw��V�*�IN��V���z=�;�e���	���/�8�j����/�<z�"�k�a�Xh> �����;'��sl뼩�H�������G�U����o�4y���=����f�"О�8@އb;+��yk����;���*s��?����cc�]5�Z�����es�}�TwDX�tn�X��F�òL�1�'S�s"���e��m5&M5�k�$�s��!J����	��n��0��e�t�9 ,!W�J�u#��_�9�Z�5#0�F���"[�IE��,�6���%g��]!=;�d��2o�l�+�ʃ[/p�� ��X�@� � �����y�uL���L)b>{ߍcBS��R��Mb�&baH��iyPk��ګ�`�٘p	���ĺ�{o�Oapc�֘�;�U��sĮ����g�st��Ɇ�'.B�0�F�~��+p���՘�4E:��G.�����a\�G3�� G�`�=;D"�k(�+�^< �.�`Vp{��B����!a��o�J.`J��^��|�<X'�7~-��J$�����|]� ���S��s�4��s�# �������R-.�ȡ�f�W����>���~]^+�}X�׆A��,�&�6FtU��]�y42@����Y��E���-/;:_I~?�W�qQȎ�:8;.
Fy��t7ߢ����ʺ	�'܉����Q�I�]�uvI���a�p`�Tɨs��ڏ|��W5bA�V��p1��)��}Q��ym��JCk���C��~Fwe�n�~Z#�~SN���+x��.�ߓ�����o�a\�$��v���uT-��;�'s:=�e�gtR^Ghf��y�O,�'-Q��  �c#f��
!l�.1qa�����=�-��(i�r��S4V�����of5�xU6d������N9�$<q�wE��/��Њ��;�jP�s^;k��ue�T�����+?\߳ ?�����9��,|jK�e�;e��ʾA���b�e�r�WD����xX�j�x���Ľ�C�L��مg~v~��m�OB Mۢ�X�Asr�ϰ�{�Q|���'y����R٪�Ŗ=��n��#�Xuq�!y�̋Ɨ�T����$b��u�-��^si�dw�1�� �[��v��B�>	�N� e�̸��b�y���2�ᥨF' a,F�,�8=�c�C�y�. -��ԯzf F�n
/��9���1]�^���u������2T��2�`Sx�Ɍ�1v_ò��)�]\^��Çe^�R�+�;hd<uJ;�ptVd�Ӳ�.t|~�/x�Yiy?"]ךId
�;��g���0Z�.�C�pG#�r�m� �冟s��p	{!6]���|�
�}q�4��������=��F�Y3��j�
��m���q��Z���k���Z�cX+�V�Y����X�W9�<��2�*)���՛���&�d_�C��7�ئ͞sG�xF�s-���O=�a7)���꼪UC�޽���bH�&�?��|���<��HhW[���_�e��+}C�LƖ�6;�b�>m����k�-�Z�cN*��������=�=�\��L�]\�_�������Y��h�D�fOfه�����ޣ�8G�13�wi���x����z���~r\��"�C~�(����=��9�����:��rsM?~d/z�W9kX^}��>?���9��o�F�ZuP���sK�o�"*M0�n�B#�	����7���UjT�xv���&�"�\��� �6L�`���T�C��5���WC��-��U�t�['xA1���+Ա�!�J�_�/+����2J����U�T7�:�PXG�"��k�w�T$Z 3A�+��J�x%��5�0%-��BM�k�+�4Wڐ��pMz���b�Y�:%�28!�[u��B�p+��N�L.ѧ!f��;�0	��
���r�%�̰����|A'E�@���/?��  r�i250R��� �&�u�5\�,j��pr='΃�{۪R�3X�
S ��ŕ��rl��o�?�^�2!��@:� ��E(0%Sd�"de_��e��.�G֟���'�uC�6���3wE�ؔ6�G�x<�ǜ[�9+�Mm��0@���@�
%�{كx&���\!��|^�0ԎA�%_#����4/7<<n���m�`��!�L��C'�}trDGǧ,�m�]����?���/��L�	��X5���,���Q�Z+C��0�eyUs3���Y�9��{2'W����׃\�X���4[�#B���|������� ���Ct��ʫ�����zG�Ex�-���|:����.k� ;�������*�KW��Ϣǰ��PsrY�����_�ұC�ߎ� ;gE�*/aE�OY+N�=�^�P+�C����F�3�K��Ɠ�2�d㿯�&�QH��E��%��M4�2.s�r���OE�/�cU^K�4����ؙ�O3���˼m���槴i˺-J���G�o�"�e���uQ�vt�☺�s����lh�(�� �a�_���1����n�E\�����{�-�9<Κ��C|�^H��IL���zɘ�]�(-�{�@S�X�W�=+��=f��m�UO❚¼��)؆��BXM/��x�t�� ��<m�7���{��'�����Ӣ���(t�tW����R�`��F�(��P�Q3�D��/�Ԃ�����ү�3!/]��Pn�4��S�(�Z1��n��ދ���V�%�b�%gq=�::P�Z�ˍX�Հ�9x0� ��}�0<r����uC�ޤѤ��u��,4!"���v����x栺;��Y:bp'A��+J���x�q�1��U�4Ko����$#�>BX��yI��2{��b2�̑���e�u<�y��������3+���ܷU�{ܳ��Ix\R�!��x.��/�8ԏ�������g���>X� �i+�f w�}� �v�)��^����_|G'eN D�L������$�˝�ش�$�>Y�%���(� y�Ń�Y�U�X�mxN�<�+�4�Q�\>r��=���A����sO�B{�F��H�y�����04	SN[�4D���������G�������/��X�h�w��7
j�����>8qo�sP��;����3+���A�����NC�h�6�,�y�PW@5��8���󶈷��ܩ`��B�a$k:2}���\�����F�C� ]Y~g@��PD$:Fg�������u�ʨ�i���_TaBx>x#�>��<������Z����g���[�IHxl�ky�ӛ�� C�K�%911�c.*�ϙ�H��:�h���-���/t�.踬o�#�����ފ�˕�w�}(��>(��	mk�Tغ��sǑ�_��975� ��F�YI��<�֐���n
���DH��Ź��兽~�8vZ:��Dx��S
a��j�so���<���u�|���b�ً��V�^ת��܉f���)~gt��N���BC�nr��h��ʬt",�aza �"p��hu4�ema���*-��Gө��ս+�s1�v�kW@���� I�T�<J���X�Z�m�Ұ��<+�cĎ�:�~?a�0�� ��1�"{*��G��c,'��[:C��b��#ʖ �2^g�H/	l[$���i����8#�3��4�d�9rfyR�&���p�%Q7 i���] Ah9��~ׄt)i6}��B�{(D��(�W�(�B `R`�o�%�gR\e5�D@������")�#���}O�^����_�����;���2� t�u��u�e���?��?0c��', Pq�x(c�P%a�RI�a)�Z�srzB�����d����+ ��w��a�9�$p�����t}���W�jE1���($|��8�[��j�b0���Z�_�������%[�/�Uԝ��ن����=ET.���1��������;:��+w�߯�m��0C��ZMu$�� ��Z���ú����`�k�I�>�Ma�����������I�Tp��n���쭖��=s�|�?�F`y���@Y�4?*Bw�;�[��V��JEX(���B`h�^����a4�(<�Rv[���"�߮:�r0gK�E��wI�VH�	���Z�C��Z�	yxxk7��I��v+�0P�f��������%]]������$ɍ$3��=�+IV�=��������Ϙ׻}q�Ȫ<��ݮ� 5���b���<#�O35U( (�\��ֲډl��Іs��~-���v^���>��Ӊ\�L�t:b�x��Mi��m�F5�e�ڴ!� �=�elڶ�$�?���ɳ= ^
��a�1�P�3Nd4A��D>~�Y���[t撏��J%���i :��jp?�:�x�j��YZy�k4�MԼ�1�i��A��l-�ߏ���K;;��������켤`��L��� ��v��B��J��l:��\��9:jdd9Ԟi7�b��桝�e�G�L�3n�.1`�K�Yq~^To��I (�	�G�ʐ[�T�xpP�idrbTX&�������.ءd��u�!�u����׋�����������w���U���O�>���-;�lʍ��Q�[���`������jd=��*]?�7���˻�ڻ�|��xO�3ݷQ¨���Ȯ�QO���t,S���XF�1���d��J�-�DK� `�|�{���]P�K`�����Q�m�;����24V0��d�DvA�?���Qi�A�J��`��$�-htm7�XY�h �ha�@���@m00q��J��љQ���p1�����=��j�U�o8��j ��W��
�w�㛟��2�3�s�܁rكؓ��S'�n�����������oU�K�V�e�V�^ZJ���m�Y�0W�:(�5����m�d�6�߾x/o^����3����/��Ӄ�7:�Q>�k��h���j��7��W��Tk�8���e����`���'Z>���6%��B�@���c�^�A'���Q��Z�����b.��.�j�c�`��Ty���	<o:=��`N�����6���ί�M��2:+��;��֩�vU�F�	�F6+��L�5�	�I���P0'���?_���=x(ә���Z����&��4����.����h�*�d�D�X)!b |A���ؗ�[�\V�^dE��^��%ɚ��m�����.}�>�X �n�:�Nf��6�4�#\W�Â,h���������G����vJʲ"���(m=Q?{ 1�?���ݻ�hQ�%�hO��c�D�~�2e�/�3��V�g�r�߁ߋ�(E��� � �����tA?�7�C�f�!?}�,?�����o�A���Y����׾������ǜ�? �`o����b�QAa@��t{�׹�n(��8?���"�|��|�^�����r�~�����+% �����5��1��ߦ]�X0odb������)�&C&|��аA�c�����tV�ol1jc�D����:�z��r�/\�/�M�h��m}"�&]�>�h��dy #G�޳n3$��I<q$�6 �xo�&;o�T������ō[J��8�R���=צ��#|^A���i�ʂRH&�_��o9ٳ�|����,�u��}oy�P���������1�c��X�s\��v0�	�7ܰ9����Ω��,"�j���Ngb�� 8��y���ӑ�.��/��|���+�m�� ��'y�MfZ�e��qzu����&>�Sv:b�ԹeT��A\�@�}S��Q���,��3�i*�A�,�{|�N7��Ý���4�N���:Mo-�Fy���@$�J�*�����������dK ��|������lV>{�[/��\��>�t�%�������^����K�`̱�c3��!�%Y��7�jtj�gJ�֝���ا���t���y��������À+7=ft�����F�	�{�|�������j�n���^�5?�;n@<8f`4� �Z7�T�oE|�����B�ɩj����h	�A�M�b�1�	w��3���4���"|��Y�sk zk��̭�as���l��wئ�#�m_�1uP� ����70,5�zT��nu��U�����j�th�9��M���ϩsgi���������$������T^�~���D��!�D�Jn6 J�������^�����`�ݲ�s+�n�SS�[@Ȝ?�hޅ�N�"��v׏w�i\�㝢�~���^o�;��k���B���'t�S��,�O]�)�/8� � ��; �!�.�t�:Eu���s�A�R{������f�B'�C+O:>w:>�0.�5`�*]3� � \o�[��p�!���B[C����BY�-��;+�(P�hm��#����)=iҴ��霾��ټ������Ğ#=`��R���4�+��C~�L���#���;Xf:ϡI�A�rt �m:�m�2��S~!��GYMv�ne������/��KF):��D<���R������4� X[��lA��s��wk�|�� ��(�A�.�rsdx!,&�M�_��m��7��7��1��+���^ g1��^� ��ֻ�����b0R�bL� �t l���wx+G����Q�B�е�ݻy@�y�?^D
����,a@G�۠�6A��K��-&�T��s2u�qH�������8����Ԧ������n@����~d��6z'p���1���]�6D��øG�΂v [���;c�`<���7,�ҩ8�շT����Ņ�:)o^���x%��N6g��2�n��|?9�q�����c��YB֨���G1f+�kS�z�g�:�V�%[���B�`�x>�`��dސ#�Gd���)�/�����M����AS&��X۽/���Ն�i��r��G)ލ>`b��]��(��i��v��S�6r �\u%��?���[����#�R,>��^/���7�)I�)�dI,p$K��A�sċ��1I8b|1D_g�i�����W�~�������Ӈrw����+m�w@O_ �`��p�-K� d�b�E�;'��m�i�8�{N�M&�tߴ��f�f�w��e9[�W ]�5HH���w�� �dc|��q�xk�捷t�^J�ɪ'���8��mE�I���������S�H��sݟ��B+sw�٘��h������bf"��"@ʏ�`�׷����	0����+��,�'����m$��xMH�R{�p[{��®��b�f�E�;+�u$�흫�d�_���Cy~,=0:;��^S��h���H��l��
�� ǉ��9r�9��}i��t��H���4I���l�Q �<،c��E���V-{v���aO �?�+I�����E�r��'شA�C���s^P�o����g����4OF[{������/^�x��X�����?m�1���s9�B>}���G
��0z���5|��)\����6��]�F�� cB���b�A�K��|AJ�X��dF�x���ᣬ��SC����w��r%���P��S2^���f�\�|///���ؖ���?�ht�旯��u�|a|{��|
 ���gP�������������Ѽ���
.<lUl��}B�y�d��2�oC�]����[����͡5�*j�q��T�4d��J<t:�t2�°���7�@af J����x��b�T��(�5���Ζ��L}��@��I]t�>�j�������J#k���iI:,�%m�x4]Ǎ�Zrf�~ad�����p,��P�cp� �6��4gz���!Y�xEp�7�Qb��,���ډ��^�V���i���Z���Y�,���Q�O@l�B�u��Xо�i��4�XJ�z�yk�V��܂��);od6�P�i���w�,�,��Cg���H�^��vM�x�Ǉ���<�u�3�qn�d&w�<���2�$�V�1՞��g�<֟=�S����p�ñn�̆�Ȳ��`�c0��Ow���h�#�^\���JVzN2�e��X �X�32@ �iк8���Gl? ���R����~���DF'��5�C}<�l�LrP��������n��d�'S)��t��V�Z��-4h�Gx�ӑX���m�k�o�ו��7��`�u��K�$�w�<HhDr}�%�-H U���4t��,����� =��-;�	uEj�������a'Oӕ�_?���G=��%D`� �`7-�����z��e\8^d�Y��(!���T��vd��Ӛ�RTo1�����D�u�����ܡрb�OB�h�����h��ԙi�^��$DN����/�@�/Z}`��@i�ې�{�s͜
�����ZC�[ݛwxS�����D�ѩ��[��@̾�����$ C���-:��ޘX�۵��\>��a��
&�/��2hK1� ���:��A��"c�a�QP�?��7`��X�3����+�k#����. w_6���08�߳cP'@O���%(	p�!x0G ����� 5���P�zZ�>:��j7~���e��0���2p�O�����LV:?3y�u���{פ��v�˯dkvB�6;R�u0�K���U�bBc	�x�k���'�����B���O�N8t	�Ɓ��Z1��� �|�����-�>JU�=_�؊�?�"��D�����3P� �.Tb�ff�:�?T,��XC�H: �7C2O��{W$�]�)���8�Aֽw�x�@p��*.ޞ%{]D��V�vd�u�ٜ�s��p�Z߃��:�ڱ�8��v�Nl& ;`�@�&%:����M�d���*1���#>b��2����D����H��i7(�L��,XWvǀ�P�1R�e�d�U0a�`��<ɓ�?�# ��gg<�6�I�����> V���MF ,(�Y`DGR��@w�����Z�T��R}\�U��� O�2�XKL�������Vz��Z2�N�<��q���Ż觙�]��_+"���`�#��и������=����Ħ9V]�(��'YB�$�B	s��-�ķ���*'���s��!~���6�%�	 �D8����tv������֏7�`?o{\:��;�4�mwp7����;> ,�b��&���4Zo��ng�H�g�%@'�g���S��{��k�M6[z��P���6]��ly�����;�)��ۃ�z[o�zaA�u�<Ucyyz.�gtfV��Q�Gd�h\+C]q,x�l2��E���1C_��Pt��|�Z^�}Mcp�u� W���uh|<#��X�&�g��1��a�մ�xy~E�#�4�����6����}i��̅0Ő���rqqN��d<U'�Q��u�^\�����{WlQ�s ��oc�	�E��X��f���^<���$�m6���6�m(���{��a�ֳ�hnbp�D�/�O���#�� �z��gt��o�z�фe�( @�Hj;uq�`��&YB��`{��銺������n���V�K�9P���p��s�׸�Q��f��9�)���au6��Qe�������l��Wkg�Ue��Z�-u��۲�:i��P���駿Μ�n���t�!��<,����J<���t��4��^I��"	���9����D����e����;��������s �PC���!�u���:�D��9�����'9�CS����2����Qr� "~�Ŝ̅�έ�n'+�Ghe���	G�@&�P��e�){����������JH��Ų^�X0w�8�Rms�6Iv��| ��ny9+� ԴP�����ÃN?���Q����D��?Ԡ��7����U<�Z��A����d��i`6�����1/6r}��ׁ�C}0%(֬Աl�F�z	�&B��P�y� ��:.X���/8���G�Ӆ;M�=9��m���V���(�v�˴���]��(��{�Q2{��,5�X~P�As�`ʍ�I�u�f�KA,3=;�'��[v�W 31���J��2��%U:���!�Ȇ �� LS0���{}k����(s��]T�%���F�xv.k�0�qm!�FW�f��:A�C�?c���u�һei��� '_,-�N�5s��b�c ���Y�����x�U�D���V*�i��$`�/���o�����u3̌={�g���X}��&�A��f��D�=Y�f�!qE&�}�4��js�G�l���v�]O����U�����k���2^gs5Ⱦ#���Q�q&>2�C��*��c�z�#���
���}���_�Orv����9[�_]���Tm,Xc(�����-[j�.b�L�)�{?�� �6��)Y�W�
@Sa�67pb2���Z��XЍrF�IL1��C�д�,o<��Gr�	z���1�m_����mVb��:��r��sg�4����<�^�{��-�tQ��NX:&H:·�W�I�ҥ
���u�k�@������2Ĺx��9��6Mk�_g�k4ʏ̍�Nx=��c���e���F�e��K�L�s �|hdR���dC;{���T��A	V�,V�vԩj}<m- lG	g�c2ؼ�Ѐ1��,��Y7Y�N�|ֱ�;@��l��?)|^�^L ���#g0I��UJ��m4���Z�l�.�zCk�nw'�5~�9a�]m�ԏ��uBM��e���A��w�1	M�%�U|��(6�����6���AJR'߽M� **�+����aI1b 4=���Hs��ΙP���ڻ��x�1
�m�|�m1��l`,/�UM�>V"���X����L^��~����AI�ǳwU۸�͒tLܘkI��6�����Ib�pv@R�@$�3���Y�5�Y�Gy�*��3���.b�d�^�����!���$~�����~�y� !o��M-�%�.#���t�D�c��1�,�9q��.�e�S��rk��AfT���ώ�Ms'��[�X�f����/��f��co\�l���LNgi�2�E9Wc����CGt Z'�����q�ƒĒQ��L,�`�Qs���ky����y�N7���I*ԁO�s�Z�ME�c,rI�4��7lT@�Y�:����b�#��$�홉�S��N�qQxi������+�c!������c�_���|�:o�Ŗ����$4�UB�c������>snq�n�#l��h��c��G
XF��7���駟��c� ��8GѮwj��)�&8�d�P�y�%хs/���ۯ.���=�`��{˭Zy9�e����p �6�/f��e.��V�gH�xpRf �1�?Ǻ�洆X���9<�����P{]wcR5�A	��1 ;��Q��j�����e"��J�N�IC�@#o�/Tfv T��9���a�F��6�� v
׫2 �3p`)�!d�Zfgi�@������\ǔJ R�z�嬯�KV��*����fm�Ŝ��߻]E]�5�SX��φ��F�uܫbL=�L]8M�kg���#t#J���n#[����鬒;=Y��ɜ@'Y8x�M{��`K�)�l���Mi���@�;~���� 	2L�N^.a��!��8�܄V9�Á_��KZV��_<�/]1�ns3�a3M�[V>�k����a-??ȫቜ�\����`����GY�Wr��U�la�p� /�u8���%��e�3����Lu��ù~�@��;�(���kq�G�m��zp�ur�ޣl��LX��gd�9�&9�:��<0g�D����3'���|�4�2Ci�ۂ�,T	ЎaDz�v��|f�Xb��N�Z� �+��cQ�`��:��,џ�6Oٓ��=���J�u��;�6V"�@�n�I������ʣ�ũeT��Q�z�@�<L���9طK�mΖ� D����d�h���8���d�1G��ܩ�-s'�~|;����v O�,�a$��u>����D9�kʌZ:�چ��c꠭�~�70��e^�����%v���Sh�@��#�$G�gHQб%<x,�|}�k����z�1�A�*71�}e��u5��%���?�T2�lԜ�/� H���.ɚ�ql8@�.�����GkK��1��`���`Rű,tn� jy����~o�Um/���x��J���g�r~��>�������3�Ո T��}��X�M"�j���N&jO�L����`������w�@�Uw��I!j�t�jKv��-E�!&�u?=��_��ѐ��V�����ޝA�H q�7�KTp�F0���O �0-I���N��%
"@�kp��Bwj{q���,�?Jf@4h�@��7w4��r�A�bM9�&��Ƚ}?��,��c��ܟwJ,8ILv�{\c�	H���d4C�/������&t�g Q��a�לZX���Y��-��h[�c�h��.)��Y����1����D���;�:Ӧ����l�P���e�b|0���E5�4'�îT�O� ��`��-+|`c	6��әL�yV�V���z��boF�
s�4������?����i~��\�����̴t
g2�.�//K�ԈJSy��ԅ�C�CwOrs+�?~��}���q���l���=�?(+<юyMө���|�� x7V{8d5l*����������mؕ  �&��B�k��/�)Ϸ��0�	���>hF�K�n^.wa]��z6]�6��39���zc���g��1k�⟝��ҁ:~S뉮��1ia9�����:z_��u_���>�t��A�xi��̤��i�o#�w*�ѹ�ޛ%�M�ǷV�J�x���k�-�5�k�k��������T�/�J�M�9�A�m����o.�x��:H��.65:P`���t�(�~�(?��'����m��2�8G���¶Τ
.�������?ɣn�ܞ,N�����w��Z�3��IS��~ sդ�&��%-�trjL��W���L�X��G����X?��61<��H��/@�+�(�2�Zm�^7KU8;��g����^o��`��YʦHޝC�w���=�P�;�)��gd�����Qd��O���@ܖ�l"á!,q؛8$�bf� ��Af	@�u�
���O��v�a���q�2�O�s�2p�ӂ�B�S��-���9=�iF0��jE� ���l��4� x8)���H
7���E�Dn֬y/�`�l_n����C��Qc�@4�/v�w�@����e�ݝG���;��6m����偊��Ɇ%�%�4	2gI�o�P��@3����h͂ɜ͕��5�{�@KOp۝��.�}=okϾn7;�;{4.cw�-�m �&� &	2d�A��͊�O���{߁ෆe]m2f����(��Z-�X�?<0��@d��面��aʘ�zpL�W&b:ZaM��j���m)�Q�j^I8[�q[Q6>�&6�Dݬ���ۏ��a��|���TP�lD�Dkxd7�ր,5d��(���-J���0�U��W^2�� �]�����G��~xH��6E2&F�e�k�&3A��hP���ǋ����4X����:4T�>	�-p�OЈ ���Y�#���29�6��n?��(۔�R�{��(3�����~'�p�.K��z�a�R�Ձ� J=.���U���I V*�9�N��"h������aC �lYP�9t��2�2J�� ��7^�`�m=���ñC�.�h�g�����ڟ6�2W���婍Z�/�Ǧ�c�

#�+�o���Y��o����xc?w��g��Q1�r��mޟ>/尮�e�nI��p@{�N�w�ʲ{���	��������<Y
��ݘi��\��^���R_+��/�� '1L��}b @�Q5���j5���/�?�>�V;b+Fy_��m��������G�G�ft��J9����;��ʵ1���j����l~@\5�Tˍ������~w�wd p���*��R`��X'���9NX���8�� ��ߙrB��ƴv�J�`u,���W���f�����R(+_��3���EĽ��ڔ�o��{K�=jZ����t���l,����d�����s�=�����=<�$��`%Z^����(Ab�$���q�?��OeBM>�>?8"1�ܮ�^�1�����H�CS[ #Ȳu��J�nn�鯢�hv���7@�y�624���`{���a���G{�m{K�x�M.�o�ҭ��`lٍd���o^����YO&�[��n�_x]*T&�0� ���˫K^�e��w�}8��ڎMJ c���:������,sPǀ$|? �+/_��`�f���i���� �&4����n�HH�����D�N��Z���M\��-��a��a�y�13J�Ѝ��|��w�L�f���L?�v���L6?��">�c�a�p{K�tM�ٸb��S��~����;M�]��b%b�n-w���jώ�� �s�%@��c��K�W��=2љ�}��<�Ŗ�sJwg� ��v,q8���`��N;K{Hj��1r��������}�n�o	L���.^v�xV�i��o�H|���9�$ aV.z���o��L���&w`g�@偄w������Ib�.���^�!r7i�M��Ɵ9%p��rs����+f�G�ZRu������'��������⁠K��Du� wN�-�=�`z6�����R�C+6��77���Qn?~2$H�gJc��.�	�����w�5��]r\�� �!���ݷ��'���;PC�?Z����M�n�B�wvvN``)�z~�ՊǄ�1D�AqG)�SXϛ.��h]���LMgX~�[4q�ѝ s��$ ���:� �AM. O�2��r���Z����6G�)���h���X}a�~��`��� k-�w�@�C@uH�ޑ���1��R�vwt��,�����C0';�u�e�g9��>w����G�օ��%�� #���iM�93��Y����~Ń��s��vL��l�ǣv?��#�^;�2�>��hL`��Fk׎�D1_�Y�� �F}D#��C�=�:��r
�\[���A͠e������̨�S�в���e�Ń�s�ݵ�C�X���w��u��Z��C:Fy�����^V�'�K8#�9T�_#8�����f����>?Ԁg ��j'zs��90������� �� k����������fm�1,i`ן�!ꠢ�
����Zn�}�b8f[x�-א^�խ��_^k P6�4F���@|�Q����l
i��ı#�`͎������O��hL��� ;�A���z���!\�v�5�*�����X�-Dh�y��t���B�f9��-�̲�>h&�>)���H�}+t��<��k�JEڴgp�֖�@��������Qv�\��iM�NWњ�JX05
���	������[��tF��5�z\��(%�2�;�N(�1� %����#`��t�2� f���f2ͥDw��5��!3�>�tj:B�#�ꗹHxd%}�;=U����Wn��CPvh��C� X��xH@	���5�Xjp{�������/��կ���W�Y1�f�8�D�	ж1v����M_�0	���N��a�1/5���R�݁e��!iG�3������B������O�v���,�r��Үԍ��Fp�DA��i���:`�����f�ڦ������5�@�Q��?�%�嘝5��,�J�e<�@���gIu�R>><������7�`[C��1�OYb,س�]�N�RI�Yܣ���+�Kחʽ=~"��S[y��l�Z��+�q����y�c�| ۞iN1�139��"��<�#�%Y�$�u�
|1��.\[:������g���~/�^��`/ދ9w���GtsҠz	z�����	��ѝ:�������ع@t3��(��Җ o�e�9��F�#$D�l�M"�*��"Q��m�Q�N��Q>~���[��r���	?V������� �F�3X6����g�k�K��xB�9/?�D���O$��:|�vdL���sU[��u��R�XY�.�ZbT�2���xY����5�m+���y�"�d�{�0��ؙ�1��@	"�H:c?'P�|��ٌIf �hq�����X��`��6��K������!��b�����u�~r�"�o�������,�/���Dc�� ^��lX������⫙�S�Q�|f�����h����:���tVN��=�N���>(������_��������e�NĔ�$y�x��7�l���C/���nk�����+-:`'�*���藌Jw��//=��;�ϱ�����]xl�:�_��g<� ����D�<��0X���}�ŗ��j=�)��i;��H��C0�R��3w���i��wP]� F�;�� �

�Q/����=�ٳ��C�s���0�O:*�Ⱥ����t���+2!`$kwD�az|����b�����ȋA�؄�1�#х	(gY�<�S]�&�{���x>%(�� :�4NU'�^����{�X�1�]5<J�dcp���R��Ew�x8nO�hCih=�n�zC)����I�H�Mv+�o���g��_���M/S�ߋs�&����q<8>�p�@��FU����9�7mrDƬY.�{������9��h�/���u猲�.���nE�o�0�0��͊`��Ѵ�����X���ݝ{~HpZ�� TE�3�����I�і�sVd��JaT��E�쒙Q�";����:?@��x�#�8���;� .Dh�m0���<p�;c�kˀ��Y�]1�^�A�Y�͡	�y7Cz�u�
�`z>�Nn۝ږ˯V��e�j+�B	жld�(P䅓a׺��$�~��T~ ����8�C�Lбf,�)��s��b�?�#�'2�;���'�H��EF��k�qX�����gr�A0�¯�%�
u��[�$�d�|�,ȯ�e_����:�Ib��+` ���hvw���wk�~XS�xvr&��Swj=�y>�`Me�������=3'�?���'�@2���T������f��������n�r]�F�����N4@N�f:��Ap�tIv��#�o�:�e��fJE<�����0̰�B";��oZ�������9�R���5%�Y*�����R���$�W�yD�X:�Ö�Q�om��T#�ؠ���n���3%�Q�����ԏd�gr�Z�(�ٛ-����9��kcqb���@g�4�y�0��S�tio�):����^��(:�O�RA{%��.���m��N�����Ad�� V$��G�	����1����ے�ʬ�.������>����I��%�-�Z���YE4]65lj�y�׃Z� �E���wtL{��C��S2�pC�C�gg̚��S�MF9������Ou��|�5V�����U������p:TGL�����r�q�~��1|)�������Tr�F`�����5����66`���;���q<)4��iCY��{mTq;e�t� �o�����:GO՞H�u(̶&�(�3�%�z0�6�^���˛XΏ���m��m�nu>�]X�xƃ�]�&*û���}p�;�׷�����@��ӡ���K:��==���hV���k�K�v��`� *L����1%���i�5� �V� o��d>#X�=�8��,�Β)0��ѽ��^���Xa%Co޾�������O�/{�|D�������k�}y��Mj�������O����<Ƹ��`/���i"G�S-%�B
��'�/Y�n�Ё��/�MǊ �	�	�o�}�y�Yw��k+���_�#ǻNֻ���V#'8! ֲ���|�굼x�p�c���;�a���V�f��p���F���%�	b���0��w��<.q�L�������!�@�Q��l��0��3������}|�����l���rY ���C�����81�����c���M�.���l̓���O4�������ѹr}, ��?�_���$D��G���E�s����Dh
4k�ޗ{��W�����m���%R��ǧ���I���-V��g�|�������3vҷ�J��}I:�8�(�2����G�|}��c��6݁:m��V4�L;���S�u( � T��<]I��_;H]�c�C�t�A�ϕ���L�i���6��,������p��,3�괿y�N��K��[b�V#���Aq�$�/�gm�L���a �YKƹ���A�p�꥜��{7�� ��lJ�'��E�YQ�T���#�����<`6�4:#�MQ. Pt|W�S���٩d˕u	;��Xl�W�7���Z�0�4Zj�_��cCx�6XE�?����=E�ʲ���7`.����	ر��I2Bn|����[#P¹5⢠��ǈ�R�%JEjn�,i}� @�6S�x���^o��<�3�5,s�Y���T��X��p���묣2�;�U6�̄�͂��'�d_�୳k�~Ly�&�k���Z�m" 
_c��N���j���s�Rs@����A�sIJ�^�/=E��D[��D?��:6�O[8w.�S��f�έ���Yok�)�/nQB$�0�����k�!Q'�kcw�5�	�ݹ\�������=B����� v"S�x�,��3��S���-��� �����奼~ۢk6"ӻ�U�s �D0*|�k1W�=��o?��Y��괼��Z6@}n��ʧ�G�c�q#�3���]��~��AUȨH=\�|ؐ�F){]{	"��i�c�v��4Ft�p��_�R�zO s���e?�P��L�r�vj�v�h >� f�P{�]k���V~Ftu�CK& �x��Q��0�u���4�3������
�ۿ0��렎�!p�'�G@w���^+ <��#fL�H��\��֬O�� v.	�D(�e6{g�6�e��s���Pm˄X�Ѐ@��1S[G@&�'
��9�v�$�.fn��0�@@�^��h����ٙ��X�}'��1��%�3	�����Ϝa�)�9��Y4O��H�iq�By�� �]�D.O.���?��n#?��$����Z�ە����%ZR�Z�Pn���^7���8wp�HӍ�w�Y��1B�|� {d�p��7���+MDT������6�dqI�'X8C�f����!�� ���$�A�b!Ùi���C�S|�l�ur�a�:�r�/K�j��p`�0Ѣ +a�Z���A���4;�c� u2���p4`Y�3� @Kv���q�{|��m���;m8'�]L���n��%�rd��o��E��Q*E��xg��ڄ�$@�e:O�z�Xl�h�[?��N8p��>��k��3|s� ��9㾱��ӏl���~6?���U���<�{���ل�Lf���x� k�&;��:_��zqy)��u/�o>�}p���O?�IVOO|�8	{�%�4���[uG�I�׿����oK��l�CŒy����fԓb�kG����?�@�6�ԇ��������1$��^�MtA�B�`]��x�NtZF!V}ԽK�!Q;�R��N�� )��Ȗ�cwݵ�%�ŏY�o�_���XYZc�r�I�_�"c6�^ץ�qT1�-z��-m����GR��u ���̞��tq�Mv;w$��ܒ�'БT����8�R}��W��) -4=q�S��⬊�Y5�{�=���?�����i̅���c�181?`�/s��_�l�xL�-VpFO��[����K���l��_�,�UG ] 6�G�����@��8f`xA�tD� "Vɬ�k�P~SK*�r��=�ۃ�zsԎ�6[c���5��6G�;N0��t�U��!���&!�߲�	Y9�!Um&����E��#`����#��k&���h.�@�6�a���C֢#s&]w�,�;fQ��7�g(\a�&�� ��!3fh	��cYo�n�(��º7�89�:R'C��
L��i�@ˆz6;sF؉-�_��WW/�ڙ��&#H�ԍ���j@ug�����nM4�>Ő��Mw�(��|�R��4���ʪy��j�`K�4���-v���8����I�di���"d�m�t��NY t�y��.��G&�F�z�smB���g}1ȿ��˾ag������p
Թ��Q�����f� QS�k:�E�Ncѵ'����?�>�#D��FB��1�G�+mژj��%C��lc���2v=�����S��sk`�)ӷGΌ	��\G��;9��Y�C��L�ծ��'�Men��1 �"Y�/7�.��[�~�k����M��8k�"��5k	�$~<���1l
u^��i[�f@_�.�O0�̸�_�
1�+R�K][+�cle�YA�,ʅ�R��,����5�9(뮱wls��
��%2�g:�'t`�BG�u�о<��o����Ll�KƔ�6��u�߽��J�\�ʠ�� �J�KGB?�8�u�j�9�]s�3��5�=���nSG$~^A`A�b�[��Ԗ�Oh=tL,u��Qot���]#�y9A}p����PV�3t��Zi,�~j;��:f�o>R����{X����`㔵u�j�1�J�(_�@]*�~�I�!��iȨ���э��6���sӻ�س[����[.���!��>��#[����	����Vh���0Tz����G,ƾ�"tc�A���1�7�ٱ� u�����Y�W#�!(��A�$aTT�΀��B#<0M�bZ�xѽ��@̾��D>�BA��؃Kj�mX�m�Ǜ{�����'��n����$��H�@�H�k�B����#��Bh��/�8K����t4��w'��w�˫��2(��vt�1�R7͌6�`G*[��T�9��^��LM��d3�9�T�Z�H;��Qve]l�,�P�FH5��r-
��� 6�r��%" Q�`N��Q�@w,���yיۍ�[�{�0���@��ɔ�~���0��%rkώ���s@�l<#�s̽v[�o�b�% �;�e�I'�Lg,-L��19��_a@���X˽��^�C��J���Y��z㶲��w͒�ښb�S�@T��) ���p����@�l(�<05��mL�I���z��S���Σ��������ξ@)��r�wf�	~�|� :�n>���΁�?��3�D�������O� 2�Q�{~��O�]�9�`������S�(i�NRX�H�4U���u/���R5d�j�4��f�8@��۰S�߽7�C���1H9d�wò/0�[q�-�
���6��:NQ�jo�>���z�w����������� ��:ƞ��N�?]�Jmf��^�������㰫[����=U���"�[�2>������k��,X�	����+X|�Zi՘D��5��hl��b�N˹%#�z��@���nR,:����¤��|)/�^0�C2���;��gg|�e�톱<����d�5QYp���N�9�*mqq��!�qM/�%q��K�Em�����e�U_����k�/
`'���ɒ]�(@� ��$����mS�2���Y�s-6R�|�uN��ڼcJo�z!?>��g�"�<�=���;��-���e���*`�+0�Df�`N�z���G���6���m=��#Hp#�U��3���1���g� �i{�aܹ�T�������֒�v�#6΋��J�M]���z3���w��)�����p��*�6�+�ӝ.�S5�'�P���B��Vj�h�׃Z��k�ch��;@�K]�_�b� �۩:>�띜���|w}�:��P�f<�R�A[^��ﾓ�߽g�K�W�����N��i�]{Aв��@�@_�쌋N16���ְ��L�����\-9��"��Ą|�+�`��B&����<��/$��u��_���^Gu�Q:�f����
qeZ;1�B(��F�t֑�c����@A`�˷�:�����U�-w
j�ۦ(u��JB���O�t����-:5ц�	�*:�1��k��S���9m|�;t���E�;�Q��N:[�B�̞�uM�ކ�P��ۣ�r	�v�ĺ{U�gK����G��$�MC�� �Z���v��ah�A��?�B;��/���E(صɎ��1�nklb��s�b>�FALtL�m��9�������mY'���>ϖ�D����s�#(6���b���u7���%��������<>-���Ħv�Z�����j���x $z��;���߾��Wj����R�����^
�;�v�.���uʦ�^�U�#�\/���J��� 0�q�m��f�~=�k�� `g} ��ݕ�?�@�����U6K5��Im��p)�Xd� ؁��lh�R��m	���3 ����ȷo޲=��R�J!{��T��@ j����H��� ��\lI�!�F�.�=2QU�?vJ�YN�5p7�_����v<� g~��y��@�1�cqy� ��7`������� ��Tk��R��@�%��xk����m�[
O���=;=�=v-k��IX��fG���Y�'��PZ� <>!�d!���p� ����s��A��`��50����������TN&&,Vƅ^M���لsa~����,�"��8C���*r�����O��W�1v�B�;���'��>�N��Y�[uy�B޽�N~������T�F�#YNX�c���� ?�"x����pHffۂ�l%g ԥ�w�i��X숌G�����AKa��)K�؏w��܆��F���s`�q��TmoCpl/5C L6:�L���G��m_m�|m��	���
�Z�?����D2s � ؙ�:,�u������a�vG}��޴�`7{%y���2���������5lo�{�N�ر�n�B���8h���-|�I�HiM
=>0�g`�c����+K50�5�oR���`T��fە�s�Ӡ����	�!��V�Io���k�<��':j2(�kל,�q���G����9��o?��'�|�*� ��7�"�����(l�K����o�$vF�Y�6b�>����6U�K?0���3�GK���h�':�w8X��{&]'#ة�@�4����ܡ�[m�����<�Xv��
@��  Gễ��r.}=�B�j���
���o^˫ׯ�4�u���?��ͭ5� 04z�V��v�"|�6�1���vc�PS' 0r�H�H0�;�w���ĵ/=��� `��^���(O+�]:�8#�ե�9�E�B��yw�~�]EEχ�u�E�r����� �$<�8������v��B� �i��z���(Y�|y%���ԃ�RVV�\;0�9:HkK���י���Y؎ ��Z����}�>�c����@�ޛs/N�q�mK���X��{
����f{5n��!��J�v<�'e˨��U�;"��<9�4Ť8.���k�ޱ{z6�R�}��=Ҝ�ݾ�dv�aW��mh])H�'����@���CϺkɼ�3U�5�t����Za�-��]7.d%�c3�vέS�#�A�b%�M�G�Z;����W(�M�uH�
��+C�&F3�vZ�(L������{M���ƙJ��{FYߩc�8;!���[m�\�]�|�������wv���-&ƆH��P�a���N�2��f6a�֋�������3t���քp`8��{��ۺ��iÍN����3���4����-��ԥVL�Y�P�@��#�&���@��a�Mb��ڶ��|AdM�xc��1����5�𷽋f]FL�`�x�<���3����R��d)(�m3��;���]�M^�AdA�4��b���O�����5�y���&������J;�'�9��F���P� b:"G�n��LF��ư�|Bv�}U�0�g���#�aߩ���3�<[b�P-kuȍ���Ǐ�����j�vx�%���i��4*FiS��lR��;���L*��>_����
�hg��2��u�c9����dL�rw�װ��gCuV�+�樂]�C�Ƕ���f�װ�RP����x ��-g	M�v>�r,lX�3c=jخ6�5���(��}�rM�ɺL"�C5RGv<�|r�P�a!�6HB����R���:9</��u1�&X\8�Hk��8 �ſy�J�ԙA���N�ԡ�n��	��F��b]D:����nǷ�w?~�Te:L#�E��`/��>��I�5ʃ �A��x��dh+>`{���2��\�ծ]n�^YP�F �����4�BK%�*�{��1��{���p(�C~}X���z�!)C����X9�ک>W�s�<f;�N!L�ݰ(C����YM�Z# �Z]���cT���s�I��JrX� �S^
��^p^����Yntu�c2v`� ����y�[CO�`%.l��Z���@\;���`���A� �=:��Nlq�5�|�}踜��\���:��3��P5�n8��f ܰ�w������V�Mk4U8]���c9[�k`����Ϙ���������a�)R����0'�c���e�o�k��jC�<[�ع푧c�[W��'�s<�Z��*sIh�t���Gp=����Q}��	�r�6�`֙�1Wr/�	f�޻o�G�^��p"�V�j�#��-�&�'�QK���� (���=rY��6+b±�N�1�@��1�-^��:��s�@$�2�R�.����	�y\���K0��j��_I�k�i{�����d<G����8�i`MA�n��*�.nH����f�q,ɻ�$��F��d����A�p(��z71��i#�:�?Ï�����(]s�e'p�Sg-�(�I8^��g�	��������]s��v��f�=?L�<�.~��>nhSo���g�> )E���t+�H1N���ٯW�/��`��)�h��2�<,��#��KMS��@�oA�`��z|b7]0����'��%;Pn8�["��f��FY�z������w�}G�?��5��`������a�ѭq��`�ZB33���f�M"t7=�Ź��/�ӵ󩱗��[i<4������k��Ēp�!۵�����{j�ŒQ♘Йu�Ͱ����؀c'��FVOr�p�NT`m�|q�_�a���L����Rm��I~��3�����Lt/F���6Wk�YY��V��|H;�
��W7.썵1"@����c�����<�9p(m���>�� �PQ�}�����arR�%ʴ����S��S7&�<`s��{��R<��A�Eږz�Q�dA����z��I�:-�`��ϳ8:����,�`چ�� YS�`�h	�*襢s%l�' ���I�*+��1�pn��<!]C��K���I���'��rc���dL��@���czf�MH1�W�k�~������ֳ�_0���T�ªƲ���ceD0��+��6�#�� 	N>a�����B�Q6��; )F#��D=-����v�D����0��a�]������V���~�𺩒('�8ߞ��s�k"nb5�A7�A1"	�_�a�U�^�1L5�zyv%sl��0I���qq�	�EM�q���ld	��YP�+3:��޼����&4��?�s�Сf��~�y���?Y�GвW�|�if��}h����	�e�ND�t˽��tsF�p�٣Di�������5o�Y1G-o�I�*��_(���+��9�#�@���،"��2�B���}|&�)�������vJ1�����vR�'�C�-bwl̙=8�c��T��qz^|����Ѵ6�����V�#�El4�����ł��[��nm�rk�0h����q��1��-���<�sak�n�[��1��D|D�`���M?)��ߔ���M��/31c��c  �ր:aY��}q�2M�ϊ���TR�ո"���vnm-�C�o�%ffL��L3��~��Y���/|�"��Y N1_�.�������F�-ڝ��r��wP�2./�>����;�=��
���R��F1@�js)��(j��TF(E@�SLX&uWG�5�;�@F��N�m�n4��6	^j��#2�O�%<�{8�tP�뽱l���:F  �A�J����%�zp??;�g�:F�R=�6�^bǻ#P������=�N�$�_�{�����e��:�B�&ԛ���w7O�0o)l�T����u6Bp�l����v6��[r�bA���AD1
���pHY�>�$ĝ�':�0�����+��nR6����\{�9��[�d4���z�׵�q��Ou�M�9�c`V�(g'S$J�a�z�5w�+�szyd�����5�׉��,�޹�e������q�"p>uql�RZ:�U������]R `g������O��̄�'���f)Ò6z:8le�v�e��$ #�^0`�Y�.�̰p�[�.f�kN�u�u-��c���� W��������r���c����tm������vF]��[�F�):�1H#0����K22-�n�$h����������J��2���Z�J��^��v���~��ʂ�~�������kә��1�L9�tw?��N  hG=�#q0�@o�>*� @[n��w���넣�|I��L#@^q�g����h���
9���y	m#h@m��}y�����z'��K����s�k6+i��lP���hS�
l��@�p���Ϟ��nA>����T��=���˰�>�@2v�*��9�����;�9������X����+l��\?�[S�(����c��(�!����-�@��f���5;8�͡���'�%`������|��6#�e	�F��#�7��u�2�?(�U{N�*Z%��6�58�tCv<+\�/^X2�!��h�@���T&%@��'fh���,��G��t-�w7�?`� ��m��[�1�����כO�|x��+}ɫW��	
�] �>f\�4��^#	��UC/G1�	u����غ9b\��d|)91�8dv2�rMt�h:0V�J�"b6�!�f���]�p��h Za�&����1$�ໂIYWcv۴9j�c� �SX�6s� �O�ٮ�q�$7�w���'�ǵ������\�u|��Ā�?2aBP��ޡmh���:�(b�ITu���hzSU;6\���s����^�z-���`L��\{����\�\���aǡ�J�ڐ1!D������w��Q$�p`����<{�u��e�%�G�d	'I��b��&�sFw�*iWFIR2�}7���Z���~�y���+�eK���"ڨ��60��5ݰ��`�!f~�����Z��]=��������ǘ"q�j�h��ژ�Y���q��:�X[`�㱶ظ鰂�����2z�w�sE�$�A�+�����/;	��?x�a�����
���ZG��������z�1�[/p���7%F��- Y##]�8i��Ҍ�>�[�:}^�`4�I���x���  xEJ�?]�y���A87<���m�!�l���ǭ��n����X���Z� ��z<q6\0�ӉV���S�l7�N-S���	Z�/�m���r�����9�)j�O���AMjH`����ԩ�HA{u�����zG1�:Y�јLH��:��6����k���#�Alc�%I�p��{Ft=W:#[T�#�de9����cK�hF�]@���M��Z]�B>�9�F�tX�������%E�v��)����0m�����$!����>;��?q^ϲ���+g�T{�XZ�00��׮� ����ZY���K��>�7f�X���m�]<�F;ɒ�F]wƬ�:f�x�5�1p�m�U��c�u<h,x�e�0W&�ږ��T�.%���um�|p#�N4�áL�[s��4XC��W�/X� ]�D����pz&z��*�t����|Zi��s6�@�Sf�.zL-����i�S��X�S٨mU�^Y�ɰb����Zx�mi��z|��?��B}�n�* �DǪF������2�p�3��T�6.Mn07@\#u� �>�,xdC�5B�	A+�7ϕ���w4�A�%�?8�[��꘼x�BN��g:�C���:Ӏ*~�ƋSv���<�W0��ԙi�n�]�I��Q��L�m�  #��� b��L��[��,��ߌq�5~b��W[=�'yP�y�1�-�w�բ	��3so�7�5 �Ȱ���4���33l��<;c����ӆ��a&�5��4$/СB�([9;!P��#�2�lž�n�k��ӽu2q�FW���{ hH��,��
���@���l1��̤L��eb\+�;��zL��3����X�3���)�K�l�'k��1f)d����w�V(�P��d�K���n���"Y�V}�p0�Z��42�KEu�
�&(�>џpʱ�R���|�:qeҜ�|(+.�ݮ�s�	^#���ҹ��p�_ǣ�L������r�Z��Χd���-�v7OM�M������Mm���O/�$�k�d���#�<�1+j�6����6��í��>QG�eȽ�M8ܹ���MhH���f�º�1��Yw2| b �D��(ŏ���ڤֳ*�. �hM�s��;Ş� f�Y��t-+=�;6D �ɂ�,M���C�ž8�i�����澇y�5�����b&�^�����N��Dn�&�̠���	�@#$�A�`\�%?��-��!����͐1��Q��MZ͜�͵��"��K�"+pY)=��<��v	ג�&Pң�|�]q�ҧ@���K�����f�����'�\�04gx<mW�����ZK�^W2���A�>��u�_ �v��>���  ��IDAT<�}����$t3��_�;�$���Ռe��!���@!}׆��J���X�Ix8�])Z�B�6�ʝk��.�{�xb֦����izZf��ܙ�2}�K�h{��5tl)�JOtW^f� qQ޶�ʁ������Yz�4���GgY�'����8@q� 4e0N��drMrKH Nc\�g�%���� �7��4�����6tM���|��'2|����b��Q��y)?�*# I�����jK�K���1 1T��^A�Qڱ|��q�*S�	��_8.�@�ן��͵<�e�\��_2��<�9��� ��N#6z`l`W�p�ʮ��V҅�$�Y��y�`;�G?��ڭ�J��@��S��+�b=Ll�D;����9`㏇ck��>�%p��3/�Qz�|�"����#67�J�֔���g'r8���u����(s�uy$�nILϡ�W��g6��9^y�gړu�11�>&}m�$����5v�S K���]0����`c����!8C�A������PzN'������}��eF�I �����3~R(]\�a&�i�\��>p�@s3�tJ���B����ýLG~�Rw�i5^D��K��.��,C�t�,Q�b]y[I�{dO�p!c��,k�ǂ��N���+�]t^�Ɍ0���!' ��z��&���sц�v����V���眀�n�����8y1����{u�wD���N`	�����l�: �������&�D��H#;+���������J�(�������X��uЦyޟ�M�!C�l÷6�m������.�KѸ���q2�S0�8NH�4�Jm�]��)�4��nr�䦣?�u�D�W��v��eO��%	�)g9���#�Mm��V"��~@��ƴi�Y�x����[��9x͎�!d0�f�h�4n���Y�p�y]��`���B�SYfI��kЫ�����ۡ:�̀�Dz.\�yEvG�O�ޱ��Vz	'�����)��߼/߿�-�6���{d��x�2W� �y�:�oon�aƆ�>�Yy��%�o^�$Pf�DG��ad��/������Nq�J��I���3"�f@ԌgE'��-p��K����=#�=�U�1ۻ�t�U s@N��lB�^���pNfz�$*��@E�U,X��,P@��N��O�=B&��;*e�Yvg`���0���s�K��q�R{5�Qy�	��}�	K�p��������'���G6k�B@��(��i�-�\יo���$���;#y � �Pz��vP})�pW���#�����31N�ڢ�qa�� 2�@K�1m���	�����3f{�no�� [��r�\�vA
7ْ% ��0�O9����I����I:Csj��O��pή-tK��[����g��zO�F
��"_Zj�dt�C`1�����	If��R<�[������w\(�X@�V�#fma �6|n����g��F�@���No�yIpt �����zMf���3s��5��VL�Z 
��.y���w����Sh��>>L��!���~	3��;�c��t��l�lb��Gm)J���(��<Fv���eYM+&�&��[��(E���b��v8�u�-�#+��p1PLY����5�v�\����?R�%�,�s��)��GY�������64 5����]�m+�H�͇��mĭJ�[M
4RS��l0� ;�	�޽��{�}�G���?���,�;X4���Q��-�ǋ�;����\M��3ے���']�Z?VO6  h��s���;��7�K������f!������$VZ,�;,����~,�`9��q��iT�����P1��%��Θ8�٘����ceglu/V�U{y�v2��Pd�� @������:o{��0�Dd\��%�$%�	CĻ�I`���;�0�ZW�fآc0��Z�X�s݃����Lx Q��.ynB��9w�b���.��(�����A�h��蝶`+�9+��s/���}�p98�>��Xt��1M�ǽzxd"~��<�_��c�Ƶ836�q�w	x���z!v`q�3G�\"vB0g��	|M;{��1^`��N��#�ԧ��ܚf���OF,O	V��B'4�p��ʍmT��{��?�,7>�u0�w� �몙f�ٻ�;��<��`=}��g���e\0��W�����gDuI1L�L!�m�U�gfmՑ8��������g	��֚Ɠu�+�f^�_��B�}/����0��+�Ų8=�Ca	��y	a_w�<:�cbn6�%�y�Mv���gQF�-`����d	q��0���"��t�Z'W<Rpʚ���F�i� w�b97�Ӷ)
���5�FX��TT�D��9�� �Q?���uC�WO��ٰ�1�M�[?!�ټ��LRow���M�v��D��K[�K��/0v:��х�uD+:eБvz1�j�=�F._i���\���.��'94tf�:��Mr5��L�Dt8֘[�+0��e~�=�v��!�v!
�q �������]� m~g�B0Y���P^�^0C����aǋ�#��Ȅ���B[��Dv��(s�`�QZ��8ڋ�1<.��㇏�Pod�2��<�"�N���;�J��>.�d
 ��V�N@��.Ne��qra�a�@��z8��B�A���>���j�߫CQnvV��cj�?-���̤����3=�0۵��0�<��[�X��@���D%�����zAl�5��2yf�N���I{\w��T�MBkC��i-�ֆ�J�jl��B�M�s�,�;�Х`� }�);�-���DA��8���:��� ��!�'������]�J䐃��wwuU�����#�p�m�53@wUef������ȥ��"mT��t�ɍ3��k��Mk��1�ᩈ���ʶ.���̮����˟������D�%(H���'[��+YB�
@�"H,����a-���pd��<�+Q0��.N�����s�݁Ǟ4{o�,\3��Y�ؒ��wKIK�]�b}A"�&�Ģ�&%�+�'$�������)�h�dդ}���m��H��\]]ȜW3�Ql���ʋ�����;vLXp;���� )X[�v��߾}ǹ�_S���

�����Txc��hv�,��C���)��Ϻ��
��kY�"qA��J��B�0:#}}d�Wk�W&�B{p3���{�щm�*��q?����2̰ %��UQ���c�"��x'�UD��C����}J����#h9����";=,�3�P�x�#�;U;�n��T�������6�Hx��}Z��ޣu��_����aV�¢_��V���{9�h]]�v�K��f�c�`��8G��ː]׬��tF�tq���`⸥�+?#�X��9��)�A[0f1ة�#�y  _'''L���Қ&0��QM1�?��2=o��Aρ¿��+ӗ��b�Y�߲�0��,�+h0���Q��u:�g��N>al������[G�;P�f�}�2Rš`�b���u�.w�;+XqF�����u�Hcn��YXN����1��t���:_9C��4�Ld]�&Ӂ������γ���C�9%dј��	�=�Dz�8�|W�rƂ :�8���1^����XЦ��z�<��Dj{��]�-9��A�w���zJ61�YwW�a�`�?$�cgX��j4���g8Ql��'� ֤���(���_<��͚nXG�'��O���,��	��|ol$�Y��x���s�k���gc䘥�)Y-��J~x�[0b�:I�b.XH���Q���������{襡p�����L
μ�݃P�K�V`=Io-=���k�`�@�z^��r�\���>��<��|o��KZOm�o놣1p�{����Ë�VGw���e*?���jDDS��{oh��C'�wjK��Úw��&~��`\�C|#Q�9G8*5	S��=��|h�y�(��Pg��c��p�.ᐅ�	Vl_ ��0c���T�LR~���RzY`y ؈G����Lf�񰪵�`�Ʋ1 v�1����D�`�Q�א#�&뚁a������0y�=�� >���Ii�]W�\y�3�tFffw~��9AD ��C����R�"{���#c#}~�x��;�9���\��;b�,��J�� �C���t>a�f���;��x�8S���iv���G��M�<�'��h�H��#����Q��-ɾ�����z�z{p���hg?�0�IgvL��&�i}��-�S^�4������8`[V���:�����8s��R�A1�\��U��i-!F ���ǧ��L�)�G1��?<�2�e�اٯ�u�K���Ο��g@ ��RK���'��Lf�D�?@݊�
� ��.=�������`�@*�\�%�D��O,�	rVF͕�%|&1#B��i}�Ѐ�����ǲ��������?>��| }��?c�E��<��AoL�+��B]Af-4a�9�戍[h[P4|F��.j���H�����@�L��[Wٽ,��td�4���%���r�22�)���n�X{���<$W6�T����I���61ϸ7p��F�g�Ƒ�%��l㯿��h���0r��x��:b:�\�G�~��t0��p���?��h�����T�d���[ݭ����sLis- VM��4:�=�2F6��>�biZd���0�ͷ�;�Aa��M� ��EJX��ƍ���Ikݦ�����k��k�s�'�Pt�|n�l�f���H<PP��9��ܺ����_&�ҙ����ɳ�ź.�ϡzl��&D�`gk����}��Q�8mX;�{����);�����tg
�k`���9��7W�<���ND�V���^�����k=J#=+v���z����>�bAɓn��O���"H�}��بi?˴3�5:���܊��X�&�Lv{K�|�f�YZWobk��u���y��[�RM��܎Ѻwv�az��mku �1�:҉l�k���Ƴ���I�r1J��%�n'�e��G��mS;(T��X��)�[��{����%�8����~J	y�͠��K��6z�\��}�����0����H����p4�I��_$��k��VVk��
��ؐ���*e+��g;��	��!����o�u�����9����L�n����n"tG�в��}���x6X����ů��JU��$V�ӟ�?��qJ��٩����p{}���Rђ
ɔ�m׏tO�Z�������� 
�^��ݮo����z|�&�ގ�Zp;
F�w6��(�����]�ښKi�q��X{���XP�W٘�r1-X�SP�Q��٤ϖ�E��[�7�:����� ��w>�������b���	�X��m1O���9;I�[>A0 �z��=&]g)1��]A0@��T����WƋl�WwN�/�p����|7�c�t��]��Or�p���Xb@�|��s�����^�[vR�M=����
�F����Im�)���k�˺6F ���Xa,6PC�0%_�8@g  u�M� �.$����A���K&?��>2�M��x�f?ĨP:P�c�ӌ����DS�?�L�K����}��2?(������Qß3�z':'�ƫ�A6�F�ڸ/�����P�Қ��X/���0̊�<�w+2�Z2V'����1��/Ǡ;i�`4�!��n��q�!�E�fYo��!���hS�Gra>��c�� ��N�	o߱X�ז�I� ���b6��l	"#� \ `0IW7�紧���)G���#�Sͤ�Y���
����-g���g�Hw*^��{�6�~�N�[L8t5_�=���~ç��̈́*�:Įa8�>X��L8���Ɍ��y�O�c�n��1M�aS"�a$�H�]�B�XO�]�'��"%��K���Oǝ��=�F�)G��
6�4��jf�,G^�=�:���ϰ��C�5�;ׁ�oݱ�ՙ5�4�ܱ���Y�OÙ$S�4���$a?����z�����e���ۏd@ޱ!qO旮S���U|-Ij vȆ�jd-�fs ; ҷh �i�����9�s��01n��b�8$������\��e�H���=��p��cA�Ĕ�F��`:<��V͋�wSW�c8��:!��,��iCo�#��Q�ZtVN��NZsh�T{�4���O l� �M���]��gi�,�x���2��ј�7k���-?C����~?��c�����4j;�h�V���{��Ө1,`�XPy�B�߬_:��y���u��Ӎ��|�cf��g폮��N����$����kUsɛu.p>40�0`*0���R���Ŝ-纒x��b ���/^�W�/	�x!���1,�t�)/L1���
�� @��88<Ͽ{���[��U��RBQj��u`�V�AԘK��qp�3��0���Cz��u���w��-���� �W]n�Q+b��)O��.Kɩĵ�����+�bA
�.����X���bc���DY����^��H �P�����	 ���&���U ���TZ��UЬ��p��O/?]���#���5pr�!ǁ��/�Hr��b�y����W���!�A�����Ê���*��YkA�T�5A�[�&<n�(�T�����)����4�x1Mf��Q���D�'G?ۂ�Îg۲�=�,G�{N��	����)�-1&�2��p	uF��Sw)��M�n�)�|����*rӈ��D��L���NW���;q Ӿ�������]�n�Vj�ogtCv�0zՕhv��p�/O_�ӽ��7IA���F��砷�3	�*s%����
Tꭊ��DT�^���ۆC�t4?�<���J;����E "���9�ݗ����AhN;&���8��0iT��<%�c!Q�����E��;2��R\�����X����`_̎���ԙ��!L��a÷�Z@9�~A�zz.�#�+�&й�+!Ca������_�PB�E4�E���+t�n�5aN��E��>(4��χE��2�YN�m�������gۑ�*y���$vݜ�݇ 3�ʾ%�'� �������f�%����6�n���<�l��E�{�q"�mkR%̳3-{��$0Z��)�]�3k�|�;���0�3��A�'�x!:�6����0�I1� '
��u�Z�UD�l�Nz�քs+��v(ṳ���k�D{��Hm�$_���$�d�C�c|�T�=r�R�B@��f�]�3��m{;G���C�*�$ج$q ȘH���xX� �tM�� �i�TcN��� ��G�젱�N��YJ����5�^G̊�t�P�yG����V,ԃ�����s�!��7K�Bnb8��jñHu|PTMCg���Yz�`��`m�J%�-��x6d���L�
$���+EW���7CQ{yy�y�Ã#�Ī�t�w���p�3��A��!����j�rW�(�3n�E�:]#:���a)�Mv��Luk	���,�7 �C�l��g��:d�6�`��ĥ���i��B!qZ2E!��̘�8TG� G	a�l	@c��3�� R���I�`gm�t1���}k��b���SZF�Y,4�p��5�p�9�)��./�w�h�L!�	�@Z�-�SŸ��0J5�[�w̫��h.���FJ��Qr�lҙ	��y��+a,�(�-7�l���H5oΈ�}ѝC��b��s�A�1g<����/ٜ`��ڀi#QH' �D�8�_�r[���Ai���=�k�^W�Hka��#xh��{��ƶ���`�N4�����m_��6E_�y�����O�{�����_��6@E��er{��l ��-�k��b��K���V��}�G`�����p�# ��n���Cv��XQI���4� $=����������gA	��82=_2���7��'>/@��Q�g��.����܆��Mد�|�x=4����>����\���ڞ� ՚ϒ���<<�7�͏����E|�fG���r�G�h�A�����z�!����w� ��9�h$P#�d���%�C�!�(��<j�4��A���r���v|ϡ9��WoY0�kf|
�f���w�L,+�{��=ٺn���3��LSQZM_������cM���贶�I�(�hz�}0Q�u�����#�׶�̓�aH��%$?�H�Ysݷ��Ts�@��t��z\3����ي����X�||o��g���Y��=ttz���O�YO4u^�o>>���w/^��>y���}���3Y�2&q'[�	��'p���}e�4Dj۔ƚq��3��L��O�c}U�Z��]�Ih�kj!h���4� Vb]��笣���½L���p����"��#ϐq�~�b�֭�Әۂ-�y�j���'�������&���k�2x�eG'��y���G>�������^0�xtz� �'��Ĳ�(N�����9�7�,��b��6��l� ���C�Дx�sFQo�\�m�`��ż�{�*�|���"6}R����#������Ѷ\��O.�m2&�2�Ck+/�b_|C�����썭�yW�����#�7\���I�������9�[��� �Y�I�g��Ի-4��Lg3�3w�v�}��	{d�B��N6���>�����ҳ�4U��z��]X��LC4����#c��������ߥS#��~�Q�N�|��6�ʀ�gwa�[��P"���f�
��u���F.���Ix~|�;{N��nJL��p���8a���T�J����a�挤��#v6mT�7P��|/�Viv�X�ݧX+H2�!� M6��l1��$�H?/H���+���"҆��5߿tK�N�o��d�D͒�A7f;���f.�@�f�+#�u9++~'���b�u[��Xh(|f����v�HK�h�=�C�XpBM;�~}�6�����u
�n�Hg �{w��ݗd`Іܔˑ  P�z	����;ݠ���IzϦh�[PCba#MMq�]fa�����g_<�Ҳ��a�GT˳eQ�)~���Z��L�a���N�m�A����Z� ���g㇊;]�	�Q��!��}f�;���'�{ߖ�B֖�����@.l]�\0m�`��m��Q��O*=�C�-
��A!�����:�T����s3��H��� 6n`�k�3h������!h��X`��UD�C��(0 ��&g��w���3��������)�y:վ� �$a,ڧ��w��Av��ʺ�8^	�I�AB�)�p�[�i!.�A�;xe,���@��7�u���;���b�	ԁ`rG"t�9�;U�[T�p��+K[w-��H\��ڔ�n"Gwp-Hư{��3K�D��=#\+��mH����:=�3;�bs�D��0��_�܅��?�?������9ŧـ(�!d��C$�(�Y��SՋŇ�R1���֛�����/�:�^�Ɠ6�;[�w�W(JH$�؂!:�ӑ^�R�GG�Ov�78+w��HϪŸU%�]���D9��b�ݣ8�k�Fl�Lmf_ 
��
8�
�s��s�k���;�Ui����{�D3R�����F參3�'�B��θ�y���� p�����l��Y��3%=,��	{Zk�[C�XS)�xmc	��;���؀]g�s"J7����ل�TT $ ���uvT��)��k���E�3l�N:Xy`�=��Q.""�Ĭ�ƨܪ+��	����}X��a�7皮�$Om9^`g���̘�y�>=
����}��V�.!^��n���~9���E1�x/� ����������A��S2`v9"��>���,v?A{bjBʦQ���(i�r]Kc�zz���)�-0K������?�g$�2�
@�X�{�p2V�q��	|�3'��q�JyDM[:R5��o���������#(��:��L�ƶ1B��#�+���\_X�>4�c�;��R����������A1�~yؤS.I�V�>ހ��5\wY�=Z���)%ft��jL�5;mȣ	���`lv�=kL�F̉�Yq�N ������z.R���?b����|��9\Y�}^���~��_ vj99"߄�,Ư��@.��i���{\QڀzYVx��Z��HT:�&4<�ljԁV��O)? F�O7tb���̵0����"3�	 �r;�9�j�x�a����Gg'�|��l���K���[�Y���߽|I��׈qȑ�\~��=�O )<�������@B#�L�I���ȅ�G��p|t~x���HgV��۬��1v����90r1<'�Ȱ� c��x�m�}�����7�KӋD��D�$9 �kۙQ��Y�F �3�vwzxLF�Ś)�\1!�Ϩ���k����NNO�t�C�y��H�AhBj����a����d�c �c#�g�;��j�3��7Nh@�ǀN�vX��)Y+1|q������	c/X�pW���3��jtj���'���L���	 ő�&����k��b�{g��6g��j����2��6��;�Y���sv�rՊ`�>����H>G��\yqS���\���y<m�����Vb���'YC�y1[��ac/��4��;��?�3\�u;��t�Y#J��ŚyR��3��?�����rv}j���H��
�{�</O_�����E���*�~�W�L��S�:x_0\|,��	*	����3ً:4K�~�tf�\Ox{j%��B\-)T�!0w���0��Q%8c������d�8��8\��t�v��md"����p���ã���V���Y���"�Θ�,������M�V#�s�z��8H�A�n$
)��A�"%r��0@gᑳ���A\�5�,**�@ ���+!{j!�`��p�p(�oR.1s�>��)��I�P�a!W�IHf��X`t��(��;pV
�%]���`A���F%R�B2dAX��y�Y�[���3~���E�}�xLJt�A��3Ƈ����N��ek֝��	���H��߫_1����, ��osg��~t��Z�!T� ��i��.P��0�6�f'��?�Ͼ4X���g�Rk��8pq@�A3��
:�u��^�6<�8�UΑR�l� �@T�:�E�-t,��n9AW�Tx>��m�Q4P�!|!vP{!ht�0�3���M�>�5�l�#*2 �\@$�x=�Y1����v�v?��#�2ȩ����b D6E��A=��mt��y=����`�}�hf+&hm1BO��b;��lSA֋�g=�gKV�l'tv�;tp03��(�:M-'\+�*�	�zB��C;Y���ۣۆ�ׂ����PK1q��U��?]��>��a���l.S�g�`#Ս�a��W۔ʋ*��s��F64�~��m�E_m����A������\?�)Am�cT��	��R�莁���'�#s��%jH�j�U�ZYL��-�Jw� ��S����q���	��Y��A�[��,;(��L:#��H-�^�_��Y
m%��yZ��JcuS
���IS������`t����gMKx_ۥ���t��p�XE�y��z^�eZWS��G^_��q���u���X@�Lӏ�u��� 
¼�>5и�Ůi����&��ϲ�.�*,6)!����mq����Nf������,��nZs�����M*cG�N�N�J��j�U��gf�&G�F���Fa�}�P��@����1��4��x�q��LNB��[�S�퐭CM#�s�����C��Ņ�>�ʀ1���,����`�={v�X��a����gq8��b�!�#����N�k�X-Y�<����W2|C|�������ۆ�n���in����\t؄q��*$'t%�sX��<8�� v;o �]\]���>��� ��"1�\ˮ�v����b��;�4߀�k�'+c�z�5��8�N�%�B�`� � ���a��ր�A;�	k��>��adTZ�e�Q6�B.S�����=_��)4MS�� +���toT��*�%�\
�2v�����,}�6f�c,!�W;������C����C����ƙ�IG���äռ}x$�
�:���7F4'�s��*����V_�I�#Qqh��J���=Y�h�>G�g��C��x^�G�d�`��%����
~`^�p����~y�&}���}Ƴ8��\{Gϑ���/@��)Աu���k�E����c��/	�B��t
C�e"�.���Ƴ!��矊e4�����XՔLp�{<ۍ�oSԎK��&�t�|���e0m�Q>���Z�D�ᡵw�yh� ��5����Ѡn,GgD.�;��_���T�睱�}o8�:�j�5ڛ��F]���^�y�����U����Q����{50+cF����>8?��B�@��ͭ�E�ڳqs˙��躇v�
�(,���	޼�M?tԉO������'Z[#MX{!c�X{�g��������ŋp�w��e)��]��8q���r�2M�̠��B����[���`����	�Z��ZP�4�iOP*=o|ֳC;��z����؁��7�҄mc�'n�w��};�9���m�4v�a��A��	�9����Y����<�z�J���K: @M݊M:�hff!�~ �`Iް4!�h�R����$Es���\�RR��V�o<L+����~>`�{5���ɀ �.0�g�zvt� �<�i�,����P���K0,����i8M��X覢�u��ęW�6�f� /���A��$:c�Flv$/s�F� @��#��L���x��@����"!+'���=�>.��'弄��F8H���`tt��lM*j����m ߠS�p�ҽ����cm�ĕ#J?��0ާ�����xQ�>��r����Uq꠴1���ژde���2FE=����#�ƣqN�_��[��3���E��#]�������d7 <y���[ʮ�p\Ĺ�I;��o�g`����rRz�{�N6�F�Y�$1�Sp�P ����F� �"6H����/r@��N��������~�d�l1�J��%���2�ńL2~&ށFG�	x�<:�q�hL��sϓY�G���Z�5)��>]���u�����:=;	'���;�����b���T1�0`���N���P���M��6f��Z!>�ay_nk&c�����ϲ�GB��I��}�Vb�.e]L4	�9�b�}at e[K��cf�t1]�:���: 3�>����Q�(��wS��������������;���-z`��z�1��2սZ�z�Qn�� �X��s�������9��y?IHB̉
��a�	@��1������t�b�VЈ
���~��;��Ho�6�=�?��'�d�-��c���2W�vX?H&�%c,�쐣��U�1c�98,|�93�K��f��4s��h��զe��I�xqq���y����ئ5�H:3`��	sfAh�)���\aQ-Cє�]0f������Ng
�)����)�]"1���F������DN]��_�00;����=�����##� r��I#�@�K`�b'n=Lڦ�fĔk��7�M��CLl�Z�qg��9����g�ЈC�x��^�)ޥ�E��ڴ�p6Y��/���? �+猚Z3g�S��"��Ƌ�6��8ù�(��1�7�;r�T,F1�/
��@�Fıĵ��#H��p��@@$-C��⵰'�`Ra�K#|���m���M�
{�>G���T�c��)�P�Z0�D{�'��VLH�ѧZ�lx/�c�����s��2�^߆�t�1m5�d_�49��G�����5�T����r���ٰ��1������Oa���� ���@!g������^l�c>f�;���R���GN� v֛{��d��fOm�a|֮�F�@�Ď�x13�ɦI�`���`Lo��ƚ%]8ņY����3���/(~��G~>�8�1�LR<(Y�o(��.0�>~�.�.)J����������l�ћ�����;� FG�Ux��8�PV�ɺ�r}�S��iWJ����)�����p���������w,&;g;�����S���y=���|�h}�<Xc��f�+��ӧ��D��b��Ȼ�.9�
����@�*3oXl�(-�moB=����/՚V���b�`@O�<������9{���0$-�67��\w0�A��?�8���Mz�Y4�٤�5����;��[k�S�|:��қ08�ɐ���qR\x�_�w�����	�:�+�H� h����95J]Q ^�o<_�� ��8z�ɑ�������e��q]f�*�q����	!�11d���'��	V[�'�*�`��dn�ؐ>X�`�����^�
��	/�=�!�Q�����Z�����5�8���3@8��W������C۳ެr�Ѯ*;�!Ǡ!�9�b��p^@�`��� 9�O���E���)l����y�s��HZF��� v�/��Y�QK�}g�}�vxx^��
�'�l�$�60��=t@'%�	g��%��������-��a�wz�i^4���pĻ*|�Ċ4�'�M�I���@�D�աkjY��,�&��ZUB,w�C���iJ��- Bu�V�D@����u��<�z�]�=9`����r�J��뇰�<��I@%ݛ�����K��A 
4��0 Hwv����s��d@(y���{��1���L���9�ub�i��^�fI���(�/�sQL�Åd���1@*П� ��C0�C̓�?����׃3Wl�K3�s�@2 D���l�u��*�m�`>��v_�/�4Kg�H3��c`ǂQg�x�F�`�;u���̗!�3��(��5d��V��]��$��Rr�(4�Xi(���O۰_\�3��oԾ0X����{(��+�7}��rT
\�K��X�W��Ǝ*�.]P�q�TU�G��M��A:D[v�Vr����	u٩���pQ�>�ނ00E����������I��3Oh���ú���l�}�*�U$$���Eр$l$�N �L� ()~c$ �6��1�[�b��D�X@7{&-�@qs��r�#T �|P}�$dْ����b-�� vݦ�4r1�{;���& @�Q��Z�X�\u7Z����;�[X���XJ	#� ��pqJ�g����{j��>���#��컙�����S�qyqA�1�zX�{�����(#?#�˜��&
-��tF(&�u��#�W�����iv1�{%םu6Ħ����n;
��;&�5F8�ք�����c�`u46fC-���8���$/Bz��A�`�u�����F���d�5�zu���T!����f��n��dg �f0�Q�<f�㑞X8�<��Q���}<$v؂R:=�YlT /,���?��]�m��~o#ٍ9���,�<�al����&Y�Umm&���Ɨ�d7�1�'qݭ�9�����cz~&���w�+tM��$a^0yuAk2��5�~��k<�vߣ&����7���p��u�R��k���X#>���� N\Ò��T�dR�Qg�Ѻ�X�=	v_�{�g-���y��)�ݘ��.
��	a���I���^������M��+�O�8���)ٜ`�`����V,~�1Z���bv2?�����aX�]�����S��7�����P�:2nH�,]ĺ7&�b�0dt�Ny�p �"�{B��/��ʸ�� ��Թ�k��e{\��X<�����*��dh�A`��<�Ph��Vp��e�3���31=�"�w��u*��~�Ncʘ��A����7C�7B� �>���H�h0d/�ͷh�-KX�B���W��E��LCV #�3x�l���cP�7W���� �W�k�����	�_`>���5-GEtFe�\;�MvQ��?�{�8s�
{h� �p��^�N܉�tM��헜��s~��)\}��>��m� 5�/�\��N9�^���rq7Q���}0��6�ޤ�Y}0��u� ��}�^�}@#�V �b�6Ǆ �7~��[݈�I��M�'SE���߅5;02��1�<�����|��>�Kߞ#�1�)4�Q���ޅw��e�_��ݰJ��5-~����ِ�����(�k����RS�XH�:�on	�4 �o�D�x�3i�VS��PVu���#wX��g �0�quy�j�������l̮��[ч�Q���E�S8�M��n�s�\s��_r\V�lo�3v���-���)T_�=/�����8���𸹗���i����!<�(�b�T��|��^�u]~>���jTp��<���G�N�-`nk��7hB!.@���6;8ƿ���eʀ�J��3*�-Ǒ{����x)3���_�=���A��N��dY��������|/�M��+�0qi�3�����%ؤ��tc��������z�-���:���0-F"O�酐�@ZڄA� -����Xܭf�Z���qb�5ݱj#��hW#M(2P����A���&����+Y؆�kV���/;������ ��k@J�Ļ�{|��fJ�@ ;�¹�8���,�|wI��hOSx�����:w4�%�o��E�emlɶH	,�4������{����k���u�$ $�(r u�6��>��m�MYg�K�O�M����]��	����@!P�,�%�L�	����W� �����8
N�1��IoJ�#�K�����^c`�`]-��%�?k��2�=�������ҭB�p}&�Y�� �o�s�3��v���x�6���`(ر h)��c�a��%+Nŀ��[&��`(�۲�a0�c%�x�`�������2�%�Hj��<[�.���� ��=�;�3��c�V�����
��W�,���  ����؞�d@Xk#8�$�,��0��3i�v5��:�s ?�Q�:c&�r��=���:�:H]��m����N4Ak�F)�/��X�ڡ0�يB�������-f;d� �B�
�����y�p�M4:�b���5��UJ\p�v��@<�N���+xӨ����((OPx;��,���������[?�mOw��HҤ
9.5�h�,��S7D O��D��7���-�̈́?E�Ҟ����E�*���\jv��;�PMH���_sqw�w�f@��D\X��Ko��f���@H���Q��G��(
P^���������?]�u���Y�n��; yE�Y�zk�ڮ�ήw�"u�]#�AmVy�=�əV����Ӑ[��)���L>��;յ�vX<w����:�������)V�q�V��dzT�"��0w��˚s��ﬓ8d��7����>VԳ� �RS�V½����Ui�1���QR�?5 m�(��(�Fb�Y�`�qr�$K��^��(Vн�8h��9l�����P�����Jg��!�@��u6pf@�B��W�n#�A�<
��?G�Q8^�ɵm�ށ�͵� d�޷����a)�J����@�f����,}>46!�I&�t�&!�Y�9 ��}��,�f?1溱b<d3�GsѴk�pn�.�m\�a��Q50���`2�o;���m�q�;���Q����%�c_��!���$m�{܋rσLiвXٌ<�j����0ecj�����YM1#��!} ��зih�>8J9�ʅU�r ������~�G{FdT5br n�L�ypyHgN��,9�<5�B�t~~}�������t�"Q�������2�����"�Ň��#��#��|��� ��?J���5�[�Y�=��]W|���[����y�A��Ew��2��M�Nc��h��O�U9z���Α����҅����7�c�z�.cASّ]�QG������}��u�eu�L`E�����C����y'ْ)�!GE-p��c�� ��u�χ��@�i��}�8x{�5��=;��c��u������sا}��@+-��y4��3i�c	z�MOv3 L���W/��{ٳ��pvt��4��G��G�������R�6�:�6�k�*6(�u���%7�	<���[�eeǺ��\�z࣑Q���j�^�$󜊪O��3Y�Gh�5����V� nl�F�%>i�}��������a�G>�֑5��ɂ����]z �0	�&�1���o�聘,�6�A󢯤���D�A[Q�cm���(s�,�lڮ�S�P�t���%A��ZQj�
5>$|�'��!XWQ�� ��9;��I���>3J:%��u��� �\$?��ı���tp$��]T̵���G�u�FTLXR�@�;��j���f���kZ	IL��*����5N�� �N$k4>p����Nî���Sv݊[mk0���uc`Qk�����g��,aon��Ho�[���o��������}G w�u?M���qmb�[ss�l�}j�.��W,��]��`A}X��v���߈&L�1�D����r3��f�Y�t���~��h�1�}�D"Zw��Q�Q1o��1�3گ~��m!����Ɇ

��Z�N2�YU�֩T�K<�ϣ��3$�x�6;��6���@�G"jk�	_P�I?�
�d@���aT�u5krW��5�H��.`�Y��n�4�XW�[�eW�Q��s3#�8��Ѵ`o���x�b�]�\�n.�N6w�r���n|��� ��Ҩž3:��`�K�Fsnr'�3@�/Cr���	�8eO�o(��gE��txla=����D�7�xx��h�XJW���rZ�F���#,<�¬@��)��9=C8��C���X�%�1�u���#c��)�! Cl��3�L,6 ���,#]�`�IB����S�C�0� �*xy��_}y�p!w'�8��z$t����;ˠ(�t���\	�����t.M��?��!;�=���f���]�ﱖ��������$��G�K��E�w�w���4&QX aR�!�Â��T�h��������쑄�����88=�u�!��O.��q�e��h��Ĳ�5~�=�u�Fyef�������>'�ʶ��,�׃h��՛���4��#ݚ���:����Ngé6@��k�g�J&�Q��l�;���!p�bd1;1���SZ8������j�|�2�\ݶ7PX焳9�8������� �V�V���n:�����r;���t�U2U
9"�9 f0B�\�3��������m�b� |ۚCV��>;����0(bF��fY��he�_�*����������p\g�5*�1c18 �NƜ|Gg5������,�;�b+�p���cd5�
+��y儳��#���R �T��2[l*����e�En؎^Ǟ߸!���Ӧ�)�p�`��U�v� ��������G4�l }d'�E�����B�Vl��;����:P�qM���X�X'G��g~�:�C,���1&�\����G����r���F�p���Lo�AgE�'�y���w�j��D���#���9`��<M��3�b�5���X���
�ń�rK$�GAs�U�U���e���z��A0-��Lx�A8Lg���^3&��Cw��`� ��d�\��e$�
��s�b\^^_jl���'1+u���w�<������@�Ɨ��PWt�L��Ƽqvh"��`զ?�Tt]_
u�ԓ||����"���d���1���$Kp	5�jsw�)0��O0R��[,�yޤ�����@�.����:Q�am@r�����.�B dƹ΃�r{�&��m/;�%��ߌ�B}�PrT$�G��e��j�bK���� �m��AS�u�����;_��@+�Ѧ\Jjx�=���9i���;�W���@%3�\�*�U���C5���l4]B$hF��D��̰j�E�liKM���s��Q��*L�3�[�;�l�6��̝��|�~��޿}L*7Ǿ~&U?\����x�	n.X���?���H̊A�j��k9�@*�5N��BAY�T�c+�8��@�����&��DDms&���ol��߲�0w���
�W&,dv�1+��)�-�u7|H�ĺ��֣�'���"��Bq��������,R ܐޜ���6n�ݔ,�)�]�\�X�8�L������@��rz"��r��\N4W�Nw!9q�A {���c�6C'�2$$A`� x:�2�lk��ަ����õ��V�cH,DfrS��3�7�254unW�`7���~���FY�vb[h��U�E��՗�i��ְo�8^�9�#���9;�cw���Ӝ���ﻜLu6����:Y@���"[�!w������[�Х#��w�˝,�.M�F�z�2�SU�WoA������=i5N疺���\��ӯ��=�=����Q�0XP:8��`��p8@Y����Lp7��$$�;�;��7�IoYl�Һ:(��ag�}��C�g��F!���X����Q��o^����+]4 ��z���ANp��rc�{J�'(��A��S;~_	I�H#?_?���b��v<{Y)>�	E��g�Icn [j�e�w�)f�#��X	-T��\\b!;vz	�Fb�t\8tx t]_^Q(�������8��.m��gY���ݦ�w�N�av�F��I[+У�n\4زӨ�f���(�w_�h�﫻�[`���4�E���_�om�v�En48[�E�i��&tv�}l��t*&�
z��[��]^zYƮKsF
�A��^ $�]`�y9x���
�ݾ��ڎ���"�ҟ�o1vL�$�[�}����ߺ���+>z��O�L��h��E��Κ�F�/}����r������b\b��1�6��̜Y�g�������Ui��p�@���`&Hl������Q5]��x��ap�*F��|-���C�o�p� �)q� rٸi��M�ш��X��gg��{0]p�#�d[5�D���#Ni�@Μ#�r�3ڊ���g($9f�fGN9�7b�E6�T��OS� ������^��T\���0>�M&���|D�T���窱UR�~�l�z�&K�ܰ�wS���K��7^��v�-`�� ;	������ݯX��,���L�,��I���1�Y�2w�C^SbTa �0�A,�k��&�����0nSf��or�����+Q�*5ܪ�c٦��.s?����Bo���6����A��\��>ޏ^k�2-���@]�G���yxv�����[ω��@c��0�e�m�>;�w*�?_^P4�çO�����;3���g�p�t4�8H zTTGc�p�#�)��ÌyTe�Y� ꚮ�-X���X�� :L��hQ�׌7U�(��|��7%���Fo�Fg��8�|�����`��r:�q�����~b1�E�hu�f���'�]�������+2�=?CF]Ϙ���Z@�`	uj"�L`?�hĜ|�Sڝͪ�ϬR>\�2�=�;��h�5�O�^�M�����NM�\ǒ1a8[3� ��kt2�gؙ-�'�Y#��}�^�T��ۊ���i�ly��p��y�O�T }8�	7��� �DF��P)��T���듐��+d\g�=O~o��S�1����Ā'<vN�;�g��m9����gP��p���߱{7d�J[�����	�
�%�[�2������8P�����T@�3Υ &���R��6�Ԡ-UV�{��X_�x`Z�͗$�@�i�F��g�5���&n�q����"�5S�4|��?}��Mp�QG�V��9�P��)/�̘�t���T�٢�P��=ɪ��ƽ�����^�ɩ<<�(F"�2�G�:+�H���@43g�@W��t)�Cx���J Oڔ�������q�n��B1��[P~WЀ�2UҦ=H���؜:6Bb;�ܟ?|w�7��H�`�E�L�RAׁu:��)�F�<��u�ƹ��2RMeb�;-����5��-'����T�����A���\�F�^��싗/�ٳga�+{6� �;Z��2�h4��\:��>�� u��E�ǂ�vǊذ"u/MZ^n�yK��z �٘�ؚ�` =��� ��o�Q�A��
����G��#�^8�ر�{�1�������u9<@"�?��֧�&�*'������8t��{�|#����Aلz'A���b��bI�9������5�����(� ��H�	N�nc0+�Ӕ@Qh�ڎ�6�Fp�!P��iJ�k���a��b���D�-�5t����C�+���Ɍ����O����:�{��j;<q8>��@���dօ0J���r�����}�n$�9�8�@}�׎�^Չ���g�0�������`�k�@9V��K��M�0.�~�Ct���I0�1l\'�(��L:s0i'g�0���)�6�U*� H�=;�g'd����KE�t��lP(>�I�	�C?�d�ԉP�P�u7�V�h���"��b�_O��7��wt\!�U$�����!�D��`(48�K�R��ޚ!�,���bG�������)`R������n^�=���QE�}K�;��o������V��tR��17K��b�1�4��[���1�]^���w3�F�����j1�Ώ�0�'�6�ߦ3J#�^�	��mpk��`����ۙ�����'����7��y�(F���Xf�1�#���9΄&϶�9p�Ok� `7�y�yz,�R����"l���"�O��_�;��0�9��|�:'߈����`����`b#L�
�L� '##����3�*S�����[P#���jc�b,���9�ka�A��c.�B����c���]gt����q'��`M��)5/'Y7����w�ہ3��`m�t�1|��6�BZT�&��ȇ�E�����?¨��M�<�mt��]	�B����4�1WL�q���EN�f��v�֔��Z#�� ��S��qj�a�_��s�5KZJaN�Z4�g���z����9�S��L�l䙋�/-�����q�����/�k<���6@�t��28ˣ1�;�E����:|��밟r�%6g̽��@�k���n��s��ݑ�agS�u2+ � Q]t걶;�<�#|h8�QjZ9�=�tgh͝�Գ��h�=���q;��ia_�`j\\^���:��!|�����F�!���E�,�JL{{| +#k��և3,����6���{�g�=�X��B&�5���)�-�\\v�s��ܤ�?{����qR�)�=�#s��I���D�}��Λ~ĢG�9]��`%B㫰.�rw��w)}V-��0�����1�7�K����|9�:{��~5R�]��Б|�T����k����#�� 0ȌJ�2 �W�k2��:]o�b��im�&}gG�H���Thl� 3�OO�h>�K�58L��6��s�ܑ_�O��ћd�!��k6.�u�"��g9N��ic����i���=��$F�!��
�����'���O2�wnx�=)mQM�p����v!8���N)ײ�t���!��I�z#'60�����	HD? t��}b}�)!�6���d�?�h����]õ�^\�=��g��ΦBFD��h���Y��Ū�/
}^%醦�(с�^ã��prpf�4��S1���JH��~�U<5�.���xCm��3%���S/���U@g�]t��Ɩ�F� (�Aq�yI$6ʵ]��� �0��֭u���cp��*.r�D�רPK篊]�h��n
>���i�=2I��$�{{�.&P�F���,(��`	y+&T��Ryܘ���No� ��i���bi� W�_������҆�tK�O���B��t�y\" � 0�3�:,,8�`�9C��k�6Aڵ�Me��H0�[��D�>��=�Y8C��xҬ���!�/Zr�D�%3������1ē��b �ϔ�Є����v#fH~�0tl�9�I��-�џ�F�s�T�I4�1|�>
O?ߠ�� �(��G��Q�������Y/
�I����A\��B���"{Ċ:� j찓�]�!�x��	@(���(,��.(�ǇG�`�!x�5���2f���N�Je�11B���!�I?�wW�����S7�����5�$n�s�2J��	��ۑ]�'ƃ��Z0�Ӏx���h&�T�,#upW_t��{[�t�ۄeZ#;)I��<�`����S���)�3.�zc@�9��BBA���5e��^�}�����,���}�?`�	#Tw%��-��PQ�;�ׂbo>��<�́j2S����^^2n�:����"�υ��u�F�f�v���E1��g�#Y��w7�A���u�Ɣ�/wҨőwi���Җ�9�FɋJ����[��
�~��P!�ےׁ��3\okh{)������!9�.4 R�T̉�ta��D�?��bJ�%a�[�Ҏ�+�,�4�:t�P��;���'1P���w���[*��g�G�l�$�Oy�s���G 1΁ݾ�N1���v|}T}���hlW�n���x�ft���f'���F� ���Z|��EHj�\&�`�,&B�N���)x� ����xla�g��5�8�PL���c6�>�m�M��u6,���mК � ���4��<r,g�`�1�u6ƊҚ�~�
��B܁f�VL��W��w~>�5xtx�#G�}�_M���g���}�6�O�z*-��Ԉ'���>}�d���8j���E��3�� N�dm�5�%�m)vZ����9;�a4Bl�֣i��pO�NLݦ��A���iM}������S+��� �|�P�Fk3���:$m�N^C���(���F����5��T�Q4ε��Es���1��u(2���}?����C3k�#�����g�� �B���-p�i�=a��#[����S�>����[6=!�p��Q0�Ϩ)��L�3�&#`�#o�D#�9S7�ɗq`K��K9bH�>ca4��a��>'>���)Y�d+�^n��k��	~�o�t<����3)$��Li:	J�f|��-�#m�����K�-��F.Vcm7?,�tv;uKL'l$�Lȳ�&���}����8I��d�|~c$��0�/rK�`������B&��m�<܅u�Q.a�hjM*w�z��Z+��<.�b�?�u��F��)@4�
M� �8ľ�ÿ0���J�;����w��[���_	$N2�y�g����������
V��G�bhYM�\��0 :�,�<n�s��'��qFs#s��ٍ��ý����yxy��������s���c�7�cw���z�$�]Z�\Z���nge.��/`�رO�Ti�V����=�Р6�`}�iK �#���I���RW`!�^���� l��iz�ݔS�i�c34f��u�֨��������\�����%E3&Ά������2@M&�p|t~z�c8=<'�a�N�aQ�Eԗ�7��E͢ ���F� }| �(�^��z�<S�=y���Z2ScppL��֝t�-��� �1��McT��,���ﻻ[ki�^|��3K,~fPƜ�r!��ii�Fo�e������¨S�������]��)�^���o���Zpk��r��u)�
�~Ŷ��]AJ�%vP�*��'�0Qґ�t^��B������p��x����#�r�_�Ͼ{n�� �����������?|����8p]a�0����ӈOъ�Z�(BoB�:�D'�V��<P�%�\ZG<rS-��"�T�7a��63�Q�i��Y�&ɤ���~cb"���(7+[���?c�JZ��;�4�� 
zs4GIև�D�NCg�ꬰ �(�i4���[��퇂g�]�\%~#q���0�-�(��S�����4�'h5^�;�����7�o�Ý� "�\�"S?)�ΑϞ��@�q��m�)���?��?��''�㷙W���0�Zo�V����c`<8<
��{��Rb��%˽%��֛�HV0v��0;.۩��6��rl�9�lrD�#�:d>vF1KK��s,�&O[�q�L��(��,��}���9�t�>0�:;�	��&�{$��i,�|��9�{V��v�&�R֭��.���:�I	R��j��I:���N1n�CZ�>>]\��t�h-��e���9Ӓ�:��ٹg
`��q-@(�`�ǳ@��� �LQ@� �I	+���Y��	� ��Ye���"�RU�s�1W��o��מj����I��n����i���ߙ��@�o�:4V���9H�O�&�VZ�x�����t�DH/ba�QD���<�mK���}}�FA0����@�-�d�(d1��Z�	�,S񻳷��:��Q����}l��q�ǓRqB��m@�����^@(L��@}�b�
. *��	�*�hE��Meo#�l�x7���vҋJ�Ba$ȫ�*�����x&%+tj��yq�L#7m��N��ƅ��]�Z���:���?���(0y�.1��&�Њ���=�	m-5���%P C� kz5��s���ٱpkD��j�JX��:|�����I�BL
���~�>1��ײ�:^��@�0�F�mD�q 1mpM��5�BP}.��  {��l%c ]+���.\h���Mk�`������b�Bn��B�Լ c�,�w�5�6`�?��A6�ޯ����(-�l����>�+�dFִ.y�N�����v-�wS�W.*�N��6����9�3��$���3��@�AsN ]�1_v���%
�� �lO 9���Pu�=���qK+{9 ��l.W�kJqbg�K��;��v�r��Rb>�٘�y���oi�LCzf�� r}�ބ�ƒ޽{�5\����Ӧ��X��M/g���Y������ɖ#�ie�egt (�0b�.�=��\L#�4�x~<i�S�W�`��kF! ذf=G���V:}3嘍F��|�B���i���/���w|�p�"H���
f��K1�����m�]��P���-��;O��ٳ��?�)�x�"�1����X��;pXt����B��)��0 �����%ž��?�?��7GV2ݚ	k	6��.KPӧ��ׁ�+J엋T3���'��x9��!�7�4�xY����������͂�A��_��&�o޼	��7��t�>^m���8W�F���F�摹-����� #_� �*�g)� W�~���fe9�@���鳬��aDNM�O?�������9�vǲ�b}�H�@Ns�o>�VD��2W����y4I��)_]^��W������ȥ�jJ� uM/��9�,α/���_}O�_߿o~��l��/�k�"�y�x70��I��#��ju1ݾ��������PMt�5o�z:9>�N�3K����!��n�r�#���Bj��b�cQd��5�F���'�b{���7��h��PuWQ� 8�����+�*:N��z��5B�
�?�������t�H5���Y�V/&3'��1�䁝��F�~0W\HT��<$��c���#!��+�8d����;�cy�3.�ł�6
3{�87�Rap�J+��p�{�
���[ru��6���&$����Sz�`��V�ˏ�

���%w쇴�*�/DKkZ@�zt��P>���׿���旴�o9n�ō �`��gϞq�(�w<�t]�4-��U��٩R��y��0<��2��F���1%A8�$f�L��.���04ڜp�n�)7Z̭%��*�*���)Ѷd���E
Hr���g�d��%�(�	���qq����з)��ɢ3�Z��ƍh��b�� �:�b�A�yt�r����"8�\� GG'}�sc��1��:6�hU����I^;���BA4��\M�"��p�%�:��iђa|�`	���j���E�3�#Bg]P��N�1�l�Y�?1���o۝�L�Լ��k�!��������g�NXn�ϣ}���n�k�����Ci�.�3�X������
��o���:9��>�}���y��	n��c� :�`@ғJ��V�`c'�lm�$�`���F��5Z��s�6LbJ��l��ĭ>���Y#	��_o]Z���)5�c�0-�LY��oI�����`�:Ž��%�E7�2���Px`����ڼV
+��i38��%jsx'!��1�\���#
�R���?�?W�X�����}���#� �b���#G���mA�(4�'G����Ã3��_|��]:�|�ua5�C��~E�yh�1��j>���XN��OQ?0ƬS��`i�r�b��X�$FT�Q2QS��[q�=�$k�jk�b݆�g.�o�}.�\�����0V�z��bK��?�T$�(����}0�At����?��{dD�>��ѥ&�<��*4�ҽ��	^k	 ��Qx�^V�gC�_�}� ��[ �ц�O�S2�|w���N����F��#�0t彳�{��"Ѧ���Q)Z�t
��Ot������uȣ%��q�LJ{jR�ˊ}�{v���q���)�+$:�)~�g�&Q����s�iy��`Z-��1m����EQ��oV0��;���JcN~�~*���,!xZ��MI�T5�3[y={���������9D�̊�u������
0t!����^XL4�d�IxJ���?��,(V������޽M߷��֙!I���,�(����7���ݽ��Tt[��9>�� ��y��uuC�=8[�{���|�7�xX�X��i ��`n�7z^}a�2{N������%u/�QԙfM4�e'VcU\�9)�A�z ���s�%�Y1�n{����Q�`|A6<F7�F�^��G!���EO%s-���S���X��³u������@���F����zXQ�����a},��!���}��	��x�7���6��S���R��lYn����8�5����O/F��(�Q$a���/�rE��g�Y~־�l@��k	�~�k C�?���<���tm��v=��$P�ll�*sÈL1˹������SQ�*������~ާ��3vm�h v��Ux<.l�N{i�c=?��c8;?�X;G��o��Wӱ�\�P�Z Q#��G頙�-�,q��3���.�g|�^q����� ��G��/����X���ޟ����.�/�I<�c?�}$L��̠֨_�@mkM�&���� H���4p���΃�O	�`̉�x�&)����p����?|�J�sw������0�ҝ�أ�t2Ayg��Z�8~�F7G�k垨�/>]и�o�ބ7��X�)�yH���kĭ�~�Ć�c�,>D��~
?��S���  +�?�	�P}p�2�� ��~i��vN�P��a<��}�?���2�)MCIN�i��|7�z�"�������Wa�g�o(,�p��Vr�����!�Vwnel��_8a��h�KvY�.�=�:��[|�$�@�`k1�F��{r-	�5�n�Ǵn޿�@wŞ��
h�a\�eL+`zE�0a d�#�����O�ytt8!0�����K��d���t���J�j���>䋦6�[�Ju�W�@�i��Ns�<�0�� �Ś������*]�������UJ�t��ý�prt�n؜"?�U�E9��h�Ĝ��|ѣ��BK��LIw�`g?�|��:�F������	�M5��� n��W�EW��]3h�Lf]���Fu'� �2�
u ;���0��tȌ�
�&��?�ԑQ��?���~���<�{ǣ��ýuf�7�z)�#iD�u}��H�BOʌ�:��qY���msa0^p�=X�4QPt��8a�%�^��@G�&�w��2T?��xx���ʱ�pr*jF��x�7Y��aJ:�t�G�x�Vf����I8���6�$��q0}6^���T�������&����!� ��}�ou�lw>������v�b���K�^[ש7z�D#���ș)�������b��}0J�����N�-j�=�g@��D������_ߦ��ܨ$��["�ώs����~��j�Hh޿�@�7��e�C��D�K	K��Il7F��bD�y�b����>=>aמ	q
�o��ʽ�F�taH����*�|�8z2�(�����d�e	�ܽYmn6MxhWa�>,��yP�H�#C��ThӀ�R�%�^�4Y���[�� ��_�-b+����w���5����z)�
������H����v���8��x�ʁ����H f�b�)��AlX�eZ2�DQ�q��ćm�	��c7p�C�� �E�lm<V�?���J�}��O���k端8��D5�C1�8�\���o[/������=E��E�b"�5m{���O(Ra�b�߈�\U��B�� ��`Ike�v��d/` �#ٟoG��H��@rw%,�!��Tn�����d��E�uĬV��TG�}׏B���[ʾ}�;���ٸ�rp]�*�:;r�K���&&d�3(�~��h�RнVa�M�D�NŮ��������ȍ9n��^Er'��P�ɱ�����h|v[!j�ލ�υo;�`������JAj�4��ֻ�\�ۦx�ϟs���oS�g�Mi/C[��x?�~�}x����/8 �4�"��=��-���Av�.�
;�|�φs�Im�f�N��Zo��=��F���}�_qT����&\����C�@;�M�K�n���uZp���-}c��uj���_���- �G�`A�F0�&�_�����drk�Q���>k���s�E�`���{Lk6�&�W�n����>k�EfR�b�6^L�T3�n�	�}Cv���i{��ؑ$I0@JʧJ���p�����N�t��dJ qaf�H>VuO�nVg��Lf!<����]Kp4�,9�dޤd>��_ �ɀ��fC�7��aEaJ0$s�ui�#�1*9���~V2H���^b,~����=��ϵ�<��������c�����z��dK9�JY��LEZ@���q�-��4eH��(�'�qwC-;vE<��Dr?M�(��ie�'�	f@�XbLPR�A���e�j��Z�7�y�I�I�v�M%aٙ��qJ�G��Z)
�yc��cO2r�a�K�%�%�2ѹ� >w���@���Y��$�����!�F��E�%FkC ��S����]���v���$b��<	�j���9�@�[+��JkǱ�b����2 ��uPJIb6R�k��ND�[k�f3�Ye���L��e#xd�����m��~���5cy/�pF����Pl�I�<���= ���]({3Ě��Sk�e(�X�Z��m���b� l�3<�l& ��7������G&�qN�т_��p���Bd�PH\1��ݝJ��߸�"�x�����.T��M�~Op0��1����;Z��ޤf�CŢs0�G��-�������)o��]���w3b�UWN'���F�s���va�č]]�I@g��̣u}
��mQ�׷��:�(�\��@�t&�,�
ͭۊ��C�i�P��OρT�~�؟�I�<��!x�H�^��E�l����0�uQ�c�� ;�fY * h�"}Y�Cv�{�x�/֠��Ϲ���z�A׈��(x�}��A� X�֯e��mW�nT����l!�Qᄐ'�8���Z�Qei�`�Ǘִ�8*=V���L:��3g��FM�h:*���\�jԫ#��8���`L*�/}q<��+����,4��$}�����̰�8&R�ݢ*�(Y�v�V�{$�5b�δ��L[���8�L�&ưRuYuſ�`hl�����!�Ȣ�@��P���ՠ4� ��iC������[�B��S藎��|�f�3�=P�Y�/�|_>	_�}�&  �z�:T����^ �`-�l��ɇ)��|AY��t������bg�qo�Z��n �d��C�Ç�0����갦"�5K(���̗�}�#���w>(�bPơ���Y�t��:{���֟�'?K6��wB������ASl��X+�:g�ֹ2=������]�����
k�PI�b̍l�J,Z�8\ �~��f��/����#m&�*8G�xA��h]�,S�W��لN�\�,�uG�~Ap���Fe~s��4dF#t�F�3��#5����<�Q9�������X(*��\��<��@�d��r`
�\É匭��n� �ke%�Pf��zcE��;�@f��pQgI���[fG}���'Je����l-1Ӹ5�F����`� �p`�w4}�΂ �͐&��wq���,��ضP����	p���E��0��S��N9�xvM��](���9�	>��~��`��k�y9xk�c�)�ٹ�Ub���cHqy�p/	I\��LN����� ���C[���g��I0'N��<8\Tƙ�ifB�Xk��X�Ӹ�>���s��O��8��?�!���?��>�H��£���G`�A�N�=�(��T�n.|�Xܛ�ؗ�(���Zc�#��,�e���3;�����种�.Ԫ=� �Q�|(�bӱ7� ��+-��ִ��w��I��
���a\�Z��6:�f�>�Q:sG��~����������T�2%���WM���,K����EjRr������+؁g�����j'%�^s�cj��k9����bMMܟ2���	$c͵�]�X�7��`��`%���|��b-�\�':�=9�Qm����y���������+X4�Ǌ&�D����C��!��5Ol���$C���ӳL���E��\�鴲��`p`��|@ ̕`�)���dʢ<L�q(�s�r>נ�xu�]󓠥%%������&��h��X��?�|씼g�b��mOC�������gI=[?�T�1���}���~�آ3,��b�|��4G�lwЀ���3!|h.v�����z޽7.Qy��km�Y�'���C�zI�|%%.��#dnZƹlɎ2U��si�Q��h�M�!�I�"q�S����a�d��#����>�q~6�ޅ�KVʬa��P)F���sU�^O����<w�@���am�ѣjke�=f�|q�&4aj�&���;'�c�9��w�{�%1���p��ԕ>A�;ļ��ڄoN"�%3Y��?n�v&�ف��(K륁V����}�_�A��`��6̎8S�d�߅O����U8E7���ںq��hJ5��۪�b�:ח��C>��`��}5ʰ�٩�� Bq&S���zz`�j� ~�����C�-Vwja��ۍ݄6'U@Ap6�Y�x�X�Bl��t0q�yp�_ޱV3Y6��Q`&/CR'^�8f��d�p�0L�ƨ~�i��� ,|�N�R'�b4Ǝ�:�S)����s���fSO�J�N4������`��{��Y֧���6
��#�<H���;��Zչ�=���B��l	�vM��)�&�ر
��`u�<H=۷Kx�hY�b��|
W� ���M��!������$>&3k������fǽ�/�Ji��e�0�1���8� �����
'H*��R�%0�Ms���
�"XB��"���Ѓ6E>Q���,�s����p �q>�i4�qG���e��`�f� i�T��kFk�'N��R�� ��
��)�c�ʝ���i0�{���R
�oeɚ���5�Ƒb� r��:[ϛ��6g1���	-Kc��n#���O�@�F2`vy�*[�,��lI{�8��Eh�?��{/����j�5�>c�Ւ�Sd�Fs�W˙�q�pyy�xO�^!��-K\щ8����)4$�S�Nr�7(:����#�]��\�Y��멟v0���_�E|�6�I�c��t�]l1x` Kס�DK�L$�j����H�k�U�d�����fGZ���@g"�u�a'e�����f�Q	�W�p����ÐJPm)�tn 6�,R�Qc]����7���6�]�<Yg>�,�	;hU$���>oY�)���ksU ��=cz�|i���:ͧjk�a�x��E$3α��^�U��q���Xk�d ��}� �	���T�������`Yjc��bvqZ�B�'󖪀�wnA@-8�X�0�3���K"�!H�s4 	�_kkg[����>,P��8��B�ဢ,ɓ��'��͋�:� 4on]+��t-�����JtvOJ�aG��'����Ղ�%kJ�ٞ���Aq`�ՖP�!�
���K�kY�B��*�Ŏxy4P@"��aG�� ae;?bӖ�v��b09���?ɷ���<*����K~�q.{e_�Zv�i�vЅf�۬�1��3��eq��0K��e+��O���y/h*��׎y�l8��$��+�a�c�N�H_ϱ�u�6K@eJ�:?����'����{�И,aKI��AO��o�ņ��CIzz�X�-r�x䠕ʀf��(�Z2x�;����P��~g�z'0��6�S�u�l&�����X>��A+�K�v?H�e��|O$lPn��I��̒G+�k���t�y�C]��K�8�Z/su�+m�Yjkl���1Բ1�͎���`�G�pdY��7v�v|L ���c~N��ܔ�l,��ؓL �|Lx��<4��e$_8��YJ�Oǵ�!Y=SW���%w���b"���_Ca:��c�'V��oln�p�ܥĸ	l0����A��j���+�n�Qk���Q�3��<�R���Χ)��2W��1��۾�S�h���6��bX���:Kg��/�Q��l�t �������:2{w;��`��M�I��:�Ϛ�U<Z�%�ðd�j��0�����P�:�_�߇�~��j�lY�B0ֻ�"y�R,ZZ��5���q�Z���$����\��v�����H%qҡ�׺]gWP�	m�P+���;Z�;��8���2�4 [���o`�&��yWn_�Qy����.9���8�x-��	��6���1�o<��C �i���0G+�4��筮S2��_Q��L�[`v�`G�Q���B���ԑ}-,��r�04h�
Jz��
�ܒM�㍧Sf����2�A���GT6ʀ�.[x�1<&sB�*�c�s[�̙�$ӳ��`���	���:�,�nˈ����c��o4��F���NH��,����1�kՔ����U���v���E��8ݤW6j�7=p�a��K�@��-�q�@u������5�^���J"a1�8��Zl86�j��b���=P�N��2�����PCY��<������kA��!<�lк���7ظ@d���Q�d9�O�g�ޔ̒�����i(``�M$���C�1���I�������)�<�("sSA����C��ۻ[f��OO�3=�#A�o�y���T���ڸ�WY�/�Sm��d�	����{ݰC��b�狰̶{��g,��fO{ [����b#���g+��Ń�B ����b����:����Q: ���M���WR\)�Ϧ��J�-�ʣ�`i$15���F����G�yA�f
��Ꜽ�=R��X���gH��	��=eA;��JE���5k�d:� :u�]c�<X7����.�C���0�+1���܄����!l��{Ŕ(H��Z
��g,�կ���x�M[D|y& ��j9HLkV� ��6~,���J�����N�)�@;^u0aR�9�_�5<P;�Q�q��m3��X�ٻ`	�ƴv�J%�K�M*�?Gk��y��	<�Oʊ7�/1�53�j��8�*���g��4���@�~MQ���," � �0�T[�{�l�Au�߉e.L/q��G��	i6�&����p�r-�NM+]�V!�o�p4�gS��r��i����yh�Be=��:��Y�|���{y5��3A-h�`-����MOJ�j�M��:�Ρ�!Pǁ%�x/�G�Tf����k��>�j_������K&D10���M������8ۯ4!U"u`�T�c*��zc��T/��C�K�
Ѻ͕D���3œb��c��w�>X�Q�M��(%g)F�.�띘--�Ew\��Q`�Ԭc�/_�� L���vL?���_�O�a� � |���ԭ�H�
bC�g��+���y"�Ql�A���
�ɼ]{a���j����N*�������-��M�=L�>���A;������Dm%c
H�n)mA+CM6�G��Ƅ`���e����sY�6��R�����ͪB�m͂��W�
���ˮ��a�P|xW�����7 ��[��A��[F@p*�`	��\����w�SG�9}��Q��$\��笔k#Ւ.��%���n���z���\zY,K
*�kM8z�Y��0����+����_^�:���v�[���w�X�u5n�;n�g��aމ��'D_��u�T�����>�c�%����$*��ި�3���6��Wu������_9�֘����?~�L���x�O����6z#�z�����G<���w���@�gU'j8}�O�o��?�5�/�y&3Q�R�ل�P�*h�}"�ӵ�!C+2�½�_/V(Ś������pPq�#P�
�w���g9�B���~�Tt5Vg�����6����p@Dȟ�s p�h�5����
(n�|�>��C��0�/!����,=��׳5*�	�/�^�D�#�����0�@�!��D�wH���n��o�P�$Gς�^�L�N�j�G39;9�4^�N�9{��g4`�e�@�oތ(�Ai�g=q b���u�h�
�ݮ�r�^�-Oϥ[Z��b�:8����J�ԪKK�G-�v8�O��D)!P�y���]���꫖����e�;>��\tN��4-�QC�x���*�bxB�L�5�uؿ�_%���&w6�����ךgtk�޵����ZC��Pܫ�QK�%�J#K�@�G�
�N([�����E�/Ʃt0�n����1����ׁp��S=�#��-�&ۃ�'��/�r����?y=}���_tp`9�Q�?����G�Wj��N\=���xWF��]66�S��(�� bv{��6����U����Ai�xF?N�A5梽�g��x�i�<���մ��CG��:4`�dg��Y]7 @�k�Y�|]��F��?�� S �Y��+0��M����C��{_�ݰ壺.Ymξ[3�N����@�"�Țp��]��������E>?Zt1-���t��g�@h��M��o���L�ׯ�2x�	
8Yf����U�����7.Vv���"U̜��p�ײ��_�J�v,��� X�I�Q&@�L�3MtLA����F©���*?�Uv
�.����A'\;������	�q���V��5���X%ad3��U����*��#�I�3O�����1�k-i�yqL*���T�� ��n+�}&>u>�M:���κ��6�4K� $g�՛<�è��ⴖ�ţ�qyW����̂�SV��'�3�5p�׸J�0����O��;���Zz{����a�|f�7ڤ��~	�n�~���^�f�l����Mڐy�s�$�+:h��b�ُ�}um��=�]M�~����U1��(�K�#"���;Ȃ�,9�в��ؤ�q��q��k���:6��=�ݬ�^�5���k7�ĴD�O'k���$Yb��\K�K�S��.��p��1��.j
�	���T�V�9;姍��Lod��y�2
S4�߻&Ic>��޾�݇�]Y�~���o�:+��-�(Mp�:�5T��j}Tྔc�=�勞7+���o�։��;��@l�+t��͹�0g�Ȇ�%Y����K���e�\�s����۰Kq�� �-[��+��G��p����+0m���u�V�Ίnߴ�|S�?H`�}��}n�g03���a4]��� �A]�,,�����i�,� ��f�I�xHr�e_���p��C^��W����Ebɓ� ]p P>���+���$]+��Z.b�NKa��8�r���^�O�;�����`PEv_��K\Eʉ@D�(ٍ�S�����kU�%L�4�;�����k�,��������cXe��رu��IW��:3	dp���?�)�����_X	��y`X�i��`l)	<�X�M���>�#7����Q�˜��g�u�p�yG;��V�	mK��h�������'0m��2BP'IT�����ty� ������U9��RpqZ��_�o�v��!��6��lO^";$�#��H����j�[ b�Jt������Bl_R���0�A�%���Q@dto��y�{��n.x�*1
��(|N�u^���g
jEk?�:D��݁zht�b��0 :��çp}�.OƢ�q��Le�NxD��xi��G[�Wܤz[�hFv�hI;��x��@@�%�O/�B+�"{�ﻱ���ʚaV�����竳��ϹY�(�7��F��B(�X*�\r�2�_L���5��3�Ƌn�C0Q]9��\[x	u�����k�p����LJcG�؜8�8H�)c�4����ʖ�+���pT�0��%)���a��iP��u�w�<�E��Q�E3m�A-͓���2(�#��k'�]����W0�9�1�]��It��Юւ
"B��̍�.wH|�:+���қӵ�[����X��������C�b,��YK�ڝT�o�İW�^7����pAG$�ģ�A&�6R�Ɓ���I'��V��̫�\"�l���I!�AA��I�FбM�ń�)�ۘ���rLNن�Q�����"�<������������c��k����������q��Ƒ%|�͹�&��>M�Sb��X��%s0;��J��K��B�Q�uv�y>��������� L�"�����\s6	���<�,N" �����K��w��� 5�DA]e,��nsB�%8�h���@��hF��k˟y�h��j��]�_$��y7�|8 *�H�7OA��w޴�o<�Y�,��Mj��?� ���n����������Е���Q��sD�u^�nuP�����؁����N�1g`�̌��6���[%Uƅ��k�+�㚝�6���0Z�;
��.z���a����X����`1����ϸx
��Ը��ҬE �NS�	WJ<��^]6�qt�a��a�
��� ;{�X�(;��*�Q	��w�{ꙴ�,)�J/Z˖5t,����'y�"��:P�*�������˃�Z�z:Y�|��;�����6��%���M����=���ޅ�Oŋ!��ۆ�ŽI�1�,4>���=ܘ&�㞕�ܰT�n/o��	6#�2�p�M��>���9%E��Q���њy�w�JD��]�6X���2[�m5v��$L6���%�1�5�F��7@�i�X���6��V`Gv��&A#�68[_r�ۙ�J�3Xj<Ú�ٚ�lm*�Ź��D��M6��ӟ����xWLv�tm�c[���}��}V�'��C�݌by	�`̹i��L��}�WC<��������j����m��L&:�T��5���o�#��Z���+~��b�-�$k
I���V�@��x�0qG���[@/v� �ii�t~F��J����Vt�� �ʦՙ��}4���s �Eww���}B���OƂ�e��G�?�[}�vR�d��M�&��-��:��c����gɤ	�<�}K1`�����C�)A����]����Q��k���z��T~>eK��@�*_�>D�Q������C��@/%�ޏ-O�߼_q� � ��}�i�b<��˩f"���_y�A���yM=�p�/�d~x�����%@o��d-#�q&��\L���?��/������nk�Np�A:��dg�hk�2['~�����WS�u��z��8`5�l�� � � �km]:�@*�gߌ�ӶW��
k� �O���W���}]��:���˕�K&K>@�9��v��c�{|�E��ѐ��5��e�U0^�m˲]1IE �1q娎��"�
ݮh$ry�$d���bK���U�G0�������ԁ'��^m(G�uU!0�IĆ$m������Gv���7I�/�m�"��_�#�|E���ph$x�v��)b�f�A�x�DMw�?~�[���&'6"C�gC5[�(⽼SNc�> @-�+���%j�Q�r@ Vb�b<���U��_��l�w��t��M�k�;d��o8u�N@�,�45����{0k8����e/a�`�]w�Qr-��e;րB,�c �(�CG��o3�1��ۂ�<���.rZ��vq�H����89���Si�Ψ�P2Z���-C!�ݙu�q]g�����X��hl�=���O�����.�6��*�xCH\���N�U#q�����g�Md ��0o
�à0�.
 v��/��u$�ҐG~>��˨�����-~������6��o+���u����ZI �HgN��!�>^O��Z�M+��a8:.��p ��"(���� 
�T��5�Y<�P�t��ֽ̻�N3w��2�:G9L�y߸�և>[�{6"3]�Լj�x���;#'{^�!.y�Q4Q<�cʿX�!����,�72c��Ǉm$�D��z6ǽe���9 ĮX!����Ͻ����܄_�s�ݳ|��I �u���'��X�� pku�ˀ�r0�z��.�sl3oF�g��A-g+���X"T�ǩ���t|������R�^���]����l��κc,��.�L�|���]��,tPݕ3��[�0z���4O�b�v�����Z��lN'������#�����%����
(���i5o,�2��Ekμ� �\�1?[�X���#˳�1����؇G%IZ�ʱ��,~���8Nt�0V��KM(���0k�z6%�
 ؟5��s����t%���k@�9��蠌:y���{��d��bOu�o `�6#����w�$��d�-`Z����>=���"�<!Ê��q�l�r�@=��քo���u�%���`�/mpQ�)�6\j,�����5�v�˂�����~�
�ߞh?����l�`��酺6�Z��
:�\��6�E�]�́e��'�q�"� ��U8��䃁���y�n�77�([������Ѳ��͉�Z	�@���d�6� GR��9��dj�����auq�U����'׺ke}����y�$���#iu�ϋl-`�g.��zڧ�}ޗ�I�C |jR�Kf�&J�?k�3c�"(��<���kq�`�/B*��S���m X䟖sX	�b��� �H�!�d0��&k�l%l�~�y������v�Hj��l�L���d��^W��*%����fx)�����CUo�O޾�Zd���U8?�[��4��7̘����L�B��J�p���Tg1��I*%.�ޔ�8���C6�ʼ �����O?r���e���=h������7���cp��L�D�6;&Yj�,q� |����w6�̒dX����'����s����?��|���&(�X���6�!朝��Ewd$�`#�����M2�
�B���2�P�Kc�CM�g��A��Yfy����Ɯ����������k�G7�%��v4@���0�n���?�� @����4\;��W�Cz��52��DiN�N��g{�����^�-��_�Z���whz�MLs+��:�-��FI X� �(�cN�֩uG�����K�F˼\���c�K��Q��I51'u���-�hX�7i��8��"�	�t	&�-���h%���s��ڎl�}�H�J���ֹ�>g*6�P���E�xT�	7����Y��� ��N>��y�Q̀5���x ��1�</t����d-�E^���\Z	��f��
���q�z�g�TFcD�	ś�X��xAp*�F[�Vu�)-��b�b���&��yg"c�M6�M���/����Aj��MVq�(�bT�u*\Hd�f�yx|y
Ϗl�r��M�!��ﱑ8�h#�v��R\�h$V&�z�`�1�h��]�d<b,S�����꼺����;����ܩ�~���N�� ����9H�{:MLŒ1�^���� ��&��*�e8f���ۣ�dC���-�F�aG�R��[�g��H���Z��m��]���
�=�����0�=���|�B�΢���K�]�\}��"̞�����3���{e�zj<��B��n���*+��ف��$8Ȋ2D�nj���E���?8 �v%�&�j+�#��HW���lTy܄o`	��3ԭ��	���a�i�դ��)���r� CÎ1o��,��\D0Ʋ~���õ��}�X���0(�w�gu�k��S�%���	(�Õ*7����ѻ,���M��j�=�f�g;SgRr�����D�k�g2D-n-Î$��l3��X�y���!�X��J��큩�dt�B��Mv��ϼ�����4�nk-�;GY' ��vi+�3-����:?ϳ�̇͌ݛ �{$�^�:wgL�`y�Ĳo���Ω	f5�%�s>��3�ףt��CX�Y�sd���9�C6ǲ��(Y{g��P3�`�鸙�;3�d�Dj0�.)��4~|���j�,(q�<?���T�)��B���4Z�\��e	V�ϫY8[�A=7������!:��L�?�UZ�Β��ך�R��V�2�#��WQM1�p^P�:w���f�F��1%�A������٠�  ��3�jŵ$���/���e�����e�w rP<GP�fP�S�u?h��3x�>a3�����`n��ڶ�v��5]T'c9���o����e�F:8X;솕���Wy���|�H@�]�Q0_���c��o\d`Aj�"�oTvk�Ta|�d�ƪ��{� ��������:��L�}U����MkC��i0��	�e�����L��VZg*�\�}�GB	DK����k0%�P_c	v��`�F�S�kZ�/�+��a+�h?�=�����5�rp�_ �O���_�����=�r[E��w����Yݺdח��u�̹�Y�5G��O����S����K��e�ɖ21WOz��mF'r;'��	��f����֝�{�5HB|�si>�%��H�����?Re7���gJ��`�[� �ce���Իi���v����g���2e�R9�퀒���u��~W�,��$b ��Ŋ?��X,�LC7S�,���9�}��4a��PP�~W������?�X���o_��}�����|yu��(J�$k` q~�5;J�Y���b`\W�`��@)�ei:��zLڲ����0����)��m��,�#��B��l�!#����&�P �����'��b������Zc��0Q�����_[�\g�i�sN}>�A1ɑ���de	��̮�]�}s����l)|!�d`?!A��:��2��nKR�� �
p�	�Y��g��ga�YB2�u���G��J�d:Ö��ơ����J�k��q|zoΣIlM����ث��W÷&�p^[�{�.�i���gy������@��;<�C���|}V��Ȉ�����!-q���m`W�c���0Iɒ覅f#�N���mV[�xx;za"�c:�7H�1w���(4��vM��LcE�Ղ5pQm���+'�g�م�É]+�䛲,_��ڷ�g�"]�Z+8�8j���т�E;�.����[v2.��{��udV�\c�t �I�Xg�xf~�ÈC��zu��&�u_@-�"�����X�b��r��i�'����w� eH-R<�Iə�M+���1�Z�1TT��jY
?˺}�Ҏ�,�G����lGs��'�	ą	{��,�ؽ����YM��b�g�q3x�I�'� 8{�o��A:c��N;�#��ώ-_RP��]��u�R7�� ;]=�kUO��?$�z�zG�=;������G�qf���p U�z���0�\w�D�ϻU�tl��y�9���Ω6�Ez�����?����5�*8�U�1��s�U
�&lɮ�YTF�["C�ӏ?S��Џ4�!�azM���C����	�ڷZ�a��0��<�Jӗ�ceGi,߳+K�l~b#��E2���o��S-��P��q��G� �I���Hѝ3�s�8�h����
�L��{�";�<��'�k��c� {	�8�y�>g����9�ɯ{!K'����{>�"�cP��x����"�=�vy��Ma��y�n�:�� ��3F0Z�ZGX& �Pr�6���j�Ŭ}@�`��yx��;J�x��g�v}�m��FK �xd�����a�u��.p���0T��9�p�F=�^��!�Od(i�ĒE'|�V��n�]�m�������삀�	��y��.�,��$�F`q���� �3����9���|c\���(���;dU@kg噠^�h�Mb����@,����Sq|m�^-�՘����B�H�C�nAe[�!��s2��zp���K�3���in[�q�T$�� ������P�:@��$�mt;R�Yfclj�(�~��a?mH���:��ϷO����O`<�`x�1��~���Η�qD��NǶ��A��I��_g?(�y�.�,s1!qdʑ0��Z���@2���U���X3c3��f>�>�-1)u�AY:��*ג���r��I��7 �e>�����7�scb�=1d���_�^��f�
������I���I0�

�;��n�ɦX� �$�P%i0����ap?ɖar~ՀNl�|���V��)�:}g lǛ�K�.�f�k�()S|�YW���NPu-��8�G$O쩝���fV�W�͉�nG��>��K>�Pr� 6	�M@,���,���o�<\{GL̼�a�����XՀ�E󙦫:6v���[�K�	�;ZI`��UW,c[�k$0��t�(����,�V6̘�4�7d�X��@�� ���{g5Yd�;��}�C�Ww�_�&��q����!|��%,��'�o@o%d�R�>�5'�H�!���ƢD߾}�ϯ������#sc�9Pg��l�}�Ŋ�hJY�R4�*Y����&�����?���
�G���_q=��������H�6�P��_>��~�(c<�6;c���01z�^$6���w�NM|p� P�_��<n��A���py}>e�����/��I��*_;�VgJ���1~d�cZ�)�2�$�żl91q�e�7�R�&+Sl_��z��pP-�J
(�R�!m��(2��Fb���/lw��1���ù����;�s朌/�3cxE}�� ;�%'
��1Mh��H�a�c�ƒ�q����������8[���IDTg�Q�:Ɵ':85^r���&A0�d��S���D�@���,��b��X��k�<@M'����P��/��J4oj���d��#�:����߃dcm�G�bTɀ!0��؟�F�Z�O>QD�5
,>=S� �9l�E�b��);����hY�j,�G����>v~��\�-���Z��Mǲ�&�dp�|��`I�ER�N� w�*8-�NS���{�[5Ts/]���~7�z�4Jp��2���u�d$:;$�r�4:�L��p�����2VA� s?5�z;��*`�\d�LJu��qصI<��h_� V���G~���_������E8��@IT׭t@�{���݇�����y�֥�iU�,P+(;$=�J�c���GŋmTV����[G�3/�uF�R,:�f�<����ɺ�����@0N�U�#� ���F!J��P������{�7F�ۄ�fVV�o
��M�������<L�ĺ���y��}���jF0�	u����?R��//�Q� � �~L=EI ��y>�立0[�����|g��1�;^$��2�_?e����
!8���{7����������F��e�4F�;��F.kk�[�
n��z��s��M�X�`ݚ0�,����Z�&��&��61v�IbRZ��o=�,[�칲��E�f�5��K;@�F���\��!��NoF/f6ϛ���T��A4�쐷��� �a+�+�6���L@�����y/�*0f��\
DM�D?eo������� eGu�����3X� ic�'cS����Ý�������>,�V�R���<.���5�o��.�<��`�X��/qb��ј�E�Ѵ�ܗ�<��
ji;�6^?X@�]���I+P��Ep�V�3^#��Cj��W���1u�#}
�o�v�f�Y>�f^P���j!^���8y����+X$ �p���;�L//Țyy܆�K��&���y[�`�x�Z�Sg�Oe%2H���Z������o�1,aY�(��T�N���!&����0��e�@�$��P|����kp��J����QP���Z��!X�֖3&�B�-Y���^M��{�gW֗�s��A��D#G�v���Fg��R�>�b9Gm?��`W�-��Ox2�@��T���	�6�C�ZT��d�3�i3e��f�s�A�����6�me\�����M�1���Z�Ǳ����@��r�6������ZG��7�� n�(�$8�hz3]��:P/p_b$�M.��ؽ�K�y6�DH%�_:��P����J� ��X"�B�8������rEso'��RI�r��K�:��1���hC�s��ڗޜ�J�%(o;��c��<�`�i��4D�A����RŪ���o1�z��`�����#��ܲ�^��l씨[wp�T�F�X���Ŀ��R�x�=��������~0_��%J�K'�u�/wO��'			�Ec�%ו5���a���̝�� ٙJ����g����φ��z��������v`���o���%'�I(����k��/���߾8CL���I��+����0����X��k��I=�'O�=�1��4�����D���"�AIC�����RM���WlS�y��G�͟*'`�`� �l]+a� 9�!�^� ���E~}�2o<�: w x��5�Op���OC8�=��$�S�zL0"��ͷZF��ќf:e����X*3)I�1��
BB8-��W�{
�|w�b�W�V�����Püv�yR�r��ÇO�O�c60��/&4uw�s�JUy���D[�F�1|�h`Eu�f���a����i�

�0Mf+�^�O��/�����7�&�o,�W(O�叢9k��B@�-*��%/T��8��qNT�[�*kd�#[�8�Qgۡ��|���8ݯ
�F�Mr��	Sk�M7�J�H�UVǎ���=�r��AםP�yˍ�ڍV��_�L%�^$�\��+yr݊&V�p?mgk�]�AN�_�ܱ�*�����w�n~����$9�i�J�Tb�žj���0F��]�e�;+۰cɆ4D0�>��h���A�:h�nI!g�|�z�R�'�A��9Qz��[KL\���� �����M�Q+}��M�����v,�d���攽�obd��^� ��Q;��X���O��8j�Đ���P�h*�C�}R��fۓ�i������"���(SP����X�{�A��\�Z+;�~N���כ;�:�}��ʥ������L����4�ф;�M����u~���ݺ9n_wHa�3$��aw�s�l7�PT�8S�K8+����y̷�l�j5��B�G:D}K��aЍٳ��?�3��.ls�p�;��u�8�j�� �[�#���9�i��%k'q����V���������q|f��=	�t9�I:V!`�3
��h�$�c��@�=�u�C�HU�(����}5p��=��_)C�׌b5��;nǼ�wa�98؄E����w�P	с}�Q�!tQ��yӚ�Y,���;�� %������w�eo�q�����x]]J����xO��g�͉}�� �v�5Se[Ȑ�[Io]�ଯ.ϙ!���k�%rZ&z��WC��'���B8Z2d&�	,M�|��	]���38�g9���',b,]t0�`�?<�Ԋ]�� ث���M��YW�%�d�0z��R0ܖĢǲ����2�d9C󋙀�Ј]{���}�g�l|�	�Y/8�p�=	H-):�V� w��K����J
� �UA�>�K��Z���%l�v�i�ơ��L������r�t�q�ٽ�ڷ�hd��R�$�&_�:]���Y(	$k���G�p� ,��:4uޛ���`��LKn�����D�5΢(-K������U�3 �u��7�|�_Z��k���Omx��xsvƪ�Ak��@`�`�J��=xWf��M���NZE�<�z���]-��⼷��ݣ�'�V�Y�@�_oo�!{கz�E� ؋s���D�ad����O�Ύ�ϐ=@�q<�=ZK�X�x�A�d����h9;,�<D]�ǡ�����)����DG/4p �zn�2�3�M���ؚ�&���FL�	���\��i,IU��
pH��V|8�J�ӽ�kLB�>�k6��O�>JG���`�]� ��3��|m���K���s��(0;D�l,�s�.M����ނ�|��@��أC�e� &���5;T"a���ɷ'm[> "f������ݞ?�uyoe����z8{���<+c����E�!9@��n��R�]��T��r�:�|�E{S���b^�M���"qa�i wp �k�`L��^@�p�"������!�`���D�|Q�:�5��::�b�!as~v�Қ�h˕���cI"���R�W�������۰V�;�NO]lK�8��<7P��U��➅��q���7��W���7��]�Ӏ'�U�Go��zT��`��]6�X��\�D�D7o�X�61I�ex��ά�������X='l��m*�r	��N��O
�A�����O_T@����݁.Y���1i��:X=Q�A�F�-�yH���Yt�56�A �[\x=F�X8��yс�б �"N>[O�@�V�����4�AX.����i� W�o�n�� p��	���D����P�i�坬��ӹ��eL*�ơ ⼳�Z�@��G9,
�i,����9����$��r�8�89�e�t���f�sf�� \Ŧ��鄴�Փ�J�-�T�>�g�Y�hH!70ߓ��9� �3�y��ۻ�;�@Z֕T�49����g�����y��1Π�!��M���mN=H|�x�\�2��+}�W�e@ ��8?/;8�{���.�/�r�|֗��V%�e1�A�z��]����Є����Kx�������s�&LB�rB��#�7b�s�q�I%@̭����Nd�wg�p���NCPg�!��!�b����@�c8D�K�Oi�9�!%���!�L���]��l	~XkL���݃��<o�:Z��1����d��<���-�D�ͦ�0HI��w�6�r�ׯ�1䌟����xI����+"�3:{XWGv�� �{��[R�iK�e�-�0+dQ���Et#��&(+{�\�t�N��ɿ��Y/e;��*ю�0~[X�<��n������c��AAw�
p��]�ϥ��N��d�f-q �`l3���a�;��CA��ˣ��U�92ȣ�Iv��x�(��C�%��)��m8�}����>��4��m�u���q��h�e���o>��Q�	�8��6d�,�K�3�+���wW����"_��`�0;�,&;�<�p��3�dm�^�Yij��+ $�b�4oZ'���c�+;+�*,+��(�wx�..\g����0��m�u{�p7�^�dz�FJ�fde�)Z�$%q*M������CI��e��S�6�b���@f�� ����C�{ӕ�����E:�L7�����:��{Ä��ݘN�~�܉�h��N�י��M6�|4�^�=�%�z�ѮM��\�X:
����"c�a9N �x���ZAveb�O�ʽ��#��`	-�E�<��ٖe�&��m޽K�H־>Hǯ��Yw�o�,:_Q,�H?P̮>M,c���VF���%FT���Զ����[�ΰ���9���f�p���	{:mX���s�?��遬�;�J��,�Ls{۵��m��L.�c 0����~�Q9
$ő�A�בї�  �@zg�bo� K�{�e,,0���e5���-���^��Y30_�}o���m�5>�	��3�`?�(]��^v��ow7���5��_����sx����s�8R�)_?�ML~��Y?��9���;7Ѵ�$����˳[^#�6~��*���k���W���1�9V�
�& �HvM�k>��O���u={�HM�.�f5e%��c�p��ܒ�,t�6�)��.�^unC�U����;�h�'�#y8�ٛ�p}���� �vdl���"�YT,�$ɗD#�c���|ܧ�s?�x��0Y�W �u��K��bM0q`�Y�ʁ#3X;u[���4����ȴ��w��%�⌯.���/���;Eo��7)#B���Ug�����+���X��/��Y�aa���*9�qD?o�����"�l��Ѻ)Y�� �& �7�j�M��8y�;�u`��ɡ;y�����o���䏊ȥ����+����4g�fԈ��G��+�?����c�{��_x0"��鈅>�tm�SNӥ!�����~�1��n+�����	�v���[�F�w����އ����;�*������d Ь���s��:~�.L�pZ��*j����y�0��#�6����R�wD$�FØ��&�P�����Cx|V' 1|oFr�R&�I�@�՜�i��J�z(c��@��\K�Ra�c�;�ǲ�Ũ�9.��` �b�������M���3�NPW��}t'ǂ,���?�uGZ����Z��* �%�z�����W������2�}�#�����)���}���c���a�FVl�Q����&/���ߊe�k۳3k���:#��}�{�O?��cvԗd�<�����M�r{��
'{	�I����c,P؆��F��ju���Fb��D]��p���uu�3����q<H�4c�9KT��G:DNYM��,x�Q��[|�0�7X+3f}U��X4�m��E 2;f/9P�ّ����CG�b�q8^A�x��Ƽ(̭��]k�����F,fl� ��|�5&q�Y�ȫ���j���6(��,�3����8��q��-��ݮ P�q�<q֘���Ng�p����O��ҥ{r\���{!� �A�z� p�Y��� �@�ԭCj~��\b0�.��j���YD2�DwVr�sB�@0�0�p�d,�� x���ΨfK��x��Y�k� N:}Kvy�yf �9��F��;�x�݆���S�s� v���������0g�������;��V )���a�^��������3 �p��.|��C������U��
B��b�\^^���)�(Ag˛���?�ǿ�6��8S�`|��3�W��C>w��5����L��Y7#��:��U�F<J,��œF�eu�Y�C	|��sǁ �n�!����@8�7|.�" )�ΩN9W(��	vRc~=.lMH�@b��-�:�ٶn6O��9���>��?�b	�n�R�z6��2'c�!(~a� �S(�Ø���J���\����-�0)�qi�˲*6������Г��|�d�e�� ґiO�ݘ�S&�=����ƘH-ui�T@"��RI��@�T`�q�L�e�x:�R@��0�xH~�j�,֦� �v���CB[n���/��������[[i��Yh�.XL�V��/�pT73g�������_ջ���y����>S��{�9�'�<�ŷ�b��5F-��Z����6�4Aog6�NLue8Z����V�o�����+�+u��9�b��U����V��rV��u�\��%I���uPE@��%����͓֭��C��~�@�# P������ta4`7�v<�<���U�Qt�+%�e��Q��v��~r�&P�1k�3ܑ�w$ǆPe0۰�k����>��}4�f�*�@��FzF��{��(���Z�}y9o������\e
�{�X���Ls]�*P��͔�'?Cj�z���UJ��^��'KΠS�U���z]�o�l��+�~�� ����b��
V��X,T�ޏ�aud�~ ��c���	ֵ�>lw�+h�@��F%�����V�w@��͚�g� �)��]�(݈�]&��q,Usg#�(���{]�7!�k�-}����1��[
����<oR�m��ј7�����׷W�{ �/[��\�A!Z��O�Ěꋶs7OwU�hT�:��4Ȯq:[~��B���l�z����O�bS��dC��D"w{(G[�,J
篠,� �X����h.���˩ՁDC:�S�[F����];Ԯ-��X�~huFw@*�P��ZW X����i�¹$t:-k�	���#�Z�3��wJ��*[Dw.2��*��)0J���@�T{*:�c2�����ǻ�́���^����d>5*�8�:U���p��4݈� 6��0wBT��.]񮡓���}��)�r���\5���C��j�WY���9�SXRZ3�f�	<e���_�55�c�OIF��ו?tu.�L�b�F��ƍ�d�e4TS+��c�(�\'��N�#~����Dꘃ�*+���:- KC�z�y�߾28��B�˕�zD:~�٩xzz&xrq}��*l�<><�;��}xxz�A3J�n�,7��t��q��[ɘ<d\���y���.��v�����p��gۚm 2�� �+S~�����3��:�W��!�Ā� M ������x�����f���Ţ��&;Q��<���Ys�PAB��5�����v�@��-Vo^-A�`�i`B�к�s ��g��Ɋ�1��`^d�p2�6d!�ʬi����!����>��m�Q���:;���|�egz�L4XQvѹ$�u��i١���XM��aST:���ت���*!}���yb�ŹsF(m��� F	~t@�ɶ�9�AZa(���߿���`��V�T%%`K	�b)Q;3a_�ꩈ�=���۹I�v���L %g���ڂ[d]��t�C�$X��9���������A`�"�?��@�b���L,��;�M(��i�#��^�-��.?[��W�vO�pwwC���&<?m��Żpqv>�<�fW����;j@aT���nvLP��?��l7�ۣ��g(��$ %�し�[ky��dD �&+_�{f�VG[mQk������;�[�NT`���~�a0P	-(�	&�E���u�JyO&`-���8�Z.�-���1_������@�2۹�w����&���yd�a�䱽>�� ���H�v��{o<�� Ew���Rd�%֌24��X��3���Dg�=�NO�?���� ��(�`�� ��۱'i� ���#(K {i�2PG�s6^�=��S{͏k��V:��y�>D��^~���ITR����(���5ͩ��xe�/;����+ W#a]�k0��Tƹ߫�0��om]�N��؁g�����wxtq9�C�}~��ϒ ����e(�80i�~�FX52:�r� ��Ȓ&pV~C-�9}C2�u�:��О�H����`@���KX*�˯E2���]����4��G1��`��
��k4��b���ܕ�t�z0��Yh�bR�"�6&�\y��z|�v�3��
���5��,0i��-a�	3��ì��� k/���˷�Q��L`��ϭ���c�̓���g;p�u��Vk�%�UQ�`�MC�A�-{-�����`�@[ˌ��f�(�3�r���Ca���p�WW��]�bi�X�L�2���7��C�S^����,�\
����^����!�{�������t��d�����(�I?,�}��{!�@�	zf>gt�����H��X�-�;�$�)x/M�<�qp� ����#o���B���J�V�۝�H�<��%��+*c���y��c�������L���e���0��B9P�.!�zB���a�,h�Pzx~��9��T���t��<�}^��@�d��yR�<��Q	�p�X����ߗ��x�1Ă�����?�4�2y�F{�@���[h�&/��[O1
�z��9U�{;0�ǽj7��#��/ʖ@s�sJ4�f����*�$���kL��@��Ѩ�E�7�S��UWAc�)�Q"}] �e؍�':��5-H�����:����A�{Xf'�?���p��� ���C�+f��`e9-��Z(���	��6��րh��Ќ2�</d#�C�nu8�V��Ԓ���Q�Y<�X��$��T����b0-�J��fT� b�ڨm��������8���,�S`��b�2Q�p-��V%�i6�iV�CQ����(8��xh%�s��N��d�Ƙ����«H�;��2�1�}�C>;m8����/?�X������j��N�uDY��N��>��X-���̇|�G�߾0�_�߆�?��}�!��k�7����o�n���!l���k�ٯ_o�/�n��6;���%�;��c0FP䴷t��1����p���yv�/���!������w����%M`�DFǣSqt�Ը�^��.�d���D����޷�o?\��q����H�bX���DI�����e� �N\�E��K��W�9�gc�y܆���ֹ��E��8��g�y���8���̴c�����<�(1Ծ��{�{���wr^ �6y̏�r��E'P�k�!ܜ��n�LP��?X=W��?^��3�s���! ��,.�	�7�B�y� �λ�.%w��Q�b� ��2���U>'>^Q�d�A��)<�,âEw���h�^����vFsg��Nx�c�{;�a[�dG�>g���L���,��(0��C���*]���_�V�`����>ۗl���&�ҹ��/Oaݭ�as`h���)������9�V�痗��A/�N�xJ&�k�I�
h���=�թC�� �o�c��?pߍ��!���{���x�xW��pqy�>��~�1|���e_�ބ_��K������!J��f��警;�^]���'���pP0@@��le���t\?f4a�i��m"1��ɠ���#tؿ��ݸ#���o� Ol�,��x@���eO2�l�E���r�-�`#��g�^�&/h���{k��ꜯ۽��Cs���1��<�����S�����;u�ߡ�U�$������2t�9�����g�^�4�rwd��L��l�����8u#=���;��G��1���#��I�pmP���M~���y-�9p�%Jf�c2�溦Xd�����ck��XJ芥�$4��k�M��X��f���[)�|��4���i���tV��-�^V���
lك���&���3���]���܎ꄆs[�si"1͌����z��l�6�����B_���]؍ů���P���J�XN_n>+�pl���qEs�`8�^��������H �ec����$��c����0Z����+�����A�b&?��A���"Ƌ�����sj�m呰B�=�)�c7�V�J$D1���ܕ�� Y��w
����;�x��qax���zNy�5Ή��Y�s���z����ҼB���=�lxm�ْ R�vמ�5���HRa@&!/jԇ1:�PZַv����yf(�ʚ��^��ڣ�6��bu�$��6�2�NY�����8æ�GbN�C�)�m��Pb���?�+���5��I��U�v~c/�Rῢ\�#}�6k(	���,ΩQp�{�p����zA:���C��h�o��h&:�*o�,H-AMW������E���d4 *&�!F�kK����U�Uk��x�>:]� Oڽ�P�%�5d����%e5yɃ䡊��	��AU\36��9����7'���_a�k|��4��W�u⼝2Q���h����6{�up8R0���a
l1z��j��Fg�,Ŕ��� Se,��[wgo?��J:	8��>y�2��ם����������fH�����e�-�Uf��������A���a�(@FRd�Dm��Xl��v��v���Nȍc�: R�Ɂ߷]�S����,�[]�.;c�����p�,%k��A�ve�(h�1-�-��J^��1T�p��I����G�_�i�Ƥ󚷨q����;̲��R3k)^2W�MU;����fV�m�4�d��(�z����6U�З�];kO뽔���d����
6d����$� ՘��E��)�!�J5��-�m7O��滼Y0�\�.�r,�"�{�5�Zpγ���� �{�#h�N!ox�9@ނ�ْU�wZ�K^�_~�8�mv_�k�:#�}��T:��]�]ZF�ݛ�Y�K�J~�V�p}���_͛��{�E�T����[��G1U@�_�9?_���ev4�͗�r��M���ո�w,��P�P�g����4$�@#;���9;)�j%
q�	�6l��}��R3
�h��!����:2���*i�,gK���ܙu�i�u�~��ûp�r�����v�?�jPy�A��8�<!(w%c=dg��">�����c�����}��tH�����)�F��������G}-[y�o�E�\I�%D�CZf�8�K�oB �ٽ��ia��J����N?2�,H}����b���
���=�����J�"��v����)�?=����� b�z9tcP���@-�M�>�q8P<�J��3�/��uy�NJꎓL�6�5]��xb.NTF;#-�ܘ���A9��E�e;�}�0�8lT�D����}���]�s�>�y_o�Qk����o��ɚ�Y�2M�g����7P`��t��ذԪ#x|�=��MO���u��4p�k��k�^��_ �5P��;��=1S:��G<DY��.,.Vd��9����kW[��Πn&Ü��q;R�h�T��;V���a�4�]�PNp�׃r�U8�>S�!4��}��}A�g�(�� �o,�E(��Q�	��Qh�[X��M^ͱ)Zzz�u�N�' <�l��q)�2�1ʼ��#��=˰ �ęg[??[�f�_Դ~��xr�6
`�@�	3��f2�q�#����d���<Φ�&�P��G���ybF��%��+��\t�r��$����i�:�R}tx�A� .|�|b�� 拳t�����>	��r��;|4ȀL���z�:/�L^���Ș����5cͰ���h���q�>���E	�J����/��t��-dۍ�8�Q�s13����:� �~vc�m�5�<�g��g�z��[=G�c^ſm�s��j�]0��M�J��	�$G�L̬��u-�)oc��+R�w(��"L���W�]S��n���O� ��W��e|[�,:�c�E�i��[�m7~h�6�Є��tr��A�Ι��1��^q,�v]G�ڈIhj��&�0y�?z�jM&�B]������+�0�2�Q~��(�s��cw0Ƒ�v�U)�j�,����@`�x5�k���'2wb��g��8N�6Ƃ�vyÄ��J�{C��>^��`�D_)��d���6��d�LZ�ѽ��|`O>u��8s۶���S�F����W�I�Mz���[���ƅM��|��ʻ�%�)���F�v8Q�	��=�t F������K,o΋�K"�Ȳ��M{f�����l�ѣ:���8�]�&�|�gk���O�>S�f�� C����#���Q��I]s?�&���!&5m�轎���S�N2�:m��F�8�M,��I8�.�kX���T�j$����ɩ ʫ�������L1����H6�~8Ow�����7�&���=��&�<�M����^�k5�b;���[H�[sx28��rzl���@�b6�*YN���@+�-���H�����c3ǚX���ٿ<�����_��=��!;��C��O�V�L�{�Q�b#[�3�&�|�DIg�чP2ښ_,�����lس]82�i��y����7��.g�|�`'!���_�sԧs���_<tN^>%8��sfv��5?a�0���6���@$ _�*�!#��2\�A�h��o�ܑ�ѢӢ�(
D=R�f�,ט��F!�,E���b�
�}l�����3��G��F�X��{a��6w��F6C���i`��LA���s �F�!ֹ�nMr�3�"2�d��h��z�O4n���r�ԾuM.�l  \�ga��� s��=Q�(䱄 �d�Ñ��h;Ks�婭rG�?���@!2�`f��;�E'q�S�SB��]W����ʰ.& Ɏ��r����O�X%JSQ���H"�^���9?k��� ������ ��U��粝�ez"�P��S��Pm���Mͅ-��0��'J�W���UX^��N�q��DG�*|��5�ۿ����y�$��=f;qw'q���g#��h��Q���Ը�$�č�g�*� ;v�%��J��C��!ש�^��LKkp��Xr�Q$���8��3b|_���)<>݅�G������/�-�Z����c��#2;K��3���O93��=6�܎��gK�m|J,I;[.��$���P�� ����h��` 	L2���ϑ_~yue�~������Qe��b��w,�˾ْ��0��1 6 ���;��	�{��:��9S�w�{�"J�u�o����$�p�"��|�v��e�Ƅ��0ai�U��4����4c�tu����`�hz3�97v�xi��J��J�,I�ru�;A��h�3��	NoB~��׺�דk�|�ϔK�}�^�D�Dv�y}��+���D��:�C]S�����0�1,�P�s�|l1(���J8Χ7�u��`:,WL�"� Nc� )�%�E`D��;��j�P�����d��k���0�����{�Ƒ[AR/۲�Qս{g����oڝ�;ݷ{����,�dl� "HIά��e�ҶD��x �� ��ۅG���hD��w7�B4m�uX`�c�"S���q��(���i*P��粨1 |�dYg5{���k�Cp��9G[��|����;�6���F(��U0��g �z�e�q�!�KŻC޳�\Ҷ�z\j�g���-�]�N�h�qX�drQ�l;�\~*�Sf����.�:��g��&#��j+k��b$�̗�s4����;V^�Y��nV�@(���:S�m��~�gM��h���AiD�΄G�����g��PUC�c%$<,�3Һ��z��`��C��]��/vT�۠�(�y�m%�jA��Ę�_�w(�t��͓�E7iU�#�y*l����h����lF<C(Jo�6�ӧ���S��n
ߋ_��f�ۓ#+�������L��?}��ruw�ޱ/�ޱ�ݒd� x(<�:��Ii?���JD�qzn>!�/y��"���!�|t�)�a�h裘�t���)�Ώ-�|#a�����*�G��������c9��f��I�r�t��S].L��f&ߏg>=#l������%`V9�f�pN�+�2�\4�J�S�<�m��q�j}�8L�˳�����Z��dԧ�K"��D2^%��YI�G&�����t*�N،��yP0�!�J4̊M�8q���-��5 � 7 �E�  T���9��E����C�'T�K���l��d'��P֯�&�i����76&��t�(�~Ir?D0���ij0���GYl@Vܰ�bw����6�"�ko���Ŕ�V�C�'�EVK/���gGSwuM*!)�G�Y��t�R��	���"�ӽr����
���9�(�'9����n��[����7�&�ֵ�2�k}��a7V{��^�ze��H�J����z��J����4�G��v��,_��0ҥ`0^�:��Q�ȡ��`���ux���X�A'��(AX��'���C��sF�r�K�븒�&jƈ]Pk���}�h#z���j ��� �A
x_@������6T�nE���5a���k}wNϙ�cO}s�Q�&+��Ւ`�9�Z-	�B��T�z��&���</�ʉJ�������!���
��T��=�e���m��ND+�F�D(�Lˈ}ɨ�~�������ސ,���t��ǧ��������3�2��!���o�_�y��P���թ�6xVx���S��ރ#��H�`���6�� ��<K�O 	A̚�u%L�u�)-�8�t.�vhɷ��+�s���E�b|��t�kE��*4�Z���^�k���iN���a�TG
�`-uA9���ٰly�?j���X���v����Z#v�K��x~�)�S�/��fQ=�\/��d�J�{P�ޠ�ۂ�1#s�!�Q0�V�s�)*�$��Cq<���ݽ#��x�Le	�I� ��>�ș���ڊI0��k�&��Ze�����!�v��y�.�В�]oS_��ͪ�Af����5R�A���
aM̴�a����V�ˊd�uS���m�`�S����9�~e��8��KO�Uf�!?� ¹V�Sj�nL�ƍ� b�:T<�����B����`����`���ΰ+@���/;Ny%Y��A�hyvK㲃�ϋp�)>�M4ǈ�i��,=]�=Ոd 3��ס�YC�<�Br���[f�#�ˠ,8����7�)H2q����b��������8i,k�����|]y�22������S���R�N2V�p�6n=V'�63o����΍XOA�S4� XKkܩ��T���9^�qvh��u%K��kP�T��e��+�WI���+��3?���s��.���WC��e%�DHo��%�z�ڱJF�+�Ps�{��ǫ�$\t���C�7e!��U���k��4v#����˩d�iU��&���-?�_l)�t<���aD���D�$^�-���%}��G�d+#r�e�k��x)j��k��U�Q?���F�H`�PLn��(�A`D�n�4���O��Q��	G�m����42�Ja�U��
`�Uci�D���[V���<��d�Xpе���
�Y�K*��H��/O�hT��c�&���v:�'s6����8�Sy�|�i�8h����c�LZ]m8�EsN:�ӗ�E�A�I�t.�{��o�޹3r˯��n�_�<!�!9�Z��q2�Q0��'��'��0�g�ɴ� �|��u�7I�XA))���<������B9'�3ʆ�Q�t�$��[�:)���p�&�&��D�(���Ȓ�H ��:=�piG��`3�M���wXo�d�]k�@-D��*�[N��߳����h��X/b#z��*a x �+�2e�����"W+�}$�e������6cO�\�����yo��+�4D�43�굚��1*jA%�����#]�5AA����Q����$�ޥ=���}����TgD]��W��D��'����gs%�&sݼx�#�m	��<]BZ�(;$:�,i��T��=�2��Gu�� ���742�[M�Edˠ��B�	~�MG/�F#���?N�Oe�u-U�i.�qzsP�$߈j�<���b"�R�F��*���/�z%<�4}Q9��I:�ɱ2����O����"����$��P�=�{��#�_�Ϯf���e���D3ޕ��j{��[o��y��N��X�9�KZ�H�uNV�Y���#�ħ�'����|��Ո&5a� �Q�C��@"�Ҏ��g��d++���:<G-�����V�=�jk�(Os��ݖiX5��Y���'�x G҉��`�z-W�ײM2��\B}����Q=ַ�L>/����h�7x0Ob7�HD4d[�ɒ��#TIA����Zn�����Lb�S3 
 v�
<�5W��1�.�y�\lh,P��;��o��>:�=��7�"���Fa�|��I�H>D�@�!j����&�m�9�D:��_+Tbʖ0��+�����3Ҳ.�z^���`�HLE�Ƈ����A����/�y�>+x�b!�&�������O��� � P���.��5#4}�Aѐ�/���,F��[�#�	�� �M퀃�^̂��ؙ���0J��)a��<k���f]��������o�<�������Rf}��C��=K[{ܱC�4-�/��	���L���t�RHC�磨��y��Gi� w�]�+��d`�pk�J?��f|e"��d�"�T�Q�A�Ńk��7L/�; ��m�^��G^�
��^i��GW��G��3�����'a��LN�|� ���Lrg�&�7�-pH�aJ�"���6W�E��fd,@�������xN���JO�T:]w�6d��~p`_AZ�}+��D:= G�V�c���y����0̏���2ɣ
���y���,�ї�6�6�@�����p� ���n�&%/��=���M7�W�P� 2�#Nވ����mg9���#K��?s�x��։���$�R�mV���"�����s�������NO����%3��g����/I��60!���z|���l"�߿��y�Ql�� W���`q�C�d��oռS(��K��{�؁r?��Do��}�����c�vĪm玂�_�)�{�1&`]s���Z�s�2��R{N|��"ż�@�:9�Z)��gE�?�(9�Q�nLG�D����z���B�JN��G�[��mi[Q�ȪO�r8�|n�\Ӯ����̻Q	�����ĲZ�GiV�(H%��z����~Ϳ�x��NwɸH��:��U�pX5����Qy�v�w��)@$�M#*0�3�@�^:(\L�"�1�K"��^�0�z"7��˸oo6r����+*�0����$]9���C7c��h5�gA>T��	�����D(D��BLRv{���@����I�c2�Fp�,��PF����Ay����3�QS��X82gS��
�V�zI�8�" Dۀo�a���G����'Œ����;ʚ�Wg��$�|=��g�{㛾��5��S4�^?��t�ަ��7��aQOz�@,�B���!�"=z���
��㽮!D�,7i�_�P�9�0�A	�s H6����Bô]n�`�W)W�ˣE�D{ ��#a�j3X�1�J77��BGˏt��]���}&���=lx�e�2� YFEA���es��[�Jk�$i��6�-�h���U3��Q�J�x��)݈���f)�i}991R����-K��8�q�!�rѲ:���-A��������PQv�%�CLy���44�)\y< ���"I\J��FA���6�׈��Q�Aj��|O�DD�@z�0,6i�N��k�4!�H$��H &���2\s4���*�2�k��6�7�5�*D�6�{֔�o�Z��mH��6^�nҸ\�4+�2(J�D�FS�X%q0�F��7V8��⨟1b��k =H��k��}���H�#�������A�Cdq�ZP䪈�!u�
XH�ZsM�Y��l�Q����\��9t��v�g�}��ĹY�X�̮�r�k�\��DK����y��K�Ի�Me�k{�Z(vυvd�/L����n{�1Ŝ�������-�DYr�h�TA���OÐu�����j	5�h�J�hx��M!���,&"����	�c7���&����ٖi-�Y�Њw�r���/��r{�҃��������4��s�Ff�R.��P!i{u�v�銟�f�|i�z��{f\0�H��0��m��m/�\L�F�q�G���
���Z�����9�߽����,' I������������#�l?3��5�O�H��t�h ��Wm\�7AO�nT ��ϵ��~D$W���������ߗ�0=8���0�?+����d[56NX H�u��7�������0]³|�9����n��p�#�޼���fꗺ\)�^p��w�c�yv�����l���`���⹫I�& �/�y�K'��|���vV��f��O,i�ʢjXoͱ��:����N{ u�i�{*��;M�d~{T�|�H>C��g4�g�����#ׄ����ҍc�B�9��V�&A/r��8����'���3�/_>���Q���G	ۭ.�ǭ7Xl��j�L�j�cw�K��+��O�%:;�=��м��BȪ/�C��܌����' ^G����� ��E(?���sŌ�)&q��f%�6QԔ,'�_��w��M�e��}^��Q��k���Μ������$�_ClRe��7K�s�k�D׈oD��{^��(��������m}����G`'������6e�Ӄ�ȝ�hoƥ��%���55��$�Q�.�'�Z�\ޤ��V^�O�
/"�N�@�
�X�  �EIDAT�'�pl	�(��ZI�H����w��B�-�8�7�PP��R��kVϨ�#CW8�����L����0���_�rģ��ٚ-y�>&� �hC,����i	 Q_�a�mpG����|�ER�:(��R�A�|w#���S���K��C��C�Hp��Q�;��H�^}�;OJ������g��$s������]z}�1i���"��|�~�c����'G�[��	��=Q�c٘�ASR�T�D�̌)f��C]\�z�լ �Z��*�Ad�R#+��ߨ��������\Q2��;�	�(s���K{Ȉ�,Íʌ0��4.�F��%=�K���x��Q�됉��g7h
w*f�/ ��?��GV	��k 3�ZyD��3�<�)H�_vO�Y��{Ls#)�x��r�ӝln7Zz��2���2Cm%���ލ3g��� ��.3LR+p�1���~I�^e��JsX�v,�I�}��s ��VQѵ�k8�>}�$�?5��s�<�ݡe���}�Q#H\�PXk%�$���:X:F�Cz��X�B��a�oRߥ>�M/Tp�s�@��{y|y���{yy}L�p ��1!X���Uz��<Ad	F�n�ot˼�� �)[y`�;yNE������"�H������Wޗ�˶���M�k�e������(.}`	h ;��Hu��J�<�"V��@)�y�Q�X��� {�> eъ��x�P�7 ��Et-Yժ!���b &_�J罼<	�]�*Xi~ :i
��w�� /�M���uP����P���YrzH,仢�'�D <A��j�����@�R՞>��2�3�$u��9%]��"v�9��ɍ�G�a+���=\�R"�FE<)�ڮ軥�rsVs�3/�MC���/�����CE2�z�=���l77M��~�^�I:".���1hխ=G�1˥����ME��;�ɴ�:�ߨ�?7�Ͷh� �z}��W���*��Z�z{#�?~ }F���J�(��iKշ�����eEUhϘ��{��:�E�J�4�,���<Epߦ�6�1�
�4�F���?�gFH�
���g������3��;c����6�ۜ"W��k+��`z�!�p�#���J��@�>ZD �J�R0U��[�y���m�ܬi���Ն�W:!�L.h?nHf�#)�0K����=�9j�5�id
��×�|߿p�Ւ����ņڶ�u���+<G�Z/��v^�@��k�MoaEj��oa�i���!XR�,?L��O�Y���9o��	M��I�e{��`y��9˽�'���M<X���KJ;R�B���Ь�����+]8H|�_��Mj�2d��ߧ���DV��6�]al��м���P/=&�H��E��?���	蠢ؿ�ۿ�ׯ_�AbԌȄ�x�lM"L�6/.�|����2�iS�(E��0t�����B�	�,\�*����B��yB��-���h�i�>_.�g�|>�s��_���pG���g
@�N#�@�9��1�YO�������'/�i�
S�)g�)M�K�XH�j%lz��p��q�Y˛�3���c`k�) A��|��r������m��2cw.�٢j�9m���z_h��Jp�\!b FfZ�;���{���sG*�H!�`Zs��,��L��Y�`?<ͽ'G�������=�H�����F���Rj�/B�g�NdB�@3���&�<��`�ߒ�BA��Ƨ��y���
��q��i'�FN�m5u�7�Q�~CyNV4%K�?5�i;x��ERD�q�����{H߹N�>�;��$��jӑ�� >��#+_*3!-"PP���'��V���呺��z���t6W7r/������6У�<s�|0���%A����I�ttTA|)J��S���>`s6�R��U��8/����ѡ�F(�^	k���ّ����M���v��iY \FJ	����+��L;�� wC�(�[��s��3M�aU-D9Ge,=�Z������;hʙ��,1��C�4/l�λ�fBO>����՘ 2\��}��ZW��.�X�'xU������UvŻ�ٰ}��B�]�j�Ɔ��QC� D�����kv�9i�0b��
`x��۴F�(����ݞ����k���t,��&�8MS��8yO"Twb���}��|0z��w+�?�9~�� �'8������_/��$�䧀�����\Wwi��<_l�>��y��]�a*�����m:d,��5�-;H��d��FS͗��ɸ&���r�c������#�@�^�vd�k�wcD�K�L�k����5�	y��9i��O.I�L��S��x{ �L9"��W�2Z��B�
��WV��ql�s>ɭ�+Y߮�<Z3�.�*J�z�򪰣&u��j��U��y׺���e��A��3v#M��Q�1���b༃3sn8�t���B�V���c�,�4=��`<?m<��a��"�� #w���k�,5�	�W�HĶӵ:Pm�5�e2[��c�E_锞��dpHAG7(��5=5;��KFq�F)��kR2<�rIu�am�S�0�E�~��W��Ͳ�ۑ˞î�iL�@�<4F�x�.F�`���)4�{�[�Ӟ�nU?�����Mۋ��{���F�XŨh�aJ�f�d?��t4��ʵU��*e΅��nC�*[ꨚ٧�������HG ;;%K&��R~YB��ر�c�����o)�n���ږ�M��c�ƃ���m-��dӚ�����KU�s�G�|��p� ��ī�U?k�����1�
�Mg����8��R�+)S�mjW~�8�C�ގ$���qw$�
y��z&;+{�f�� 4�����s\�GT�H�0rpQ@�IaS?�M��<w��o]�2P�۪��b��� \@���7 k���exYh՝
'ִ�A��XA�P"GN�N�<!��&�^���O�M��m�r�{����c�����Wx�(4Z�c$�O�9x<� �:_�~����)!����ӧO�{��z%8Jb"������
�q���|!6?|ѡ]��zI^ϏO�D�G����ZN>��A�ѸiB��O���z�0�Ҟ� B���r�l��Z�Y��P��\M1e���,8��-ǜ^�+䘱��{f�bO��7��G�Ry�T{|�}�$���?έ#���o/��v;�Va�7�1�Lo��鶱���_��qc}!�s!?�^2Fb�\�ko�r��K(�#�S"�/�UC`�=<�T�"�i"��	���W�d��(��@�N���P���}靨^�`r�Cզ�b[RP��ED4@r � ���
�(qn��d�޾�ȇ?��w���nk�=�<�9�w���|'�;u�c��y�u.4�R����l=(�0�ץ��=�He�k�+z�����*)O�����M�_2�ɀ�����
�}w��>H�:�1C�Sd�
"EV�� 06r�M���r��g����ۻ�P|a��-��w�{zN}�d����Y˚#��a���B*�!�f�H�K������TȻ�������D��RYa{��F�|��Aӥ2��Hc�j����*�����}~���s�h��^#��=0Zul�j�, �nԊM�)R��a4�M�/������E� ���q���:@��:��ٰ:�H(u��%�Qy�K�]q��/@���qO�Q9D�|'���>��S\h�����ZAJL�f	��MfC������!$ h��mP :�f\�a����{zyy��=~�� ~Nk��=|�/i��駟�� �������4瞟�S���}��3��Y9eW���,3hj����.�� ��햀����u��<=���Cگ��(�:�7r�5A�k�%3k��8D¨��I,��ä��@a��iH�#jĔ�՝y���aE��kB#'؆���t��ˣ���"B	���uu��N�����+��������F�͉�$P��+攥��TCD� *Y̷`��r-!�@�����K��x�)��P���5S
1� ����Fp�@���&u��"����	�KĊ�hw��&<F�נ�0O�`)E���ƁQ2��Q+�:�X��X;݀rG�WE���Q�`5>k�B�N.k���0+�Y��J\������hD�
wF�;[�63Ka�"��YU�B}��:o�h�a9�V�l>� �����;�hÌ:�x-)[:������%��5E�T�UNb'������I�>B���jtZc����Ŧ��jҒ��ə�佒q���
Ϊn�x)n�����W�(wҍ9rf�2��Ad�di��f#T�$�ܚ�����9$9i%�s�E!2ƥ��:Z�لv�m��͠�p�� ����ubh���{6'�ȑA��^~W�w��D�:���[��٨���Pu��u�P�A&�����\j3�&�\Ƥg��p̜9\Ma �V��2΂n�L�Fۛ;������b��Dl�y�rqY��y�m�e��R~�9��n�N�8J!�
^�r��Q�- �@��������Y�8�r�8V�Tk`�y8}��;����ż�]8�ߏC����c�>�`�.���*�w��5���ie8�M�d�P)��yLD
qn�˱�`�un�L���@z�z����@(��v㳴!?$������${3�o��-.xO�$��_�7�0V�̱�rmF�%E�ރ��%�w;�z��mW�͵rY�y�����Qf@Tu�Pͱ�5���kڞ�]��YVT�j���(G�:ݢ��n�R�N���p��oYK���}gm�+�~-�,��Q��='���S?�	��s�����s�ٷ#�u��Ej@"�#C^Q���D?��v�'{�f����Q�A�凊��� �#��EK���	�4�G�]����d��@��)�a�I��\򼩉��ل+��"�
1%[g�[=���«�y*WWK���Vna(ܬt(0��:έ����,�&����c;�Ɍ���qj��SbL��F��03J�X��D"դ����r���Yh��6�FA�J7��M�N�9Ԫ��I;H��ls�"���쓢��=���?��O�?����O��<�S[��{�i�Z��=�x���Xi�/�ǡ�^�3˜���^I�R7�q�����Q���0�1��5g4�������
p@��ZJ�~^<�XHsw����7^���6��l�ݫdH�_A}��G]� �S� X�U@#Ǽ�b)�1Xꁨ.���gMC A3*))��FpU���)F���;vD��|�a��%�=������h��I�ѩ+Y��f���jS���2՛A��;�z��a���"=�e��� ��O������H�����<|�W�:������_]�: �=��!ᱦ�d@��+�h�Bq~~}R����L�y�inӜ�ATT�.���0:�`�5f;�w�	�T~�Z��N=#��3�Bu#��#��r��թ�AJ�|�T��Kҕ��g8��Ղ�[�ЀJ�Q��
QR xz��Ty�\�����pAߧ��)�!��p���y �X���(Df! &Ӱҋ@�x��w텈(T�Bz#1��躡����^��M!$���s\��tF��أ9����Ͽ�����V���xEts�7F̌eKQ a��T�c�SEή4ӷ���%տq.!q��d�^�v��-����{�4��	��E�=�ܫ�Pt����v��tLi�g�`6���n2��\��0�a�v�VU�?�z��F=Sr�6�Me�f�x\���Wo�N���"a��k�$
O��̒�i���z�����lk��B��u񑍖����q8���==U42H�,tvf{ϪXq�0�;s��F}��AO��6m��JDRc+Y!4��I��$y�~�g4��q��L�jNy��Xg �Q(�ubz�Lն`Ք�� ��rN�c�]h4�P?'T��� �|5�;���U�4�C��PYn��r]YE@1P��f�oW>����eQ���s�|�0ϰ3p����Y�"�MH�k�rs%W3�`7ds�i
(� 
$��c�aՆ��yc�l��=}�,瀟�LK�w���O�̼Oe�7��(��z^�
�Q�Ӈl�f��d)��U����EG)�8��,��,�s��%ΕLLOo����|�B# ��?� Ѓ�qh��S�rbTj�#ӿO�C���Ԝ.��B��iU����O/ʝca��zY�����h�;�]�f�ѽPq~^#F�f�	�\��g1ή_�9N�=_v�:�C�y��i{��`[X�8ˣ�A^BQ8���f,�_nʼ�Л;�������׻�i��QC�z"�=+4�xm�@�ʏ�#�Y�8���h\ѳ�3��a-cT�	#Dw�$�1�$p�t �D	l4+�<f��K���2��ۦ�c>$�?RY)w����Ɔ�����$}�V�	�A#m�A#]�����u2��ɠ�!!�ܡq����HO>�;ZE@���	�E�/������Wn��Q���)Y�Q�W�MO���-��$��ط�ք���Z��=���K�7�HmP�Q^��V��p��8A��W!"U�@����������_�,�������R���J�Ic�A���tVL�B�3�
F���kp0�A�H`����g�;%bQL�}��0~�S��|�l�o�7������Z�e��T�g1r�%�_��r��Ha�*�u�����V��yc^п(�4�V��}Z�(�} �
�]i�l*oNd(5��Vӆ`L��3�\�cHɣ�l�i��	 �ޥ5�L%A�*C��)Aw�K?o4�%��b��&�_��p�a���o�B�Κ�zܹ�|u>3�$���*^INaNk���<}y`�8��Ś)������dX�������V!B���o���u��"ځ����+�mF\���drMDCuLO���r�ݒH���F�@���O����:�4�}���Y���ͻ[�;��D��KC��0챣�CŊ�K�ĕU1 �]Z�B�߾~�
؎��.p"��W���4G��gyzmb�^#��+% ��-IJ|M.�ev�"
�J���p]w��Xz�%4���J�H!���CKVʂ�N(�}�� ��� ~.�An�A����/���� 	���!���:Gv@y����� [��c� o��t�EZ�ۛ[��܃�B�Ǯ+4�k��xr*��y�jϥ���!Gq+A�� [SuTE��<_!�ζ�v�G,�뿸�+=ֺ��� �)Wn��iy����)�<��]��Sj}:��Q	�{/y�6@m�G)c� ;
y�����=j�>z�N��e�N�x�/�w�c�{C�Wu�a�h$��֖v�ޢ�E�<(n�f��ֱ�mh��264�1��kػТct�Ao��F� �@D��AcM�`��Ƣ�&���nakGɥ�u����"d컌��B���a�yV�p�=?�#*8��ߪ��)�~�<�
|i���Hg 9�5(� da�g-}���P�[uH�kT7�:-��y����u��W�_F��ա}η�]���d
�2�J	�P��l|�����W�(��t���J�͌K�6To2�*��
��s5��X>�/�L^�I|k�:,���w�~~����c�8��Y��=r�&nr��2�&���lw��"���_E�ķ��2T���-.���@t�9��:��jTrJ����
y�P��z�-uG�Zpʣ��z`y���S���|�����_D�M��7@��P�`1�[�rm���Z^\�{T8;�ei�V˜�y$<�P�+���%��t�7�[Z5{2�ddޫBЛ;e��""��g��#o&\%�B�5��Ā��y5
t���	�j�P-��㞼�י���*����R.qy�Wve��>9��w&=�<���Ǭx�o�"n��LZ����L{�<���������G"�cB`��5�Ϋ�#��������r�;K���C+GpD��-�a,/u�E�!�[B%!�;7��2�Nno���|]��ǽi�����V�Qp�ȟ2d�z�uT��J�zc��� �!�/�RGz�,w8vT"�M.0l���R�2��HC�0~R�%e��CR���k�@Rd����ImM߸���O}2��ۧ�`�+��5�����_?ɗ_���I>��Y�" ڨe�7H��^p��`^�f�����0�����q ���(�O.V{IY�.�<�	wI�mNn�TBr��\>{���ᩡα��H5�M�e$ئ]ɒ �h��4���+��4�//�S��2�h;���eY�UN!���`�rP���鑥�_�V��s�����m�d����9�CIݨ=ק�՚K�<���F�(����㈠�/Mj�͇mj�J�/��|}|a�,*����N�������Y>�U�F����Z�>��H� �~���r�Y�È��|���l�����P�d���'��~��9�����6 -��x����\�g`$�vM���ˆ�U�4#-�L��j��7w�����(q&�]�g��4G��S;%E��w�$4ǽ��_��$�?�P�$[�)X�С�	��4�p�k�$^u�l��
�jT�h{<N��1&����}G�n������ʗ�9c�@�FS��(�0}r�}h��Y��)�Dp�̴�:��� N8<������ P�{��N���{�ݍU'�$�:![�VSEvԎ?�����(tC���z�$ 5AkYm�6�|*Y�PC����fB��c��
P�'�E�=E2X���V����Ԫ�f�i��bKy��^�ط�̯c
�GE��;��H�6�����P8��-��0��2���&��@��Ʊ��p�#v���32e����D�`ߌ�ϝ7��T8���6Ҏl.((�Ŕk5���E)c�`����V�C�(��A�;�<�i����ul�v�dS;Q:�/�L��}s`Z���9�i���W�fL���6��\g^IK\?����ZI�q���wi|^>�g�5'����l��yUU$ZI+����h���z�"Ѳ��w��$��ҁ;_�@�c�*����*ɒ�&�j�����}�v��oBe���4�̈́I{�������d��d�%	�H0Z	��᠍�b�$al��T� ��������(mM��3���h~��4�j�?�X6܌�z��p�:¤K���ZYc	%�
�;���C\��{Ko��Y��F��+@�m��Ү���v�ܽ=o�'ь�0
qdyb`�������tabVF*"e����O9*���Je����Fz���v9O�^)0eӜ�Sބ"<=X��������9��R�wA<4yP�����л2�^ͺϧ�?%�a�G�L�@��ؙz�y~���;��Y�=��"��:���g�]Z��\0Y]骼��5��p��Y)ʁ��wSK��q��Vi�=wڏ(���ǖ�@� $y|�����g�Hr<�ih�>�V���Jo�f�qe&�|8܃c
 �Gp.-%��F�7�A����J�����J;��`H�%ZG�	,�R[qc5^��`].s�F�{چ�R�����:$<&��< �j����IV���YHTM5T;�1��B�P��썻��U�C����9�*�GF�/+���yL���dp���N�������ȳv������HMM�H&|���y�]��Ǖ����;ae,�$��Q�qg��9��9'(@6N#)������r� ��*k�z� �] X���l��1ʽ�z��&�/O�ě��b�?��u��j�6n�F�!U�=b~Ge�g��~�'��\F��1�m�|/�,c^D��H��ʿ�N���!~�rľ�"2��Ld*��?��tD�v]/od�nA`���%�����*��z.Rr`\������?���\���r����Bh��`o���P���_��y~~b����&+*���+9����ǧG��~A�U�o�� 	�Q#�w��LXB)K��ҦX/�7�MbP�'�c%N��lR_��W�38a @\7ġv,7���4'��ڱ{J��ˁ<;�Ϗ$��g$i2����4^�����-�F	z����R���TM���L�{�!Ŏ��ɴ� Xb~�]���ʟ�Y2����'��'��{2F������5V/Rf}6b�i���@9���Y�G���0�Q-s���/4���o�*�PxB��<��>sp�up��ȿ�G��ܦ�~�W���Wk����J�Ce�k��;B�-�V�\��r+M"��51X��-��e�l�NS��c���ie��,�U�N�����T��(�6G�~���%�΀�q��PB��X��m3/�VXxi�X�7<��j6�㐁	Ok��maY,y��2�3͆��}����^�u��,�+*��9A[0�SA�L��#Fm��Hv�K��}k��ƪm��P�^QNxUk/p�>�c;D�Sֵ����{���ra���;P��%B�8	I4BK�{t�KcM�or���Q	��՜G	� ���7�G�y���H��:	��B!�v�!�tO)6l�wv��SD����C���� ���U!GV�����H�:mP�� 0�"��&���[�����<q6`!L��w��cpb��F��o;g $�)�I���z��!�D�((���t<j�PX)��8(a���v��k0�7*��Bik<���Q����:L�?��SO�d�'�0g���:d��0�x��{��L�lfH[��VH� ���b �L��\MR��PM�o�:~�纖�pe�)N�����<>�y<��Ri�8(A����co
Z�ƪ��y+k ��ߓ��t3x'�X���XI�����'���o�tG�z`����8|4�hxCQ�YM£O�]?�Dy�'������H/��+}z������_]!�4� (�6��=y#?sι�����Ы�[b��bC`'�v��r5.ȟ�"q"*V)�X��3������n=�1��ejeDy���I�,e�HVF�*�u74z�k�J�ͱSj$��CY5L֨U
�k!�7�P�g�	�I��z�`i]p��F���b�(�o�vJ�7*��X�8��C��W�������*~��,W��"wFS�D�w�*�L��s2�È���#Ɇ#9vD�ḳ��V�i��w�&~yL}��ilXd�h)iD�ܴk�[�Kcr�y��ɨ��n��"	IQ� y()>�X�i��ӎ��Y:�'Ry����0aE�!�wej���d��֤H6.r�[\Ƹ>z#��hDO�|ŚB�ʠ�'$�i����홖��]�{L����_�� �#�%)�Yl"�T/-8sZS�Qʛ���X�1�b�4"�O�3��Q�m��3TBk��r�a�h��FT	J, ��yT�N��ۑ:���8��U�q��0�l
9��U�B��6���Ĩ����6��hS?��q�~���/��'�V���heզ�=���n�}�_������=�c*����]�o���Ϗ�º�xG��F u�n���B��uG�X��X"�\��Z$Z,[\��|��m��1�����ե�0(/CϊU���f�9H�:��	�#W�� �ȠE�FS�Ѵ�v�I'��C���p���W�����E)^^���Nk�i'�Y���9i��ź	b7y�[�#��r~�sO�?�.:�ιHyP�)ι��zT}����������td��`�DdT����7~�%F�7
Ҳ4�<��"�)j�s�S�}�/��&9� ��~�*o�-�}�Ӛr	���y��R����p_���Q��$gR�FP֥�����]\͏n���
�7�2��9�UR`�-D�(ʎ�L<��Pބ4qnH���Wv�(�;�A����+Ba����N�G<��y�
�2��/]��&{��d��I
�b���b�p�����~m��͎|��?Ie�vY'�{�gm�v��7�3�Q���ʯs�<a%�;4dg�T�g}��4�r9������3�K���Gߑ��j��/}��+��z�b��`�1��N������_JA'�a���Ȧ�G����W#�*Q{I�f���E�ű���2�[CNxcc�vޭ~�IT=m�C�d�lЉ�L��0�_��nM"��ө��u� #g7��j���*Ii��}�-�Zno�ɻ���n�p2wf&��z�h�X����i7���A��:��xJ�����w����y������mk��TȎ��	h��@=�Ǟ���r��{n�A�єE	F
����b�z҃��S%�� �3�)�Wr��:,Y@ב:���Ρ&~})�ū��yci)��F�P�;{hl��`��QtD�d�u�!�"m5`=��l F(/%�CgK���i�w0�)��\7�N���Rzx����������o���d����A#LX�u�f�|k�?������?*Qj������W�F��=k�:'��f�{�ՙo,�1+���	�ݓ�ji�F�ѝ�Q(���:��mZ��� � )�Q�GQ��=�R����	uġ�Ձ����; J�[��$�]�������R<8�3K%oʢa������y�R1Z'7�'�����1$K^�a�)Y�n�#�F����\ɡSPG*��ˮK���]2�4��9|Z��52�'��^ǹ0��B�$WɘUL���sT�D�XE=�R^�^�*��C����m�b�  �~yb4�r��Zt�2T|Yt���*x��tT�����4���GV��4��ȡ�-��Ȕ�+��p�	���3hd�c��Q�ؔY�Ӄ�]5��7%�YIT#��N���-��6ru����HP����U^�^���D���4XJ�Wo�,���2Ĉ,���A��47Q&��G�邨���K�n�� s���Lr�������ސO�; 2�R�V,���Wr��H�U�=��2��XE���U�X����z�1���b}�bZ��Ow$�޿�k��"����'0�I>���������g8������( ��3��U�<�bV�4y 
��kQ5�:��\�^�?o�n�G�JR}<*�̨K� �X�Gj�'��l�Y�ԩ�R˗�����{��F?P����2�m� a1Jqo�%B7|�� _��I^��  D���!�fوh�����W�x�{�K
��c� Lc岗g*X$;]p���3D�`�S�3�p��c^��m2pv�e��8d�@y#���t}r������n�k�� A��pT0�{O��dp��Д��AAz�X�*;�\�;`�Z}&�ˢ,�1B�k��G��@Iy^��ǒ�b�e�r�G��@����>��pL]o���"*�#z
`�5�̀Zv��5��bz�v��֎��ж�#�@�bZ��T>��ɩTA����v��0U�����d��i�C�Twu��1>�΢�b��[�sè5�T'�U�2`�������O��c%G�g�ƌ��GV�p4P�+ ;�\�Xf�5&C\�
����[�F�H+�/��Z��f���&߭*2�v�	��w�n��2�U�Jd&�M�Q]�/��/��/������Z�;���o���X��bV��2����:��:;��&��~fd�toAt#���Ndo!���Su�f�0T�KU��?/ �a�K����q���Y]��=��`<��g$���7� �h�{��!T3i���*&'"\p{���?ܳ4&a oH�M$���� Y�g�B^>��fӡ����^�g�y����%Z���S �<�	�s��}J�e�5�N��k^�F���Ҁ��D?��FYP @���T �t�{8�{��G���`5d&{���_wC��o��)�ϟ?�b^��W�Ԥa}m!O�%b�����	�t�Km�I�2lҝ^ω�G�iP}L���,�j�����}H��N�	�����
���+ހ�J�6&�j^�d���ݹ�%��n<���p�Eh2ta\RE�ӱ�d��z��u$��-���^"aj��sMT�P��c�?��b�Ih�W0�IB~�A=�6;J[Ks����]�q`gt��x.�߳k�%�0+1�'�z�B��7��D��Μ:�N�%tvF-�`�`�t���g��Ǽ�n���-��.b�{�d5',�����
���*T�n$���þ��-1]��k�]']V��a�|=�V}�3�n/7>�����0o��/>�������\Vj��t^J����_����@B~�8��t��[�1�w2��0P,f3���h��VcԊ6P�$��I	jY���;��X����i� �啦�i�y��ks�r;wa��մw
��8h�`�E3����r$s$�|$	.Iu��ܱ7�[+��0G�&Nk�[��p�0�$]s���E���������VT2#��('Ԉ�p�������|v 	J��
�>��=��z��m���։�jNL�.H,��I�𕗦��dֽ�KlO��d�A8'�fRrrx
u-�.	��f� Y�^'�zBE5?#��𻕆���);�FXqO'�v��һ��y�s��pR��1�k�hG���ݕl�������1tN h;J�#{�hQ��	:o|]���o5�8o���e�0�,�*����h��,Ր������� ��9�C��F��co����1��v�:��y���942��X�j���@�kPdIK��4��Ο����w��ek�L��N�cpBկ�ψ0��!#f�k���zJ�uj��R�Nkz�(T�ad�������(��n 2����8�	�P��
��vP}��m�u���~���Bkc-�A���IX)Z{��}�~=���1�hq�3�獢>��s걭ٳ~�1_���z���w�Z�� ���M������1������C�q���>��Xb���v]��[m:�;�ж&����瓬��B��'� �8yz_��;��c5/�f�g�#E��o�ս˽�b�K^pC��#6��j���ĜMZ980%?Tm�J��`z�EN�v
�)�'�o�C3y�qT���\:�d:��H�=��t/�_�A�	��_��1;�3���x$�:��@�j}W���.���Fߘ^�뀇�˷_���y|�gaD9F���1r��T�UYvK�̡�z�y��9���0�=j[R�8>6!gZ������>�������찣�|���}�\B���a�����	��؉�z(f`��Y��@vII�b=����5�R#^�i�aA,$R2��K�I5 ��{g@�|Mz�ļru��%�p{xQVI�^��/q���~D�����'�S��H���P�p�X��V���ᇳ����&��z�����)�hD봩G)N�Y�W{�X��yA�5tQC,�fb�ي�^a4�Myn����[���*��R��2B��Ξ�}���U�CЮk'�B�	-^�ڤ�EcZL�I�
0R%��0f�u��8rXi�'����Vܱ�s�G�r囅���wCV�(�3����	'+�����Zh���(���Tx�C�s.4�ф|��ݿu��=EB���n&���4���5��/^xs.c�ʜ3�\��MÀ>���}����@�����"����E�FGS]~��MW��cV��Mv/ӢY�����Y�Ə����^Β�FUG�dٳ����(�΢!Z#2�gF��D�!��'�Ÿ5�����U��5���a*��2J/���k)���
�y�jHq`S7b�C�����%��A
�����l�AL��t/#	򀪼�	P���F8r��9}�^�-8t�|Y~D//��^�ڐ�ok���a�}�e�)�K.�K�ѪO��ؽ���$�a�"(2��|�>9B�Q������3�<����QJ�VD�4��Q v ��� �9�`����e������HA^�w����<=<���=#��GS�WL\3r�9(;����������'��"�vl�b���Z�_L�bQ>>�BoC�If/����ZY�q�7�S󷢘�.2F+P������8|���É	b���f�>n'���Ԕ������ettN�o����u��d��X ��'ׇ�l�]�py����
3|����{F֑�40�~�wW�MG�;�嬆���XWQ�Vw��c� ���;�oU3c�7+��^��uKbiN�4:�ci^;��^�"� y��*�4��ˣEM)�,#D]rX��q\1���:~�
�iI��HT�c9���q�uH�jj�ܹ�T����/�E�x�Oc<
z�����Ԉ�%�T�7����^�֊��q�R�C��b�� E���i��զT�1�������!y�
W��mW�բK�]K�f��]_�:R�k�I�kv
�N���X=�L��F�K�M�	�<wP�uC�mB��c���{R��5��\���O����2%���ـ(SUMf�NbB9�z���3��i�'�m�;P��qж�c�6;N��k�?��k�p���30�0��A���y�j
)?��-}�+I{�e�Q\�p���YB��=�ƍ����U�>X��O����7�z���o>��r�T��>5����R���	����]�!�˦����$F�N�M��OIV~������A�쌦�t����	ޫ�U�@n����v�;y���7��؉�Դ����| ����"w(�T#�ŷ��?H��1zĎNv��%G��0�.5tI�����c.[�|a>$E	׿^ߤ���j�,<a�+({o&6�m"������!xqj���� ��%�������|���wx��=����V�"�A���m(q-��!zg�g���8
]#�n9^X��q��	�{��#�����l㮈4%������e/;c�mb�#&:,j�qCId:�s9Z��w'�l��[���Dz"�Hq�ᄃܱ��CKa���RwI��)2uż��[W&B.��l����,��������Mk��w�n�Z�����"8�Lb6qM�.H��Ǔ�}��_��1�r:W'�����zA(����ȝqr�S 8���=�y��ҹ��Z]E$L�*N�M�[��,'�V���TJh��)�4�!ϔ%�6�5���U���Ԏ���M{��`Cg��V���2�^��)�E�00PD{/��G�t��>8�u������g�|���E&��ʆ�hzBK��S�΀�ͩ�7��0��6��c�ɚ�L���(̙#wF��uO �S0d�ūx)Ι&S	�����i��?��N{������i�C�KK�?=�Z�3��������'9;M�a�\I����8ǜ��)-�� '�L��޻�I�Iz��ݑk�b۸��G��Յ�o8��W4����r���Ű���2�He/	�aF��iX���<��� ��w���vL��fCW���(�*4��>�<��:q.�� �i?�2�8M�R N�x�I���S���H��B9۔T�Ƹ��r���VJo��VF�`��������!V���i��&~ӑu���<sՠ�oT/,�3dZY�V�lǤkKd�;�GC_yc�t��gc�Q�^��ysl�-�cjG��<,��];��(����o����%�G���J������"5�l~�)��5�����8�����z�\�N.��-3&V��\���c6Z'�7��;��>�$q�&��N7�g�������2�&�l�=�
h�ϵ$oS�2�瞥 P�7�]u���鼪����ZNK�WV�8�Wi/q`ķ��}�� ��h��]}_/Z;��#����쵳�� {[f���΃e�-��I�eg4�}��.�������@]џ$�n4:?�7��=1�{���/�D�ĮiL�� �^�����nN�s���1S��C��Z��8��M�_O��O�AR�<$�OB{�`����z%T�mBoa�S�g�۟u�U�=gx��z �EìI�����:��{���7o2�~�n��0·hFB���J�} �ҁL��d��C�(k)RD���$�i��P|Q�!���qU�M��f�������;TKn ���<���B�{���K����|.z����	��
*��Ez���+8(WD���i˫��e3�p�Je-+C�z������`����l5�_u꽧G%Ԟ��7�1��"@=�+7��#MB%����m�_>v���+�P�Y�܀�\Ea�����+�*�:i��Zy5���T��(�mS=�����X6�Y���g~߽���l��5z:��,,���F&Ϯ�VM�.��1At#��*�:��B��X��x��;F���M���s�q��$o����W�u�J!���W�G�X�L5m6|��߲[���9c�vO���fD�h�A2b���5҈�X�ʘ�kZ��`����wƻF��J�y��Y���� 8�E-zN&�m\�感_MJW����o��7�����q�s0��s@�忷p��6�e��^�{�ARo�˕WZ�E�)Y��%ϳWP`���9��;"�z=F�`k�ޟyO]GA��GX���W�*�
~!�D3F�XT���{cr
\g{V�Z��ީ#v�
������a�û���w��޲Z�~X��)�u8ЈŘ��:����F�����v��[#�E%�\��;X�qsr�c�pǼ�z��*:�vmu$�{y���ޝ��K�r�ԗ#����/c3���W�j��n���l\M�m������K�WXI�Éx}{#W�W�V�w1����DO+�H�[��#3����x��l+��S�3#0�:���se���v���Gm��w����";wi{'��,�N$�n-2J��-VeC�#R�����UPD�+PQ0��
Z�s�	=���}���fz�x�F�����^�2������1˛��ޛ^�G����S�!\\�b[Y<��|G.�-s�W�IFg�T.���[G8�k~Nu���A�<�2]�lG�Hh.�=Wb��U�(��t�ϡ8ak�ܼ8��윘��7!�[C�=J�������a��-���M�Z��̬���+m�8�\t`M!���f-�e�y	{�i�V�e7q"R�;h4ʥm��O��L�����|Z�"�M~������y"n[�����7FVL`��g�S���E�v��.��2�3���_�&��o��?J�}�}H��,Y	{ ���#�[H�К���R|��Ŝx'���.M�Nee��k�6�-H׮�td����˯�{�o���`�����n�����6��vK�负Xt�-��v�%}� ��2|����Q{���s<�@�3�P�<%]/]�N�[��_;��
�uC��㞼8������~"��������όh�h�t]xHƘ�8�:��	�������1T����шIO��d��$�Q�M���
IsQ��/��k����m�&�8�8ϴ!����p^d�:�f@�6�w:�G8U�k߭"3�]UR�_�jP���le�(�%ܳ�d��a�Էr�2�)��J{�� �0��Ƅ����ڐ�!�}�'Uc) ���WkW,�P�6ԣd�[*S��� O= �g�����_u�6��dr�7�	u�v�){�V-�8�`���X��xE��sH?4.�q(e(E��'ʜ=�����g��g]&�l�h����È��i�5��yVF1B���%N�iX���0�:W/�iߞU\���.=|,R/���૦9���^�M�ԁ��&QJ%�XW�"f̍�2r�)q��97G5�z�+�M����1�˽Z!�킋���,�~p�ЙO��s��9����I�LȎ���5�2��8V{�=g�A,�< #,Ր�E?�cD�Ɉ�4�I_�^��w����؍�/�x���/�:$�f��3˖�&-�GVZX�5M��L�����9�|̊������=wd�Lۏ�m�Dx�BA�ZC�<����7��Q�?D���m.'��U/�jrT��sW����҇
���B(e�!�F�|8�My�X�g�55�B�K$��G��}��o?JK�P��%qra�+F'� �w}�"�7x��c�7rq� ��x�g�����y@�ȯ4��Ѥ��e�/P��ՅǓ`�r�K{UN]�zo/�yj<=�C}�=���I�T��N��F�8���U��EB��l�Aj 9���ɴ�{�\e����۳����=�s���s��0��M�ׯ�.���O���+��8����׺N.Yw*���W��=�cCݭ���=!G��Z�K�o�>걛��Gڟﹳ=�m?�m�|���;0�O�j���>��}�uEj�>뮶^����$1Ǿ��Z�_�앐�I53MI��X�s����._�|�_?�U��o�nY<����N _Y�Лb"�Rr��¤?F.+���#�]�u�BN���o���x7x Gc��Ð��n �����J��h�X-�=��xlZ���\����94B����[�"�xc�T�x����ӣz1����C�sr?=>���7���#=*Mg�NӖ�DEG'N#.�@��礆{�E	�Xy#�%0o�9���Vv�Gy�������Q8F����?�@��X��|c4��(<Ih�1� vP�0W�W*�Qe�.)ɧsorL����47l*9[��
��\jzx�	쳳���ʦ������m�m�Kc��sAS^5�Z}���3C�#�B�%�qp��xB☿�v�����6'Xߖ�z'�h�\Ou�V�dE�+��a���ǹ�6��|����XH.u��b�Q28*ż4�y:�w�%��e�i��jܳ���kȽ;1X�Xs�w?pT�P~��&/�n;�t�q)2�k�IJ�W4�j�o+_�Eo�@^5$�+��z�
�:l��y�[�	�����7���|�Ty*{�<ՅOu��=�o�r��+�ﰅv	p%f,xJ�+�Q9N�*�{V���3׏�;1��ƒ�`���6yn/OG	�������N���ʚ�~��ҍ�cx�6���2%�����Q#B=Y}Z5q���d�l'���3@r�$Eqs�%ɷ﷌QS+��}T��@^D#�b�(p�@�k��6�1hE�{��d�9�wf���	s#w��_��{"������x�6�
Q��i,��R���Z�l8�x��3�
�1��w왲N࿷Z��)܋�xa4U�)�K�z������\eF�J���>��C����	��p�熦E�F%��j� S��C���ģ/�;Ve��vF��J~�e�gT�{feT�F-�ۈW��uи^d����B=:>u�B�������
ؙFb���'~K��

!�*d�vI\d�T�w��>u<ř>5]��:yko����E5J_�,o\K,bƯ7���8�J�&'�9�{��>?N����B.���0y��:!���������uh��R���ߵ���&G�E9�sta���u����g��{�����e�|�t����k{C�]���g�v�Ӭ	_N8�"�Y�;�;����x4!tYg���f����QvI���g��lD�%#��S�<@&o|�1]-�;�!�k=gvH$�)�Z�3��ٽ>3@�*O/��=��9'��^�s�rpV�7k>b�U��7����#�r8:Uޓ�:r,�^V�B�e�R�\"�	��a0��<��fP�V�r¤��F���l�޲4ʀ�A^�X�5��iN0�A��I�￤BĊIq��%-=5�Oμ��g3���4��Ϝ7����U�4�}� ����W�_�����/���H����-�8B��-�3�,��-�F2�N?T�̶��J�+�"���O�2��u�N�[p�z؊dj��bN�_��n�#B�^umڳ:W%p��8+���9��Jj�j@�A$��r�9N�T�̜��F7��{��,,�7o��y<�DS�I(s��Z�$�'a��+6qrᲱ����v甑sG~��!��Q�Q�${�����P�S�gMx\*&�3��^�n��_�6
 ���;�|�ߟ���߼����S'O>�/��Td��+HQ�P�P� '��w{	�>ɟ#�D���o v��K�N7ߴ�.�1yG��1�����ڡ̣ZW*�nJ�hV�d�m�\l<]A˹����+R�T;X|�9��{��������|H�C���z�����yZ�ز���r�.������1��y�S毷��(�����u.o^�B�L��Lq�|��J�Y�y�JRzM����U_\�����.U�1�^�!@�$3N�;<���F�v�Y��=KQ�� �gu7��ncӪ>2:��5N���
�{� �� ���K�o����êѽ]���F)%��'�����X�Qk%���T�q����q����Xj��g�#��s�E�9�NC�}<0��U+���R�E��k�/_�ӥL8v�����i�G��N=��e��9pDj�D��B� v�Ǖ���q�U�e�G�>+�A�t�x%R-�`<Ƀ��� :�T��h+n��?:�s�NN�G����0�r/�;�'��߫~T���ֺ��R�"Z�N�/\Ǿ�z����s�n~�z>�Oԃ��|�r��#�?�����rz�z��A���+ˍ�9&���=m��rz�����AK������?*}�{������e�w����l˪a�UDg��mGc���L�jڬ?�����̝ⰡD��;�{s0�6���V�vwy�������>m��Yw}�)[Z��ʶ��5�NQ�����L��X�P{�����j���yI�/�_�ׯ����#��#N��HtpH��w�f�!�]V���63-|�l��:����r����������U����1���jҷ�!��� ��R�� ��t!r��ׯ,
c��8�G�4�_Y����;[�l�	�5á��h��y�u}�ļq�3��F���bU�f���Q:{�@�N��t/��������� v�ҳ��4�{%��Vqa[�F�����B���Mk��������qA#�G�;��W�c�l�5���|��R6��g���o��곢4TJ��]]6�]�W(H���X26ꙂY�T�4����j^��wc6�Z��X{�ɯRZS5�ȓ�{��~L���3Z����yp~��P{��Wes2ʩ�͔�e:_1��~( �E`�_���L{�ʣ��|"�������*`j}��<�����G�r��BM!ܱ��9�+��I���%��F�J$�O}���U��s��I��[O�y���)c�&����U5+!;V�w���FȌ�٣6��+
=��2�$�	Y��뎮�����5G��^�������E2mt��?���A�q:�E�T��OZ+j��u�K5w�U��z��;�^;)�:wY�>����s�p'q�L�+�̜~�U��У�1c =�N0g�Fn�� ����� k^�i}>y��h���yf8�A`K�1��(v9b}��>�R*[���O��S�ܥE,GU�a܃�:�蟣>��4��
#v�1���
8�(�-�ҁ�[��g�����i4u�ht����*N�-Y�?�޻�q$�4(��#3��{zz���������Q]*Eh�`����U=��|L2H���r��uF�R�'մn��<��1m33P��Y�}�w㚰7y#a�x�C�k�@�g�EJ�+%p�����뺟�u�5��� � � ��s��q��D�a�+��<���vH�Gn��8#�|Lt'y �|��$�ߡ(�|��@�P�>���XvK����g���Zu��7��Z�&�J��*���nVuR�u���9��\���Ɍ�(
�W��!��d	T�=�*�t�zyy��_9ΐc�ʑR͘0F��}r�ya����rɿ��k\�VBſ�Ü$�ǎ3G�N,:���|�!�:�i襃��˫K�~���o�.f���%yخ�ly�����P!Glm�h�����(P\'ӣ.�1��j�MO�7�W������{|}�WL.8�r ,m�;������@6�����l��%�� x�'y�������4�$J�6`Z���|�� ��W�=��q�7z��e�B��=�$�A���|zF�lz�x� ����g�V��������g��7 �ч�;�x�>}���V��s��,U^�w���S��w�0�t�0�(������O�����������i��-��cs��Տ˾��^���8{�ڏ2dd�C�^I�//�^�鄎N� ��U�3%C�0!u!���@���r��r���3>r�L�Qb���`kL�.Z�'k"���ư;u�������n;H�NNBS�6�z�h��G��4V�e�������P�A1�ؽ��Vп��hĸ`^V2Rc޲B��5�o�=��B�6�e� ��2��X�a�O��]�z]���t���+������*H��UW)er��]%���, �����P����!�T�~�� c�NT�V+��L+�6]9�>�0]QÎ�\���	$�U#��$�
Mퟛ/wa�]���^�@d.�!@�a�ݟy��8����R���Vn�L�؉{������$����.;�v�4U�{��^N��P��BS�KE��8"$��.Q�6�3heb �()�Zl�\S�Q$�8H&S�b���bd:�J�ޣ
a���B��::em�螅��V���	��fHlI�j���P�<�ѢW���/�K��7��y��������>��w�тυ�!\j0װ�d�QN�F���ǅ����[��[Cr�I��cy��U�b�����l�jPFSL�4ӝ��7��F1Gq�Vk�Y��),H_��/f�2	�$NRJu���ă�yW?��h� u_�2��/H�P6���?c*G�}�=��ڙ�x��1UZ��s6<|O4#H�^m�>m>C$�i�yD��w�����S��R��!��aW�$ڪ)�	e�e3V[�b���ǆY������@�]��I�eR��A�C �������Q�0�U0�U���mi2+dHG/�)��ǫ#�{#��ʊ�80V�W�{T��:#Q|�֯D��@������7�9h!㕞�1�@%�uo��'/9ubO^215/ظ4tZ)�U�&���,f�����x���xA���Й��͇�`��X�C�Q�W�,��t���`3NY��;���F;Â4熳v�d�ecr�����9��ݐw�z����+pƭ(�9�ju�Y[Ζ��)��$�@"K�Er��LON_�k�z��_��_~���Gx�_�z~��0��"�UTq�i4Ph���ܣ��̑��`ؖd�Dك �qTG��Z-潌��`ɇPvt�⤣#���>�~�������ޮ��u��gxzy��-���0�W7�9�z�)�f���^-����+U��g��
S����m�΂'+�n��`�4o��͝6,��L�y�j`b/����y������#X�����?����Op�xO)"���]/�pֿ�l:�E`w2z��R_6&��p�C'���o�� �ۍ��)h���,�Z7-&gN$��/6�$ܛDHK��B�+ܥ!&/z�P%�o#��(�Pi���1����Y��? ��:�{1��?̺�A��nQ�����4Nocl�d�I�or��T����Q�-�.�+��xZ��3���N4H)�ke^	9U=rf��%�a�Y$Vb��I�P��s���da�ʗ4;�x�J��	�L �lM��j(����G�g�����4(�pp�Py���Q��Б��^*q����hm*O+yyg��$(� �l��=��QF�yDTz	+HT|G�7�NDQ6l�)��k�̌ǚT&�92F�+4��A��)��qV:�{�����I�&�G\���g�/��E	�n�T����ޘ��:&���8MHtcS?���u-7�|p�`F�t�N�qF��Cz�K�1��� ��V?�)��Ng���.����q��ǅ��h�eCp[���#�Q� <$��uS�Q���-���*Jȶs:���Ly����K�zTY���D�ȡ>ǷG�"��i.L�	oj�4hH##Ak�tuQ��Y;�_�e5�PD	g���+��=�ʺ�vHC�|�rC^�{N��Hk"8^\��!�����/1����.�F����;Z�Q��Ӕ��:�s76"�2q/�"�z
[V8�B,"1 ����*>�wG�:`�K�L=�R��x�b�2���]Ue��n��ْ�Jy#+d����i{�ώ���]��.d�<{w
j�X(�}�㻬_�]Ɗ��Xf%hb�0��%P>{�*�{�R�ڬ��3� �n��]ph  �񾩗��l�D��๸P�����lF%�I���ikF��ږt�	S
�3�*�|Q�E�3:�N&��8�~�.���`��o��2���ˈ�=�$��@`����ǋ��G� o@:�����^�]RP�L���#MOÑ�]\\���<�"��#�L^@ ��\xrO95��!�� ; (������()@�2=����m�
O/�����|���J/��>B~u~~&G�;�!@�R;�4i	���"�(*i��e�3�D>x�h����Y
�f�c�1N1z�4�fydY��/Ί�t�򈙭�����\�ֻ��S��S�Sn� ��d�@%�� !aJ2�t�Z��$'v(�S��~�)�nϓ���р��� �/�����r/f����i��S�Ŝ�f�F�>� C���Ѩ�~&\���?�������_�o�_ɨ���^�p{uggKʶp!]�)����L߆aj����P�z�	C�E�zq�㏻��+S��z	ʫ�˟{�Sz�Y�#Zߘp�6�k6�G�_�c��r3��fLB��'�H��,r!�꾯�F�;�(�		�z�GM��(<���ci�Ep�L�a���A�_��he�00r�`��f��.������
ώw��h7B���i.O��}�!A�� ��J8�B�k���R���fr��0��1�.y;�(&�2�tqp���p�ע0Z6/��.����HhVO��K�Hg0e3�G�N����P2̸R6_��1� ���>F۩�b����^H���k���a��tK��	è�?q�3�� ��R�}`ڑ��5+�OEE��Bp:��m[ݻ�	���+�b���7+�3J�tς(R:yvMa/�-bM�B+T��.��xB�<�P��eh��Y�x�@��ǅ�W���QtG�?�=��B,�G$ˡA������h���a+�����rY����eWx?��"��`#5�-$�n�Z�O�+&9,�L<���棁.�a|���0v�ӑ?��V�4PЁ��b�F�؈i�ZMP��$��,uفЀg�c}�A&S���!>��"+5�@�ٌձ�Q@O���!�-�h��k�N��_4�d'�"�(�u�g7�py0���c������<*�i���8}��R�-���g�`�戆�o��i�jzuNvu�����L��5[U��z�[�"���6��H�>~����֩��փ��{x��yLe�5#y'�|�\!����i�k���^�̄�#e=��F��s�J�^��߲@l��&�d
�D�968�֐�=��it����	���eR��f�S��a�d�]ֵTO&C3��99lt�_����H�/�5z��H�Bc�~����K�g�g�ҳveX;w�[x|zb=��S�������l�2^><�uF� �J�$�؄Ǒ ]:��	|`p`�Nܬ%�������+<�<�S��0�׷gxۮ	����Q3+�bg/�H�v�̹�����rzA���K>P�f
$BEA�g��7f���T%����Y_9��\]^ѩ@x}�-v赃74z��Rd�O[��C)��{Ύ�삄�:�����p�K�4 5���P�O8�!a:�ŞB�Zq�b��-��]��H��ƄLM���"��J����/_ᗯ����?�?���Ͽф��f�\�e?��k�/���^N@f�	 �o�tX�F#4����ڈQ>�#n����uT-cR�9V�*MH��r���<HF`�+iI,�������8������:	I�ORt4u�"�?3�/�����.ߒFwE��CN9" �k]gF=�#/+�%P��ͅ�!	�1�f�(m�,I�$K:��� `�~�/S���SD�1<=Q3P�?�ɖ��(�����1���~�������"�&�"�c���+(�������<~�8�eO=R;�e����m�A<ͻ��� ���(���'7ُ����9W� 5�D(�m�t����Y���ˏ�i '<��(��l��n���n��y��G��]�
��e��h�}^"��D��&| P�ܲ�����k�Í�i~0�a��ZUt�bÌ)��δeX��M	iR�"c R6Fʺ)}Î�0K|�ZI(E9�q��e/�)c��yc�n'�Î� b�l��KBToO�jƵ�]g�揻N�5�3��Ȓ�W@���m;gةV�~�3ވq��DC�ʜmiB�~6
X
u�4`�C�2����f@��I8���B�"Y����r�:��������Џ���t�Ğ8d�Y��]�9T��w�	<���V����	��`X�!�eW�99���i]p�G���l0&/�9(䡑C�$�����ydϜ6y�7m:h�{j��<=rq!#���?�'�7�����}l�#xf�RA�����G$�c�f~��?�V��ɯ���Ưhl�������L7O�]��u��lG��ρ��7��]S�\�m����
;�d�#H�w�i&�g��N���k2�{���L/��p��N�[��V���|� h�i��f���y_h������A!aKϖ#X0S%�wuuE�&����̓t����,/}��
�>���-;�.0gQ$̽��R�wl�c�{ �Ύڶ!�9փ����~�߾�BƜ�����E@����w�/����8�9֍v�8���&��3o��u��CC�މ������-<�C>g3!���-�������Jґu���u��4r��覧"�I�`�N�g-hB�b�e�A1xv��?d�A�Z�C����gxy}%�a6�-\�_Q
vD�2��b?���ʆ�k�+�R�n�/�����8!�=�u�tO�rO�g�L �:0���?}��OȜ ;����Xϖ��hQw4�hú	ʰ`�C��c��7�}�	����T�ߙ��5q�& ��@���(S2$'G3&�M��F�=Ѳ/�aG٘vhM���E5�D]��Ԯ���Twфz.B�����[�g0��Z%�ƹ̓x�g/�d�͊�@�1��^ø@N��4� R7��9��N׀*^��	�O���ᴎ�yt{�!ӌ;f�2��2a K�D���&j|uj_а�b&�ML
kLLZQ���D0:nѽ��G�0�E.�/�5�Ӵ��(����F�(�e��JaC��d����޵�&D󏪠Q1����~�A9��N� p�LwF�~ �����P����YܚV��.�8Xv�c>p8��HT����5���*�/��'�v��A���=������e�H���&�)t,S$RC�?d�id��oM�tb�~��vC���&�Q J*o��d� �������*����"z솆7+����q���QE �X� hR����	��r���5�PB�ըcJ~Tڗh`<D3�$a��,v� ,i�?@ɀ��m%�����K�k�?��y��aYd��lM�˟�_�����=���@���y�>h�� 6:7��;	7۾��~�2K�_���61+�l��ϩI�C����� �_Tc���e��IF������F�{�C/bL7ɷMt� ��w�λ�˥�1O�0f��L��wk�����j���$�Q���j�������)��a��X_>Hfm��!��$��1����eO��x�v8}	�Xe�d��"�Ƙ},���ql�k������>�������}��K��k`ޏkuc�ayz~���%�/8b�B��ob��˫�=�{==_.�z���O$S?<ܓA���3�ݼ�>��=����������wt8aOˉJ������{��Y��������5��_��I�|#!W|�D��E&*!��\�P�~�:����F{4n3k��F�t�� Ӽ�Wmjfv%�N�z�- ��<v��E�>�����Wx�;\�⪧7nf-�c����i��a����;	����	<zw����<4�l�x��W-��������p�@��L�*��cfB�5�'h�k��NX�������W��_�u�F^;�o/�~�o��d���C�ւ�]_��(S�x�)2�;�l��F���
���:���D��b�	�QN����DM='���J>�ׂXֽ�y!J���\p�^�+��$��5�]�H##����1�A����t�wt`�a1n��
M�$R��XE��r�n�
;�@��(�2�"
�����\2p$a�)��8k�b �A��~�E�0���&c<&�0"�!��.��I��Z�T�w�}W�6rC�K#X�C����8*h<#-��X��r�f��h��|*]e����ZUH��M��~��m	vWrsǓ��֚�\X�#�p]�-U�I�r���e\��c=z��8�S_ޓ�����&!ܯ����bz��mC?E�*�����#���G +�2'x��l���V�d��M��0Հ�]��O�?����g:��,J30�a|�</D ̄B�ňe�*U�b���Pa�%�I0�z.h,��9�Ja�T�3+Qb� 6�\;���ma�_��.�q4�X��x�r��ŞJ�R��:��w�T9҄ ���V�u��l@}�̃'�A���(t�l�c4\�xL&�C�t9�L���.dk��Y�3�"{�:Q������]:#����L���x��I��ɺd�"|��y̳ٻ�I}�*q�g>3�j��k+T�!n��'�e!-'��%c��/�G�G7y��� ���h|�?���9�1�*�̚���8�8hb�Щ�N%@qq S�z�5U6���'9y���m�����q���Q���E�����b+�+mJ��B�ɾ�H��.��~q{1$(�mu�+D��gm��*�]��c�g�=��}�v霅♘�;�X�Z�J(>� ۗ|���r����/��z�&�}��$J<v-����_�W����Gj�Q|z�r�ȃ墽C�.��ᢿ3P��U���JCN+��x;��/���Wx~z"#b侬��6���:};1�[pR̓�� N������vО��)>D��hsҊa�p`�@Y�3�B�$��4�隙KU���9�vn�o������;0{(��oV?@�e�����16�ٱ>���M�T���X=�U���ųe1�����/}��v�����<'���!ܞ�������m�d�y#��-�)ۉB�������Zh�Co��s�ӟ����?��Ns��'�/y��ek��`{���/8�z�,[���҇�~v����B
؂�,��3؜�Ⱦ��.�r�ob��[�@�߲���$�٤�S	�S;|��ƞ��˙�˜h&���BG�\Ԁ	���jE���Զ�y%F�~��xc�ք�v��y*\<�pӡ@�m_�6z*݊Ќ^�"�u�Po&+����KH��2��|�l�הX 9�xwZ5ǌ��7z9A�}U�Q��ֱg<�x���3) �b��  ��}U�J�r���k ���(�
*�
 �I1BG�����3�l �1֖�P󞮌>��X�]ֵh�Vů*��l�;�H�z�IaZ;�{����|��?��B~c�^״��!�|,�e��kf�J!�>�..�B9���BW���o����Q��s���|���rw�E����⥬w�";����%������T��ɑC%�}E�5�3pi����A� ��-݅ Ȩ ��p�$��,�3�g��6�F�54H��40��<^�ɶ��~e1V�f�p��+�k�ʖz���$�u�]��v"� ����/����XŊO&uF�D�D�{'d��Id�����7�)Oi��@p��}BV��v3��@��� �=���e���<T��Rub�~��m��x�5"�� ��.�+!��	^N�V�2R��C�ޖ�.�B��xH��z������k���_��ቌu14B3�3�d�����������o��AM����C�~�ސ�IyA'R����3�f�u��X�+�6+��)T葄顦e ���ʱ�d�B���-m����{�+?t�rwH4�<��VrƩĹSф��$�B4��&��b����ʘ<�ju�^�ZP��Nx)��6�ՅŮ=?[A��%P���<l�_�I�F���aY��+2�`v�����w@bt*پm9q{6T�n�!�7��X^\��g�_�\�ai�\@��,���b�\�;B�,�K��`��>�טP���3���d�0S7���e�~�R�����NTHB:�m�����nn�j�F
���5�q���l	7�}�$� ���|��q�<`�\A?������>N�b�`���o)nN��B�YC�I3v��''i����b�Et��H�i�6���F�p;���p~}I�RO}�=|��_���מ�F����?��׿�\�_�u?��5
�o��ʇ��2~h}�R���ݏ�BŔ�h�r�����RN�Щ����,;��0�S�x�C�YH&�_R8�Z��v�*Ϡa���l�!Je̀E�!��>Z)$�gq¤7��ՓY�;a�* �]:�xs��ӄ�{r�q��7ԅL�U�7�=�Р�XL��ϡX4��z �C �!M9��1U���w�b �"��>,*�P��}���T��
� �ݕ/�p	�B��.��F	��]rM=1���I��^(p�����k(K��e�@=�i�i�n8m���-щV����^���|n���&�|���E3�`��Kō���EWmK�֤M9ڕ5{Z����)ڞ�[*��z�]��󠟳/�V(���1�>&%o�x9�_,��$��I�VA��N�{�!�C/���^0��7B<##+��$P���덱� ٜ
`L���~�4�1��6D1�a&��@��-��`�|�X�"�1�ɻN���&�N[ײq�ҰO\� pSk��)��veV�#�	���[hB�F���_���+]
�;P_�>�V4�M����P�`���A����ԟ�n_"y5����̌:G������YsAZ���F��xO�t����;QWC�y����`�37����ʲ��QM�!��Sm;|V躅j��0*F��(r��L��P�z�q�v�b�25�5�Pv	��@q'��*7ũ���S�iZe/xy�H1�k�I���y:ho��<0+���+D��9�	��[Ĩ�:t�KRT��Vn�T�r^���ć�����u�6ʃ\aE�G����p�vp+���)�cE���`�K��+$��f?*}ID�g����LÑ�L���A�"B^ƃoz���+�/.�us~E�1���@�>�<�-�f�Kp.{����&<�_������_�(�	�y{{��Gh�yY���l&�)��@ ��ո'�I#z�f�$]��w34�-!n���^4:���Չ�w�Ǆ�]�����"��.�(+����(��	rί�+�amh z[��F̤���x��ef�m�0�	�r��ۋk��_ߖ_)]7��n�����![��ę��v�(�#�#м���_^n�S�����P)Jq��	6m,��#n�R��BW�팖�rw)�^X��I���E��n�/d\B���Q`��Ū��G���˟�?�~��Պ o�'2B�N� �ݠ�֬\�#�ڷ�R���h,�����
�'�`'x���"�p�1?��p�*��˓���TgH���~.�c+u#�J�b朞#���F;����za&�*�g�iO�|�i���4H�
�f\	�hig���Ȩq�dRך�N�pa`h	��ja0�k���$�`1�4+�MY���K+�;&��W7�0]Ҕ�7�p0�����ݚ�Fsk.nrrQQi���	���s�r� D���X�WJ�6O!c�$7x�kL/-�.�Y�w2H�o`Ś	*�G�lzr�RoJ�n2Kpz��_k���c6�!�WꍧA�-E�}��ݨD���[�>��~<�p����{��Owf����Q�rJlJ!#�2�O+�B�PF�+o�kLteP:���C7�n/~N�<&��c�\''����tP`E�.�7w*���d��',{^��Q��TT�հ���A�&��ST�� c��L���48}�gA�JL�^fn�����JR1a�Y�;mM?
?���S�{��}�nt,�TH栒�P7��i
�":���7�Y�)�����֬�B�y���{�h$�� ��`�kH���La�L��cue�}�ʯJ�
e����d��=8.ӌ��%��<1��+���#C0̇�%9D{4k�7�s;��Yý*&����P�	� '���l.�"[u��,���)�l�5ҏ��d�p��7[�y�L�S���۽n��o峡�sX�o��+�mj&��`�?g}):��K�4*�ֺ�tπ�.O�Ǯ䩖�nef@
y��r�ӽ������:ǗCg�&�ԩ��{���ݾV�~/�Q����ڥ�{����	-W�vu� �mV��T!S=��m�t��bO<���P����ۛ;J�}��?��=�$Och)f�܅-� � �pwG��||�7���A�Ѧ���������H��z����4N!����ë^�����@1�B_�2S�L�q��mK�/����p}��O~��?����8_�d�Z�a��;⒌�Y�}//����L5콴���3:<c�x�@�g��)Ơ�e��ۋ+�����}��"��䑂7�9s�Y�|�!,���c��E���o����"1TŢx���@�`h� L��V,�5vF'q{�j���A�G�S�ZfYmpVW�� ���<=?�4�9�����	�ڿ�ֿ��KX5�^a�m��p3���Î-��%�<G�d���}�_�w���[� r���G�	Íf�/����I�	:c����c�#˪.W�mo�d����c��}�LЭ_^��m�:#��6cJz��'RJ>e�~��m�<r8���U�28f"���;��)B�oeFM'��W���lt�<��\��=O��T��b�	F�>0�4�(��y�(��)�֗��������P0,����{���=\O�T@U`0/1�c	���+H�քf�2,��<��$!d3Zڐ���g^�тtS�ߪ� R����\�*���;>k^n>z<���Ǽ�!��Z{�T��c�u�m���/������2w�)�I��'������N-���|?Qh9EW�Z�*5��>f���耍�1)U5��L�^���{!��O�UIIO�W�1��In�]Y
ec�T�jdR#��r�6h�[c�4`�=�t�WfR�j�W�s�M�i W�_dPW]�@�eo���u�B�u�{����ﻲ@�~jV^L��X|�ND+c����wW������#���Y� z�,�Et]�m�=?��[����-�����˜ݫ�Y�	�!����<t��T�c��c-(F�<���d{5�-��'m�E9���sg��H8~Odmq; Xuտ�J3�[�q���r����eXt�V��-�&:9&�HQHlۺ}����|ceO�~d� k�ѮJ�R��?��;���ϗ2E�O�}���"��cdr�e��FS���8���ء6�����"Ĵy�>���(����.�������mqC��û�ap��>lI�D'����¿�V��s�����6o]��ZX�3���Cr!C
~F�r&�VB*�*��&����ra�l4�W/~�ۭa���L~��W�c������,�z�YZ�\�g�>e�YM
����m�d�z���k�|Y.�d��w�򩺄��Ym���vuv�n�o��>Sxf�x\qF)̫�X.`N.Lg��(��|������2JF(N;����k��j����-�!��2.�b�h�/A��e����d)�,CL	�x�e�kEB�رAS��Q�o���~�di�`�(���A�A��[q�>��؇���o��Џ��|��
OϏ�
�.�
���Z#9���g;l�
z�v�`g��#�{A�kF�D�1e>� ����#��OeD�p�����H���ө�2F�YǏ�s�oC&�8�2�Ƭ��Y�%�FTe��N"� +����)y`�cU�����W��p���7!�z�1g/X�L�h�ᄪ������w�VeҪ�f�[,0k���|�$� �c�"�P�=68\�m���E��h�_|�I�,��8f���b~{�ͤ5]�F��;�`V��<��1XM�8��w�w����{؜���a>�o>�֜�x���C��h�M��(X�J`}�<0���Sc7�tQ(�a�Uİ��P LhL�F�yJ��yf
I�œ���ae��EwP"y�e^3Y�ܪ��L��LY:��9UV-4$�;�$���4m��W�����?Ra��L�ē~(iQE1)�-x��if�����1��{���N�1�/V?�a���v�Ʃ��W<���Ab0��kV�F<v4;%[i��IՃ��I+m�؞L�e ��t,�Ȉ��W19o�����eơZ�ab-�S㠆kO΃���#cy@����1�k�����QX��OJ�u�~�@o��gu)v�����&'�0l�h�n�CgT���\tS;R��l�e��i�T��\=H������?��+9s`�:�\�z8?0�*���l�\Rl��J�>_��.�0[pX5&,���q})9O_w��Y�#=���#|W�@I:x>ӉwMӰ�
��{�����[gC8=Jv�<������'�����rI�:��B}�0�g�&;�[<��/Q~B����gsF'��UK�h�	�Q���f��TY���]�����5�p���{~���qM��h���@F����a�@p$ȕg����vG'y3X�|�Y���3<��6ɪ���KPك���h�#W�Fۂ�Id�
�"S�E�i�t�r�����و��������?��/��/a���ۏ��^Jm:΄E�^@�i����\4��5�?=���a렷���:��QK��X���v���\mN�-G�(��Ǌb��I����ڒ�Q#��&g��?��`�������J���Q�Zb�N�1P%TL����g�B����;�f��L���I�**U�jd2���wC����'����˔��=�-U�S$�r��>����&٨A�7���NR���ek��\�}v�J��$k�e̠�H��z	&�N�I,�J�g홁pd�#�8=%1[�'���f�+�ߩ%�=��,��%�+�+���rD��au�!��e^L]�[��ddE�`���C$;a'�z�Ũ^C�E��Ӿ��Y�)B�g��{8"o��O���E����U�퇘�S��a�(ph��W��!~���Og��9�WFl����oԻ�䆹�q�S��a�S/�-S��|��[Gl�lw�Oc-|Wu%7�{���q@��_����SXrd��ڷ��)7"{3�������)yxr;��5i�٭���ʻ.�p��w]^v�����Ƶ�_v�苊:��aj�O��rc�����ÒC�̉�b����qy��#Ɲ���3잉>�LP�y��r�����?e��J�T��h���{�9�p�c��~�䙋gE����n����Kf/�6�5A��!�Y(�@��.ĩ��5��%9\P��v��F��	cz���W��(ٍz��`\���h�.0顓�=���b���
�������n>�9�8����S۱�=�����{��J���2�$F�7��u�bR��8[�_�v�j_�Ȅ��}�����]����-���m���2�da[ �����sp���n�Q�7�] ,�c�~r0�;�#���Q�gLW�歗���I��Њ[D��pO�~�qxx
.�;Y�j�����ß��$\�ڹ�' �}�/k��͞,��ҧ��{�*;�Q�����y�ɣ	����k?�� /�	t��Iܳ����NM�:�ʽq���D����X(R2�d�EHR�窑������0d:�¥��D�qQJ	b��T�FpF��_�)#}'i�:�%)��b��'��$=	��ow���{#�J#Fz?� b����U,�~N:B�pM$N��^#w�g�	�)�'H���!���y�z�r��iD��P�m�%�T�s�HЀ��n���AO8�;����CN�{��}W���45R�p`��)f�\�1(���y�❮�6��Įa��G��xe����A�6Z�mBÒB+�lT��{�-�x2��NN/ƴ�ĳ���2�ٴ��J�!gK�4��u�XčӖ*ƭ��P(�� .�J����2V�-�?ʏL �[*��؈�4 q��ꏻDM��U�� Q�=�S�w�pw,>~'���Z�*++?Q��ݬ:����������$��e��bp�?c����]���	m-S6����%g(?'<ά���b�!��I�"xd,��J��K�S�ڐw)�%��M�}�Щ�g�(�U�a�k!_ۏ��>=T�*=��n�/]�#k1�&Oh����5Vֹ
�� �)xG�ȶs�<T�ppU֘̓�2��v
�t�k�y�C͏S4T_�Cn~@u�l9	�3�t��hBc&�Jr���H��Ay4g�+8_���E��T蠱�2]�3�k����ͽ܌F��+�̜g+ʎM���QAlަ�p.�V�s�'7��G���!��9�`��<2Vh��8��;2�����%y�`C�۽x�n��0;a�H�tl���x`V�/_���:�������1��]��8�v�t��ۈ=0��c!Z���[��7/��V���Ǿ�l���W��LY%pp�t(�ahyǰ-��E���b��7�k�f,�"�h$�ؕ�@c�PL�^@ �T��C���	ݾ�= ���rE^:����?� �>}"fB.[��c#���Qg�.�C	3i��4GAuFxh0Z�߿�Q�o����P�4��{q�J �b�c��@�2-�(_"ʵ	,�?�h��u�ݧzD��$���-L	�ޝϗWk"��Q���
��O1`q�g�Q��K��$�v�M�K�C�K~~B^�zjh̩5܉W1�D7����%L�#����|Be!�reN�����_tJ�QRV�0ʜ����#��pؑ�U�-��An�XHCJu�����O(ҕ<{$��kn�	�v:Ŏ?W�u}�mt�3>���C(>Wh�i$M�:�I�������n�ڶ�����xo�>�.��	�2J��#��&yx_>aD��E>��\�#u�%�HP�N�f�wpO��A��S�iN�P���~F+c0�432��S)/@�]��3�$�<�ڇɩ��r
�G޷JOG�
�ϕ.e�d2�_�3\���*.'��~;�x<��4r�������4O��q}��)������tJ���<õ�*�a���c@gLv���� ��
`��<vP�A腘���k��P�K���EӍ�EZOëҍ%���I^G�V\��N��0\X!��Q���'\6�#�j�"M2�(6I�tk��"����Tx�aN2�f�3y>�*���"3DI+�3G��w������|1f/k�%�)��#�,&|C�2�I�0k{���eKN"hع�����Kr��Ъ�r�4�Ў�kz]�9q��K�&X�:��d�F�4Qf�W̐�
��	��2�M�0|@�9���zf����,ڳx-gpsuC�:�77�7��0��`hb&0�&�fu3���Ќ#F:�5<P��=����.��a��4y�����)�sEam�J���!Jw�7��LĨ���@x5���]����*)�i`�9%i:Y��D�^������~B����A�}�}���{u�U�dDSF�&Ǥc��:��4�8Y�fN�7��p{uMqohP�����G�l��%�����5[r�&�tb,�c�f�ڑ����o�۷/���[?	����ɕZ91��H4���p�6L<^�SH{D�����0EE }�w���J㔮>/���L&�,֙�����o(A��>��"�e܎0'�`̄Ԗf����d�y值[8Ai�Wܝ0�zE�����O�o�v/LN���+�r��<�.q�}w�ok��L�v�\�Qd���s��h��SʞN!�W�p�=c��"Ś��{�p��k�֖g&[(�;�zW˾f�Г)eJ�}�'{uE9d�`a21�����{欬5~�1.f�Ӿf�%�3hY8�LkN)�V�L��@յ-y�<��;�ȑќ�7��`4�\�E9	��̉`,#o#a���ȡF+�HB�32� ��!���5�ͩ�������� U;�uwx^D�:%���I����%�~�7z�؅�@�cZ:>�����R m�j�^����rO((ｎ��,z����4c���u�	�)*�0��#�B��*Wڞ�y��ڐ׮a���ג�e͈�Ǯ�^�^�^qopUC���YU��3q�7������H��T9���)g����vx�v侼�����C���~~Mo�,3����X�y=�<��B���}پ�R&��:%��d8��^z�%����� rM Ix,;��}3�Ǥυ���Jd���E��3�X�>�������.�\�1��ׁ�g�Z¼/�6�������dO�3��sќ�,�كP1�0	�d�oߨ���掼w��靲F�E��܍N%J1'�<5l����&�ι�|�����J��N�adh���a�1s�v��J�����+`�W�s���r��1#�b��t�XN �,}h��k��
���GNy�W��p�חg����ud�v1&F�$�M��-�WL���y-��Xʄ�a'�1SF��ܨа3�H�<�T��i��d4ӏ)�.���;����u��p{}g3v�B�$c8l��s&8;�M��D�Lx4����:��^vo���~���;_��c�ʩҰ--+a��ޢ����\JĄ+$�/U,
A>{n�(�L�k �I��+o�xTW��o�����#F�.�O�3?��D�=�iL�_Ƒ߃d�bK��x*�G�m�VF�>F�O��sy��4�cH��3�X�3#�~W��aP�&8v}�\r�X��N�绯prK�y�I:�{2��;i����
o�����B�0{�D�v��H'УU?p��'t������3:Y0�d�]�G��&�S;״��q�Ռ3"�$�⠌��p���_����W����t{8o�4g88*�d[q���R;��l��e���i�T�4���R�a�:.��>�A[Ks܉��d�A�$2�]9H12Z����z@��@k��sHm��U�]��P�:9-+�\3�g�?4�!����<Ct��Ю^�rZ��`��P
�I�w��1:#��o��g&�T�v�ifM-C�25�$�!Q����ߣ�����1ÑG��Д�~�ɭ�`:���4�#rJ妩�e�8S���Ͻ�5Q�K��/��I.T���z/�Q<���y�Xp�Ԑ5�NS��Uvg����(O�E~��r��Qyݳk�GVE�F���ˇ�v�/��1��2���u|��({5�A $��0yk��}YGAx�
�bO����'�+2���ZfIC������	|�~eE���`z���3����H'/W�L�K�w=������!���@Ɇ0b�o�	+Gk�����ق�*Z���u{*�@����1;bFm�B{Gݠ��Ѷ�`dF�Nͦ����x���.�a��6d�!�h����X���-a�a��v(��,y&S�e�F�D�(Z�2O��/�ޒ�����R�c�-��}qy��wdؙ�t�� K�'��_i�&&"�����?^�.h�6����n^���y�  1��dȠ�� �=�BW�O ��� ��D����0� !zڬ��рD����~GF�;6�$m-m<],�$"j��%v�(L�p0�Ӎ�D`&��oG�Q���ґ�q	�a�Ռ,{�,V���I���nO�W2����W��_���}�ǧN�8k-��2�N�|��F+�$H%���%�K�'NUg��0AA�������	�.� ��
����Hv��c�ۧjh̑��w y�Ԯ Y�Rc�����2�D�D�n��\VR�Zֈf��wn�Pu��E�'�����<��B���U���1���вJ�����sUg�2��2�_��_O�	/ ��N�����mO`(l�C�87��HȆ х	�P�d$Br.ib�����g���H�<^�.:X����r1��ޡ�b�Mш��Eœ;Q�p�(-�R�\��__���~��b`��������.[��?"�@�F�_�)����J�U������T1�0h2� �2z�"�E~��ӈq���zab�P�3o�(�� �a�b�;9qA���\��>�H
�V]�N�,%e���N3R�.y\��5,�U�czľ�F�Z񡲼���P,�L�)��	��;�vK���k�͠ߟ"\Txv�6�+/�t����^�K8B��xW��i}��J�bul�Ҿ�q��d��6�EYȡY=!&��;�GuqUڮk�IFU6��%��0 '�	���a��O�C��8ʠ���ySj8�ա�,?nŜnK7O�'1�#���UV�Bwr��>�h<� ��y��$k���y��gF���М8J��}ʟ��Q卐%���������*L�D��!�9��Iۦ�C[O��>����tJ�(;ҹ��?�ᣝ�/P�������#�Z����Ccr�EC����.>r�V��A��@`�g����w�v�7�@y{���_��Ï�~>����7�#F37�ۨ�_��0�,&A�JOKаsw}C^6h�A�!�n�ň�����ͼ#3cs :8E���;�/��������%�q���p�6^����6r�ַa�����3wp�n.�)�և�OpuyC�_0���i4�W�fi�R�뉕	�;aH��V���)���(�:b��d��ơ��$�d��p�1��B/B��!�5�Me�ݬi�9��Պ+�L�-��k'F*�l*V�(���q�������4u����A��w�/:�������p��=
��CGc�wd���~{�J�����:����� Xd T�"�z�М�r�
7����-݅�6y)����B�9k�T�������19������	�Ro�������@Q��96>*��g� 1��Q)!�P#� ���H�mτ�� 1_Y�{zf��C�fr@*?Ɖ_��p�Le����	L^����� ��x� !Tuj���'�PD�d�!���]��}O�blț�E�M@�=+�"����w��a� ��$��N� �N8�"�,�P��L���	�x"`�cF�/UҴ%& {��I ��	uG�/���_%�:�Q���x=n��W,��]�N�xu]�[ܵ�B�d�F�t�.��&�3>,ކj���ANo Ϲ�e4|O��䭃�<�pm��؃^g$
P;�ګ���h�-6� �aҼ����h(V|���?_��d,c����!�oW|g���Q��]�|������!d�**��}G�R�%�7l ���r�d��<�<ijK���T��C��O�8�����HY���R��i�Uz�����W���;{`��Z����M��2톐�ͤ�`�9]��";�99�;�x���2���v�5!k�JO�s���ۨ��ZT���y� N@t�vH�"}	���~��J;��[r\x��k�voL�	O����s���4�z8m�<����Z�A$�t(��f��E��{ύ+�x�������L��wk]%m�=��J�Ge�+5�.;�VOf9�6����ʘAx�QB���8�8��� 2Lש�!���m
m�z���9\]^���,{Yw:
�j%LS�ݨO���=����m���B�/��!8�ݎ^h���ٚ�T�	��C�l)�-�H=v�q=u���;��e�kfp�������+��֔2}���|-�2��o(����5E a[�C�&ӽ�~�%A�6��2r�&�����K���#�x�����e�B��O?����3-�d�Ac	Na�����$���mr�4l��سE_�y���(�s6��Lx$31� c(Bˈ���e�7m��:m6{C�Ɓ��em��n˾��Ճ�}!84�f������bʵ��+<����~�tO������c7�����F���:�m4�QN�:IG��W��?�̑&2�Ig�}s�����҃22_��G��*'���I����[�R��i�2bQ��N�,���UҲ9u��xe�T��?yՍG>ZU)e���?��*gXzRJ���Y��H'�
#ccM��K��X�U�;hsD���:D���u����t�g0C��.�==��Șj�a)�=v��7�u�$<�Bc�ħ��b�b��)����ʏ�*�"�Ԥ����GՌ�և-�):��V
�'�~�H�Rg����Ngn��W/�-ا�*o*����(}�R]�a�|DWMt8P1Z`���� �����;�sw��)lM� 'PZs�*�<�8�;���PCQ�yZ�>c�M'��{��m����4MU�CO�X�caR�EA�Cs��Z����4��).��M!�|�.ث#��	Ze�ud�E�yph&�PY�Et~�]�W<��[0��*��F����p�it4�萝z��d f�����j�Ҹͨ�L�~�NKKU���L�DR82�Mr��T)�tq�EFKkC#���V�� ��
/zb�H������,�ZǓ�ر�Ja�#�'�k�b<~1��2�I�l��A�[KϾw�G�#��R��ӟ���,���1�B����#r�	���v{[�f���i�k��L�.���n,��M�a�u,�h`�9��SyZw�CEB;��j  ��>�>=�А30�de�� �WZ�r���۞3�d�̨��.�u:�j�A�v-��z�v��8_��ɫ��z������f=�Ͽ�L��~��7�K����0���&�#E'�O���n�6͈��y ;�oa�*߬�����0��e�sXP�vثH��FΌ�eS�Q�2�-#N&�OcԊ,B�9��;2b���m/�o䡃;�BZ������+�����!'9Q"�	C�b#p"9͛�J,8���/lb���!��5]��)�	g�_~�A@L��]_]�u�@���@�6{���::��=��;�'�X�߲qg���sfC7���FY��3i��d����{�����n/n�~r�Y ��ח��_���|u�����/�d�9v�iq1���:��(ņM�gB���Uy�РrN����(k:do�|�F��MNt�P6-���q�2�&��箬:T�\Ѹ\�q�s
{2F/ L7=�ē�8�D�ʥ���+��?�n�L��&e��ӄ���.��%#�����)�U�&��v��$W�������C�1������=q��Ǟ���m��'�ӗ��M��� ƀH�$�Zg��_߶���3	�l�I4�*���y��bֻ�S�98���ɮ���q@�|\�����Nb���r�t�"��G��/w��[b�C��^\UXt���Y��^2�rx�PN�e�E0��;@t!����J����	\QN�r�N������^�"�~]$3�^����u�Mӊ��BD?Dȉ��OG?T�~�x�u���l��2I^P�'N�p�q?yT��%�%;�$~�q�5J�N6t��vPWU0a���TqIk��e� zE�K��8_�ce|�tc�hp�5�h��h���\��2����:kD�����z�d%:�KǤ^���՝|ɺ��5Z��P&��d��9�߾��i�ѩb�g:�<$�gUg̉x蕴�1�4�ߡ|����xsi���Fi��xӃ�>vK<��1m�EAW��Ƕ_�xʹ�^n��d�d"���g\�=��A��{:יq��������:R�9#�7�ɫq4^���x� ��K����$��V�b����Q����yHz����z�|��nR���bQ�tDul6|	��ҟ��\_��F�D��S�M<��p�^V@��߾m�l6�tqE��g�=�<'���P.����7��G��8��^>��Ѹ�w@O�vߗ���Ŋ=�M�O�β���G��w��u��k�4${Mi+ٽ[J0�ɚ^������<uЮ������./.	0���G��A�Nla���C��o�������V�Ī�'�hYG���%y�|��?�}�_>}����ֿ���UCߘKr���?���ta��\ȋ���t(���Y�w���.v��>�J��Gvπ�QD�Aa�lr��CĶ�s�DO�7��Wg���0䬟���y��o^��������O���kG�<���ېUc���_�ⲅz��X�ٱx�,�!�<w8���f���N��ރ��z�J��]�;��S���M�r����V�L	w�ϮXt�)^�PXI8*pզZ[���cƇb��h���W�Y�#W�.@�� ���PI���]ғ>/��ɶ~78��oW���$3��|c(���^%��/�z:���!���?�#c�t��I�B\�x�����l������V<yA��E���(�jM'L<��z0���O1�h�[����jr#��5��]�![jP�vgυ�Aۿ��rWO��i�~O:G��<b�YQ�W�ޚ|�u�*t8-���f3,'jj<Q�]&�3�Cxb����]��o"�2 *i��F�,΀x���x����]���w�B���T� ���L�1f8;8(��Sl���0M���*�/5d��9�Q8�Zټ���wnw���K�e]�t�� �y9�vYu�I��ʃ|߆őy�-�F� ��|W��q�#p�iS�'�*���/
"�Ԍ*Y0�D���O��smH��m�����ɕ���I��"�W�Z�C`LR��9�?���mv��������eؗ��/�H2e���[�0����Na6c{��A�3����0���:�t���5��� i,*�h���C���ԕ�$팓s����~�e��~=}�^@o�����}ftG�l��<�ϓ/'��"˛���*c�!6�0S���؆4��G��T6p5�5̼�Ш��'�
Q9�~�Kc���L�-��մ�ی��(�>�2���3,ю�s�K�׿�3|��@�
'�����6��A<�V�/���9;�#����W�ܲ��~6�ȡ(: c�~�
��CsHڏ�'b��(�Fq9hS�P�f������a?�|������...�_�>~�3�1�A3|cdy,G�Qh >b��EP0+�;�{��W%�l1��%|��F��5�ǡ{�C��p~ɖ�L=~��(tin�Тa�(���Ia�W/ �bYm�ݐ�s��'j����A�dQE:$����,V1�?4^�^��[�y����O_��>�L�Ȝ�<�����#v�Y��N�����BoL~OM'��7&A	D�����|��1{���1X9y�~5:��XHc����ƃV)z��z�]�l�{9�2���*dPK�,�a�P;WM��H���8���4j�Z���7��b�w���z�)�"����K�����T	~]i�v#�5� �P���遾{��L��7hPyE�Et���ټ�E̮')A;�0����|V=�\��~�K�:u���;bl���Y{�X���fʦ�O\��C�^:;��S�n����i�u��/G�X,yQ��`ɏ_�����y���/��s�SY"�� Q-;&z4\vb�i%f��69����`�[��B�ܻ�2o�nQ@�������i�5�ףQ�!��Ap~��1x��֯���6ݎ�x(^��L��GBs���3��]u~�`c��~�,����Ke�%(�Tr�X!7����҄�����V��O>zD�\���<z��5��fn���8��]�W��m��֌�-��|{P�Ё:-P�TVZ��Z�w�7�_R�t�6h��X�Jt�;Qj��8-����&�W,L4�в���� ��k�7X���������0=��uz���GƲ3ښׁ'�F��`�L�g���+����l��莬�Q�i�گ����W��$�3��8��n��+�g������(?HY�t=��U�R���o-�&Y"�a��\l���LX�+W��[ꌵ����t_�beiJ�������)6�� �k�`2���	�t��|��v�!c���0#\��DG=p��Z��A��5Y����k��z�<z�}D�=���!�����y7 �d�E�3��Gv�!��q1	N��"x|z���G����<���a&-�Ϲ�����[���|��\\^��`Fc9W���hV]H�Wm˧rt�4����^�-�C{o>���-�ׯ��m��/�k��v���psG��R�#�2�4G,"��5���mc+��`jB�x4�Y#�a��;�T���E������l��'�}�o�|}�����7���gx޾�l�$WjdBi2N��V�7��h:��p#�]��G}(Ĩ{_�Dއ8�2Ӄ�_"4V|NG��4vJ_�[�~7˚��wxS@l�� YH��d���I�J������e�>�	�J�9��e��5*Aϥ�!V�
c0q�2y2�ìz���k޸�
Rkk����R덵q����a���P��'u�>S��F�U�PF�����{����i�)�IY��q�c���l	������_m�*"���rم��%w����	���)i���r'�V1��w�cQ�z�ģ��Ϲ����O�&�����c�%�o�N}�̉��9f�Y�,8��yO+!��;���L��� ѕ�_wċ5VjT����hء�C��B�[��u��!�\&Ɗ�(�/�<�}�M��_��+��J���\~'}�(0�S�ɚ�G �W���^(�3x��,��B�/W�>�b��%�9~ő�#���qx��nwQ*؅~���WX]r�������b:^h��Cn�:m�R��z�i&pkg�Z�ɟUM�g��V3�����4{ض;P��n�0_bV�2],(���=��ϞG�ml?pf�������]��YGjR�Ӱ���z�����X���@���!�W��F3�&�8鶌ɂ�X!�yO���@+�%�v��O��q2�;U(�"�����3y�d���F�����ш���^�����Ts3�V9�h���b�͓����6�sF��ϓ��%�����&Ѱg3nh��t��i|������2I���Һ����ݞij#���!�	�����/�5���_���.�gpyvN�D7�W��Xd�L=�D�E�\;l�I� � �ngdLL�r���Y�~}���M!��$�j1��lտ/���	�И��L�:���I���?������?}�|������k1���C20t��=F��cG�\��/iɜӉj�JD��?���_�<��xz}�|�O/O�򲆟~��o�~pv}G.�bu�o�` D.El2�ѨS/^�ddӓ�i���&E1Ҝ��9����ܠ��������^�ׯO_��o�_�_�{Dj}��s�:rW'��]ϸ!�a5�6�@qΨ�,>O�D���;��}K��;ɐ!����ĥ���Xg�z9%����}�1�� -�m*��.� it���SRӔM>IkO��`��)���=�(�u���W��UBS'�e�.�P�cY~�0��b>ú�`�����//��/�]��_�V+��|\��
najy,(U��Z�f�q�f�T��S2�e�ة����B2� ����߷f/��=�x<�I֐��Yi�Pfodt��]��#���s�!�)�!�S�jW�,��sd����-��	,��v��-��D�+�Ct�0k2�L�x>��)EA����"��s�I׸SK��V "1	d���`.�S7�Lƞ��]<��E �}�E셛^�:4��PfН�GH�.��4f�Rڡ�'&/.�$��(F-�{e܂Sh�6��dQd��7��]���-�L����Z����Od�m���>q�e�����/by{�԰L�x��Q`�ƌf����7�M1��E�B�f����f�݊!rt�U�4�-:M�ˀO����
*�'�8u��,��T���AF�4@��Lđ8l������~�WSћ<)Q/קWF.h����B�PY,����+�yZ�.�)0�����^9$�=�.d����d��!mM/�'B��qY&ϺT����#�!6�|��yn\��6>��-�)�`��h��3^3g����X�ڨ�tB�=��wt��o#��������F �)�}z�=!3d�2c�ˆ��ߑ�[>	�tAe��gMYː1Cr٨:oUK�t�ġ,?���*ш�X}���}�ǧg�:� �ü�ж��_���ﶽ�@��\�+�x+��QC����0�a�D�L�%�`� � �72��?<�����h �ou��˾�?|�H�Ow���V�5+|DҲ�7���T�&�g�I���̨�k�6� Z���B����s�|�~��~������L=���O����	>�����-,g�h�J6,��@#���ɂt�ě.��
#j?נB�\Z�uo\R��@
f��ĕ�N1�
]@{��~�AxE��|~�����f��Æ��:���1��.Y7�`�N���<٣ɉ�#���V��}3Pz�X��c�5*}���:w[H�[M�	�� ,���^�u�
Z�p`��$�"�Vm��� �g�;�7xyq0_�tbL@ԂU@��V����m�-�袚�VZo�b�d�������:�DB�r����Mh\��	�4���R�aez_�$a�����D�TX��GWdm��թ��$Շl:�q�Lz<�rC{�?:�k!�X+mm�=��HC��M3'/��8���Q\	��
Ǝ�Fq��C��:J[#i������0Q�����2`x��������t��ý����iԕ!�ɫ6�y�ޗMi<�_7-����O�(�]dªt& p��צ�	,����J��|�M>���)�:`L�x렧�� ����v�A��4�9�n�;��h긙m��
������"��cӑ�ң��2*���*��|��y���'��������C�v�D�d�|�Pp��R��XT&>M{멼��45�m�g�c}�!��*�Lh���e'�H�"�B��Ym��2[*��B
Gږ�]�ѡ"��n���0��j��A<�Kk���5[N�ު�0�z�~ξ#d4样=e�����e�?�Ln)�G�V�O��h�C�),e�	���|�$ޙ2�2v����<~��<~�\?��O�������aٌ���W �1�d�En��H���N�ܐ�+톱+�)��V}^ �-��y����.3Z����Zg�઒�k��k(�c�]2�u��l�G��m�VjI0⦦u�!��8���X)?8F=|��U���'� ��7���U����u�7m���z���B�0Bh���S�����/Ϗd�\�ȉ�ru!��3�
;���N���<uf�^d���jS��]��;�Q�=�z�C�F��՘���D�Lk��S�#����|��	���ʹB �咼�� c���e��8\H/x�g:� ��w|H���i��D0$�*tZ��dܹ<������_~�חWX����@���78;[2�4�!/�}g���|�ￛ��g�ᥰ�MV '�������5�Sd��}Gn�A��צ_�7��顟��v��O��3<o^z!�@�20嫥-�`H
�Y$���4#)�e��F�i�����x�?c�C�<g2M�=����U�<�BhA�E��S�thUX�Ȍ$e�}����>E�]�m��As��~;�re:_����d�FE֭�f��ګw=v�p]��N����iJ���>�[��jF+ �Ó����k�r#��`I��ݾL6s�+��lɌ=��&U1"�XdI�ݜ�3mIu��P��G��^pPfRƳ�p{b i�K�ڮ_�^��U#��-�Z��lݸ%k2 ��z��\h����~Y���L_���8�?ȑ)i���e`�E�wm��q1!JЂ#bN�
`-Zb����q�x�k����k�T�V�7�.y���\k���z!��3P�>��zU,�Γ=�(v������`i>��y�x��`]G�*����E�sjG"����)x���kIٝ��q!;V.�<����s�fe��v������) َ=Dq�t��>��5��梔��>9l�rG��b�L�`��	�"~�*]�Ko-Ȧ</8�R��o|8|��r��N4Xӄ�~|�)o���Q��=~�����MƉ�V����4xf]�m���˸��Z�c�(�z�ZL1����?˗��r���=9� �)�*`�˖�3��l���N�Gِ(;�����Q�Nk/t��`��˫GF������xl��Vi��:N$'���UQ����9�v>�<��)��5�nX:RAq�;��*�0?�3O��Muϡ�^j�pY�P�ga�%��ܓ(�<rJj�C�~�5\��@H��e���L./ %����H[�ӽ�����3�Q�J�t������/�bN�a`�,(��`�0{�73�C>�a�P'�n�]P^��e�e�Ŭ����wzhz|d����̆$%|�?>�����ӧ����@��ޱ�#V^j�$�2ˈ8!���9Hܶ��-�
M�;�/�s�uɱ����?�����V�%��͇z��==<|������/_�/_N��Ȯ`��b̏%�/�`5g)"h�0*V�:�a�b�J�t���Ï}��������Ԑ��h�^�^y�J��~�o|c��(s�94zq���ݻS�&a��\����T��M�f�,�!K�	�U�S:�8:������'�뉡�L�����刺����#k��9�EE(!�)����i��,��?3dCd7c�vyR\���� ��� b���M��U�k������E鍞�.�4�	Ɏ)ieVy�3i���4t�+e���* �/U�C�������J?�v�(�>��4p�|{��x�(G����%m�M��8�#s��<q����x&����q�p7"��3���%a�����0z��T{��Z�cn�5'��R���	� ����G vBX�.;.s�c2�o��DS���st��g>'�H�@��({��i�W�r~�Ĉʅ���vR]9��F�I^ ]m�ޒV��������5"���q�vf�.\��XۛiZ���;C�mc�W�t[�
�J��>�LIP����F]o8��ד�.��b��7���e�]��0nMð�9%��H����";iu�F���f���+/E��i�����f��Iw��;������S��呲9:C�r����) _`W���E���/�g=.�lZ�5̅|�,���M�m�����<#c���9�l�@(��^�7W�K
d�`��Rx����j�w'�����"b��}�O��r�&�d>]��y�P��zt I��m���V�{�c�J��dr��ߐ��SD鳱Hf��0�	l���6���yڊ�J�6���quMM�����z�J��R�dU-���U�'��γ��1q�g�.�5&�I���w�up���[ȉ�#f7�w�sփ��n�5���v){���|,��9�l����}L�u�F��
'̩��Uk%������	�
߅�3�7[�
���jhсC�WE9)E���^�Wzyz���z���~���Ϗ����3}��@>�]��s�n>_,vf�X���'`9�2Ø�(sf�����_/��B�_�_������O�����,������ӧO���g���o����HnJ�H�1�Q���^x�z۟{ �6� ������l�T�vw��SK=oo�8�a���'z|�E�~�<}>���+_��w�t���3�-+�����>ҡ8 R�It	�J� &>�V>ٜ~�"��g����T6[�^�8Dzy������'=��8M�92�B�ge���^4~��g��Ezdm���h�7�x��0�]�����!���,p |iZ��I�O~���Ѵ��X���R��{y�n �*����¹���_5�����(���w: �����w#�@��B� �Ł��4�%�U���5#�M����'�~6��gO��E�]��5 $����X	A`�~u������&�0��#��p�
I@�մxQ恝����{Q����� ���L����j$ }7�'�M�0�Nu����W�)U��7���7��!�j����Vc=�o�1�;���3\��y�>���h�ɓ;zQ����c�b�Z�ɩ�����0hհ�7���1P�Z����_���xS���Ô(Z�:�5A�j��mOy��)�N�^��6R��cWk~�Op�$z�`N��f�U��{�{������H�}��l-�7r��Z����'9Ŏ���:�Q����U��?�s��1�vU�@�$ÆM2�"6C��M�����4�NX�A8˲����on�~��V��#�V��/ �h�+Ϯ�b���\4�M���cg1,aV ����Ν�*�֛�xm�?Y���ٚ��kEG;����KJs|��*�|ݬ��W-��X}��+�3gi��Ͷ~���/+��[��(>�{����������lj��jH0xU�����`
X��&8�E���|vP������Yy��6_N�뒊0R.�Ǧ��cR+!�*&<��$��/D�':t��N���z�����lxRN�+��;�Vܺ���"��w8�����m+���_�o��p`����[�����O�sJt���r������նT���mɬ�F	�]�6; �h�� DCᚆY�Aԍ��{�#��{������{}��������7��)��]{}~���*�7{zw{G�둎�/b	���$���F�N�$��T5�L�pШ,�A=����A����B�H>�t��7EѲk�4�����:����k�5f���t�g���mA$��0��Q�5�##0��Q D��M�s(x��+�g�����i�pϓ��?�Np�D�#����A���������Vv׮/7�{�����'��Ԁ��wuW�Κ��+��3ܪ<3I�W3�料��T����Z��	���òS�
�ږ>������:8��p\\h ��8l��5��
� W��݃�Gj�n�0h��#aRG1UWp�?��ı8b[���%ˢ�Ŏ�9��ـ���I��ӷӏO�����/�=^���_T��;^H�fh:s���}����O���s
�y�,�[=^67�N�ea�N���%��<�z xu��
�����g��w�o�.��D ҲgES�~��9���{��{���|jǾ|r���Vc���+v�8�@fH�F���mJ���"�Z���FqQW���'��Ψ��F��c|=Wew^����f�|��N����X�l�8ϥ��S������b�x��>�=	V�1�xi�Z����6<�j�=��Fj��β�R��mU����ְ���
X���JZr��M�|_Ax��:m]�5���c���mxA�OWV�9�(ۧ��#��F�����,� ����MW-�M��9L'�ٮ�A	���iŚu�JNaЌ�C1֟>�'��ȸ��Z�d��d|���y.�=��-b��AkÜͺ��x|�t�V1�ث��׭�(ǌ��wU���9�Ʀ�W�1�WA�h)�,p�Z�$k[�^\�����K-_^>��١펉}O��YH~��_7gW1%�x�1ܞdV�?4K���2�Pȏ�(�S�qVe�����,Τ�����;}���>|���1rQ*�!�n�&�t��ꔺkC�����Ȧbgɺ�FJ�T�P�Fdf6�H�݉V~�0ч{	?�p��C����vX\@&�?���U:����S�߲��>M���"E�[Ʉ�<��RA�����?��/bͳY�S��X�S�Y�]���= �[N6���(v���n���&����` ���]҅|�Tvے��c��AYƋ�Sw_v�xk�ڑ~�����B��9���b�V^�M����^���gt�sNW�F~Q��SXx��2�~��y��t�%8^&89w`"T3ٜ	�F%7���K�q��b���]���7<f�;�S�/g65w�k;5���4 [��e!�@���W���|R�d��j�#&�B�'�O���*� ����S�s@7'e���,fJڲZ�$���d�K�1��|��k�8��5�����[���1��{�g�[�=A����D��B-[�[�hK�J'�W%��o�0)�w��j��aBr��S��Ks�t`;����*�?#�/�SڗC�7UqiQ\�w,�����+}h��
 ������箾v�J?���6�yb
��s�i����j��ײ/1(;z}�Cx3����ܾX�!qK/���sm)m��q�P�d�rС���Y����ѭ��r������Fl��$(�����C�Bi� �>�m^~�_7�:]�ɫ�In\�<ڹ��\��T�H����5��Q�N���UN����i�6�k��ר���y�1�_�Ƥ����r�X�Ʒs�o�}.�U,��r'g]cK[�!��
>yI���U�#>��ʭw��b@��E�+�:�J,o/~3:�^ md��e���[T\$X�l�0�͵�%ˉ��U���r�*W���b�S�:P�|��b�ꉟ"�N{v�R,f��[O�9<ws��g'G蒮ÊA��>��j}]�:�V��ooo��L)����e�'���-oqD��~V�S4�<@j���aQԟ:x�˝��f� ���_=H�ʞ���q�Y�JU�h��?y@�A(��h.�v�&�$*����O� N����_9�h�v����8`4�q\��T�/c���@ֆ�1���z�R��s� �����֋)�(��r�+�8��PR�N��d�7RH��":A�R�kSO�b}⅃^��k��҂��jS��r=��e�ãm�！�5��e�~���C]�s���}.y�Ŏ�׵|n}����9��-?_�Z�0�����?��͍S��ZN�`7%"i%W��A��y��\s�Q_��mU`GD[-n�0Ƿ+v��NS�K���*�<n���߻4��mM�@���r���"c�?or��,�L��'�N���d@3u�W[��o^���'���#�y��"��Ds�lt�8��Y.c�{����P���Z���B�[-,KU�B�%Y���(ة�?7ϭ�D���kL���3m���q@Gռ�kx�)�.������=V�ᙬ5	�e���Ə_s�M^��;������@�b��
6�0��cRW(C���9V}r��Ӟ7�r�-�Y�c����[��+e��P��j��c����=�u��\�)&�vn~{�)jM)����u���ZGg�i�v�)vګx�M�0��ֹ1�z�N�o�k:[�v�s��uqo����m�x�\�����bD���v�.�T2>�m]m�e�ZX���4sG���jץ�=�=�٧���,mw�2���%5f�A����fE�f i�^�ޙ^��(ʖ� +ǩ`!�S�Dm�j�����;Օc�	�u�"�z���^��7,�̪��ԇV��#Ӄ���KA�cyY�� ���T'
�̦�r�+�	a��Q��nG��N��I+踊8�*LA@�w�T�5t�d@3ՎTj���L�ͭ��N�r�8Y>f5U��I�|I%0�8M+(�N��؉�M����e-�EQi\\����ܷ6M�ֹ�mB��:#�j�+�p`�@��y+�.�i�Րt�s.)�F50���q���L��G
�|}��@��~�幙u3�~΃_X�Zt�n�c����З����vK4dr��=��~��Z�<����lւ ��?�Q���= ����P��V�� v�8�J�lP우�;�9���wW���Wim�8�5��+z������~ڵ��L�`�ř֫#����&դ�A��#A~7<�բ��7{��0�̮-P�xQ����D��Ư�$Y�������2^��2)�(�h#�v����; �R'�@�v���j>�f�iW�N^i#��KsaS���5m^�]���5�	��mOԱ�q8R��=��������������O�������#�	'�+Cp�Q2�JF{���~�CQdQn�����o:��X0W��๘�V����(����Us�kƩ!�!��s�f>P�.]Q��:ަ�J� �� ��8�V�״"�����Jԫ҆bg;�.�qE+����c�O�[R����T���K�"'����k����ޞ�{+x�Ŧ�.Ϻfd���Q!�������(#.�srS�=�z��G���E��Z-���	,����Xذ1�>*v� �T-�%��\c�(�G�~�l��Eٳ�[(���,�`.B�C�<��zw�=0��cmWq�\�Z^)�L.�*��czJ�b�J�J[:�Cc�,��68�2�@����$[u��D�J`�Y��ʹ���#�������id(w%Xb����׌��{�Y8�w7������[詹=j� �'����4e]� 0L9�K	;�VM�?'6vJr����h7� 겑W[�%=��#��`r���I~�꠴�V2�&Hh�Y�1w�e���̯����&�,z��H("D�b�q�z�21�A�S��k�D��x5�&_��Ll�#m���4��Rn@�FbJ�L�������;|Ø����zq?*���H��F��'j䥐W�w]��m����Z �u��@m�8�!j���
y�5���������.焖\��/��_��N��Ζ�?��ҙղ(��^�⣭�n6cyQ$Z/�~����?�[�_L��vDT� .�w���r5�tv�h��{���߰l�QuX��j��j�qD���Y�jԢVѥW�;ܖ�N���frY�_���:��o`����G
�r11�(uɛ�~��yt�ji� n�kC���+ny��Έ�I+����e����G��ו�/�8.��I���F�A��Ϟ�Z�n�у=��ղ��z��d�KS�s 
QV�\v�ΩJ����V\V�w{+�Z4�����I���eߛ�۪�"�������E5�̀-�N��g��{�M���N�>�(H�R��}z=�������2��Z    IEND�B`�PK
     mdZֆ����  ��  /   images/49e5ee10-9185-4279-8a25-10889e7bb4ef.png�PNG

   IHDR   d   h    U/  0�iCCPICC Profile  x��||eE���6�ѫt���H�w� �l6,�d7$٥X��lv7��l��.  ]�4\�R��4������I���̝�x����/�}�Mδ3�|Ϲ�^��3��¹��I2o����I�{�wu�W���o��$��,Z���Ց�'�~��ǒz}���J��~֛9�h I�W,��K����/$�~♱���%z�ѳ=zeǓӛ:���V�)�V[:0}��$���^�(IV�O����y����\�w�@w漙3�d5H$�=wɼ!��И���>'I���xv���=�:c�\�GЭ�m���������:���L�^e)cͩlf���:��������C�6MT2M��4�9�5�kʴ\����Ӕкdx��v��{Y��"��t%,I��ݓ*��,iƫĿgZM:��d"^�If'��|�'C�@�m҄v��5azHf&�k�%5�R��BP���q-`�%g)F��I���ןŃ,����͞���M����5��$$�͹�^����OĶ��r?��μ0Iڶ ㎱�|�$W<�$�\���$Yc�$��m �ۜ¯�:����������\�\�ܖ<�<���|аj��a��7��pm�C��ZcT6j�CF]6�ѕ�;��o���ό�pL���<1v��3�^1����#�=���+�_�+o��Ze�*�Y�
��Xyՙ��q����Z�e�[��k\��Vk���Zk}o�O����9x�q랾�V�ݼ~���lp�6��U�m����xݍ��d�M�lz�f37�p��8����䋷5���-W������j`��~m�k����[}���.n�ӼSm��{_�Kzov��� �s�t=�t�)�w}u���qh��w>�kg�\6���G'�c��'m�k[��׏�풎�:ߚ�QW��K�/�y~����q͞+�������'��3��;�2�Yl��sާq�ṿ�����>=�ˢk��_z�.;�u>�kr�ak~�u��[s���vܣ'�{⸓.<����O?��g���Y�t�%�w^��Oλ���-��+/?���?k�z�k>���q�~9��]o�����x�7O�y�]��s�}'>pȃxd�/|��O6=}�3>���_���ޯL��n���Ƅ�v~[����}������bE�W��h��(�v%&6�6\7j�Q��zc�L���1��=p�z�n\i��Օ_^���9���a���1k��օk_����>�ޟ�m��7\k���ɞ�.�������՗�/}a˦�-[M�z�6˶=��gmwY����������A�,�R��M��q�m�������Խ���-l9|©�M����]��Ү�|}�n�v���'ϛr\�����J��S����s�<j����o<��W���o�����0c�@�̹��f�?�;s���>�{����=4��o.�dx�E�,nZ���������e�<�3��;7}��C�=���W=�z�8j���<z�1K�=��?8�ǟ��\u�'���kO����O������'g�{�g�z�~t�9G�{�y���K~��'��w�~/���.���	�ms��W4\����_���G_]�f�k7�n�_��[n�q���9t�_|�Q��x�ٷ_|�տ��o����w>����z��w���������?���{���{��?��������;��>q��{r�S3�����gv�v����ϯ�¸G�4��[��_]���4����S�xs�['���|�w?��&�o�����}t��ϭ������{4�0j�QG�zg����������m6�����\��%������Ʃk���k߼�=�>�ދ�������6�����	�_���'��֗�m�����v�z�6ӷ]��C�;����?���{�ǳ�ث�m�oՠW2��5���[��r���'��-&�z���]��o'=������V��b�W'�NY�u��u�����1���1q��{��i߸��֟����������fN�54{ɜ#�N���}��{���濾0�o��-��mK�X:g�8nٹ^u�m?�������숶#�8j���?��cN9���_zܵ��r��?x�ħOz���Oy��WO{���~�����Y����><�s?8���?�����B�8�������o����.;���8��î:�g�����Ϻ��k���_�q�}7<r�7=�˗n�ǯ޾��n�ܱ�7��ֿ����w�w����{f�;���������?x�C�<|��}�GO�㩏����O����?y�SK�����g��e�gwz.�k���0���_��KϾ����~�W�����q�k�__��%o^��5�����y���`�������㙟��H~���0�ἆ�GMu�h5��1�c~2��co����W:o�i�l�ʫ�߭z�j�~�g�y�Z��}�:��{�zO���V@����Mnz�f7m�Lu��n��K��<|��[ݸ�Cۼ���ۭ״]��_�'=8;���/W�[�=�Q������0f�uw���ZG��	��:�_��Io��������=:�M�є[����3�w�ԁiG�qў��빽W|s�o�oO�=���3f\1p��������9�ɾ���l^���t-��o�����x��_.��?����A���w�w�~HߡK;��K����Ǐz��c�;v���Z��<a��8�%'t���~�CO?�G�q��ǜu�����sN<����8��~��~rÅ�_t������t�#�����]~��_y�U���ȟs��לr������]�7�x�Mw������'ny���o{��7�x���fŝ�7��ݫݳڽ��7���~�������;������Ǯ~��'.��EO���iO�磟9�/�?{�s�����x�{/���/���K_���;���?����o����o���޷�y��wO{o��n|������~壷>��'� rX4��< �8>I&�+�jŊ��N��]e��X���I�J����b�s�_�dʗ�D�^��$��t`��r\�su����cV�M������M/�v�*�N��d�?��ν+�ܷ<IF`��'�utT=`M�?���iI2p�{�94��V��@���uK�j�^	ϯ���������v`�dc����ߍW��U!pS�0�0{��_�+p|zT/^'��L��g�Ex���F�6����?ݿ_�ߟ��S����|=���+����;���^���h;s�{�
L�K҇���������%������2p�8d��-u�~8$�������}�[�@�K��I�ecv��2�E	iN�g��Z�� �A�[W��c	h��b�O�9�f��)�ՖLN�1f+���b�s��oD6Bm�	�|��Ԃ|��Ѓ����?N�iG2�nP�n�^��	Υ~�C�S�h��|�Mh��\�cMK��}��Y������'�aӈ6}�J��d�>�����\�$Нh�>I	�L����$å�Ɉ�U�?�2��ԇ�M%�'�&�4��O}H"Ȝ�O��$��?�ҥNzK�9��V�0�tY$�@%��C_�ϛ�~�9 �6C��h��c���o��Ѓm�ܩ�/�/}�1���|�w��Ŝ��;{�y�Z�T&���v�w�N�6��^6wn���Ќ���C�W{��g.���^\�?k�����2��}R�䖑]g-Z8<�?��������6���ӿ��ٿ��L5��K��d�:Ј�������v���T'��tu���X�i�<���ob{g_Oo[�$1ܔή�I�m{m�sjGo{cǔ�jc��	}�Í�ޖ�Im�}�{z��v�M�6���=�x�:�U'b�s��u/h��.��`�s��}�B3V����w��6��Kw[Ϯ���S>�	-=m}��o�X����jk��n�ȻuL��&c�X\_��NVm����̘�jmMp�XZ�R[˔��4V&O��l�h߻mb_���4�6����X��>�mJ_��޾V0L�n�m�2��kJOO���6�T�І�����胈����Bo{*�K���ͩ6��T�[��ՁP��U[q��gV�Z<'H�Ty��l�W��Ϭ�'���Se����͝8�����6yb�ܕ)zں��A2˳>�THqBGK�n�B;�G��6����o����l��Z�Xٵ��7��x��}_�Wml���tN�һ������]�z�v�چc�6N��m�{_8a��5e2��}��V&O���݇�����1�����'�����B��[�i���pJA�������u5ɾ=ݿ{��vB�{�=m�=�L�sT2�v����Z&4�#�dk�Sa%�Z�״jT-���U5�Së�ո0�����|��OV���g�"X�E�1+MZQUvSߏՌPR`M5��Q�)SVWtU���/c5�,SUY��pK�	&S!*&J��%3�GGX8��S��ظ��~R�D&9��(-m�*��J��t,�,u�gBXj��GF+�⺒�И�?v4�yVe�k�a�c��d#T��Q�Qe5w��"�i�0��2��T^�b���Yn���2)-��M���(;��1���"���L1[5�$�}d��������יѴ���(Q�T�1�����*V(3E��A�d��8F�4V�Ɍ�c��:�d��wj܎>K@����u^� �h���F,˔��g	�	�&B2�II)�
���DZF����f������D�љ�)��ĖZwdҰ����X��L�-�z6)T�Å[�)�Q��pH���� �ɌT�&d��Y-���:S#�z��!�&�f��c��3���VO` �rͱZ�o�Z�yjmN!�0jR�z�՘4�\b��6�*�ak�����$U�,�*+p��aF�jR��	N��\#�q� �V*���he���5�2)�r#`��=PY����	I�]O��X�m	��b�ؗ�}a	Ο�贄PX2�P9U#�ġk�R�
[�X6�hN;�#�feʉ�ڹcq�O>�s��#��I����N>'��N*h��,�B=��$�!�Ԓ|)�Nji��n�c&ͬ'���(�p�b�Y��*�5o�uDF��Wd��֑��d4#����� mWp�ďȝ
Rc��0h������ؘ�QW3�0PZ���P�
���{������V0v�c���P�GW�4��)X6l�,��.�9X��
�!�
�9�[G����9~��;l�(HѺ�f�S-S�e�)!x p�
6.!j�T����(��?����g�(�����"��U���6U�TBR�
�#�g�k�C�GX�)q�>@9�(^{^G�PEi���p��A3�6��[=� �i�������a��hH��K"�:�+���疤
5�)Ed@%@�f�0�Ԃ��@�pĄ�2�+8#�j�FZF`|!Nj{���6�8Z���7VuA��BpO%N�W�)��J���F��* M(��JI��p\���mf��RZ�@�H�X�V+1�_G��Y/!��R2L�,ڈ
,E���u�$G��¬�z8;�pxX�2�����$M#,�(nY�$����q1����% �T��qdX���i�F(%�:��f@V
SK:@& {��ZJG�CiZB?&9��ٚD�68����#��B���Bt *��U-
K�YOh�m�f�U'U�ۑ�`�F�wrHaL�>��@dX*2-�aF
VO�&a���dH�Ҍt�֎��0Π��a�a�{p+`W�ϑX=��4�גpp��wX�EE���!&: u�"$\�%,��(]�5D�����ı S�c� ��)����W2�>��E$geK2��[��4�I��L�ɠD�ӒL��H~�4�L
���<p0L�_�+Dֈdڥ~��5���e{���*e����8t�đ�U4���u�b2M^�B9%��W-�=:��Q��:H�'���j*��b�����H�#+ ��'C2���U}GA����#�t�^
�uI���(B�(��(��g��z�-�'�X*2�|]8aC���
$\챾#�#<�Qsʩ0�Ó|3b��%eq UC�AHڎ�,EŔ�q�9��!�������{8VSVȉ'�����J���LX*/Q�(.8C�����<�BF�E�!GqQ���cF�f$�.Z芑%E��! ]�<���QM��|ᨒ�#� �t��
�����[�*d�xc=�g >H�E���H�tMZ,Ք�1�����Fy�&B�V1��Y��%�֨\J���nIu'�i=��u D�����Uj5:f%�@�`�P=red.��paι���� eU�:p���:��d��/�� `d��i�@x6+�XZA��?F$Y\80��2b��T���9e��UB�����P=^���c\*��8xPޒY!]� �V��Ǒ
��"�{��b��2:S��& �!�:�hH�(�� V�-q�EGAZ�H�sN
7I�V�Ҳ�S4��"'g�z
"�U�Ҭ�g\,"��J���L��|�
I�GV�Z?�MK�F�\�5�r���K|kT�T��|�����@��%�5�pF�.��\��\GU����\�l8;CU$��'\zH�=���EO���\Ru&���qFs�U���%�=����� ST=�j�EONY���*ydEU ��1Z�-�:~��6p�)%��r�YL�d���b��e������9a�Գ��{6v������M���'+�& 08���34�=y��D	Q��a�������K(=E��B\Flir���irƥ�lG֔�{"IǏ�'�Hwa��o�T%�&@oq��q��ʼ8_M��%3�ۃ�b��V�9��&S�l*+�AظO��lJ�3��L=��9mI��R�|"	@LU"CY)���be
0@CN�ƔH��
��²��b�p����"�p�1V�5�e*` -�s��6N�SF5錕=��� ߗRM2/��:`=\`��g$�p<B9-U�Ud�J��%^3�SQ��rߔjT��D�r�J�f�d�v-�Ne�ڒ1]�5�JPq�lؐl54����֔@ˢ'U2*i#OE?
��dX����k�U02.:OH�Q�N%�IoyiS�l��xIFu[x�n�>H\�����)*�k*�"�PO%��J�Iт�)�r5Fኍ�)�`ٜ�)z!*N�*�@aX)=yL鑘(�&QBS�Pw���fS������ğ��fya3��ss"��<y�����%'8Nk�uC@���� Jz�����?���\����l6��T�'�/����^II��i��lѓ�}�]	XC@N���e./����?9˔�G:Lm1���\A�	T>���y�U�'�,�����9HZB`,�r)I��5	5԰�
���5��ꎰ.W��*�ɍ��e)|�I��)0r I=%�������V�5�
�R9^I��=� uTCr��X0C���2Ms��}Cڢ��R�l�}�O�Ӕ���27�M����C��
[�oG����U�YQ�Ӑ��e�5�Q��<5ݏ �q�!���[f%�6��R�EO�$=p��D��IVҳ �
�vT� �ߑP)�[�K�m�	T�b�S�`gy����S�[��(�
hKF�`��=�Td��~����]ʧI����Jz��39��T_�G����2Y��>i�,/=��J�?�GOS�ocO*`[Jv32q����0�Q��I�  F�ψ9=n��JCB�4u,.Уz"C��j��V�a�L�F����B�\3�S�+�g�%��
�8��È��`�);��)^��O{��y�f��H�4^�%D�J;��pY��H�M�,�a ��E*3����jUYRU�kK�\:w��9���.U�����n``�0���m��}���7R 0x�D����C�C_�!e�BX�	˥{% R���(��2Oغ� �]�/��'�YHH�С��p?Tc��VL*���0����H?�!��j#�I�:�r?�8!������TN�tY�4ܕ�'�7-J�1�r{� �	��T==�AX��7�DQAf�f�,.�U�&��݁�8�th`�SWa{�/�_����{����IlXn��ɪ��ͫ6/v�a�g�=V�g�YW�geD��A�̬�<��e��]e2(�"��0q��o��Mt�HS$�6�I�뚳`��9��v�74wY�__2�```Ѣ�js����;?�ʒK���$]�l�� �_�C",��wDh�<���<�"��H��D�R��j��_IC�@�='-=�p$ ����G�9�JW!$�$�����9^
�<祼H��'���+��+F�k=�s��N]x�*o�H� ވ��l�G�fb�Eʠr�5��ޘ���P+B����v��k��f�/B+���m����I
�������3z���ؚ�e�x9�;��U�.v�$< ���E����t���%.��&�;^�ң{�j3�X�_��Ǖt�%��@��������`q�"���D�%JO�=��"/R�[q��wS�׹�H��׫��p�����|��@�E�v�����mz9@���f5]x ^'�|Ct�)O���o��
'	�jp��'3�å"?��,\�@N�P��?��,U��8��d
'�I&�\�8��r0Ny�1��9�滩,�ǵd�"���ML��6]�9� �� t�!�,�2'9�����,y�U����J���9��̜�g�rx�,_��t�&t�0��"oE��T�Q�nT��y�J�V��'9���#��7�M3g�:0�Ia��`��>�\��
�'q*�wp�=@�o���Oj��	8Mq������b$�7�6Ua�r��w�r����
Z�n�������;Ƽ��3��*�&@Ϋ�kw$>F %�,#p��z��CΠ �
���	C�[�L�A�&�k9YL���F�kS?[F�M�@
Z3�"w�y�5~C��D�B�J�*�F�á�@�Bxڕ�fF�"��T 9�ۤ�����2��To��H�H��5�5*'j��9��vs�ӯA�
Qu��AP�n�I�ΰ^R�� ��@��2A��s��4�VKK�$����e��(�*�KR-�Tj�&�!D�؏LR��$�x��ZI��rT�x^���W�r�A���$|�'	;^�
T:�Y1�^y^l��u	g�ݞ�I�X�y�Y�V�(H�@��%��r@�t�0Y��:^�_��V��1�i��-�#Ӧs2�ao��29o.r��_�&�r�X�0�8�{� ���������Z�{�d��&¼�~�F孚y��B��Lr���x���=#��`�^XJO�s^�a<�da0(��,�K��V˼�2Hʟ<���z�r�Z�O�׋��{��z1nM ��2�,�k��'0,���9]~$O��y��[e!3���$]/��䭖{W2�����ʹV�!
2+Zݵ��W��W'>�]&H���ؓ��CLE�@
�V@f��܃x���bo�&�lP�p�p
a� S��0����tC(�a�a�χp���HƼ��s�{��d΀&�/���y �7'j����Ѽ"�N&�������>܂�ޤ)8y;��0c�pƆ~B+R.�[`��B?Y ��<b�APpl�s1���=o�a��Er������j1G���ұ/���-b��f��@f�YDé �=)�7�Z�x�0� Æ�����)���a�IX$=��;���y�������2�\y�0��޻6�Y�Ф��FC�
�t����
�ވa��`�ظ1����-0���z�.�#���-0�R������S��1ś���,�&l^��@�S��I3<o�0\��H�4D��h��EC�e,92m�'�!t'bNɢ_$2�p,�	ڏ1���nd���T�����72���d��H�"bN#����K>CX�[`,=�q�2i�ڸq�/�-0u
˱Y!>xu�y#��ҙw�����0���j��]�H&ț	�[`���/�[O�b܈a��� H���Af����#d����7b���!��O
�~�=E�0�򮂒��MD�<o�a��x -�>��a�r����YX�~܈a M�,|ؐ�nOb6/߈a�C�>$��@���@�ў��0�L�H΍��1�@?��f�͔.Kz�@M���Ё���-b!�}�W�,����T1�롄���߅���x��`9iX/BO8�)�y��`9,���0�=E�0�>� |*���,"��夁�:����-"b,�8 �� u�JK9o�a�j�wb4H!�7b,Ǌ��*�P�\2b���:��4��c<o�a��Y87+-ݴ�>JF��.0d�}��Bb�2bh���ܧ�T��DF#�9�p ���˽?�� a�6������A�*X`�R�'!4/��a(��Ɠ<�51�$������t]��F®�n��r��<��Ðv�4����:����Ǟ ��_�\�P@�[`L�|R,�Qz^x<��"b�� u��4�!bI�KR{�L5��d�0��W�ƣ
Ƃ>D���"�*�	ѝe���a�Cli��q�+ˈa$}J�Ҋ�k��!e�0���ab��FN�7�����6�XVF����F���%��7=BϾ~&#�A��ӂ��&�_C�0h�:t����ч��]D�)DP~\@	�T�0��n��e8M��y�Ì�$���U*�[`���TB>v�"�Q�|�{R���T�=o�a��F*�̇E�H�y�Vnϼ/Q�ٴ��T�0he>o!?ώ��Cy��P}�ט��O�h0_SP�(Ƭ
XC�nZ�Z��F�z�WPY�S�Y�����a�Ӻ:�,xp�|�P�(d
^�0����v{�"��G7^a�S־N����Ӫ�a�(­"�����[`E�݋��|��9��FQ���F���+]�'ވae��W�\��_k�[`
��#����^�"�Q���t;'U���(�C��C>�x�-0��7����C@A�1j�͈a�]���w�{#En��7bE�A���t�<VE-�R����.�WE~'�6ԮT�0X���ڇ��k+:b�_� *W�[�OG�<-�nE�8'5]�d���0�� ���͔���6u�0t- 2X�	�����a4\���G L�RG��"i#�^�Zy���P�g�4�7i�<N���n�ã8F��E��:bM�M�C�I�|\G�� ���Z�`0��F#�
��b�	}ݐ_C�0�KLgc0����|ܛ����p\��N�0��Wx���̯!b��AXJ���Y��SH��}ZG�s�S(_/:c�? (��EG�)�w+Z��O��7b�B^jxT��FG�P��Tm�#h�ĝ�F�)���$�ЪC���`
냰F��}7d�ܯ!b�B%4���H��1��~�F�p�pl��00EȻ����}d��1��O9����yhU��!1ZUP�x����-0ZC�ӤL�y��>�<��"I�-���m!^�M�0���'x ]��yC����(��m�DC�Y��oy�
��M�0���=���.�h���a��	Cw;��Gx�EC�ث����:�����-��y1T��{�����A*_�6�^<;  �!��Z�_o�0h�<8���>@q��I11��R>䧀�8d"��
��c����!�2�ա�`"��O�zwep���Kco�0�����v��1��� ЇR�a9����-}l1D>B��}_c2��a头�Z�a�?3�P�#�4h"��;&b0��
9A����_s4À!����g1��-{���ᢔ�]وa�!��
�}y�N���Vz����rL�g�B �sΖx#��n
0�4a\c|]�Fc��B7��u?>^؈a����-�p�ҭ4�y��2�Y���������-0���3�!�)�-ڈa(5������)[l�0t@,08�H΍`#�A	�R`��-}������6~�(��F���Y�0�|��Kxޏ+�T�z#��OVa�B��>�yc��&T������1}�0LA����+9���0��t#0�P��~�F�)lV�R�H���ڈal��X�� ��t�y<Z(�~\�&Cn�P�!��ħ�o�a,}� t�Y��1��.9܁��m>���
{����LO�����l����C����~�
�Oz�������`�Zlh�.�����$�?N�Qh*�   	pHYs  %  %IR$�   �eXIfII*     (           >       F   i�    N       %     %      �    v  �    �  ��    x       ASCII   Screenshot�Ē6  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:exif="http://ns.adobe.com/exif/1.0/">
         <exif:PixelYDimension>1190</exif:PixelYDimension>
         <exif:PixelXDimension>1142</exif:PixelXDimension>
         <exif:UserComment>Screenshot</exif:UserComment>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
�QM  _'IDATx�����e�u&���r~�*WWu�@w# E�Q�@�I�PqL���F��x4�ƿ��A2���4��E��$J�(&Q�$@"���+�z9��o�s�+�� W��U�޻��}v�v�A�_�j?}�Y����u�px� ���s��9�N �n�P�R�R�q��!LMM"�~� o���x����ȋ��u\�� ��x���ˑ��˷�G��~7��`�w��=��)���@���z)O^��s����m�r����m�˼���׀��-���ʷ�����Gt3�V���G���!D��f7˻��ŗ�`{���NS�S����ێ��w��4')I��j	�Vn��i#!����y����*�Qzun����#����m%` h	��#��#�����D#��ݥm,�r������\D"���x���2O^H.����s(@��]����/_Gz<��{�y���d&����i��>���H�o��(��X("��;N�[eh9�>���|����.��>�c�����x<���� ��$��"��'���^y��&z�5�%8d]/�Eqc�`�`�z���bcu뷷�o:�X_]�Vy��KX�m���h��ب��Cm��r�c�Q��8B������"8�i`��AT�Un6�f��>�-JT�HEH�bX/��PM#\t���?�Tp�w�ܳ�`��N��v+[���r }��q����%�:�y�:����HO�����<���!��.ʭ
��'F��m5[X����WWu���?��X���N$�f��V��0X"��N������sO�Ca������9�SY�	���
ڨ �q��m�y �^a%
*��Y�0Q!�f7o�F�YE,á���v�ET�+xu�wT��z�pA�D �wzt���]xܬ�]rH��
�v��o%У�Gȁ]s�n��P�Cé�����(9;h|_D�����d2�=�?~��(�����V��=����J�K��FQ[(!F��$ލ��\2�B��`����]�yW�x(�={X���F�JM@Y��Q��G��"_ȣ�LR�]2bK��:��2d�F���B�j���{v�x����|�n��L��t��/V�	���-�E� =I�A���j`w�H��b ���E������͛7T-\o^E6;1@5��b.v�����'6%Jq����h6�<�[�o�12��.���5���o���d�4�Юp7������)��x�ᇱ����/�AB��>I��j�Z�arrRkssc�h��:�r����m^[�}"����Z
幆�J��B���L&P��1?������(�$
Ky�6ʨ�+p�n�.=������z<�k�g>_T�4�ud2�l���5�&S��&?�PĚ=�@*_bt�J©bH��9LTIO9S^���&7��J�����W���Q��j[\1�g����:ԳUJg"�R�1�$��!1�"�nK�'�_�B��	�l4u��\r���{\s��Uu�M�TJ�n��ި�3-4�M=䑑��r��)�%(��j�!	Z�y9��N;�M^���%����˥�~NU����4`�;u�"=�eT�5݇@����R�JcGԡ��������:Du z��'��Y��7��ۭ���(�� 1eS"�bH�\�H�\T�&�Ll�p��pq�MBHAG�@��0��M���_>�7]�/\���u��5�h����O��v�����6EW��(9tEQ��=E��	d���F��f�E��Ԁ���޾2�|h����WIT9�`� JٷyAp�%H��5S�ꫵ:5PI�7�y�d�čf��	�؏1��x���L*�pp��O��r�O@U�sϽ�������m�Z(�Km����\;7;��Q�E�р������'��q9̫W��8xh�r����!kZ������ ���\{������9ğ{*m=AD�gTY�KʬolP����a]e���GU���<3=��R�Vl��%cݸ~G��zM!\~��z��mU�vHTx�o ��u�h#o޼��uv�>%��ذ��m�'���Q2䞡�c@�wr�.�������d<�����o'�CX\�EݘU8|p���_���2�}�e����4Y'�{zQ1ΧNSB$h��,RT?�}��x��)�!�~�H�=��\��-��ʥ��0ff�� 3܌��3'���)��r�ģi,,,�;��r����p�+jkz|��"1r��(�5D���?�G��6��	ID��/��._��}�f����R���:��C�(u<@���=�LR�r�6�֭|�k�&�ĕ1v�w�`�
�=LOM�^+����o��'����C��>��/bk����X*�!�����<s�u���	�F18TMQ��<�A��'�8Fs#T�]�^H�Wxt��,-���x���H��jSb���kh����O���#��v�2��2��|׻��Cz;�򕯐��ó�j��.���o?�o��ǥ�q��y�8~���M���S��e�a�����3Q1�NW�QJ������{�`����T*<����?���ŋWx���L+a
���A�I���O��'I��^|�D��AǨ���'�h����_ s.���U_�R�������;E-R�=*#�J����'>���2�"^z�|�n�#�Օ���� ��ҙ��!���a$y���?�y�;q���T���?�S<��Gq��	|�[�����O���P�
c$�����
Da�Ŀ�w��۷o��u�y��%D#����<���-|�S���T@A��)�ϫa��>�	���C4~E��øz�2��/P��q��YJV����DU���ۮ:	�k������WH�#��$�\�I)H�a�q�,��x�g�L:�@�X����'>񯱲���>�Cj��zm���\�t��GIp��.���Q�:*���/��7�ĭ׉ ��`����y��,QZ��Mr��>��O�G�6�G��!���C0B5R��<�/��E�T�C��Qr��ϡ�/`�����pǕ����O`jjL��y�5x4�}�����>�Ko��O��|;;!L���c��1�,-�Fn�ݑ&W�q��|��R��P��?�{�:K.�}��/��W�����a$����(�h���o��o�,慗�+W	�q�3�8q\�������?��ΐ��я��×��O���E������$�Eg�r����74��/�/��>����\�z���G\g��{�kz/?���.��[�M}|�	?����>��������,��s�#D�����/<������,z0�|�mx����=j�m�2��� ���"4���v���/`}s�4/<��7n����T7�Q,.o≧_B�Tñ�4�AΫQLŸ���k�W���?��x���ͯ~�<O�����_x���*RT-b��h��r��}�ӟ�}�{��J]��� rڡ�������ۿ���/�"^x�Uo�<EPbDE�����w=�N��?=��n㮻߆Tfo����/|�7M�9��9D5*�����6l��y�d����q��n���5J�g>���\F�I�΢�ħZ[��?���W����@��J�%�t���G>L?��ߑ~.����.�I#��f� ����C���ue�*�#'N㝏��n���>��o�:u7n��D�|?���������a��ir_]| B�j�Rڥ�����E=v gi��W���$��b}An��_�G����*��]�ve������+�x�٧xͼ�+���N݉�g�����]|���P��Q��V�%����+�)�:�o��
��	�x�'?��������@��.��_�%��1�A$�@�X�]X�7��M2ٟ��]����.�-�R��`����}T������~��s�
z��s�؇?�H,�O���A�;1�B���w��]�8uU�1�{�u��ֶ
Tk9�����)�NP~)A������g?�/��7���oý�=�zySo|�}��������r��TL�Jh}O�,u��¶��&u�_��g�37��� �Y[��"��Q{s�OށX2�T:�n����Օu�����DHi��Oࣿ�q�艧�E�j�������B!��M�H����_x��{�vo�j�2��/_�/���C��#��!L�=r�(~��������gp��4��x�x�s��+�d�6O�	�Ø$���[��O�[��>���bi��8u���.Q�������+��q������/���)m�v�^�4�������"ш|x�����i�y� ._�F(�0�����}��m���\�%��S�D	C�"1��?}�e�K;�!�Nј�=� 	L������j-B���9�}������d��h˪%���G�2\0��j����'�$.��:�6��Qe9�D"�Θ �Q����k���7j`�����UI�ѱqPc���
�g��Ѱ����1�,'H�>����(�������,�8H'�J)�#����ډ_%�[7�i�?��}�������Ԩ&�Dc� Z�Fơ���SU���&�l���x�G�H���(.^���"@�y����o���btb?y��X�q��;	!�EKHB�����*������h���~���<�<�S,Fn|����W.�X��$�o <�J�)a��e�x��/an�	���F=xy���J�2����./X_*�*N��3w���c�~Ý����}���D���F2�Ņo�����޼|]��\v1rw�Rz��<��M�ƱSj"��؝���y���E��38O��i���S�r�߼L��ާq�}w��\%���6��ҹ�	���#��;�U���P�L>D;=����;Ͽ~�ܸCNi�;?|�n�z���7iPc�D�z��:K�dRC�R$�x��M��>�����埿�:�_:=F����j,���_� �}�܅WνA5R��9�^��Y<���t�6�I�r�*>����G>�K��M|�K_ㆎS�%�M�#�*\�޺�M;�� ���s�y<L#��3/"M���|����!.)Bz���M΃����+��c��qΝK��N�Os������O����G��*!����\��*��O�z�h�Q=�4;��*�b
I�6�>�]����ʁx�I�Q=�0h�����t"����q��mq�4��ſ�����D��<7�$��7t��&PF���\�z�/���8y�X���D��++$p����|ϻҀ�@�*��.!r~��{�>���#4��B�P�K��uL��!�Tr9�M�;$�l�OD��y��=�ZHPM��?~�y�<��K��ƛ��G?���6	/pY�F�P���|�N�;�|o�q	�kD���sc�b��^٢y+�k�ܡK�LdԮ>������.��X�ʼJ9�Z�җ��k�tv߆W^���n�&!�0A�7�Ik��$<"~��vg|7��_{��O?��=����W����S��Vn�R�z$�[����.���m<�ػ1{`���+�"O���h�j夆?.�q�hJU^�궛�����>������?�v�D��G����r�����p��䴎:��ʵ�!��kׯc�������-�ԓ�ރ�G���W��m4(���{����e���2W�ܼ~�h�6����q/}�������?�n���R�h��X��닄�R5��Qְ���g�DcaB�Q����H�2�ڣ�ܡ�>�b��&t,g��<1�݅7����Nk(D��s�S<��x��m��9�g������j*%��Ө��6ַ����ƈ��xU&�Q4#���o�)����/[l�n�B����!H+�R���L�_(���1u����C�����ښ�\�?���;<�ťwLІ�a��*��饏d�8v�b� �%͛���$�|�:^{��%�bg!�Z�i��������G4���SO=%%8r�0~�����[*M"�f���3	�~���E*�o�N���&��&*��gg'��_�_�hJx9�E�� 	3��<��ьFJ	�7}�c�Ї?@����V�w_G�FPB'��E$�������R���P:��l�3���ѶlI�W��L*�� �<����R�U��~?���%z,@T�u���~��
D��b���x�FCPf�k�j���ٓx��h{�	1Ŷ���Duu�7bG{�.^^R���~?J�M94Kzn�/>�%�>-��+2j܏N؍�ܒgrPAE(|G<&:-���W_���r#9B��XO��V�X�'?�y2Kr�� ��d�D�DW?��S��c��ƴ������0$��x���Hƍ�5�6�������c�C��y��;$w2FU5�ͩ4m�_�H���ց5��'jJ��`(d4?+��Cf�,��T._�G��f����ۄ��ڲ#��:�P���2Q���W֖1E��%Sx{q�;���\�O�]	�
#����	�ڒ��Fy��P�*��s߬&�$�-��q�^��m���	���ݑT�H��l���|�z�\x�1D���^|鼪��<����,��~�$~jsa��`!?�a䫯���b���>B�;���W���1!��xAS�0�&9{^����H�������{��
�˚��X�1�x�W��sz� Y���7��nW�h{W5��X$�v{�����+���(�����Y#�]շ���~��)(���E]�f������Eu���Z�j)�T]�E��T8��Po�z(�:�Ĺi�-��q���&D_�i#��]�4�􇛐����ǈ�����b[��$B �I�P����&���8&c(�Ė�IB�l���a	
�޵�0M��O0�~FurhMR1E!` �XW�R��Z�F���a2O"Rc/�!ɽ�M����> D�d_>�|��6�U]�f��!A,FKqyw���bj�s[y&�_�!RLm��|^?22j8�3�*�pσ������S QJ�����D�k�5<�FE���MՇhW���g
����OD�^�Q���4����G�/��ŁI�S���4k��)���|\5�gD���k�lΙ3w�=ب'/5�ٻc���A�7)H4��JS���g�Hn���=P�{Q�n��w�F+��K��F]AIb,���E�J�/�xbOgzoY���^�`/2t��w��g�L%B*Yz6�ag>�)��B�'�c���;�<e�T�4��+#n��k��lK!�@U����:��5_�(��C->s����a�XcYn8�����-����́����8NG�)�e9R�A=����p�����~�"���l��X��$��p����:�p\M�ch\����u�����<p�FH���-vP�h<L���-i��{��t�/�-�q�k�ޞV�F*ݠ�
��v��b�~F=u�`�
�e�(�PG�߳��	=ǈ�,@`Z�P�p_"��c�`��>7�+�ƍt�Y9z�R��:f�z�B�"S~��0U"ZH!�|@�ׯ�:���	�5��_S� ���u�@A�b��R�(k�aLlI�f���2� ��Rð�6�&����բ��u���z�H�a�o��i�Y�0��\S��d�z���F4"x��=C��F��hb+��58ڨ!B0��JGC��OoHX���6D�s���QH2F��Ј���o�ڒA�翂Vq��A]��h��z?������s��º�R3����R�U��љ�*+1F�)t�Z��'�*�*U�7pm9�)����"Zo`�`PD�j	�K[?�l[5(�ּs4G��O��զkߠ�P.���{�<��6�V\��eBjI]��u�������u��f�MKg��)H��#��Ʀ������B˒4R�F)ʵ�QX[Q "K�{�A��.���4�6�g([io`v�J�Bր�{x���;��Bؐ�Hk]��MJ���p��I�g8���6+�Р������I�_ю�S��������Qr�4�����$m�u���]Kq)��1����zU�Qo�qNZ6����W	S�"����x����]ulKtҒ��A1*�}-t�{�op|WB���-�f�km�c�A>zZ7l�d@����&шD%Z��{e�<��E4$eQ���g�߼7h���$���EQC�94hC*gL�D>�H³I�BE�0�~���P2��Bu���؊P4���.6*O C(J��Th�,���x���5����d�v]{/G����d�`m�`(S�����T���i�����
Z�&�oD��C/��T*"��)�bRa��BE�"!���>�8��vQ�����a8h(빦b��w�c�-j�uL1�����J�r!�t������ħiQR\�NZ�

[z ��Q����QY�Pj@������w��O����RW�d9��}+?�o�m�Ѩ4y��_k�F'Z��WF���a3�����ڍ.FƲ$��.=�G��a�C�"�J�'P�b9]�_\��(^w������e{c����8����yo9\��ֳ��,*K��1�d�)���D���!���~��ö�o���iN&��1����i߲Tv�}�vi��9CƲ��gY�J�2�X �	�H����M�F�G�ǩ�ZH$B�C�Cc��M{�D����	����^�5Ҟ�-��k�!<�LY[��{0��J�P�q`U���ª��&%�����^��=�Ѓ6򍽆r��j��5k4���]T+�DV%���J�X��~d�ǂ�<�	�{��������n{��BJK�"��	�� 4�ti$�z԰�qk��b��0
Y�It�Q9�L��#�k0�����}��o��XlP���gC#���z׮q���~bGZͦ�C�>R�h���p=�2o@�nת��4ĳ�N�=�I�`'���Z��al�4P(��p���������w�a�ֳm
&7$-yb��4�^�h2�ZZ�����������Ъ�H�s|np��h �O�"�~෉�P�T�Gl��՚�X+7�[�Wlrˠ�ahe`
�k�$�q&i�^{|nҶ��׷��=UdB&��.�l�t
gON#q��RI7(N�����o��dꥄQl!��򍾉p[�����6��#�ۜ�`XbJ_MC��,{k��1���x?�ݍ��E��D.<�Kbn&�����є�m8&��'��+��W��N/�u�L��2#�5QQ��H@#�����WH�i�K8ƨ�H,��+OпHhY�pq�"-��Զ�HCd5��7L�W*A"�b}3oS��Pzʑ0��|���|��SI3�j�T���9@�D�~dª/Er���!ɻhT��zƮ�$������P�\@�Z�/M0QJF�
���!����1�$#&��d��g�&�u{i�V��1�����MM$��bfȝ�B��k#�j9j4��h7n���sTSR��D�ޕ�|5��V&�D���^͆!\�X�`] �Vl����Yd<�w�'M?��Z��gі^�6���:���8��:�ծ:w�xT�O%5-~��������؍^��U�gF�[h`g��='� ��qTJԎ,��h�XZ���]��}C#�g���y�z�����70NA]i��=�Z�TD9���a�NZk;�f�V�H�&4�#e�RHO���	����F̻qI:Q�k�*�'��+�vW+�At�%�aw�F۳Ϋ�������}��_E%��Qe����9�b �j����m"��@"NF�߻�[���A�����Z.Ï3�3��n3^M:|>�3~�V.�hI�^"BU6p0���ԉi���ˇ���s�kc��������z�B��;T��P4��a��,N��ʎ�ue3id���,��c����iR=8���hML��}��!�V2����e� �5h�C����w��"7׾�啦�A���*uV�w���w�����&��X]��}�I�CԦt!��|�^�4v��Hg��,�1�<�8��P鉡�mZg��`D2�R�&����8��5�!Դi'd��ѕ����#�0��#�ʁ���!̶]��+*�3őK%���5mC��*jH��\�[	ls�Y�AM��Bk?����JР]���R��Bk���.���j ӳZ��O%���=�D88�|@���?�\�՜���Z�4���ժ�y��mG]Tr�m����}��NM�/�M|m��F0иo����I�ec)�=$���D�ެnua곌/ !�e�Z��ORi8�u�I�6	R��M`�<Bc(�$0�G�&�7���9���`i�
�5͞�em�xg��A�"Z����o
�aD�._%���	Z�w����pM�O�9�pb{[j�l0�P=O���4�c�=YsO�>D�0:��m�mDX���0D�Ʊn�T��:e����HzP�,(9�V��zy��vZ9FC��n����jn�κ�Qk��7+Z�_��]E-~:w���w��/8C���Q�r����	,?�h�*�O�H�>L���4(���|�DR=�}~y&l�ɮ@P+O�`T9RS*ׇL3��-z�Ė�F0���̠���q�"���|%�p��)lW�J�u"�7�"*�W��W�ֈ�v[$�GZ=�$��^��ã��U.�"2"6��HDY3���~@=Vs	�K?��E��@���M��S�5�f3s��/5�Gj���=I�d�0��j�t�h��uT%z0��x��k9��=)p0Lt�*�&���acu>݆�2if�C�7�pc���ܸq}FbHڍ��K�p����Lxhb}����� ���!�!�h`$�J�ť"��)Ҫӧ� �?pd��e�L�'��A�-65+�_H93��zay��9ȏ�Yx-_)6Mo���PE���ӓ��;tX�զ&��)A{�wv$�=0R�$ �Rm+\O�3�.W�Ӧݡ^o)�z��Q'	.YG$b�x��ۭ��_S.��m��w�=�L;������-t�v�҅�����AX���e+����Ⱡ EB��X[��Ч��p��8�vI��T���T��`Mx��P�5�Ms�[��#h��8z0��7z(LM�x�#������`/N���IA�����t8����}B)�&��ݹ�$�\�h�٩�Sx��MT��C��rP�� Ky�{ш���\"�J����+חq��4�җ�u���?5fgxMI�_�&�ڮ��&���F�Y�( ��O�`.�E����"�i�fu������k�J���1��Xp�Ĥc�Į����ӱI����nM��봸�)\��Nq����q���b�A�\���bn��][��@=�`���Ja�FQ���Y��a��"!h�~ݔ$9<x6E�7P�H�[B<��1�2!D��E��{}m�d��,��X����$hiUq��x��<U�7*�
�O{�c����ЁV��9��'���ub�vI;���t~�ȴN�3.sJi'鄁��a������#X�LR}�\6E����i���c���#�Ih0q|2I���&���׊8sjV�{eY^�O�����P�W�KOv�������u�� кV����y5�A[�iS�j��TaR@ �ïV����/���*+?B�p{a���F��J��T�!DUMN��/��(��J��(e2+�j ������S=K���k�Ju�6�g�������щ�H���$Ѩ��W��G�ӡ���u��ٟ1	*�Lq5� �Ob/%�j��e�����v�T��D����Db���lRu��zw� �� uh�F�E�{s1:NM��n�H�� 䜛�\zG������R4K�C�*3��z�TŴ�F���cT��َ�qQ�D��7�~]Tjmm=�B�]���p]e웜ԱR�����T-AB�0�/�����vp��ZtN/]^���<�4V����=]��������7�v�I8ǭq�yȀ�$T�Z�D�vc+�mK!ܹ�$��:�K*Zuң'��s�"s�+��l�nO���_��荥ٱZo���Tڊ(�]��0�,�u)���
L��jʵR����. ��Z� ה�?��>71Ľ*:����g4C�i����l9�RńB���!�.j�0@����`s��{i�ȅo�܄G�xeU�z��kiu��o��JU�ѵƥ�k�O���P	�����}�XZˆvj�4��o���Oz��sԺ	��`'��� �ƕ��	"�� �:��C�(�9���j��(-�P�ȍR'��ّ�MU[�6�w�sJ$�,��To:AN��b�ԷzJ���6�!�l��=yZ��*&e�Z#8���Di���J&R`� ��HQiO�C;*5�R�$a��mL����n��u��ZE3H	���0*�[$a6h�5~v��a4:]2"Xɫ��y���:�Yl�淶Ph�P�1�����5�#�O�t0�ۦ ��C�d(W��e��V�M�;f8Y�]��lЕw)n>�rT*�����K᱌=�b�옉�&B�H���=XoS`�|�u �
F沈A���S��=B�pK�tGG/�ܸk�S�L����	i����O�dB��!����KG���:�d��N�0~��ՈF
�����*U[Â� �MK$�hWf\�8�qڐ;�'J�ҭ��h?B�i�wH (�O&5�T�
�ı	�	r0�i $��Kz�c-�D��h�Q%C�ڤP�͈��炈%r<��RT6�8�f��#ciTw��7+�)��H�@���)�FVL���M�2h�K���W����P���F�iY� ��u�_�i:�`��I�`@UU��l�`�p��B$v����u�q&���p��v��
�+��l<�-�˷W�`����:`��mR:r��zC2e!1�u�.N���A;�����:�%��H���$2�T�j�;Hõ��WC���;Cu��^�@j�����/y]1;�C����Y�)X�*;M0F��k#0�����Ƚ�2A�i��<�T&L�M�6N[E�M�x�%:����H�iKXuV3R90����I�9~���T�ym�����r���x�:�Yt��ё��Q.ޞG��4�^�P�k�sJTM�"WD�!�l��g����ݣ�Qz�r|��!���12��=�Ņ~�$�����#iL?�gBX&�m�t�~5AG���)w5��X�n6��o��W�C�[���L���#H��W}٥�b�Z�3]{�Tөt��d������lE�@�\�k�T&���V�jM.>hT�D͍�������Ҙ��!<�@�[Õ���+?Av̔5i0T�\�Ѡ��SǢ膖���H&���A��`�&S���(�k�frHfC�uc�^xF��Ĥ�=���פ��8ȘL�t"joL�J�����鄚ܺ�8ÆLAZ�3$�����!�%�8���I`�̵���`��ϒ{�6�dB�SY�(�2U��:�o�6qG�3��G�$FtV��C���g�ٌ��~��؅����B>"1:[ү�xd�>�k+�0Bdu|�	+2BJ4Gp`�s&F�Pr�P�z�>�#_����7YD$br&��Oh8''3jL;E$)��~[��I:V
�h!�����'�Hg�!�:�$�Z9�`OC��4��W�k��__lDӦ�$wx�f�
<�H�G�p���y���
�� a�Gi����~Ҙ:Y$L�Ғ�)�NGm�z��f��*��Ï�H�tv�8����lG�-�~1��:Hvt����whrN_�H�����`G�NC��pA2���Kh�!��i�L�P��A=91��`��d)��&%S%��m��~x3ڢ�[Q�k��5�~��FTmP�5�8������Oj���
�X0~�$�ԇ�� I�J�49�f�L��d�TQ�J$h�Iu}D��~i�Y�ek�&�JO6z��iW��T�)A����´�ct�+kجl���R�j\+���Ii���4�S�6Z5$B�h'8T�����"&Ɖ��B��������*��b[cD�6U�T̽��z�n�$�B�ީ�#2l����֧5���X��������>�>ϫC�(�+��t��1=1Bf�R55h��j�$�$a!	���/�M�s�5l�?�V��۩k���/>Z����q*;�ceW�얶qs=B�G�SUf�}	e��Q	K>r ���L�ϐ��2�26��q�k"HP�4y��)l�HU�f����Bkϖ��J��hM6m`��m\�+y R���̳�2���-��C����۫�������Ri�n�t�ã��>[�VVJ8F�zH/��`/��C�{�侤�vU骵ջ�}0	)	i�y}Ǐݩ��jmcN"��k�yiR	���4h�i�=�1�V0쑻+�|�Ag2r�7�*��ɨ���g�!\�t^J>_�<ěW6鄙�Qm��ܽP���#B��	�WE�=�x�2��t	�mf�^.]�Jw4St�ز$�V�'i��բ��72��5� �p4�uh��;�M*D����56>�k���l�̸�a��ݏ8�Z�M���:e��MT)1j��'Ϊj�J��8����|S��69�]k!�N����D~'ƒ�Ϧ�yr"CL]׺����;��H�������(1�x�w��L�]gh@��.b�W1��a}�jF�d���a	��S�����5�w�}���D	����Qf#YmT����tW�*S)��h�|%S���ʅ�Q���N9��FZ,�^����Ȑ��8n�o(|ϐ�"�:��@�"�]�]����_e�';:(��"`W��wP�����ɼ����$NMU&�A{ҖѲ�Iݾ	;��T�JJ�͈mM�B�o2ܐ@BQ#�)lue rHs��OF�T;�(ſ�n���ac�J�$�\�+�03�R�8ʃ�[X lh�S���!�h��ئ�d�J$���sW��Wt�ב#y��A������g�Z`Q�$�B�>��g!5�ժĜ¦ЦoS¤ENb[aT`ccS����4V6wq�p�,*���[��l�d��S�ȴ���A��u7zd���8��ئ̍NQ=e1��@糄���6VAxb$#�N#H���r�NaP'4��Vf��M���핒��BK9��)L��/��D5$/��b�����Z�*�L��J��g���U�ak���$�---`�s�kh�8�������/!Fn�IX����S(Rut���]Fm�����M;����b�R���fYs=;�e�� 2#2	��r�e�E�k�I�����r��nU�(���MOĵ௛ �0��|y���1OI�z�<*��c}�v�(����T܀����0;��)�Ҝz8W�!1'))m7j�_�N�0�u�!]ݞ�Ɇ�Պ�G{�����\�-˥u��|[�%�y�n,T��L�1���b`��Z\!�%�o�`�RƔK�#�u�ˊ��GҪ�:��T��5�k�`�_}(%�yUc�rg��,-�Z�P����tm�	��.����|����x�SNʃs�j�L~:x�ܫ(./!X�5��ȷw�U�L��T&���'�S�_);hC�E�+K'G��mT)�"��m�5�cR)Q[�a���L�%	��ͭ���bq%�&�[�@�8��M��9~�}����&|����z�פ��E�!pV�&M"��T_1/�Au@��~6�֦$S�2�v*��G��+J�#Ou��}A��bMU�L=
I��-i5U�"=�����z��DZkZ��蚐�3��O���pj?�q:��ࡳ�clt�;+x����֋����muk��YF*l�a�=�zǒ��g2Q4h�G�L�'T��'0_�SG���g�5	�u�9�"��vˣnmo|��:��"�U�"��jӌT�����P�l��}ztXթ����d����j�!��
v��� �$u��X�\��Ri�,�㒞�A���a��$4��F�
"�F���-Th�[-�b3� j��=����'�� ;3�*5G��C*�Dh�'�t���U�	���9r��K��L�:8�Z���R�,U���k�ym%��XK�u��,*��#ݯ}=�H�c�N�!��"�T����p S��'�<��զIڧ��9��#�g'GQ�_F0����vq�N]��lx�S���-|��Es�E�N01��֕&� ����y�����G���Hq���'�ٕ϶4?d|;���p2gd�H�}nf�[���R�ю�����D%U=y�r��9J�|.�:a���%���^����-%0��@�pQ��jx�X]�ՍK���x�(Eæ���e��fH�9H��	�(�;|�q�&hww�-��Rh���:�Io��z�4�P@s:V���V�^�Nep����i�s1,�s�)���Ү�
4�6��iU��^nӖԪ-��`Ќ�Ғ����f`������z};�¯J��X����A�мPU_j�����u}h���}�� ����5-ͥ����՘H�������he��
����g��$��\UOR�!�b&2%h�k��zm$r	B׮Ƈ��3��0���}i�ݦ�v���k�GJcFң��Vʴ�(� ���ŕڃ谔uXqi\d#���kn }+��xN@oJD@f1F��&��0"�P*�����ŀ�l4Z ��"�T�/�r[K���˄N��-�B@Q��y��Qe�L"��G��3o<��j�UB{����ڛ����T#k����'�X4����}n�!a��<2� ��uo
�^�p�'uK�,���a���5����xo�ZűCT�94a�K�M�p���[$����܋�!�5��D���L̨��>BQ4l׶Ӌ�>���Fc.fgG4a$��J�o�09������Up�DX���H
D�cc9ڐ��(��͕��ixӓ)ܼ����neO]���EĨA^��,_�F�nq�F�ќ���稾�}f����S�1�Ƶ,��=�"��ݾ�r��\SPO��3�����i�cGbZ���phX�w:u���8>���r���8~|W�nֳ.�q��/x@�&��!;t��r��@{�b[�0Q���u�ð���Z�eJ�d����4�\q�BA�0���� �cKK���G4�=M�VF���F-
j<~xT����7q��G��B"����1��S�N���]:�V�m�S���%)�x�U�'W�Ua�(�O�f��Eb�H�@X/(N�z�"p�����u�5�w��w����66�kj���P�*VBR�Ur���r�9|nf�r������A�ɘ�Wa#�����-%umo���4r�1|J�Ø�K;1��M9x7���P�����J�>+�jgkKTd�=CE�SKbS�6wk:��\���
��3	޻��x9H��ę��!�ΤP���g� I����RG|�(�*�l������ [�m행s��&��4�U\Ñ�j|}���ߤ�3�6'��4�url�aF���E�G�������g�ܸ�u��w�Z�:�~�36�<y�p��G$�#�5xK5b�3�š�EQ��5���nL'�U�R��fJO]�PDu��L��U����U5�6�ʺ�M[��A���;�S)��.��<����)�ږ���ג#	��A�ϴ�����M������k?U�x��XO��(�O9���K���F%A;���S7ҁe�G���f�#�t��iU�%����v�%�];����M1�7�+ؤ�#e?�����H���?:����y��D\��my~�T���ƬQ�V���;f�~�������/Ǵ_�k��y�.�-������SJ�����}ep���2f�&���&�i�n�q��;������
�t�l_���Ƈy�uf_Ө�׵�Vφ��P39����C��������|��ަ�胦J��m��@G�d�L_�QN�x�+��� �S��6��^}�͛7�Vu4m�������l:i4hB�Z�(�?�`6���f��(ϱI/ǯ1���6Y&�1i�;�����_\۬#��q�Q�Uic�He��f\��R�ˍ㾃wb�5 �+
EH�)�biK�x	������qZ8&���X��Ke����:���0Ѥ��l���T��Mԛ5~�ɕ��k)��uEB�Pvmڣh|>w�L�;+�=��o�y�I�$x�%CBڹtKK�Z�(�*������^�����0���L���O/vT�m=�m��!v�	y�퉔G���3�K���R�>��BWo.��c��:G�K�"� tL�oC`�Rw�4��r��ՊJ��[�*�<&h+�MY�y���!�jǖ���6#�Pf���Ǽn��\z(�E I��P�(abf�'�����ɒ�9xhZ��g^z�F���N�jЯ�D���3D��]WVyV:��`�Tr��i�\�C��������:��LCl�{���I?ާ�����i����Iup���Ci-��d0c_MT�L��*���C�2�k��%#�+�2-Z�:��ˢ1���(n�\�2	Z�fӤ"�n-Ix�H2O�4#�-Ily\l���Uju��z"�>�:r
^-����>^y�nܼ�G��n��C�pwie�]������U�)�n��)2�'��m���� ��ı��
��5��D��?�,:��&��>��%����Yh��']Sm��Q�Q�����p�ZQ����zyM�YA��i�3�`V���30CȆ�˴����� ���d��_�!4k'}�V��F=љ�v~ө~IJR���d���Z2����C:��[�$d,cbbR=���m��ej� �2��J�c�����m�Ul��X�Xŷ��]"�:Y-�s6J[��J���$$]u$+�3��{���5�ct���$Hp�Gdd��΃Sg��,n޸I���O�T���{[ձHE�ɡSm(=fg�����O��SlV���N�KQ;x� ݂��íW��E�0�����J�a�:�
�L\���W��Ĕ��E=�֪�ʔ,��V�7L\Ďp��.�@�W^�E��0�܀T?J&��e�#DPatVi� �8�*���+7P���1E?|�����Ohh^�)�����:BO��{���%c;�9�b���][��:~�_wXL!!�Ly�@��N�R���~'L�S<��2W$d;�$C{ U���ڋ(�*��Ҽ���1.n/"O����T�z64/�kI���}`lcC�}4��Ҡ�M�G8��>���,���K/�ꥫ:g�|�U��,	vxr������eAH����r�r9z�qd����X�hT4A�cS�S5�A���pDob1�:�������NH�{����3������X�7��)݁���t�'w�={Z�_/_��mU	.��҃��D����ܫm:{�dBH���Zt8[�5J�/=��¶F/v�۪}�������Q4,��}=;�5��1����|�l�@��ɛ�.~���䠼�8�ҩ70��P)��c����+����9�m��U���&Vv6(��1��I����s�d"���M��������Be@��췂�O����^@~K� a�)�����)y]����O�1=>�R�j�7^G{Bj��NϽ�<
t<�u:��.=+N�*0���f�Ρ�j��/����x��v��u+�oE�ڒ���,t}k���2��XxgF�D$��(�J��,�-a�茆_$�"��������葈^�<j[ V"$l�������F�^�LNz.B�����kfݺ�� F�K(G��M	EB��&�+�p4��ZD"����a�2 &��v��
��M�� k�|%�j����y�iI��n����m4���i�R��uv,�~邎x2�m6�e�h"`�c��P�7��!��D�n�Y0��o��J��jc��R��jYu����v;j�%G�	�F��9��Gh��I��#�	���l��r�	�p,b��.})2ZUt�py�׹E'�� ����L��pZgІ��U7��A���h�K74��1nU_����<�N?	0�TkJX8Z��)@s���*qn]}��y���0I��`� C��azKr��[������U��3<a���S$c'c�d"6%���7��:��8ah��R�4h�i�͓��]���p_.�1��R�j��HDJ=Cn���P}�Q)Ut}�g���<lU=��hū}솔�[���f�<-�p���
W��5r�ݼ�N�q�<D��T�Nf]K�DV�d
y��\�~M�#j龳��M��A88w��G�n)�=x�����R�v(�+Ké�� f�{�<<��o4�bcT0�����s[�T5n��J��x,���Mm�����/k�jnzF�=w�:Cc#c�ԻE˻�Y��N$½s	d��%�,I!QJC*n�����-ז	oR���lH�Pn�<���p"��w�GXq�M&o��;M��O�Cb46��ҩ�_����ғL�@r$��VJ9VlQ�f(ŷ���	�"ר����J ���i�naWt�<z����M�3������ht����M����	o���G���;x�&r��R߇�̋/b��".���>g\x��#Z�a����K����mD�yO��h� k��g�������Ğ��ё�ڦl&�Hе�&��L:�
h���ȓ�� )z�bp#V��E�n��r����A%n(�Wq��M$�'��I@�G�VO��MMO\#����pY�c'�yJR�h�����%�2T& �J[97����ְ�(*8'x6F(����|q�p�DA�TD�t[�y�� fE���I�p�t)��A���9%��wh��k�y_���Hb_&�=��Lc騍�ZC�+7���SV&�@K�U���$�8��!�V44޳�fcc���Κ�h� �둟C� f�L����a���P�F֖L˫�a�^�(%i��L1C*��gP�$_�NkS�ބ�R�*k�0��-��D�ig���@L\Ǣ,4N;8��/��I�a�Ez,��DSc�x晗Ѩ7��>{�,�}�Y5���YA8RI?;=�8%$H8ۤ�i��j���n>4�F���%���ncE��؎���Y]j��G/���LQ��b��h'�s�x�Q����:Cz�ߊf���9�@݌����v5h�v~�LZ�Uj��'b�������79���F�^c/��1�똾{{}j��?xZ��?OO��`�SGO��r��q�jv�t��8�2Ν;��D�Q�FL�b�kw�l�y ��r�h��@���k_
�P�h�-�֧��15P�ʹ{SD˞i=��vx�]� ;k��у�k�Vچ�6EPn�)ˮ>��X*�Z�����#9������.�U�����-J����t��u�1/���G*�!6&L������=����ٌ��V���@g�Ӛ5����T�����s'��N���#7%Q�lAbw�<����-�v诸�Ma4j���`�v��t�_�n���xei�b�/�w�r)�/�L���b�����{]?�fJ�����5��봑iډ\.G^$�����Xn���e:R�(k��'U���J�zO�t��w#��lW�D9T�~p��"8��3�m5c���p��k
��R�Do5X%�Ӱ-�Z�)7��t1h�~��rQ��õKm#��ax�L1v�����\t����u�i=����cgU�A~/�M��c��f��>G�h�У�"O�=��Y��-u���`���,0p���H���D΍������X�+)~�«�+�穉)<J�J���6g�c}k�h'S��C�q�F4l�p�6��D�J��3��	�e�O�ᖗԵ'b���;���W_U#.9�q�~�ZY7(#$���G��/>�.} ������~���e|�r�c9L������юV�:�J-�]-�%��g[x�N�F����m�(�C(�/ s:�@F]d�S��>�/
�k"5��ș�93�c�`�>���$n޺���r�$!bI�xb|�v{*��5���5�>uV�z�g�qr�Er���,w�s7iQ	���s�1S�?��1(K�}|��:�d(�"��/�C����!���'u4�Ciye~WG��s�*պ��%5b%�p{Q�b���Q��n�u��:��3���l�����4v����A\�v�`dGS�o��d��:����p�t�����4W��x��3�g�	�*w��.��w��5@x;��J��B�PR��������6� z�w�/��6&�`H�$��M��V��\�����}LZUQ��5QRQ��mB (��c���vf�]G�x0�^��93g��G�w6h5zH�����Q���(l�P���U�\!F�hîg1���C2H����9���r�ԤR���9:���V-|��⅋��d���0�4�\�">�|��S�t�yP���e�y�#��|.��H8&Y���&�d�yZ4OT������CC��!�X&���C�GR8��ǧ���ژȌ�T�`����J��h�x�c�ԚX)o��:X�`��<�΋�P�d&�>�t0��i������I��'�-e��-�{���0s8\~RE�y
c܀Vw��>�;z�L��9d\�&={&+�=.�q�afz�kτ��h�{���$B�5jD)4f��cf\9�=��7?Õ�Ej1q������!&�򅱘���n`.�(�0_����\_X�_}I(��F��1��]���Y����f�Q7۳`Fṹi���!]�(l@؀k�RQPle�9nޚF,�[�9l�x�o����fs�����b�T�( 	�1�JZ�Mc>����v~�����N�[�[��-i��7�GU���'^��Q'��)Y���.m�)��+5D��T��%u��~Q�5B�0� ��#z+?��ɢl�z�>��A����vW��k��Ko�-aaj����"�8��������D��2Ow(m��Lbso]@GNL�4�q����T�t5
�����oiZi"�k{�A���I���/�4��O::9`2E�P�N� ��	>������O�	�}rL��a2{�at�<䇜]�7Q��ឈ�c��5��.��LP8���w�F�Ҕ�x���K�3I~j�������C����DP�z�lʀ{ӥ4���Eڽu�B�I�pL����C�^g��x,�:�M�-l���S�,�Bcn���f�b��E��qer�ȷ	��l��1��[%�A���+r���pGi�����AG:n��􋖠�D���r����#w�/�K��(�̽ʮ�3Nq#Y�{#���I�fG \(��W\BVh{H��iQ��W�P��{R�k�g2�)�q�64����.=�z�D`�	ߘA�ܕ��?E�eɏ:��|�^d��c
_5긿��/�U�V��&hxYX����-�������]5lFS������o7�*����f�W��FU�j,�A����q��r3���dk��E��S!H㾦l27�{G<�������OW�HA
Y��ː=�
[xXT�X��Ww`��ѫ�҉M[�&��T**7�"�d�?慩HN���"Bo�ID�͒�|s�>C�m���~��L�k+�����mT�I�L���>�"W�`q!���ivn�j���U�`�N��ͬ�F'�M���`3���Ͽ������D���&D��5?y?lcb2����.�E"6J�=�o���B�&wn�$��$~UCWy)ֱ2��)�_�K���-�8���2�I�UB��%˧��e�"����D��u��DQV��rT"�q
��n U��^�;|���!�a�LG�T�45aA���̠�"�W�Jy8l�gw	X�n���8��&a����_9�7��\f	�V���.�d<��G�2�����X~���ɹ��Tqm#���	Y`5�S�2��iZ�Cf���Kf�J�F�5������>�E^�.Q����7�q��|0�0}cJ�������������6�J����m�|��v�lX�x-$`���TJ(X��r�����Jq����S5�a�L+�`��J�m�	�33�q�#��z����iZ���G���\�    IEND�B`�PK
     mdZ3��C� � /   images/cff7cff8-0125-49f3-ae91-9e6ccc0a4cc7.png�PNG

   IHDR  R  ~   �,  0�iCCPICC Profile  x��||eE���6�ѫt�q�"�����ٰD�ݐd�b	!��l#[`a�.  m�"M�(E�HS�. � MP����ܙ;�w�������w��L;s���;�%ɾc�,�3��$s�-�<��Ǟ{UWz%���K6Jt���-]]	~���{,i��G�i����g����a~���a����_:`���'�}�s��Dc���!z��G��xrzS����
:�jKf����d�:�Ë&ɪ]�i�=<�2���м����3�Θ�$�A"ɬ9���>�Ɯ;����I2��E�ó�dm����}F�5k���6)�L\R��~��.Ӻ���nU�2֜�ff����[��78<4�M�$%Ӵ)KӁsY���L�M�M=Mف����n�ٻG�e�'+�iIW��d��-��N�˒f�J���֎�5��׭�Y�`2���P2�l�4�]�3�M�^�����gI�Ԯ�� T'~{\ˁs1�Y�ѶE{oR,���g�����u����C�f/��@����jM$=	�Bos��;}l���-!����b�$I�`�!������d��c��$k��$��@�y�S��������������)�9�%ɵ�m�ɓɫ��6l� vmاaY���6<��ڨ5Fe���:d�e��]����G_<��1��sژ'�n6v��+��s�wĸV�x�y+�v�MV^��C�LX�;�<Va�+�:c�?�ֹ�]���~�z����rͳ�Zk��������:����i�m����w����~a�/\�aۆ�耍����M��ț�n6c�7p�c��_L�x[�_j����O8cˁ���국��f�/o�����iv��k�}�/��u�|~�8X�Q{���Nݮ�ӷ��C;���_;�岉��>:�;�<y�]���~���t����ԍ�Zw[�}i����O���5{��k�7���ߞ�w��o���)3���f>��}���y��_����^�xs�p���]v�w�:����>��#78���s���vܣ'�w⸓.8����O;��	g����g�t�%�u���Oν���]���W^~�{������|r�S�����r�W�ܺ�����o��󮻮����N|��<<���?^���lz��g|n�秼8��^���]_�ፉo���x�����^�тO��_�?����ڕ\�|���pݨG6��3p�{�ye�A��w�J3W����*7W�^���[��5�Ys�Z�}�:����z^��>�p��&l��&{l�x�S7���W_nL���MZ���լ��ns���������=���7�x�XY���כ�-l�v[5�~�vޱ{����������^8麶;w~l�K������n�!;w�2w�q]��vo�+�+O�j�.����=��/���7_�֊���޺�}��͘3�p���3����{�~WϹ}�C���O�W]�ɢ���/����Z���c>c�%߹��������#�Q����ѳ�Y|�����q?<��.��U'^{�/N����N�|�����?9��3�8�Գ~�c�>�C�=��_��?�`���h�O�^<��/�x�֗�}E�\��U�|�Օkֽv������冎w����C7/�ղ[�����κ��;����~s�o���߽|�w�{���������~�؃?t��w���G��g���������'>�������̎��n������^���F�<�o+�����������vx}�o.}��^����<��'�����>��Ã����n���c��_���a��Fm:�Q���Yc�{����ݱ҂��]����U�d��V;~���8u��ֺb�׹g���{q���0z��7�z�6�}��7;a�K�������Ҹ�Mh�r���n��6�|�'7����[�ro�x�{��-���JfU��v|u���A�زӔ�}�e��C[O���kv���Gwy���]+_���ީ�N���{^�6f���'�����W~����ӷ��{l�&�dm3�����x��C��{�~�Ϲ{�S�^_����٢�Ż/�}�A�����:��e���{�*�m~8;���ݏ����>�S�=���w��p�9�铞;��S^:��察���>��3�;���>�чgp��~x�G���@�%}���.��%���ν��+��򰫎��q??��3����+���w\�����M�����o�ආ�+w����~��o�;w�]�]�w��Y�ιo���>0�����!��c9�ѓ�x�c�?������'yj��s����������em|~�ƾ����x�ٗ��ݯ������?.{���/~�7�x�ތ��ݿ��ƿV|�����m>��x�'�$:�%�5Lj8���Q{��{�}��1?��7��m��+����U6Z����V�r��V?s���<�K׾v��ֽ�����+�_�x�&6]��M�?S�ŭw����O8g��zh뗷�x����m�X��+��˲�ٙ�"q��Uݣ5�ؿm���cvXw�	;�u�̘����I���z�?M~�}��7��t�޹tʏ����\��	���L?b���͞��⛛|K~{J߬��?}�+n����3�����7�>�o�9��m��������?|���.^��%���_?(9x�e㿣���C�]r�I�_r��G>~�kG7�ޱ�/�k9��=~0p�ܓ�|�)�N���CO;�G�~�ǜy�Y��踳O<�sO?����~r��_x�E����G.��e?���+����ّ??���9�ڳ���/.���n��������7��WO��̭�����o���?�͊;G�n�]��W�g�{W�o�}�����������w<rˣ7���]���O\���<���O�磟9�/�?{�s�����x�{/��i/���K_���;���?����o���Vo���޷�}��w��w�n|������~壷>��'� rX8��< �8!I&�+�jŊ��N��]e��X��I�J�s�I�����I2�KI"�a��g�ly0�j9.͹�g�G��1����Ã���צ�L?h�C'�Y<���Z�ޕv�8IF`��'�utT=`M�?���iI2p�{�14��V��@���u�5x� ��������������v`�dc����ߍW��U!pS�0�0{��_�+p|zT/^'����gԅx����xm��7z{�~o�~��ܿ�~��W�zF?�W�3&w�ok��9�v2�@���z�3��i/VJ������hq�>�[�P�Bp�OH%8�����/���� \�������p�e
Ҝ.p�j���|��n]	��Š�o��?If�����W[2%iǘ���|�|�En����&��[S�p,D�2�:�L8�=Ȁ�Au��z�c8���!O��e���7�} �s�;�5-�:��g��?�?�2�\�M#V���+i��A��"N��tm�Aw���$%30����@f$#:W������S�7i�D�� ����?�!� s?�4�@;��J�8�-��SX����e��|�I|�?o:��1� $�)sd���2���K���gA�qs������l��g��A�s�"��m��j�R��������;����2<k�9���9C��/�?���?<kpQu`v���м����������ۧ���:ch�������޶I�ƞ�E����Uf���N��$sՁFL=�����������8�����e��JO���m}��;�zzۺ�'��vv�M�n۳h� ��:z��;�v�u�uU�'O�n���tOn��k����=��mJo�q���E�ա�:	K�ӿ�kx~S�u���Ý���7���|]}�{v�aܝ��zv�6N����Ll�i�k�~��J�(�[OW[kowKGޭcZ'�6;���Z'u�j�5�eƤUkk�k��j��Z��e��2ejwgKG�^m��z���ٗ�i�q϶�����ImS�:�����abwKo��)}]S{z�'v�y���6�TİgGGD��=ugz�Si^Rm�v�����܊ί��D�ڊ�\48�z�Т�A"���k�fk��?oF5?��Ξ*�e5�Xm��a�����)�J�L����=���Y���H�A�;ZZw��!?:��)=nW~3��sw7d�������.�8�����3��z �jc3���s���]F0u������Ӷ۴6K�qjWo{'���	c���S�4�T�2eZ�Ķ�>ld����I=U�E<����og:��JOKgW�S
��n��d���I������������#��i��fZ����A?�c��V�2���'[�F�
+a�ҽ�U�jt�W���^U�ƅIU�����~�������8���R-2�YiҊ�����~�f��k�q����O�����2��~�	f��ʚf�[�O0�
Q1Qz��8(���8:���'%�JM��=����&2�9�Ei)h�V)�T���c�e�k<�R��<2Z�Hוl�����AGͳ*�]��(4�M%�2����*�)�s]iMs�Y4�q����u�r+5�`�Iiy5n�E�م�Y-�)�@g�٪�%�#�%�_������Ό��Ԡ<F�J�J��X�05e��T�B�)����U%�%�1rנ�*Nf$3T/�i%C8ľS�v�Y��̬#�J�F�-6bY�܎>K�MX�6�1�HJ�H�U��&�2l�p�4[��M-5�$*���NA�� �Ժ#��e�F���ƪ�fRn����I�2G.�R�H��
<P�C�G%�Lf��5!�$��j�x�י��5��56��@���0�)l�8�z�k��~��R�Sk+p
��Q�:��Ƥ�ր�{� ��)�T�[��^G0��$��e�TY�#f��p0ZV��dXOp�T�9��@H7�R)�F+s�u���I)@�����r�
$�tMH:�z��mKx��ž�K@�p�D�G�%���ʩ�%]C��T�
ǲ�Gs�Q6+SN�����~*���L���p�8w�9iwRA#�5f��	%�AX���K�uRKK�uk3if=�Fa���K��*\U��y��#2���"�'����&�q4�xMl�i���'~D�T���@+G�$ͬ'������ ���B�%�ZU8|,ܣ%ͬ'�/����;�m��>�"���N���a�dA�t����,U�YUX�ι�:�^��#��0�	`��FA�֕�0�j�:~(+L	��CU�q	Q��u�Dq,����p���?CGQ�h������?�>�����=PH�?C�_�?�*L���ʩE��;�:��*J���+58��Iޖ��	�LC�d/n6�FC��� \��_1�?�$U��N)"�(�4����@���#&��I]�)U�6�2�)p
P{سդ�������z��� ��
�C����{*qR�JM1�T�� �42�U�hB�TJ*t��b5,���h;0�\��Z�F���*p�Z�!�:�t�jx		,��a�`�FT`)��| �#$9bFhf���Q�ë�R��%ͬ'$ia9Eq˒$�TFp\W��a�_G�,Q��$�#�Ru怈�HS5�@)���76�R�Zҹ 2�,�R:J����4��pE���$"��(���p�_G���r��>��P����j�PX��zB�n�w��0#�8y���(�؎$�'�0��C
cB�"�R�iA3R�z�0	�o� $CZ�f̠�p�v�u�!p}�5�#݃[� �Z(|���	x�a�����G��j ,*J�d1����%!�B,a9�8�]E钬!Be��'&���2� h�LI�gD`E��Q����.8 9�([����
�Ԡ�O"e*O%� ��d:EG��e:PFX�i�s�a
���X!�F$�.}0�P�9e,��c}G�U!(kd�FƁ�C&������ܭ�#�i��)�%�j���QĎ��8 ��A�=9X�/ WS���wD<Eg9X�?	��=�ȭ�;

� ,���{���P �K��x�@*�@� Dq��<+֋l�>Y�R�g�C���	r�W �b���A`��SN���D૘+��()���@�vd)*�������� ��)���BN<YuT�Рd�Ry��Dq�jd8��)2��(J9��*3*�0#I�p�BW�,�(���)�T�j2�3G�tQ ��W��(�G,U��bV!����?C �A"�/�-wE�k�b��d�qF p�d�>0� 5����%�*V(��F�RR�wK�;�O��g� "wnX4�T��R��1+���[0��+#sQ��+p���W�@(�"ׁsd��Y�G&+��x�(@ #C^N³!X��
�W��3"��yXE�3tP��U��)����������TE���U%�R)�g�	�����
�е��=�T ,�ܣL��(��q��5 aԹGC�F���pl�{,:
�r�F�s:P�I�-�J������Pmi8a8��Sa���f%=�bIU��gR���TH�>����mZ�6��"���'��DO^�[���"�g�[����� ��(q�Q�3
v�%��(��:��eU�b`���� 	E>��C��YVG.z"�d 䒪3���u�3����w�(���Ѯ~(]-����YVK.zr��T�#+�����jmy�񫥴�CH)ὔs͚`z%+-'�@��`(�%���%�	;��e��ؓ���M�@�=m��=Y�(4�� �1�p�䝡�����KL$J�����մ(u^2@��)�T���2r`K���fN�3.d;��\�I:~$=��@�{�~��*�5z��t�S�V��9�jڧ.q�q���s��"�	U6��eSY���}�eS��)�f�)0�iKzFϔR�I �`��J�+S���@ rZ6�D�ŠU~8��L#��� -���/!o�ی��-[Pi�ϴq��2�Ig��D\���j�yY��y ���%=#A���i��Ǩ"CePڧ,�q�������T3��%
�SOU�5�& ����kAu*�Жt���U���dÆd��	dwH�H��Z=�Z�QIy*�Q0�&+���%^3���q�yBR��w*qpNz�KӘ��`S���K2��Pt��A�����OQ�_S�q�z�(iNV�M�$&H	��1
WlDO	� ��L�Qqr�Ty
��H���cJ��D�7��(�J�¸K�0�0�
=Ed�?'���4��\������`t�L%(9�qZ˭��P�3���� �!����U�'�g��g��=�}�f�P���L�H�EO[�f�����J�r���0�(sy�@���Y�t<�aj�9EV�

M��)���r=YfiNF�G�A�c��KI���I����U�HV��q�Tw�u�J'WyOn4��(K�cOzPĀ%H��H�)a��\�,���B֨W��j��J
o���Y���+�g�łzl��i�S�`���p�����e��}Ҝ��g�'��	�h
���.
�V�;r�p�6��fȊ���,3��	�
���~��C����2+�QT��/zR%�S>'Ҹ~H�����V ��* ����J	�J^�o�O���(��;�×t�R��ۢ'E�T@[2*S�(�I�"�0���#f�̸���P>MZ=DOU�3n�����:=Z�甔��2?�Isfy��V���<�8z�{R�R����K�?�ׄ��ZP}Or 1:F��q�TR��cq����A*0��W�e`��SGeR5��%�z䚹�^=�.iĞP�Y�F��SN�9�O�}~ڛ }̃7K]D�H}��J���(!��P�	 ń�"]D"l�dIt��Đg�(Rq�Q\d�V�ʒ�BfX[
���1����)\�t�����vȅQ.H�o�,�Ӕ��� ���'J�����)[�
MȨX.�#(�ڼgF�L�9�x��=�|�t=��BBz�������&�bR���a��F��q��PyM
�i��!�	I��F����pʤ���<O=	�iQr�q�����N(���)�)���Y&�
27�dqѮB7?���%C���
۳����ڭ�O�[��Mb�rÕMVm�n�y��Ӽ��c�y�u�yfF�~�mD�Ȫ��]:���EP� ���!������&z�Dw�4E�j�������.�=�o���Cs��1���s�.l�6��3�r�VYrIR�\�����$��uH����!��-�G:^�g\DR���ݓWJ:^M7��+i�Ƚ礥��@�x���8�Z�*����ע��b6�K��缔���$2c�tňx��G{�UѩOZ�	��2�-����Ll�HCT�=�����jEh1:��N�|T��2�EhE`t��������9�@��9^ZB��rFO�s[�/�uG��J@�@��Μ��;��?1��N=���%u��RbǫSzt�Zm�]x+��At����n��A� �����,�W�7;���D�I��'qX��E��}+��n
�:W#�V�zU~��x��|H�HԎ�~rAѵM/�@��٬���Đo�n�1�I�9?��x^�$�Z�6�df�r��B�疛�k�I�
z��0������9�L�d<�D��Gb�\�	"o58='��|7�e���,#_$] �����ߦ�3"�d�9��7$��V�$�~�5Г%��*52�Y�u�6�p����,_B� ���U�nЄn��x�Q䭈�~��":Jߍ*z9�SIתa�<�$��|~!��f�i�Pf<)����s��]�kuY�$N%t�����Bb�0y�I-�9�)�r^�?^�V���Ҧ*��X.3�^��`��ZA�����r�_�s��z�Z��yu~������a�s]�ru��_A�xA7a�v�㕩7H�D~�#'�)4]��ym�g��iH�Ck��Y�n2o��o��S(RɜW��H|84�TOB�r��(Z�V#�
$g~�ty]z^�_�r��MV� 	�)��&�F�DM�9'�nN�y�5�\!�N�<
��<	��K* 3HV&��|Λ�f�ji	��6���r�Z%z�@ʠ%�J���7����I
���`o�\+�_�� �K����V1(�w��/�$�c��"ZAx�J2+F��+ϋ�٠.ጵ��S9�k=/9k�j�)�u� (�t�d^��N&2?B�+���
}��a��;F:Mu���v�c�tN�:��PQ&���E� �˱��@������q/�\x���>P+saϓ�z�D��܏�è�U3��PH��IN�]�[\�g��=L��K�)q��0�g�,�"��|	�X�j��_I����\�X�\+�i�z�5{O 2�^�"��­	�2V��~��� �e�_:�˯��7�y�,d�ݵ��D��e�C���r�*@�6tC����C9�*0DAfE�������'����ޠ�{2]|��I�HH��
�L���{��/�� p Y�ܤ�j�N!�d�y��t��n2��0L���u [ɘ�![|΂yO����������0Z"���D��x��0�W��đ����0p�և[�ڛ4'o�<bfl���OhE��yC�@��Z�'��1�GC�8
��{.FW��-0�7�HN�7��Uy_�#��Ⱦ�C:������EuӬ yȬ8��a8D�'��&�V�}��d�0}7�9��1�#	���p~ǰ�=o�a�՟0���1CF��/���{�2{�~܈ahZ�Ρ�2�Z��1��7&�T|���6�WO��er�Y<���_ʲ0��>BrJB��"��xx���ӄ���[`(��a
S!i���+)��H�׳�a���%G���$6ă�D�)Y�D��8A�q#��p�ޭ�L�ԑ���[`��F�{؁��WD�i$�QyI�g�y��g>nR&�]7�����Na96+��n=o�0X:��v�]<� 恷�0Xm�r��y3�yC��T�%|�IY�1t�� �t�6�,b��=�a��>��F�\[�#$��I��ﱧ�BR�UP���h���-0��2��T��c1��[r�S�1kU1�i��R��I���1}އ$��U�5���ɽS �¹�"�z#����,���eIoC"b����Z:pR���E#$���J��] x�*"��y=�T������[`,'�E�	gA7e3�[`,�ER#汧�F�'D �O�;�֟E�0��4��U����ED�� w�n\i)�-0]m�NL�B��)��F��X��_*��AF#�_xCY�&z��-0�>�f�e����GɈa����̼��TH��AF��2���T�j_ޗȈa$2'�}���|��g2b$����&�t����0HWT*�$���1��a\��x�g�"#������0U���x��H�UэPYNbX��2b�n�R�Rg���0�"������K
�y�)�O�%9J����YDC�\�NC7�9D#	q�@j���F��
�xT��XЇ�a��yX$\E8!����1"w�- m�:�ce1��Oɛ@Zx�9��FRu1LL���I�fàՆq�����~܈a�¸D���G����d�0hաbZ�:ݤ�k��R�nP�2�𵷋�a0��A Ï(�㐊FR���`��i�3�[`��S���5ؼJ�x����JB��`��U�0��/sOʀ�1�J��-0ZC�H���С�i=o�a��m`���%�>��������-�'��W�u(�[`�����w�i�k
*bŘ�ABk��MK_�P�(�Wo�
*�}*=��511}ZW�����*b�L�+�����n��T�0���+}���	0��uZ1�E�U�;���>`�y�(�{�!z݁��>�Q�(�[�ިXx����1���?�ʐK��k�y�`AA� |�Qt���Y�0��3�a�*t=bEwȳ� |ȧ:��Q�F�9}(�=F�1�k}~���xo�ȭx�F�3�!X��Ǫ�a�e!��A�@�P�V� �����҆ڕ��ޗ�A�p��V|mEG�+}D媠}p+��a���ح�礦˙��FY�@א��R��ۦ���D�=�?71��k�{���)�C�atV$m��R+��:b
�,�&�&���ǩ:bڭwx��T���WG�黩�s�9i����a�d�^B^�C�<>��h�SAPT��"���k�x���`��l��?�À�{��X�Ky݉F#��O�#���5D�"|2K�T 9=�p��`
�Y<��O�Hn�`
��%@g��@執�a0��nE+���Iz^��FCS���B�J��a�
5��M~M��sވa0E𓚤Zu�Y:bLa}�Hw��,��5DC_�ࡄ�¹�}~�#�q�گ�(N����y7T3<���lz�c"���)'?�:���8d"�A�

Co�2C�R¸�Ak�{����5�bW�G��5T$	�E]��-�뺉�Z�Ã��89o�a���!�׀��͛�a�5���-OZ���Z=ޡ'����%��1�� a�n����/��a{5�C��X@Z_G4��W���W0o"���~oàU�:�!�/H�k�&bËg�=4T������pև(�:i"�!��^ʇ�� �L�0`Pa�z� ^7à5�>�X�¸:�L�0��Z�;��ri��Ɛ����4�<7À�P�pB*?,�[`����-��GHz��kL&b��3���6X<��g&b�{Á��C��x�D�PP!'�q5�k�&b0dv�CӰc��#�1�e� ��]<\��+11��Z!���b#o�a� ���z�J2��[`C�)�Y��z��o�0�M�c f�&�k��+ۈa,}Q^�fC}�����1P�!��.Z��f=o�a�V�<�����]�����{Ɲ3�!7����E1��a�p��`0�c�����Bɹ��l�0"!B
̛��/����0����o����(��2�����xa	��q��_o�0��*�W�����<o�a,U�Āj^�ع�b#���)��R�y%���җn�7@��Oڈa0��
2@*��5R1��uK��wA��<o�a�G%����K�d��-b�3��ᰃ�4�x�-0����n:⃔<&���%�;pt�͇qrPao�XCߐ�I�t֕�r��Xz�x���[��Iϲ��w�Z,]��֥��Rw�$�_�Q���d   	pHYs  %  %IR$�   �eXIfII*     (           >       F   i�    N       %     %      �    R  �    ~  ��    x       ASCII   Screenshot�lK  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:exif="http://ns.adobe.com/exif/1.0/">
         <exif:PixelYDimension>1662</exif:PixelYDimension>
         <exif:PixelXDimension>338</exif:PixelXDimension>
         <exif:UserComment>Screenshot</exif:UserComment>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
���%  ��IDATx����b+Kn$����r���f�����f�i�m��,�(���@ �)��3�ͦ�D��2#�@ h�駹,�y���Ҷ��N�T��/�0���Q^���g]���yL�O���g��>�~��?_z����~��{�z�=�vl���/����>&��]����c�g��K��>��)8�+��ֵ���?ȱ8�y�����t]��+o^녟����k@�;=�<�{UV���Q~�Uf�)�;���������b��8w1浭��k�\������1��F�n��ֳ�ɦI�D/��+��4�a��M����M�,��g꺱��up|�5~�{�9��ƞ������>.k�k�;/�x�n�-ϝ�<��a�	��z./�I���k������^>�/�k'��/��<!.0��%`�.8��|�ȟ]�g)/���V }�m\�W^����<���B�nB�
���(�~˵�X�\�i�r��m�g{�׮�*�n��"Hl�s�z���-� Pci�3�$���P��j�Y������`��Y�� �uRl��
��s^���k[}����4�5��s^���|H�����Y��=��'?7{���WS���1��%��ǩ��nD�{��n�=ޫ�x��!��s�����L{yPy����ܗ�lUf��q@[v�i�޴*��S�vv8�oi��_�j��K ß����(����d�~˹��(�z��1�d˖�k��h�5?����//h�����! �8����R�;���ႁR�K� ?������G
58m��B�Z��n�<�	���j��MWe�8�U)�R��4,L��?��)��)����T��� N�$��(���ܸ��
���p����}�����s�+����m#���i�Z8[���D�lw������{ �ֲ����"'@^[d�,�#���^;޷��k�{���k�/���6�y�<.�ւ�З�g{��w�{C|&���u��o��ۿ���?������o|ӞgS3H����c�'��� �`F���Y7&|��X��
H7�NVo�q~��<[ V�Tޜ,��z�d85_߹�r�s/�c��1	��^u�Y��έ�iD5~|������aT+y��O�ʺ���f�ǹh��GL�Ȧ�2�j��\^ݨ�����|۵���i���T��=�k�齯��kǺd�_�K���l7��wm-�kV������6�|���]������w�����8��rk�-0�vn�sE[S�ப�V�b\-��z��߬�K�Z��>�=j=�����_�O�Q�����p��{yi#�s�����5��%���r�Sv�l��i�s���n���X�u����j�v�a���	Hi�ft��K q�Z�7%>�X��ސ��e��}\������?_z���fs�����=�@4.s�y�f�����js�ڶ�o������Эq�;�kc~�ҹ��o���S��֓p{+�.[�d[�������,�:,Q���9ߗ �K`�?%9=��6m�eե���[���2��XK�{N�w	L�g�ݗ�+(��qG�� �k�*�V�z}�k_�Z��Ā����D�@ʓ"�:�����۽�1�����*͏k`�?�__{ϥ_��㵽�;��ݯ=�Yp2��+V������U��k鋅��V������g��va_s���[���}�r���}S �_Ӽ�0s�>����`�ãi�E[5@ҕU��LJ�!��9^WWB,؊!�J��$�t\��	�?��.�g�_j�����Vhy����w�z�cE�����ϥ�9N5�.���Zq\~�	ەh�r<�N���<??�?������j�� ��Y�����_]x�I�M���Z�[�Nke9]�ޮ����]�?�o�&9�,�8�8��{/}�{�_�}�Vvv��h��r׬.\>�}k!^;��{��9,@*`*^SD�4P��"Ȗ���z��=��ɭ��&��ʏY� j`����Z�[�����P���p��5���⸎��7�n����Rz]�ȑ()9T}q�/?�ŵM�T��۵�aU�Vr�ĭ���o�z�~H�<�	,�e��+@���ɟ��ׯ�Ŀ�z#z7��U�eS>,sp�[��53>_߻5���o�����߽���O����um���)7�-E���^s��0�f�^�k\[>��Z�Ǿt< �C����kns�3S���]�K_h�o�Q� bx`�������
8���K�~e����k���������3�%���#t�M��ſ����Ks0oa�V0��B3
 ������?|/���hQ|�߾�ͫ�h\�5���M��M�$-O�(�_�|)����<��wy��ϟ?�u����o�1�y�d�f{[ �fM��[^7/���������-��g����}�s�&l������|	���T����9]Q��D%]�����߷�l�� U�iT��`�}�/��z�ƾ�t���J~��wN���[��Lpk�*p���פOЅR� o��c�y.�7�YH��+�R�V��D�=��:���� 8��������[����������bm�������f�P�������{&����i��N���@1���|������O�������/����xL���% �����e����v�̟�<�/��[�,�j}~�g.�|�k���5k��ud�k�.�5������\�k�5�c���cѵ��5�f���Tt�/9�)}��
��k}������I���3(��j<m#H(r�Z��h�E:��� +�\W�A28��]���փ�Au����9�6����[�
��������A@���S9,�#����l�jL߻��6�µ�7�W��'L�.;\wX��<� 
`�k����(�v�ǀ�[`�.���|�^r3.Y�|�%���?�|�f�~˱��sڂҵ�o��K����K����t�����k�@�;[K��wl5�[�즶l"��,hM�8�9Rr��A�O��r���c�f�͓Y]�����9 �C���[. �KPŵ�v��7��V� �H�8��0���1���XO���vӸ���Y���Ҹĸ`�������lN?~��\��sMA}����X?,�mr�����=$x��Iw��' V(�F %��g^(/&�y������3@�w��@���U��G����k��%0�f�^����~.�k����/�_�^�����2���ZxϷA�Ks�7�ɬ�������۱��K�!;���1�L�4�8�2�b]?�%0EVT���V�1S�U�i,���(�L5G^%jIgQ�֖}���΁����<W��(O� S���\�E���>N���_�"�����W-�YzNr}�l�%uu�E�oR� r�t��{��xps�h��.X�E]r��m���3~�[�@���\��luw�k����ϳ�a[+����e����.Y��6�Kחݳ��l��K�|�\��˟����f�G�:�Ų-�Cω��I���E��<�܀^�����q�	Ƹw�.��s�k JnځT�$���V�<�H3-�� ;��W�w�1QtH��Z�d����F@
�	��p���*��_�B����Q�����v��`��	���^�e{�(,�X�kq�\Z#�<��i��Vf��&���Z0�I. ���������w�iN�j!x1h��H�AVYH�5�E�W!ݴ1�y4�^}�U��)"����rIULT'�� �9i+�]-�q���Ť��}��|��)i��-������@�q��Q�"���@I���>��ܶ��������ww�]�A^"c6�[�q�����"���:��"o܌�F�ە5��3����'rs�3�<��%���(�n�%�F]�xv]XB�-���� �tVeV+�9��t�_ɽ.UTh��'���yۦ�u1����Q��K��R4��߻�b>v��J�s��R9`QzTl#�Q�}�s�d>��+׬Z�h�~�]O���HYxD�⨹���0�vlU)�q}W�[�ꅠj�s��r.S���㳸��>�ݻ����$� V���-��$�;�QO'n{6ĵOT�]3D�,����iA�_����?���_��%2R)��^�L�����տsʕ�P��/^�t��I���r�粓ส8�g͚��D��A`o	>Zk���B%�3G�H�����xE$.�m\,����q2�.���;�Z|X�zUD6�:�:�����\^�@��S�}/;/������tNހ.�t�G\�|�`��r���r�q����=Z�L���x��2,ݻUw6�1�]��l�J�4q&�%DW��@�/7鵋��%F���B�a�X4���{Q�h�6_p�8�����=�\����3q�x�"=с��5�+xb�XH�gb��J4������&��f@������9�x-�_ �����'z�Ј��p�;1d��s���/<q휏s�N<��l��x��������������OY�쨁Ù�����7�r4
�՟̒�*�֪]�cȾd@�	�믿���������?�ub�,`a04��ˢu�{^�"��dd�_&[?�F��P��@�������V|=,��U���t�67��|��y�Eۗ�2��ʀsX�mc;�����gV��1&&wV��cnn���]������J�����p����\�h�X�&��.����bjOgD&o����r^8���Q@��'ۜ��agr��r\��g�P�ƣ���SY�B��p+����mX5��,��QT����y(��Ţ˙sZ�M%,��\�ae��Ƚ:��D�X�@��u�ߍW������
u�U����\��w�H�7-&��������Եt�k�b#S���5��#�)�4ʆEQ���(*B�����ƌ�ȓW���o<�5�������h��6q�
�
��F�2.�����'�F9����
N���{��y�0?���8��~o��A�Ԯ�V3�k�|���N��_�o�k8 �+����H��E:{=l(��)�� �H.�T�Z��A ��ڐ\ x��鯿�Z�d���.�!7S&=n�IM��tu>����d֠�v�q�`��ЬĐ��ݻ������?���u�1i�]'v��w��n�I ����K@�/׵���r�K>'�N8̱=���q}�D����r��)�NE&%\��[ )&�k-�EKւPm�ܲ��j=ʎ�'��\����T�`�y�����ή|��w�qM��NT���R�\�2隶�c�~<?�eAcǵ �︻�),��;��[���C�V�.tq\Xj1	O��H��Z��4 j.�i��ԂýQ<x9f�,�Zh��$D*��`��[�7�Oq�Zʹэ�	�?,dl0��5}�t�X3�6{ә�8�}�^��A
�XE��s�}�W��a�Yօ�����4W2Ns��}�!�A �[�Ê"8�U��w;y���{\�����9�fe Tc9)k<�6�c���e�vK4h����*�B��������������1�$�f�	zN���`��/�8�1��fhM�em�:==�el';�nj�<k�-6�v��*7\���' ���x����_@�m�5 ��?/�ݾ�	�Xz���2�9����Ų�vbk)�_IA�	����c�����0 ���Í�V&�y���E�3�(x*���\�-�p7����,��I.���ݸ�������r	d�zvz�.x�w��	��q�������]�ܟ�T�!u�.��t��sc̰h�Uf�HĶRwJt�8�Y>����y�Bw�y9�mo��.s���nnj����:X%s�0�]���F�C/��kx�t�ټ�'��~T��*�� �eRY�zϭ�W�{��4��{d_��{j
�1&������\��,�N��Y��܃e�/ks$s���z��4���� ���NU��G�	�t����|1�a����ʼ��}	>3|+��5fh���)�0�u��ū p�:��y\�r1ޚ/��*��Dj󎻾[6�[�4�����˸��&���.[�!�9i�+���7ޡ��>Λ@z&�~�,�������ٹ;l�.�|���I
Z��n7L..���ﰨ0��� �#��d|)^��;n ]*LG¹i��,�O �e2"�@�V3���l�o�-_�.���pN�Tª�
�T�����Od.��Y�j�+ ~]6'<�g�Q���_��X�ߗ�~E�د��u!������2x>�_����<?;�M�O-�
��/^ �Y�j��g��C8_|?����tX��YqP3J��8W���M�Z<�i0~\i	 ����<qH	���])�+[�'x6���GKQ��,�έ�v�W��R��)f=�}��bƼ�XBM}�J�:��;c�bQ�{���㒫��������X���|��B������&�� oB��s�w����ߋ���7�W7u���Ÿ�g ��`G�VL�e�T����ͪ��w�2H�vIj�����h-͋�1���.@{g�����)f���'�y�c�(Ć�sU֤]O��\�Jw������c�� �".�^n��;e�H�h�%u��0H�X���.��eq���-���?L<�@�w7�X�}�w�Ggّ73K؂(�5a�
w�E�+��d����.��k�b 7��������f�Ҭ�����(���f�H!4l_4ݪ0���p��Z��w���������o2qZ��1I�;��^8��U)��1�O�X��S�@1�!�%J��ˤÄS>\-/	&}��8��i��y���� VX܍�	�; އs�Jٰ����+?����+X���0/H�)�����W����{�y� �r�O��86��x����������<����\	�3fH�h�������|^Y� ܤ�(��ȇ��#��ViL`0O <}���픑m�/=@ ��oI��u�t���4������p�ܴ��R i�<�	�"�~XE�{:٘H[�"��tTSb��>W���Ov}��'Z��8u�Z�輺�?���J��-C��zh4a͐�ˢ�l�2'�f���D?�{���_S���$��w���VwQ��W%E �j�H�뱝ޅ�EwSXn��oL(��N&���4��l���jQ����yH
�� �ާJvsq�d�܈E2��]�'��؝l�0�p��ss?��t*!�k 5��1+B΄��8l��y��˧f� ƞ�w������P �Nґ��t�צ�h���PЍ�@똠{��7��M:��P�샎�͝���"R�ND$Q[s[=�t�Kc�, �QW?b#� �	��̡��ks��J���������X r�đD������V�S�餯M�@��2�m�K��z�R�Dc�6�D������D�ʊs �5��\<��븩wb�1��ʔ86O��-��w�۝ݍ��k�!��[!�y�@�Ojk5q��x ���U���Y�,\@����NoQ�������Q��Z�x�4w
��rW|�"�������"U�Ckx]�E� ����_�R>�~��@���(�0wZ��p~P�B�9�p�����?�M�HA-r�EQYvS���%��K�r^X�p�>��I�ߋ���I:$8&��fh�������&��^�9��WKe9�r�ɸ��� ��N�Q�*��5�a���ir��%�`L9Nuc���z��|j�=sqޝV�0�Mp���H�1��-�b7kʠϢ���Y�lŮ��&�N�,!\�Ԙ0kJ^��n�s���s��@�p}#z7*�!��W@j�'�Ż��&bR:��+7V���`� �2�b ��� p� ��R����\e��J�R�pKq�l¤�X� p�V�%�v��~ۤ����u�z>0T��`o<�h u���4���H�����eó]����A��ė�n�77E�[��l�٢�����q�w:���%.?aA�E�I�T4�J4�	|�#��6+��j�u� 1��]'\�G\�&�� ���Y8IR	ʙ��2 ��7}X\W�Q�����~L�]�a��G$�Tk`����hgsC�I����*�����{��r���e!VP-�Mڗ�Ȣ��y�I��E�� �y><(?��a��4�9�ɤ����M<4Тꁮ]��l�,� ��W����Veeҥɬ�N�Wr����e]��ﵕ2@G9���c�,�we����ǯ��È�9<9�A�-�&)׃~�<W"|��8x	�ڂ$ͨ���N`�;?('~R����o��:��jZ����ѧi�8P�#��g�;}	��Nܵ�C�_%�P����7i���k��=��\�5���Oi�5)H��g�����5jr���Xy��,�l�V>�z�:�2�h��B���f�7����Z�;���v�ɢ���EJ^�r�;#�%�4���g&��]�8X�@�4�K��3J��߼VZ���4I�~c�s���� ��]����ν�t�8(�bz6�J�gJ���ANº�>BS�6��dt�ܢ�~����g���4��$�d4��>�7��Xu%����<M��u�����vu�޲X�%o��ZW$a��X�hx���m�7>C�oZi�l(8�<�Ώ��,�#�nl8bɎ�G�u�v6����GS���r�B�D���+Ξ����u�(t�A��g�<����m����p�SA�Q�LK:W��%)1�j�{Hml��:�je�ǖY1�"}����ϕ��=�W���u�q�5"w@Ć'�lq�������r�Gq�(�厫)��v8h:'O�|�=̚�����ãg#�f��%&�,��)R�XuG���s�ӈI��8Bja=�ƀ����>�DA�G�9�S!]bn~%�3�טe;�({�E{6KB9���D��e��� � �����Ь"U��U�����&���h�Hnj�,��63+؛��(]�n��F����>XY��,��`)ugy��V�����5�4��yn�腄��C�D��4�Y1��3N.��$P��k�ܯ�=X�'w���u��믿-��,���1"��U�a<�s6�X��{��� #�2 m�����Y����p^�� 7
�s���x|f�0S�*�nE�)��poSp��*7{��y���{�(9�9��֍S���h�u�p=�-2,�T3�|��W�)Ċ�f�Lĺ?{���ʴ����;�M����&y*���#���EJ0}#j�rP��/��E&ԕ���s��Ee)��f=..�ނK��� S�KD�6�1uy��}��ew]���&@�I�dL�[\��;�t%��I,5F�w��gia!Φ�"�"Év/��4��d��2^s��E �IWn�gW�ke�G�7)6�tA���Z������}����(�=��g#��L�o�{#V=lt�I@|�0�W>:8�
?�����bs.80Xb�E�u,)���ҹ��A��{s
�5^w����g�\��o|>0�R�����-WK�����RF�����{Cr��7t��.o�s핣5�^@ײ���������s�^��H��1D T�#2����i���G�}]�s��B8l��v���=׬�,*5��JhQ+A�Z���v>���j��4%��ܑ�c^��5 \��i,BO��+źtci��w��Bg�5�@�A��n��ViH��{�ʟ5�?V���X@��ʭ�j���b}q0}�"U�xp��w�Y,mT���(���WΛc�&��E:��"w��Y@ԄԚF��p*���T��2A�1 �U<,�2ɊEtլHD�L�T�s��'+%*X`��������H�ĸ�HI	��]F��F��V�2���`I����Y�Q-��@01q�,RKR1qݪ�8�4\B���3��RY�p����D��o(����΂߳-������΢���n2g�:)ťX�)�<؂�v8�BaU t��7�)�j�ߙT�\�2�R����?��P�v�@?K"�U0�ň��i���;���H{I�T�F�饸vl����;d<�77cX�C�s颟����W�d�$b����hWXM�����P�:���)�F�>�j���N�A������3��h������z[ߐB�kB�3�S9�弻z5��G��'�c
dAUּ��0֞:��d&�nm��`2�u�tm��M�����7���|C&^gS�N����.�*������_?���V3o��o��T �D��CuTy���J�;���$�fՈKb�[�ƩК��s!�[dTS���x4�B'����h!��u!����K��+~G� d�$t����W+iΓ�	,sG�=E��T��VC�����g�	PGը�V�	�6��F���k�T����,,)�;�Ɠ�.Fd}��-F��XdC�J���R�=6�\�LK���Xq\�I�;C���E��z�M���g��v�`�Y2�&qh����j�����`��s@j��N��R*�u�NI��#��0J��V��7n�3Uz�l ��,�-ad������Vb�^e�W��mSWHH�A'�@�.0=�X$F���%QX�7��,.?Y��˭���4EJ��uT2�[\�r��7<2G���Ez	L]G���)\=�|	�t��b�Q�"KK�E��Rɓ�Q�!���E�o�trkV��a�ź,�nq���pm$U�`�MѸU�b ��Ȃ���H[*���!�q���"G�v��q/V�B ԕ�|'�,�K8����T�F�����������82����(�H��:0p��9�F�;<�1a��/��Z�`�z$9D^�2y���?	� ��F�Ct��]s9\�\���Wǆ��@��WV��v�B���Ϝ\�	��@$g�c��3��͛��T�v�sg�cP�E�=��<{K/1XUZ"n�+W�o;�!Q#g���*/��w���w,�䆍{�h�ws��\�D�l |�9X����1���XO�҈�M��97�т�b�@\�����h�'\dۄqg +X�4�ߎ�Ȣb��H��t���*�p���{4��V���ݔ�u��ؕ��e^!�l��KV��1�?��o(�,n��0�+�!��	�­�<��5�0x�L�^ ���}��u�7�������s�ZN�P��W�|�Ny
�a)��u҉X�@A�IGwe3Hc���\���,�M��f�9\�b��@�,���ieV��&f��r�9F7[P�rB-������W��|�ʻ�;�wf�<���r����.���ad>"���2�(��)M�8�Jk�剎�^N�iLo|��]�|�jY������\�4�0��4�Ҽ�^u�X49�7��������)�����fM��ߤ�TH7���h��Tk�=6�O=��Ѭؓ���=�N2�\��9���~���d�q0MY ����2y��B��lƣy6)�P����Ò$�B+��Xs��qTl��\��-GJ�"k��k��A(肷d�#{%t����{�#N����D
��kuR�à!��Q��Ē^�Js@���I������Ѓ��o+p�Bxp	U2�9I�*��e}`�a���R
xYt�TaM�X,�&?�v��12L	P�2��-]�:�QW�N=X�yN��WR�B�Yt����3�i�3�Xr���O9'�v�)G�׋d��Z��ӓ
/Ƣ����̽�H}�ua%�S��[���M eAV�R7y(ůW�?�hI��qZQ:��Y��`Jc%�%��@��݈��q�S-QKv��&����F��/�-�_[�杏/�W�~ P�����\��3�r���%;�[
�,���K l�C�u�i�b1gw�=[�>�{I�U\ŢT阧�I`ρg���Uҧ�P-6"���[]#Q�F���h`��1�RH�[��i���p��m�&� �3��<��{���:�u���<�+#<=�d���~ٵ_�O6Xu����lN�7լ����Eц�%C�v+�>8]�� $f�<�kf`��뗯�9F�]�ٶ �)%�
��U֊�u�n^G��J�U>�&�t$����N�>���8cӤ�!� c�͗A��GP�)[1�l1M�ù`q�w>)2���/,D�d>�$��jVR*L#��U$֤D��Ľ�h����^����wi�p�yNV�lE/z�=,>�G�Y	���|@c���be=y��3��{\/�@j�&��l��>R�Qi�t`����l!�)rO�{�fM��3�MJ	"�Q��m�iu�3����5hG�ȍj��J��w���-竅N膻++�r�EPh��C�`̯�A�Μ�`R6S�U,A�Ӻ��������
ߘR��u���)m�e��K�u��Tk��������v��^��d�Egu���r��g�1Z|��-l�W��Mמ(Xj��쓆@jBw�529NP��5���u(��M�b'ǂg��87t�1PR@bpb��+���=V��o�0�Vid��pcΟ�,@�,��dգ�:D��\�]�.Ό��k�{g��8v���1��d�E�e!-�딲U�2�H����'Y��~PW�$ORXD���� �[Oo�9��]��6�k��q�|�&�ʹ�4Zh��0o�	u���(0��)o���u��;6Nl�qM���� @o�l�p�nM�U.�@��1Ƈa�Q����Qa}��[��e�H���y#c�>xU�W8wՌ>ʆF��vjQa��z=�\�['d���jU����$t˜[*үM��)�ԅf>����cLG-�"��Nl�7M�T��s��^z��I�N����aD�u�InJ�d�<.+{�n����ϊI���d��ΛrW��e%�z����8��A�z�ld�H��N�:�6"��8[a�~�1K�k��h����U~��]W=
��!���]��wM�S'Wg�`�9u���z�(�h��^um��8gr~¶ksT,�k.�˷�h��;���i��*7��c�B]�H�+V������do�z)`k�uUu�1� �� �ǣ�8�Jj���"
��x�.�)�A�J��<�Kmջ��?�Y�CZy�< �?� �B����	�zGL�z��廏ߋ����</�S1`�nS�o&Q�1_;M�|R��5fa!Dq�,JN��<y��}�(�w�ڒ�� C����|�.k���cI@z0Z��Q^k�3�$�ۃ��a6y7u�%��4�FU��,�X�A���"�4C*��+W�T�v%�,RD�ihy�H~�z��Z������r�L�	
��U�ȸι_�`�Hg�71��zQG��~5�ֻ����8^D]7.�e��јt�[�.� �'.�I�-���{���:����6.Ց� bGС6m��b-g��)���ּl��PLN����b�ձ�����=���E�^FUE'��l-Oȥ��dO�擻kl`G+OK�=�UK��2zͥnl���4�����h��ڂۉM��A�� 0)����`���Ǧ[E���q%n�zL 6h�s��G�\:��;1���3���𜬯 T�<[:S �|Z+l�!�c7�S��hp�qa�EZ�
ƵG�w{&�d��C�ylNz'V5+E�j��pݣQM�)�qI`��1��#jo\*-��5� Qjk���i%#X�ˁQlL�9-��Ѳ���jG5ـ�h��$F��^��3�7*R��jgJ�� m���޺|̰`�8��dԉNv�0�v�e�?��� �,��}+#�+`����+�|��3���[�GѺ��/J@�&-L~K�QHY@E�"�D�.����e)3N��TR��,:���oZ�q8x�s�����I-��zq���4��uU����$y�*��-C�u+%�nk��d p��<�� 0k��cD?������H=X݁[[�fF~�Q ��9ϱhzM& hb`y�K�Y���+/Ӧr���Q�jj5.'����b�aQLN���,���lW�|:z�F"݁{�1
%���$�ι\ݤ"[k��&�Qm��hiC�0���$dHu�G��3M)+ҷ~�O�*�L�A+6�76�T�rȰ48vS�[�bxo���

��k���4%K�ܻ��͔�A�{��=^ǵ�������WY9H|v��=ߝک�"�~)֗5mU���oi�j����d|z� �ƃI�Kو���3zpNL�Y��q��Z��˒%�h���!\��5UO��]H5�;}��En̓e�0XE7��(����q����P)q:8��ߛ[�L����Y>9w(E������ߍ��)�	���P���dV-?�yb_l	�,�,vw�DkYw��R�2���Q�1'O2z��}��t�GK	�Vt6���F&�&V�;4�Y
N/@�q�~�J���-uQH���;<@�Q�x�����W�`���]������������1S��mL��HaT�ܺy�g�$��8F��AwS���0�J=�1��2uS������,X�n��V��ƀ����
��b�bĸ��ܨlɖ�[�9�Eԟ-0f����-/����<aHV�g����q�(��Z�Z����r��
L�.�*ӱ/aP/��Y|G�H��=�B*ы�B�D(58�=*�$y�0$�<��W݄w����G�E le�f�h��9vF���:5�%yb���&I��f�>�&�����R��n>�%��S7��AK�ꝵ+p�xN�o��c�N���k��XA8w����P[-yGk˅ģ�:�Jkͭ���Vm�B���g��7�l1�YE?y!�;N�$������cX\���ꏻeUp���k��A��� ��nR�{�4γ��6� �s��xc�U���y�X�s��j]�ʶ�u��A�k�4�9s�+Yފ�� |�q)M�ͪ�ַ��Df��Z����A}�b����c�ƆŢ+���f]��RF�J�,2��f�'��FY������l���Y�ō1$j��0Ƣb�����^RF:f�S���U�Z�h$1+�����̳d�5��8��Tۚ���VH��Q��-0 N��d�W�@qk+�/���0t6���� �\{J8L#�.��Z9$�彰T�O�r7�VM?��a������2kA��/J��J�Kv�s	��{KM��� �1�Ѣ���/���՝a�5ъ���X����;=�E�e����X�|�.��qZ��� i�d�3H�*g&n�l�뽽���Ƥ�5	��I�{��0
�Un��L(�? ���8GX����w�z� ԭ14�U��c��/���&<(j�Gԛ�F��ei����2�E�95�7�T]h�)=˜N�(�\��������:
��y\vև*m���}�0�D��2>��Z�{���v(�(�B��EjD�`4���~�����[��� i�31ù�q�B����N��7� �;K)�x�q]U���p�YmI�NZ0�����z� �~jBWT�˼lB� �����`��:����gԞ�Y=�3�|.${t�W<���+ �&��nQ��ݬ�6n�r��ɕ;�B�q ��	����C&Z��n7{��%Z���,��[6��ƪ��zDo�H<>}Vyʤ��rJ����}^����k~�O�/3�0W�y�k��	ԭ@��Z O�#o-$����1�;�;kJDV��X�+�DZl�C�Zڤ�e�"+��à�.�g԰
>+Qy�q#�����h����x<�z�t����T�T�� �D�����_ʓ��x?�4{1,���RWUH�,��VJ�'%>�7��;knҥW~�%�� �ȝ5sd���<mEì.���f�^dk�{a��{���;��"	cd�	��A6.�@��U�vο�c L��e� ]��b;��,�<���Q��NXJc��n�	�Z��d�vֱ�Fj�A�0K��:����jӞ[л*N����M��r]�K �� �y���f=5���װ�eY/�c�����k�6|�\�U9)�l)tQU&�)�KV�v
e��f���Y�r�K0�)�����Z�z�H����D�/�������4S�m I�x ا�Hy��
g��eAU�]Ŋ�R��@��w���K��VO�����9�k� )�SJ��Z�J"��Y�T�7&����Bp��E�gY3��tk�QX��ts%G�ւ-�ъ~,��_�_��/�?��?�/?�R���ߗ�֪���{F[��sDe'�����|�/_�3�j�Q̀S�i��G�g̀(5no�zƀ��)�Am�`J��`��q/03Mn�)�]���{&�Yu�Sa�I�j�"�lC�tV�[�]��9l�W��3i֝|'�+t,@��֊_���l�2ԊSy��McL^��S��<��Ϫ��(L��ܛ[O����h.aOT�m��"JRL����lY�B�9;�2}��D3��Y��g�B���'��XmaT�!K:�.�f�f�.��
�L.L��z�|��^���~K�K7� ���
?X�6�#��h�.�H�l�f��P#(n�Is�5	 �`��T�B�;˂'���'�,�n��̈;��i�I�`N�W���fϓV��� .�7(wi���Vζ�J7��.��9��N�L�G@��v��㣧�>=j�nB �,�R��tc�10:�{s�q2le#R!���TV:��π�dӉ̩�6��-Zn�H�Rq��*=��
��|��]�kp}����Ze�U���q�+�Y܋�0��b)Rg`yb�b3Op!�נj�ɏL���%��0���8{��������%n=�nz����N1����֨�+"�>ͣ{�DşE�f�2�ڸ��.��ծ�����}^�D3ff����E�֤�������4�5c�.�Z��Kr�I^�<W����D�����Lg
�/n�8?���0xAj����U0z�Q�Hd�<.�xy�^*g#-���NNO�J=�Fϥ8����T�j���P��Z2��1d�
���/,N�F!�3�&n���#a!ª}�,.�`Z.�Si�ڒ[d��62��STC/v^��d֎���h����|�H٤���A����6�q��ĵ|����ճ���H91��j����¢��]V=װ&=e7)�;][G8��Ӑ:������ާ���1�T�l�,�ϙ�a��$6�\�����ؐ����C���*u�,n��_�^cl���`�֑Qd8.��֩��G�Q��9:3�^�he@:,ލ��d��9f��-�
d��r��O�0��&�4�7)�����t��ǟk�M�2��^c���Qi�:�*J�i���L�7��AUf��	=s���6.�4D3}`�ǀ˚X%0�W�_|��R��~�W�b�u�'w���]Z���lwf?��}�:��Mz���.P+óT�r����Uf�7-��ohU���цc��5Y�Lc�U�m��&�`���O�N�f������?�`����i
���M�q�B.���m,m��(�L�nj �a��:��Lw�^���dAS廿���g��o�����U�f y��/�$���%�j�U�u2|P��epP����#�f̖
L��,8�w��+ 5����J�����\48�O?�, 
.����HE��s��A"2*I�T״L}��!o�ns�@R�Dv�H��to���d-3��ʸ��M�.#�b��rՠ�@!t�I�Z��C��y]�y��B��x^�esր��M���~��8�Y�P�����`�E(O+���z�s��u4s�X��Y��	�x4�k����,�UZm��E8�h�ؔ�TК�u��Q$(@�4�nj�8��-���"�G�������0L�

���g���嶀�cN�7�~[�ԮZWB�P�)��t�q���lLr����Z��fK����8M�*��1�i��za�������W�v��u1z��N���0V�ųq����hG�c-Ց�~&�#um�:���S�@-�.�bF��8k����[?��借O��#���X�X�5��k�E�g���53�q,�=��,�Lk}+�ք��DjsX���d�)�!�{t�p�4d4�^X����Y�.ߩ5���>�N���T�a�W=�I����5�9��U���,KĜ��#�ߞ���.-�� ܨL?mr������Q���m+kI�k3S]
l���
��XV�{/	���ݟ�(wH��9콤|���xD�Z��\b��Qj��s�7@*��z0I�M_�~r)B�j�[U1h�iDfu=�v��Uu���b͕/~�e+����񇳻h�s���qe��(��A�c��t�f���'�8x�(�@F�%ɓF��J���8���I�����˄�F�(Y��e����X?���D���&s1���A�@�g��_j�f���Q2�f��ꃖ��&R��� �Cr�U�f]��z,`A�m��u��бӂ�8W\�ϰ���u�m�*^Z���tŕ�iV���D�ժ$q|��И��#�ުE�Z���'jJb��o`Ѿ{��GX�����
��8&b�Z���D~o[*�;كbO��O�R8&�[��ip��*�SA�\X%l�é�N�`CňeԅEF���I��#�yK�,�"�>A�@��>s�Z*����'(#�ͽO�i���։w!����pe�&�0ŕ`�>o+�8���<��aH�@V�d5�q/��-���+������9'�YM��k�(2�Ze+�$k�nb��53n�B��
Ms���`Br��1�T�}ZU�Е���6-�'E�z���R�(e�D�jn.�w���0儤���,׶5*}����h,�§VU���^R��`I���n���,X�kSb�B��,��RU��#��/�
�Q(���7�����\�����//� �K��%*4$��,����2�S+X��7����/���T"����I9�k?�6���!���߂��
LG��3K����H߿��)8�ުJ1���\*�X�u���A���-��l�Z�ٽ�\������%$��9W&sW���Qfy�d��*�j;/�Wl��g��/�57\׺ �I[����g�4Cm2�����I Q��䛼t���0̩ R�Z�&�?������+�UvΝG�c-g�U3�M��Ґu8q)L?��{����
A]U��$��ie�
��.|��2��V�@���w��5�
P���^p��1��߇�#�D1�s�QvlX2�|��m��!��i���FN�_�-���y#��Ux�Uޙ��\o�]����V��BP�����+����Q�:�dp-bLD'�闉���S�^h��*�ٜ��ֽjmյU��9�?J�S�pm:���dp��f�7wB�@�`�+
*cӑ�I� �	lN�e�V�ѽU[r��	���~,�BE -R���"�5�DG�������/�������
C�?G
l��Ŏ���,�y.�<v �M���V��'��E��J~s�}�r��vQ}�Zе�k���v{��3P�uD�i�jO'si�
_ZY�i�	�XU&�RU�V��k] ij�X�ww�N���;Z@�-�iE+ú�9�L�TË]�e�R����I:,`^WQx}^=W>�d}Lۙ�|e����W�?���s]�d���Y�\����u���j�P �Q�����o@h�������Ug<����m5�V���p��%4�&��}�}�r��Ҵ�OG+�i�����e�P	� 8,�&����&CK���y3��;y�ܓK_�-�f<r�V�{���#_��a�nY�8��"���I�b�,��%��~!�Xu�s� �ј�[S"!�8Ǖ:�Z�ɴd�R�O���=+Uͅ��p��R#ʂ.����F2\o�eWҞ�Q����nnҷ�f֒���M�"�Qu�D��*U���J$�?Y�G7����:q��E������1�w���&OLtP��F~�*�?�e��{�˵b!j��N���+����i����{�R��d�B=��U���7�H��ju���E�G�r�Խ2���6~�|�\�Y�U�aډ��e��#��<�)d<7Ԉ�:�kZ�zs��y.U��Tw�դ"�(��+��cʂ�1�� �E
�ZJ,ڊe��9,����l˛V3R"�7��t6e�hJ�`�Yp�E�,<�
"��A�O�H���݈�"�-Tmf��a�����0����ɭE���wnA=��m�j�@6��	���X�6y+
���!V���/�>tڳ�ru���l�ɩLv3��n][T�A ��L�0�j�)�V�g�!�ՙ%��<'����o�2H� ׫�'�5�1��k���5�=�ԥ��Vyp��b�����:��B5b]&0�*6�۹wŤ�,�W�cq0�x���*<5�)�k���i�JMѲ.������1�;u�m�t�X�khr��:Vk�*�5�G�@W��� �a����P��8�����!����Xz�ss/���H�z/k�q��œ�h"� ���*��8	�h��¶�2(Js�P~�XQ���:�t��}��xx� �H+dI��Q[���h@cwc���<�U�#��MC Ъ	=������R*Q�~'(��p��hP[�"�VZ�V������h�7{�v%7?	��[�Q^�lhў�>(�:R!�),��:^j}�Vst�<�$��`%{o)A����¥+���wI���ɳa����[����M^�])�x��K���C�N@�q>?�����/�N��S�D���P,h�nB6�D��nH�`��2*>n٪ԅ��bv��w�;��r�W�0~c`�9��e��HCɒ,R�Y��ŭ�u��2GƜr᦯�<kk�k]x��p��|p�y||��8����K��h4�E�[x)~c��=�ִ��Yf<�n!�n7&���q�W/SD�9��c�W��7Q�y�>��9/`����]��-�t�e��9u-���)���rvCȩ���;V���xHa�be,�5�CZ[��d1���t�[D�p1WMx+����1�p�N��)��&�6A<e�p㓔9�9�O?W|��u{����cU�(����"i+�4G���Y��(-�!����I܊&��[�J�{h��@�̡�f��of�ϗ$6��Ra��֥��X�a`cD��}�PG�,�GNX,Q�s�G]ʺ9��Y���8H���+ei�P�E�Iq�t^���'��h[u[���ͳ���Γk��	{���d�םɆl�s�P �l���x�)�.�͓�#��A��Q���0m�˿G"�jSXA�zJ��*��eN~��.�_��]y $�&��5�U˲[+֧"�:U
:ywO��a��xqE�^E]j�Uhdp��&a�7I����,u����>��C�����>�A�Fˠi%��|�XI�C�3XXҟJgsۦqW`��{=���;�֢�t�d\�A�B܋؛Y;�7N�2���Xe��2x�.��C��:2��Ff��l���/GQF�Xx|��`��xr�*�֦~Zh瀯 �9��i�.�cb��, ��3�hyԤ�,��"ܨfQ$hKj�Ӻ�={F�Fn�(�.����A
�U-`�|�Ȳp�;��Z�&D�FD�@	dIё;�nխN�9�l]�Ǩ���U:�
�p�.
���l@�<��	��FtZǲ��&C����E�b3��э)Zѻ9�$���ԅ�Gv�ޖ�xOS t�:��z=�T��鰪E���`�����o��&���տ��^�~���@4���{��k�o͉�C껜�]��e�,�\��#�h~T������*� L�>�m���kL`	�����2������,���:Og<.�ֈ�<@p�
>�z25:^�|����-�qL����+�|�؎*���g�Ï?x��Y�^37��vnN^�gK1 P��^���Or�pY?�?H�i�����I-Z&04�-m\�]�G��h�Q��U0p��7��/��p?@�:�i��*1��|8�WQ�-'T�p�9�3
��3s?��IY[\��NsE�|��(w��\ub?-M�@p�Χ��`���2��ë\��9u����Bk�>\Z�4�bU��"%�H��(�{˺�;18�ef6Z9#F�uהh	��qY���R��b�vsW�E��b���jD����qF�KK>�g�0��誅��F��&TJ�H�d˗���4�Qǆ>����os�ݵ�aZ�9pts�ɓINzue���'������0A�h���4�� ����Qg\ ���8�k�v�Ĺ�@P��2�plT����O�����@@�2�p�C/�N ��h�tb����H!�X 	�/�H?K3�L��u'��6�L��Z��QM&����O� [QG������*T�,���� ���yC��O?IU!���ڪM� ��i�2g2iͽ�U:�I��ڑ�XTV3v״��N�-�쓼J�Ś^[���,�.�, `�J:g1���o���^�H#�z F~77jϖ���"�lI2T���"&"����u�E{lԭ�A�"���5��ɁV��}2#+�!��h"��p�(��Z�3���wF=�FE���I6�\E�Y�q�Zc���	��Y�N�̖��[��]�7�w�PR���	�4��3c�T�y��ֻD�/hY�7@�iXU?�@�}NM+M?;��)�x�&��c���亀�
x�Ѓ�ʀـ�.��j�v��tV+�5N"�/�BB$-[	g��,"'�����U�����w��l�ȑ�~Sۻ	���v���zʧTR����G�q	�h>m�h�O�� �r|��7�+
u` D(@��`a"��h&7�%�����L�/�`�Q��{#U��PK�l��Z��.u���%��\����	]	��G�Dp�qM���n	�x���ԉYp�G���8y����K���{� ��
,�_�Ż��|�l���]�Af���=H�����廏��&=I����vvoXUɯ�v���{:�$%�x�������9���w�Ǔu������n��&\�X1���>O�\�CJ����
�J��3�xn(��Y-�z[n��ճ��x�nmv�?C��6ɓp��;�B$��N,�y����}�ׅ�I0�C��H=-R;�4��a�:�:zH���C��]a�M-���ֳ��bra�m��0��r!��:�NL�¢��άOrx����O̪b�G)��xS-�܈��_~v] �Ѓ�R{�Rp�DD_�<U���Dtwv;�k�����E�y�h ��"����? � <�djd��k���,����e}-�ը]ʀ
?�RX�O�ZP+~�\`�bsf`u����~\�U�� Rђ��t��#P�}���} %,;p�8g�����4 �n�%	)c!��j��Υ��[kwV���L��������}c�b$����g�M��F����-v���Ng?�d��a����<�@�|�;��Ki����Z���:�K�֚�5�|Rg 5�TE��b�.e��	q�j/���h���3Zؠԃ�V)ӴRAhp��rE5XrU�M7�y$A�4@�,�c����4�,q��=�A���*�M>���b�±��V�<PX�8�u�9���b��Q���$j}�N�7�5�&�D�uJ�%�F�t?���$� �O
-7}��������̇@�ߩ�UkV08,Bd���X��&�~^@;�I������Q�K�פbύ
�"�-F�B���_��W��뽀($6�{��g�FD���6L��i�5�b�<�4�)��+� �p��#�c�i��P3�f����R�p�)��D��֪w�����Y�&b�~V�h�[�2!����.:��C�R�t�b4��0��|�˿�M�������3�7@�·y�l]�.&顡��:�X�ݘ'�{�g����ʻ5�R��R���� �w�w���0���ØP~��:���`��>��*���	^���Q��T�Q���Z�оBiG��b�.���ޔ�	!<�j5_���F�d>���Tp��"��͍j��kVE���'+����]*iI,���OKR�pcЍ|o���Ւqm���"�>q�K�2!���E���R�쮑q��v�K�o2IKi-W!�X�Y�NԬ/<��S��V�9��S����ϣrdg r�]~��JME�t+�p�Ά�Aq�p30�qs1�-��5�8���̗;�]$�mǯL� `�+v[�*���]>�9����6Њ���R�8����UF��m�`�sZ�f�N(�޳W>�2��ƅaQcB�c���
��N6B[�@�rp���kĽ!7.2m���-h�M���`	|�Jy����$pz�1w�i��<+E�2/�9�s��h�wP��.���\�K,D�����A�,���B�Y,�Ӳ�� ���&�4�:�^���}�ڼc�ޞ���ƚm��oG�K��׺1�f�)����}�'� i��=�������#b����m����Y]m���쾦f�5����Rd<���>&�R|٨m�U�b/aqk��8Rw�$i�d��*au�q���DW/������!�b���U0N��,���E\�w�����E����]��������wޤ_ˑdM;�Kuc釻X@��<���֞�Y�e�b��(nם��p�*�6�*D?X�#�,�O��cY����Z�$��ϼ�7�XȍU��\��NN��!@f�\&V�^'8\0<<3�h��Η)�6���dd�*���e�A�܂YD��>���-�L�k�p~b/s�C�1�E�=ͳ�Qg��&n�a3#���Ζ�v�x�=H����4-M�7�?$j�xG���:d���2W1��yRۤw�I�`�\e@���+bqE����xܰp�q� RC75���ܔ4��h�Ԝoy�ng���^�y�Tk��Gs>��ɼ�aEG��IAɛ��'�Z���p�Ck��dј�9*��,��V��}2��&~t���xl�6��`*��k�T�A
W#i\.�A�dň[_Q�;Z:��<Օ��9���4 ��
]�;͘�ϝX�YXJ�^Ӕ����+˽���+[��.������2]��n=��w�� �<��"���#Hoﴄ��.^k>4��B�+]ױXI�y��~�Nݿ�=(~+�o����y/�}�n,Isi�bU��j�=�d%YQ�hc���p�q�n�����L6ĠF�gPy��$3�"]��	 �a���\)��՟�j�����?��F�s�XUQNN�\u��ffɄw�^����%|}�"Jd;�>���޺�j�r�bsu�{K�"�f���h��g,����mndS��wV��J��Kֱ��σU���Gi�RŃ�h�GZ�5�C�+`���zb\���X���a��˘8��R@�ڼG���jy	>V������(�X��:�ǳ�rKxs���,)�Xa�*iE�0Y���}�s��װ��½̀j��k��6�B��L���0Lf�Х"��Z��}�!y_�동%z�ψ�/`ڞ}biq����j'�(6��6��o=�Y�*�W e�r)���[��Av{���}��|�o��&`��o��`!ii=8m���]_��	�������ಖ�5D�Lj���I����௿�*���_�&էif;d)@�|��I9�`�3�3�PUt�U�A���d���c��Xf	Dq����"���E�,<�VЧ�^7!��o�MAՊA���叿k�ҏˆ���X��ِ�xa�q��R�z��r���x»�}�=e��?
��f�4��Sa�d�R[����R��^Ưb�QՀy%r$X���z ?e�lo9��K)���1k�>X'�I� ��Nb9�
`��,��~\/��ϋ��{��M��f���:�2��FO��F���"`�7��3ZS��e^Z��{��8����5�,K�2��Ԥ��Ȧ�F�d`�cd��`��F��c�R�B��ˀZ����3�E�5Ϻ�Ӧ�v#�,T���"^��Nƅ��0�JY������`�>���j�<��j�P7��b��%j��b�e�NV���p�]vL , �g�|zN�8�d¡{�˿2G6j����Vy]��C77���H���]g�w\��;vo�M��߫��N���0b���+��������ɤ<X�\�HɒZB�<�mϋ)~�i��\��|���d��BP�a#��Y��)YM+�ͪ�l�u�S-У[��4�E�����St1�/�KeQ�ײ�2�Gk�J"���_�1�qy:>zYA�)%N,��H+>k˛��(M�R�;t�˾ؘ�(~P���e���.HHY�y6�F��`�eЊ%����&�R�\�U�V1�wL�%���,O�=�����}�_o���|c��Y�6@�_��6�ɩZ�x�Jg]^?�{���*��lj��N�#j:^X��ǫ����֟�h��6S:�s1�Y@�:k�#��E��U&�7��b������gӊ�f�D����ȿ��7
�:�%��k��gI�V�������U }2@,e��"�`j�V84�+�O�ĞGI �=�Ϊ��Z&�^�N��ں`z�@�Pf� 0y�3\,�����z� RXKHՄ�@J
����m����ZvR��U�?��k�r�6�b��H<!۱��b�9�h6���'��v�¼q.*����������}R�b6����o�L<zDNI:rh+��E��<��rlyz<�<���3���/�)	ܠ�
6�O�d�$��9���l����7@�g+�[��$)�''I�/Q�v&?],ӰV�K�=�(�Ǔ<�nn���M!#��<�1V@�j���oZ(5m�\�<�:�H����v�k��t�9���5��Å�J�x�/p׬Y��v�e�	�L�/����m�	GUe�oP�l���v0���}X����N�*�{=�Ț}W6�*�òz3=4�FMND�z5�a!�ߛ%y��m׺����#�
7�V�]�E��Ӣ�l�w/���oJk�����8i��p�O�Hv�|���5���� �k0K¬u���d����y���C�����?>.���$\�dUŊ5�=i@%jQ(�=\���h�YEs�(&�4x;��;õ�l�,��~0O �:��L/�C��Uӱ)hK�*����9x-h|t�+αiZ�i�z��ì�:"�nX/ԁ��ZV��&N��!u½��a3�c]ב�&�"Sy�O�\���C q㥼 <&u���sN�yQL7���w.F�X�E
P����kCN"P}��@kؤ����m-���^ܤ5xne���Fp�`�*E��}Cb/�!u��U��I����Tq���(;�h XU��o����K������U�U���:G��s�ǹ���e�K�<�i�h-2A+�)�mJ]��5��Y�q�S4�u��yʩsy����D���u��w<��Z�uU�8.?�"�9�%7[2V4��3�sD憖J��BO��N�@F�6�f���Ho'�*[ �s�e��%�j�S�I*��|��GѼ�vek����՘;L13����6`c!o�5NwBH*a���d�Y:�j*+�[����N� hXĄ�@�8��nj,2ȸL"�@	��*(wC[�*J u�y���WB����Cΐ�J9����x������1Z��Xm�6�&��rR%v�^[4�G��eN͖�X���V=i ��/d�-o�T|���y���ۘMO��u"LΧLF��ٌ�h���?����U����ִ������T�iT7�--�Y��Ά�d��ڤ�jY���"����9 ����zi�굽�F�|@������RU������,��i���n��BR����q����(��`�0�sC�L��2LO�W���11!~����n�j@�+f�s�z�t�XF��I���Vf��je,������h�p,&��1��,����"��."��&!�o�>������'�}Y,&X��rJ��Bd�I1�$[�,|�MuSrէɀn(6��>�jB*O�g<�/��r]�H���ʳr��u@�Qg��C���b�}q�eO�i����V������SaOx��YyU5�g���d
P:Ʒ��Ⱦ�cm!1�#�����Srg�w��F���<+R+R��D����1ڜ��c�>�1�4��6�3���uf-u��o
�֨2Qp�n6�:��fEYy{�����u����щϾQ�Pa��xhj:5����+��mj�*;G"&��2���!�Ɯƕ��Ճ���ӷ>Z�(�i�o�A�������U_��k�z�]H^�����u(�8���=Z;�:�<�L�B���&^h���!X���q!e�U������'�rÒ�SS�m��X b��|��&]��!;�<{ƌ�ܢ���Q^���r˃EZ$z,"��w� `�A2C.�AlO���I��\Q,row�i���y:*��,-��
Pj��E��d!���#����xJd���eH�r��)�-��d:'>���;����`��̠ U�V���mE�04k� �uT��4M�� w �f<��F�������d�9m�l�GkU��0���	d�z�5ǌ:��V�l�g"�C�(>�&Dm$7ٝ���?l?2;�a�b>���~�f�V�������%S�v,�@X�k7�D�b�cށsv�L��Hq������}0ts#��0��e��ӆ,��S�;G��֛K��y��ۻ�=�Ju(�V��2}��� �ǣ�(c~P���ޢR����@���ft���Y�F�Z}
R�$cP�|}�\]e���y��|'�����Q��JA���R,%����OU-��źā��*5�E���ɲ7����{ʁX�]A���\�l�C �e�He0��k�w�b� ��,-���,O$��i��V�¹���1���,<�i�o�-�����I�Fǡ'��Ⴠ�6���2��n�,&��kC3��B�0���6M�e7$ = Ǯ*�<�$ޫ�`S��J��IrD��ZXf�{ �ů��" 
ks��\xxH].U4h�^X��>�����r.¿[�����g�,��8���l�|�N6�/�ƚ��gSOX.���⫝̸�`R�J$�̡��A��Yͫ�*���k~Dm�㳼�VlG:+i��A��4est
�F都5���59���,E��]��Ȅ����r����H�E:9mPI�6�v4��cQK����%ܜ���+��Q{|�{�Uq��E�� p� �{��Q��i�Ө�R�SI�Ԗ��G�Z���w�mč�N �#u�]ds�h�"�W����,4惣en��9jiD0�`-݉&�����|���2v����Q���\��`�x��
m�z;�Iw_;�N�#�[��%����{'�9珬�c��l:r�Lb�¼2���5N�2��EB�����>Z�� ��w�x(=�\?���Jz\[�Vlg�b�TJ��E�4d��b�!��wH#�J�[׈&�f��p`�fFf�6��ڍ@�����w�{X;����XT���(�x��N~+:T���:��	�
Ny�^�%Vn>����1�$,N	,8�"�N��| �|�:Kj`2Yj%���t��F�"3z�U���ͱ��&",���8c�%M��{36�;�h�j�UW�#�s*Ni-& �0O6��-{��nQ�F[�w�P���e3��b� �R��-s}*��0��B
*�2�ޫq�&w�ש�`�;yW����jR)UPx�!8�AL��v0p�E�j.ގa6�z�G9�F�A����Ң��b�ܝ$R+u?M�'���x�"����I��e9�U����ֱ�O���_K���kv�M`z�����?-��r���í�uF�t�����wk�Ɣ�dY�J�c�1�yp�TZ�ًwP�P�fB+��U���H�{.葽W!b{���ƂMʱ�w*#��HA�,�ld�@*������ʤ���UIU��1.y�=�F(��Q>p�NX�8�gQ�ה��1�ai��A��0,�\xy�l�l�<�2��/U;P��S�}�R������<{�U>����C�@�պH�QG���K�o\�(�H�\�&�#�\��	X��V�V�͘E~kYO��>]�s��_7Y_����t,]s��z}	��kJ�5X�M-lm������]�\Ǒ�-3�zC@�C�/:z�����:3g$��譖\byann�7��M�R�U�D�ů�����#� ��rրٔ&!����X��hbrڕ�x���]I��+׽0������d|	�4��Wm�<!�S�?\������{�^RB_�t������;o�a�=� �葪Ur&��	,�x^Ҡ�]�!5j��9N ��=0;��X�l&&�Euj+��l��بxl�zVj&���U�~e� m$>������U�nt�mLz�RRY)�_<��i�<R�'�ў�M$6xRi1#j�}'v��ÿ��^��-\��������x�0�',�-�������xSN�Jm�Q�p.�#��������=�0��`-��xN%��L�4���)3��41`�#��&<��^1:�BoA��2����DI@$���\��o�-ś+�*F�`fm�x��r�"!$�,ym�z Ytb��y��y*�c���;��wh�����b�(z�{�Q�[�����D!:!`ͅ��^lY���bc=���M����9�'�R�\t��y�j�Õ�HfMb�x��m��b��u'p�KHoBi�~w��,�}$T�8������exXą[aO�L~R��ٿfy��w���O��#U�T-r�9
�ڨ�uR>��T���>�����W���Aԩ��?%�7J��YL,$x]�a���y�87�iEuR_"b\J���V6T$h��ԟb2��SP}��:�Z�Á�'��f_ �\�3$���d'��6X�O ����a�'��.~�s�C�.� �<I�e���(�['8'�='o��G�vq]$Z�q��X��K���s�)�a�x��&m��=�j�:��5��7"&��!k��{B��t��{�
&�ޫ��ދ�jb��{���tC����BnҮd��rΚzP�h!�J�\ͼ��.�"�T��cN�^�n�Y�v!�/�\)m�܀IV��]��WF�ɓ0��t&����z��א��K̸�H���*����6���/��͊9��yW-��eF��QB	��h@�$�WKD�u@���]j��������d���Ζ4��,AO~'#1K�t1\b�D��@윺���r]L�јY��ML��=k���v��m|�:��Q=?)#�����&iR��c����Z�۪�7�6!�F�$�'�q��(]'p�¤~�.J�D����hS��~»C���_����~?:u��*��2��COvDh5�3��Kv�6Yx�+ �g;Ο%C,��$��~j��.�qŠG{��J��>�����y��Cv�8�t�d��~�I�,
����&��^r��ѕ@CӜcm/ա��0LQG��W�ܸag�L�%U���*C�h��;��=Dm��؏�e��cV����3 �%	���G������G[O;{l�;��m�EO��}��?������0~V+�#�dE�ɾ�t�S�o[B��0�U�V�Q��Ѽγ�Q���/Rü&���%�����^[�#��8�B�J��:1�D�7�ʆ���A8��c�,�`@���_�YV����C��Nk�;��1&���8Ąѐ�V'�'Z��Ε!|��!�ѽ��j�:�9V6Z�ic<�lf��g��G��9B��k�q!����<�U��2�I�E�AY�,�GVڙcd���Y=2�ΠP��tj�QY����ƻL:O�I]H�:d��E>�:Db��)6�H�*��nL���������:���,Fe{�ƵQ(q_��Rm'���U���H���*����zD}����������E����YQ�'�"��jG����x�Ӕ8��m�c�7ŝ�KQ���&������~�-Ϻ��*'�18�$��H��LS�S�;3��\���ȳ�,����x}w׽���x���b:/�/>n}l"�F���'R��5�E.Ae��Q���H��֠ׄohE��u�i�$I���Ʊ��
�5/������v	�ur�L��9xE�A�F"-����Dw��z��V+ؾ:�e�,|
C���E�Z4�����{�F����P����P���!����N����1`tL0�Sy���0��|���o�GPӨ"��e���"x���h\���Ԑ\'�#øj1[�F�u�uV�t�Р��mdb{T�g��H|�����!u1��Zw��8�����9�oܠ��O���|y.��0�qD[~�.�(A�k�f�h1b�,'���1��Tm�/�,�G�j"5�SK�ļ�U�d LSUW�ռmw��H!K����pA���o�!ݹ\bx��W�P䗨�XU�e��,7a���&���vvj�'�bm4f�����V�����2��v�urm�GSvTм��6G�N�q��n.�n�֐>��
�R�v�4��Y'���������^8[x�E^!6�S��Ͱ0���駟�+�LY���8c1�qN hN-y�4�r.C�2�@6�B�y�&xE��q���E��e�^��7/�h�V��5hZ�;T�((�(��ׄj�ucb�T��^�{� ��w�f�U��86�Ň�p;4�r\zx�a�[}ڨ꫅�%�4����.�b	�՘���3o�Īʺe��?�C;zh\�9|������0O�!�&�^�:�K\�H�E�:�;*�g��ĴP�a���Yޭ���zx� R���k���g���&�-(A��=����p}4�3�{V#]\�� �?e�w;�#Rf0+�XյdR���klb<t���}`�	+�Z�jiyT�-��<�'�b�\I'�e�"�����q�[;�ｙ�8��6�/b��"�KB[ު����|~�������ܣ6��8�������5U�]�g�g�^ӧ�	j�L[�|�9E��"�؏A���*�!�a�H��h2H�0�lPw��&F���Bc4� �j����y�ڜ�l�u�
�'V�D6����5S,�̹��9���0B��%<��3���3C+lr�a�x�<y�F��Q^_�M���f���Ä�_��1c6���~Rub[ԙ��L�a����B8��4��Xlx�y�&���VB�c��/�BcX�z�Þ�[N��p�b�{�����5ʒ���O�����f�L��CHu������Kld}����`Ʌ	?7��S�a@���!&sp��Dխ~���eyȉk)~�y�N�7�������*�a�OJLL�ǆ�}vu�l>�Et~-H��X��&�CLQ�M��Vp�����t�f�?��T�O�s
��*���NC*�#�P�h�H�s��S����������Z������ap���>b�M�\!�ӷ�H��u��joTɚyJC��y�m�Y?9	b�^��3j�S�a�>XK\��� 
s1����y�p?ۂ2�$�F�ܱ��C��V9�p2�h�f�I�o�:��J�q�ZiL{`fɤ�ׅ'��C��'ǌN���X�0Qᢼ'z��H_X�Q,���v=�΃������!�8�%_��ҙ��^z)�Ѽ֫H�J)Q�(CȪ�=&�ư՚��Y��;5�"E1u!�&�
Go�l^&��Ki�F��%�/k(�d�#]X���)x���5T��Gj�ӔUnHƿ��ѣ�ѓ0�.�O�9�v!��e����l�؇Hs��a��?/CO��� ��v^=�q.�T�F��[�e�?�qM���z��7Zĺs'�q#n���k����3xR����kO��7�g70Z�鮒�sC��$/Űϕ�O��F{���SײTc�z2����=o;��\�p�)��[��o4,絥l6����8�ʂ-����}��8�pih��գ�ˌ�RJ$X G�j���s�%�w,-�q�C$ar�HE�=���|a"�O������YX넻�O�9������~�(�I/��bJ�����Mx�
���'mS_��̜�d-Q^�ۈ_���Nx�mRA�Fs�4Q�x�5��;O����q4�=ʚ+,�����G~8�87����$^�d��[�ko:^(i9�gQ��lrgU,��Pˁ���8JE���ǽ�R^�Fx[���%�Ue�Iq�j?@="̣��1���=ǌzu%�m>��>5������q��:��ļ̾�V�&\mQV��'S���e`cF/:����Դ9��.�zݠ�}
Q�������^�+cT�
�J|���M��еp���۳�N*eyh���9�4ȕ��o`���{��Pڈ���]��Dn�˵�!���y�۵�*���|�X��`"�������6�c�K�%z�%������J/�T�e��jG�T�fo�oebf����Xě�}r�S.��4Ҡ�i�{��`���jD�(;#Լ�0�x�]Jrp����� K甴m9o?��Y�"��/r��� �}9��'�"ђ1�Xm�˘�tƟ[�0��prN�ic�'����B{f�S��,ܹ*hpQ��0�����x�m�Y�	�0Y���[&k�x���81>Q�X��:�z)�s�)Ts�a3٩"�V���$�����;+�H>G�l^�������]�޽�L�P������LF��6"��C����sw�v��Z��9����>D|����Գ2d�bS�_TU�E���k�HPS���}j�*�ѕ�k��ũ@%
��FK��_{�_�R��}ꛊ�y��N�X?n�u�p�W���[c��%�WSM��j�	�+��{*�8f������������M�l�)	i4L:0V��l"�}���;��%W�n�k��G*�K�2(R����[΅-&v��b�]#��ő�u�Nh���g��_أ�K��1�s2��if=510��7�7���0/�Bc&X�k��܌~?GV~v�p
�Y�*O�)��
�8yr�lvC���������pb�y��z�B&��1�?��d��+V�*�F=���aT/��d{���+�4��F�޻��$=��% ;�D�i�O���0���]�=E[�@r>������bc-�d!D�W�K�|����PL�0���³��2��Gt��,�e�f~���A9.A�R��T��Y��־����Bw�����d[t�%�|�S����'F]F��/�׀��<��_��_~�8�|Mh_��ֿ���pÖ�8gG�}��6H<���bۺQڅ�&d�t�/!h��z&�zE��y�\�0d�0�kV#���Z�UY��q
�<2���pu�]��� ~�(Y�)NpyP���1/Z=��7|1�d�`���AӠ�Ӳ�&h�����.\��X������%怂�Ml��/��=R�9��L���ǸisTa���<�#-1���L,�`St�s�:l7�fP�hs5q������ߚdX�g�&)�M�����YZe����9[�DG�06<R$�f:;�Ƴ_�{aD��ߕ��T����z���}�v'~� ��1]���.l�r8̞@e���˙sH�U�p^�����T�'�Z<I�CX��mo˾c4���I=�[�杩J�uh�$��r���e�>�����������:��(�^J��x����M��.x�ʵ0B��1����:y`c��C�Y,�<c`-[X��d�)WCeH����:����6��������;''���%���I[��j�[W�Q��H��pJ*��=�ND��#eѦ�f49/�5�N�W( �?+k��P���P\����a��kum�PD|O�[{
�_��k��6:=�ţ��Z�p?b JH�dp~�j��hԉS��W�ę*G���q�T�S~)k��*���:��Z7A�(��
�6��e5��<+�x,?���Ex?�
�CC�F���Z{
�b��9`,��e�rث�	��D��v��6�$11�W/<6�5��4m�[�;e�hC�kQ	�A��XlC���.�Ö�L@����[�Q�SJƉ#Ne�^�Y�M�<BnV0����84:7ICD��r�K���Q�w"�O�}gc��������kXM%�`�,J�]e�u�@u�S���:e%˟	�Q��*,�1}��!����+����/�#*l��]�a$n�/T���M��Kq��:I;ym��
g��~��*R�������R�nW�\I<T����KPEwo��j�l���8�*4@>�T�W�YaPA�j|Iaq=V�k��mʀ^���`[�����-��K⻗�14bVTU?*]f)�,E���6T��;I�0Z��t�2,��^ᘕOa-�gpu�u�!J=���Q�n-���$zA���M�88������a�⌆���+z�4�T����}0J�"q)5v{=�*��UҒf�<��j�tt�V�����`.����ګ5��A]�00��k<rB%�@5G�9Z�!;��0N�)[�d+�*��]� �<�M1���~���%��v٦?-�;-�r��.7�j-R9�%��*��-O�j��{��S�U0�L�u>�>.��(#'{v8�wz�e�
�����Z"��7����?-Uh�lߢW]�ʰ��d�l��ڽ�`Cr��g��c�A�Q�3�rq�_x��U�[c1Z��Y��#0"$cA`�C���33YmjiR
������j4�]�Fx��%�1��*oSkc�5��A�Fqlhp�T��*T}Q#<�����D]�r@��/����gB���96��%�C�ɴ)��>UX4�x?�i�i�
������>60<旸D;J�(6����֒{�М}��r�4(��}Q���Xm+�E�+ͽs��v���#}��Ƙ �?pAq������=�����	ii����9ۄp��ke��������eV�^�%�.��M��U���H2�{O�8�{��y{3�{W�W�fZ=��&	a�X7�Y�7�P�n����>��bÇ����QӁ���y�8F�d]�e�����̚��&��B7�5�HQ��1"`�V.c�D�̐���j���7:�u_yֈ~֨^�Hݻ�|�j�3�����RtJ)#:5�{p��y��zK�d�4��I�ZxOYD�J�����㧨�)nr
r��z��Q�1�)��B;�ir��l1� OmH8���:K�H������/u͉<����ph��X�ա��&�ar~.7:\��p�?������Q�X9D��ũVY�<>� b�Ȉ*�=�w�!S�wG/FJU� �k�D��>�
WG������6��Cn�ݱ�27�˲���W��D�V��VO��]�
�����_\���»#EG-�����߱���U`���a=�橞� /��C��������f��x�/�cOZ2��E-�Y !j��^J����)BK��@���q��^�!3�P��0��#ᲄ�t���b�R֤����,�ōxmrF����6��/<�3���S�{�~��6�[��Ux�8�
Ee�m0��3�>x�ų��B&��8��3����ԃ�%Ԝ��I�,�d>�O�t�F�:,F�:a������6��C5R�i����^V�Vɬ#~iz��þ$���-���` ���w����m�|M[8.��{��"|w�D��gñ����sh%�V���x�B���$�y�Z�����vUE�,��0H�����B,�ˬ:�O�����7ՠp�(��^��ƌF(�Yv�;�w}x���g�6'����Z�ŷy����y�z�р<d��5�Nj'��ҳ7�c��e�C��iC�Ϥ��ͫ�:��J��r�V:�Jzw��<*/����n��c��x���H����1�J�l����tfƙ��1hs��	,(�jE4��hE����`�h0��<U�9C�֡�5����t�w<�Ns���G+���y�N��}�2稒S��%#��=��ĺ&�ٔ'���J%_�^�!;'6J^(��";C}�|q*��{��$[+3�S��V��ճlLXM}�֥:��{�Y�^>�p���S�� �]'�?Pڷ߻G�ifu�ɐNSbZ0�M)a|EybR��>T���:q�֬/(%��3�3`�O��K��R�p��c� �E9-�=(W�Q5�_<�H.�O�1�>gӄ�؄��җ��E	���,�x,j��ɵc����xn�_���X��U�$EBT��A��ۅ3��Fc�n�%�|9����#'z��z��r�Y�E�(*H9$r�j��=E|��zP5^P`&7�y��1���|IE`*�g�p�Q����.���q�m�#��;.�lXJ����S8?������'��`�L`�+�v������k��,��z�P�������y�L0�p�0{���]�qza������Տ��s�#AW��ɓ�r��;�/�oSk��j�57�H����u���[{�/���*��S}��(oD�H�p�L�.�)�2R�U]�^)OzQ�`\���1�}X����0Jd�atL�h�3l���8��:a��AM�v�O�-!�o[�M,�z>G�[�]YS1x��G��,�EC&O����՚��yj���Q��������}�]p���?y������e�F�޺��Φ߸G
�"y1T������C������&f5:\��ۇol|��po�V=t��g]�e�;X�Zb�� %BzU�-�mR#ֻ��c��a����s�,{����E|�x�Gw�l��
/�/���;CW�؄=q����"��q&��H�5;�dG����#�I���j�8�G\�WD'�u���?�P���d�0�'���oT3;3Q����א�X��OB���X���N]\ Ƌ"��L��P!�cL���	j� �A�Ę;#������6�B�sX��P���S��3<��jc��&���g��T���V� �7�1�1��H�H�`�Obn?:q�?�.�H�2��i8�%2��9y^�gF���~c��/��4��u3��׿n09e��]Q�(����L��E�ߌ����1�R�Z�٩��Y�K�y󚟻,��d��{S)}̼��;�� ��
)�E���0��66.�;]���f�����I┲��n���N���&p��Ơ�K�����f��.�e��'_�A�!��5D;����D�a%'����om�gf������A�xyk��P46/��Ͽ�l��9P!ø�7j��3���b�/�P�3��2����Ӓ�[�����+���5K��mq�s`�[MV&�|ѐ���1N/�B��14Ou��D�Ԟ�~ �����e���i��{��A�R"eT*w��1����5�H���W�Q&�?�:	ѐ����=�X"�Q#��`��yd�b'n�T�5��}��U����iHk״�~.i@􅢌�d`y+FQYo�9֛���+����y�0�*0L�ѹ_'ǽ��)S�d��~g!��:��	�{\<��wʴ	��N�]x)�`���Y�ƅN/����Z=��!�r����|�M�!u� �|�#C��M�<8����^�mX�z������NbO�ؽ;^���D��0�6
�aE����7yph����L�5Ż'.��\S���Z�'�2[��uS��s�Mc~�1w�2.�yIKIm�Kx]0*=Og?���VS�������o����1[H�m3s���b�EG��Ѡ
�s^���~˒ԤNe����I:7q�>C�:)����m��TX֏�N�6��~�a�Qm���jG&*�J�����Oj2�K˽�0ܼ�6��*�&���aZ����E{g&��(;U�-jYmO����NU#̰�Ru�����dlaGa����>^{��aP?��r�6/zƘ�@�y��<������Q�Ð�y��<e�=��M��dOr7�Íp�^4�������-$�͒�m<�� =�ʾ�ln�ML�r���Dm,F����Y��DLa5:�g����d��8��_ܠ
8�D�zS�t��Qy���K��>�/����/-���A
u��x�*N'1�l!�0���˛�c��S	C*�S�k��r���G�F��{��&Bz���/lC��bob���`�7��W|���e-_<Ǎ��(B�D��=�9O��D��z����LTc�{�R�r����������P�b��8���+�g\ǎB-��z����d	A�S�����Y	��5�'�Kx�C��a\$Wi	��D��8l�	����ޫ���%�UF*lB���䀩v��w{�|�z�3��;�O�@���5��й�s1g�̉#t|�`�`���zmH�K,���Jks�o�?��\�>�����T�L��40���(1�4xt�w��7<Oa���PWHe��wVJ�״�f
5��ryW�V0��!	0I��8՛��a6#�J1�p��Yܣ�! �hL2!z�E-:�@/Nc-�,#
���/�����3��N��U�m.��i�J`��	�:8��)���r�6��2�T<,S��^6�'�p������Fx�֮'����[1,�tB����:sC��%�����O*X*wduZ�^��Eo,S�9[���j4�m��6_Cd�J$���dD��_b�K�F�7�zC��!f�I���Ŝ$���� :DjfHu����U)yA@��1��jh/���)T��Ս,�܀ޯy�M���/�ϥ(pɾ�:u� JoT"�5Kf��+Ѧ����dᎈ���ɚ��SZ����T��Q�f�?/Z��PJXy<�0�� kM)\\Q�X�}��//��7N"d�1p Q�alY�o�c���/y�O/�5���tTJ7��{��Q�(b��7o��]���׾�'�F)԰��[g���P��d0��E��ް�H�'o�P���=�.3�u8ӵ��K'�*8p�cп����\~����l[<���1�2�C��%�Wj[]bC	�z������.��F�jh9�%� jR��
Π����R���5�𭋵�܃qҚ��E�J ��ߥ80i:���ƒ��|��Y&z)j�Rx�f<'�2.F��F/�<[�Cu�(�`�G�!3�<fe�go)]T��3��D�����3�e:��5<P��@���ָ3)��̣��sd�	���	�'(���I�D�A�����6��)�f�XUvtƲ%3�W��%
�֖��̳�5�I����z�Z����*�+��C��Y�����fϦ�xj-2G�����S���B�O�f�0P���.�;$JI�a�ؕh-BvIؖ��VC>���ۄ!������ :���0�2HN,P�#�G�\��FDF<�h{3��������`��B@?��`���kEbc�l7�}l�;)��6�wVf�ɾ����Ӑ*a�'��Gw�*�@�^)y�X!�kA8uK�,s�~O���&)[�;\J�nӒWUAF _���xYhPsF��/7Zk4>��9����tP�RO�����l����p������$�C�J�l.�*�����hU��Kx�T@�v1CJ�sDe�"od�UAm|�_�ͣ�c���E�5˦�iɲl#�7,��A�[0`4_���^�5���Mi���%��1���&�7�zEk���65;�V�1<oi����u�7��o߆��9�&�O!,W	�����P�5&G7����J:��e�S�T��@�kr-G�5Q���/�G�Q`Ѐ���?�:�ym����
X�FG�E�8R���k�*6)�h�&I4�F�*>���]#�������ų�<�aP���%���9�_�Y���7�|c}h`�@���{����}�"l�A�+1��hkR�j�ӝe�]�Lџ��c`�)'���J��ᆆ前P���e�}����K)W�_��T�\KI�)d y�ڈRG#1}�e��ݣahmۅB��f��.>���#{s�����A�sw��8Gr���P @�#=�w�ޗ?���������?���s]߳-ek��&�]�+��1b7H�b��g��MGB^gaD`olŐ�n0\ޓ�>/kؕ����������?�S�{��ŗ/)b�8��Ƹ�B?c^�="�RL��YNV"�_�P�9��b��W<VL��J%�H@�~��N%��~vo���(cu	y�y�S۷]�M��(_a�� tʕ�D�V�N� Y��U�H�N�!�Iv���6��r["��.����9���M[lEb�xRJ�/߮���o����?������u���6�0E�-u��x�����iؗ��>��("�k�.(�J2�7�2y����� �p�6 :�F��߯�~5o�.²G� ���}K���(���7r.6�j6� �dR�~뉦R�� aК#���~�UUh?{��Z�섑;)��(��FΦСA��j��3%%�:�q��� �,����Be�;�ڎ��5�Ю�39�X������eRy&6�;+ay�����簔�G�i"�/<�r��[�FKf��e��^���Z^,�?3���Ǯj�����}�{z�g=gh�����Si��R�rb���ـ���j������S����H Ó'���8��kJ��b��Q�D�+�a�4��Y��2���7�����u2!<M�8y��2����n�y��N�!$����0xƭ�
"U+)���J�������H`�~��5����yx����0����iT�D��\��t���R��nz�j�a��Rj�dl��F%V[�%1J�1VݾȖ��K���V@Y l���ٌ ��yA��b�fl��������h�0
|]N�J��z��V�vC*o*�E����2ň��%�tx�T�O�{4�k���L�JZ�QZhT�C�LQi�eF���fE$V	�Ⴭ�c�h��!�AN���\3�A��;��&�����>���*�i��WUr����?k^�v:?�8?ɲY� �#�!�?�o,d[H-�,V�h���!
\$q�̮�0:���x����TگD�œ��H8H���L8�ơ�O��9Ws�ugbV���`��^n-DEp$�NbR���Ya��PQk��9)Ǟ��jD��s�4��Z�n4�ީ7f8���(eE�����T$)�ͦ�jUR�#E(���?��_=Q(-���������,�����}�wkx�/�`�#=>E6�d��s1zzФ���\���MV�'��Ï�P��P�0%���~�nQ)��5ԻI�ʊG
u���+�Wo	��ݻ��~���l�Ta�a=��E��>����%S���?�`�����qoOV���^�z��������qfV{x4B�4����59-�T���Qk��jۧ(��|燽�w^���Q�0�a���(���0LTfS��d�1�f�5�Jl6���GG������k���m)�Ah\���6��*� �e�&|�a��䆅	\�W�ְE /��[;` {<Z��2��#(&��p�����B�{O�R���j�R�V`SE��#��R]��s#��7J.q�g�-t���_Z_����\C1�ʔʉ$������դk���p�5
?B�Ԩ/~
�	Q+5e�M���d���G��'2=)�&�:Ϥ9Y�k2Au�S�#0RfY�8���EU*��N�_���=9��0ޓ���C��K��̋���k��~�K�ʹ^QHt�T���{��|�l�� �����_*{'���E�1�K���axjH��"�Uޕ7j�U<�\S^�M�<y���
�a���"��}�O;�f�>�F����&�g#1g�c��J6��V���s�����n=��.m��d����4O�����]P���\w���g���5��5�}��C�\��Uh�^_�0^m`�dWIM�	"��$g��8�P�.���j�*�?y�T��.U>z}P�E��C\Պ�*57�xԼ�j�?���=���ڗ�o���l����A2�B�D:�^�^��/��g�:#�Ā����xo'%]TՄ�`f�\�p�����������]+����/�j�'�P�����K;��;;�%�E)U��G-���<Qy���\���q��	���sZ���A��o�?&�両QoVO��z/��"�i��RR�,i��8cIƐr�=HW<��M����s��P��<|�ȲN[�^���Q��!%�4j��9�i8F�s���XY��T��yD*���Qk��.��6�p^8pj}��k�ki=����Wo�h��2g�����AE�d�F�����N�U��gS6�-��ڐ2A+1�M}l��}��x8O��ٵc���զ>C%��(�9��C9���w�/25_�����p]уڱ�\bǃ�������>���d��̀b.�$cy^f/�X,����H�6�X�j�[�(� HFi�E��$m�4��3� ��?�33�F!ZԿ�ۿ%Bэj��$u�1���CM�T�d�j���o��mA,F�Q�r��tل�x���=z�iЃpo��l�:f>�Gy�u��W������g�y�ӺDH�<�4�U�Q�~�`Y6��>�+m]�k�l�k����56�u�F�F5�l���/S��M[ym2��dK���-R�ғOYH��z,�%n<���f˵���t���t�.4���,{�Ui˒P� ,���lE���C*	J��{��9�S&3�����M�Ç(��UF
xH�{a��Qs�J�,����ֺ���b��!O��f�ȸ*/�WF�$�g�����J�~Y�W��N�Pxs�^Ix/�p�҈j��̬� X��ݦs�H���htSyGm\A䕔&d|���?��&����Y>��C�����aSm5�'���]P���8�<0��γ�N��VZ�X-
�A.�k'�D��EZ6����������~�۸x_��-�1%W������$�zԡ����*�qK��[��!e��5���}��os���x�����o?��%����ŀM���_E��8��#�����*R3g��:3�]x�˒xp۶��ԃ,�8�5���I���7r5[�V�Ϫ�g~~)��z.��,��b0j����1A�	b�0���Gz�p���̵���wV��"T�*Au\��1pYǉ9E��"�ݶE��������z�=W�@�W���,_�T��yђ�y:g�T_21YfT���>�u�\u��m�`�cc�<�&<�*6�����a��g�ЛT�q�FM.�D�6��jp��;MJ���,�|Ө�����Iy��CS�g
U{y���w�)�A���u��A&��[;`LL���,��t��d�Tߓ�|�����qRx�&E*�N�0�Vds��"[�TRx����ʛ��Sj�k��-*�u),y���CYV8��{��c�	L6���k|���$�4��ήC�9��9�/�Wɪ�4������o���{e�����@[uq�-�EU3o[B)����|�ј
�m=�a�)��m�EV�Qk�<�}��O� �"�X�%�_��ˎ��ͳn$���^g�/�<@Uuw�������[F���6�+%7ږ��(Ө���S�K���^v�5��.�w���H��b�mS���]��5���%�QTs3��m���R=uTR�i��~�'b�D�ׁe�Y����L��)ڡ�ЬJ��RR�Ι��	������>�^�ad��O��t����g�=�0}&�K����k��u����~��(�w,EU4Ž�4���W ��{;������8����ѡSP|�m<¦$�n�6�������<�K�\zf�Ϭ��޳�uN����w��Ѳ5O5���e��f܅���>������y~�uO��_�N������9X�񴰼0���>z���S�]�s!o�`�Bk���)Zc�'x�ƍ�:�')\ͳd	�ͻ,��(I<���H��d<�ǭ��Ә�f�I.Y��
�dD��J�Y���=f/g�KN�|�g! y��n쬍��Ƚ@���\�����w�?2\i[�|zAQ��9Y��}uF56Pf��l���2�c�q�QRK�{_��x�0� ݁/�0���]���S{�I z��f����.<��m��jj��։��k!Λo�N����1�gAx�΀㺻�ǣG�hj̵���C*��@;�ܠ�%{�,�i� �\g��?�5U/�,��#����:�������mq�/����G�),�ijH`)��[��g$� ����_��z��D����F0���H����a�f�=�a-A5Ed�	�����9��;Ab  ��m۠�,�N�`jT�D%���:���e���,ڲ3�`�/���<�hH3�F���:ǿ*!�(�to���GUx��n�`:�2���9�:��&h�����춢�z���X���� [タɾ��(5����zM/��g��
���}P�z�Kl�����T�I� �yb���l2�]��|���A�������3)��~�'r�՜��E��$z(�l
1���t0j�rS֛�ґ��/���:��Eh�R�G�Yz�2_�D&�\�;CƮP紤q�P���fk�6������^��ɇ߿d�4�ߗk���<��Ry>���"$�?��5�N|鿯�v�Yt���p�嫗���K+��]3U*O׏��bSֹ�&�!Q�GIFZ�d����^G��=f���������ޟ{�v��_P�߽��b��9]�`H7Ft{�ͧ0^��*L�s�����۶�I�>��$�������(�p�!��=�H����	�6�U�q!lD����F�Q���L�.?=�-7^rz�^T.e�I��=�.�B�]�=ʠ��5��C#v=��ڄ<��9�U]cnO�jK$~�����o�_����B��}�*�a�ݨ0#��J67�y�!�Ӌ6�|�e�.C�.<��������@�Y�˦�\T���)a)\�2����S�Mc]o��M=I�J�\��2����#D`|�47}����9w{MX�8Ȼ���}{����Du\[�y�y�m��*�2�����^)u)%�w�ړ�[Qa}��t����ڎ׼�� ¯2�q-	i9(PJe@����'�!~
o�E��Y���z �j9�f�S\�=��%&���K�Y]�/2�$a�	̒_�.�
�����x�'~��m*9��`#-�ё& ��������߿3E&^w�JTzbݰ�ML�w] �g
Pj��!=k����g��2�z�ԙ��)h��&4ɍ zN�Tj2܆�	%w�\�mUR�
��p۹h0�ὥ�w�+��Z�� �r!<2QrQ�jC��p���~& �q��Zy,v�F��:k��?�j�����=�K�qO��~�Y����_#=Ϭ�W?��1��-���`�>~�3#zO1���\�2�� �:
��Ȉ�5l���Si�d�+W��M�>S&:�����ob/TPP��_��'�imD�ƴn�7�����T��8��������s������Z��[aR���t�q�φ�zj�I��ٓ\M���N�n����D�n � #�k�ɸ۳-Bk��l��Ҥ� �#�Ab�a5}��m�+�	]��Cx���l;��7p�~�����ӵ0�ކuMɹ^�k�����t�`�4��L�Z?��1vk�:�~kH���L�xf?�N���\�7���6"��+�� N n������E��5v��f����x�:@I�����EFpI�6wy)|ގ��}�w��j��g~΋�����>�Mua�{�YdH�#�������nE����o�9�l�h9���>DThw�c[U׉J��Մ�EFC�)���,ah��{��e���)�k��\Gj[�?{�~��p���B\[,�ox���Ǉ1��u��K��6�_?�ݶ�Z�6{
�Xb�0���tlX��i�:/^�0$�@�Os�>"�C��%�-���j7�Z��T	��E�D*S���\@&2`���3��|P	��q��h1!�	�R�=I��8��߀�d���2�{�H��⎈�ެ��2C��� �º�
�\d^���Xn����|�Q���ŸBHd_I��k�k.�x�}ˌ��-�h���U��x���G����^*���;/N��2O�g�9+���𪖆j[c�Qᥳ����S�j�#61J�?4��9|�Cl�S���	��'��z5��k�������Qׁ�뷭����gHf�����rx~���xi3�$lR<�F�	>�yB�2�ʢ.�@l#"���ʺ遂��2�Q]Ԕ�<R��7����c��S҉����S�uR{�)x��QJ�I5_l�/A`�n�y��E�j��k#k�ƴUx�8(�~����N�L:y�3/�!��.=�E���}����32/�g�Hޝ�m�Z�2�rc\)���ы����~�'Զ�%�6�Ѯ���g7��;��( �0�x`C����5�ľw���b�Ra���4�d� #����YE2���i�s���6�k������ݳg���>�_�w^���C��u, &b]>n������hS�ή���h*e��	*���	��A�`[7*+���}�����zzn�9�'eT�u������Fg�C��K0$U��<N�����	֙r��k�^�r"� �����k"���;���~�zޗ�h$�����q�ޤ�6�x��iv��h�v�����~�}�5K�� ��7	��d�it�j�ثطx�u�=��U�e����i/��B��8k5���G�7�F��6�^����$�\#Ֆ�fX���6ɤU𛡽Nؔ|�z�����#@@��:���i��n#Y�~��O�`�Ïߗ��?��cB h|>�?=�0�0�777�q�GIVGI��B	
��x�*6��z}=d�.���!<ٛ�ߕ��D�}����DS|aY���;���w��tvR�1c8�3�q׽�F�r�EN����g'{/�+�wN�i�r#5˲��Ն^}U��BC�WLM��+�~�N5�P��E���f���v�ۭ��t@����h��H�n��F!���Cքc�]F���)ڜ%0��~Jc�ؽ�6S&�����WC��+�����rv�����6�밐�)3�M��w�N�X2
�yh�E��Ӿ�0\ڲw�'(��8����E��0��=`�T꬧<�ө����7߼1�{�N����l��,�����!�B��MW����RaǙ�O�[g��,��6�+O���3K��L2��P�o�H�V��F�q/�*>�>�¥/"쒘N�Ŋk�*W��	���I!6����%���)<4�C������k$�,���w�J<����ь�鴷�%������wc�����	���-���,� _6��ڍ��ڪq���R8�a�=-�z0İ1����G���D�B�V^��p���]���g[ǯ�R[�p�u�|����ՑD��a��x���i�kFG���B���WzU��[ٸ��D��]�n\V<��{	��Rm���lLl�)�#2���Zu�K��������*: �Ǭ[pϋx�҇`��<x���Ѫ�umŪ1�X�GI���C[m�-F�Y����~����Z����UKl���`�K����_~|ޘn&��7��!u<G�I�|<F�H��j�n�%q��i�S��R������l�א�F������x:F�a.ZH)B{�,������o*+�0Xʶ��=I�<O��?V�&�������������?0��TyHV�HKF�s��?���~.�%��.��nO~˘
.�gD��.{�[c�}6��˦����w��:��Z?�-{��3���x_0��0��#x��޿3�K��`늻���e�N	<h
�
|w���q����Z�N��]NB�fztE����|��&��S�M�T3���'��CH*�#��&�0�L���S��ĺ�G�L+ `����0J�:H'�5��gc�Y������_�m��K"�l�s��5�z��%�V|��wM��+���襂5.O��ZR2���QkV����M?�?kH9���	�|p$��K�g�9Jʨ߄���'M�ݝ��AkI�!��в��JZ�!&��W<D�<����vv-0��;�J۾�a����j_\T�Uow<�$~�����(
����W�\4�OL@�z�"-Vi�I�eIuv���|ҧ�����i�~iq��m�s5�j�=VM4P�Ҿ�\��Q�YT��g:�yȃ!o�k���
�y��[�&���a��㽵��|i�#�v�@$��ʏ�+C��_�>M���?���[����D��S�Ph��q�}4��L��H�@������]�h��j��k�T��x�&��F��
��+���+�z[�D�ΨOԣ���{B,�E�S��B�m)5�=�{�/>����C���({&<���
z �%�ǣ֊s���|���_V6[h/l�	��8+��W2@ p�(iX�q�e�I��{�+7�G"<g|���ntU�{�����+xv��xdHS�x��Ű�X�a��P`�]E�z��N%�b��ՅNA������WqA�'�p-<Ykr���^m�8��]�x{2�2���x~��8���<�*i�;@�K���,%��k��¹Y��ģ$��;�T!��W��dּ�bg���v�l?��'"���}��	����%�ty���9F���.�5%� �O��&	VOz�F�J���N}mbB��r���*�n��F�i>5���)���&�(3*m�'Ƒ��K�\�S���QF~ㄵ}�����]�ѽ<Gӈ-�l�v>^����{{/��T�@�G��F��!I�hB�a�N-u�4�M~������m��<cH=y�y��� �	�,�a�I	'�H)�
��Y����8����;��kh�ɺi�$߄A���\8$q0��}��ou��?�P��O��X�� ���io*�mk�,��{[/��\�>�ԑ)0���:a���`-�����j+l!���1����}W�X���&��Z�z�2<�R-C%k�R�o9�©r��$�ԙ�O�1r!�uk:�/�c����j��Q9����?~��ĸ���>��C'1h���F7�C�eI|L��T���G�?��PQ�a���2p#ƥu�c�E;��jc��gi�+FI����u��$��1 �|�ڛ]�6/Fܻ�2ECΗ10~�(
�`��T�}�(��ꥺ��TSI�q?b-�ɅF\
��~q�e$��E�^K�	B�q�U�ᯚwQ0q!]���1�k����J��`z�7m�F�f��a�˕u���My!ie���n�H�m��.:�H$h����X \��.G���;V������)������B�}q@wMلL��5ǯ>酵 ��$�����'�FM����B��<�9}a	2�ܻr�2����@�� .��
W1�tro]���[���G�~פ��&y���!�q �]^q����b�}dI�6�,/`pzp�* B���|c����r:3��}�m��~}o�u7}4^�%��6��L#&���u����:ϴ�fJl���z�,��&�h�\�o2ۙ�e��6<�h��Oc�H�!a���!���ܰE��U�u��a�1��3�����@d5�d�ԇ��j�N���s���!��Q��	`�F?K)�{�&�_ّxY��@���Z�3�g��9��M�}��k���'��5���-�4��R�B�q��'��B����]}3�v����������=/^�*/_�`�����1�>��74hP�G��1Kltz�7~Z�{�!ԅ���t{�4��u���<'�5AL�K}�C�����fg���:{��PxX�'�pqC�!�H��Ґ>�w@9�o��,סni3X����.T�|�,(�IpN�0����c��zT�xU��m.H��~[4�CT��e��}���2K��a5պ�,!��,Y-���2ySA+�`��r9/�SX�y�U'�,O��?�����W�S�8&8[Sf�ü,�T��vC�gC�I���������z�1up��%>\���͕�vN�e��$�ޯI�y�돲���6�����|��Fa��7��L%�]�Ԙ�oݙ���ƞ	�&�W�.	�W���M�t&J}���7����po���2ʵQc�_��~�j�ƴ�W�2zҜl�Z��`c!Iȷ����s�kC<1�h��vOH�y���0t�G�νRS�V޽s`�@�Tk���<;�35����Ƶ�c�7��)\H�^�8��"�q��Ę��{��.��Zg[8U����Y]��U��_�����5[�:�b�V���A����ǹX�e9;�6�W^D��6�H8�-.��FK{x��0��a$^y��Ǹ��ޕ�>ءz�y\P����#��u�{e�^ǈ�θa�,�Y6�	��>j���a���l�jm��so
f482���:�I���$y�6V�'�sa ���]���y�FW�?[��S=���\�����������~oUf�G6[�Z.ꟄϬ�~���!�����Yu*�h��r�oy�dc��0�{�tB��+ê��-Z�p�+���4�_멖���:=RW㩫D��M���X��`����#4���)$W��fg���^E��
�6��=����ً7Jv8=+r�D�T�,��K*�*Aөj����~��u���wi��B�~ 	��z�[�[`���^�@��t O����e3�u��TF/cMf��:����V�$=�9�>S�A��i�ݷ���ܳjj���I�ѓ���6�I�hK���Ƅ!
4^�^�[&Z0v0� m�����u^'㪹����Q�`�p@�L %������nn�M��:U #�C�,���]Q��Mv��23�J��[#����Z��ֿw����K���*�bQ����2�|��}�*��}�=C�y}ݯ�k���,듪f��}/�={2���@�������o�i�uE��� @�r1|;�߬wG�g���qaT��V���N��+�q�S=�9�s��[ҵ׏�6�%�|储�+�N�m����8�V�<K�uR�)�l��m�8_�3#ƞL�s��wx[^�zm'�4e���Ι�e=��Lw�]��`Sb1՜��0ػ04š_�"�b9��2�SQ����ߛ�ђ�xK����g��K�W�(�Kũ&CW��6k�b��mxV�ѸAgJ��O�ir�����_�x� �S�|�� }��˅�	�`'��N�^)�C�t�L�������׿��OѺT
�Z�#��SF�nm�1�%յhL�͉`�zt�|	�-i�E5��s2"���}���~�N$���cv�JcOyE�ED���?���$�l���8�^�p��d��`�`�T��'���?��V�v��d<�������h�[Mp�I[�}펵!����*#;,���D�"�T����'M����u!2�6���4��E��{�Gy�����I�))P�;���>�x�ڄ�)}�))aצ*/sw�0�y�3d���m��3�h��@9�t*�|�@�/k���@,(7�~_a��H�:ƺ��B��'6��ݧ�l��dz+�"��gI[��ڂ^����7N��y��c��4������B6����M]����ˁUsF���v��Ѥ�=C�ٰ0�
W����8 ��9����Eb�a54�}����s�XcqN�:�,����a�	��:�2�0����Z;77�9[�+��?E�z�P�\�
�K�5h��OV?Ǧ�]z�W!}R�+���8
1�l�������6����_�Ay1���(���+
��I9M�Q���A ���������oj<��{��lq�H)[�}�x��{ͥ���Mh߇��p��@��ZKM�Ab��a[��(�"��$F�p��nq�Z{1)�������h-��!�㞛�~v-�_�ק%W�J�C����;p#����#�(k�;�7�yYͱ�ǀPw�BU��L?Oo�m��,|}�<9Ί �"2�g_\�#P#��'�t�dEދ��p�R��0�d�����V����3���Ɍ��j���:T:vˤ�h$N�hۨ+��C�g�s�0�ҧd��Us�s����i��c�j�W��T �zx�{�j��:��0/J]xh�V���`7X��v5��*r�=���=l��bks�.�������A�c�غ�P+�1����4���C'�O<���=���1�Z�'7WS%�,ٺ�"V+lD��&�l|o���b����ԅ�I��*cx5��fj9Ep]��;:�eb�S}yK���V��۷���z�1AH-��~^���z�l߮��#Z#?�x�0H���ץH�s99�S�v�(>^�mj�<�q9��Me)_�EI��?%
��	)z��;�'��Vwb��	���t&֔�S_ͯU��k����C�iT��{����)����򾖪�o`��bX�E�zz뺤;ǌ�8T����S�0�%��B��4~){�6��H�Ń�?%�|�1JO��(�［��fkƗ^�����=��~����N!I&H ��x�U���f������O�Y�tJӃ��_*�<����� m4�D�ǟ�:5��/)K�z��n�o��'�� 6Bx�Lj�������2���6�r|�<�u������U^"���Bo����'�莆��*�0�5�Æ|L�bd	e&mz����y*iHc��4��sat�s�3���E�-;�*��k��5���,8�h��;����d�_�_�P��~���{��|�͛��Ո~�z�߽�f5�k�#���%/W���yU���1���桰c��p�d�^S,�X�i�*�{�ƣ/^
WjM
;��KTN��qq'�Y((>����g;���*�{XXC[�u���J-���%^�CB���*n`c�-�L%�����
����z�P�!�<R�-�sÈ���z��S����#H=��V����灯�m�|;�V�h��M}S<�&Xݙ��nnrI���.**��~�:C}�ϫ���?����𾝱h���?���'I��t�pn���Z�5V%�;�R�a9��l�c2���?�d	e~��/�xv��0/�~4�=P����9ߠ�$	_�
YB�<q;L��U��7��}[~��7�>-a����00'�7)�ū7���+3��6�/����7���
�M��[5�"g슀�*(ı�%<@?(п�]�m��F����Ê�W	�[�4[�`�Gn��#�󪽊M�TpM��<������O׻XvQ�𙱽m�@��Y�h��s���0�	��)�-��3��u��}�!�HN������fh��#��l��(~�rs����Eg�KTm��@��cS�7�}0��50o�#��x!eP	a�5Zb!~\k{�A�܉���3���gN��ԸmdG7Q_�
#o�ﯢ?����X� (|�#9qϬ2a����k�F���+�)(B7�����Ƀ�I>M�eS�l5�2C5$�(U��g��0�%�)x?BU,�l��/A	qҌ/
|o5�	���dg;��{�<���pn��@��9DeW�eo��ɓg�xhL�B�j&�R������4U�F��һ�߫��ՈvٗI"��>�@���b�v��u�+�<ކ-�1F�e0��}�6!�[��s�r�BfPD�Е�p������٫�nn_���!Ex�Ǳ�Ͱ,�}�ߌgeH7-�}-�&w�큃�do\<<���0��1�B�n�ub�/kh8S�z�0=�^�ڽe���n�a?Z�`<�Z�4o'&
�Sk��!����؂�lk��:�UvzNU��z`s�f�0����.��uYzz�翷�-*����!�m&�I��tj:�`�-�j
u7�g����U:�	iU��3��~E�]G��]=��־�
�TZQH_y�T�P,捌���U?�.��
��gi��t�T�MlmHEC"	�&&���N{���D�=Vs�C��Y_���v�ʫ����Pv�d���XI�z1���`q�z�g�Oمp�ทԨ>�~<�:l�:��'�F����ͬ�uM�ai\�d�S)�Dq�)8�x�`�z��<yޖ5���g���:f��	��K��V�|�{7��J�(���8���ɑ-�q�6&=���Oo?���J��I����<�j7߫x�γ�G$C���臜
(�z.}�m)��P������[� ����^ �'�(Z�P>�_���/�%zI��y����BScks��`��~۱5L�fr"��S�A�����p)���%v(hj�#��ΓWJΩ����5��h�Q%���^��B�j����W'����2zM���IUjj.d/-7�짱��i��r�(�����}�-K+!�#�z|��G��"Q����r����a���QO�L⚦�;<ѽg���-�G�N�V����S��5�+�=>ϸ��V�p܇a�R;�Lh�C�����n𺢍�] �����)_��\"�$�u��a�U�*�c�Њx�~/���W���p�Enc���{�)�0�]�]�*�������I����j	G��[�,{��K��D�����q؄��f�ø-����{�
���q�-9?�9�'�J�k�G����tj��"���ǣ;�h�~�$��a�8�?|�p7��=ڤù���|��5ح�^��ic �n�R&��P����>~�dk���g���h����(O^����4�KU��oڐ�Đ1�<?u�1h;\�O_����ԟ�GS�o"�%3�x�ˣ�I��i��~�¸��D6l��C�<�Y:)�6z-��R�v��WC�ܬ�~���Jg[�OOHS���H��5{]�x��-	���:mvUO#���u᠑!}��r�'�W��6�M��1G�7�_YH�k����M�Y+C����1�,	t�Н%ެL�6����d"o'��Xx����l�O�0ɑF_�����]�`˒����[�1��w^5t|���F�N%g7V�3n�]\����3������Õ� 
`�EC�:�BƧ<�An����EA��L�P���7�q�@k$)HKZl�&yX۽�=`����0	���XԹ��9��}�.d;�ѽV��m�2�UkZf���K=IO�����x|֐jQ��U�o�:]�Le��+��ԍ�"pe�8��:Fj�������$G?�I�8�n��V��V����[�X֛��Ӟ�"$+���%n��@�fPu[􏶈���������Gx��|s �SEH�?x	_c<�I#�P���2]�T�q~Fx<���T�øš3���{I��lً�)}��N������6��i�f��v;zU���m�,4���S_"�SF�a��ɉ�VZ�zZw�Uc��VY�aW�d�Mbn�k��F��g��Q�C�C�x�7xH��1����r*lS���e�H���w��Q�4>�2K$Xk�Ѣ��:�*����Ō���p7�����w��h�<Z��Ǭޓ'G�	-�Z�[����՘밆���Y�嘱���Ko�����v�.��=��ߧD�`,U1���X���kS����:z�7���]D�G�ߒ�R� *���;�u.�<M�S4��:.�&1�a�U�ʙ���S��I�\H�8:���U+��z�B�e,� 3�a�R�ur��1�W�1���x���O����@�J��+:tpm�3>��TWd����YA�Ax#@�1�����A���U�T�eF�ZN��|k�%Յ��YRĿ����{���F�FzL�ǥ��5�扸���W׀n�����DJ�̧��@���{+�w�r�n�%�ߥ��P!jI���U���K��6�v�{<�~ps���7���-]�`��˭�z*9��^����J1�M��õu�>OA_b{`��3YǇ�z���t�~��mU+ڡ����^�W�b��L�g��rн���b^7��w�Вp���6j��Im%��|t��IqҺ�k3B�"�
{��G����hb9K�7+}��<�GZ ���VGk����v%[���Ґ>�MS�c�[�M��bbY�Kc��E�-��h��I\U����p�N��F��BY*��;�(Hn^h�#���1�N�����3�xH����P��\�KQ3T%ImM�"
��?�!m���\փ���[dT׹}%�ߵ�!�R�Fo'q�h�#��n0�[3o��kO��c��o$�V��٣A,�t�ħ�,϶��#Bz7�%<����1�41�zZ�,��.��a��%����dK��١��I0���ς�/��&A�<^`���}]��ɬ��z��#;3�Q[g�%�B���rI�Q�?�&��H���(.>�w�5���ZAd�%K�gF���=�Ti�Y��.V���hI-�����B/w�=Rwȼ��?��E��Y7Xx��P�	PZe_Kt��D}�i����U�(D�gb�aR��A��3ި�Ɂ�&�o�������=;��v�<�L�R�%�#��mSxN��ncd�qS<q�y|!�r-�?|�
��R�BHxt�Ulʳe�3�ә��dۚ�):�ȓ�$M[��a|�ε�RL�C����˹�� �e�!�2��^�Ņͩe�]D۰0���M��?סE����W�5B!�/J�F��S[�+�-n_��x�H��Ŋ�J�^#�}�0l��Z�D�!���6�mb���#(�g��KR�z/>��G<ؖ����1 ���z�;�j|�a8s��g�m����KU�X�/Z�M�}Œ�h��P׬��Ɠ�S�A<,Ό�=	�(�&`��iCpO�@����â��<97�q���4O����CKDrqp�y��#aH�p��՞NxK�'O<�� �[x?;݈YA�p�ԇ!�\!��$8'VIN'i6(EX��&��5Ga�E��ﱘnt{k+94��#u[%�'���&X��<�a���mTZ�C� ��=����c=[o}Q�q`/I�^�#m������AE!��O^���}L��s�-2�&p�y-�q�guk�D,���qL�.�<Ѧ,�	��Y_�j��7��v̓�7T�<`Fu _�1�4֣i�5������L���+z2G$���M�9�D8ӷ%��R%:JR�k����Uy�vJ�~#�S�z����j>y5\�D]+\/��p�%��G��ݝ�	�-�v�EL��P:9˽��K

����M�`�=�FtF����AuC��vgǋa�ޗc�:l)�9�ʃ�rB5\+;~G���L��x�B�.W������k�0�?���о^<����K��5�&	���0�S�N�BY�pwwon=x���AR��Çμ�RDG΁%���]mW�*Rk�߽3�Gx1�>����w�h!T��xd�|�zM��^X)�+���w�ɯ�Ŏ1�h�p�_Q�)?;���#�K)YC��T'!70l��Sk F%Ų�Q9i��X�}�3"y�A)�8&�"q��Z�|��[X��JO҈ձ\���!��;���kg@�ˤ�l�f��¸��0�:�>���$<rZ�)	�f�Ή��W�zZ�u�\Q§���4�Ȉ�q(m9�5�����Xs�&~��U<#�Ak�� �7yѮ�e��f�VF��f�A���
�F0-:�a����@w�P5�Q_�e�O���h��9�=U�G7�5�b
g��L��,��z��c�Ԕ<yĥڷfG�ߗ�JnV����oF�ia�����_���K��*Eo�$�:T����M�ӳ_{�ɸ	������XH{�P�Q/�K��{��?:�������877�P0� ��F#��bg����Gv!�{��ޅD���AaD���k=����@�WtIˉv��X���i^8��g���l;*F�_�l�V3d��ʛ0v���.�k��P��M+�H*� ��w����TF���+`p//_������8 ѿ��_����:%<"X"�Fp�8�������3zrI�yY��<2�϶BCu�%�����!�|�%JK9�s�-&�������sd��{�0��C{$?aws@Q�1P��pD;���ߟ��<-����V7�Vy�l�wrQ�U����}�zDI�B������]E����{V���L.����G=1�AT?c�d��١�?��˥��"���c%�n����:�{d��Y)<�R��(�~�F�l�u�h�8��V���4�tl�=E,�gc���ΛgY��XX�I<�N��`�����7o߮^�k�p��G�c�#��1�AV�����G���7�"��Q��II�=x�Yc\?����<A���K�����c�i�nd�x�ך>�+Z��ٔ(����!��^eL��Z��4���1k����!����`j@�fLCX%����������~��{�P9��r�޹���߰Ė!����SON�W+�	��,9Zs3��*ˌ�^�y�ۦ���:�:PT696p�7m|.�O&�|��2W>>���v �M���D��R� [���d�� $u`a�\�Q�����3�����jp�����X����,����u6�?qo�`�q$	F�* E�%�L�η�����B���֪%$�:ޕ���f� ��mi�u�
�ޑ��nnfW�$D����>Ӵ�6�_���3ez�>H�8$c�)��qmV�Z��Su{B@4�6���RJ3��d��usV�5 X��z��R�[�!����G<~�G�/X��W��u�39�����dAU��s0Mio"�8����3/b�����t� ��3�0�ҧ���;rG�-N<�#n����\���7���~�C,�S"%ā���?���ca"�ÿ!x���1(��<壖yC*��C�M[��ΫZfk�����<�r4A3�������7��F% ����ِ��3�r� ��R�����;�Ϡی@��o�-�}��5#�_<���O�}����������Ⱥ��}A�(�vk�n����<�Iu��,j.�J����L��z� �~~ޘ2_�VXq�o+��\�MW9&,�Ƙ�ƿ}@[p@��mZ+�a��xL���ѡٶ>�]T/ʯ~�uz�Z�}�����g��!��I�
���B醜{v'�s'��A��q!�-f���X��&S>r�Ћ�X���j��2���PR�`�-�5�9�*�";���y�c�����<�Hۓ����D�j����&/�O��Hc�7i0'́vCߐ��B���4���v�.M�j��i/�-K�B�����
�<��Cn4"�s��m�~ ����\����?�Ok����+��S��T��� ��^3R@
������Vi�I���8T��_dg���x~>�hJ!�^�~]6�K�=���*��]L��F�}��5mO錴����h��=r�C��պp?��_���oH��2s����on�)�b=��S�|o޽��v��A=��a�3�`0�̋�_��h������Q�}Rz<G(�����16�h�aȒ�\e��p���>R<<w�k�]�8xD�s@B�G����V�mh^��{��6���#�Z����H����DSt�ƾ^����I�iӠ<Ƙ���GV�VFcr�l��qm��{���6=h�Ur:'�U���/�9����[4���LU&'�d��+˳Y#z6y��^�':����{dF�`�I,�~�?�$N}�04����?�H�J����1j>�?�;q�T�iF"*c<R�+Oާb����J�T;��(>�[�6�0`n�[eA(;��SՎ�X�U�ˎ)67���O��~Ɵ� �����9<n�4�&�A9(��E��Z9�x�������]ܧ��R{�,�&��z��q#�b���A�ԗ��h<̽x~�>]~����� @I��+lp�w��!����:�����c�]��l�����#�P)�x�N�$��J��4=ʹ��t�
?�U�z�d���L���2%���7�9�r��ߦ��kt��,�D	�]�H"G�P<J/df��(k�A�CA�W�|y���k��Dq\��Bk�Sd�A��8���!1/�=�1����6�]YVOd��I��"��r]2z���HXce��[�n-y���g����M�뻪�Bv��9�K6z��d��{	,��ڗ���3e�u6�E2W��NcTQ��&��'J��{^�����k�Ë����Vz�������=�#*bF�Z~�Ġ:�!�;����{�]�,����O�߿[3џ#���詍4_��H�#�m�R�T���n�OK3
°�Tg���b/��Mm�<ސnR�Qa�l"�XX��Mg5|z^s's�93?h�g�{�lIM	�rd��U�~��?ň��Ե�/�^�nDk�`���T;��∐/��������nt��Q
:���v�w\�3���)*Ԭ�}��{�W�$1�)$��b�Z�\���lc\�ZFnΛrA���Ȫ��[��2f��O�>����J>�m^�R������m]�E*�S6�kmȇ�2�Á���ټ���"�W@p�D�6ڤ�l �1���_|�5�X�{R,"�k;D����=��,�H<x���O����}v��THQ}7�i>tR��T��l�~(�j3�NzuqGM�Iy���l{
�N�ysǸ�J�>�x@�6/>���HւƆ��+}]d�o#�Ywy�ҲG�Bs��WkI����n�_���@�GRe6���9����"=s�v�i�r�5��A�h���k�S*>$�&LĔ�n�کn�P�\��Y�SZ�Ţ�����.�+)�23�t�����(7�8������O?�_?+��M���`f=!(�[��Ys_I��DY� fp�����4�"�9 ��L��pm�i��o6YJ7^2H�� �@���]�<E�34�2��:��$����q,�|� �Y��/����f�G���dS�IcX�7T�8�c�4	�-m/^��}���!+�h�3�q��p%B'�!�K��"�ĵ��7{����տH؁�"Kƃ�S�JY#�@�m^n@(;��e�<DH��Z�r���y�U��Ӈ3"�~�a��M5��kVJ��\�_�U�[���6�OR
�=;;�+�7�=���z#xj�Ԯ�R��!'�2΢̘����p-�����܇��>NN�]���De	-�Bi���6&�/__3ꩮ�j�M˥���-Wn/��^e�H}xG\��~���f���^�y�i���>�UDj���|d�#��uO���A��>�Qܟ�l%=��(����0ZFU����/�J!��g+���B����kX�p㹹��m��b��4��ī�p�����xnѷ��-�4��;����OB\nH�@�g[��d���~����:e��S�̹����!�A-ڷ��� �fveo�3ek��z's��3��)�JZ��ޖ��<�We�,�7ia����{Nՠ�7�/����'��M�i�4�U	v�!� �����x|H����8o7�k}�s�kԅ�'�v���� �C���\�gi���24�pq���7)Kکv�w����{B�����-��s�n�s�b1"�b�F*r�A���ިI��;6�M��@�Nϙ�:����ʘ�.2\�P�| 5�"�4j9�2�T�n
GY���mW�YAH)լ�n�	�I�,�}t�*�;��M�����{j������{�π&�N������q�O��12����=B�x�0�Tσ��^�0}�=jvl$�{=:>%��{]e��Sl�l0]S��k�����fecY�����61Q7i>�0H5�p���QRٱ��!���4���-�6����?�4�ޮk=L��sBi����.ޫ'��9�NM��c���{T�x�!�Y2֭�E��Ԟ����6�¥t2�>�}�{��r3��q����QS|(t]�R56b0��k�w���$����46��$x�"��0������@�ߜ�=��Y��"�DT�x�x���V�̦�S�9�
������z~�3�JPl���s�& #�N�(����;�N�h�Zr]�[M �ϻ>�(�;�}�V���w�:(�bL�ʙ��u"thăA�Yd����Ԕ�վ�'������4\�ƹ=_����n1Nd���6�&v��.x��&6�9�/փ�Z|���f����7kP���^���F#E8W��4��/C)����@�`&��������^�F$��L0��L����I�n��O�Z�T�]^�[n������7d��,�7���=�{	�&2�����ʩ�6x�P+ݤ;���8,4߼}0	g�sE����d|�v'M���m� �Pj�Y�Z�)������T�_�q�";��O8�"�����[[�����i��GA���*�g���n9�{�� �03 n��������c������{>���ށ4UH�(]�d�.� ���i�L�Q'���9ڃ�Mdf󼨣ΠlФdX� ���k�nx-}H�q� ��,�2�c��ڌ������.J���hl����7G3�xed�k��x�i������@�f���gE���1�GF*l��S��x힟��xT �Q�E�ꪂGTm�4aG
�ǟ�Ok�#�c��Ypx�k���W/��,ܦ&h��^7ҫ�)������/����Ӱ�&6��}Nv����f�Ζpwv�d ��Br����K~��G�Ƈ���W�E�����H<��e��f�i4>����);����c���Ư^
��E��E���i?������J�����	_��%f�[�_gg�tI	��#�;4�( �lo��25G��~������x-�.R2z��F� p�#��,��^�qP �?���7>{�|%jE+�L�"��F4�~�k��y�'#c�y����׏�bK����F9N2�9(	���)�j��p'�P��\z��J�\m�,<�CX�<�[>>�bz�C������v�W�� ~��.�lnY�x����_D����W�رP5��+l�H����M��q,f��,�ܑ[vV�WX��Q���  ��IDAT�j\A��4�އ���Ɋ�e��N*�^�:SL(���%�C�����놎 �n����Q���b�g����(-���Y�?c@۰!�S���������*�����t�qܬ��2ޛ�A�t��=�Y8��Iy�RX�2� ֖��G��#�����Z��<�>��sj�FB�Q�acX���5#��6L����Z:IUT(�x�Y;uW0q�l2�a�9�X��0ݒ�~�b������B�lKX۸gw��b�G��w���� ;�z!%�=28崊�[&2���H^��?��u��y�?�?��7�H�\��d�X@rd܉�*�q��2Iź&C��S�t5��s���ٵ�iP�'�n�M�A�9��dx���t&�]�`d��F�nr��Rg���� ��iP�"�̬йMdȝ��b�b1ὁC&(��S7�pQɢL,��nt-�hL1}�A����_)KJ8I�Y���yfv��o�	���@�>�6�cV�ҩL�'*��k��d��ë�laa�y�QC3Ts��p���娍'�	B�iʱ#��+@̀k�C�R��ɕ:�'���޺q�+���& J�	D�=�,{^+�=�����5�=��j2Ξ�R+~����-2���JG�F:<`�<��������{˹X��:���x�JSA�w�6�̾�h���ޮ���@�0�A���y� �HX���x��l���2[4�}��^�W�f#G�f"�L�ȶ0A"����IO�� Ð��!�H>&�S#<AK�.	��iq��=��zʳ{�Ѝ�\OW�)\��V�r�י�e�����]e�I%q>^�,����r���A$|wB�����h '�cR\�  {J�ܼ޺�<a���%���鋛|7�%>˕�Xt�Jd���үsP�:|5L���@�cd�S�)v�{�`H�Sj>�3}�Դ�_����}i�IT����	��@�>�lO|��͛7�0�� (�I\Vttt�)�u��pREBJU,#��9
:yQ�H��	i��yI�f�,��f\�\0�1���I���=��׍���w�Z2��������_��:�D9��%��c��0[��X,1�����x悢�����cU�^��2\�r���=O��Ll^�N"���fʦo�����̠�{�f�� |�7�s�P�IN�fu�E��̓<fUT�G;/�E�q-ll�����G��Á����o�M����ʾE��k�T���������3X�TwyEC黪p��V�)��1������N%;��B����	l�H�T=Mq����L��u!�y�:���<4��9Kݍ:��蒖EEE�~��E*���I���+PR`.t�q@0�d�J\ǀ:��̦���r��55�bZG�����ΨF��/���#< �����4�JƲ�.�-�Pd���Ȯ^3�wo)t�
 &� F�X*�Fd��׬�L.AZ/Q�u6P`��N)v����sZ-��c�m\����-���9�2L�qe�&�A#���ƳUH`�3�S���F�Ȓ�5<P�ny��L���n��_��:F����H�@6�7o�C�m@Ev���� �Uȧh<t���2j�s:��u�|МT&S�,g($*Ӄ#����.��p<���xh���<e���o�7VM���k5*�����!���5�����1���L�����Xz���61'O��_�;���S���̮&��N�^��@��$p�)�inZ����?//��9G6��	CZ9��������kje��0h�5f�Kn�]\������eE�4/^�����8U�4��ct��5�i���|����=��̑m>�'��=Ć��).R� C��Uû����pi����-ltE�Ҹ�!;�|P^�麉�E��8<��� �v��y?@� �TI�˒S�*5�Tv�+�M�
�q���^Җ:e��v�ll�f9��8�{�#�s�y�6]t��i���9�wg1�j���e�of6V��b�����!�1y��������D�C�v~����;���ohrML�L�%��G�<������/)?���z���l��'vr����sv�c̎��`=�u��0����qD�;Fs*+���ދ�CW�I������{ �Un1^�Y4Ҟ%4����vIw�s�q�l߃$i��TT��1�����%��U0mzBei�W���]���Y �򣒃�Y�t��TA���e�Y�,�m��9ƣ���v����9�#Q�pOO��>�^�R*O���i <7��.�Z�#���u���?�����G�Z��y��D���n�AN\��B�_<Oo��u��������)3u��~<t����pٜU�^B����[�.#�B�v���-7@:}^�����ݞ��δ�|&tXq���g]����5�.��΢��}���C܊�n�܈T�B��y*�����8��2=iNW����=x�?���v���R�|�EzM@ ����N������t#͎ME{LZZ׊�n�!@�ݰ��n�W/"���a���^��'��=�=9-G��$��)��,��|i����(�p��_��)l��Ie�N׌G��1="����dS\Ĩ@�H��o����߱�T�Wѐ+�C'?��0�������῀Q �J,]�"Z�/Q1`�R�!� ~H�gڮ�磃�/S�������{���δ����n6iO�QX��>'z�u��@270�} �C�$����(U&�Aa�G���$�c��͌4��m=OD��*���S� d" ���¥���w�}�"n"�Nx�?���j�[6�v�������ᵂ�h -(P2ƍ������1�mf�Sz[�.3�As�4�2��ͨ t�XB�0]� �d�;�ht�� W�?с��N�J���K�A�seQ,��k}��!��\x�UX/�ی@��mN�%�[q�Dr�{�(��D�?����T��D��ξK��<�!���ᷱ>�p��e]�U���ݻx��9���md�w�M$:^\_�}�bx6��ț������F���Z�>��;q��q>�]_3�ب�z)2�g��l�7�B�'M�6zf�gcȄ����DD�14W�BS���1M	FҴ���e8���
� ׆����g-Ł���5��H|��E��gbq�O�Y��/g��J�ַ�`
�����ũ@��j�E��:����j��l�4��倬I���g�	�IX��'66&2�m������{A�;,�v��
�������'M3�i��ٙ��(�PN�T�	�l�4��͛M,�ql�M�>pj�̃����5�.9�&p���΋� n�QV.�m��O�w�]R��{bgL9���[�ݖh�LC��������Le��0]_�aNp��
/����i�f�e�g,��4޻�nyz�z	�*��%�2siJzu�u��^S�ȸ�G���IB�$U�%�3.x����=�)Ԡ{�aX���0\�j�{�iQ	�w٬��w��~���Zd����oޕ�ݻ8���Տ�K?�����0�ǚ$��u���U��.eV��^=�3��5����<���:�������t%��J�ٛ$�8��,����s���Q��YKa����H����VR���5�<}�0�$�yw��7>�����O�0Dn��X��,nT(k<����rgӘƬ�4�_��MsS�,����ѿp����o�$bI��4#��.�PV�>�CZD�h����t��l�޽{_ǎt���6[�"�_��3�!�'F\��<FF�&��.���Pe����`m<�O�M(��g}V�dWz�ᘐ��\�l��t!C+X��/}�˹�"�w֜�P��4����Am��f�v�G���57���5��x�,�3=f�Z����+ �\7��þ>�g�lL�`l��P4����?����6�LLn�9�N�1"�$�� ��K0;�-F���x �	���0�9��M�C��a�A@CdȌAg������r�vڧ��d�K�䢝1��"�dr��؇�ˬ��Ԇ�BR�W�0���^l�����x�
ѕ��v�	�,�#\��q�A����4�)s�w�}�����F�q��"��v�������^������*��Β� �B8����E�e8�q@ ~��u����ct:�'~� �����s��N���!�Í��{k Mw ͕�@��cd�n�-�r������u�
���8;�8cB&�{z%2��I���Gn�x�:^�מ�ާ���E��Ѹ����3�������x�$V'���y��c-�Z�.����Q��6+����7�>$���웛8�Lg�'-�;}�%��K�S}ςr�"���J���Sx��]|�]��P����)�KxP�`�����p�1u��l���O�
��1��%G�<�5мz�����&^� ;;{��=�"ϟ��fS1�9o���Y@���˸��a7��rl�4U��O��ʊ@��e��C4./�Ĩ�y� �iۦZ��w<S�٧2�Hz6��Jj�:#�z:���{����G<~1����gU�J��y����
�>3T�j�,��z؛�Ƚ�=.ǘ�0�cVOu���Cuֱ��ٜy�5#�Uٔ�8�)Y��9]R�L����|�4�UB\t���)q�C�a�QUʧ���S�¨�}r�X�ȷ�>�@�j���P�H�T�4vh�PH5�Qj�1)>��JF���r�,Kds��4����bZ�N��(�;,M��< 7�m�I%d~��_�o��Ɯ��<�\��Z�����l��Ag3�)�h}����aVs
;��Q�T�C��Qg?���^r�
�P�B@o�9�Pv�!%~��C����I�C�ּg��z�hT^Z��$����&���@w��8(X(�;���7$v�*�%�sY�eLU�M�n/�_�u��E�k��pS*�(����~N���(���^��H����繦=y�l;�5t�ٜ˘�n7J�S�i�ɥB��|>�<��Ct�7����C��4[J�y¿��㫤� (��a[l64�Ѩs��9dN7���?r��ɖ�"[ec�PKב�K_��(bQ�ݦ\0�J)�I�L�����NA�pCe��y�'����%;5J&�8��ѭ0K=�Z�ob[E��P��(�����)�C�7|(٫�dj�t�.v�5�j=�c�_�j|~���ˀ{yO��30�[�ۮU�^>�PKD�/����eo���/��O6� � �x-�����B�_\c)m�4�Nj�D��իxo_}�yK���Z��rj-�/m\�B���F��1/u�iW����l��2xnwヰ���ݨu���FP)K3]�(�euQ�b��"�ʱԁ��,��8�zS�W��(�>��oo�z:��0yϢ��=d��L�ޏJ��0��[��F���DU�����������<[��&�%X&��s�Hm�՛�R� ����f-����#��w�%�mf����`p����F��w��3�m��/6b>��_�Fq����i�,\�r�
m����9�{c#+]εy�����K�P������s�A).�exaFCO��9;�x0�1�8�F7���szeE�#�l�q��Z�J�1wn�����M`�+\�S.i��k�G���������#���U�ڂ.�GIl׎a̦��+t�] �0�I0 ���d��	RB/Ѵ�B-�!��Ϯ�gt�c=?�:�������X�Vv�o�^{!�8Yf�H�'L൙�r�`Ȯ\���L�}�w�s�Ჾ&��zB�0�e��ե6�t�XQ��H�N�aB��%�Y���s�{�`�T܋���1�\��>J?o��g��_��j��ZB�\�i��{U����Ѽa��>�{�1�'4�g���|N;$�2>gdU�s.Ve`#��2c%�Z��a�%��\S�����7��ￏ1�(�r�[3�_46y
��4}]0B���>=A���ӳ�s-�Z���3�N�����aހπ{��@6�+��/�uV��R6p(��]������|?��2�*��ޠ�,���3�G��of��~U��IHA7��}���bd�'�X��(��p�;+�>iu5(��fD�7]����m��Qy3����=�������c/K
VU'x~�x�'f����嬩�;5˶�����G�:{�9���O�t0+����l��Q)��1
���t�q��G��s�N�S�A��B��%2f^@c[�3jk������F�P��e���{��{��QSh�X�����{������2�~e UF�~�ϊF���SV��HB�a��H|B��ף���a��R��1��w��t��m�T��S�ĝK��(�������RBͱ_B�B:5A���Ҙ�&7!o0��}N����Q�\��#����GuB�Pلr�E�g��%�C��8�B�s9�ij%�&~?��͔�c����z�b�Pe�<�<��TY�L������3&8��H4G�Sږ��Ĭmּ"��S_����1�|^|E��cx�yFv�q�w�cq�[R|��,� ��A�eZ�3*��hpr� X����c��=�mTmc%�p�5���������x�8\��#��# ߼�5qWvp�:��`�%#�J:��#.H� _(��a�e�{䁊;5��_v0D�nB�}��(w�=fۣ�ݔ�{r~����8\pPڐ�b��<i���X>N�\e9cpUCx+����9�me(�Q�p�;��t��:�u�r�ZV����c]&-��ԾϿ�1~.��#���l����A8-Ё�ۘ'�7SNs!?��%g:��s}J0���tȠ��6[�����R�TJ�����1/(�VU��S6d�
쫗H�-��d�I�8M(Qʳj����1nX-h,��1,�y�*0·�徳����o�#��]�FaZqO�H�����W)�c�������r�#tE���MP�ύ;�y�ҁJ��Ԕ�݆��5`v��4������T�и���$4�n�v��/Bݑ�q��UUZ���b�ڼ�ݜ\J��&��=�x�<:����x�~�ז�����LX�g�ꐥT�7�԰.�׽gO4�&Py��Ô��N=���}b��	�����nH�C&VE���z�׳��OB?�G:@� ?iƔa�pӇ���ZL��� ��*@e_A��TL�F)7e�T�'�NQ}!	��W�������8��"�MiL-��1�tQ������˥�UFZ��O�!��kd����b����垀�nwN�;�]��_���]d����*>
�r�\5���V��� ?H�N\�F�z;6�塵�(�l(�σ#�Hi�6E���-��-�#>o�q� �	v�E(G@�w��&�,j�=i�Tjꮃ3wf��m�%�NM0�����|%�p/��qp��%�������e�Ǎf����
)c�P 9P��js�Q�)j��%�S4q�ި��8���j��8d<6`眗��
�>�A�n�ڇ`Vȋ���L�m����&��7(OXs���(#?�����\p6M�A2�J������r�=wG��!�]�b2�� ޳M?��>W�XBi���Y�L� ��x09�0C�DNgһ�����!�7~�Y|с�=�=�,y9�2
*$9�!]�S����:�szC@bK��W�qV�H��
-��B���pdF��w�	�����k�ee�/��RO�y��V�:����x���M�bFK.�%7N8���� �XZ��0TR5���{m�Pf��?u�!p��"@�{�K�P�����h]q�,a#����3Iܱˎ:��o�(v��ZP6��j�b�4���0>�B���Xz�(n(�3#�n�����@66)l�'�����rB/jf�MCI���0\�Ѻ��t|I,�jQx�5�L��Z�u{I��t9�D~����t�4]�q����[v;�!e�Y׉6�8o���3)a&�#��_J�����=6����q���i"�i;^���]�3�����Urͮ�����CE$u
Kxm!j���BH�א���$�e{��i���ʄ���
a��;V7���J|�~��E}�/S�ZN$���E�Z�h�^s���>隆��8��o_
���h�$>ϗL���	5�X��p�J���Ѡ��-e1d �D��|�2�0���!�	�Y*ۘ��r4��BX�G��?_�_����E��!�3�<S��?�zU��(?��Ͻ	��P�!L�"�gGXM,���u���Ը����� r��������(s��zf�t&h_#8t=e��m�OFz_��D����W�	��F�Pcj�G~1���7�ƃ֤*#���r\��?��)1�]u��1ѝ�N\>��|ݲ�ܘrhc�b�Y��S��@��iN�I��	q�"31�]`uU)V��#������c�}�˄Y3�N�΂�#v��B�?����Db� (:Ճ�E�\L.�&0$�w�%-'6��jz�]�%e���+ߚ�C±�6��-�um�罕)�������<WM��x���3A
��eɑ!�B:O՗8̱gK�y��)�%���%wG�������|bZr�3м����%ٔ�Bt+E���qX��F��Ŝ۴��B
�c(��7"c;�?��z���Q�韙�t���mb�������������O���Wm[�j%��0�gR�m�M�X]��42«��
��>�9~�r��N�:�����������x8�Āc���Tp!�g+�rB�%�w�l��R��R:�BL��a��U�O���Lل�Bi�Lk/���O�!Fq	tIg�����MY"5Jc�����]��a��廏�1���ȶ1Y�-HP>�j�I
ZM���4�5t%�w}O�AI��ˠ��4�1��i��ω�{<�
�,)�<��b���+]�$Ss��l�Z��^�� �i�a���a���.q�U�8	 �x����Շ�,����ZJ�7q`��J���(�փ��o�%���{�@N�T$7�������|^�y!;�6&/9a��p������ns��BQVGu����g��Z�/П���S�|��l�'��Ǽ�Y́o��[�9$CdFzmc��,�MdtpQ���sm /������s*��De��!�x2?[��Q����_԰����됐��]W�J9���Va�s����g��8Qj\�
M��W?����bX�ǂ���#�ۧC��uh$�/�{h���]��54�Y����9!�g��.0�^N��
��E&wr��%���l<���ku�=�)�;��.Sy�J�<CC4�,�9����ơZ����C�ČRC�vG3����c�[�şqoBEt���A�b����p
Afe!Ǣk�(7,��تa�3��Rg�[���Dȧw(��w�N��͕�^k]!�ڿ�� ��!(����:�`#f��}�ǚ�ʏ�gE�J��,�7�����m�݄�������y�0|�V|`������)ب\���x}��K���Z�c�Q��"�#�;񍱗<`��{�HkR�_yt��/�t�G��5�Yا�x���췴8I_,]���r��$U��L3Z���F�;NSv�q!�Q�l�����Y͟j����E�,E���D������˿�K���')*J�6�lO������&X�y� �GC	c��o��>�(`��؜1�qsT�rLuFˋĩl����)�܃�sQ��}����bea։�첝��v�� 6�~a�8r����r��F��������-�{����x�F$�`{��{|�>4��&O�"{��)ǛZ�.�{ġ ؘ4{�!lp��gNk���oU�k��I�KWK���tY�� `�����n�"�k��Q�{ś����x
fs�oD�ǃ㖗�4¸�g��P�օ��C�	�����z#�\մ��g:��{�]^��#���a���5Fx�i�Q�u��z���ě#�jz�{8<� �դTX���cr�}@_�3@
��Р�ܢ�J/��2qH縠b����}p����}5_����	��<�Z����MYr�D�/��Gi���EnB��3V�b??>xdk/�'��\���V~�8�D�Y�����p4���������% k�S7y��d9.�6@j �F�T5�O�� e����Mt���Q�Ar\l4�ؔ�pѱ�
���AM��0 �ѭ��(���mw[���V�O��	|Q�f�tq8�\zPM�\�WHk��i����N�6��ME6�k�.?6�[�s`����׈�͑�!��B����.�~�B�4��R���D-�J17�"�N�܉[������q�w��ۻ��N8H���=�|j m�|���:�_��9������ب�7F*,��ڢ ��{$
8t.�SAv�A��m��� �ݚ���eɃ߭��{v�L�0a�X����N6á�i9���1���"��Qm��^r���������k�~%�T,��7`��#�l������������s.i�]R$fO`�~���8xZ�:��U Ŭs�z���K�!���6��ޏ����o�G���F�/Α��+�ÿ�¤��m�t�V��}ē�r��`t��,�3;�$���D��ɕ��(SW� ��]WUD�J�E�O��|j���I�<��Cᢌ��Ǹ�^	Q<z�عJS��D��7�؂���wmv��.�ki���8ib%�<n�W��p���3i�i��j��s2cVaw|���|�����ׯ����C��;"-�u�k�Om�$�c*P����&����	�x�`��P𡑶�MvU	5^�W|�m)�����Q�L�g��G��*����y�؊�X!���4�{漮��!��/�7:\Nɚ���.tB)�<��멼}����w�����a��c���Dbw����\G�8��#(i�d��s�R6n�U�M���ʳd���s��Z�S�EG�~����H/��-{��koL����#7��}c����7j�I_M��f͝���p'i���#��K���E~�ˋ70o�N��3����� �}�@�m��S|w �"ri?�ޱ��4̼��:qxi*ۺ�Fe��x+z�e�u��R�}��yMR�8Иa��M}iT,6�%�sNvE�2�3��XI�JM��q�kz�~r��9,���I�:��33}ln4�����T����TM�cvq�5�	O��bTg?~N�Lx^d�}牭�ܤx1>�����p[L�Z���$�s��e6�U��7f9��q��Q7DL`ϟ���[� ��g���5��E#�Xg����r�Gq������2{<��h(��7�_�M֢�g��rZh<���Z��٘��5�zU�3�N#��X��Y�ƕn�JKW���BW��o��/�F���v�L�Z��_f���k����=8[1�[$�V�ܦ�	$KI�l�#4��P�ؽ(;�]ՉO1˽\�z�N)M,���C$��')���0�қ�t���4�c�C��M�F��1ƣ����AP��*Ӈ���T���ث�H����ϟT��i��[>٘}��y��,�/�G�	����w��֔G�g��P�������4[��AAC�a#f3!Lg
�R����do�]��Q�G_�&�d$�q+��Xw'݃�$�08�s5Pњ���D�E�7 �M}x�>>�|t�#K���DI�uWk��H��`7��S/Ϛ,̹�b�&���k�T���P���)���ߧ�?��Pi��W�ք)
gOzX����k_�KӨ=-$�ϵ82e���n	pM8��`A7�iߌ4��:�=��C6{��)�L ��߻�@�C"t��!�.�PCo������!ƢT6� �_6-�L���4;�CU�d ŉ��<�v;�9{ub��)O�HIk���"�C�,ߦʁc���y������e�N	)D��4<�@J��8�Q�z�����r�V?o���n��?�ø����(h�`,	>K��2(2P��� F~�N�i����+LR�B_��L�75ɳ��6�L=�����C���O)����N���U)���C����$�^�xx �4d���(G�pFGF�@
���f�C�Ӝ�p���u�R���eP��yJ�y�do�)�ǰ�[����^�Q.A��n�`�R��X�R�B���F�z�gk7��������E�Ǫ�������f@�����s�׿�i��瑀��ϣ`:r�H�&�A���.�=t�'1�ݡ�N�T	���i���jrժ\j�4���Q��Ժ��!����U�:�*�0��G�Z���9$v�2�)�5��u~�)�G����G��b0��iɧ�0'�R�ύd���F��9{"[��%3�&ѢM������ba��&�13dΌYRX�%�����2�X4C���8��1���:�����^~��+�Q��.�bq^�H��"1�����Y�Y��_~�K����ğA	�m��e��D�F�&3��b��K���pֺ����ׁ��L�`<ݥ�;�Q���LK!OtLΤ����)),-���3L�w"-�n�5�����f�SP���gKS�ݞ��+��9y��bc���=�/iE��Lb�jB�0<I�c��)5�x�����C�͖ţL�E��w�ςA�Q8��
��_eé Cu�L���f�v���A�l��;�4����0�9J��ի7���]��v��Y\9�Fօ�&B��#;�χB�ar��`�$hʎOnz�y6����)�yl��oX�WVF�͹�20	"ͅb�ɩ�.���^�����id�S&���5��At��������С)u]�58�<���i�����������ߟ�)�쥧tiB8V�h)KC	*�d�E�Zӣ�[�պ�*쀅��>6�Q��(7���L(}4���#�z����nD���	�}�"�T xo�X<�`/�%��*��({�u�(�9K����!Eg;LN6I���=��'e�������f����qU�%��@K��UD=[���w�&~��jr(�F�$B��(3r[ٍy=��j�209�6��t���nw�TI�,oa��`G?P������3�M0����=F����Q��̨ܔu6ۇ��p`�2iO{�%#`T�Q0$� �eA�+h�Bh��e�}��jK8(�,�<M	�:����F�HpY�1Cޕo��:G��w�:2	[��.�4���}��hw7U���,��'2�o
Z�R���=�t��Ǣ|����o �g0�M⢥\�@6�`�W�:e�i` \�"-��H�V���u#����Pv�K�T�Ð�Sz��E�C&�Ax��A�1(Rab�����Z�bEc���6�u�;̞�]ދy�O�(�H�q!Q��.�ٻ��#(>�{�.)��N�-���m�I�jfaC���cf�n�~fj��cc­�.�q����3�7}���Ӡ��H�91Zl<6�ٓ��o������2�,G�ɩ��a�X3��6��z���	�ݚ8���M�떪�G?K�1�q� �ߨ)�,��}`�E��r��Ma�?GJ�T�M,g�{$*c�w%I�����HI��1u\�#G3���ڬsG��>�~�f:��2O9t�Q�,T����˹�#Q�E��[�\ީ�|*��KdȋꦮƠE���o��{笌�J��L�B|i���xz%��_+9�7��N3v�6�°d$��W��ZA���6Ҕ��3h�@jl՚�O�@y4�%3RP�`�L5ԟ�ׂ��SZ��ցy�]P�"���e<�}�����8x�_�|Y^~�R�Y}�YF*h�����S�zr�J�����^H�5��\P��{Һƫƚ��:�F��6j��s��{;�.�x��:"x)�O��tH;1��aq����k&���&��{i��4¸-�)��R���������೸��LG+��(U�8Q!��I��ԽF`�D�&�B`��,hj�q<hz�e����{��̢�s�3�Ѹ�T����*��$n��YM>�Uͺ}�0k'�*]qM�M�����9f�Ul�6-8��%OA[�^��e$>�yrQҲ����6�9�i3z��$~S���?���ˀ�{}�T�F4}��:�r~�E���/��긶/C5%��>�)��4��a�;~n�"���Q���gb���X���dUyp���M�yH[��a@��`�pD0M��ha��~�L�$���\�7oh�w9�=`��nG�~�\<72��*��d�4��t�s���l��xz�vI�����S;ez�k�ZZՅ���U����&` Wu�4 ��d��^�L��;�GSi8#Y�OY��qh� �
&�w�ְ���Q���@���'�V�P��"e���ɝ���.S�}��S$�i_���ma���<��e���I�gM5�����q�OfdC��ݣ@�<
���8��+��6��PP@�M�����J&��(�Ϝ����A;~Gzx㎜gE��E-��;7�5��s��9X!���`���Њ���P���Xe��	t^�~��`\�(?`ܣHf�J��������@M�&���(��%f��c�T�\�_���i��$��|J��b+2eO�R׼tT�	�1&x����t�� ���E�.�Y0���X����1�;.~�O�I��1�tC&�����3@*?<�����a�N����E�n#J��6!��jp��5a�!e��еi���:����2mU�����X����в�E�_��h��uF���_}c��f��ݻ�A��{��dp���Wk�r4$�~n�z	���.4�E���L,0K2�pVc�u�~�������}#����z�02&�߽KF �iQ+A���.���y��9���� i�}���O�l��oބj�Y���e�/�����|�T�cT3��ٷ���'�9��:u��\oBz-^~3����ԭ��V��k�I"�^��HT=9C��$��jBWnA[��y��:��nX���]����Q����/=W�>8�h��yW�y>/<F�����������)�Kk�r2jb�������*6_y�5x�M� ��e�jM{5��䘾�-߮����F͎��4N����zc׭��.��{�9G0%�T���/�L4��	����N9.�A4n�h/Tނ Η%J��Z]�8��C$���T.;ϙ��O�cf�X�W�eq�s�l���I�;�	�M��:[����{�����~-0�x��AP�j]�_��}͊������s��gr
��RC�1�(�ޒ�d������k�]sR�T-�u*���!�C���zf��ob���Q����&v�����Y��~�J���V��ր�xV��l�O�p��l���`
��hT��I�!p�B�|=����ൢ�h�?��<`'8��/�������
=��<�-x �O,�dӗ�ɣG�)�W�P2]R�Ŧy��yHG��O����!9D���"��T��ap����t�_�P���´q)�,���,U" ��^���S5F�dH��{��b��^W�ѶYlĢyN�)������b	5>���cӓ�ڟ	�G�6�\�	���b���<,�ƴ��]J�d�E�>2?�/&�#��	���e⡎-n ������D�v�n��X�c�N|?�8�����Nޘ>z	�v\�
��;�krΠ��vѥFP��B�rXb���C6"*��K�6O�5��*��ꌶ&"K��gͤ!.��F�-���8U^>{I�����0y/�w`����3���my*��k��yX�.��U]$L����hY�y�$��1��4���b������ߝi�����%�Fa��o����B۟42��9��>�kd�5�	��2�sJ�Sp	튏����VyE��(cܰ�M��(�Ү��(�������KR�ĩšV���N�l��9�����kD��ֿ��`̭�4d1����#��\f��M�8��Q陮
��93�(�������lr�%H������<�.��?tE�8�}��i���icȦeD���̹�~��ۯ�����^d���u�tW����5�h[��U���`� ����St�O������oٵ7vbɰ(���$ۄ`�Y� �eh^�'�޳��;n>6~N5��l`a�ൠ�ƅ����p���8ت_0��y+��bd��u�F��Nh�(Wy�E�-nt��iקf�x��6T:Dm��Fd�oww!��q�q-��Π��}A����OGL/�YDq2�<l��޼~CK@2��~�Ҙ�Q��W?{٤@ ��N���SX5��"34_e7P)�}��Uu��M�z�Aݰ$�n��ǎt��anbm�����gF���;���{�+d�����ee�9	�1� N�6ȅ��&��	�����#�:���`��N�L��X�//Od�p���3�C�0�:<�<h3��$=�7��x�K�q�{=���u��D�	�~H7�οW(%a�c/�ى�D4��-c=��N����0����cݜ/WI����e����9.��\��`��|g� �1�X��Q���}5^����k�\�'�Q: z�4�!ι �ǽ�y�ۃ83w�RG��P���^<_nt`}݇Q���$�j���'(�1+H��1:zs��G�5�y.[�M����T��� ںe�@q����c@��M�8k��J��l�3��D�i�i4���%���[xM=������\Ap�a|��2��=�lU��?G{�z ��7�Kғplnh}������%�B�l��ETdڵ�3'����q -���^oQ��t ������S�/�X+Qr2���`}Y]��bH�х��D�sC�9��Cڽ.��O�������7�+�â��/hj��b׷��NՃ��.J��m�"�/�||�]D1�ؘ}$a�,S�lOlP�̃�`���;b��m%4(j�у�%�v�	�x�{k�q�1Lu3�&x��m:�?�~8����_�"���OJ�{O�I�,�A��뱔a�k��|J2N�	L`l���sK��,��"�h��?���6�q�I)=n�w��@��2�#f1�s��4����*�?�O����\���m�gԔ�^��|�ds��U~J>���]�6��zrm��}(��Y�s[�-�4��U�^6�4;8lhA8�\޼}�Q{��7�|�	�'���L���GtP�M��/��|�k5}#������HsJ�а#l�o2R�Z�!������t���
��dD�M��N��2#��%O�c���ۓ �1�ۻ;f��#I�XS(ɷ��H�`�lKgc�c�nY��
(�?��� ��`���t?���#E������w�>�Y[��$Ɩ���S����*N�}.j��T��}�q���e�g��pRj =�S�@쒝�eI�'�e�s��2�T<��$v�]= �������z8��[v�C�+�DP��DgTƋ{eU�M����	�Nn���|t���PZcg=m�I8f�Ј$6obn8��}^[[b�o�8#0e��+
�Pg�R'���;(w�)�<^�;4��0��2&��ÔX�	f+���N4�1^�?�&Cʦl#OluLS�=Ԇ��Y$xR����q�)@�_�I|ɒ9���;�� �mܛ s8��/1/(:�}j�M��J%v������]HRw� ��l�����4�!S�hP,C�6鐟�Ri#����C����>ǛT�Q�p����-r��)�l�1�,���Sc���x^J/��yxZ4�JQ�d���d�}=���	���5�NE��~?�3�ɦ�u�99���̢��8V�2���2�1�q�^7m�`19]A�����
G�u���z�~��8/M�#$�rU)6�!M�s��fa��/�6h�$�9أ�h_~q����V���2��۵����Q2�}Z�7�gw�?�<�����MK����V���������hAW��p����X�7��8VsYq'1�`Q*}��12g�V!xpvc��774�؈l�j���R�q����Ŭ��'捌}�an�n�^a�M-�Ge�|]��j�3�M����O8��=yp�����x��������m�d')�Ț/�9u��Y��נ�t�}17�gR�Iɬ�$ek|�~��\�����������cuB�ы�`W|�%�4�b�kGl�jՃ3�����RG��s�Kof��۪M�8�y��.KTA!;@|Ƌ��p_�t�F6in�y��9�Q���!�	4�R�R�,k�#�Q9�ψ�4��f�DU�K�V�}�!�G#�t��D���e�r/���W[!-��}@Y���:�
D����U�a-���|��$����J6ע��xq�!p`�v#�NS_��zK)y`�튰C�Uȭ��B��ӱ�4�PyR&��d\5Y�i��_�O����c�ϙa�ţ�h��|����Ң�)��Y�|�ߔq7f�՚�0nw�fUW(���P$N̹���9�@�AP��as��_�%�hO�!�Z�,@��WLU�D�pn
�v�� �_����(�F�d�L�U��Qw�T�ǧ�[��^��hnXmЫ�Y����H�!@�M���1>�t�~�+�	����a�~����JdcX�Muc/n��������wa���ȝ� z^S��is�d�>��4:�ض��颬p��eI�/d���)��Lǥ�T�Ȧ4a����4�=�χ��V�2�Nc��gK��h�xl�骢sw�ِ3N�{�I��@�D2�V�H�H�@�n7���@������a�̾U�Ͳ����4�[ȋ~�4�麇 h�ܺb�����,�&-��@z�h�^6���=�g�,�ڇ*T�����8���:J.I%uR�Im��Sgm�ߤD��D����ʐ�T�Q\��N���%�k�}e����+�Ď��K�����)���;fn�k=�9&0=��?��(��m;g��� ����q������Ғ��P�A��]�;�=�a >��C0f���e={)~n�j&o_�=ຄaI�����G���O<����i�1�Z��*礃�R2�������Ç.��	�w�]���C�~���6����m�'�ɬF֌ps'��ĉﳩcX�%�+"��!b�l�*��G@_�v&��ϩ�$�o�=�T��3�-��NC��G
3"�Dŵ����#��(6J���9��4���*����
h-[��݁�Ҕ��	?���B���o'KwC2m�pC_�ޚ������Iσb
H��Ǔ����y��ɢ����
����b��������IQ���C���������w�Y�'ŽW� �_�4�'P�م%"��a襠	��.3���D\�;�� [QHJf�� �Lj�s�S����f�Әת&��������b�j=�5D�nޞ������r����}�i9�L��3d)vxږS�F�7�cf�!67����g����d�cOK? !����z���Q�^΀mI�S���n�l4�v)v��{Z�	�	�׼䢏Fƍ<�\~#�bT�o8����Ⱦ��2��x�~0	*�PʯJȀ�����od���f���zS�����ڷ�
��f��L]SH��?��$��'����2b>~�D�ᡏ�������f��p�~���Ͳ>9�X7�6	�o�S�̰fei6)NC�`]W�5PG��/�*�_5��'��w�<�&S��5e��$֎=v���L��Lj���:�����?������A'3�N����@֎��L�S�A�qe��c5ʐ�Z��i|�B|l�jWq�&]�^u�L[�cvGy�*ބE��Ԏ>tr�k�5A�2�cf[�n�"��$lȣ�'u�oB�w�qg"6����äFK�!�GYtW'^`'2/�6fj�A҆����q-��]D� f4}�q"��ָ�g�S�C���� կ�A���p�.�iL|N�L�����u��~I+,H�I�������5�cf\+eb�q�Ry�i��)z�mU�~��������P��ry:I-�Ϻ=n��F�M+w�o2��x��5��]t���]�n�@�?��{���͊���"�c��Ʀ�����^m��^��x�?���;�r�ɖ^�#���e��0~�����4��i�x�R�E���'�_�	�i�y߫��2Cl!���+m�u*�<�N�0���U-�+���9qddHo����`�򺝓A�r�M`5����7��:�}�{b�hMJ��+8���N�k�c�_H'CB��C��u�ĭ��߫�j�T�2jlk���6|���_yt������ĉ�<M����"U�xn惹����[κ��d�k�Ig�y{F�@NoP`�x]K
���et�=��y��ެ����Bd�,WM�	+D\4K�H� y��c�{�M�Ft,|8���y��7��1d|�l:��}ǟ9�cs����	����%�:�����~Ō���~p=0Q�w��}Ѕ�;���s��0����b��xu�F9��DS�04������1W���XL����`�,
��pAd��5�j��>�<�q��h��I8�!D	KP�L��<�]I'��n)v����>֐q^�>��r̪� ����v]O�@I�˗����-��yT������c*����)����Z���zƛ$�c}�A�&����6����Kݍ�$E�"ke���k�'ܻ�ς�A�1���%|�{\�����d5�aW�Ql�L���ȁ{[N��q�0��T /{�؄ډJ��{I�Ac��x߸Hc-�>d�S�b�:t�X���Q�R�h�`Z��+�xZ��;�w� ��s�K|���٩_7���M�K��fbG���$��%Zכ�WH���y�yC?Jb]>��ǩ|fp�N�0��g�N��{И6�J�EΙ0������6��
f�����3�#U4���Ej��%I5�I��I�zC�g����b<͆ґ����i5�����
no�'4nt�I�#��c��n���q���΋��~xJ1���Fc^.�>�@Ut����-�K�n��Ls��?��u�Yl8-KfBf�C���	��)�:���F:0�jCK��/8�[n��*��5�b�Jm��߻�9q�+��d�d�4'
�d�s_�i���?��жu�}�P{�̫������:�R�9�$gu������|�T�u�7��"��)����ڵ����]�8���p]9u�:��x��)�[�Mb����j�9>z}�?���3ړc��Ì��#m�<;���A?�]�5��Q?1nJ7E�L�֬!Y3�;������p��}�TcfC�q�M�k>у��\<l�-�p�b6��S�pn��I	rI��C6~lm�p3��w����۵|{el�w���y�	Z�������&����z� 
b�hA��Zv%��x�'��1��g߮�'�5�������&�G�`]x��z�U@Θ@/CF��&�d�17/N/20a=�y�������5��i8���%��m�=�t�6��І�դ�s�g�'V��۔ٶ���;P�S�۠8m�?<g�?������,L��Sa�/(��0{*�4��9����o٬�5�6ܸ�����[y=�u�/j����e)R�����+�MP�nh �e�t��Z&M�2 <��gwZ#/�9��?�#{�"�g�V�f6Ec?�����>� �h�������s1�t7TW��IHh��
A��E�Ǎ&+��$�;ޜT-l�p��O��̮�d���_��P�I���~q���n/ӅA��$ͷ�.� KzΝ.:A�mI}B3� J��FI��%KMs={����H�`8g����06r���'������K\�~��r��.X�S���z1���{Z�y�3�"*��}�J����*�N�P)�/��pRИ��n�����`ia���������"Rג�ݺ�(�{�� �Ƞ��d�嬿�R�����#������,)�K�fڟ��z=6���'��x�_�H?��D��� ���9sN#(�q7q�)P��R�j���r�t�l#6��
��?�ic�Sv�����F>��A�����<����O9.Ǡ8�Ğ�q/<D�F���1Մ��f�x=��Y��c�_̑H�8�p��L��VY{1S`���0���׿.?���HV>���]�����O���]���(B�P8���t/R���|}Oyp��߱S�5��e�jReݨ@q���5Pq����J����M�F��C�U|�?����͎^Yi*����k~'$X�Y���U��b�sl��=�;nйf�����b���h�Ah�E�	;��p�7�4��M��G~�_�����-:���Mo�1"�σxy�!�)c�����Ft:z��R��	W�K���M���}�LÞ��̓Iu�P����ӲMe��V,!�I㊙���f���l��#�]�NFI�\ܼ*Y�]_n��؉�z8��4W���M�-��im��uQ�px��1[�0;d�شl�<�o��J��]��ON�8�� �vC9rc23l���<ظv��[��a�G��*�`���vbִW��cx\��������&N���s4x;�Hǆ�E�����Ԯ�a��*����N��~O�t���3��UFZ�jkg��RHc��%��`b���T�E�"(����ep��z	*�|X�0�>��ϸK��?��2A�4�!�a�/5�~9�~J�+��1�~���UJj��/g�&�	�F=�(�s���tw'�0+��ԉ���7�f�],rl�ʸ)C��/�����l�s�[��c_3N�K�(Ȁ~��#79�s�+�և�e�b�"����73k����të��7�1�U�˚U��J)���$���ުcn��Gx����ļ��z����v�0�y,�g
M���.𙱴N�qQY{+l�@�G���oF��]�� +d�`��3�Y�f���g�;�˘�e��Aj�����>��ݦa�V� ���ӣ�蝘(sZF����c�)�}���� j�y�5T *�;av�}�]���� �u�&�Yt�cTJ4�O ��(�V���{/F0Y(]�k����4=ŵ(�):�����JY��{~�쇅P۲���˗q���!�Հ.:X*�M��7�|ݾ�&ҫ�^����(ZwJ*�u}�O���փo�O���f,/u6��X$
8�^��:֓μ����y�t]���oS�l
u#U��?���7�ѫud��ε1�E��,0�&R��q+�#�"=ǅ��=;�kw���釬'8}@{������
��7��;n^/&��Hy2KW�Ɩ���J{�����coϔ��po2��WGx<�����υf���R�\O'Y�.:�<R��y
�	��-7Gfpb08�GP�Y�~Fl^7��G�"�i�fT4��U��x�Z��aҼ�sc�SHS�r�(�s:��l���ٱ3�Td
�y��aFRt]B�+�T�6ҩ�B��J��7�,�7bH��n]XO�@�{��5U�9���"v�em؂��B�Q�i,��*��	��2�R��>�h'1z�dvMҁ����S��w�H�����q�pH�v����σ���ˬ3 ����!��n�:�ヽ�7�~~�s��t"`~NU_��T/=E ��]���+��&=�Cŧ��<u��v�71��+"vm��j6�f���K�q�y,�,�I�7g�i�ZJ��+�Ĳ��m\���r���'��G���s����|>�1�l�(/�,7?��#��|[�[�	G$���j��"�ۦ�dqy:�"��yM���{Q����x�w��則�F(aK-u.�؎.��1���� �t����V!R��.�WP�G�����������y�1Y��Ae���PnE0צ̌tK�kRC��j�z�T=���2���7����yv��*��W4�Oq�D�Ce3�fM|dc{�j����ml����^�U&���;��9�|7�T������=���ZA���G����L���2�_�m����w��"�{~UV�
d}/;���tN*?�c��xl�b�x/�9�7���P�8X�ܠ�}���	� ��{����3�-Zf�c��N2�mzf<>����C�AX�C�N>�:�g<��}PU��w�ƞA�����?M���@���]��Ȧ����� �K���'>?D5O5��O�a$���E���?������Q�6�6������8ii�p���ό���$����s�3�JwO`ye:�P�e�V����c����RHPZN� X���4Q�������uRf?�N4m����$���2ȃ�O'O�4�b��%�g�
H��{2G�(3�E4�QM8&�v�,{�����"�&�E���ڲ�V�k0>܍�.�.7&���mO�c��Y�R(�KA{�mG��3�Ci>G5Y�%a�j�5c),j`�]���}�>�7�,0��>���~=��o�`��
?p��cl��b�l�����,�v�H{s���t%���ٜ.�����%:�/��B���/8�h��8�wn���Mv�r��'%1� ���4�&i�b�H�#�z<����dD7s,0���Su'C�9\�񲗪���>���� '�"��>*�8�!hI�A�%�����(tJD�Z����U�����^��g��s���(kW���ݺ�;�������3K��fw�I�es��1B7�=�aSrv<��A�;+��A6�)�CU�+������7k�p�yo�@�:9�ce�C8�[���~~~�:NU����G#*Ǧ�r8��>�⼪<�l�S6�↊N2,��2 ��f�1�r��<��$�9�S4�P�,���E�L����su�CTJ������a��NX�g�{4�iJu�i��9�M����H� ��]t����$Í���>�r��Vr�B\�+��f^hփ�^�=�GmBNv�AJ&(��������yv�	A��b��ce����B(����.�i��\x�������Х�PGL-%+�(qO�hm:c,��"�R+�iʪ���h0��
�dѧ�����;H���kr��S┡份�k�.b�R�H�s��!��.0Y�e¾o�:{M[>�G46�̢�=�=˦�؃}s?�=�����1�����FS����z��b��%���
P^�(���*�n�) 9�g���
]=(���{I֞��¦f��9G0��8�e�L8�Kn�kY���t�;�(����O�$��ϯ����"K�1Mģ8��x���e����3|�קQ�aK�K	]קYt���i-5�Y\ü��/mo�%ɑ$��G]@����!�-g������a�4n�*���X5��z�o7��BWeFx���������s�[��*P���^clO���
#��3�e.���$�[��1�U��<7��wZF$�i�����s��B͉�x�(�E�R%��2x>�ª��������$��k�R��:xѯSPO���EĜ�dY�V`E�C)+j��WI�y�':텣��M]rf�b����!o�$��_��2j��b�x�k�](]�NC�=�^԰�f�=+�(��@	�� ������ |��±lbj�s?�h6
�q���6�	-=	�e�N;��H\<��sS5��$6T5a�Ƞ��Nec���`�H�mܵi�H�C��N�� �l��Bo%`$Y�������������`��5���ϱ|zlbZfpCQ�i!u�EF m�o7
A뫯�7�~�6,�(���4M,�/cQԾ�xl�'u߽;F�og��n�Rd�AM��ei�k'ꮌ��;+P�<�
Q�|3�Q�y��i�T�~,�K#^y,��w�5i�^+A6+6 ���0���D�T@�e�{��Y���Z�����4Q'�}8�5mf�b���$w��
W�LEL@���}��V�ؘ"�����q�(SO�ȘIQ��@�n�x�Q�#����m�q=�F��
�v�4=oə/GT��6�����/,��r$	>�(ψ=��_?���h�� �A� ��W_�����,����C�V��@gB��1�ĳF��0�:�d��z!����P��o�f#��Y���R0��l�`������ɵ�&�m�E@9�� {	<ԃb��<Hf���u��Ҥ�	6L�K�{&A����Hܹ�R'.�qդ���))���m6�i�^~n�L�Σ��r`P�I�]d�V:�)����h��%}ǩ�`y�xn�gk���̱��#p~�����߾����6�$<���"����t�
*lh;�i�2�m�b��z��K?��w9�����r��_�Fy�����+��߾��0�B(?�r��0�qʖ�C��{��ٮ����g�)����q��I�'A&��B�:�]]�D��ҽ�����>(��D����G���5w��Ð��N���b�"	'�*����O���YoNl���G���>)P9C���ޔ��u&���]X7�	��*�t9�4X�n��/&�~����/|<�R�����"��k.f4m��N?Cs�ۀ`p�[js��\���ƴS�٬��$մ��RT�Q�P��q�!㎲~|�2��l�@��f�H�=d��Hn*�Pۚj�%���^�ЀQ�T���C@{9��!�0�<[/�Q�WQ�!��_�`�F ��]���e�
֘��f�=C��;][z9(��Ǎ���bŉ&�gw��Ͻzyn��*N@����:����x{vqF�a�Xl��V�=O�<Z�>.ґ{��(f&��W�H��6�~�>�#H�?|���[����_b�=`:���c�f̀z�E����z�˱j��g�yMk9?l����&�I&8`:c�w��F�(��X����l��bs�;�#�����l�m*K��w{mJ,�q=�y\Jg�,�p���}�Ld�fJ�Y{V=����4N'2j��� ������Έ�yhF�y���X�̀ץғ�J�<�e
�iL�m�<@��x����3��5�}���yx��8i�W���X��kς�N���Y��áʺY�������^���7����^�{�V��ƻ��$t��xS����Z��RQ�w{K�P��r�Jχ��bܧ�ѱ�����!Uy�6��#�1����E�n��,qlT<䛕��I1��L����r,��<1l�뛄���|��z�ƛ�����.&Nc�P.[�DF:*#����]����ﾓ�{R7{�	��,��!Q �'w>#/�����9�}H���?k��c#��F���������n��׿2C92����E�.2J�u�BN�4 �u��ʦ-�A��tp{w[��Ue�v��C��R�O�U'	!FlXa����^3�K�V? �B�F���E5 �[�aVm��'|��[�Mg�9�K[|�_|�(�dҺ�Oy�.��q`L:��+0�a��<�k���ӟ�k�ￋg^���8���l|���E4T��|��j�@��eUPj�:��z/l�n��9���v�x��X���%��5|��;+������������%��A�XO�7T��Wg�\6��d��5��{|�*CG��
� |����u�q`�3 ��Ž����z:�`���@l���z0�i��V�4�d���.�h&l�©[orl�3f��t[8�7�x�W�l u��
��h�T k�i~rH��I���y��DX���N$:FL��e|y��?1K�)�����v��^�pЄ���t�I=F�yL�
۞E���f�s�p��v?a �����������E�U�9%�~�l�����m�X�R<i;a�{U#��x�; 1X��[Da,�U'��b��*�rF=�a�}{i��B��D����*�^�e�Q�8n\�Q,�;�Ԝ�Ⱥ�sނ;�∺����#(a�%
��:�˼$_��Ui�F��wӚδ�e,�b�Y�o)���/�U0X������4q$��a�I˕I�fB�S�
ĵ��S�ߖ��t��"�]�;
�=�^�Qdh]<,+���Lx{��fa�b��2)tӐp@���_��yVmAPu=��.�,�t�~���=�����,��i�T�[�O��'BR���T�r�|��k��8	�� ٭ȸ�I��'k�,�"���:7���Y���,��'���t�R2FC?����Ć��hb�5�q����C���Q�MN(��^̄q2�b:�J�^��=�u+����:�8Q���qt�c���di+V�x!�I��}d�8���pJ3�l�4M)��������Zό�)~���Ked-���&��s��R�%��T^.P�W\�����"�R5��e���-����t�"Zp[��L�i�=��[Sy6����ZF��u����DB���0��|��C���Zl�&���L��?�#[�鬑%/^+�7�3�~���pJ��0�wI��GzD6�$ӍIc� L�̽��62�4曦@mK�FJ#�������of5F��W���޾�Hy�� �7Ym��{�,�{vH���j?�!�.8���/�|�ow#�\#�_)��.�Yb2��$}��l#*�`BL�J=��لrR�I���!�K[�2�|)�hv�������UȏC��U,1W{�6���������D�$~�(gwi�J�u=vzG���κ��a|�@����GT������b��Cq2Yrƍ� ���$G~�d\4vv����q-������|�X���nh:@����+H�Cl�3l��<�rn˼*|r���������M�و�
YFf��!�M2��S�\��&ס�L�eO�rpw��b�lE��TtO�˒� *p�����~�g��w�E�A�^6z갻�剘)!����ݝޫn��}|<�fюI'4gm;��NVb�6���xֽ�`T���f�^2�j]ྛ~�^A��z�R[���*��@IH
A�>�R��f䴈PSi�Zha2��H$��1&[�5`!�<�i<�b;��Nr��W����k�e�X9��H���y��T�������Źew�Q�i�3c�$Hͦ�@i*\S���43M���f�WA�E�y�|����aT��e/G���ₙcY[���$'F4JE�r�E�� ��䚑��Q
�D�.���ӘW4*����|�M��G�W9K��*�ӹQ��Ԍ�i��,�9�Å
��X?��ctd�	�������j�6��Dq�<�.&�6m�Aq	���N]m��ً�S�@S�[�\��o���[�̬�X�!����ُ�\���
^$P�X���I30���$΋�@|^��_� �y8�q����gqρ��+��r2�qm�t#J̾�No�jH^&~��v�lǇuT[�Wu�kgE������6���1�����nHo��)۬�t:Qm��OT���!f+x���b*�Mœ9�Q�3�[5����Tw�7�/���Z��JJcG��b�9�qh�k�PPT�:����28yև�^�m�I�33P���r�٧��R2R��9E�3�L���Nh�.+�v.�K'�m�T�}�f�L(6g;V���}r_�Jg|��;��J�(�҅��M�/���:'`r�;��o,f�fp4/4R@�D�e�#�
���ݖ�qq�w��1�$��R�i�H�Ji@�Gf?�����l�sI�R�=gY�FE����d���X;.��Ǣ��b˰����2�1ć�C�lCeYO�1?�k��m�ב�"�ޠ���w�\c���ƥo�mf�8p�3c��D�+��d�ēRMr��Y"P"S�ӟ���˿�Kd��m���.O�.D�&�=N�%�#>�ς�NX�af]��⾓4?&�j�[��@����C4v.9n��f� �0M��z��{�m�aJ͊�~�f�FجĨ���tO��Q�k��4O�(�����){�F��<��;g��sv��	�'fJq@��P�JF_� ��oD��NA��KN��!ݲpݞ�6���uY	Ն�N�������2�.�ͯ����Z�M݀.�k߻�gb��NknJ��`[����Mۖ~�_��e)?�t�T�ҡ1�����ڽ����kx	�*}ee�l�󘭢�*nD�GH;��޿��D9�nJ�%i�^����I���3��,��@����+��3o?OW�}j��O9,KC��S�L��96�KJ���Jn�Y���xA/|D!����FfQ7��h���SH?F��I��H�(1�j+�q/̑�E�vaI�qNp���m���Ds�h��pH��I����n��_�5,�br���=:�RY�f��C&�r��.������ ��H���%j	w��aAVɜFɸoab�N�o��L�7{q_� *�B��24�jC�Mr}�lA�Rs.�/_c�ف��[4�1��CL�4͹v�j�yW=��gc%�V-S��ZP�8@LHf@��{�u̺��;���I���%�nfB���y����Gp��+xw�3d��{���%��+^sf&�R��oT?�ҥ/��Wa�q>-���0Y�,�##uB]�ir��]��3*�����4���ë>�8� �|M�2��� q�4m 9��_*<ћ���m���UI�j�s�s�+#5-L���8�d�MbHX��[���"�1��/��es�5N��<+96� M2wpF��-4։^�N�+f:]��a-�4�6z��z�@Kd�������������K����W�J
N��=7є�M�y=�T�՜��>���d�m�7�(W`}�������xV ���P�<����w�4M�tHCeu[y0p��R�H���0&DA����k9@���9�N�e�@CF����J\Qz%o�LW�w���ްm��Ѡk?����e�z7�2) F�&�C�� �5�']T��V���&���IH҅vW������T Պ�倸�����%�k���!_�J���_|)��C<7T !�>rM��%�^�c42��|M4��8� ��<�#�1ӗ�@�r����x*���� tVYǸ^�3͈��"���Wd����3!�JJפ���������*���(H�r�����e����n#kG��7� �W+N΢��I=[}�����M4t�Mn,���v��w�������S/p�PoL��.��3x���:�F�V`Ҳ�42�$b�g�pa-�%7�f1T$xQ�ص���7L���� �cVxש��9I�M��ߏ��[@=ׁTʝ�$�/�d�xϿ��/������őƏٔ�Fu 3���@���SaXn�ҀƎU�E�/��s̉��Uކ�2,ݶ����g��#G��ݣ$�V9�:���ζ7��}�2oպn����A�e\Ot�qH��"x݋PV�͊=�z�gB���%2�+Ǧ�tWդu���̎#�G�i�(>�h;1q��Y~�e<�A����|X�C��D6I����_��w]�Xz�걼_ġ�Mz�l�y_LMv�eyv���x*3��b�cmWUn�&��q��V����v�U�;�kd��>� ��T��Q�������Sڹ�h���LS`�;��J��)����.�Η꿥��א*l����ԫ��>N#Л����=��z����gƍ�f�n���S��7?m%�c�z�$�ԝ�&��(E	dc="�~|`�?��u&��� |�]�_c����TL�X8X�p��R8!m��ak���Y��P��X`PK=�i?�Q������`D5��;�\�H����(^��#o������l�n��/i����+g \���iRb�L8�'^��ɍ1\K41�m�h�^ [��*��48^���C��9�E�� d/ �= ����(l;3�rmωi2�Sz1<>=�&$���\Q)�hޑ�iB:�?�<KV3>���uJLv�n��(�a�̭�����D<&֋�x9��&�R6eO��BvyxN(G	{0�8���(�O+�h.q�5_���d�ltbo��E�t�\f�i�zn&YYׁC�s҆y���FO�v����wU�0%���s�rh�ݤ�v�'�6+�o�wLI��)�eR�E����B�mRƚ.�&h�[.�ϱp�f��l�P(h2�g��y�DBw�t����ܝ���t��άH����Ԛ��`�a�����)Xp���4�">�C?)�]W0�QC�p���%�&)����q̬�e�4�-+2�t�r^i�pT��fe���Yphs�h=��v��$wR��o�J=�)���햍"F`s�<�n���'kʣ��d����
�U3����A�F�A+�B�0�F��lm'Cq@�s����ʃ�MfǨ ß�͙�sֆ_ �}�"�ДLO���r�����1ߩ��h��j�2ˣU7m�b����n�[������P��4�V=a���̊3;��2������i�pJ.��S�
m��'ǐ,�)ް��Y~���;枳�O���V�v����m(c��!Kg�fk�Yp@�EK����*���7����wS�S���П��1C@�8����`���1@[:T%�Y�ˆs.��	3#��8����97�OxS�U�3�wJ�J/�2��KN����.5G��('F���z�'m&�g������\�<7���68�Ҋ���>2��T:�'u;#�u�F)�y���0�X����"�D*�kh�=Y�%$0��&A�뮨GyL��Sc��r�(Z�$��@��}f`��̴� �4pZ5n.9\�^�? `�ؠ��"f�>>�������2q��������X-�5�1����~U�7~��%�k���jp[6�i`rQC�n���slXVFR��EIKD��Y�3��N��qO�%;�k���|WF�D6׀5PH�0�6���/6H>s?{F�K}�{�v��Z�e~���w.�B�w�RPPs4ɜ U���M��koa)͹Y�|��59��Y??�ǌ�;d�]6�@S��,J�J�>U�������r�m�`�KF�R�&�K�3g'![cP����S�����?c���tb7�K��S.��Q�Y�62���4��c�1~�H�X�m[H�{M��E؉�_c�X�6�����<�5n#�nU��̥�G��8]^zzfdx�0E^9���3	�����玁'�I�*�!切���;O�8P
aL�9�����s�2̂��X�-�Q������D���� �88�02x�ψL�R�M���:Kj���`��[L4�����Q��q�q�Y.�|��:$��|uô|{#� ��Ө	+L����ಪbj�Ͼ�l)�:]8(�����4	quHx��Q	M���A沖��]Q3����\�A��?��;%8����\��:Q*%?��%��@���E�t��K6��k���DcpV���[�r�+�V�d��{kM����Ep����p��G�ԕG�j�)�֯� [J���7yA�a1�~�@�`j3| ��	T+�����N�,+yZ���2��Ix��z<����6q|�����ȑ�ƹ��pG.S{=�B�m����`锞�)�<z͓?As]D���he����"��w)_{N��� �I�[�1�qd�n9}��� �gc�jE!qY���(c��N� ��-4|Oݣd��7#�n��g@�q�Q�4�=��d��>X����|`^�.�q끁r��f�\�͉�svs�U6G.t�w���W�o9r^���"[%�=CWi���w�=�0�FM��#���^��$��K� /�B���m*��������6��4�1_zH!��.�_~�eN���8d�us���,���,JIn_�Q��T���#����g��G�_������;b��cjH[V<
��.wͫ��f����\���E�&fZ=+x��6��+OˋL���Ձ4Ae�*���ɂ�ê8�q�:��-����N���^8��Ŗ+2m��)��ۣ!����Ҹ.�EZh��Q+>�5�5u�]}g,(&�T���1�?��!�� ��8T�l��u�m����*l����Y?�M�،����K�8*��נ<0��X��ٚ�m,�'��Xg����%��{w�?~|l�_�}X]��añ������a� 4�(���q�����ǟ�xp��Sf��.Ql����d?ٰ���_g�沺J�N��>U��n�%~�'9[a�̼��SJ�s���no���(q�-����F����.l�ĝ�/����s�)3�h���З�����J�$���9G�3fb�����Ҍag	G,��]w�t��bmc���0L��X�bu�iT�lx��4�ȴ�ݴ�����I������W_4�)����)��~��.pX��x{m�}6$�R���	�iҫ��t㰩����7&�<�F�}x W���
��]���v�|�)�c�+3G �%��7��г�C:����@�,iȌ�;�/��t׍eH9,�jsT�ms�Р��K�,���[�}���
&o�N]�y;)���o�=��+��t�i�̨m��[ß�a�z����{�V�lxJ,i4���g&�Ɗ3�e��V}Fv�R�6}Rsa!�/�7*ooڰ��Ȫ�`np/�$�cr��|���>e��M�e�� �*����܀<�\c���3����a��������Į,�F� �؟bM�x����י`���q��
@��Ph:����և��u	��z��q_�6y��&*5�rT�%����ͻ�-c~���wKc��ujI��ޟ��;�K�{�-�%4���`�/�M�b _�p����՞t%ܑ}Y��=)�w�ްq�>�u��EXm���l�:�������,e�(2P�z^$;�O�p��(�t�4��q#�����N���p��&�����>FT�4��|Q���j��P�M�sc�����1�1�"�M�moZ{�DK�}_�ї*�7�>T��+�eSloQ׵����B�97��z�a�@=�{���mT�س�NZ�����ѯW�s( &0CU����&��-���8n��0�o�,\�䱰ەl�[��`�S��R9�Ҽ���|�j�͍��f�sSSB��vr%��nJ����5{���~W�{ˮ36�4Wt���i�lx��A���������g������Zw�(s��T�:Q���1�ʠD�����i'8����l1i_�/��,���j&�!��|#9��5�ak���*Yn[�)Z��֓�x� �	�M4��'A{s��C$��_�^��=�S�%��Զ�RhC�������ld	n�(;D �2R���r�6���	�f���DB#�����`؊	q������4.8Ci��ҐX�uĀq��wl�7����RT�_����GfT�������P�)��kz٠���C�s�y�|��R�_��;=R�{%��6�uƀ�/������+��`�1K�����Gm��{�L<s��:�{�DV1�3Ͱm��f�"�dT,���22Wx��kUҽ|#k�@�á�%B��A9gn�
[,
-X�1�'#� >���u_�70Py��D~�R��8>�,�X��.���0�d��m���-�$�>aR.�C�Te�ӳ:��8]� �:�%��<�>�}7�J��͈0�ޔ&sm}�D}S,$q�M�2��C�A��}��2���|PvU�j���&3P|1#�l��(���ܼ����<�������]J�J�Ru���L7�C����b�:Z��~
 ͓�ޏp}�����Fu|an���x������@�.�up����1�~ l�:6ö�!��0�0~c�"GZ�Tj�U&5�pJ��涌��i�B]�D6:�`��N���q��_2�H[��?{���-�󂾗��L�삞����O��cÍO�\�Ӑ�52Ͽ�}`y��ϐ��<?W�0���(��}YqOCࠒ7�ޗ8p@c�2P�p�����ͻ���D�S!|����p��qzo�d�nS5<'O��z��D �O�/�M確��&�~��b!vWv������5�1R��{̸��{=(3��(8��?Sz,a����+������>j�wK2yΠ>$��1*��:�����Z��'{�:ؔy\�+��;�����jLm5�[e{-�d�.��u2D�}tW���ܧb����Y}���r��y�&�4M9��%���[��
�j0�������b�n���ԙ�L�0rs	/b�,��б(��`� ۴ 8Acc���p^��ƫp.J��W��
͊�R�M�a��AϽ�A��G�뉛��B�F���,_���u�����L56�v-�N���-�4�<4���{��,�sS��:��)��0��e)2��� ˒2TK��9p�M�q�҅G��>>�K� $���P<��y��2ݗE���E��!���D7ő_���2��܈'q\a�;�^��93�������Vٜ�d��
���>��XT|�������[�-˳�A1�(���r�6¬#���TLpxcnf��Ţ1"8,�o���b%ם<)&��;)�)o���=�zu"��d�{9��Zk8�U]�GK�F6�j��(��WY&�R�Ӆ�Y,˹�8�u�s��徃�C��޴R������ٓ��(�d�kS�&:��lBf���_5e�������'���2�Ln��F*L9k�	X�(#�,��ǌ�v���ƬZ��,~�4�8������F���$wbww��>Ǉ\J�	���=0By��)�m7���#��걳P̓�u� �W ���5���a1�����*��Ә؛ڭ��M]2�L��Ӷ ���:��^�.�<� �N/7>7��l̋ڦ�A��4Gw��@�86uOef5yѮ��0�f���C2,�C��+0���߯g'Y���n��"Sb��#����d����5���ϨƦqMlh^30<�A�>p���X�1��FlPC`�"*3;5z�>mL\��)=u}�v�i��㙙�@��!�_#o^�r�4"�/�41�纕�{��` ��BL�f�7�^���U�YU�]��A}�ϰID���䁽�SB�u�9�nNA�iz�R��:����L��06=	�ROO;�@�	��%}�?���A<c�91�zo��e4E����5%SmMm����H�ԚGF��8�"+@ E���	�p����O,��������_8��&=�}}��ߒ-}�x������6�^���0Ͻ��fm�7�-��F���$�_M�5�]nv�ƽ�=Q�ƍn��i�\`[�7�h��1�d����?���m,k2�*w�Ѭؑ/Y4J/N�8;����8���_ŵ9#9�M\��ک���;ós���!g�tS�f]S��r� �����ր���Cʺ,� :�\�dM\ {��'��(������?���x�~�1~�� �V̆ɚOWј���>W���H,81���3c2�׸�ڷ7t#��6G�)4%52�b]���R�nu��X��3�1�X�?�+�6f��,y�3z���=����F��
�E������N{1,N�bA�@G�g<�Y���GAp���^��p��z���Ax�JE�����U�������|�!�v�c�y��8�XK�0=E������´ƕ]gUΧ9t���+��P���yvٙ6�T����u���%VL�~&N�(���H�ǆ�/N*yZѽ��C;��RWd���r���NI���1��E/������'g��ˉd��X9����4	����4-[�a����z'�Y���:��e�ъ�]5�JJ�]~L�k� �!�]���m�Nnȵ��M�t�r�i�~#`i���A��bq8e/|>�)i�U�&ԃ}L�->_�͵�T��J�'|Q�J�a��,(X��MX�}�k�4��ڰ�^�Td�;gI��n����T/�M�y,r�e�Y|j��Wj���-$����#Fȇ���_��p�x1���g���{b����~�d��P�lb�i���Yn��]i�n�H��ɺ�7L��$��.N@5Um���&qfS�z�~~Nt||VkR���0
��p <)k�,�"-�T�;6��M���T�1��)��aQ��#�ǌh��):5m&����ߨ����5(�����/�Y�ϛ����s�����A�����Cxo���w���8E��Ą�S�r�Y�]fk[�>ϓ�� L��`nY�*�S�������Ʀ'�Xa�pfԛxp��a�	T���*ɁcE:aeG)����>F.��~�/e+J�[e�&�r��Kq~wr���8f�Nd��������D)��uQ��ܬ9u��v���Pe�3��4�Ep�qo��FCI�`jf+&S���;V�q�T��>/mn3
^���������ʺ�kr�~u��ָ���5�VKf'�UN���,���BZ��X��oOm�)x��!��ao�S�Ϊ�F˖D�[��L<�����2J��4�;�s���98�7����X��TT��FD����U|0��ج	��|����$+�S�eC7�i3����I�7{1kl���xP��I�T$�sJ��9m�񰽖�ּ�O�گ��x��4u�Q����rڞ����Y0X'�pX�ᦛ������b��@�}�}`���؂&"tG�S�f��lY��pI4�.�Kb7�xQ0��J�oH��@̊
R�l�\�'�"�p* �OLM��k�gPF>>>G ��6���t�o޼M�2�~~������M+�nw��]���{��K?<�:�#"�h�[2���;�Yc	�>}-��'� ���_4� ��{`�LIg�^[�%`݅	�=9���98āՐbi,)�Q67�3e�y
����"�{�����R<2� j�b6P�T�é;%f��n�d��F�d�T�\�}�ad�^�i�����.����UY���&�|AәŪ�L�1�t��o������Q>M��r���I٨������PJG����!i�3Gw��!�S���kAL�i%*q5P'gnBN�ԊK��Wq`������3���m�at)��|]��� J�X��nڼ����.UinP/�y(qJ���nt[Gp�i���h��,{>�a��}�9�T�0�d0�9~ߘ�%t�B&�ō����`�E��)�~Y8�� x.~3���5y�y�9�|x6fYȓ�c�%o��ˢ<����?��|�Aux�g'���)J�Yۆy&y4�@0�TJ�����{�9@�,��Feea�f$�R��ᛵd��V	�1C2!,C佚��{�n*��mw��ù��g	�$�������([�!�X��9�-��kڙ�i��51��oZ̝e���g����gLh�8��E��c�,�ָ��4B�y��tU:e6��tj��A05�c^4�`
Y蹂]w��P��%��x�$z�%��巌��y���DP�l��Pr�0�=�J_F�d@Ul5Q\Vb����,6���1^sQ��:�����A���eucp5l���iu̓���H�oZ���<�H�ba1v� >?��F�w�)���%� ��C��h�ݦ���>���]�H��)_����=b�&Jh^�I1j�a
��'�N�o��~j<�&��ܯN��4��h�=~�p�8�<��?�1L=�Y�a#8�,�;���y���]wײ���I%�����^��D�iZ+���H��I�.�M*\�(�=ӕ��3��Z{*���.����ŴLX>�
�,	�2���	��EdPZr�k0��� ��:n�MZ�������au������1�n�{%��w��<��{i��d.�3��`J�V�gѦ*'�_U/m�\�yT������R˹��]��πR
 nץdf��W�L�W��3���)��7�:j�GT[��B\۪_p��ppHu耯ej�ِ���⩮\P��7k�1��� w@s�H쬷mϴ��4��]36� 2�@>CH��Q�y ]��"6��;��m������:!��Q8]�KEO�Dn�M�d�Gv�Tq2���a��"c܂��0#q �pG?���6*ֳ,�z�:X������������K�����N� �i5tش& ���d���aP0�,�&%��\�Ў�/6>(�����j��┼�F��7�X����G��O?�������ⱽ}�/�z\�>(�ѥ�����A��%�~�̂"�+����G(?j|G,�˰��#�/� �>+d_fk�P��������)j2��r0y���<>>�̚���U��i%�~O���C��!'�YY�	���s~�o�Pז15I�V�_gY��d>�$a�9�]�'�,,�u���S;���A֒.�|EYT���D��9J�k��Or��V8A\���E�/�st�=�k�;��=g��f�i�-wrXZ�����3x��eBc��c&H|���A��@�З�wa����Nji2���^
�1�CH��"=���h"�s�̋�>��
�w �h�������xsQ��}�>)�@���cD�qB����~<�g�
Q�	K���x~���ũ����nB`�D �F��ہ�!��"���y�5-=��׎����������Ο~"��2ԛ�U�+g�}���q�=�o#�n��<�n��|�IG���ȝ�-�e��o�&��}��7�Ձ� ��$[6\�R���2�&�fTW5r�?g��y����sVW}�3R�0�T�y�l�cd��0�e,Ψ��5��M.OJ�N&0I��̣R��B��G�\d�,�=+9N�k�P��N\�6�[1Ľ��� ��o����$Nko��*�2~�TA.�w�t�Wȴ�Xq���&�v�z&N�C�I{���)�ؤ��wf׬�� ��:�RY���N�꽫��T�2��⻚/��U_M>�%�+Dg���Vu���49#� �:#-1��LF�@ڔ����
ݎ��БG�T�ߍ-����VG���B/�ޙCKG�_?b+U|1�n��F���W�X��$!I���J�b������u������x��aC�}�۝�1L�0`�$��pP8fX�vYo%+��D]��,�?�d���J�5^������Q�"��Bڭ���H佨b��'m�/�S��3�< ���/��N�/ۆ����,Ɠ֤��|�1)[x&����5%'���������+g��(K�u"��F�q��5���|Nbd � g�Ee$��;��im����̦*���D+;��E$���l#��y���I/2���D���hn.A��9��ZΑ��]��9�YI��x?ާ�m�*�y����m���'fK	fיJ��=:��r#C��!7D��}G�*3�i��w܃�T�1��s�#ڶ�/��U�����zN�I
�?ǽW�|.���u)�u�n�^� j�>I�0<� �Ĭ��K2< ���I/�u���/��.�#8�)vk|��N�qN��eе
��4s�J���/�
�r�����H}ّ������7���E/����駟�x��<8i�Mß�=��P2���E=�6H����Wo�����n�P�=G����S�O`%�� Es ׎נ��)� #펍������*c4/����F��b�� �Os���ŉ� �v>gC��Y���x&���L��M8��$�A3��Z�� ��H�?oA����;���D������1 ��}0��'���--�>;!�3�E	��t�#P�@	Li_���H��SR����Ħ%�ƦN��=��`�۪��{Ѻ��m��~'���)��,$��1���[y<p�Oߍ�����l�B	��T��n�u���!
�ag����\S��o'd�ϱq���<���^A�G�W�}�5��0g�4<\?�md;�2�^��|�����J����yev<?_q[���^� 21�t휥��o���d)�2��A#�q�$��
�����p �7VQ��&�7H�	�X�%����M���HX�H�h�C�w�2 /
��������Y`Q�K�["�k�{��ft®��JWS�����a����.r1����.6���p�D>���[��D�;��@�׻��n�~7��d��Ɗ>n7�*�, ���ؠ��NGI]P����;L��.]���x���N�q�+�)DzR��\t��^�>,NF�5�0g����(���p�0E��Rk@���I�m���ta��ȥ��ÓuC�����`����[0�@�uT��^dYr���j��ˢ�޷�J�Ms�c��M#Ck��ڀ{�!�?ws8p� �� ߿���7���6���/?��������ݑ�Fl���(���f+���-dk�M!HrNzN��<�x�@p��/�}�|����~O�7]$F6/dN�z���a��@;Ӿc ŚG��s�o���=F���Ҭ���7p�9�9p�4����f�f億��|���~;>ӽ��Q{���{�͟��&l�f+�O�۵D����眢d�1�`]5�'�%�L�FK���}��7��8���@�q��6�b�L��y|d�q�(��5'K��=W�Mq�*b�Re�:�<�	�onL�_���g�l3�L��t�)m��F��̛>"x��lyҖ��iX0,�E�^�X(� ݨ��iO�����?b��|q$�I3~|�t�6jb�KwR��s}8Vc
��)p9�{�.�X-��ԚF�;o�Ԏ3r�����(�E���P�0V�z��yFZO�$��IC(��%��L�cPf�)ʦs �`�й�/�TwUZ�ع��XfyM����u�{�1Ӫ��\0he�(�o�SG��x�z'Ïm0���嶆c愆�l�ز��b���hH���.q�e�rNyl&5c��j�e\G|�ܦ�:2�(�#���!+6���g�X���S�+e,�=+2n���=B�*+�	��!dm|���(Y��fI���LƳ0�N�F�d?멘|֢1g�x�8�&�L����XmIƮ�kM�+�֪,.x�K�h��s���X+}���]?F�����JW��_�is������--�'���%|%�t����_w����B�n�7�yYx�'��^�R݊Bc�.w=;�zk�,O| �Z�T�1�AJ��KĦ�M��4�?+zp��09�6��%\c�vuIղ�x�v�t(DMµ��o�׊����)ʖV��9� ��o�gv��k�tcbv�9��Hd��,���[��������oqx��͙3���@�y:����:� �N2�54����y��V��M�o۹,F�1�]ݥ�S8��,���أgڶ�� ��aHޯ?���־��}�yL:����`>{I`=�q��ro����q/A�3aj�b?*����M"|��_"X�M�G���NH�5���<�zә
���<�Ij@�g�C��#���_a�"���I�׀o���u�ָKޯ�=�>���U��iK>үb΁A�c��,M��5�rI��{;1�@)�1��yl����ۃ$�Or��l��ķ�`�k�Y�wG�%Mmm
VZ��?�G�2��"�^�Ц�Qzh�@��$;b��ֵ��u�� r�b�f�x��ڮK�Q8׬�t�1��q��.�!D��L7%�p�j.[�W��v�q�|6.nD�D��.�%mſ�C��RG��<[׹c�I�\��ÿX:�ylL�/��+�*���&3�V��օ�]����a��Y3�,R���F��N��ۆ#sM�>����U�/AɄ,�ǭĆ��?� �-�Y���f�`��r�՝hHX#�7�=m�I_鰲
-�O�({��b4��3�l�b��(3/���9>�YA�����M�H�'�=�)*#���3z.�E�P�=�2�ԝ����d���:��Z��1�Q��rfFM�7��0a�I�(�T���=�ۚ�I2����k`6B64͞%�5���;�a95�����I���/<�b�{J{���B2�]'��c�b�Pp�'�)�C��(�	fC�f���T/i�����;�g7��^��j��ŋ������T-�I­2��-K�J��XO��,m��=�nyN��>ưm�\��:&�x�,�Zc�������j5]öa�|����/i���?G@���m����5y*K�VB�� ���P�s�J3���A&�k�K�FiEcj�Ņ�(��В9�^�l/��I��69�wH����"�����G6�os�a�>h;e�ͮI�cL˒��x�d��T.�T����{dg�q#[�����?��i��
�"�rh�GC���nnL=���D+�pHI����Nb�ΰ���~Tkm����l�N��xm�*2�ݠ9a]2Gf�0��º�tд�,��/g�O��@�,
g^5��q?q���1>ײ��ʡɔ\h[�uZ?��������hY.�g89� �jÉ��ɋp�sB��uK'6�;ChC�j6�j��2�!���*�z�Y�Ћ_�*#�"�q�4�~'#m���5��?R�Q���n���q�	�M��2(���y� v�悫\�U�)�p�_������^ȸ&s��k[��{)��"a�"�b���!�>��
�qʽ�3O�#O�M��  Q���v�,��@`�:�0y���,�f�9��-���Jn��3E��	���N:`Κk�9=�����ޤr�c|˜�Ix�����Y�̳�"CG�f����	�*��t�7
�t4Q���*?C��� cMT����6�u��A�ʵ���Z��:8�,�!� �� ����/#��J�׀_���	��v�M��k��NW)�y���Q2SNкS�25�-�](�.E)'����T���J�S$��w���pf9'UR��|`�9��N	��қ�Ik�<��'�9��Mr9+ZT��mIJ�߸'�$���s}���A���:}I���@eZWl�LM8j܄U4xk�|�+��$��h�|�{�;ߺ��5m�E�R���w;��A:��u�)�F>7��7Sb>�؁�q/G~݉���1�<�\o�"�ax�S�6�0�ȲbH�a�s��Ϣ�Pl��I��$�"��T�-6M���}p������,�����
���͑��p���>%l:f�_���tN�f��&y^�*��3=-��F�-b���2\n��@RM���OM#�)�|ʶe&��K�θ,5V�HRI��׹a" ^��&mS�x�0�"�~_e���C�t�?Ŵ����j���f�&u������8c�fj����wsS��<��4��7�gl�s��m�� :��9h�om2�Izo�c�1JЅ��A�mmoWfs����5(�YG��X����-K����KBqe����l�Uc����`Z��1���VAx}���z�����?�6�T��%�$W��j�Ӓ�f����(G3�X$�/��9�iu�_ ���P�͑PCIg��B�D��$�o�0Ң�iub�
Oϻ|�,J u��@�a�(#XV�j����s�lx<������.`¶�r�K�_`��2]s�c^37�>�3V�"礟�"�l�fε��ޱ���|�,�c<[��R6��s���]y��E@��_��u��+�#4��bY|�ή���$|tl�ؔ}�U"��o`|�!🃓����n@�y����=w6�H��#]͓9٘f����"���_�mp9)�El7D����*��,�U��(�×a\3y�X����<)#�Y�B<�p�K��^8{dG��,'�d��]4m�B���V�6��4;�[mSd�1��5�"��t�)ẫYMn
{�#x\�y}����J@3���b�����������_�o���Rx� �۴c[���=�&1�>��f�N����"˙��QQt�Nr��g)vm*�Z��w�&~Cn�bYݵ�H�C:;����3~�,��u�ڬ�Уr���%�������~i5hJG8�C��of����jzj9d�2��-���;���V|�S�lR���]r�S��0�����͍��K�YT(jq3�t:$���~�&q��Ab9_,g\R��g+�*�Nh��נ��1<�.M�Xm5�iG�����8�p��+�Qj�x�᫮�<J�������ܗH�g��.���su+iO�h����`�"��if�ߋ-��;����l��ƥ�hx+�c��{�`d3�L ��~l󹄓�4�~�V<�U�H(�m��k�%�l�ϼN�+�BU�nwJz+�U����m6���X?YǱ&Va���!��B�S5�K��~P?��*�����/VϪ��
�i��UÆ�t�Y�T����cP����ܸ�Յ����Ok��MRVa�ȳD�|㬓�%��d��$��;������D��"���[�c��/��=���p= δ#d�m�V��U�Z�~/����yJŗif�0ծ{�Y9'Y�9�����&��<�!殶��v^����P9<�<�i4��RӾ�����	��z��U	۪�߫l7f�/Kf�cG=����P;DӤ�	E�͒�*+b�#6�F�x@b�YS��>r�{Q|V=��R	;n/muh_x�j�b��3 �9���.�b.9$ig�hvSVD������b"��g�-�-�94��ac!ʓ��Sf�f�Օ+L�<���T�4|��?&ō����t�g(&%�C&Y\�i���͉�\�y�OSʭ�@`}a]��+9eYXWwu)��G�^����]:W)�^c��W�����z,�'Y���d������0�Zƌ���>h^������&%�����2�t�yr�F�A�9�ķ;��?4:Ѭ���ǝXnl<�).�.���"0��,-���ŉWFR�዁tH\�Q=��َ'gR�p�&`=z#����I�ڙ�e�ă?f�
�a`Xˬ�F-�P�|��Y�Ɉ +�^��b-jz���C�
U�I�xַ7T���R�z�C�u�Y��^���vi�m2|/��PVm�)�tx\�����6�X�!�M�N�n�:�K��B�!�
֭a.d��5�a�*y�5�:�]���%��9�nI�:~�gfuP$��R*<����ɽLz��>:����w6}��j9	�A�=�
���ʒ=�ص_�N<�4�Q��Q�8���KY.����'�y2�Y�	+���y���a��?�`��R��1�H����ddĜp��+7�.2]� ��W�Vu:yFэd��-u��*BqY�P9.��׵�01���4G�ϟ~��)�<��$q�(s�&�ӓ<I�H!M#o`~��2cf���M%�8�-3���<��(���h�ݽ��Ha�dV�4#mx��)��=�5*�V�iF��F�4�逫�h(q���ҡBd6r�r��.w��+?1֋�幡M���H�%��Y�0���d0�Ф8�>�d����^�^g����\��HY�D%�lR6K���g�Ua}��)�X��I8 ���F�ޞ�>��C�,�1�Y���8м6����cn����.�5<�sg�l@��!v�fH�����ƣ�{M��p�w�s�ؘ��8��v�n"�N���=	�1���(��u���T&P�)|Iθg�a?n���*~�!���U'ALh֝wW;�=�'ko�G�3R��LFZ���H׵�F�(��61-gFy���߸]�w����N��i+��T֮9��1�S����3��KGW��b,�v��\ۈ^Q@�Q�A�|��7GF��R�cH.��X�%)%48�qY4�b�U��1)��%����ʱ�4i �V4�LkuQ����̾>���xg֗�w7�l�|>�$TA�ԉ�����h(�~�:!����@]��MU�A�]��i�^�t.�쯊�������p=�O(�}ݿzhrw��[:��~p�fW��5qQ�bB7�1��P�g�{�p���ϋ�Di��E��ڐ괬��5A��H#�T���Z�Z�h�?Fè����9L\�xM�o�g�����r"�	"���0ݖ�k��Xi8'_T#�y?y�5��v��|�z��`�{J�E!�]i���ԡn���7��@Azl��'�[j��a,��2V���h	���L�烬J���Hݵ��r��t�@�H�f4.M��W�&�]���z��N���7y��&�͛�G�t���.E��kS����Q��:�TSQ-�t`�h$����ȚsF92/J�zZ�����o2h��ذy��3��9"��@�S�Ȇ�D^b�V�pZg�x�Q��|8c���E�YT�#�7?'��C�h�\^󠮳��w_�`�at'y"���# źa����B	�^0>� �?᱊ �V�/r������J�q�8��ZB$mǉ���4f0S@6�p�s�7{A@�j��p�f��w�4ظ~#
/�=�Q��7�����b;Q��wM�~�#h�n��й)��A�~~����43��:�#��%6����g��,��0K>s�ߢ�vDw���'7��m�-��\q�C}��ۦI�ʢ
�6[$�m2P��6,a,��$Ţg��jf�i�����5��~�?}^��ry��PQC�I�ۋl�I��WY�$l������(�(���5|/ܫȿ���UWC����F4����(�'�t�w9L���f&E�$������ѸG�i���� �����EG]��;)5`,�sSc�膇��+#�����И�ؤm��8�CO-&pw<i,&�����9y�,1	���<�
3S��s������?|����C�8�1o��Ls�Q��1�#�:�$�%�mG�����<���k�߾�1�����q�@#nEU9�]	9�"��C	=��l&����^����;�D�����2e52W�}Urj��)3_�!d��u�ּ��ٸ!b�c���z1R&G���<�rݷ5�N���u��3�j�e���9�$^���l�XJ�U{ъ5�xcf�n0�ss��.��\s۵\J3��Ø�<����@�89����m���q�}����z�������#-s.������S��6
�%��.F�y�n�ǡ�瞢dyN*1��2�Y�k���~?���.O�S��`��U�!6[����[@�
1N��_�x�\Nqŉ\��є2hgvΡ��T�s��}�gp�Ol��]���	�/�ɻ�)֘���Y
�4~Xd��/F`c�@��#�w�ϧ���hr,��P��̚��0�ǁ%�NF���ڥ�g�m�J� �~�9F5;$��]��ҥ�WL76��:\p?(�z[�<���6�a{]��Z��Q��j�b7�X�]���5Ny�;���(�L�k�q��E�2����Y�S��8ֽ�z����J.([}�TݔP��"�RᲚ��g0�T|RE����	���@'��|����a��0f%���TS��YE���$��:�4��$�Fت�Q��_QDbC|߾A��m�N|Xd0�h8�l�MǇ���%�K�����kܰ?��@4U�:%��F+M�R�0y��%q���\��?�>�B���V����>�n���1ҏ�=@ևR+��{n�eN܇#ug��paE�)�U(�D��(�?������{�ͽ��6�7�>Sȸ�t�[��!J��?����/��~�Y�8��,ИXzf�?1��S��	(������P�|O�u]��l�x6V��KV5'���
�_Q�1K�f�mbd=bH�3��:��STcy<�߹�U��NIu׾@5Vi.(8��:�R���D21���m�c��T�����T���-Y��<���Z�W��488.�3�|A8׈ς�2Z��\l��B>�!ACZ����r$HV��*ύRq�Y �??۵���w��e������|����ϥy�ল?��.QZ��I�g��.�ܜ�\jM=8�
�ߠ���J}p�Y�E�8��F�x6_�7��<7=��p������
�� �!���A��g�+Ӡ�X����������}�n���Ǳ���ia{�w�Y���_b��z�@�&��f�w��u���<s|��¹�g��
���r�u���!��o��cR+��ѐ ���>�(�n�ϰ*�=�ߕ���~����O�3+W�a���D���լ�!�����L	�1����g�J��>]���wE��k��xFs�Rlr�L�����X��@R|=�y����X�'�\씕�j�fIO�Ľ��1��hj��C����/	�Ovmܳ���tM*���!���?�k�F�,;����KQGէ�6a�j�J$��_'�y�,c���6R�Ikz�9��`�w$�՛X�.2��n$E Ս��Ba�	0W�� ����G�U�zzv���6e�VH���)êo��!3fw��6�RЖs�8���9e�x]g�����=��x���"c@ Ģx��}\�߾��j��F-7~/ot�줢BP����Ok�EA�d�`������
��qEc��C��b"f��ms������8��S�l��A�8����x,�?��?5?��8$0K甍�c�+B�2�Y�S�N�k����jҽM*�TÍUB �zwc�@.�| ��_B�7��_�n��'^}��h:֕�qy}ג/MV�H��akwwl| ��7���g�����YwI5���|��3�T�;�7[u�EW����%S�,F0�.6���c������W��F��~G�aQ�*F0,ĳDe��#�q�G��{�
�P�M&��X4k#���t�5�d��Ȅ����T�����l��2�G�pH+��*y�D�n��pp�H
��+g9�dGv;�O�@I�����C��Tc�i��yCyHFGUx譺w�ZcSgr����r:���X(8�%}knd������75GL����|Y�`T�z�46~X�_BF,�zTm�6Q۷3/*X��0B�bx�4΋(c,�m��,�!��3��[פRF��	ev�ۙv�=�s�����3�ڬ`ڒmj�2<�#�nW|f���Ʃ���y������9@LA=_�3=H�k�g����wYJ�I��.2�.���GY�iD�F^�����>&�`N\�
�*�d��4}/,�� $�1iQc6��<U�*��N�L9r{Q��� �t��v�g� �S�fH��x����� �ٿ�Z��]��@������ � �a�w�A��̛�q�<G妜�I��h�]�Ls� �W�z����� �2�^�A���w�lZI�i����:���u�>��R:�>,�ǐbC|�ݷ�-`�����L���bEF��Rς-�L�Mՙ;whw��Y6�o���8���� �g��� ��mt��f��u`��S�휵�Q�3��=;��� ��1�9cZ<ὐ��0�A��il�G/6��,==���������o���)�KM-㋱��=|9r��*7#�w��V�D�aq�h����2�����ō	��>|fo��vʵ�o�u�2�1u|ſ;�O1�`�ܜ,�8�3?g��lM����7o"Ƿﵫ&߷���\8\��p*0��u���A��ˑ�t��F��_�=r)o33<W���Y�#���K��&�ۦ�����+B�sc�Z3'���r�eʝ!$�3D:��D�����n FQ�!'>H���=�'=k�ׁ_���cNXH+ɮ�l�\ }�w��H�iE�)|��8#�Ƞ�/�axw`]��UY���Ͷ$�S7qcQ�"+�����w�'���`'*9������q��}R�h��!�Nio���ܺ|E;1�0pZQ|#�DF��tr?�,�Xl�J����3o�m~���tDv�Mh�����ɺ�vlaG��@zHɨ1%c���EC�xe�����Y��T&xw�9��SP�s��R�X|��j����u�:������m\H!��}?��J��>E�,���;S�8���ӡk�/P�G���� Ɵ�����US��A����h<� YA̕��c|�6ȱ�l��]ST~K:�S������{xwwUQ�s^�����d��O�T`9�fُ����v�~��<�,i�9�ye��_��J4�<zP���j?XS�V��tc�
L����>臡���F��w��$���,��H7���o`��Du6��o4&�])�t[�U�%��â�K��̍��B�(�}���\O�@U6�y�����O��D^�=�jŕ�si;��M~��J=Q�ʼ��\���ܘp��t
��Ȧ- ��tJ��R-cD��U�|]<ɰda(�BJ)=3�I�؞2�K�����PAi���Q�$Ϲ���\�>�N8��c�5��g�A�j�t*�YӖ�Q��!���a����>d����+�Cs����쇾��׼g�fY�e�V�a Ҵ)v-R_6��5�q�l�-�N6�I�2�9�
I��iԉ���ƥ3��W�tv�g�5g����Su����*����[���d��u�����a�书�e�H�}EoE�G��]��"9���n�d��4��T5ú[�~3A�U�k-�������k=������i@�������WKҷOvܰ59o���kf;���Rqh�!�Ӝi9=/ݍ��v�Qvb��?��f��L��x�k>�5GU�z� ��ӟ�����.���̔N�ũx<U%�>�;�\�/)ر��o�ʐq�]��1�qId����P�	��.dʖql䜒���c�7�y�>�s8���P��@s�B��]d�Qht��מ�x�6e�)��Ý��WS���
��H�AI�T���qlu�+`����@!��)��ԂL*\�|?:��t�2��R�5�o�<����*<��h\�{�t�9���]1&4�6�+V�>g�Lt0��ᚇB��%��V�fPQֵ%��I�s�Xm`=`�(^f�����V~�3TK}�~t��b��T��R�	����vx[��T�R�b௸ok�D�3Q�u�}���}ԕa��pFZU����w�������pY�N�:�^K���B��M��ۦ����W�ZP1��Ï�@Z��$��� �R��21f5�Ƅ�|��V��7`p�j�Xo�ԸIdB��;�s������ �	av�kL�x�%�4���Eg�����x��x���p�Y_e����f�H7�\��!�G� �30���Y `T���}<�_P�>r�ߗV�eΖ���2��+��3Zn�$�[���^l��n�������}��铍��<Ϗ1����9���ڄ�h ����:u��؄�QΗR���`,�ğ=<Ce�D���	��^���7<����ZW�#6OQ̀1�v�)�Oy�~��9d����|��6*��&�s��c>;|�y�+2��S�K��Wed���h��ˌ��t�@�y��	�\S|���'TQ�M�C޸x8t�qH_&�%qcO� \0�<7�+�����_���0݆�p�{{�N�R�h��w��}�|����m�d,�����sL<I�6�&ڄ��+�uu��H�.��R��̉��o`�?�̙0�r�rY�H8O��s<�i:'�}fz���>&>��T��+`!�(�t�3i�����?څ�e��Kצ�q*+@w��E�C6�Ω��������g؂�g	-K1�5����W�u��/��v�	�AO#+6#T4OO*�Kw�\q�\t�o3 x�0#=�ZLoH|R�=�dZ�!�Δ��"���˹y�ԩ�>�z:K=p�!d�p�tq��V�C�|��93`�Q4"�8\nb���Yd���L����V��B����ߩUx��VP�f5y=��$Ok\�m)�L�z8'+`�/�}<��X�̀�sc�Z���єH?$t�f�]����+0H��\��Y}��@�ۍ�l��Ou8p#�D����s��6%!�M��w�����yF��BJ�J+��n	��5�a���fa~8a4��~֞e���o�~-��&��ɇD6Qxg,_��ùEGv�A��e�xmQCN8)��d��A�9۽�x�A���e hL1��aF��?S�f�\X����:ȸkZ�	��׍��o�s#�7 �gQh��# �Ok\A�Ԯ��39)�k�[����s���1$FxR̌�s�|`X�@�6?s����u`yt�31o����߿�~\d�lqx��������w�b�1l�B�R��,�%1}�ZS}:�wUc��y��&�AⰚ'�A���\7��૔�%_ԍf	����yj�ck����vc��g!ue��vcj|M��%vs�gA͊���4A���k��Dg�<�o�z����$��}��,�ss������͔ں�,u�:��՘p����/�>m6�14����i\�EL�E0���9j06$p"�*�����#��8�+��M������ت�ى��*��+�ill��h���Mtp�w�aL��3������������7�va3�)��s�`����lW���A������[����.�����@���gq������쎂P��z�f|��?��YOfCs���]\=O'P)�N��"��>��؀�ϹY�*(���E��D񷡞����9-#���QLV��@����k�����ϒ�sR�2ci����v�@yZ�vئ��`�2���^|�z�����N4�@K����GO� ��b�����̍g���K� �ذ�Gs���@;WTaN\��)J�IJ*�d�
��~6��
��T#]��zV��A�%���4)a��{�sM:������.Sa4�:���@�+�O��]���`Q��$�<op�����*�	A���'g�2�B(�pb�᫯�d.����aY�k-����B�2�3�xs!)�$�櫚0�΋ȼBN.��C�� ��?D6���,��/�����Y����^�)NamU�z,46Z=���:���>U%�
�s���E%�Ͷp_7_n��a��_~�%��o%ǃ�G,�������h9����Ad�ܩ�r��6N�a m�,�`Қ?/׼JV.�O�|e�L�����Q��Q��F�+���
��o�����k��~���u�^xvo��A�!����U?�j�<U��Z�,zg�a�jm����-�a:~M���)�i�����\6�D�M�*��I��Y�ml޼~��k�����؁��J/��|)M˄a*>){
�VK�iJ���=a�s�����X�'P̙�8Su.�Ԍ��.�/|��_��nV�Q#*�k��Z��d��/�����7_!��{���5ӥ�I��Pu#���o��vZ�G�%g�%�O��4���^w"_6R�:��������j��ʇ2����*�N��]Z����Y
z$ç�}1���,!)�]Ӕ�u���86�L��������#�n��q�Z��k��g�so�Q ���]<��3��nP��Sg�vI*��k��P�����3�M<��1�3��[��9����7�x�2�f�!,Z�-��,�a�}�ЉCF����lVaTU�􊢴��;�Q��\͜��Y�^�u 0��X8��YS�j��ЄG�v!��Y}ч�~\�2����F'ϴ"nU?U��ke�0yv�X���?^ދ��q�T���?�5�C�T�Y���&��JYf%��q��mq��_�޴M��H�<��F7^"�������3ϼ��F�D�諮��273��@Q��T	@wUVfd�����9�*I��2�����3��+=h�,�tf��qx9�
ㆌ�TT����d���\������AjT�(/u�����������s�繜43E˴�&C���1C�{�@���`lE3e�5�Q$l�a3�OY����y�3Tz��CD�� aT��3R�"f �U�lQ�7+1±��J^�_����H�Ya^����e���snTm'{V�QJ�,����q�ㅍ�g|9��^�����ބ���(K��Tx������v����q�_�Y��c����Ȟ=�
��Ғ�2�/,���)�-|�C�y~�Sx�D�D{���-%�F/�3X�@0Wp�7/n�3���d(�s3h�vS�ʼ���Ȼ���f��x����ja�	" 'ϛ��e�fn6�����ȫf~:�����������Q�uqq]S^���$��ݷe�xëP;��=aMk:(S^:�Z$t�a��<�a�\��^��)q4\��^D�
���_օ�<�<��<1��d�ڙ�u]8�������Y����@q.,���&�J��:�+�-yu�w����FF�&ԳHazF��iCp{�Y�$9��-شBB48k��	��ث�1������9�Z<�vb���uB47�ڰj�;t���
5�10��D	5.nvVe:o���O�A�YȤd��& ��!�|!{*�Q�]��9��/̗���Z%�R-�k��N)�,$#�[u�)(��������9���U��l��$��>!w��W���x*�j�XOF!d�f��\�����TI�J���B+k�*��N��a��C��V�9{�.���P;�����-ͧ���kl]jcI&�b���QlӔ�x�=��[;W-{Ѧ������=��ԥ�|枚��T��4���_�ƅa��H�n�f�e�rF�#[V�������u.4�֡�58����W�aX��p��2�N4��jz�1�o�S�����&%��ū�l+�QL	p���˙���غ�m��C���+o��
O���W�%����f⬲���#d �ք�+�!6M�h���?��fC�[ukdOx�!Rr��Fd�*��!
��b�c�����&�����3ϗɱm|v�尗�
�\:��KY���g˭6�[�%����|������ oG�S�|�Mк��{���'���٦�<���z��˄����!ڥ�Y���>�:�A��!E"'���&0n1����! ��9�0�u6�mϋ7�.:ֵV)`�����û�w3��}S�xP#>2G�C�
�zX$ɗ�p����.�(ŵ]���4+�����.��@̮�\�,f߸p�VL�{�B�!p��)C�z�4�MV����X%��WiR2V���N��:l&R�"鴰�[��v Ī�ڵ�0�� �sb!aA���|G�k�3�e6/��aN��;Uuj�	�w��!)lx���L�	z8��^��gс�k�9�*l	��y��c8��L\�?t���úby�H+d\�:6��	�_PJ�~���uL�2�F�$��X��`��`�34Eql
W�g���Gs�:���h.'\6ROg��ս��R��}z����+�4Ա?X��M�愦H֖�X ��s����ً�'�9p%1�Cx�1���ڪk-6lz/����yn�'A�;��{�L��F��ȶ(BN��nY2D��$�hs��*dS9jf�Y�9��S�s��>!�C�S�l]1)�,�1�:>˔`�)Q�B��m���
�۾,�:��sn �<���8�-nv�8�V'.��zuba�4��X��~�Kc��i���x�����~�E	�ޮ�U�xF�m�E/��$u�Cb��1ZHAn�(l-������}Rg��!&bC��V�!0O�|�3ͪa_�'ɏ�%P���sk_��*�c�Q���>tHI�~������'K�O���u,�ZE��?�׺iʧ����ں��&�i8�z�s
���h;�e�6�"�ҖUG�q�N61L{�c͒E�'�$��t�+k�Rv��'&ux6�� �wֆNf��A�~z�}0 r~��ދ��>M�8f��^����6����������F=0<0�o����n�1���P���]SWT��o(�O/RH��m&�ʒcgE��o}�Ǐ�Vp4J�j?&d;1N�a����)y�I�2�@��vR��J6N�����t����Om�5 V#�q���%�g|��2��	�?�^��9�J]BDz����e霱6�)��M�4v��(|�x���3�X=�6��G�ԩ�'�`�5��i�5�����w{`���z��Y���og��E�푾 JP?��˯�� jQ'��<=�PӋt����#B���U~�!��$	x�����TIA*4�����5�{���0�tg��M�R&��m`�~eY��ҫ�
',Rb�wz���Ԁ�:�f8Al�^]*iy(V��B��ob?���x����P����;�c0�-ϗ�I�N�2s[�eNM��d|��n�ǡ�)�@s����t�ӫ�Gj��E��9��l!f��D�h+�{(C=F��C�/��ۤ犱0���?ܪ)E�y��HY�
�Q��!4��p��F�w�#��O�j�ٿ�	;W�A}f��_�:��js>x}�>�97���I�O��u�"|�L�G"m^B�0�s~����tō
/h0�q���懓M]9�a�Xc;IM�y����<��{���$|{��"�Oڙ����ϡ܉-A6�?|��r����|v��M�!b�N�%<����"����C8�rᛱ.����#N�����@R�!��:=;����h�dIP~��
K	)w	�c%[�opPWrԶsz&.�m��2���0;����uL��Ͳ���d��BV�E�7`���t�m�׺�^��!�'���:�Z�+k��q�QR��7\�y0M�[�
a���a�꦳�7��\�Q�M���B��ѥ�Y����c7
c�M��� <y+R��~�ǵ�,��}N>m�5qJČڶ17���y]$��6vsN���B��
�x}��Y�
q#��?�v,]IC5���|x�� �#�?�y`<�n&�;�cͷ�
��hH�r��ܤp��3��p��=�xƙ�l��]��C�-·9ڭx�Z�i(Ð��i,ٕ�6��]��&��4����"'s��*���gA㨶�j̆D��B����*S��U� �VR�5?�<= '%�Y���k��"���TDb�]\�!�c36y��/v$׉[��b3I�wV� �k�F������z",\��:*W�ǒ����{I�$^�I(�H�_���%f'R�ŭ�t#��� �Whª'�0�����7���ز�ay\��-'�BS��c{���p�,�Ɇ�zI���q٘o�$"! &B�[W�jQ��阚��!��a�0t��N�lܣ�֯_�$�4��T�Z��&�B����9�9���}y���|���/J���Fϡ�e��&dU9�S�qE(}�"#~?w:���\�qu�M����?�K	�Y��
lv�VЂ،9�T��⊠F�CN�E�6'�Ӽ�$.�؈�F�a'�¨��Έ����D��F��	��+�=f�Ž��j�qAGؠ,�hŬ�bf�^D��[��d,?��~��?P_�#�\/����CR����{P�}� <���������F��u���1J�v���}�8!w+x�]f����C+��qg���l���>k�h�����j�48ie#��=�~�����x��
�ii/~9��$N61�m! ��F�o"�����������ڐb1�ر��m6������;D�z)����Ƭ(�}҆��{s�p��@�Os�ڑ&MG6�y���l�J�'�����C�=�C��>���X$��Lzα������4�����GxH���`�+���z7�k��O�G|6�~6��Mr�!��.�����U[�V|�8��J��hI�X����am�)���!��3oŶ����K@�}L��F^3��P?�j#��H�w��{�_ڈ^4�!Ǹ�*���! �>���1"�\WL�cӗ���<�Ļazx̸&~<˓ۋ��
�ssK*��E��k��ٷ����F/y��B�R*��7��$CO���$Ey'&�f��ʁ[I�s����",hA*�.��;������G�p{��/{ʘf4湧�}xq0"�e�)� J	�8IԮu��
�E�"��7A�Z:�=�����=���?�9��KB�4���R��4�r+%a<iH���U�8���������ur-<Ү������(o�xF�Bf=��|L�',p�0��RD¸�����a�J�'��,-���ƽW칅g�(;�l���(��MY�{悥�u��c�㧸6<���{��FLx ����󰷇�����K.x�8��M�]r:q_$g6̻�[��4#e��8lwF�%�Gy��H9o�p���ԵC�Z�����^%eɞ�<7�B鵄pD�_^�/�{�x�~��X�Dt�����`%{�}_�\�\��ց��g�������-�c��V��M�\�]�D�z���(�����:|ZjE��^p�{ka����`���t|�}ӟ~ǉ�Y���fV4��H�����<��3~tƬ�_4��b۳͒?%~����P+#�����bW}|���J���I_���}�u��lw�����/����p����Bn0\0NAΎʭ��2n�&W��Q@�#U��� ���_�3�Q��^�w��1�w�U�կr���$ak��x���K�tH���f��;5�;�~'��j�#���}nL�|[舙hOp&�h��ś�S\��^[��:�}��p�Z�^�z�s��8�Ɇu��3�#�����B0��tD�z��q�F��g0�Pu�H�s���|nx��y$,�|���"�����6���
��3[���s��3�p��i��y�}�)kM�ڜ6��Y��J�Ig�C~�xPB����N��M��s�7>�v}�	�(�ё��
�	�k����L���>Wb��p�]��ui�)�gt�DD!X�
\�������ipNx���e��?����S��#K���#)+
�u$����0t��.�,��Y'_�^Pi<]%^L
��T�~l�l��0�_[\X��=��H1���� ��+g���Y]�oC�Y��<PS� �{d4�
��5ٸ~,60��޿̾;���8�}r*��y��Y�ܧ �cr���w�V�_U�����ۑWiO�"�̺�MR�p8:��!e�z�6H.�Ov��s��(�8��A<c\?�@�p�0�Ѹ��N�7������p��y��qk&��>�u�y��q��[7:��pٔ��*Mo9-\t���L(vjW��}��=�e����?f���-E\��m�k$A�
�s7�{c����7�>��t�X��S�xb���Z# ǋkJ�1��O*� ��x���d��T&#�����i;ȟ�j�<��>X8�29zҜ���f���t��t�L�C�S8�O�F߽��Y
0��xi��_�5��B��iH?�%�YW�ᬋ�iR�"2d�@�n�ޛ��^0�l�J��.�/�6���|6T�م���7����ɥ�!�ǈ�@�ʿ�뿖����H��w�zo
���燞'<�*B<�mh`HY�|��(-���v&�s7��s�/�8����?���.�c�,���Yp<k�V��[���Þ�O�
�>EΞې:�7�a-Bǚ���!5P�hV&�;��	�)6��ۘ0>�0���q#ևMx���_"�v�Fa�����T
������%ädU!�^�0��-���0h�!�|c���D��o�(JR�~�m��w4����`٬�x�k�k� �������>K5#d.E])������ex֧Iz���	����B-Cl�Y0�;fy�N�u��W������J��Y�4f�;�:�3��%E���Z�Z�d F�O���gF�Q�J�+q��ݻERSus�h}�,��.g�iHO�4���{�<�_�C�����f�M�n���-3e�wp	+u�Z��풡��n���G5��\m]�=���:P����r���,�v�+���XE�q%S��ј?==�'�ٛ��!1����.R�rxd�'�����>����@!�R4�L��g�o%�8Vs��9�������+����ů��'s�g�R�H*	����4�e���.���R&�o�#~�"�lV8�^�}lf,~X%���a<
qPZ�6ϕ��)u$��γZY�5=�،ѓ���j�0ޞZ���)�'��ߵd��T)�����k$s�@�EGu��n��.�&�w3��Y�kVߊRAd�*�]b��	!W��eC�r��9�ÛH��9�ZxO9��C���$������ؑ=ĂB���f�Y�]���k��?:�i�t}�M���j��bs��wŨ�_[����Z�̒K���ͼ5_G�9w؍A��Kd4���J��^�?���p�����N�VIQbjOV�ƌ8�V7�<��BɢPY��k��Hz��~{#�T��>����#�2�O��p�mL$�S1T��Xôf�9Fx^��k�n+��6GiJ�Au��7��U�8��]>�r�x�m�6�΂�"���-���ׯc��0��.���`H��ѕYg\�FtYx����]�04�p��GUU��&�����#��E.��Ԧa�ƀ�Vv ���[���Y��Uy�6�}�i�pe�BS��1>_�1Ⱦv��N�\�Qt���Oɓ���AB��C�z���8>j�����<��HkC
j`(��Q�Wz3e_�57G9�O�xZ�Kb[N�I-s��u�Jgx���6�I�`�x#�dk�:�(R ������{�Y��Y�4���y��]�Ǉ��E��zld���b���8��8���0}Av߻��a���'�hX����� w�=3��)C��<9\�C�׀�~�؄3�!X�]:	���Cx�H
�8ؔh�q^x��_�ބ�|���Kb�y�E(O����>>�H�\�K:>M�؋D)+6( a��wxn�;�㐆Tp�F�W��s���j=���W=�y��Pa����*:�J���uL)��18��G��w��}��> �"[m���3���9������x$^ѽ��e�>��"TuB0���
�Ϛxl�L�n�x�^	ZYe�?W3�V��s⩧�����UHC�7�j1�5�������b� Opb�ھߗ,�h�7ʀ��#9%6��3��-Pw��4'%�R����;ʐҋ��#�P�@ϯ�J�ׂ�V븁Dq�iD�}n�Q ��ĵ�(���������}��Ҩ�U_����v�	�Z����qK<���ڒ�S	M�!����/�M�{L.jY2tv��:7sy$^Ȱ�C�,�y���ق�����G������TF�u�ᑞ���'�`cpx���pzw�H��[� %�u�S�1�������S��IM���)[�Pq�}�F�^��|E��L.\����j�	:��A�<Ր������%��?i�U��'9�,��i��+�f��5i:�� lT�/��^���:��e�L��ފ�{wR��O���u��M��{x�a�T����I��XZU�Y"��ͺV5��4w�E�vA�W��a���6��m���ʢ:�1�K�Q�|��v=p|���H̬�1�����u�n�HbEj����0y�� �
�M�Q����k���%%�,W�W-��s�7��N�NԿ��8^v�G�4e���e�S��吶I�6�?�V���Ϥ?�hN2�j��R��(\[�vN���ߊ�K!Ȕ#����5$�vl�l�+��K�$�f�h�BayQ���6���~�m����j����
s0�Za@۫�e��9�'MP1p��1���'���vL��(��+��r���4���3�X�5����&�N'�mc!	�
a�j�&(����:���MlŽ��v-mB��O������_��Q��S$jH��(Q������e�&���$ի:�43�}&����8�C2"K
��-K�u�'�H΁alLp>$��+��	�Q|S^'�w=����!��Ƙq��gG���g{ޘ��Jؠ7�����7��>_�/1n���u�#�j�={�A�R+h�=���G����>$w�7obְfD���&�_���Y�	B��S�#��;e���Ny��qp��jdwS� �����UHy�=ϸҰ6�i�觎�H�Z�̈������J�h'�C��^)xB�|Y�*/��Q��Jmy�څ�$i;F��N���	��N�=����Q�6V!����ݜ����.��@�p&q�O/��M��t)��O���ł�F��� cf��D���|N�uqia/��j�R��k��ժ�)��������*�ɞE������Sd�7�,ܐ�^���8w4������ ��b!�e���MUו	�ƻ	��H�&,̱�@ϋ�4�)a��rx��^1O��٫2성b�8z���%��(|<G<�,��L��v�+�]0|�bH<ֲ�0�6��D*Y�غ�8��"�l�Ĩ|h^8��0�N���0P#A��Y�F�ȣ��(����{�a��Ο�q�7Y[�����W��P%����%��!�����Y�f�Q����vS�U���D���))N�M0Ֆ6A���D�f���"�vYj{��!����i�@b:V#ڥ�l�#&�� ��{���-L	��m��T��+_d���Ζ�,�"cy���9]�y���6����I�QwJw�ă =ɭ]�W�M��l\��r;Ff4�qېz��l��������0�`Hc-K�S*���;>�	��K������m��SLث�N
N�!������|�<����:�(��F=�ߖ_�%ƚe��u��jH��}80ׯ��*
~��m<;?��6&�~R����n�
�0O��������"׻G+�ǧ�.tF�z��H�ʻ�:�+�(,}�ถu��3�1�eI��G]�e�x~�N��W݋���T���W�?'x�_��B'y�e�G74
��MF�A�M�����Z�;�%1v�"#�S�1�*\�  ��IDAT�#|T��4<+��_[\y͒W�p:�N����b-����<��y�'���>i>c,\�����,K�d(c#:/<R�����#e�ܗ��Q�z
OUw��F/��=�0��6�ւZ�T��E���h��܁�	�� 5a�6�E�uYc$X���{��M��d��<�m�����2[�!�!��UM�.N�6��S��(Ʉ�r�I�;d�6��������$���;6�,)�+ZI82�Y{_��t�fi��@���O���W}�v�Gy�6J~lb1Z�!����̎�S� _�W���X����e�xƥK�<�ua�Ӱ�D�t�!b�W5�h�cx�������^�&�$�l1��$yF
>�+�p�.ѨP���7Z/j��0rY�=�<iE�w��/�������j,n��띗ZU��Zk~�*��ߍ�&5�2���.K^�8r��u��$����2*�kDv=_�[Fc@�i��s��49��x�Mh�MᬌL�S�S�ޙ�Ec�h�k����kz���.�e���~�;�kQ�ep�Â�@����1�s�ȝff�fo��Y.�;.P�������Z�ϐ/kh*���g���Վn:�:/U@b����+F�/mc7L(B��ɲd��j�9�ٓG����>Cu|tY-�=w�u����{��<��1�n
��?x롶1������I�	Oq���
*G�!rB2����>F�ޠ9��6.fɍ�Z��V������ўm1���Ќ�������h1���K��kR;�Y��'{G$m��ɶ������C@�w���ï�c��9�Q��"�/�|Y^�=A$�0�U��$���R=$'���ê�>�~�8�LC8�n���p�y^���? �d�����"�^��<e	�F����'�	N��?�ujS@d��׫���"�Y�]UeƭV�Xg;m��h!���N8�N�U��.�=	�*/�5g6r#{3�'G����������6�ɡ�fxN�,�4Fq<VQ�")8��b����}_�wm�ZN�)<J�'��W������r��ަ`�_�5��N!���Jf��6~k����NaP۲L{eX4nǲ>f�Y�x��^��rEQ���n�ʄZ	
T����~'�VÐF�z�a!�rȅن�T���И�ziT��K-`܎����lWV���}��!�B5����,~<��s39-�aoƙ����)r��֙@���1��S��o8DS^F;����+�j��",3�Ė�w�%�x��1���M���/���u�3;9����S���1��x�==H���JT/)�s��ج߫·y���D�������1����؜8�NX�y��}��J�eͱv1�O�vjn9;V|-j�E ��P�vP�L�(�e����?��Y�ȕ�7�ƈ�����[��:[Q��(f�	6�k��߅��O�'�������x�wu���E8n6�����bń^��\�J>��x<{ gån����M���A|����㨕9��[q��V��D��i�;"��W���&j��m�b���A0�[P�־S���=���&���pʼ[O ^M��+t�(ٻT�
�.p�_~��E�$4"L�G�ؐ.)H-֛0�7���m��1��q�&f���y� T�m���&ww�d��*�
/g���OE��H��X8�
x�G7_S՛���[8����o���÷�r7���Y��::���g���S>�AIU+tv�,�����^��l�����p6�>���2��S��-�=��p�����M���^�Zwj��SSAl�ߤ 8˯{)��>c�\�s��T��Gm��h��LVA	�9v�H0�P�������V
b�E��'�qH��W���Ԉ�j�@��8��b��\��F�0����g����1����1�=Y���0�cN��y��>�hJ �|GNx#n�Pq�)@_,ĖZ���[����𐱣�/]RS��D��#
I	5�3�������~�L`�r�Ȉ��	���Q���̥g�Z�Q�h�{o��7gbI��FK؄]{y��.��,� �e���Xi�`�1����0�-�߯r�p�sxH��{Q��$�QY%��Js�Df�|�~�8������u��m���!?��[wq.|�5^�h��E�j�K��C̛��l|�W��z{6�f8D��Se��Ð�yo޼JJY��n�L�M��Bf�	�E��:ot��P�A�,�8J�f9����q�ដb�w�6������&������^��Ý�ga�9���K�2ꤡ�7�$�I�9�b?6b@(+o��r +9,�� ����D"|m�}h����� \8��_c����-�$�+:4N���L�j#��1m����G{H$�爨�R���ܠ��!���]\�J�W��h�Ti���{���x)���vN|����G��jw���]mGڄ�b��Е�����/�oc�-ὓ��k���z� �-ͅ���ED�$�����(&�[	lDE�L�4{ۭb��H�fޞ��� �H�F=z,�f%xf�+3<]�ӖI��^7
ZS�5([��zm����$�&oj�D{��5�n�xL�%UM�ON��tX�(�Uxn��'6¡�K��c	R�3� �ީ�5�C��v{��aH7*���}O�lH������ta7g�Y;ǂ�^l��4)=���׆��g�T[����������^eE9B�c�R�ׅ��wGO��:�+�z]d�#k}w/j[~�gI��MR�T��T�੧c�
�Oz��ӄ9t:f�,�n43=ϣt}O�a�G͕ʕ���#�y�N���>��]kA3�� 1�Y�)ְ)bv H�B��ӺT"Rς���<�rD������{���e�nb����=#�V��<��}l +m�ﶎ��͢��=�Ih��Z��q�/�⬽���ih	J�/xqWal����� <H��\f���I ���7�D�s�2h�oq�K>�e��<��φ�ݯ��#J'��]����/�F�t�Z�ͷ���(�S�7x7m��:�xO������x{}6lq���!l�Hx��=�p��Ja6��؞����&<I&WN�}p������[��0�!*�wՉ��L�mE��B
C
oH����I���c��?��H]�����
�N8^�_"�q>���/I�:A�b#|?|lc��p���U3= �$y�;$����O�^�Rj�`�5<�ׯh\#4�R�}΁��6��B	b����1�����J��z!��	9����H�T�q�k���k�:= ���w2js<P�&%�NMa=!yd��KL�t��q���HO߷Y�@��������Y&����]Ipg,)�ͅg�n�8��Xv1��agC���iO�<�k*ʕ��֨�9�!#\+���{�}b�޾
|�p��eAh�Y�G�𮧽).���3�Y�"����s���;���_6�'c�a�N,w[z��W,BX�*�4��׻�w����p ���~�79gX:��^���N���9CTa"v�l�p��j�M���Q!z��W���A}�3�����5�>V�������B��ߵ��ko��ʹ�$�G/�/K�\1U��g�)p�&�Imp-�+��
����J��I����X�T��0�I���TQ�Q��UO�}��ە�*[�Ӡ
1^;9ʆ̿$�Uk�-�����^+�K�6¹��	JV0U,7*b���{z����<`-+���ی��}3W_]�x�A�7����s�>�a�s�)GS:5���I�%7Y������W�{z�-���h^9,V��^4w�\ys�s���!�m�mg'�mEe8&M0�R�J&�;���Z^S4zJH��˸�g�o;U����F�S�=j��3�ȯJ:W/�΢�T2~c��x!��˗��N�"��<�����}����QC�i�\r��0Z__�4^���Z��AF�����9L���S��D�MC��4�ßib]��9�w6�Q�¹i���W2����%JH�<�$��A*0�̬�+��$�a�	0��+U'�����)��l4f_�/���g5�vJX��2�A�JB���$������N��ǆa����> xmG��z����E�J���b�����]�o»��E�OlN�1�Saˉ����]�C�1h�T�I��]�U}��<�	Qa��[K��V�3���kh�[\��1��+��.>gXƟ�3`, ����9.�ʫ��fo�j��9���ڃ��=�����%�c����t� �.�l����yc��oazw�]�����,xbE���H:ME�5��s�,�_�ò�������Z��??�g�c|,�ec�z�ܪ\2f����H@�E�&oq/�����^�Տ�t�y�}���
z0�hP%A�]y�E�p�IJ
�[]E2��UTX#��K%=��m��ڿw%���������s�*%�5�\4R��{��2�L�u�����Y!��
��]��=dE��_����taHݣ�5��Ɏ����=����z����n��>�b� �y��U�����	È�8^I	��,���s%6�V���N,�jo,�R�viǟ�^�~�&�^?�Ա˞R��=Hպ�������G)�՚}y����{B=���)�C�f��Y�,�xА��'��b���7�!;EL�̆x,"�'r]�e62�W�*�h"�S�	���I8;me"�JO�nDd[F0�Nb����ؗJ_�N�#)�7:�'��W�O/Z#�c4�ѧ!�bsws�h�x�}��A_{6�d�-X)�u8gN�9:y���[�����ː޲]A���4������ ��#= Jˁ�y�1OO����r"���|
=��ߩmn����q��2��D���gA	��r��Ԣ�����?M$�pf�C�˪�Z���+��n+o��*�)�u`򀒴��m(���7a\p�H�g↳�� ��W��*V�f�:�?{�meӤ�k�ժ�|.7ě�)iR�Ԯ�.�mȽņ����/�f��,�<KB�3q��Nm���y���]�fs������Ɯ�@�Ø���@�����G@d��e��.��wL<�,�gJ#���v���G4��׫vQ%�6G5�c��5�wV=6�ۆ'��8QG֟qT6T6~2cf�ɘ�z#-[&�!�RXB4�Ԟ�'=������F�B
�l4��4�Ϲ�srq�ui��-\��x���)a.b�N�	H	��t_�r^��-X&�G�A��������֘~�0\�w|�gS�f#|iփ7Qgv�;��xK�2<웋�␺ �t�:똸%���~�	��AA��\Ðx��hO`���)�����Fa�v�s���2���x�i2&y���+u�r^�eNo���W�\�%��ߩ��	��{U�P��2h�%VJ��c�	�_�8	*3�P&n*�m��7&�2��D�seuǈ���R�k���c���;q�8���?�
Uj]
�HC^�y`P���?������a�&n�o��{l��D��\��\�׬E�WBԪ���흈��D#a��k,�A����3���ae�6g��z���n�����*�@(̽�J~߾ߧGm��k��5�B�)�xR�P��6�V\r,�[ZJ��3L��t��q�Z'�`�n�)"����L�a��[m:q��~���Ԉ�o2W�k����Y�]�Q�F�+A����z�X�]�(v�x��)ۆ�Nb0�̲�^�� ٢�"�PsS]�!��V3�Q�p�J�V�yjTV������Y;sW}m��))�6��n�㞽����:ra��j����J1�~���^�8V�g��僾lU�Tg\e��DlS�[��u�a���Uj�����a�w�Y2�$�R�����t.>�d*r8�S��Fh��:ذq�#�~ ?rTr�%���X�U�K��?�;$?��x��AX�A&I��~��&����-a�Pܯ����1|h^D��[I�H,{� ��z(��+$6��1�BX�[� ��j,�f%�v����h�`�vsu��Ҩ���T�����е�u�����u%J[x��ǅ׾<tKB`�w�� ��$�А���Q��^�e�x)�f��{^=e�)oSHi-=�9�	C Q�)� �����u�^��FR�,?�~ʈ�}������1�?aF/iQ��L�Pۍ�wq8d�8为�J��!�f5%R����6pV� ����CL�t�� �uJ�]�*�G|��`!`�ms6��B�ºU�i���h����܃�=��Jڟ�I�9WV�?�����08�X\ ���:�����7�������J�"�u�Q����OC�L=VnJ����i����\��v�(�q��U�=7���!u���aCꌆւ�H���{�Q9�og���r'P���00���"<F���$�*�Y<?%�`,�%x߻��v���nH�}�M	O;.��66ni!��n�#"%u�E��iO�s�߁���O?�����(\������u9��G۞�6����raQC9Idz ��E|ǩ#%u�Z��5o�6,���w���ĵ���u)�l��{-6�1DV�q=+�T=O��q�wmD�ɺ���?�So����PȿTL�G8�1���b�ن,2p�"MD���1)�N˹��M=E���bu ÏʲZ�
�xH��O�^Xd.���je �xw]���iǝ�u���#���ޒrR��j�Љ�B�7����
���1靭v���!��4�C}�
y<��%&(�D�~S�94^'���cq�PЧ�(=�`91�g"�Ԫ�4A*^���p�JDo��ÆP���(O,td�^p�����	�M��=��-7s[C�ß�:#N��xA/���+���=#F:0�����@j�����T"jQ��u��"W�ƀ���y�߅��5w������2��z��?�JYt��?��tkAN�4<Zܳj�h�3/1T�)
W�>�1�����3���T�N�j�\Ga[:u
h��}N��s�G�"����!����ɠ�aχ�b�*Aw^o��4UN���{aJu��.��W_h~�"1�������� 	�2e�2��+«����ċ����i������K4e���a�%��jA�+x@��}��mϵڬ{�_Lrx1�$r&t6X?|�cx~~��d�Ub|���㝌�cY߹b;���=&D#���UJ�n�����	���%B-C�1�uC ���X���Rc�M�O�8rGV�=7��mFW�����3?��S�ن�F�P#K~�Q��B��P
�!H�iι�bR>
4���J�>i_gX���]_��"��A�w���lz�����>Y��lr�69 
��2��)��R��gEa�L��d�萅0��@☞�U
��;C�T�P�;�[�؅Wy<d�u`�á��7U�s�c�Q�BB3���x��X\,�chì\jU{��~p��cG�m+I-%��1�����O��S�~~���M��`�4DU���ou�"+Cٖk�Þ�[2`���}Ho����#TB��X 0L/ϓ��o�_��/!�*�_�=��۳�6U���D�;y��^�̰�*8G�D0i>d����\jH����s�� ��U*���8�7j�^B�d_���sx�_��Z~�����/�J�X|�8����h*�T��[��ܪ^�ի7g��FE��e��!��Qy��N8D5�X<l �7�$Q�f=��'�&N���f��sa7X�	��z��eN]�ˉo=Tl,���Y|S��=�y#�i����x2�D��/�=�Â����'6�����0�0��}WWM&d�,"�X��h�(m���\=|>��ꈾ�Q��g�09&W�B�rr�qu�_@�p�I���A��f�ͪߚ{��xV�?=��:UN�Z9�(ȗ�)^��=�G�J�L��z�k�Π4��.����|���"����:6���f,�?� hs4ϓM������-��Y�Fk�掰��vc<4�٪{;���8� �-��&כ���ӟ������(�q����&��	���R�wP���*!O�
(�_˜'*u�қ��Ğ�)O�J�h��SU��y������˯�~p�,�J���?�!�=�V|]X�6�!�U�lo�=��{�����P�w�(j/'�����.��v�%�^��p��,�wYj��j8��j(H���kzb�a�����⋒�����Bs�	c�^��*3��*QF�P�е�^�'�S���Jd���#\�(J��}?�ǚ�o��N��y������%����}`�����Od���&�r��7�����@�UĢ��ŒS�hJt5V|��I�����0k���
��êO�B�xHƁ:���XK'hq;d��H����e����PW`�	�8b����6����n��#*/:\at.9z��Kבk �6ڧ-���u��co��������1��ͻ˒ڤ��E&�S��+���#v�S���tl��G		D���0Qs��΂+�a �dT�C�)x��6��p]�_\�3���:H�xR�zj2J2���Ҁk)S���F�jN!4�ݑ;/{R���)N�P�7���(���%<=SU�{��.R���N�X�>K�I�̳�o��g������gV��$v��/+}x�x^�.x�~/%=Y��F(�D���+���B�8n2�>Ӷ-1$�W=C-ЪV-˒���P	���Jn�}@�����}�z�i�ʠZl���g����k3LЋd�g4��u=|@<�k�WH�`�㑡1��OU<�fp��=��K�H|�h
R���O��3�����ؿ��)�n�8!�t:RM?��?f% �hb�Ɋ�	���z��;�*:��d�^��wj�'��&XC:R�-�<U��G��ڕ,,
oX	U�x����?{t�	}�1ӵ��}��rQ�խaY>�^9R���,w\��%�յ�{���t>��8��˕BAh?�?2��8E��{�i�1��B"��)�c&Ƌ��*5K,$�p�4���7�R�)�a��ٮ7i��Y���"S�'�W|p�)~�\�gQ	*���0K���>�Y�0��*(��b��҆�<������`D�k5�^�Crc�Ɉ�k�%�h�⅊4RwWXH=�p���~�-Zͱ��%_�z#��?��+y��>�0�]b���Aߒ�6��wL����dV�ͺ.�fw��køU���+җ=Sc����(rs�P�=�a��?U|��~W;9Z�*��ȕR�GzL��j�&��{SݘD;%�MK�g-J�zw���:�%(������J7�D��f&�"��:f��v�vPu���:�� ѐ���8|ɋ�<�,��x��
�����طj��ğ��E���A�v��S��}����4�Y� ����AȐ�/i����Q�<R�BaJ8�I�_r��.CZJ��孄��nČ{��~�wUm>��¨Vj}%��C&T��6'aH;?X�tSb�6���	q���A'��D��uŤ��B�^6�d�A�k�"n�!����% ���	�LM��j�.Ѥ��O<t��C�a$6��i� ���ÏaHq�֗�^�jl�	ho/�=�[@М�+ M�U������!�`;Q�6���:<��Xy��z�QJ*�)l��:�[X��LR����DH?�.�Wm�Z�JR�Ϫ��z����mt����z���gjUFG��#���9���_5,�h��jۍ �Kb���lq�h�B��b.����u3B%-��V�V�U�}:;l�qG."���yL�u͛�Yۋ;��bq���)�#��52�g_���sU�|iغdYl�ѻ�Y����8��r>�ի��\Ҡ.<��7@ՖU��J3�N���>e�(tb259��IV'W���@��M�l�YB��Wz�MB$��WמRo� �ը���cw�'x�I^{!����wl���;j��IƦ@�`q��jm��T�$R���ך��mP\�	l�ݴ,�k��/Ta�W�E��H�D�<�����.i�f*'��������Э� ��8Z��Y�V �dXUi+m�'5js�N�"ʉ��&N�1v�O�Ns��i����4pc�5�gO�m4���.u>c��[k��qs�LY������_-�go޲W��{�r��U8VQ��{瘙RD��j j�4_�0�!V���R�T?U5,G�lO稗A��?�@;�<+��OT��ss��E��f�	�2��B<��wh��>3�%�j)õR1m-v����/��˄�?����_��$T�M�d�n��-i�����b�|���͝����lY��fi��c��P��+��`����	�?pX�$ȓ��"0��f���RK�ξ� �튻.�)�{v�^�-t���	cm]4/���wV(c����>G�����fN��]`�F�7�o@2���< j����^����ȋd#�	B�	�N��1��mx�䫂�c�d�����Z�w��܆���n��nj���ޟ�E/��ۓ������Ǭ����]���}��#F�<U<]s�2~nx7J���+��]�MH�/9.������@ev�3�ctr�5��hP�������J7Jn������0�!C��P�T"f�ip�u�
Ǿ�q��09�}�37�=ΆÀ�}R�0A�k����e�_����g+�b�c���3��]�麓q����/�ѕ:��x��:?��s�5���������S��<	*^x$ލ����d�(#4�z��O=�uKf�X$�F_��X,*Ró)���!�g��mkHC}�<���ؔ'-�Nٵ1&ZYJ��);�+_~�%��KV�����Ґ��aR;�9H�Z�>�$& D�q��)�r�>J7af���k��6ɡulf�o�S���t2`�?��s�����!�� j�	,Ӝ0aM�!f�<�Bڮ�w�F�D�p� ��1Rh�H�<�)0ޢyG�@ߧ1u/=��_�^L�����
V,�vXLL�z\d��ac������%���ۮ���2�hpna4����+AmB�S؞�����L��C�Y�ǭ�p�w������P+�0�'�`�u<�6*�(ƛ�=K\�%nCR�b�T���2��X��H�F���� �m����ƕ]YG��Q�yP[��i��&��X��a9ϓ�z�n.�(9������s���c�JT��{��$���G*�k�.քqL&�٩<�I/~���d�&��b��	�F�u���8v�ISJ���W�r������Z�*��+�J�i�P/6���L�y��P��k�M���Ťps��o0\��=>��8��wY��hQ<*Q�!u?�Y�?����] ޸e[�mo���!�p�&�.�-���p����5�۵�=�>)>��������8C\�l�V
Y�&N�&���u�
���5����k�]�9�%������a�c^`�Y+)HZ�-:�̚��1w��b� '���v&0��]p�b��̚^��j��/Ƅ7e����ɪ��˵�QX1Z���bݸnY�����:�~���7���qxNm�9D��I�,4j�B��{�ӄ�vZ��O�c��F-�T��1�%�z|�z��(۞M8b<{ZϷ�/M5��]S��Ŧ�n����-|������ր������%v�נ��ؗ�q�2 ��^ ��{69�Â}{^�V��FWȌ+���g�6�&8��i�,�((I�~�^<�c$>����q=��2��p�e�ɐI��L,d�
����b�k�^���F=�4� 2�0��n�|h1�j�aD<�]��K��G�7q &�t_�a��9�ڂ��n�.юE���]���3�^هl�WڊB(�m���]��`6l����	I�~h��Z&�{TLysa ��e�e��"x��䢂S<�h�|������
g���a��?W�@���unzl��.=� q~g���ܨͧ��;i&t�^�d�A-�Ik�,�����veу�:0��/l���@ ���J@T�¡S!������8��D^8�� J���{]zf!6��D���*b��X.�Z��T-mq��V�]���Z�*��f��+5��>�]&}Qn]*�9�Կ7^�9|鑦�O-�m.���"�&���^�]���ʣL�|C�6�!&1fCWJ���?��5�/��>�iý�!}�6�W�'���rt��#*>6��1�`̉_|�D��	I.������$�*M�υ`�����:͒�P�u^_3��%���F��ޑ����&��	�����<)`Ha\.�р��]a��$f��dޥ1�i}�K	���A��u�s��:%��V��Q��SŊIzw
�&.���� �S�����w�}�{y��:H|��h���"Ď��ń�Qz��7��ECU������:��3Q�U����<!�׵������v
�Ǳv�!_��b*�.=�w.�鬀��٫4� ���\I��l�,�(��z��N�̂Ȩ��OCJ~rm����(�r�z�Pdg3Q��sB�]QݰnJX.��.7�e��H��la�y�3���\b���Y�*�j�>��(�����@h�؝����DH����yW~���^F�/�?���"�K�6b?���!(C�O�%"GB�mf�¨���(�0G��:��\{o��U�H��aD�6PM��W	���a�!��]�=���U��<��8����=��u�^�������<f��a����9�C`c-^\]䤋���"NLxӬ5ˮ�c�̗���w�V4��v�1&�8n�=�QO���0;#��ڱ�~��ʟ����/�����ߟ����%j�D��-��ya._ebf�9��687�mO��W���7�kH~Y�X�9'<��:T�B��X�qj�Ԑ窱�6i�(+ׇ��?yУ��E�k�cw"�Џ_��C�ψ&X߿.�Qg�#K3K|�N�-Rji�Q� ���!�?h�j�QUB{̜��-�5�;��X��s����pi�z�v�@�ȱ��'�~˘ڑĿ��xn�iHm,kVIF�|��c��Y80j�;y�s�9I�ng>(5YN<kTH?K���_��؋��]�.�;ӫux:��P���,l~�
6�-��p8
;�'d̀�锕@�-��Φ���c�x1�l[H��|�S11܀����*<������ۼ�mtZ#\�ï=)-��q�>�GW1&�z�6��R[cL�x>��&�&��Z��;�9�$u�T������ ޤKR׫J-�r�qx\#6��~$mM��FԼM#w��w�1g7�u���d�1`��lI��S&jB�wm���Z���0��0dnC~{�u>��1�����8gx[� �4���5d���DQ'��T���rׄ�t\��a9�+
B�e���i�ޚ����z���\�0iL�3g�m��cj(16��ѝ7ݒƽ��I�����fz�u��j�����9#<m���w�G���I7�X ����Tt�Ĝ�9,UV�J��MOJ �Yx����Z;��$�-��`�Vg\I5�e��x`7L'�Ԗē���ڄF����]0Bal�^QG�l;��C��<�NG�2���6t��á&S<Y\mj�CM��Q���>�cA#���~��5���9�4P-�����<`D��@��Ľ*�XŜ�.<_z�OO�������!q&uJW����d��5n؊WT����&y���2$��>>=�����My�S.F㌭�8�}�L�ʬ�7ShlD)&��U���û���%���@��Rb���MR�t_7��s���)N-�cQJn
�Tɏ���V�Hr��c���� kh�荺?(�D��]#����\F�tvl�F�,ʹ�R�L��
z�u�5�^�,�3Ų�Z��5v�1�=���Ο-�8���G�Cy�������/�!59��@o��3��%�kV�`p\�B����c*t�}I���䬊0L�G�H�7łR��4R��؈�	�,4Z;�p��c��Oj�<w��s�-ʱ�l|đGz��&�צ⚵�o����S!���s$[�\���}
�.�"��s�q�΍�]AYx6P��Y>0�	d~�"얆Ø���hS8��|�a�e�M�m�}�0�51����cR}���"	ջXO�L6���P���.� �'�yK�!h��ύ)�Cͥ��(LI��x�M���v%��N��`�IX�4m�Kr�������P�W[�͈��&>g�P�H���4E�Պad���3��K���N�l��f׆��MF7�w�JG*��<���:[�x�Ш^�~��+���B��g쀾���{[��)C�)c��7�l>J6�*'[��R��8ln�U���n��s	����Q;4��м�p�T
� Y�\x�7��c}������ L�$)/�ΞH2���#�0�q�P��Li"p���^�d�eV�t��Ŀwݓ@C���>~�@ӱ�cK�7O0�)�{1��az}��0�I�P;�O|�S�k�,�j�%�[��wݳ!o�mi\К����5n�w�Ħ'Po���eN�]9[>�P���8�����P)�g�89�[_TY�8��·M�B3��)�}�=��s.~|���cvZp�i�Cw*�e�͹u3���$˨IۧQ�<h�]��߻���a��������yΖ���jIcc��I����N�#�m�`Za�Jw��h���f�KfP˚�gZ�;\��0`.i��
8MtL'�tݳ��L��kD�Aȏ����S������E>���t����槉�����b�NY���+�H^wC�X\'�����Ʈa��[ɼ�㸻{�J�&�d��V(0NXP�
�7��Nl��#�d�S'n��WL$��A+j���h-�����k��n>����g!�$�9<�q]�����*���>���������RJ����k%%#���<�ΕB9c���'�ŕ)4�g�>U~��3���B����	*� �dfx�l}vYq��8�S�\؄����8Ϥ��s�w��{��c�=�K'�~�)!"�NDW�n��!�A��rb�������>NI;k���^�!�!�k[�Do��N�� s�4!\4Hv��!�ә���^�6l�1�`r�EM��ԧ`UݦX��etNl6J�	m�Ĉ��ƚ[��]UI$��!!3��֟�%;���jO�y���[�:~a�筗�b��1��.x��9�&)`:�'v�����U�Y:�!r��u����d��T<:�E�?��hMA��jCi0��B��u�y��� ��"t/�Eą������cx.m�����5АSOs�x�v�
����XO����U��%�����i8�%�V��[�Tȷpnbbh[|6��AõP�������4�NT7�;ȣ��$�T����(W%��)$�,TL�k-����C�c`ڛ�=�>cc��<6�s��Mm��h�Rv��gV�{��\���抱a�����w)F�4�ږ�C�[�����6�e��.V���5�W;��	={{�^S6��v-�c��?��� ��:����R�xļ&�3�)ӐVV����ۂLUK��e�JW1kϝ`H��m?�Dx�R�7���B:�$ �?ƒ�+a�}��R0Ț�Mɧ��Z�2���EP&wO4�p`x?}&�ξ4�S&���e}iħ*7�܀�8�7�6��QF߆���
�l���l��4j�B���q	�7EX�hO�!<x`z�-��f2��`�1����>�w���x	�&w:L(���G��̷��F]�_�믬��f	jx�3CkÚ���c��j����hX��&,L|�>�)h7xe��U[i�N�8�s�_�����ĳ|��#�������4&,$4.����g��C\� �
��Uo�?߮(�a��8� 	,!L\D���i e�4��6�g��B",s�w�i�Gj�%�N��W�9 �Պ��d�E���P�(����F�����՗���<>?�\ņ�{�Gj���0�/>%�I������=:{�Չ�^�;�:i�*//Jl�P���Y��d�a�h���[�pVՖf�������C�.��J�7iY�S@��_��+�P(�lOl�����s��K83�A��X��>f��J�R-����=6Et}���<�\d$9)��D�&�K,�&%1u��~5�4њi�-��O�i#Y�S·v��d�1�g4Tъ�v"᳢�\x�np5��y�Þ��o\q-ò��Wp+�Ns��8��Yn$tb�ܞ�c�&�`�/&�"��n7Ys^/�哕F�^Zks�UL��J�dZ��Eo-���W%��s� ڸL�����5Uy9f������ɞDr���I���	1���Z�.=agB�0%���z�V(CB�ٙ"Y�H�I����}[����X�)�I�<�?׉n��,�,���l�k�4^����}ɤԣ���ƍW�NDm��Rlڰ�1=ρZ�nj]���R;@��!p�=2����2�OZWmrG������^�|6���5�(I�E�\��o'��'͋��	��oRs26=�ٰƔ��
q�V��ܐ�F�sc�i�%��r$PΝaH�)bϳ��#�O�KD��H6�՞��+��B�+=�������f�:�Jt(Y_��XZ�]Q�!�t�~�͵X#����'j��*�%��o7ۜ������#C�٤Ҹ7��9<G�w��E��J����g��]���$T��pت��T[��<ܠ|�kj#�q���Q��u��8:|�A�C��-�*=�넦��&;�z�r(gwj2���]���8�G�r]n��C���������'�D�����A��V�L`{��m��K�>P�̂=����d��@S���OY��d	�x'�j�)��ߺ�ƔF�%�W#�$�d��/�z�+��.	Wd�>?�iJL��6G����z8�$,6ɞ�-���ܐ����!���}ØE6�6�Q��+��j���0��n�ס�V�����@bh�oklS�P����>a�`�`}�3?G��}�6�2�s�jU4
�M����?{4��K��v�Ն1]X1��7a�5�޵��c8�"t��[�ͽ�1	Ri;��zюꅷO�x��Hg2��Fa9�QԦ�3��7EX�������s�2�ky����)D�Z=e"L�V�?�%ӊK'�*��h7�k�V���aJ�'�3���x���?�|p���>1�.�k�ö�=�����9�����|����0`�J�kӤ��E��p��}��Y>��>�_m�c����zn��-5�GT�ŔΟ�S��7{��Is��:No����cR����0w���"4��N�e�A�3I�U�qt���⇀��;�Ic��
ٸ�	��&���V�a�Y��L�+�vx���8�?X���E��so�Rc��}-63����h�2�u����l���vO���xu�D4]��_l )��2���#�ǧn-	'�?Ҹ��%�r"��+��Y[��4�V����L�;\\I�Ek�/w��X����vCM�[����Y���R2���i�;�K�R��4��&�ۉ�� Wٚj���P\ؒ�aJ�I���j��,�o퍆!�Q{偍���5��ԭC��m��fL[O����D2/�_�sLd�]�f�d��će��cۆ�ٳKx��>Ss8G.���6	��Y��j���T�ۛ�?�b�"����ʉ2\<B`�B�ŭ}+�~^��z��G��:4�K󻶅t�w'8�@~у�J-]^.֌3�����5>/�4�udϽR�H9�I�vw��R�d���G*�
	�h���@z�6"#�`NA�,9���a��ب_8���1������.ʴ�?���c���w�����r�bH�͍?;>��3�X�Bkh�%EI$g��
���|��>4q�O�Ĩ�'�-(�c�^e�'}'�7�{��P�ڬ�m��~�:�K�����B%*��/�]t�k�>)�:7�j�� ��[3���h��ᢗ={q�䡚�`|�����¼�m�8�z� ~�I�a�n�-�a�KY2n��{i�\H�G02�*+�0�KÉ�=}��;s�	�}�̀d�6�u��vW��s{b'C�?$�`�����-�^��?U�����e�}�wr5����=c�E��X*]K��^V��	�Y�:-��&�:-B���0�J�yCB�m�L� �]�Aޗde�����%ǒ��ߚ9	'u����JnE�.��c�\�Y��1�#��t�A�zڦ��Sn�|pT"��1J"�R��_~M��9C�<��t:V'iY�ʬu"�?�_��\X�&�R��zm6��<4&��O����P$��j968�z�L�;�'UR����oO�أ]*Qג���~PT��d��X*4M��<<�L��>�+X�O���5)��mJR�K<W�7��{��v*�@g��+!_���p�VV�>_��\G��r:���$0�.!��ʢ$��I=��JQ�mfg�G,P��!�>��(�C�I
я�̭t����:�Df-8ˌ�8Cq��&	\��L0͙h �p�@�ԟ1OO�}-͹9�}�p�c�䕽GG��D��9���ËԢ��rb}�"�&O;���1��]k�>�Xd�l*o�!� ȋ�Έd���P;8D�4�jϿi>;$�!j���xմ�a�\�u�."lօu�֮[�L'��^9�꣇(�èdߨ��Rۍks��,�[T*>=�w�4�+���b8K����v:VC�?y���3.�7���'�WL$Њ�`�2���c���1����g><�Ա.�*]f`S��U�A%��_P����<�p�׵\�a.���~��ߣ���؏,,��}z�Y8=R�+�ӄ����6�*��6��f�~�u���Q��Ami0Lt�rG��rU�ɩ����V��8�K$��i��Z� }H���s������t/�k���#U�����H�EZW�/p���00��Ə�i�ᑺxW*-�<�j��d(0�Yu!�Z�5z�M��TKm��T).Di����4���҈�5���KE��'v���c����oYN0��YRh/,}8�*���v�굧Ę3RS}{&���x$q�9
&y�Ĵ�x	
5�P�Sl0%��p��[��Ð���0���^�y.xܜge�}o��>`�ḧ���������|�*��pS�/(��Q�P��M�ki���z�ckG���kr߄�"��v��z���;+_��kl�wY  J	�ZԠ������;@kZSM�$��ةK뼛�Ђ�ɨۖ0B$�NS���=�����XrQSL�A��}~6��=���<�j�;��N��C�X{������b��n�PIlR�\M�Y�NgƝ�6���#���r<ڶ��>f,ϛ�#
}�9p-���(��ņ�zv6���y��l�l��>6Q��zM�p��7z��ڴqGd
�y`�2��<€�\��ax��x�!;qa{!�]U]Q]�Q|`g+��1O�������D�=g������ M��]T"���&��<���q�P`d���hq��Z�;td���MǴ��W�lQ���g�NI�Fx�}���S���9�	<߹ψ�s8��ߢ<�������;��R�Yf)E�>�J������lU$(��"z������0 �dzg��X��(%��+)Ҙ��dM�fWĘ{�_2����Ō��v�m�v���j��>wk��ɂkA�;*���'1�5��@G��k�SI���c��A�o1�9���6#��9�B��:z��Hx��׏1@&��26LiIC�$O���"�� 1ZQ��Cp�����3M-���O�9�_��*d͔ͬ\�W{e!�!/�c���LI�����%���C���rzOcN�<�1���>ƀ�dW���4M�dO,�[�����\�<đE�_��y$�d@]d`ʞY)U��C�z�Z���Y��\�Viar��!��9����z��I��0Be�XG�+�\&\� 9E׉����u`ua�Sץ��1������Y�^����%��߻�',��L]��-OaHƧ�+'\��	cI9, �D]�8�{c��b���	��Ѵ���PY�|TJ������S��VMG�=Z��b�-���h��>5�Ƞ��!��9��	o�c�8�g�����&v�H1v/T:
��ٞ2Ѳ�Z���v+Tq���P*�*�˓F�l�M�a@��a0�n�N�}Ub�m�M�ǽf�xb���<�"�k�ǡcL�q̍�] �d���5À",Cś[�X�����4�T�YCF���r��-O���m�m�s������Z�,b*=������ʐ�f�^�xޥT� �j>{t�Ӷ�B�W���IZ8s)��)ф�tٮY4��k��Z}�&��i�l?��uz��Ǥ�!"�<il��SW���d������F~���'1iH/5��n�Z5��z��8a��2I�Ĥ�aD�׍�I=ۡ�����^�o%���6���t"�|�U���T!"��At�ͮ�u�8�^�>e%�e"ϭ�t� n3,�����"�;��h-��	�SS��Dɾ�P���x��Č��=t�W�1���?�����J@OY��ɓD��5}9�Y�g�92أs�k�b�Xe><2H��lD�}M-,a�7�b�R����'�
 �5#��PiZ�~�<�3u�����=Z7��
�-1
&�g��Uc����&X���1�*T����S
U�2l��n���^��mH��)�>���"#� �x\YV���OqXN6B����L��}^��c�p�.�����h!ɸ�jZ�Y1l�^Vn<�w�غࢤr�RrZ�+p��E����׶
���P�ŷd"�X��ڪ��̅bG���Ӑ°G�c�$1nBx�������n	9dc�F��~�����?�=C��8��X�!����u�Jb�@��oܺ�֢,��8���c�H�{�G��f�6JM��vZ�yڱ���]����(�P���f����W/㦂�DI��I�"dΎ���"��E�M{0���o���5����b�b�vʕ>O+�[�] ld��M�P�x�K(%�օ�c�g�&s��(���u6q����`��#��w�WQm[�T����eJ\���՘�cV�g��Y�o�T��'�Z�ܐ쀷}�g��{�{��a��<�B�*>R
1eg�����!���5 �8e*��B��vR��:���"����$Wi9N�y>H"�x_5���=�}EU��.�	jm.-�fѼ?H����UM��_�/��KۛhIn$I�f ���L&�LU�]=�o���d�fgg����x�yD��-TUDU�Ar��:_0"#�p�z��H� c�-�Y,^�-P'ఙ<�9n���
�C��!��F0���F�2gY�;���
őI�'�^���ŠtL�8�;�1fC�0/d�-<'x���%�g�ὲ�����0���3AVÓ. [Ԋ5'��#��'��qf&���,+�X�u{�%9/)V�6�;�����`{��J���7,taJN�s���9�F�b�K��XyD`j[��~�V��ƲN�%�W,+=�~,檎����*��ǇE(�� ��$���Eƺr3�;�x�l�p�v##����c�z6M݆��HU�۷�csZ�M�	��h�\�?<��9���h�~��{��s�J���-��� #A��~���EAC��l���h	��2�s�..0��/A���JLWc����|taʲaos̰z`����PL(6C�r�VU�áB���'�5� ����.s)!H�HQh`�iX0BA*p�Px��� ��o�����gx���$s���P���]�;;��O>��F0Ut�������X�V�$��h��jޝ{A��`���\�HJkݿ[�L�k'݀���e5��e3�%�"e�ʜ{�T?{�[�����Ơ��5���&z��4���� M%w2{j�6k�K�
#`�H\ͤ�['���	�j���#?���wa���"H�$�kI�`ֵ3�����V��;}�����7>����=Hh��z$dD�a+��β� ��<���{���Ԣ�|�}v�ms�VɫW����:OG�� �,w�N�˒�Ŵʴ��z���J�������_����FC������=�w�X�������2Z[Dh��#w�$ԇ�Bo�#�'�9,OW�k�N�Z��B��������[�����%!!�w�>z�_>;B'$��FV�ћ���ͪ��Y$Ĉp��b�G���)>˵'�}�F:-��JH�<Ú��D�u��yB���/�
x������3@ѺS<Ql�=�����r_2�T�FQHO�X��)��8S�&B������	�l�f;�ҙ�M&G,�� 38C�����VI���K͸�����U�?���O�U��L��z ��֨���4�,�,@��c���.��Z�����r4F�2Ff��KN�ΏYЖM~�n(/�%~�����F�q��"��Υ�q�k�U\/<n���{���ƌ��N���rdǒ�ws#�.��i�'d[Wv�G` N�1n��ͅ}�_���U���ug���Q)�I�uBbg�{k���ap����A�Q��{��`�!\(���z�����a�L�@2�& L�,�^��ك�y�0���ғk_�Z��o��@5�>Y��iã�u3��`b}2���!�k&�!�ҲX�Iaq�`��8�dT�߰9j�>d>ڂs�Pĥ!|e^�2GͿvG������G(о�A��aߊ8�o6�r�L2�)}B������-{_�8T*�b(����%��U!y��k�s��r������K�|��>d�:{�ó�;$Z2�_}��
G	�u�q����[L�L����n��a$����,��j�I�����m��b��p��l��
{�Jz%[G��+b�&���ȧ5� ������wB�?�����v����*����MkBF�v$n<�u'���h��{=��Q ����][��h�&h�5��Tm���M�_eװ����2O����R��o֗������HY���-GKDЛ+�ݬ���M"&I-��o犕	5q�"a��H��=v�,x�*=F����}��o#�`T��Y�Mt�#�g�I%9����^R,��3���ֿ֢:�{�2���<T�jJ^<6)����|�����VJU{^�*�Ɖ�:y�p�G�l ����`b��ڸF�� B�ģ���<���`�rl��4�TCG�A�����L��Y����_��omS�˿ڗ�-�;m���{26���;]��DK�S����
Ɵ~�IaK���ɻ!�tg��[�7߁2�Ww�\����˟��'=t"�=p?~4�$XP�7F`�\��FID�̢�?�`���{��PJz>�}L�,��q'I����T,P��m^\�i�R�;�B	g��=�A7�T���#�R��1hJC0�:MH�D\Pvu�J�p��DC������d#ʆ�t������sI"L{1I�-�"�N�eiĜПK?�� G'a�A��%�hF.#.��g��ޒRl�3�|դ�,�s��;�
���(��]wy�������^�'�<����e�=!��n}������0��(˴rYvL��4�����h��dY�h7�ϞA��k5 ��T2lA�<���t�9��@�X"�}�R��K4�<"6:��ϓ��^�J�a���z6�M��4OΔ����}���^z|0�ިxi���&c���X��ͣE���A�Ma*F��A���?�Q���o��\�A!Qf���G��z�>�`�WK�mS&�l�M��f�nZZ	��9���zXXz�0f具�֬�����`1���7�}����}#��\��,5}�Aҫh������0��\c�C���#ɫ�z�s��}@��Sr�f6�0�LN\�;+�T���,�rO9�����&/#��xm�	26\��Br��tĳ�=��*���^���̫O�w�UA4G������g�B=؋�{��;iZ+�{MY���T�H҉0
P�p�;kX�����Q�?��N�&V�0�5�UE_T!Þv;4 �v#�����{���׹�W���{Of0)ֽ�-Kj�\3�?�O->Z
ɷ-�`�y��YA�|97�1� [�x6�z��}�	b����L��A����ȧ�$W�џ~�E�����[9�!
c[Xzk���հAo]A'��Īo@|����Ĭ�g�&�н��#�l����m��~�
���:B�b�ko��h1*d��q�&>hC�TV6�h�����Ou�K6�%0n=�C���va�Z��.�n�a�-x.����wj���^�a@}�$�8	�+>����H�P����9x�^G�"�T3�u��+M��b�R��dB��W�l֧Ÿb�G�	T��`�rH��8�F���O6Y\�쭐-����R9 ��x�$�b)E�������xWX�c^j��~U|��Q졋!�yh_��B��B`��X��L��zz�L;�����?֊�8A>���D
�RBI����;�c_���*qL�2~��qo��!K�:i����C1e�o�p!��ք��(]���B�h�̵�a�H�AE�W���y���G�;m--�Co��M���'5��SΌA��Z�b���,�#p>�.O8��&�5����y��b��č  =����4X�D�+G��G7��?]{X�� �{�������VɑJ�լ���+��ēy�X��Ԣ����1O�G�4Zyƅ���������}<��0"�	F�]����:ks�V�Κ�����/�Ю]=A� B� dURBZu�{��$D"ݑ�3�,�l�(Y\�sl���hTp���mJ�����i����ŉ�p���������ʶ����,����$H�ZEVE3�@�;ͯ36�Xu^�<F�56i��+�(��8y��9ؽ�w�Dr�7��m&hX���U)9[<����/q�3̆�֖�y�Z�'���5� Ʉ�Q� �H*6�L eKY&�r?�A?�axI)��<{
�ц�#��%+�����$L�wc�j2d�<,#�<3�� *�s�-҈�.>v��Bc\Yh3���dq�������'����軛u�ǩ�.&T	��^/�/���f�>K�sQ����k�/bŶ_o�p[���C���\s-��.��� eN �S����7a��Y�����f�}	GځK] &A:�t���lG�����1���2|��b��'R���~��>�J#���#F%���%����b���_~�I���\��Ɲ�I���(JDE��_����ʵ�|��33ky�]��Pq��g��!�EW�Jل�`$�T����Ųn��c|�j[��JP�:������϶����;�� �Q��p����CD+9ן��؆��ƚ5.E��z��2���7H.E��XEUѼ쵶C�3Y��=|| ����4�=�L�ޢ���F����\��2r�l��$��d�K \^*xau�Ⱦ+��*jd���Y�f��)R'���<��E�X�gO.��U6�"�	[q,�(�Fu�u�_-�����@Q�k�zP�#�c0�ת�ޡ��G�i�Y���N�{ؙUJ�m����5����q�a�5+\����5?u��y�_�{V��uO?�9�	e/��u��V��yX��{cθ��k�s�m�t+0����^S�4eڡIݔ����*D��f؅u2�3�{����O�i��*��T6���"�Q�Niٱn��TLQ:
�l6�h�����s���a`��V?<Z�MBs���D�YZY�h�*��^jP��z Ѳq+�7�r����d=jp���v2����dC}��ԧ&Z���r��NYZV��Fgj� ��ϫ���̀m˒V�h+�����$Ðl}r�������D,�x�\Y7m�}CaC8EH@�ȋ�~� ~�Љ�� ��ג�	#0����,�*jJ{^ѹMH���BZ8�.9���#F��n����������[aa(c^ܘ���!�n��'�N~�[�P�g�v?�e��(*��u�}Tc� %��� �c탊�+���R��D��9�W�@8�2e�O=�dY%��Ic!-���Xn�Sĳ�C=Px��d{��V��kr�4�	��H1QE��J=	�Ń�:u����6���ѳk,��t��^���KT��`ت��|τN�dd#�� .�|���V�L��(�(`q�<��3ar����V2g�$&~�j#�_���"O����8�|����h�G����ߠb
�A2>&��g��g!���b^;�v�do$@�P����9�a}��Y�Bd�p���UŨ0�b7Uh�{���%�L��n(��zh��N���y5��L��Y�ރ��t��g�,��dGʓZ;����:���0�F6�d�!zDwzUTd��3��}V�H��uJ��hYt�b���ո?��O�;�u�rR�EH������9~vog��U^Z�Ғ|���e�/���1]&���i�_��%/�ڔd܇��f��<>N6�#��2����a�G n�D�s�uB��>���G���q�ބ�I[�?3,�������C-��>�3Y��io2ϰk+�B5��Jrj3v��R-'/���E��dC������oz����/	H�o̥�fr�-�j$���v"�R&+fꃈ$��-h�j���b��
s�BaV����������w��6�']\Zf*��� �\�)a��~��Z�O�X\;R��p�X��-��D���?�Y�+�"�=x���(_���	;
RyI�K��[L������������Obo��j��!+����*��1�L3V��rv�5���ʄ��B�_Ą2��*�Z���T� �-BT�	�8�%���4Y/'=;pi����B�#I���c��ڊ:c�Ζ�4�EQ:��w�*!�Eq�B&���H+_n��Ð����y�D�[���{��2�B<���`�=�.�O�GZ
	D~6����,�:@ߙώ�t�.h ��9;��)d����)�BTz�W�&\����]��y��	�R'�k������;8J�g���]VM,Y��	�͹J�@���9�{�����}�|~��K�{'@��Dh�UKMZ�~DUC���V��������z��[�ݠF�w�����U9Y���G�H׸B�4�XI��tm>�@�bq���BDsߑ��1z,�ӕ<{E��p�G��ev&5�7P�����I
T&q���"T�V�%�,,8��ꮣ��������+�Й}���mtv����[��ǜ%ƚy\u��p:���	,O��Q�����U5q���Y�Bܨ�Ž+V�ӳ�ʏ.�8�ږ��*��� �A4>�`κGX�̛7/T��P��[y�X��R�L�TP��s�	K��KaR��	Y3g��`_.��Zb�D���Z�S��ꨒR��������1�8�I�m~�3�j��=�V�9y¨�.����8N�+������@�hr6v+S�K�Z9�t��SŅ�|�4@��l�{l�W>Rr��P�~���&[f�o���j�=�~�L�d�Q��/V�=������v��r�e��0 �&3+k,������%��F�6M-�Z ��0�ota�W�|m����" �ĢءJ렚ٛ���t˾�A���&��y��*�`/=�ֱܯ���Ջ���׊H�l<�\/�YL00�d�ф�+�lo�oQ�
�u<��d�@Zf�-j�F]5����#�������h�v���
-�+;�Cc;#29h�[�n��݌�5#И�b��r����,0qr�������#�uPP(���a���F��y�0g@<�P�FT�=�b��� �k�$bł4�����TXQF�1#��� _,�-�]��I���E���V��N�:�T[9Xυ�J{�c�6ﲍK��Vj�7S�D_����49/�)g��Z{6k�B|�`���zP�=�1w�p��Ͳx[���So��s�53�ß��̣R75C�:(��! �⺪�t&�z����r�<Y�!?��YJ�P�$"�ƀTY
w�����䬭l0y�|��ni��je~��7�!&��\���a�,�ʺ�*H_i�_>O�z� �,�-��%�G�9yTK�Y}R��䕺'J�/�O?���̬(�^ܘаB��������Zg�)KE��l x)Z��Zo	-H)�@�~\	�M��F����ϕ<F�/yN��",��`�Q�m��I�=�f�%���ă쓧u��Tx����0��{��V�K���
�'��ܡ�� ����\��l����E�p�b��2��k��=���*Z�N�T����a$_A$��}�oad����=,'���!%�� d�҄��"��1���3�� 2�p*�Koeί���4�[��b�&VPr�����u�0��`E���C��ߏZ�vꬿ�������SBBܫR�lT�V�,�V�ٹL��
(�wN�#��,֐����B^�D_���4��p4V�q,S>�!L�{YҋT;@�(d@��
ȝW qR�]�;3����>�e%3-'	�=�����O�@���'�x�,���Y��I�j��߿�b����OWJ�Arz����j�K���nIW��Y�֞��H����9e(g�˗�l�WNֲ�>(���~T+�ɓ=�8ِ���Ma�)1�j��'���YX�E���jUӢ������i�����E��۷�0}����fX-�G�"=ƪ��ԪF
�M�.�5CZ�+�iu��;�Z�"HE�$�!�@%��Qh� }\��*�,YW��}"��X�tDa� � +M�Cg�I�Ғ|7F���+l��	V����
G��<��'�b�,���	�b�7�<ҫ2��}1����xNƮ�� 觰�̼�?zW�մ�;K���!�yr�;�a�P��bg�l���L`} ��Z��g/	�5*1n���,�]b�������$� Hz�G�ĬSnb��gX����Bm���Ls2�^���</����Z^Y�f�t@@{[������vU�Cb��.Td?#(L��j��yLP]�eh�8i��Z(�{Pk���}��$]o�K���7� {��8�O#CpL�Y"��"�#��m��Q��8�I+�}��tj�p�O������Ζ�V�p8���'�*Y��� ����4kN��=���%�U�rL��F��9|ڷ�%�c	����``���_�E��ב���3[�<��m-F�Ԡ��a��i<�Eݫ������v�	$�Da@j��#� Q0�	h� 3����/�0�Ue����P���y�����5�^'���Ei�RN�����T?�3찎��Aޤ̫x�浡>�L����hY|�`�,��	,�e�;K޶��q|S���V'�0���d����'���YĲ�Tϯ{�!{��wu�aE�r#Hj�J�AY�xv�ʼ�ⶵ�Dn2x� ų��R5�����v>��I��C���T�*d^�p'$0Sfo#ǳ��cL�*s�IY�'�5`aU�>6"/mK�5k�K�gf�\p�O`���2Q�q�y��Y��|B\m�Z��R�/�b�3�7fuSU�[���2�2nc7yFLʨ���?�5E��(����i�
�VWQ�b�C���^�ҽ[4�cƕ��.�:G��R �[�B�M�Ig#�xB����=����Ě����O��8Ҋ;v��B*��u=�TY�ü��<��K��#s%����=<�X}B5#���@h�X������ƦwTD{��4��̯̏(�Br���}����i�H/&�� #�Z�׍		��e�o?[���?���?�����{��aU�& wч��:;�g(��mL�і�=ښ����Y��#���Iy�hunULmI`��� ,�:��b�
D"m����u�v�<�=��F�\�
�����޹��/>��(���YX�p	�c�1|)��m�M[2�m��sYae��Hr�����w�)��&H��d*�I6����w��.��{R!	�������r �-��7��_-hV�ui�-a�
IDb�.�nr ����2��8�7�{��в��wr��A>[�3�~���K����JY,�LK2��g'�s1����h�n`�J|�]�41j��$)/�*QXr`�M=���*�����zP���,y���@nTÈZ�+�Ti���Y�����*Y�>8�R�$$�˅>�8�~���Y.w�{S�6O:�fn֤�Lw��%`S���,�����5L�����>��?�L����ɞ��`�4��T+��	�C�%������k�����_�����r��.������V!+�+灠R�A%H��l�qk2�ZMBjP2�xn��kѳ]9|Eɼ~���L���:�d8č��MdV�	�u��~���F���,��!�$>%�5Y{Ih���ū�k���s�������-�����E/}��QRN"v1Dd��^?G�Os|��ެU���O	�1xٌ�ς�7�Fzݵ6W�*H7@��Ҋ�+E�7��e���Ԁm<8#Q�[�	-Ж���ߔ:�T�8 �vk<�2�ĉQKE����'h
FuG�8���~���\R��Z)���:�@j������-���@�>, ���u��p�(�3���H�4�����B��~>c��Gk�_��J޲d��K
 ̥	���3�l�!2�����Tb�POS���;Kܦf�W�Z�J��R]�f�ǌw�K1������Dc8�rn�sT&�ׂ:�����'��L�O_��R�:@�@[�ir{X^śj��sb�O;*_�~��$��&�Z�l����4C<��'������\�6��6�v.Ժ;F��%��)��`�C4��U�]��uO���/�?T�QJh��.��0�]0?-��Hq���f/n�������� �	�/~�Dd����5Tv�C�Q	U�+	uXTB!�c��]�*�$}�T�<���m� t��f�	�2 M�,v�,�ͬ�Z`�^	⎃7�B�$�_�l,Y kdqX����)�sAO��l�=��O`��R_�$2CD;-���Gj�e#Y<l�k%�|V�ǳe����+���	�m�������B#T�ЂXH�Y�G�:����T3di�v��N��\�ܯp�� �=����~��!!J\Q����	K^��������	������'�s��|��0�*��߁��	i�十��%�� �HƪɅ�fzJ�i��?x�19������ot>>��F���^���	�,*5|%Ș��tv<�6j\����V�8cYzP/@�6��0�����'3\����YY�X�j=�s��A�70�{��L�f��gI�Y��6��e,D�����Q�B��:%z/��x��hB��9�b��#�<�Y4�b�k�(!��|��z��.Y��>�:6��"��qc��%-$b2.�L+Ӻ"�9ۂ2&$�'tm���?���,�n�k���y�E"e���AFh���ZcM"<?)�K���Q;�/����`��̢�H�;�0+%k8$�����h�T��[two��n"����O}�w��S U"|<����/�.��U�BT��|SǷ4_
*E7��h�_�i����1�f-'���<���b�/c��a�Y�V[� ^�ĉo?H��$xW�&\Ɋ��%���Vw�|�4o��V�gз�k���6�%�Oel�dԟ~jk����_vȎpI-̰��.��`@*0�`)����nҘ���#PR�*��3�ǲ��5	N���ʆ� ���d�B�UΌ�Gl��]q�*�o��O��s+r�Xt�g�E��B�,�d�d��:�]<�PJW��'~Y��R
�{�3�;W���A&�<����Q7.���2�����i�El��ؼT�tD��ܦr)�1d���pݙPe>��£���Vv�^f�ס�����	�at8�U	X��y�k�rK�ļ��-������TC���w��bN��8��h�=bb" Ξ�4��)#;&&�����CJ���_�V޼7*5��5�� ����t�g8��^�
�Q�<�1�fQr�:$�Xt#[PT�p��<�G0؛er���-TH�0��n*�����n{?htS4�PͲ�q��?�O^�Ę%�I���V2N�3#oE	��Q�(�Gt��"�0�{����!]3K��"��y6�x�������~��s�b��z���X�ۃ2~U��3Q���c���؅Ejkw�J&�/"�IS";��Q�`�[���U@�:�+lƨ��ep�ek�9�f����jz�ʂB���l���H��ݒ���Mv���+i���]V�T�d��W.Ku�;�k�0�"5A����i��,�_�%�x
�8a� #��s�~Ql+��
���0����"9�"��I�y�t����a�{�D�ڣ!�ջ��u��K�J�En9����K�2����!�晾R��g�ɉ�#As2ws���G ���Ѧ�V?J1��oTK� h����Ы��H,�w��s�AeJP��5tPGY�J�Ȩ����rZ�Pn��-Qc*���n@%�>]�X6�^�&��HΜ��B5�O�q/և� ��~��X��{���%%�;����(� ga�%xX3��?��0��G(���Ǆ���n��دG���f�XU�q��9�*�h�F&-��Y��c�]����̏�d��X��FR�	q�\٦�؋D�|2��u%/��q�&�)��&�d��I>�X�ռ�[/B�	#+ ֻM�.u8��*s�Ks\%ٛ̽�s���ѽ�x(*�����b�}s�nq����a��rGh%�	��HV_,�^^s�3�W�Ԁ��f�𴴕�]1,j�4:π�=���H����A1��@����wr�&���z��>h�ݽ!T��hH´$�1�sri�V��Jez@B���<P����o���3覑��/���b�2��n
�^��xĦ�/f]_ί��Մ��#�XX8L?��o����ަ%.�nX82&[}sZpY����(0"�Ț��)h����V�q�֬|��C ��D,K:�T�o��]f�XQ��)^Ԫ�ȶ.Q�Y2���Q�-���us[���:/��{���R�) �6��[ēiQU���./��ƣ�qߢwc��}qq��N	�_ {^fk;R�
�;��	���ppK��<��t�>�2���݋�η��d�I�v�U���Q!����x����$��L��=c��X�u���*a��O��MY�PuD�zf�Y����݁�������Tt�QK��n��pH�(�_�zR�c�Ϸ�(o5д��\/g썶=�ƒrv�rxBo-�[����N�<��~Y��5))�����'�=0��ރB�����I�D�0�~/ D������e��N�+x�dmIkB4�F�s�k�~�g���{���6���5�@5	-P��h�e��E�7�̜��X*ndҵtV�u�|W~Y��L����J[�9��[ڌ�{�0Fς�ӎ�(,L@A���Eq�倸c;z�`KR��u�m���&5�ӣ�)���o}C�yH�X�B|��a�,!.�x�՛����^�������>��G�Ӓ���?�����J�L�Z�J�;lljd9x�b���7t���Tw\�3O�@E�[;�OWwZ�i�� BF�(�%��Z(h�lɪ�;�j,h���3/�R0���&L&+�e����#�_�.H�2\�/��$l�쫯��À=o�����A���{u)պ/�5|�u4;J�S�Y�L��9c��="/�e-��ZC�{�ҠK��#`�чޚ�ɗ�#nQ�eBX�*V��s���,ހ��Q��p�F����w�6e��`1��#>�24"�^0L�<��ܵ�>DX�����N{�YL$�w@�<�6R��()�.����}$�l�d���ߕ,�,i�3�H�O�"���^�Ze�n��T��tBك��� �HA�l�b]����$A&@��I� ��KҊ��F�p��ks;��Ć���A7!S|s��*�H�`n$N"p�Z=p�p �E�m"F�D6�d#��>M0ka�
!X$҃PL���Q���V�s�
���T<�B����B������u��
����ߛ�#�M�x"`b�[�l��|-��Z��Nk�͵�����0K�m����/é�B�x���7f�����S(��6�Ξ��݁��%�{��;�{��>���J��R%Hx�\��B$x�9{6�S��������~V5�,8ם�*�;C�6����Ř��"Q:{�	�/-h⻙@��~ډA[�<X>�@x�۝{g�V�����}G�6��k��9�;m����v���3�P�s&Z�a�h�nR�����e���U�P��=DxĔId֥��g�|�;7?ڮ��!2�-
�J�&�9�ɠ 5�^�*d#p!�Y�uT�2->A/�MPA�Y����
�D��b����~7k=�Z��߾��K��%q�.�N���ɿ�WȑXdgQ0Э1��Z�w��Z jѭ�P���=?w�ś�'��VC<X��U/��%�#����|x���r��
5٬2/��ن�H��a� 2�Jx��� B�gi8&ց�1�*��bm��X-�#*�e%Ze��pԄ��,/%
�FxaB���gp���`�:����,�/
��Y;��!
�n����KWe���uʹX`�s�11�J�	g��hئ^�7���Jf0��֬�q� ��1���o4d4N�̤��R���Y(�Z᪒�%��ueB�!�?W��D�S���>R� ����X�e���+k��!�@o�֘�J�E����[\Y�42�3�ع w2ժ*a;E�!/
��d��PK$��uc��V��g��]��zx͠�[�\��8s6�GFB�hWK��2� �!Ft*V��4*.+/C�-YM8��C&��b��:��|VX^��f�t�m#���c�a�~_�q%�75CvP+��<�`"�Q6��* >>x�D&S�c$��z���5�b�ˢ)�=��XC<�[v��
&!uw�I���8ʃk�YI��3�.����+�H�M1)��/�(���Y4��ޟd�ZW���؈��m�ЋIY,LPB�Ï?�@�a���ʦ�X1yB^���X�ujfS:;(J���Ϻ1Ņ��RF��:B&yn�	U��x$�r�$q�?@I�|� d&�ӳ�^�5}�̲|'�XP֗)\q��Fd�e�h��:+~M�ݼI�X�;!��&yi��f�JI���?"�y��8۳F�����v�� ��H GA�%����gX�zn�������L�3���Q��Έ�����ep���Ef��`)c~B�U����(��i.HY�nݰ���\
s�����[����W3�c��&o'KYI�Y�&�ѱԕIS7h�f���D����#b�̑h���qP?�KI�T�!9^ٞ�rk�'��(]5Y�4g�]������j��k �5�tY�L����ĳ�`ƀm����RR'=eԊ��������W_~��̤��������/��(]��j������L�Ӄ�׿�M�.�=�tvS������$��V�b���1��b>\���,�2��ɘ����
������Y"tۊ��h3d��[�ʸnJ@�u�S������ʿ��O�?��/�T!q>A��S(� �Y�պ,�����^2G{�CZ|�	�`�;-��Ib��W�N񒂘�$k�����-R�'�T��B2�q��{k8�X�倾�KRaK`�r�y^]�]�nqxi5�ݯ�v�V�|�"�����g����|�ͭ	Pُ����ٱm�ģe\Qef �\�wo�`���F�#k:!�&n�4���x\��L�����c�n��Yc��Q=��l��r��۷V�W���Y���'?�T�'X��l�H~ =���P�|T�閛�rB��5<d�ŋOTl< ��1��˺���k ϳP���V��s/2_�'SjR��ȭR}D�7�u���:T�SJ�%����$H��-ʈ���y��2KC�eA��L�Q=Cn�l�$XŐŕFџ�M�͝������Z{�ŗ_@�[�P2��5�:��b� wИ�!O �%��1H���/�P��.`�HR�y�]�ip��6zɬ���n�7Գ�V6!���*Dr�A[�5�;�99�Y#��X�>�^��>�����:/_�%B��=(�2�L��/���)�D��:ˬ���(�kl98_fbb�-ɀ��M��T��|B[B,V;�ʜHi�h�<f��8��v��i�Ͼ�[�@��2a��C�ϻV~�|���$���A��/�|�o� T���;g&;�;:��Ԭ�s��Y'W���d��6a���M���`��{�:Y�܃0<9�3�?����=��?Q<�|�}E�턎�X��H��lu������p͊Qp�_`0��k�[mgJN��ϫ�)��P,�=VG4�����{nb�<��<�X�����v83��G��#k5��������ɧ^��D:ˣ/�q�P$����d;b��,h�¸O�������fF�ENH9Ϭ�%�:.+P���)��j9�#n��4ެB���Q7����]`)b7k�`:7f-k��BP�U���C�P�^7���i�#dn���CӮ�̍H ��W����X��v&I�.v��4�̹2� ��J��^5%%�o�ӯ������Z�(P'�7Y���MM�(�@VQc����O 濽A;�Ul�Eߧ�{�>��+,�q�)���f��&E����{�[�MJ���H3���+��z=����]�^������+3�k��M���5����bu	W.TB|���A��13�Vf<˂˿٘P1�ɝg,p������p�^��ɕ��%V����L�	����4P~���5B�=�j��PX��lց��+�ȹ���e��
�a�]f���XJ�|c�'{��r\�Pv�J�S�O�2�|�
e�K.J�����K��p�Vi�28���*H���"����K�s]J_ɇA���V�uN��x)6E#$�?���Ad ��]�X���q�e��ز���1��V��*n�T~�5���X]��U�I㹗�����k��u)�1�ԤҒ�N	�w�)~T;2Ni�F���{��_b7hLL��6{\S�y�9\��8���?��������V��<����7��'맘?D�o��)���������o:G����Z��NNj�hx��H�w;�CM{�rI{��3�+��h.�o5+y ?�HA�����@�cW��u�1>��T��l
㔌C���}��^���߮n��k���ȟ�^а�szx2rn�ɲ�b�ҢȢ֬R�I(B���^��XV-�F�^�ú�>i�I��|#b~�g�]cB��ʿU��X���²�`��݄ɽ��XF�o4_�~R�	0�UxJ�JHX�u~BՓ�{Բ�������i!{R�u����;;J��3BK
�q�Ӯg��@���,K��w֕W�{��u��h�x���d_
��
A�h.@8���|�'$��h᪌o��"�وW4�2Vv�e�����l|2⤔��aXs:m���	�H�&a�L�V�ŉR�����j�+>�F��>/�;ь�6w�%EZ�h|���A�`%k,qeVRƧ5��8e�������a�M��1����|$�5�}���F���`~XF+��)-ԮƤ�Zm[��٨���
���Z�e0��-���Y[r؍hמI	DX�� �9�UG̈u��gnƦYcp�@{����l��Ү��b��0/%�X,ƽ�5�"IC@��'*�Bv�@��u��H��mHƴ���|6-�X��2�X����-����Ck�΃���(��=��흹+�6�v�i�a�'�K�C���9�T�TN	|nM�3��H�w#��G������x�u�P,S���@'�cU��aT!)�f�OfE8�F�W(��s�=C�rR�����=E��90(Yk���>w�Y�hPˌca 2J���v��ن��Ͻ�	�hx�����i�`+�>���/>)�[�Wu��.������N�dec�Ĉ�! �
a)v�h5�(�=��S�Y��4���������Q��e|�);���/�d��D���]�B�gްYd�|�bR�8Fu%�;�� ��(0�/��F��M�q�G�G�M�����H�����"dw�=�=Íň�p���a< (oqM�-���.��j�g�S/�&����x*�=�ɗ�!@�� �!_�%��\-Huɠa�k�jX������B{��
�bG�\oΙ@ԇvŚ��̩�R��
�|��<G��x����&�Ș��ڼ�L~��k����; �5�	��;�����َΈRlbJ�b�A�4˜[`p.��p�+��S�����f�E����-�蕊�[-k���n��|�ֻ�b���rU�B���`���npV�M2�J�qL^�T�l�L&4�q���ͭ���kr��n
��-DC�!
&�),)�2�#�����O�9�V]\����&$S�L�X7R	"�d�z+H���s�V�~�ړ~o�]\�6��apl2g����O� ̪�����b7�X�V��Dٛ|)�e�E��*
��:�{Vc�`�v����:�z���&��]%��6eqx�'-�nn��G��������������cJ�.{c�gu��m�pб<M�W��M�����a͚r⊩ U0j\K�Ssw�ղ��?dϕ�\�Z�D`�ߧ�OP�nJ�3�%�*G4�[p�>��m� 6���R�p��AF�9���� -�����(��-d�'�Rn�krAK��.��m-���k�k�d�y;��b2w�3R�l�*q�iVAO�AA+��K<=	�#�h��"��;��E�F��Y���4
�_V򢰅���Ln�OaDb��^1�BMa�(2k?C�	�����h4��"P�����w;XG�@/��P��}�yfAJ+�?�Ӑ:6�r�b�K�7����� hAZݞ���\U�#�L��A3>+�$vz T�,3,�܊��lu`i(��}�Vc{F�yA���R�=�z��V*�B�z/�w}��F�4]�	��R��E�����_��#���Wak[��J\42�'lOM+w�~��J�I8��*�3����T��dr��2�K�at�dg5��0�����WR��z1��
Kĭ� �f\O��,��l��ϣ����?�l{8)Y�D��Β�dvz��@"G[A#���-^�3G�UM&�M�1�"���3i��؇u,����jB��T\�Y���u?5';'֓�������1�.�2֛��9I�e�
q��M� ��yr��B4Z.۹d�s�ZIǎ��� `\����F����3B;3�6GY�� �2Έ���8K�	60$��G��G����ix��IJ*-���$0a�ig��û8���2�u�[a��lxI
bR���x�j�ea"�Y�(����)���pH�>���� ������j�*�d�n�zD��Es<=X�e���0�97Mm\�����6!kD��3���T�
�|E
��:w���+��� �̩\�P��.!Lf�D�ԟc�zpi�����,lP��ն+;w�8h��i�]����`O��Il3z��%�4�+8�ꦡ��Yc�6�m.�j�*�uk��3ѨE�޲Ҽ���5��8�}�QgG�O�b� vw;�#A'�X��?/5N�A�ȏ�/��6����b����5.�+</�+��п�~�Z��h��]W�H)��+��Y!�<�d��2g�� �l-ޘݨ	,��K2Y�/�8%
<kOm���hk�*d9�)�#�RJF���p���z.�%5�R�L���f�F0�O>�T0!8���S#��V�e-�� �!�l�2��}��'�q�53�A{�Da����$��d����s��(�/`ot{��Xˑ��xU�,�Z�'�,��D�''���G�8�]���#�꤄�L {�Lo���v ���;+f&%�@L�2몙M�adeiʨh�!,�
x�w[\~��2�O@�"�ǧ�j#|6+��|���9e�A�\��b�wt��h&�D�#-V*�n������ŐH:�D�8[Hh4H��|v�e�kل*�[�ė�mA�)��Q��!*�ܵ���N��gzH����g��.=�ù�\�=*�&E������,Hgߗq����*������{2�c�/���;�؆A��N�2<�3����IA*<���G��E�,H8��p�I�X��	�l!������X�ZD�'~c򑷠5M�;�G�W�D�s��%�m%����{�Z� 5��/R��
ϟ4Q�Є�4�:?��['YkA
�%����͑Z��8�D(53�̒3I���(�f��jGs���BMۍ��� �b2Q�u����>x�|T.�p{��d�hѼ7�E+�<
����U�����gW6&����ǋ
�B ���պ��vv�f�I,�k�ĄEa�m7�#���-�����D���3���q��vc��AK�k]J(��Z��J:+�0א���Ikb������K�ٳ�(��/m9���uM�z��Ƀ�!_�gX��V��a̝3��?�!��et+D����=w|͡��1�Ӫ�j����H�>	Z/1#Db��iK��\h�D���r�LF�I�m��-��[+܀VΖ�����{<!F:$4�52<���݃�l�x�c�]k�&
���f;'p��S�)F,H��� Z��(]��ap@���!��-�Z��+��Al�@�7�%�6�`[��!��%�Yנ�g�b��*�:�o�`4<���Ye揙����$��4i���R��pB�b�
B�YZZ����	��jь�bt��B{#�C�������#�L>ǜ��Pc��Y/&�'$:HPc���x�!AN����u�Y��?�bY�%�W((hMRIx�
��05k8�l�@��߶\&/��T����.pS����"��P^���y��:��p8y'Z�k荒Q;z���{_�������Y2�Q!�[�5A�ѣ���.&l��ͳ�빓� k����M�z�i�l����`��~��5��b(�:�6!��F}�s#��#�?<��x�-qyэ�%ҚTeo�d�1ob�O��2b�����1}����/��/�/�������?�q�%����Ҝ�����`���"%��ڣ��8����Ԫ��C�ԯ.�6�jmM�x��]G`��v-�j�6�ט���#K*�0��\59�)��4f
E-��i�&�^�&@)�(���s����y�gGV���U��1�΋�-	��B�P7=CZ;Ʒ��!���e&���`a�h���n�������>R�{H�Z���n{�.XTqH͵���MFG�bm�;a�:ަ���d�	�.|��ܽV�����z"�##�l$|6�Ґ�ɞ$�sVg=d�b���U�%.�v1
�7��bVii��f�<����sT�Q�f�Ʌ���~����W�G)�%���oj`���u6�4�7�XlE1����|�����GŘ6�����5D�i������M���	3�T����+qϿ����e�-��ߴ$Q(Ȟ�M.6)O-�xV��'ب?`q8�f���n?��9"Nf���%7�-ښv�����R�u���-l�/܂�poL0�e�n���t ��_�\[��O�⬚t���"!B!���P�DC(�f%!�V����9�=y�Ň�2�[�OK��z����Z���(p�������R��7X�YM�hk��S�B!sֺx+&�x�}�R�?�� �h��&�U�3�Ë�x�Y��tA������g*��)S�����ka�4����`��Vl���[�q#@=��� υ�l��gB�-ƭ��E���B�*�k B����n���D��K�4��8G� l�Ҥ4��Έ�z{p��,�s(D�o�[��A�4���
�mH�����S��5���j�Jl����QZ	����������)}��	X^^d�і�s��W#�˪��pA3�	c����ƴp(0;׋^"p.�D�Iv��t����P6�M7a/�K7Y�C䥿�� �[]�^M�������h�%ǋ¤���/i�y�
C�����BEh7\����ܨ��5��h��ka腡fԏs��K*j&�5�c�\��'���ҽ�<>� L��a�H
S�JE,s�T4H3�Q#:�����'�d�<Ȱ��$iaR x|��1N*9�NJ(osvrl�0�I����;����߆?�kL2lB!��łZ8��>"��j4B��$	����]H�E�\���d�u8��/�a�DW�a8P��^U�HuN�E��e4�İB�G�D_��U^��/����"�C�Di��7��m����,ز ���������Qa�8^q�il��W���]�KƋ�TgP�g.ġ���+]�E�����E��G:+�Rh���F0o�뉣+
�� �x����������BL+.�����������j	��wZ��
o�����zR��K�"ׂC���w�[8�����Au_C\^���Y��H��p�	h��M����mU��}�"ͅ��9����� �6�S�2f���g>7�е�� �Qa	$�GuIC齿��_�65�����<o��3B]����<Z�˳�zM9���䜼��^,²n�&�S
'[��A�-��u��M�vmDW͡<����$M�WL���]{��v����55���"P�A���pp�āV�c(���b���@�q�ԝ���͵qLTS?'Q�����ʵ!]����ڞ�ϼ�<�|��5z���&r���{C:0�����t���a��°� ��j���L���*"�=���mT�Đk�����_/���}w{���e,�n��h���:b-��-:Go��\��xN���Fk�kT�FW�3y���e)1������Z6cʹ'�9��M�J53�\YNjw}f�*��5`�[W�p,~r���औ���VpvV��o~G�����k{��['u�#�3�"F����� A�?����,�(L����m�ľ��I��LK )�I�;]��e΃��_���o�����7���0����$z{*�M�D|�po�˻�j ��F�лu��~�������^�r�V�P�����Y������!�������G����E���h*�qAZ	=Bɥx�"u��Cd\6)���M���:�k�C<��{�ֱ�}�ѯ)��TP:�C�U��%<�8C&��IǓ%� �)2�f���iaqt����
��l'D���*P/H�@|On}2,���n��ˤ���W^����U\wZ�����ji��a'�,y��͡OkB���~�ן�J�R�l��p���u�1ǪS&)t�ަ�јy\�$�b�9�^���g|iKR$��P�"ݷ���d�;��o��V]i�_�\����r��fp�
d���#�:o� z��
FU\K�+��JRD����^.#Ӟ�*�n?����O�Y
�\����{^S�l`wE�	��zb&(�|�������b�"�&�-�0d��Pf�$���Y7�[Ʉo�q����f�?g!���	���`!<+��exV��u)i3$I}խw+�����{ŚY����Ą��F|-7�	�-m�9��,08�W��vG�u;C�e���ee�wo���k�?y�� �T�ҽ����a��
k��ΊϞGKmB)�E�-��O ���<���o�}8۝!�>#?K���(�;Oo���z�� �g���	F{�q�8��n��z�M�u~\zCC�b�i�u_ ��\_;��"l������2�}��% ڹ�c� �3��V�0�(��Yr�Gx�G� �%�n��$�P���W3��=W�E��� ̖B�����Z|����ul+��#*�w9�85��i�n%=+H[w��?Y�n:?�BT���p���c��q�YP�|r�㙻���0/����6���愡���n��k�[�Ʈ��
�Y���������]���Bp�{W����#�E���<g�!A��I�V���f5�;�h�Z�=���%�P�.+2f�ՓJ��m��n�!P-m�4�U���wo���7�J���{��䁻2n y*�&���k#�~�U:�F���V)�(KT�X%�M�}�6��#�@��(��ý��{1���L;�4	Y���n��K����Իn�������=��q��(ka�tx����o$�[Z�e�K~�Ί+�~![��}��#&i�e����Xi�����-��<���Q���F |�{*�th�ƹ+�����7[+�&w7)�k���[��8�# ļ���F��ϰ�d�1��_n!�u�`=��&Ɓq�ｵI�C��M�����}�Br�i}����s����"aI�_�<��A�Y�n�XN��m����PX��`hK�0kz�v!7��5��]����]���Ш����6��@��ȉ(c4ɣvw��R�.p�Hs nH�<km���jz>_0
Q�3Iݜ|��S�!�Zߵ��%ָ�[Q�}%[�I�*�t���z�C�L��m�	#į�qRu��%�$	0fηI���~1X#��6����cw�@	K�>�Pά[��8JaX�ST��/e�����""`��17sۖ���Os�U؛���8H���x���5���[B9��֩uQA�=#=�O����τ�6��=��E�dM��"?��VJ���S�?a�]����S�
�{�r�[\ؽ�����-���%�a��n�(�)�bѼ�P%Ƭ���m�r��e�[g v�}p�:S(o,���[�|���TZ1-��t3���eK._h�^�V��*绤�8�K���߿u�ʏ�ٸ�	�Ą_�/J����,��O���F�iK���ª)�[KDh����,&6��|v<��I԰�<�g;[Q��Ԓ��[I �bU�����u�(�+��oXLi_z��a����h��}������JV[Δ�}͐���J"%IJ���!�yj<Zu�&[�4��^<�<�`L��q7ɽ��'��y�>�S�Ҧ��8%Y�Ș���9TNK�}�6QP�y��Ԓ��	������ٜ�Eʉ(%V%=@~%�l'b~��Á��bf����7[�=�$���!Y����S�|�3+�kWX�y ^ؼ:˙�[�@��C����^� ����:��"�_1|@���}ٝ�ˇ�-R$4p�D�u�cx��T�	*)G���=殭�ln��N
��#yF���������=���������S;u+�a�t���1�e�?��.l[2*Z���g����a8��K֥�k[��E"A�V�R��wI�v���מ�?F>(��+V�!����+�钖�7|��R��
�Y�N Ş�O���5<�~�f�%1�_tw��Bcm��?�nO�^��Atޯ���x���>]�a�,����B�٦,\�k��8]']�nB�6��V�w�bz.҅�9�6�-n}S��aUl�� ���y"í����?'��"�ԆVNZ��v�1�!���'��Ei��FK_~�4��B4�-d�f��[�Y��s�c�v{���SR����ׯiX�����b+Lu���^���B����<j��z+��_�kӴ�au4�t��Z���g�S5�h�j��$�`@ޘ��/q������B��"��-]�Y���O�vV��պ�Z�r�jٔ�f��%�uV1�!oȬ��X�^r9����v\!����O�����rfrc��E[��v��n�������X�k����twsś,�3YM:�3\�\Vm�tqQ�܃cI��\�4(�K��X?>��m�D
��|~��X�$Q�G�ĵ�v.�W�Q�aV�PH����y,�_�D+=)u[GVp���\;s���1P�w�PW*�0�J兩����;�i�H�Uu�8�qi'���&Bi��ȃUR��8��LI��d�1$�~��Ы��<,f���)9��C�O���l�h��V��w�����R���5��p�ݚ��fhy�b����`�)��S��lx�A�K�C��h�{Av�����/�ä���w*�du������-	(ZE)��Y��~�qZ^<������6�@ݘ��ܧuǓ�r��_�=�!�脸o~]��h��w*��F��6�qʘ�s�Dh��fܤ.����;�|=�|qo`�0)h-���K��LI�۹��5����)����S��u´��u�qEjr���td��K�6�y�R��Ya$��kSh������o��#������կNBw����3N�gW�����!�qmV��8��U'm��SJ�t��@�M�qA:�c$�'�E�Ԫ�'�$B:�-٦פ��/-S^ޯM��UhӺ�+�!ֱ?9���~��`�'�����r��N�qi����͊y0\��*��?S�4a���t?Gۧ��	RdZ�ɂLe��pBh��+.?hf���A����;�(0�4B�ҿ��cU���|{Jr��ݔ>e�<�R�'j�=�\(�)�)�f�m��jnEWO
Ty�`M�K���&���l͛ݙ3����?V/��f�NA��ʳ?�rvk��W ����p�@�,\��[P6ٞt�8PZ�<��[<�Y�w
��5�Y�!԰��T8Q�otK�o�=]"���-�޾��пek<�X����-���ow%C�sI�PI�%K�VV2�x��!���Y�u�.���4(�m���_->���|�=��Ŗ�B4�Ҟ�V�u�ֲ���I��H�z9��ݷ��l��Y=�E�� ���/-n�g�c�����ڸ�u�x��Z��w^�k1�xM�n�����~�N�EK�ژ�4���}���ܧ��\�(!D)H��u���2�����u����Iy�������2����5&�F��I~MB���[z�J�	V4[?D9���qP�K����u���kSS/>��(!{L��(M�J��3�sZ�nusZL8l��U�����a���"5��� w���'�\����qa��Ǫq��İ>1#��I�m{w�����CQ��7���I�n_&�m�<��pqm��vi�a�Cދy��l�$v%T������ۥRF�Yq��˽�<�e���U��NqУO<��3��[��D�*(���t�vm����u��ͬ�|�� wQ�Cw��p�M�pZɋ',�����:����Rx�\��sa�Z�E���+��e!�E���smQg��Ù�M��r�/j���b��	���A�ܒ�$�/[,mޥ��g��O�H��,S��"�����E�J$���,{�j��5�9�DFE�"��ܵo�l^T|�����%%[m/DC��c07�ZaI�R2�2B`�����L>6>;溃m�٦c�L�ﳡ0�S�������\,��j���i����I`�DKqX�������z;Dꎉ7�bF��n�-%<n����;���c2���e�!-������N���u�?�W^���;~Q�O��ȷ�����c���,�z�=�ikN���:K"[ afY,���A�qE$Tx�)ȓl����r9�ܷ���}��ձ$�b�f��k�7N`�q;�<a�,���K=r��;��K���++y\<\�����i��|mEN�)>���~ug����}�B�_���k	�Z�1�lV���k�0�||�n	���!I`Z���gi�2]�[��pkj�xfH�NM�ckbg��,T��R:>k��6r���I��~���}��ڟ���C?&]�ӅRz��1�X9��38[v�N��\�h��y�#�J��m�,��ǥ��L��-�<�W�f����]9��w>kkݒTH����,�Ycc�VS�'�5&���b�].:7
��vM�-h*���+yM�^�i��qc��e�Q�ogE��r���>Y�or<�s3c�Q��V��b�箬8,�Du�^��Ỿ��R�ӗџ��I��{�ſE���C}������;})W�������DQ"u%���Ȑ�d�*)tIl��tV�v`�1��	v�K!z�:ޮ�ż���0�v���9��z�R�O���qq.S�T�f�Iıq�X;w�2$@��#FW_aq|���%�����������"m����,/�l�/���[���+�\�Z?�5</((��:�F@��Յ�t�zi�1����`Y�X�pH´nƷ�Ʀ�J�҃��u!ƹn` ��ir��]���q���:���j,Z�1��㷛��jZU���tm���L%K4�-I��:TXyqk��B���Ic��ֹ��0�Y��Ć���p�A}:(;Ko�lg�m�}�N��&�u��u_�X����Ւ5��3˗,�N�]�<������v���j≬}�3�V��~c�C%w���~����i[v��d���0�/w��0�	�,L��	�NX�$H7{�ZLۓ:i�n-Ү��!�^���u1�����__���V�W���4Ǽ��˂8�B� '�(~��%�����E�}m�[o�ør��r8�^�m�)��|����|Y�&��J����
��kI{B�:ۈhr�P
�cI-ea)�bK	�5KEL����r-�Х��Wo�_�o[��IB�2S\p
��j��[q~W*EQ�ll�^�0>3�Eg��Ǳ�
������h����+[&&ٺ�eC���a��s31���o��k���M�����Z��&�j�Lŷ�zX��m:� �����}��6��Xp�I����k���T̽��b/Ș5Q�J��J,e�[��[Ӆg����!>���!9��2��[oT��Uf�E�>ځ3[�I�of�?'���a�9��L�����J������g����k�:1� ���{6��q��\yI�1^r�;L\QfIK�Mփ��65^��ݮ��~x"�����f����zw+���?�彳`��P�za/D�s�s����������!�_�����VO]�G��ʢ�m�P��j�+��H]�B�v���*�!����6��5����^l��i����ic$��^v]���t��\Q���V�@ɦ�%7İ���v[�XZ�8]@�9�GJ�A˓k��](�˳���Y��ޜ�팴M(D�H�Y-�r!L��U�q.�3y�r��a��M����^�	<h��B}���5I�����{�dAJ!�f~����r���B��P��O�����f����6�m��b�C�ܪ`�J����.6$�z��ݿ�m��{�x��т���'g(�7F�6����6?��__�6B�ʥF��S>9և&
�L(�p'�3�_ 䨿/[�����̷d���u+H�)��x�n�%k����Y-��%�&��a��ܤt)DH�+E-e���*n�&�`�:�	>9��D�5V0�D�Ō������N~?��0�s5�\p�D�/&z��ox�Ͻ<��~���O.[%�s�I�/m�p��t���+�l����[����Ȓ��;�8�����ZZ��/�ŵ�ۡ���3�L
p�H
���7Xt�j	\��M�ʍ��Au!J�(���\���.!_C�ۜfM�{�N��R���B�Sم��-ǔ9�[!��$��nt'hZqNLޏV\ý�P{�Y'^������P�;&pMh�a��9W�ׁ�K������3Յv����9�4�y��B0Ϸ�Gz6��?k��<Oc��t��p����A���ds�^&t�T��
�笵2(���/�D7��Ğ�9�'�}�5h������4�k-��59���g���|ie���v#`�5o�w}��R��H^�� �n陂�2u:A	��������/{��¼�ul������][�t#w7d�C����.m�.f�l% ��\���� <����۹�J0Lm-8�ݵ��F��8:���*Y��r�����y�e"b�C�R�_�I� S\�;��3t- `}n��z�����s��P6��gb~��K_W��X%�z����♙�c�_����Tz���.ν�b��m���ykj���6@����q�S}��M@���Ak=��W�aN���8�s���E���k��:�{�:�\��,̻�l�B����ac�O1�R����|?�Q�1�yp}?P1˾� ex�|��b�4������RP��Li̍�F�׌)i/HC����aQhL*L����M��i��?
jZ�҈���$�пG����7�~㤂a*s=�r6��$��k��GO�kL�iO�%�qު:%u�N�Q��T�&�{K&���-�S�z#�
J�^K_=H��/-�x1(�& 0}�L��p��X�9�u*�bB�2���'߭@]||o�bW��/�W�9�fA{�.Zy��k�� R�%!��讏��<�_!X��L�(�f�\���w]g����i��#t�����wm)���7�Y;�0,X�hlX�ǔc����|D�C����ެ�|��]�~^������M��Ú�$���6B�Z��?��F��l�~�*�����1Hդ��b�q�)݈���-j����4{;z��˽��m���,Rlt��"�ԛ���H�J�i�0�p�p����&>�K��<iF԰F���0��w�a��#�:l�j�X3�~�E��q7M�KyN[*ڣa��ɉox��p[bc�U7-*��l<9�#���a]��"�`�iU�8.b09Ⓗw�BR���^�k���7>)�R��:/w� ]g���ѐ�Б�ϫR�8j-	r������}�DV
�iA���	���=� �j�Ε��>-��=t��B+>�\ׂ��i��ZW��т%����<;l~>�]�=��^����%������b�&<0�����P��g0�C�W-Q0b�t8g|�E�'����9�=���ޑϟU	��w���2�U�2�Ie��1=��ߛ���!� �4��f2��Q��b�L���B3��H��dS�����v.���P$X��6�bjrs=c\JG.l+�����@�T7�Xn�P Bi%+�DN��o��IK��،/X�� ZH�T�,���N�����, q��g�5Y�ys�o���b{�G���f=)4�dt�U&nּ5j��<�)3 3�����g(��roʩ���q��Ly�r̹��J�A�����x~U������rx��xx�?��
� �B�;�I
O�cd��{�����l��@��)��֝��!|�J�s��R����y,N�>S���6��(I�3iz�nQ6D '�g��d�*�΄��k��ܢ��9�H�WV�n�|ћ��a����N����-��$*,&"Jb��0���C��j��0�S��$�ݗe��bN�d|�d����~��|pC����Ĥ�6b�ɡ����#�N�IU:��QK�W��)�%*�B���!⳨�ƹ�{�J��a>�Ε;��ٞx��ђ�1�T�q�m�����[i�!�m�dj~0��W��V�rN�>�sţ���[e�9��zc�J�/vó�o�,�.g�k�F���Q�a/ip7sR|�B!�1G5a���YvM�خ�@���اW<�{���
 ���|�!Lq���M�6��p���+�a�u�v?\�����V+y4�FK֫�u������y���n,����is$I�,h�GD�̣���fEFd������ٞ�#�q��=W 
��YU=-��"�p�(
s������R���hǞø���up�^�&Q�f�+y#��а���l1��W�I������@�{���!���Y�x��O��&v�Wl�h���t�3-����FŒI�dz�\�az�p�Ս5��j�j��*��5��h�޲������έ�w�z��E�.<Vz�������7C��rO�Ets���{}�l�Q�t���5^<M����\?_`{�w��_�����r[:.���K��X���6,�&Ԑ�;�Զ��/2oM5���<�ͨ���
=�>����hܣ��m0�j��u\{�`]����P��)8���'��=�
�U����h��T����`�r�u���}����mY�xT���P������M~�d>�rD�v
i�)oO�6�����Qjr�c3%���b�������x��;C��G�e�X[?��'�>[ܛ�j�稗�IXH�̇��k���-	W�s��^fw ��`ה�M�t��+���"��"a��"灇[bY|���I�=��A����8���o].�d���Ȳ��iƷ�T�w�U��U����[���9�y�{�ĿG��Z���o�q��t#eߝVV,�X�r.n�w�%��-�L�?2�����}*}�L�m%���Ɗ�s�Դg�0���l�IR{�m�=Ri��KG�&j��{����3Ȩj�������$_8�������2E����"Ch�N��	��NM�Ƙ���o�N�k՛�	%0ѥ�S��x��I��J�c.�j	�V� �]����Rx�p�k������gb[O�h0>��ǛP�׼ 	_���'�y�Wc8�s�j�)�*���p�z8Fp_Ǐ�"��6a>����^W��C���W0�Ϻ�҄�a��f�L���u��1�����H~����㗚9��nz#��p�<.����4��a����_�r9�y��dcd��ƺ}����H�u3���Ҽ/��dQ�0��
�
`I�hF�!���k�<��g6n���`���:Qa����9��~��x�)`:y�I��}d>��J��wb�;���=1Û��W'0���9iHڦ0��H�R�Vq3LLd�5�[�h;{g����Bǎ����݆�'#'��t�jo��x��N�f4�5]���7�X����P��U#�d�q͎V����J���z�FF���������Ch� �f����ލ��s^,�c;��Z>�yN{�S��mc��ĴZC���C����#��5t�V�(�H"Ft���0O��(����Gnj��θe����U9�y<�'?������a��~�scw�A-��㭅cza�l��Q�=�ŝ'�e��&�cz�;iZ���,_kJ~�-��U'���ϓRH�ǁd{�n;��;[��R�U�8�>�|�v^k�4����u��ۊ�>M������27?%Swm��!*�5	��E����K?A~�����\'~g�����������V�<�G3<pH�_�d])ah(�~dѭj��� ִ�J�����'�<�f`;3���/å�y�`l����-zb���f�O�|pѦо�WSk�M�ළ��ɆԎ �Ӝ1֪�o�y���\�T�c28#"��ݫ�mi��ܰ���C5~���>�a>�k��<�H+���t�3e��Q�i�	��d��
�ǐ���y�@Ư����T���׶j����T��dL����� 
�j��>�86˜�Q{X�^�b�"�z4U� ��K�����N���qW�g�R��ww�+0���kyy=ˀ�ܮ5��;��2�pBj���x*����+����/(��x:V��8�����/2�([	q��yNѲ�m�=�&cYo�p���Y��q�^��&UCf]�8ݝ�����;o��D�-n���Pŋ�����k��R�R5�=Y`��h�݈��߹S��VPQYXaT��ZhW������bE���t�z)w�q�'���{���}ib)�Y�^��I�M�;~l��^�/c��`�D�#0{�`	0�f;�y�H+�i-���F�v�z$�ء�m%A��N�ӂ�8������+9'�����<��Ś7�k�j2�y�Ѡ;c�h�Afw����G:p��b�1�Q��Y�[9�/���7Y�>�� ���C��V_|�v�]��P�f�����,ľw�׭1�䍲e���1)݀صv�8MX�ًI\�z1JТ�{0��N��ha�$7���=P߽�̣,o�j)^J��>r_0��a����� ϯ��i��#è�(h���P��`n��(�x_�x�~͌B6;t�w�Ig�E�+Ƕ���=�\ڗ�������&�TcX� '��6km�[x�o�����0��}y�}1�SZ���8���%ъ��;�����ی�~��z���%:hMG�=�5��_ܰ��D�ƙ��\�<L~/kw���d�~f��ܯ��<�"p�A�;��`�yBRP���3-�<�����|>�o����v��E�ԐN>e11�RJ���>��j��^� ����H���G*���A��d�Rո�ܒ�qf|GU��X��q��}�N�&)m�!��R�E>on�#�@)���f���Is��*=�|�;Ν�H�!�]T!:6��M�573�BV�?�#,�a�E��+���7D���;K7�7�a	o"��z��nz�/o�LM��ae�5�B?>�4Σy�摒�>K��������tާT���~���2��1���.�F�օ�lcU:�?������#8hr8��^.�r�^�7Y�R�m����d��ì	�:{gL$Ҹ�"~�c�(��Z�i���Bb��lD��&����GzΓ%s8�z�~&�+7Ӄ��g���4<�ͽc<��nv��1��@���p+A����nz��HI^71g޽��%rc�Q��/ylQ���?^�]R�~`���4�ؼ����uP�X���Y�-Y�dh�d!����2�֒w�)����1y��a8�[d/���ƞ�9����%R��wx�ك�7�ȳ�q�J󱩴,<He3��4ݓ�WR`����y��Y��&*?����g4��8���Lj��� @7.\��#s�BN��\S�zDX�V�o�2)<X��H���?��J<yJ+��Y}C/�������aWLN�{�Ѓ$�	�p���=�E<�)�@�=Zۛ����Mi����l�� �k-���P��2Y�{�����B�h'/@�ƛ�]�����5�����Ʊ;��o�L�E.o=��PLp���=.r��sՊ��T�--<���z��5G4>��9�98I���7��d��H���pU%���"c�wo:P:1��O�ӜS&C��j��Ox@�9��{
�Ժ$�[�&u�kl�L�Q�J�u��*rĈl��d6ݘ�1��W␠A��ܢH#<��g��z+Xn�b����8/j�K��,���Ui��kڄ�>߀7��:o����o�7s��z��Jr�Vh3�B�K���fQ�x���l޶�������	�P�}K��������c�헭+̹}��߅8u�����[T��[C�F�����.�g(�n��5�nHØ��F�V�7u��`}G��A�8Yt�	�)wS*3uO�C]D[5����ڝ>�~6u,��"'B�6X�`�.�A}�8H�	��ͷ�8���v/�U%q�0��ǘ�'��F���`0 �e�6VH�q�ym���p'̪�����$�3����H�\���%iJd��Qb%�H:�:E�&�6�HhrR%djHk6�QeC�ϷЫ5�k�Ʉƹ��t馓R���D��rc��1]k7��!�0�о��q����m��r��xj��Λt��zc�9��go�d��6�����{Cnr�
$�Z�ļ�AE����N�Tɭf���qJ4ɁND�����1�s�kU+�v~�G(��7r��t%ɵ�`�R��"��L��V�1->�tq�JO�'��:,� �1���ry�څ�#=J�Җ6���?}�W�T�l���&]��<���n%�u�|���H6��sTC�
�&�������'�	�L�=8�c
�~��-p�tU�1XU1�|O�w1`������q
;Bi���wg�5�wa�m�4
�$�u��j��,���&�N����W9P�6�.SF�x3.d
�=3�Z6���lC�|�1�H+���f�Z�c����hq3��M/�jl=������Glt�v5N���i2B_5�I�%���ޛ��ȇd������'�e����~}�X�C;�;ʪp�;Ҷ�gq��"���%�b{!{eY�P�'�-"��X8����J��ݵ� _��:3vH$Cl�L��ր��<0���E&�浓~r����E@3�wS����C����\�"��h�7n��0�dd���Y�<���(�Z[tb�b7Ő��'4�ܦ���`�@�I^��p]���ɯI��YP��I�Z
3�h�����1(�
��*2&5�8��HqAf-6c��bx*����Q޴�ދ�{x�)t�����
�7x����5���}�Z����m~��qv�e޷{�o�¿%OH�1U=�n=��u4�3%Ⴑ0r=�OR9�5C��ᑾY��+퓌"b\�=��9�g�L���ҭ:*�J_�����x	cB�f�9�!�AU��u��t)��bʊ���%��@�b�c5왏kp��X�)´�K\�i.|>�0�q�17Cr�a��e$�S� h�[�t��.P=�U,Pή6)�G��!�U�Q�U�v��z"s�<5.��,�u������[EGe����z�P�м�����4�w%�?��z��k�HxKf�0jY��OI$E�3�PaHn�m�s%����PNB�^��ol����c��u�rX'*)$j,7�<O��o�	�j�9?���w�'�/|�Ͻ����2���[_��8vy��n�)B��2T�4h 6���!L�p���p��dl�|j܂M�_s�g�1[��|��}O���Z1�01p��5AHE��"2���['�4n��B�x��[��>�rO��C�����#�7�P��*�o&>Ұ�%@]��!��Uj�등��KBGX�i�y���<RN$���$�w��>כ�Иxn �J�/xx(���؉Q~4�\��4����)C,�T�hf���8@SO"�1�vJE�ND�(�-4� ����c9���u.7�\g��F���,��c�O�I8-(��\M�K��j	��O�b�y����m.n>>�Jݿ��8�{P�1N� 6���o<]0�Zx�#�DSa���z�>�{��*{�\�������8�`�Y�R|ml��.c9�a��������1������e�I��k��g-�%�G�=o��b��7��A���p
�TC�M�z9_��`��PU,P�~=�-��i!s2����pf�X�m��u�{��5��)m�����*��^������g�qX�|=E`�6G^D��S\S����,EEџ�n��7}ǐ�Ɣ:I6�VȻ�����i����M���!17�P
3}��I�_|v���Q|j��Z:������	5i��a�/������V�� �}�n�T�W'�y�X��C!_�)����*k��yo#���m%yڴ7��2��޸nK�;CԦ���jrЉ:�ag3�H�Z��c��m��i�R���i+�ޗ=����!������[���|�3���ւd���Wu����e��T�l�E+h*-�{4��C��.����������x�#����Z:`���*c�E�q��1���"048��L&��9��C�ܟ>����$7��'0~��s�ڝl�٠m����G��\�Ԯ�Q�Tf-����0������y���m>���!�C?E�i��(	MM)��	B>�OR(b���۶D�/���S�T�eqT�	�t32Ђy��#�n}L���l^��M����	�V��O+���$�4q�����j-�:F������'�}�|����kzH�0J�Zk3����ń�n:Q����Jx�@6�:�]���W�Y�p�$	G};m��(�MC:��9��S��}=uV.>���iM���X[�Y;�l��M6o���Ynn�B�B-ئE'�q�)�5醻�"!|-[�:r.�2HZ�wj����e%���B���	�s8L�U[��][���F�����W�qwh`�B�dd^����Z�F������{/f�E��eI{���Ң#��\]BѬ��w�6�j��uɞ��.�I��f����:�mҍs6��i�	c��������g�c�ݔpIg��p������mT6�]k�!p���&M<��~������s<���h�F�"�(A�H�s.}!�P"d��+���[�ߘ �o��Q��#W��,c)�m��u�F
[��a4V鸯��Y�1�Q��״H�����h�g��G
��u�ʵ.Q�UM�l����-=oFFEľ�7#���Fm�)��v]�aY1���L �[��7�%/�<�:��c�Qϖ�=�X3��q�m���O�y�6���\�l�ч:0�0��!��O^dA���k�YBWx���?=<�ǇG1�Z�t���ÿ֋z�X�K��'*�N���71��Ċ�~�������)j]��6�)Y�k�&���"���1撠�� ������u������T��Q���/p����Y]M7us�I��~]���z_��Mx(R����o�4�sS�����W�@)yD�}�A_�<(��W%qrh\�)�e�w�V솊Ey*�h��U'�
��S![%s~S�D�>�w�<t�����V�o~A��N�DR�Ę��o��v��l ���"�h�d]���'Ch �s�pz-50g���j2l�8���(y�׽�͍�!����(̀I������ox5�7E5d��։&��1��\9��Pq�Y��C�����LOQ�n1�-`�*e�V�����9f���\�4n-y�=v�]�l3r#�������y>���nH�$�G��g��.9���t:����EئhS<�ٸ7�?w|Y:�}׭0<��ë�)��H�u��:�a�'yL��^6�	��{B���ɫ�l	����)Zm�!];�?��Ѵ���j6m)l��:P�n��M�`v	t��08������o�u,Dnx9rN"��kv��Z�a��/�K���\�wߞrb�	p�D���͡n����L���4x|,�?��Fy*1�4���ކ�<�O'�Xs�{�i�_�h	2ҿԫX=�u��Ĥl�/�,-ص����?�<t��ɹ!}lH�C�_��Z�9���[��L���ǋ�=NɅ�#"�2�V����6�蠟��=l��W��z�gO����D"�?�BӬ�Pi[��G"�Gx��ON3�Dq;���í�vÄ��1�W��%r��^+����`y����=�o��������[5�Ֆ�PWp��J]{���i?Dp�2��LʻwO�0�����(��h!}���A�Ks���~NQ��tYR翪T��I��Q�z�ɒ�5	��m���}�:�B�(�1X��h�n�!��<���t�:��$lc����?/�.ɵmq�ژi����^0�%�򊐫w�}+�8�8��݂�ZKN��S��i"(>'���11��Z�jFv��C:F�αɎf��5h��m%nv����r��6Y�Rh��A�xX-^�4��@�v��*R��Sϰ��[K�wx�6V��>�C=<��tٴ	�7���go��1O�ؠ�jIj�[��қԝ��� ͞,�3�3_1���z棆泊�݈�o���b�Z�p�Ί���|PĘ�w]c���*���0�`��'�$Kn4@����� ><e������\^ϯrZm�wUq�pH�)Q��=X�Vɕ��0~�yO�$<Xї��;����Y\hH���<�Y�xuP$�/q*�r7��b��ςk.s�;U*s�&3
�]6[ t�����T���v?�n���*�� ��/f�.G�q�����r)����^bb��E� ��� \~u�h"����)������� ��'>8\���Ky}}�n�Ѕ�Un��{����]v�w�qc8�U���ls�%0�[?Q���ϼ����U�k[;cPn�*k�{L;��t��*N������+�@�u�4��Wk��mo��޳T�}s|8��X)�!���S���S�98��f��u]5��#��p�D C��/�C�=X�x4���Eݯ\o��R�	�c���6��{�6�Q���Z��`��Q�߇�Q����_�hJ�==�ǧw�Ib���|��y~ѽp�:l�kWC� F�TK8�Y�$D�SV��XGeg�J=r��ޖN�K��Ѕ-Ns��v��ƴ$�I+��9�)%&%y"v�$8q[��ٓ,��>4RX�I�ٵ��g3̫W)�7�gcS(�xG�d���-<�������3l�&�d��A���nt��C�\ݱ�dZA�1kzeOO��d��.�$}��Zܐ�"e�e�d�mkγ�LC6�\����q�!�Rb,�œz�*�!NwB���E�0
a?cc���H��0�!��҈F��p9G>D�){��N��-4��A4rJ�jQ������F�!V��%'S�f�0�����W�A��(I�ꡋk9��bL��S狀q��$]v�H'��a�!&s<z�?�Q�b��j�N�����Hk�������q���MUClN�x����`ى����;M��8��{�u^���~/���L�Z�f�iH�C��'�!����dУ8�i���A�|��x<�$
��BaL���t��K\ļSV�IW���(��А
=����U�Adr%�D?n3����&��&�8�B��և^Y�0�0x�R��M~
4rT�h�?���U<��݋TC��1X��G/����-|r�iT��%+�U�A�I�aBY!W��A�����Ɍ���$�!o_���Q7R�/��׵q��P��N�����R7��L-aM���ᘻ�:~�b^ø�G�����6��+Ly��y��<�A�.'{�}��,�j�{�!'O�;z���1��6���a��n\/��`��7�������;y�˾>��A�Yts8�-�I܇�5��I0|vvbdm""�(�бT1�e��9=�v�q3�_2X�d5(AԬ|]�>�(���_�e���
�����>��-G�.`�bF"mo�^��3bqb >}����?1h�V�����<~�=�0�������}(�?|�A{y~1
�R�a��)���BL��ӹ�	I����mnɐbR�*�O��w[nI`��KlDCBٻE��p���U嫄�� $���E�0�O�w���������^���˳�%�3�ٸ~Ś��c>}��U�c4#�58T��iEq����|^��F��?㤪N�!%6�B�}s��8��z��6����Q�s�`�o,6-H�vx�H���b<}�G�}R����m�,v0h�U ��24){p�+;֝rS��@��	.�W��bv�dQ�L�G��G��_�e�Z~۟0,�������d���^����*c��O?���姿�$k�����|����vu� ���[e�æ#�Ӈ���ֽ����k�Y�f��}b�;�{x�N��k��k{���������lZ:��8�:�s�v��~����b��#->G>g-B���} �z�	l���?���~�������ʏ?*xm2�lO���O?�(#���r��<�{ŀ��|T,�h,ojݙ�!h͊2�v�Ԟ�}�#eA��&���� $7r��s�Q3��}��ޞ�����o�ʷ�����lsߔ޾	���'K��O�>��O̛(����i��wb�_6����b��C�oz���p���y^��l�{)��SO��z�0j�lph�@��+��5��??�:U�b�sz8������w!�����G�أ�֞�A��"��{��`�8`73^HhH��oV?Y�S����Ō�Ѱ�l,e-,#=��*!�a{R�&�ڮ��s�1ߎ=����G��3��Z\���ע����c�����������|��ɮ?}��B8O���dH�PgF\��;��!�l :o<<?�"x0���@D���"�I������U��{���2R�_�G���2�He��4.����c��V�I"����#c$UtR�2N.6���]=�OHÞ[y��,�m��������ᓉ-t�LT6���jwxf��]��X��^)FoUѲ:>祥�:
D��.*X2�G���!8g�X�3��aS_�
�`��A��$Ԥa��ћ�:̂'�x�%ޝan�v��V5R�/�R���H={r�
7Rº��M�4�^��7@5�kZX��9�`qÃ'hF�l�2�Ԓc̩
M�����`쿻�F���AhH�`��s�#S���4�LFn�mrLp��-�Gy��p�/q/>�C�@։ϛ���e*��"[�ZsBb�H(�����U���c���
�~4x^����u��gK\\�>� u�������r�R4��!�F�"Z��c��%AŽDF�x���*s�j2�N�t����ԦUpឍ����=T*��UǠ�a���M�Ի�3���Ih�Ϟ���!���?5���:�<U�.�S����<������������+p���\r��:Tz0C:	cݗ�S���.�-e2�|
>ʤ�]�)�u�[bߑ=D|��R�9�r<�e=��NQ�G�b'j��3�a��$`O,P	���w"�y|��8h��Ռ؋Q���r�=V�(���\��)��*�ϖ0*�F]"�J�_��t��p����]�ȵ�3��y`(�&^Z�nHcQ��x�����E�Xly�]�BJrjRc�愣��-�_�rDMa,�,fx�:d5��n���7j�����9�[Gwn��G޼�f���ݷ���T�������<��E�ȋ997�b~�T��5����8@��m�9���!�i�Q>��aH/J]�=v!�9N�e�ZU|Em�;&y��J�E�๪NK��Mvג�;J$L���%�]��{�?1�A���ΒC�p�|���똹�T�U���u�_^�5�b� �(�
���!E-q2���g�h�S�yO�*L!8^b	8md�ODl]Y^K�a�/���`6��'�F2-k��O:|�p�C=��&�&�N^����F0�݀b|x��]��_������>��J�b��RbV�*���!�iqc��?��m���(���qS�_������ �������|�E��Fr+�/q�th�#e#��5&���:�����7)�I<(=��(i�<��+Q�Jg��lГk�g�Yb#�Ԩd�ݥ!]Yqe�ˆq���נF���H�,f��+ƪkkp�e3C~�7�c!I�@o_�}-�y���kt��=�Ed�5����񮁙ʠV3�e�>��'P�0��9hԛ����z8=zv&�/��Y~'���8����_#I�'�	�O�R�CS���s�J�=��dG��l��Q���N%H
��/)a�
���'���̗�(_�K��b$N��n�?�e��c�Q@�$�d�*߮��?�MM�d���XӶ�)\e9+{��*�=ı�hW�H,vꍗɿO.��XV�dց�	�&	>p���z�������P7��G��Ȯ�m�n�R���)Q� �J�_öJ����9����n497��3�{xx�J�^�Qw��9�lw��I��}����9n��W.�u��dΩq��6c0�S#�E�݌��ǝ����b�r2)�O��m5�{�l�l���b��>:�c��+�����*�����E�&*m3���=�,������/��
a��/e5���E�A4����[U��ƍ|Z|Da����a��sX�pp:<��iV\y�<���c�3�,ɻ�������_��:��\�DL���~~�#m�O���67��w<�7i��G��۽�ڂ��fx�U.�Nh؅�篂���b!�bL�=�t2;9�.dbD�au�!q� �U>�L^�nY��I�S��D����I����F�F���c7i���MZO��J�������sx"�E>�ܷ!�T�),���i�!T�b]LX�Nr�~�^���BX��_�xtWgxʦ%�D|�m�`��Hn�]q�n*���լ�x���#�K&��A�Xj��f��<@�\Z����u���d��v���TIB���&LpЈWvVO���>g���S}����7�MiDy�I�q�z��-2/8�����I�FAK������j��8������G��j61���4z�I"7!ѻP�y��,��97����e������^4���If�x��ι	�#�P~�&:D����H��<�֭�d�����7�z���d�5.�$#�i-4��]�x��i��Ž*�d��=��@��F�P�[�|�O�|���q�M09�M�{�a,6!L��Ⱥc���7�-o�L�r�y���r(��x�-YiZ�������ӧ�f�aV�|�r��h@�4M��`¾Bl�1��y�-��U�V	�$�k�C�d�?~�Pϯj���F�Ϙ��ō䇌�E>G<=;X�y���0�k�9ε���!MۡX�Or���,�=$�F���o4��Ҏ�&_�	���v��y8�a�
����'r&mb-m����pzsMMf݈J�
<=�=b�#K�1ڿ���"����4����� ��7��6���2O]�L+*�"J[�(Q�?F,ǣ��T����T\��/�3We8M�mƞ��B)E��<8�z�NL.�$^�{�k"�>h�j2�F�  ��IDAT(�aQ���#�!������H��rL�p��\F�L1|���T��U�q�-N�%Q������1����Rb�F�q�s�&�z��04�ѱ���y�Y؃O�
�0mf��\I��]�=�v�l��Žϩ�"?�;L�_�;���/��ɸ�g�J�!��T�G�G�S�FL>�F��W�tU�ep5��0���q�ظ-㎃I����q ��^@),�����Y���Q�\��BGA�m`I�����l`1��u���V�UÛb�P�ƑBgH��� �g��5���9�R��2��ݶÔ49`��A��t:(F�q8��܍�վOp���Y����n�%��͍>d���Ðխ��rb&�nr��ƙ&�	5��>A�-���{gd�0�e���d\Y٨����OX����I�~�a��-�DƋ��\N���k]����S���P��L"؊�!=4�j�7v��Ho4;��5�#M��w��?N6�"���la[VDl���C	�b(��ms-KO`,���*�?}*����S�O�0�!����I��O�5��6�]u{��n���y��}���ӫ&v�0��l��92A�;�:<��s��u�
��d.�� o�J���\O�E�\FjP�7uUM��#�<*�G#�8h�A��ɥ�X�"47��}�0����I>�+¸�_?�������`����p7��vik�Ս-������������7$����s�+~����XIfj�Kc�;���<t{�D�Èk��sN\�<���5T;�q�/��}�9�p��|G%��
���$en�1�	mK�HBN|�R���d~����Zx�x/H�R׾�7�*Q"��
%����Za�j�bo B¾�'
c-9�w����4y�#Bv�l��B�ª��~�m_K_���OO��8��� [�KC��
�������|Pxg��xs���4Ҁ�K���5�Ӭ���W�w���b��?#B�\�����?�s�ր���������2���f���M���d��.�ѝ�/w�=ޕ��M�l��%{.Y�W3�f������p����q�-�Q�adH#Vc���j/z�P�/�X3��4�G���ٱPO�䲬�ү4�/6<�Փ��Pl�]�c�da?I(�y�>��,?��6��_�(��L~�hFH�����LmL�_�s:��Yq�bz�c1>�@�b�������_ZoD�v,y�qW�8j��g��zY|8��ϳ6;��%x�0x�V���V�&W%�@Ė��;i>�(�{���t;� �����7�}����zR�m�T��~���y_��0�r ��Df[��h$�f�����X��
皑��d����vu�'�>TQ}��rgA+�(b�'>�
n��$��'ג��>&W��`aJ���@&�)�N��'����E�Tk���j��چ�Q)5Q���H]{���֖������c��ݐ���G��U�^��?ݳ��j%�����g駏�7S�@�������q��7*���mS����3�s
�O÷?��Η��R<%udu�e���)4*����^����g�����>_d�iS!�K��܈��?}�h/�{�4⯬�ޯS��}��#uQ+�ݪ^�E����]�����wØ~e�������I5�;)	��U�	�S�CP9�7�-�G��D�R�Q`�f�!顶n�f�b�ɀ�]���deV�>sd��-���FeN�F�{�Rا'�`�P�bt9� |qD��IAX�����xW���?�u��g��RR$�=Fy+[��d�GoU=��~��za8�+|2.2�M����<�sk҉X<�ZH��}� \�1nl�E4��w�Ϗ�[&V��kP����!�=��n����K^����'O/I��Bt�@i)�^,2����[��@�B�y�����$���#���Ӎ�!�	'���7������O팧:�g��j�#^�>��8�f��!<M�Dm:��ƶV*w��WJ<2��9����t{,T�"��D��!n�9�u�'8�������a�F�����E|�8�Խ�b<�f5�v xv��(�*�*�*u���fI�Cx���R<H�����i�V�yS��n��c"���嶣	
J(�u�C7r&aD?��Qx����(��i޽)�|�����U��%���&�Q9�jH7����.a�x���%�O�u��\�Z���i��)Ҋe���~�\/J�y|2q���֮ςJ�r���G�N�������ua����t|V��,���eJ"��L�R��T��X�,�(�L��I\��M֩e����[<	����V�͞�А��(�9��E�M�d���a�Ae�>��^��l�G8�,�F%ԇ�zh�~�)������͇�����{������=��Y8�?�?��*��ɒ5*ް�������s��b�%iY�Z��C��x���Ԑ6�cB�N�3k�'%��q*������"��SH0aS���ּ�3�_��<[�':N�&�p�_>�*���P�=sêR�R��+�QN�Q�s��K����a�7j�0��$�?j��%8&��{��^��V*��&C�,Y� ՛��س�4����Ud�?��IgdPђ����>X�IK�:�嵑��qL�s턈�s<�\�*'�a�5��=I�u�p�
�7�ֿ7�5����d8�0 w����I�����ɒ�����<�ށ�U��I��ε���0Rή�tͥ�X�29�j����E���+������s重A'XCGK:$2$�����k�p��Um��������`D�s����ũN�vv@�b8Ǿ�CT��̠�4'���,�ɉ�Z����#����d�}^��E�N��T���먅�~3E!�Q�t� �nH�R�*1�~�R�>��1�$(�p��f̬�*ݤ3�����R�
!����\��"��'_H�WE�y�[Nf�����?��_>�2NM�֭t�qzO^�#����&f�dQe��/?�"#�P�Z��c�a����@�PZP��0�2��U�_�TeId=� �ֵ�ٓ	�"� ��5��ʁ�������8f��F�h]��.]�L0#ſ��/��P��Ƥfu�����ϟ�U�����Ce8Ǩ�^p�g�7j�z��˷��7���@�	�A�Z��M������f-7h@��m�oI��\J�e=�`f�X�v��y�p�G/l�l�(��J��S2�z}��g�ޱ���F���!�E��M����܇���������!�R��s-��CR��%앟����ix�rt��(��֍�p�)�߱��5��m��$�9u��8�۳!�)s����1�[#�{��i�]y�u���I	)���m 1�F�Pu��gkU�]�췔e��^�)���'�X�:/U1�(�PK$;`p������^�U<2�"|���er�dz�T��=�	���'x�P���G�}�����`�jD�������OfKz<�l,"�"t��Z2��h
_(���O�)k�W!�_�n��]��a��c@̳*�� �⬙j<O�	��c��ƨaH_L�t �3�-B����\b���#f��XT�9�ƽEϮh照����=��L��X��d�[5��m�St��N��Ʃ����c��Eqf�-y�ԕ@� �]�%�E�\����h�&��]�L���9O�g>
c�E�uMH��Gx����mo-yÕ̍�Rp���32���6m>W��dFݒ&�����$k��k���B�u���Oz��ʆ9�B�p���yZ�uw�O*h��B�u=�����{��rk,
iN��u�Y�P���o�Ye��@�|44Q�vR��8�I�t���/j9�Si�ߍ�Y�ߑz9�C|\�ׯ_$)�m7N�߽>��Y>�W��:���e��dNVBY0�i0�K���J�Qx��H��h�VJ�kٱu�.�0|��gfE�_A�bC�u4��Gz�%��Be9"Ssz�m��)�	~�"
M�qp���k�BX���US���
�l	h{e���i�Ģ�w0^��[�ډf�إ��_S��Zo+��I���fFP�mR�����wL�9�@��&t7هK��л��R6��J���;�>�á
F�e���&#��{��G��6k�-�ĎD��TY��_�*׃�KR�����6NO�G�\2�ץj�
%��p/���U�C,�?0����O��@��T[��kp��5?M�Q�c���d��dڶ�B�M[Q<i��Rj�������Ré��$����Ɠp�{�È���{�\�|��Ѐ���e_�ʣѾp_���aKT��b�Q��X�Ij�.��{Ql��PI�.Z�c/26�s�T��Z{��]t�Naf�1/�%�0'ӱ!�i����z�(x�ŧ��PxCd��� =��J[�o[ŏ�Nso�c4IB<��h��h`���m�n �S��X-)��}v�9����q>�~Jv���f�B��m ��*�}7�-�q-��5�V2�T0I2F�)v��o=Pi6stn0�l��m0O��Du<TpdQ�e1-U���`��:E<���m�����.BWk�)զ��#��f�iS�#:'���ܨ�Nt~Uj�� �ѓ�����ɸ��`��C�2��L<�0KI:`���aSO�7�J����=_:�U�
R��g�?4�>���`�}q΀c���U��&��U�y�Gg�2�����AoFg��j��a�5�p���(+r]X���e2����QzLE�.I����"�Uct��	HlOjܧ����U��h$
N���ő��D�5�A��{�hK���篠 A�D՝@������ڷdSE����8B���<*%�F!W���qEpS4�!���/hOtfu��кB�r����5 �
`<V�T[�i�c]͘�G�%��>|f0z�� 	��)?�f�Kz�R�j�S��r�A~63"��P	0�(˵�t��$�TŐ��)�����Zy=E�Kg�|kt�b��U b�#�G���<t��₯j�oBkB/<�P*�=�I���{r,���;��R�E�*FL [��a�7srD(����x�4�3J`�O&��ywN�q<#�!�ed�������jT���U���.I�޻*��tk�A��R�̺��X*:��}Cٽ��j��q���S����yk�9����e[aj�@y�|@�4}Kf�J�|�m"�#��2�A%Ho��R��;zULP�~���^Y��S��B's�Z<7�GR�Q�X��+����jNx���{+N����~M�e��ɿ5֐7o�M�ʆ�:[$�(3T���wjZz�Y+����g҃ƍ}��`�rX����U*�t�	�ޖ�{3H���ZJ�����>D�k٠�d���P���b<b
���QHjm�5�o^�!�;��ټi �!Q��x�E'Ka��>���(���1q^sӡ�<�x��ڇh���z����zc�1�f���+�3Z�O���OW�Ru�K(nZ��J߫	&����+��&�\��Q�kkߞ��H���7���n�}�lָN����q��s�,�,3�Ÿ\p�߽S�(6�l�)�m���������o��vF�a�z>��Vv״�mz'�7���GO�I�#��������8�[�K�u����\��U���M	��j5Ȟm��Mۙ��#�`�(+X8�4�d��G7mӪ*�<0X���>��@�&n��^����}Υ����*@S`of4�����zS�[5�����G�K�Q]���iꌌ|F�L�=�7�o��Y���U�"�roվ[J��ci�=Ɖ-vrW��D�����"�
b�jݵ��X9ׂ�i=���M�ܢ��`Lp��lO��O�Ol��uc$J�c7R�o���n^���]�������6ڰ��T�t��*Uj��Sz�,�&��B��՘8 �#��y����
�g�X�}�l�LN���yeӦ� �]�[��݌�x��M)�˦z<F�1����
�"~�ԗ��Z���}UHk*��p��vN��Z�H����γ�d)�N��C�����+����:�x���@���*��Fw��pc����\�1��#94�6��Q��D)i3G����P�d�#b��э���D筳sPA��a��,��q�6L�P1�Q=X�e��N���EI̚��^ǌSJ��Xo�L�ζIyBx�-%��5B�،Ψ<�D]���@P����'zyLv�CaHs�?�!�Ù�Wcr�= �3�?G�����j��MW�V�kS<l���U�Ӥ�ެb1_�*��<�IOi'n���b�,���Z��(`��ex���e6��bD��u㝏&�	�
�@S���A��4B�0��SN[b,����	��zF�Y{/1Q��׆�����������<�R�D���K�b�o��}1L��h	@���oE(\�l�Ų5�V�34!b�آdq.O�i��SR�Mw��,x�!�q�s<���ä�NNp�/3�O'>�ҳ��U1�V�EJ)2�e$��j8�r�Ǟ^�@��5�Ѵv1sp�G�׺����}7���ܪ���4�u����	1�>V�4�s��e8��ʹ�!�u*�D�1U��6��6�m|�GHơɎ��G�%aX͍9I�j2�E�w��NQL�, �5��9�l�z���k�@���u=ߗ�^K���2d���ςh�h	92"<�������z�k�y�#�g�Q����)UL���C��UK1|YjH�"m�Ӌ����CI����T��{���l$�JZC�?~��hI�A��68�N�+C�@=|��k�ڊ�7SVk�+vZѺ�`����g�m�`bI����FCB�H�8��	X�4S~zg��RvH/ъ���� q�����${ T'[K���갉��I\��z��RG������>{K��)��frKy�A��{���!�^U�m�Tn4����R��R~h�y.��S�ECv�uæq��d��z�kִ�����0zľ�WJ�;6F���H^N~0�Ţ�&,)�2^Z�eݺ��$�b��1��53��q5��)�^�:�����}W�'��l-�4����Yᔢ��2���T�,�%}����ZUܙ������giqc�5�;U�� Ts[M��(���y��0�%5aH�n��©n�ڣ�@FT��YP�eޤ\��_��币��a��1���ō�K���;,:q��7܄����1� Qɉ����G5��U����1�d\����Vh�x<�0N��4�E�F=W���a�dJ?P���О�B�@gC�������gk�Cs,|Rz����]�Q��~�1���I�1;Ob��Y�sSR®ʄW)��,�?P9���%Ww�F��q���4k�� �l�d�B�o��������Y5͆�m�����&���U̬3�a"���t@���08�c�,�s�u���J���_�K%�-�5�\3F����Z`t]�*�'��V� (.���e�F��>*vX6�9	�+�:e�KY,܈�����p�0kv���h�+�)�=KXԾQ0���f�͜0�M���by�6�li��F�R����sc�/�c��]�$M)��g�&6�͞�FOim�U�r?;���$�<�o<'[��p�XJ�����p1�w�M:�Wt�B������^��R��dH���5������΁R$uC}�>>�h�PJ�������5�.{����8qPUoJ᪇o�cB�
��ɠ6�1�%BzϲZ�!�j������Z�,Īz��E����%�X��%�xX��V�^�U���i�k!Kߣi嬲p$�@�Gj	>�ҪSn��41BaiN�J;����W(J�|��[�R䟹:L��qn��Q��_{����B1|���kr�D���FT&M�U��>���	�J;��������8�Exs/{V�Ұ����~���	�WmϬT̃Q�L�js�����=���%�!��#%ĉ�`��d��Nޏ�)�|a��Uh Ӡ�}�?!]?��s�Y�h:�a��X�á<=<ɀ_��ȶ���b1��4Ŗ��·��}�<>8A����=���§��
�b����2�'��g��w&��*��s�@��.�Ҵ�8���P��Q~oSVo=�ߞL��h�� 	a����$+����e_@Z.���*�#�}fM^��m��r�+Ġ�f�0���,M���`:��W�C{ETe������!?<j�$8�����j�R-m�jg�T��Rs���C��9��[1��X]#i�:�����ۊqF3������mD���״��z�x���ׂ��,a���d-�g��j"@����"齚T䐔�6��|h�Q��FO/Č��R��y)��l��҃9͠��4�#�1`r^o�*���Y��{��.�;�j���j����Щ���L%����jnp	�)�v��1�P�K��y�.ë�]M�C��$��Ӥ᥮��Y>Q��ܖ7_���7)
������(k{�+B�0���I�����f:Z�#'"��M����9�(�i���n� B���J�ߍ���Z�o���M�6dP^���GA�a�h�c�q2E(-��bSa^��yz,�s��x�C�FO�ه��*T{T1�&ɯ�GzWKNmV�µ}P��є�1�l�9O�a�ч�M������o�ä���Q%�mhDGr�"\�V�G�z	A��Z>��Q]A9�a�Z$Yv��}5���xTc	[��V��������I�����D�P�1�����dSxV�zc|���Qc���ۚ{F`�5i�2���m4^H��w��C�l�����,��`���SU�c�tX��L����K��-�3a�j�+ 5�#�MOĐZ)�"�����hkEZ�X?��4�H�2J>��jҪ� ��d�*= ���^n�|�4�E����
8`�וЊ�g��o���E��U
y�pް���������óR�o�9�ժ������	����X�m�^eFu"�3\�+�MQ���`�T�f��q�t��G+�<״�)���3d�L$�ʖ+��So��nH�=/�Q~�Y~f�T:7�«�Q]̨�PĦ*>j�Լ���{� �Z�G���!-~�����(�s�� ��J�I�ʤ���]';(����� 	.SWp��Swj��ah��}���˾��^Η�x<h��~ߨbD}JB��E��Z���
������,�s��I��}\�l��/�'�zY����B��*Ǉ�X��-75.bH�>��4"wJ%~m扎fL�P?�Ʈ�;�T�]�O��@��
I��6nY�\��.1�ܓ���N���X��Z������õ�߬�vh��Z��71��eσ���p��D����R����[x,I�M�OK�!i���rLi�����F��MǶ��!�1Yl]g�(�K�]���]QL��4�i�=��v���ֵ���8J:��`9֨x��Zh ��W���n���C��}�њ���E�2ȑ����B��5��m럛{��mt� .�qp�V�\�EJ�0�1��8P��0Ŕ2�hb�x=��*�Do�*��#��ʦ�.��Dn�8�j*A�탏��`*G�&z�.��ƞ0��x��S�q�k6������z����_z��'�Nţ?$�g�eMH}1Ly2>�������Y��R3@jd��sk��P���`)���H)� �E��^K2�&�i��a���-�\�	����W-�[�ӝGZj2zz}���A�j����!<Yō)��u���[�7Z�lpΫ�d	�#�!�Ca�������xh�M��h[���*�`��,�m+��T�Jb�����W+J�Aov5Lu��|Uᝫ�d�;�Fd�8��E��{�G`�U��mm�a��hQ,0�0M��U��]J��ɭ>��	5���դ_D���ZG�A#����m�A�|˝�Vh��
i�bP�(�.������$;�^j��5B����l�X��3�#�ƖR_��/PQZ��{�fq_�|��RE�'7.��5���ڎ`QS!�:��eČ�J�M�vM�g�y"�����Ed��d�U�M�]` K�Hk�1zM��CL`��G�A$��P�V%Q��?�� F3{W�����C�������og(��@=�����o�trB6(Kt.ʰ���q���Fq�Az�|�I%�����A	�7+d�X==�׵�Kf]��V;�j4��ã��o)aFn&�T-B3z~��)�����L�D�7�B��uH������e�Y�f�S�Ha��ǋ;��`���t(�"�e�aX�{��.�O�˥W�N�$�NQ@T����'S�>����ċ�n��k1Q1�=��^��˫�$�{,��aAHE��M=�q0�~�8UNL�@@B�KD�U�j5Hn�+Z��|�Y�i`��)lm�Z��76���k�/�I�릘���-�,	����]�{�P��Q;#��Ⱦ�;��}D�uxrb-3̓QI�u�
�n��/���m�����U+	����-�C�r�ʪ�8w$��ʖ��CͶB��֛~�̙/��˙�ua�U,M6��!���=N֔��������E*�{(���j:�x=���C�`6�&X��}��Cpk���4,������2�̧����d�Z��j���>;�F<�z��:��3NcC��� c�1��n9�Re��-B5&oj���W�!��٫*��Y����rP�������(J�/��^���T�Ζ.l��UPG	�WH�]�`�P
�kMX���W�����A��i�dh$ýG;FT�Pr���_e�һw�c̱���J�,5��d5 ��)�m	5�/��f����d�1y�7i��R�}��t��<jK�:���v�＠����������g��Hݰ�P��m��#UO�RO��(��_~�E�`I&x;#3���>X��b��7��~E�#��iXoj�2�~BC�D�"N)���EPG3.'+1���ż@�_�񽸆��U�J=�f˛�r�?|�(τ����G��â��F%U�e,\z�� 5f��v�4�1�%���jI#�P�s.B�P|J,zR��p3"��j
��O�<u�7O���xh[�t1�l�j"Em���W珸�����(p(it�W��K��+ŏ� 7m�
����%ONf�5�5���Ƃ�Z��ؼ����*�h��֎E�W�O�1�5���˯��"����� ��Jj�B�N�n@3k�g[�ë4b�H�C�j��r�����T�lT��\j�KP�&0q��_u�Ϯ���.�M��_�����עB�B=]�CU���l-�ci��I�����PoC��x"�z�5��T�Z�i�C�{n&�A�<"n�5�xH}��4���e7��e��zz��C�a�ELFq����uY�ۉ�Y�?�	�	]Mv��b'�Bƙ�Mj�4�;����?���m�n7��A�1�⡱�k����?2.q���zޫ�?��5)b�����s�O��ū����k�4�j�DO�h;�� �m&j7o⼱�p(ݸ`��b�-��H�YKo@���iZgH���U֣����e�L���-�m�V���K�1�w�v�41��ű#�a��o��!�s�9R�X���⼳��f�<3�Rμ�����u+���b�u_Gg��wV��yI�+`���u-֮=x�wb$��A�ĳ��f����
[�H�Dg�lڪ��՝�:0N��+X�P/&Ծ���uއ�!��������=�k�	S��|b��H�d���F�� m5�|Q��t�MC�,��T��������y����PA��B��׉�'ʖ���$$&��K5�JR~!ћgT�঺k:(�P�U��kׯ���1�*��qCZԸ�l�{�ꘁ�ߛ�����i�	���`\ԓi�Z�DTJQ�9���we�ٰ9��XIi�n�������7&�b�x�n�量Wċ�%RZJ�ϞT�O6#<�!U�S��5Jq�]^�6N��Q7T��<5����H�\I_,>i�P�.��R�R�V�xEZz
���v��X��?X��� b]<r`8�D��U�RA�u&�R�H��4�����״�i��'x�b��rh��]�z���7�a�w�\2�t"�fr���ږ��"y���Q;[9�t�R���'0TD|��x��t;S��l�0Po�@��Kf�pR�����W۲]NY5��A}��@l�^m)�J�X�]�n1C����v�Ӗ�I"^�J�Z��0��:)ߛi6%�qd#��y�P��\�0�8�U3�����س��0/�ْ�S�Q�FLi�Zc�v����W�4N��'�Ji�UZX_�5hYQ�0l�r��R�B�h�Ӕǹ!�Ny��oL��+�(��<!7�C��/�	G(����o�T/��3
�k�j�f���ސQ����3���?����sd�D2*�Rt"Z����`P�.�E(b5a����.�DSA:ʾ:kc+]m߽+�?|c*F�4m�>�N3�L:�fHI园clW���Vg�LIht*L�߫���sZ�]w��BJy ��'�f=�7<H��3Ƶ4pQ��`�T�����Ū��!0W���ئJRl�����já�!�����K��6�w��/m�͋��m�L��n��J�� @TJ��Ҷi���e4�W��*@�,x�Ha&W�Υ{��u���;h5�%N�24�B������OdD=2���������V�x6Q��Neo�l'�����0����4�[(��,F�!��;	�᭛�|v/O0Kc#CI����Ѩe܌ղ��������Ca�h3e��24VS��N�[�U�a�����?Z��}���˦-���=�9�z�Q:�����
[鑆!%��@#��)���L�ө�H=�X7,�Dx���b�n��+�e��~�_5�%dt� �=��ì0�(�'�w��"iz��\�b��y����=ca:E��p(��I����Q����}��_���?�mn�G�lи���Y1y�H3˅�3�o=R�rwƱ�Y̷���j��[k�j�M�(~8h;_����)Q�n��ꕃ��.����7��oK��q�i+Qן'�Plc�h+GA�U+C�ڿ�^LjP?�O�]�ͫPzEm5`��.�$���/]�2���Φ)<ق͘��1��H\X`L'�c=��3�C�zrK;t�B{b6=Ofz��C��%K�p3p�`A������emH)�C�D�( 	�����"�y�����I��[iu2�;�E��|Eb4�u�M?fZ�H)I^���wQ?���F�;1��2��<T�d���G�`&������*�r�ar*��������L�_=�4���KU2W��H��Ƃ�K�c3,Q�$0��Z�%��Y�)H<Ѧ�.��j1E�ϫy�����Y���.�'�۪� D��S*�j�'�H�`�OD �:\7�)�(2�W%��-�a�o��S���;g2M�{����eN����!�P�H�D=��GԳ�V�0���4�70�U���`#~�Ŭ���48n��w�%�&�&�$f����j��l��Q3�}%�bGʨnbop�DK�p��A	���;����xM4��|�����J�]ʇ��G�Y� �01�5�[�ɐ�xR��h:�u��X�K:8R�,�/[5����g���]��������F�����z|\����C��b�q�RHzу�����d�Ӑ���d�zJ�U�����|0��M6���-���MQ*�V����ĈN���j��Ѝ��HkQQ�}�q<���10w�/���S"|n% ��j�u��� T��O9 *��͕�T�I��(�Ŋ ���G7XjH�I��X6܊
aa��!�3K�^(��^��XiL��i��>���ʵ0L�t��w�T�a�R���	�h���n";)�^�{TS7�m�ʹ��,e��O���mi��Z#�����aU�~����b�OM��O�{5&z����1LL����LQ^y��T=H�����H�4f[����%��f �Ι7���\B�S,����hl�SP���q�Έ�� ��Ma��=�Ź��?�&[l00X�~�c!�Em1�+X��'o%p�U��-VP0����9��@D��R�o�-]�ܯ�������Ÿx���o_=���+�$�k�*,��ãy��x�b�Ce(c]/��+B��M�J����J�l���:�)ITU��b��d���YՐ���y�h�E����8m"ƣ�CE���u]��8���K��[g�L֌�&\�I#��j�1~�6��t'��m�a��p>ԛ=�sT���#\�x�r�*��������ٰh=��/_�����"M��B6�ꑑBOG�WXV�]�u�|U1��A�(�u�
��z�/4q�}<���*3�GG�|K)�B��Z;�V3�az���dh�mf�2�?0���#�i���@�i�Z�&�Cy��zɖy���^�����#I�"r8J����c�Ci :q���Mc2��������n`��eRY��}�e;&zT��-����v���o틭�e�a˂ـk�w6I/��W�u�QO�p������ӏ��p_�[K/W�̮W�~�=�x���E��I����B�&b��X���J�sex�fՏ�b���D�';�4��}8����`�~�7�Ҁ4٢��,�2�JTiZ>���P1T)�02t�p�e5��(��K�Ř7fH�}Q#�r[4s�6�øfN�qk\��b��XPN��tVo����سH��B1�! �|,�ǫ�#��������gŅ:	�U�'�����������>ȸ����A�k�b�X/�~����͏z��umy-���݌V�㠐���Z�o�*N���x�}�o�Zܠ�/��"�-S��%�w��V��Lո�z��(40M�$�`��;~z)o�����gZx�t���ܪ�ʗf��U�4L���
3>h#|���5�nlc�D���XX���'��|2��<����#�I��<3����JC��yf�6%�ofH��z�cKb����p��h54$�y�sY�[�k�n�6�c��4�t�����?��O���?H�
�X	����U��?��,�=_J��84��9�)��'ث�tٍ�Y�M�Z=�H�RjFxoH�_��ؐ�o�-��e�s����$R��7�W��Z�x����Д|�&Ja��xJ��Q<m�B��M���#0��M���i��W�*FN�4�Uc:�uVN/Hv�i��s$)�������ہ�CL��,�"��jQ���{�����}D)H��*��?�]��~�8��Y�&M����&~Fet|ch���{ߑ3��������vs�OKy?��;��]8�6Z�7���"QC�kReP�D,�&2��"��][Z����3��]oC{���u`H���~�v�{0�՟�_��7������K)ZY�u7��O�5��;��<5,B�r���<˖ԙj5ڍ�
�4Ƥz8~��l�z��ܚ��J,Qf�Đf�up��w��LcK�F�������:3_����M��\��c,���ϖ�G�$�&i!�A ��x�e�="�<T��E�����CT���ry8���I�v4���ߜW�Yr�LpW�U��U*����YaƚvQBGc�����-�I{����.�G�жf	Γxc,)h�X�J�MM�Rr���I˜��L��b�Đ��ek�\��a؂{ �����'�#��
��g���}(�?~�q���_d��o׫g�5IP�NF�:C�[��v�Ƅvb��~�U�ᒯ">����|�$��YD�:����s"X�Z���Š �a�4�?)T3֭��!hs�=����h]"z��zt��Y&�%2�3Yk�at[�����m��LhoL;�Z��l�w����xs;�>v�ZW	�섣�Q�H؈0E�
�bj��&�x2	ɸ�Vb�^��S�!��ʷ����+�$r?�S/A[n��b�A��&
{P�$�b�� ����7��8��"!��@<Si����x�2�3H+6�EJ7a@�U9Fwt���vՒz�=��'��J1%���k�<�CK<�jٿK*�d�J2�碛�4�&�{tC��0uS2�0^��h"CiH*\qxÀ	���)�r�5L=̲xf^�2�|Ґ�#n�#�<�e,�a�<cO*Y���ma.�J<�B���)�g�PH(��tM�K��֦��"\&�ޤ'&a�C�����Yg�~�۹��aӹ&^�u�L�T=lD{�)��(颂4샦̍�Seu��}?P�
�1}=�,{o�e��9'ՄEߤH�Jc����8�8�Eh��}��ù	�h�j�7�	'��7�����"�B5 ߪ��h����EB�}�D1�d.WK<�K��{V���s�v���h�<��"d��� n�V�(�I�ϥ���3�LR3jƕޝ'�������]~Ag;e�Ԓʁ�贿~��_m1|o������B5��}�o<G�X���UU�����_��p�G�Q��τR��x��|�w�r�'{O�<�(�T�d���_��Z�IgR#r�y�&-�� ���u�M���0H��oQ��D;������8,R|s
�N���Ԡ�
�����FՋ:���M ��a��Ć���K!�f^���Y�2��Y��t�b�`l�����b����R��ݑ$G��� 򪬃����?0�����/;�&����k]TD�<2��o�De&��������;R�.d�\����z��������])�'��E���k�]{I��[Ș�=A���a��o��lr�ܔ��J#f�U���9\�����h~}�O����.#��J���W��
��aѮ��^����
�.�އ�����Yi�S�yJ�H�D�5;�3��	����v*�fbs���,=�FY�����h`Y�'�L �v���X�I�R ���43��*���^f�K�5���SF�4י8{w ���l~����vL��
��k�h	��c5��rMR�Zn���7�9��pL_TfK٭���Р�����n�Ĳ����n]*],�0dI�ȼj#������Z����-�����	+��--�K��4�\|�i`�i O[������eC�h�A�Cp�9�e��@ry�i.WΤ_,��'�&#�I�Jgr��Yκ�C4*�-�\|#�ȝ�O��l-?W�{�B����?X-=F�2ܕ�C�� ��?��z�ʻw?m�����)���0�!�̃�"�<���<�pZ'�h��^�����k����z �@?����a��t�Wдޣ� )�m�CLzx�����v�����N��ѵ���+~�C��u�@Js�SIO�E��0���C���L�ӯՇ�>����?�H3#m��A���lf���	D�y��A7�,�N�;3��%L�޹؛�a7�F��Q�,��i��l����=6�4��t�w8���nU�����֯��
�7�*��-1�h�!�Z�]D�vF���=���c�Oκ.wV_�����s>�'u/������eGsjd7�D?}�F �G)�}_�e����<���}aw����o�����?�}���mz����t*�MU1�>�枲Y���7o#@������Fm(Ϩ:��1}�z��t&�r��N:7S��v�4�p��L���sr�un�X��NP۟�p}�_ca���D���s� �O尖��c̓#�����$��X��9<���u�-�"0`M�_.�_���;��H##�5��A�zӴܿ���df����wp��kՐH'�Ӽ��t���8^sO��nt8�eL��͛&p��9�6����0��R���%��VQ��,ý�X�V_`����Á�o��a��w�޸�6�}���?����wi�.#�۱4�T���:pߒrR���.$~�©��¼�;Gj��1����8�MK.����ƦkY��+K�l�i�%��Ve�f<���BXJ�_�,q�M$�mf����}�O�-�z�X�\�b�h�,`?.�nĢ�먛]�oA�������7e��tX��zՄ��|����LK�7�&�߂h��Mf����;�zh�=�Ad���
%J�q�>�fR�M�ދ�1694�:]����+��'�Ӑ9T
{+�,7����Q� v�k�de���=-^/���.��jRIOn{;>�"|�/����ً?|�#�,+$�+Ma�KT�� ������#X���m�`x�Df%.݊U�����1ف�.���6�������6�ɱ�8h�����3����J��=.��Yi91���\�l��������k��c9��^�D��+�c4���B'��=�q�+[��͝��?�;�ӟ���3R;t��������S��D���yU�t��+���O��JA��6T��vA/8�ۦ�ʌ �bEAT��H3gP��v'��\ѣ$��kn|�NK��5�M
J�-H�l,*e��UW�a'6؎C�l�n���Ȱ��	(I��U3�([��	���>��p��G�1ɑ��8��X�bbD�m˦�o����ّ�|�t�������*�l����?�/;�J#��GI�	J�#�\�;�J�^<l� 69����n�#�0�M+��j._.��l0J�LmY��^�J����<�A���4Z5��8֣6 �^���qb��~�\gsE�t�7�@H���Η��(q����|\�qbEC(��c*�A�����{��U���>'�b�9�ơ�uM��xj�uXĢ����π��
 �A�O�[X�ကi�~/88��2�n��7ǉQ�4�G�(��y0T���.����R%��,R��K���g���?X;��]+���s��av�d�yR������e?/����Ha�$�@�׃P?�ܛ�N�Y�c
"6�r����<yl?p�_tۍ�@�-X|:�l��D�ؘv,^!��m4��x"�)26֘;ŵ�yD��4�fQxfe��&�n{G2o��F!���ow���$<��&1.����R�[���K��_�'V�Y�5��^
��,�b̌L���V���A_g��2��H��ImsR�=8�:��q![���-�?C�S�ݭ�]F���|?��dmv�ﷆG�,�\8J�AZ� �Z�E�Lo,B-�1�����Q�2k�8��cs˻��E���������+�O����e��P�������W��O�JR���ӻ�}�>��c�S;׼��Xm��ٳK��W�伕~�n��5̮���H��-�`^2��p�[�g�a�'��i 3��8�\v2W�~��Hϲ�:��$�����o����˟�L�'����x��yIB0i?%O�t\)%���p�����Yj�H��wYe�u�Ԯ.�>S��ߟN�]�Aw]Z���ԍ�&�*45�֤}�>Q�e�b���
S�j-���^�vS�(/ڌSIHV�;���V�J50nM<��Ԁ���)~�Y�����b���"�y���M�=
�)��CF^%,�ospa��P���YY�,��9��u�Ԭ9<�4NP=)�CH���dH��5��cA�8�������B���ɓ���u�>h��咢�s(��p̂����Q�����C��dh4O;6��QϮ$lJ>�d_�9�W���m�a��O�,�Q/��,���C�����؅*� �榉�ƗKޗ�	��Xc|����ᢱ������|�K�x'�1l�y��I-�c�Y�D���v���M�GZg���X򍱑��TF�VJ���1�fV�,+1�og���y�9h�NT~4���F]���öR^��|9{��I�l�La��ŀ����`��Qj@M�ۀMs���gd�m�צ7��^��- 6t�����.��1tWr(��ţS�,tQIn�4�mи���eyǒ,�FY�R�*�g�rO�nHq����4�<����C��Y�E��%�� ӣ��jd��o�d��H������vc��и�s�!x�7���3a3>|�(K,�ƵZ�DUrf��������qH��Y�ڨ`��5� ��a���� �@����UT����ǿ#8˶	22�:�H�r����BM��l�с�\3���h�g�#`����Vt�����&n�-	�f��S��-3]E"^`}�����������P<1��i�
jU�Ċ�]j3�<v'lv���z����V��w�w�����X���B'I�;���Mf$��, ����XG����{7$F�b�@� �v
����yz.;m��lLU_�!7��>h���[k���K��O\8�C%us~�U�/;����!��42�X`[G�[��\� ���ʚ� �va&����uޑ���#�h�n_��h�d���]9��j�9�e�8�l���A����z���y��3�M�O!�|H:�ihd����an�x���
�\CS�d�J#���Aԥ�Bgs Tm�z�wwz�]�_�𻠰_g�T�/�w��Z}�wQN_4;���p5�����\gɡ9yt��#<:��$�t`�[�̾D�������T�3��볭�����S"��zX\7�/#q}�n���xnc��G�]9ዯ1GfJB`���%u|�~�=a�j��{�VS�:�{�ZhZQ�����y����z��޿���WC�T�v�o?������Q ���Q��ZjF�uҡ�F�7eC���n<�/z���u���/�9�O9�{�E� ��<NQ����1$������q�7/��Qb�ӑ�� ��^�͓�Hrwu(^ˋ������Y� x���:��w4�62��p�&]7n�k�� <:�u*��v��L��|?��W)T2#�f�vE��B,�����H�������sl|�ldg
R��H��E��$v&��u��wx#}-[56� �;�����Q�4�84��
)9�����޲[Cn�N�\�'�JX��&�����c�u�.)V�!PVeշĽ�!�D�%��������Z�#X`�Ә��j��ُ�Hec9/��3#�5]�����=����q�W�mG-��:�z��f<�Y��O��h�:�T�]D	����`\������s|H�kf�*���iS���Ã�b���\�� G���k�k���'���v��q Uv��
�u�m���p��id������X4��$��bI��dwo�^��}Hn`(l4v���э�m^�x���4^��F)z�k��O�c �'��~��X)��<w���1��[I�4�g��MPe���*\�D`�F���ޤv�7}�mY�+�%s���s9Ks	퉤��ՙ�7d/UZN���ɴ���.���~��.�Yu��,g+��-c�������(��|怽��{�6I�x��'K	{Y�͑��w��$�x�&qI�Dru�sҽGA����Q^O4|�qͣ>��y�f#k80c��A�ް�����;MX�HW�A	��{��	��ʽ8*K�fƃ�2p]p���ߓpC|Y��C� ��~�ܿ!)O�dB��i���۽��1ꮦ�l5ǸՁ�k^�8�����u�
n�`�c~:9K#h����>�
x(���$�����ת���71]�뗌�8���Ĭj����:Q[�j�Դ�1*}�{qu -��]֠/Y��r�((ݢ;�r��mGpR���ݛN���7^�Y�O��Ҭ�xΓU
���M��d��1��:�榅fy�W�F����!0yJ�
�i\����3�ΜG�=ǴeL̘�#}�ad)s6\<���G��+�d3��%�����A�����qy�@jQ#�s���\��Ȅ���QM\c]<k*& 
�ă����c�k��&e�*�W�L��u>�����q��t�%6e`��F��.=����)�!y��)�2P���+�4Kus=K���� y�e�r~i�P�y�C޶�_댡^J��� ��-Mmnb#�p��8�!��Z���쮲hFׁ���� �G�H;~��Ǹ'��8�6��yu4��Q~�����"]�b�V��dU����r��@��^n"�Gm[�@���������o�jV�D{��]eJ�[�1�{h$c��c�K��ݹu]����������=�X�-5�\jc��GQ��%qFf���]��s�Pο�J���Mcr���V���	*�,2�ZC%# �T[�9�9Q*� �?D�B���扇��;�&@Ykd���X�5p]�M�1D�جS�[�`��(�,\f�Ɨ�|?��H*-�bT����%1���K����|��5ARp�y7�r��A����<i���d�uh�����w-ŗ���(�i˵���p�e>#� M��>[QW�����y{<�(a,k��>|L���� ��-�!�%�c�8z��7ԦE���}Yc�ꑎB�R�%r���x�j�Yc{Q���T���Y�-�Ӝ)��,��p���@�*�Q޵�=6Ia�R����D
����Ʉ2ҁv�P�q]�L(ͣ�)$��k�6ÿ��k���(���}	ap�ĵ�z�Z���)��4ơZ��g��,�V<.<���1+��g�"�-�Yֵ22<���.d'���zt6���7%�:'����c�u�mv�9��F��)^��2k^��k�"�]��U�]I�~��4�rJ/�DZ�&�~¼��N0э(T���w�(_\�A�����CH`j��p�k�3G�?�s\Lb�7=��8�pL�����]�yɃ���r�:�����:y�qZf�z�ӴW�!�Z:����ǇtU��ꖙ��������������+�<�Y�����^)s<���gP1e����Sor������j�Y���þ�yc��M�B4H��%̢����17cwf��Fs�V�2�;e8��"�r
B�|
�%+��X� �iv������XP���APP�9"�{��^���$fI\5���T9�p������^��%��pf�x��UR��$�׫�7�2QȊ��N�dӯ*�*˦b�����jg��A>����Ϊ����1H�SA�\{C�?>�c�^�o�A{7���l���x��q�@��ْ.���JS�7d����J��1���]&4u���,��C<?�҉�y�"=+����Ę斲KI����FW�������Vje���7;��2��i��Il*qH�-ʱ$��s�-5_�躯��/nN|�^ԧl����L�z��?�9Wd c�f.�����m�r775�Z���4p�[�Q~]���Q2���
,�&ۦ�LR�0�&Ӄ�8lط���� ���,�v�����A��K���Y�ڵ�����Y��J���Nv}f��J�x�~/���U�����f�w H�h��oqRO��Sr��v�^�8�j��s '�@�5I;{|�/0X x��m)Rh�!�o���V��p�5]��ƹ9�HǒJY\>>(����@��b���g����X�]�N�'����zph�XGa���9��Z	��G���)iejܪ�h���q<�lyX<�r��ˎ�w�������vXկ�:afw�R �}�F��ZLJl�?f����)��~z�����Ac��+��1
l�[/�-�:��ܲd�S_���_��C���MY/&CV��<e�!i��F�M�^v{K�9lřV�&�@Ja!ꡇ��䑣��?����0��6�G��-;��{���A�� �%]�{���Y�kLIy��WƟ�	��9X�=�ˬn9�Y��ṏ��p�!�Ixnϝ�@��S����T�gC#ș�(�Y�~u}�QJ�Gl��e���ln���I���q�`�\�cN4��P��U����`��ZCe�k2M�]�G�>i�|h��i����T�Y�3��ʸ!	��YG X�D��,Wj&@�����3#�
�b@rcmNH(�z��0R��N�jVM�6U�G/E|�|�x���J���1�ov���i�v0#�kNӍމ�~`�����=F ���訆r��}�Tj�>#���CǾ�~ٽN��Q�]F��?�\�e $w]���d�D[v��{��T,֯_w�As��	[���{:�Ed{>`1�zy�llf�m��ʛ�JZ�J����M �N��:fyu��Bg��7�Z഻S��#�H�Df���c���3��c�}
΢�q>���':��S�Q�����ѣ�C�;�R{�F#`���j�q�Aσ	�y��`��.+�����<�8����<=>3�GС�7X8F~f3�f�3����Aoc�<;�Z��Y��W��#g~������?�5W���r�pů߾8��#a <�_�(	h��H�JS+�fY>�=u���'����8̿�:�7A��,�B�ǫ�I����UFQNc2���]���7�F�dҎH?��ⲗ����{�����0�%���	� 6J��Uc�����V[��x�rI�i�|��ȭ�S�f���FV�j�c�z�\�����i2�'КA�.�5�tjxC��_�%~
5��=!�Aՙot&������t��7c�y�{yΎ/�`V֓��GNK�Ů��-G�4��0nX]���Ħ�x=��O�IKd���{�y��UT�)L�nA9�f��J���%ɸ��qV⛙�,��.5E�|�1��.60K�.�X���s����-��j�9��dHe�dv�tO,M��	��D�������%���������uh�{P�����G�w̆�x���\�K�ן����w�ބ֚�60�`�(�Aխt��k��W��=�3��$��i�՟�����,k0�I�V�͝̊�X�}�2�Q,�UA����\�Fj>����k�� >��7�b��I�Y[��4��׊��}<D��T�%� �pu���D?�T>}�\>~�P�����?��X�v��g0M�Ti�Q����;��׈A��Y����Ȳ�,�ԞʾZ��F���ɘv�i3��lD����0�f��4&JϏK\˻8�����R6^�dk���qk_'�yh�!��B)�w�����O����1p�HEc|Ee��D���y�ωmƂ$
R�� 8��.���l��[T�$-�����o�\Č�:`�XT�.nGy�[�zJ���۫r#��2X��ܟ_U1c�31z��ˎ������]�&�zDݰ��b�m�O.M�Fa��"����i��J�O�4<��rh"�"�	��0�wJ�y��|��	'||a�e�e�_1����{�d�>5t�z~�[\���XcM�����ndi�Pw�fh�M��v���F6� �%��׉�Q��A�C(C1�V_m��qp��p��,A-6��]����cTfݧF��5�i��K�=_>2D���'����UڧO�@�Gdc�w/5��a@�o�0=��R�����f�>8����k��0��ب���Rn,%�l�����{	�Z;�h�]ǔuM�J���>=@��Z��UJ�U���%Fp+G�7�$���!�Sgb9����f��;V��yޫMW�R:��(p2�LM)bXq��;zؐ1�B�9:�=UR���@zJ�!,����sy��t�Cc	�F�Jn���#�/���u��D�_s]Mբ��H������s��n����. ���H����e�^����Zɡ���*�u�!q�i��aᆘ;��޿��"V�x}�៴8����p��)��á}�h���eӇ�tz�~�`{���nZ8�pꃃ9/c�?��m��3\k����y������V��"o��Y���FUQ7>ab�S��glp7����d��)=]�56�i
Co߆%2��j�2�~� �g1E3h�w����LJ���*�0ǭrz>n��`�%����7���O�j�rKp��!��H��x��g�F�(X$E�c5o��r�d ��4��lٴ4n{���dbs<m�|U�=X����#4�)��c͡j�>���=4�z%ؿ�*G�R��������UD�/5(�%?��*�^��N�}cc���R�x��徴�t�k��l=�D�F%َ�'���A�}�.�U�N��bn����X�A]�{ʂ3ep`�� �͚x��?���n���Wh���3�q���T�~�ٻC�窇�zCX-|���pTUM��g]��d㭨�1W��p�i4W��t�7���<6����X���F��.dĞe�q��Y6A�QY4��(�X��ۉ���by�e�kC붧 q�Y~�H��u�vҦõ#�J�/M��q�)%���Ą:˫vVݴ�v�Zl��墮}��1q�h����$�uR�R��%��9�<��ڊ���E&}b�4E��2�V�:����d���0#��p�Feૂe����������ݞ�k�ɺY#��y:����$�F�U�?�ت
ɒ�=_v�>��q�(�� J��1Fk)���y3g��>��O��e�{��_x���^~?DА�3��k�A�(zI ,!�F���7�K|ă���m��L�3m��-��`�����g���dԙ�l��/�%p뚳|*�O�]f�IL;7y���&�鐴`U�`0�Ùl���������oV .:X�fǛ:��ۢ��F���,��B�����T��#� jH�.��$��ق`�h��)k�͜�F֪U>���$�ɦ����+ ����Ui�&��Ȧ�ϊ��Ƴ����[�w��s���ɲ�J��8��fɎSl�mVQ���&�ϴH�"�ŝ`_3g�{j�K���gЙ�0�s�S���R� G�nޕ�%�t��{��0G0zt)�7w�|�hg!FYt��Ӭ�LL�m�5kfY��L�s�>��[���(���R�3H�g�E�D��F�P��ɭ%�,�'1��s�J��w�
���O�YS����ÕRiJV�Mf-E��%���1��pp��������q��ܬ�~��dN�?v�@�Ct���������Z�\�}��((�2�ը�I��H�l|�b�j������Q�k���_S��� 1���׳�cW+�m;�b���aǪKm6��U7p��0iS}� 5�,׻&�u��74X����bS�f��M�(o�0��t�I���â�:�$��,�+o��_�ZL"\OAs��l�a�������Hc�ȅkML+LׇX�+������8�<�uQ���Q�"������֕���#�͐r
C��'�}��a�s�O)�>��D�A�Z4&��q9ˏb�LX��w��Y��C2|o𜸖��q��#;�,\ʽ�T�^�^�% 8���m<yj�>�s³����ޡ���.��[՘�Ds�r\���,7(ӡZZ-Fi/��.�&����y9�fW��hA����ʺm�<��~�Nw�P�����լF�4Y�����:[�1�`�Yo��P�H�s�F#h�Oi���R�{Q�����y��@�
�V*�3diW?�
q���r��*��_�,�ۿ~�Nj4MJ��d_!�e��#�(:��T;�Z�s�f�LwR�m3`_�(��u`�p���m�`���%������G�Ny,owYW_�k%�CV�I����)G"�ɰѸ]�#�BN��^Cj� ߁g��xe�M�Wt��e�'>�\�jFd�M͚��Kl~�=<A��1��M
�~#^.��[Wy�e�s�Yo���U�m4��u�5�E<��CT/�	lbb�$��K�GŠTF���/�ds��ڗ��"h�a51�$�IB&�=X�zJ��+�A�bjk�%y��N�(Ј�%��?�yS��@��{9_�E��f��q��J��U2U��� ;�A���x0��`�\�X�h�ь�d�Uto'U��]y���k��J����FT-�w���ws����:�S6)�bu��p[��g.r��҂ʅ�@��(<d����ώ]`M͟i�Y9��������t�#��o��d���ɨ��~�n_�h;f�!)4/2�m�6�Ng�@>%��A`�5<o�_�g�7j��y�p���s���F��{�a�b���\��:�p��w�c�{��M�bǼ��/�yIE�4Uyfd �\�U?���i;�*h�Mˣ���)�� ��I*d�8x�q��3������u�D�Xk������-��(:��*	ƀDg4nFEc�\ٺ�9��� F����C?РSm��[��1�-����t�5���3�z�y�p�E�-^�*�/�h�|��'��h8�*�	" y�EKZ*���]E3|S3�"ik�{ �9*>X1�fJ�t��!�1ɕs�fVt=�EŜh+,�&�^b�sd^�b6�SB�{��M��ؗ��HYU�fl�M-���:�C�������F�
��"�� I|Ɔ�B�ldб�1\���1G(���<�R�8��2�F+I����8e#4d}Lb��ٗ�ۗn>UA�Ppq&��%n�u��\́�f�GV,���E5���l�X%�>����(���>df�d�8���T�@��1�s-Vl����:�� �4���ý�%�7q�ѽ�x�(%�����y4��4/"VS�.�s��S|��>�|wX1�cP��}���<�@�~�� 43�ib�:�x/��^ơ";�S���@�d&���j���R�ɠ��	���o�<ש�y_Ƽ\�GY�r����Aّ)��4�qݪ��L�.w��E�:8��{g>D���N�pKH���_dA�y��F��9s
�C�Ǹ���דБ�A�b�tHH���]��3u�����������3��$�6}��;i�PlYgx �/�﵎{i�Ӎ�q� �Rl�G��~(�7�\���؝ɼ��{23W�xZ���r��(�Q���1'uQfp���=�,2��-~7�%|���(��\*�=+>H�
�����&�L�cf��AA����p���nFJt��k�$�f�mݸ���~~��y�n*�a°�g0xE��RM�W��t��&3���ڇG�9�k�����yx����0�7񞱠LcX�xX�ɗt�ٟ���/����m`�q�U���02����m�O[����V���v��b���H' �n6��0Lï�� �᳚^��<�}��(19DNs�p�e*=�v�������i��7ǘ$�.1a�[�k�������f>�}V߅>�J����Z #�w��_ޝS��g&(��"�Z8���<�Hi�Φ��A��`F
!BAt8�$z
3����RLWUZ�6 MY�B��3���]м֥R4;�)�vY10�*��u���*�^Ѥд�l�+�ѻ+���m���y���4��2����iL�K��r���v�i�k�>�)q�n�:�2X8�4.jL��&0W��lASX��?_&0EME��k�v�n4����d/�zeײm�}���{��������I�.��Z�B���֛�"d6VnB��Q\;u��؝��=t�-��쭸w��#�1_v������zTu�yM�Tbd	L"�Y�o�5?�qoc�Ƴ����F&)k!cL�^/�X��zt�y�.�!�Ri͌1�D�?�h�8���;�I�pG��E�{�]O�����F�3_כ��CC���Lp�֚��.)G�l���$�o3����%����	��nG'���3S79$����ł�ϭ �~��cnrf�n�x�D������E�}W���#�t�)�k��"��@Q�lY����>�����,�N����A�Ǭ�Y�Ѱ�!�I�\�7VZW5�Az������ׁ��]U�k\�)xw	g).�F.�|A莋_
�6�J��jR;��t�)wd�u t��*��ܠM|�|_\h�8��R��|j���`v�'�dhJX+=+�!E�z||�)��U��i*�P2O$��ƀ���x�� �ΐ��n���4׸K'f�O�V��NQ< *lpkoq��t"�	]޿����������̸1�����N����e��r���i�5j&޻v6F�^�P���D �R�&*I�[$��h�ވ�I�視<�S��hL����3H�`�t�e����UH�p����ƚ��� ��)�JӾ=((�B��vɹ��|������x�ǫ�����9V��*/f< ���_��c��ڊ�y
��M'�2D4J/W�4jP�o�����ڰIzȊ��*�z�z	�ε�2�Ai�k�!m�A}��Z+�?>�zxH��Y(�k���M�a!b���DdYN�0cf���������PN�k�4VD��yW�e�J�jD����>�V�	��.P������Oq����MA`��=�	�O���]��
��A��aP�V��Yɧ n6��[�$�Ts櫭]�"%}��6�ie��G|*�l*�(!cOG��:�囡[�ch�ե4��$�߼(�g�E,��8W���uG.���O��g6�r�y��v�H����x�a�`�>�z{�+�k��3_2��ŋo+�MA��b9�9���H�;��C���9��^�6�S_gqx{-�%�.����|�M�t�P2��J*����Fv�T���3VT�L���I��T;��iP�>�f��=F�Y~�]�QԤ�x����/��WKYt��mnZnТ�� ��12���%���G�����J)E�Y�x�����Ш�5��՘��x
�=��/�8��|��&�h������kI�B���l��u��Ց�.sML*8;��,�:���w[Ȏe��C���3�!� �pU6���7���m2��e�w�KֻR_��i��I53��ն��8p���<>Q�	�|4`z����^����~���&�.����A������zj�z����	�k�B��<	�<e)�����.*N�V�`�΁x���p��9z��ˆ�o�t
����!2�]��P���4��l��6"��(+G6���:��*�#��6�}w�=j����+8�6��7�N�a�2ԕ,����@=�ڝm�����q\�{=Hco�._�M��U5x���m
�Z��}��_ML�,j��A��0{(��`	ʏèk��Sn"g���pl�%�h 3�^�@U�n�ޣw�ۯ�qݲ���!��z�O�|���O��9���[�JhMz~����N���X�'㐂hĊ#b�P�a�iAc��sJ����XaVٲ;�'(��'�Gqm������W�c�
�<*	�*�4�r-��WT:���[���ل]�7pӵk��:��5Pa�:Wʟo�n�<jCJ���Y��w���jS��'6g8��X��۝ܰY�l&/@�M�j�Դ1 �1N�Ǉ�(+��q��3� 1�����:k�\צ�#��m���iH�b�L.�TiZ�sC�F^�F�RWe(�7u=K6炏��+n���b�r�.�B].sd��c3E��y�}o'p46h�G3kZ�㩜��M�R���h���>(o���#�7�]��]�^���ِ����Z��m}:1[0Ab�����sRrz��[�c�e-���X]Ib~\7��٭��#�l�3��+�L����}�qM�P�7S��l0�PXc�����C�$�c�^F�:���$W3����?�!̔m�KŽ��!,�^��� �O?+㮬�'���T�7�uK�E�Nd�&��F�`��`��������Y&E��a���TK���>�tÎ=�
ٓh�`I�Hǿ���G�X��e�Nj1	L�r�F#b<���YK2a���R�ŗ��j����.ЖRR������s�`J���FI��8���5U@|�*��@z����K�.X���0a>т%:��n���v�SQt��z�)�'��eW'��&��8�@j:�Md��h�7�W�!�D�*&��[�<='A�J"��<)D0�ri����!�LM�?O�f9��ݟV->�"��V p�(l���nРM:�2�8��)�(�#'�E��0�XB�H`JP`�����Ǚ�y;Ȟ���{��4ω㽄�t8h�� �"O~sX]2[�ڭ,���ɍlR<�&�&~�3�Šr�k{&L�C�X��JCR�G��Q�5*�q�g�Y%M���(v�!�"+�5�\.iHeF�Oݴlh��ow�^��v�)�	���(�쪷ʘ�Y��E��y�
a��J��$l�@:�3�Œ�YD+ޘPC�l�y�\��,�ܲ�j����L�*X`����������Q0�5�秤.�`�A8 "ǻ���d��J&�Gsn��'wZ�wu��x4Vſ�D-w�ɫ����X�d��ڡ��?�㓴�_��.8�<Ŵ�z�l�9;���.%|��	�X�p�H��\&�:�g��vx��<Kg�#nd��c30�R�.v�t�L�H�K�R\�1{�F�`������"���0āt�ǒ���{GFa���Ecs?�����N�����n�i�����5�'&�ݏ������5�{䝟�Y����l̊)�d	mL�g�[��}ɮ��I��
	��ri��lks`&�?c�=�������{��"��R��}�#�}��U7�A࢘�9F ���4&����q��Ш�K�FG��$����'�6xmX�Y�`��� \�U��Ɯpg�kH{1� �@O��df���`��.#���G�����l���)�M8�A���A+�)I�D�&nʌ��pcSd��;�1c�
�̷�<�N��U[����g�Y��σ�.���ϻ_�Q#�*F��q�!P�M��n؋���|��-6�iM$y�wY@���r<mswu�ƿ���� ��t:s�rMgz��ѝ{p��Kw� k,�/��]�Ez�o�]�4Xr���
\&W�m�`E��c.��N�qΠ�fU�3�q���4맙�Tq�I&�u1,*���RV��Vxy3�`�rw`�E#s��-�hj��xM%��V> ����O0I�������x-��(2"�3un?������X�bg��Z���ԃ��a��Pח 冉��Z#K�rG6�<ΜS$�Mgw&�����l��!��]�Gݟ��=�j��K�G�/*	���k�}R�l���9+6W����ӻz��O<�0N>����6��)`����Rs��.ON4�/A��ǽF��b�WC�x�N�7a�mc!{VN������Y���.3��&�9�?R-��PV��£���=|�JNZ.jd�X���bsyQc�B�fIf���/6�l��ϳ�xT}�Hޞ�rk�hT�Ø�G�G~���M4�EZ}>N
ڕ�HI%3?l|x$R�9H�[����c��4$�(sNj� +w�6d�P؜B�%����]g��E��KG\��!�3ZK�jQ>�ݭn�^�D���P��@0�"���a�"lS�8� �_oȠ^��ڲ���V����y��FD��p�=�v�0�boD����^NA|����Ƽ^nY����tL���XV=��Mì�vm�x����+�W?\���`V�C�d��;��=�	���)���7z��N��Sz�kr�G�%~����i��m�� �uű?��bd�A�oB��p���0����~vӵNq߾y�U<|�E����+d��'�N�J8Goļz㧆��su��:��/���!�oЂ@���d��L�g0g�{(��] 5���Q윭�x�ϧ�*����`�&�(���$ʒy��@���7�F�|�ǿhG 4���<A�i�Yb�?$�����-2U�S��4:e�?��sy���(�@��ж�,��i�͋H�/�m����Yɷ�R4t����e"�%4�x,��1�r"G+h�Z��.L�#u�d�R.`�<鸵�I��(��<v��Q	�)r4D�k��%Cb���Uv�y��4�~�$	�~�-�K@�ۙ���;����ئ4���-���X��B�(9ֻV/�F�Q���<�#����,��FF���)�&4���l��a���We�U�h������h�$��c��_r�ʲV?Lv�۸�X��#G�	�����RH���Yh쿆��(~+y�X�*�(r,=$HG�S_I�/و:�s(�_��v���(��?�Q�	��7p��F؛����_��_˿������?h:�����.>n��--��3(fpDG^��0(T�A\�l�[';C�YsI)������V��@V��5�Y�_��'�J��d���JT��	*x�#��`��&���������X$�m�L�9�o��]��a��Es�(�tZ��*!���es�m�:�Q��#���@�-N�����K���_4�Q��9��X�ӀL2���׽eh� ��2�Sw���R��wc��\]��+̰9KΘٹi�{1�H��,�Z�	Z�mɥC�z8��.�]hg���AgM��I����r����n���B��A��ٞ(������߷��"��K��[\�V�ʺ�ɩ�jc���p�际�D峖�f 6α�r������)��;���f! �����kq8�?��G)ccb� 95GY��5a����)�:	��s|��Ici.��:_��wJ�q�cP��o8
��e���)�xO�o�����R" 9{w80~2aL$@p���r�"�W� f*���U�l�|��޿]~z��&��@�rp~�NG]6J	�`�c�����������?/�kY���ګWo4��T|���.��{M�u+j��n6]7�R���3%��jU^h�{N�v���n��aSi_;VĳL����#m�����`��O�y��}��I�4�5H[|��MVT򃯆P��'����x#TP�����-(�2r�3g��CEo"t��B�c|úLA�Y�[5�uYY���xy��m��
%��m����|w�/��$���E��:@��b�yv6�MVa��1H�Mǎ�U'~/�+�fj#*���)D���4U�jcc��\
��˷�����@�>�u��7[�1t�ew�#MhH3�V�v]�Z��-8n�[��Z	k�F� �	9c<6�m=����2���Q�}���D'}(W0zz�)2�=�:��w^2X�<�Na�i�����D)���bqo^me���NhԬ]P��D�h��M��XS[5 ���Z�{�j;�ߗ��_c�}�C�����/�}-9�G�<<r�*:�`���F#�����ğ�IPI`�:��{6�^?N$�*:Xa���-�_~�u�}��޽����z`C7�n=F�8�z�}��A�܍ʘ����V��%��X�Ț��o�������3�- C��ʰ����⹖�MǪk���q�����2o��\+ºTity��!?J"�7S��3ZsH��f�X6Z�6L��,[�)���I�����8�K�ɲ�$&1�� 6)�v½�V��ӌ���YoY�z#e��rߝ�yT	�aR��:�í����kt ��m�73���$z>����i+޼~^���	��ϐ<�4K�����Ix �M��|t��0a����S�H1qS�$�E�Q�k�������.n��%����ڂhh�g(���yY�sЀ���}�ҟ��o������m9�K��x>���t���M�n�����)��o�x�~�2���O���K߅FԒ&�x���n�g���)�����i�\q�@���@̏������o5̖1�~����C���6������(����so����*��p7����_~�����+9���h���K�I�Y�?Qm�޻�8Q�SE������� ��K�w7P�u�@z����9/�����K�1�h��@f��*=����䙃#��8
�u0�e���W6��]׮�xݗ�s��^��@�4W@oB.��˷���{�ödVW~f��G
"N��jTA��@:O��s�UI�w����Ϙ�R��E9f5Y���^k�74�na�� ��Q.6M婉�c\o�v 	/�Aq��8#%=�-��W��^c�����[wZ�9�"���'f�[0����%��>��l$d����o�7���?M����@zN*���<�OIu�5<0]4����Ag@-2�-9mAb}�C�95�-k��sl�w�^��#!�V�@��?���!����S�}���Oa�Z�~p3<�>p��],��n�׺vKl��rbd�v(-���K|�N�3����[@yS~���(���z��t���v�##}�@ڔ7���m�����QB����wRf�6�����˿�e��������ӑ�>�sd�ӈ��E����c4N~���@e�n���ˉ͋5�i����ś���U�QU��իf��z�chLt�c+!��脪�
��/�v[�NCT%?m�_������#�iD��X �Ϙ~K_<���m��/��P�{:p���<�Ên3p�E=�C EF�eF�@ʾcW��D`	*�N�6*z~X������V���۶6����a�x� �@JX��?�N&u�Yaܶ����Sf�L`���ç�ш�d�a�:��"��~�i[�2n�����f��k�hI�����fP�����(4S.���/����I��^k￫8,���H۽)'�&J�Kz����
�]��6z�=G����l47&�RvdV�]�.O!)tgm���X��JL��s~y.��~���"�SL_T��w�۫�C.�Z����ھ�7����5�[�C�Agz���|�z�r3H����Q<�,ż�F�&�O��!�y�1�<ؤ����Jk���<�S"��̠���m�j�U�bNz-�Zl�]iM.,��wB�8d�(	�>����o�y�=�c�������i�D0LQ�c����:^�����m��0m��8K� Z͛�~��9>½X�IЉ�z�d��a�ulb��N�3�)�	^W:i������W)�N����iZ��֑+��\hd���(�(F�fqǊ5�?gf��γ�IC��NF�0C����X1-���|�"8d?$�=�������}`c�Kiuhp�1f�0{;�NW����=.j�R�.]�Ĉ���&����k�t�5��K�+E��h���N,��Mpu⋳���a���6��?呺�'��h��߲��aG����N��ݰS���Y�96�^�VG|H=U��W	gopT�3�\�J'����*Wp]��,M��Ը�3��3���Wuc	|��9�	W����󘔞1�5��A��g�������`?��l�R�j���k�ej՗գF�� �f��[w����݃�$��P����2g�u����ܵ�)�}ג��nWg5M��Ϡ�l�����B�`�ؤ�)U��f��LFDP\N�����p�o5n���ǪVy�������=m�]�I3�<����ء�R�M��t����W?~���r��P�u�K���p:_�a��f��]���[�"��M13M��9d��T�gL�0�gC��T����?g�flz5"�7
�	ԩ������U�,���>_���n<U�xG�"�z���jJ�FT[�hc�j��R�����Fd�K5����ņd
9�6TI�7-ſQ)�;"����?�'<7��9�{��B���Wq�$�	A�)R���J)��m�K�Q�������j�$��kUI�]͔Guɉ��_lQ� �#�>��L�"TA��bnN�
*iT�.����!�|I��&5����@���� �'�~_���Y�j��ēNH�̣d� F0>`�A=z�i��Jk42�8����ˋ#F�>xTӐc���YV9\�+����o��Y\=CIn�x �C����������h^<2���_�G1�<k%�Ǟ�L��!>�u����|��AR�>+�p��5��ף"���4�e��L��e�ւ[uc���|Lk �x�ׯ_���\�B�ɖ�TΩ��u7���\�M��8���M���������H���ש%+@�Y}x8��l|�p���z�d�����dFO��]\���)5b��Rtq�B��U��b�'�i�
�C����	�h@v��{o�gN0(rs6�=�9{�&3��1Z17�v'��.͈�0������^�s%�{�{V'��>�4s���i����$��r����V��^�]�K`�R[�U
s����<+p��qy��F�|�5�����Z�0E��A���x~��i��l90�:�I� 3��&<|��]3���C/$4����<_scǂ��}���3m:��f�_�>w0�AOI�3o
	%p�i�]��bYY����a�L󒙳-аI���=E����C��ô��e�q�����)��_^�1���M{N7����ks��M#Jl��2����qP�M���\!�<.�|<f�ya���CH��jf����}hB����a�A�����L=�G�꾶���TZ�B�1��"��A��n|F�9S�O@��a�ϵIr�黔sN�C������[a��6�p��Dubl�'�2��ӶN��D"����}!�-%ǌDU5Oym��A��J���X���*٩�3�i4�3�CS}ƚ�����^����t�u��f����ˬ��9��n\
1{\4��/4�F��M�����pS��5�0�Ʃ�3����j(U:gEĢLҋnU�A��1���{�pƆBV�VC`��"�����B'�++��Ў�C��?~������pfj��n�,7�M�<hXN�ѝ=D���51���׃Q%6��m�?>�Դiw���n(��u��g�����z8� ��FD�����^�;��,F;�T�� LàU�5�(��-��r8B��^�9\�il��|�v�@i��5��7^��P���2������9�~v������m�|��8��2X=�ʞ��P��euPxtr4à�[�޸t�Z�Z�qEײ6�o�.�q`b�c4W�T���½9��U��w�fmR?<�X���#_�F[�wm��i�ML����ГCj��dw�-9�P��19����YZZk΋���<��H��Y�;������6�E���m��b��Ҿ�d��ǚ�i�;6��6t��	\����$�e��3�N�4Q^�β���୪w�q%�Pq�.E�3�̼Ff��j��]��K4^�m�Çn[��.H����Q���Y��^wY�:���(������<�!���j�ǅ�/������k�^8�?sb0A� 'Й-�{��)�.�y�E�)u�n������8=���~vL�P@"�,����%,���I�A6x��iH����v�0���E�,~F ݂l���1 Yed�G��)Ue���<�{�`�v4!o���n��!��i�Z��s��:ˣ9x:��Y��X����6 ��J�ƃ�uRd�}'��ܙqxZ���8�T����w$����L���Ȝ!�	�z)bdظ��3TJ�K}�U�	P���mò�Nd���ύ��l��zl�-@������a-G#�H��� ֔�Mc��ʘI/3c>��63�Y�	�n麄
�edc����-���;)��'���>#����=BZ���k�J�c��,���H/��:�#s�r�vl#�@�N:͈�4β�C��5q:R*_42`��vZ�{�B�f,H��8���N�A��ҵGJ�^��0�8IA AY^Y�������E�����lP>�����^,�&��ʝ��wHi��Y����s�!��t��%���O����`��#K�x��l?)"�����ebm8��V��[nv���9>�R�vI������Ꮟ @k�U�n>�Je3B�%c��X)`���e
�f �M���Õ�(lukX�ȶ;n��H[��4����� ��`���3R[c~����Te͚��fR4˔4/�������?`�H���V���>F��ږ����l�q����
�:Q����dBCW�>36V�W�;oA���n%��>끙v�N�2���GŬYM���s��3Ҩ<�hӢ��)� �v�HW� ������O��8i6�ܽ/��f(mj(]�w�}�b��^{��0������n)��PQү����[��<'���z�w���Hu㑐;%��P��$bG���'bVi�- �[���#���_U�]�"���>�{0��%iHwHm�Nr�:Q�23��k?����`���~<9�hɪ����(�	�tS#{?�%���1�0C?�����6)b]�#x$�mg�7N���La���"#
�E�E����[d!qM�����a)`3s�����z�X�`3hfX+��j��13��5�La���zq6j+���1���H��u��t��\O�-'_[#a��oǷq/�:���n�9ع6�%��>{��V��M=Ⓗ�|Ƅ��3V���o�k��~�ؐ����`h��~݉��XҴ�"����B���¦B��u�������x�Z�y�����tHKS#��f,��o�u[;�m�[t�5%�!���߾��I���A�]�i)�X�M����>������6~�U�j��ƙѺ3Fm�t*��� ��q�:�@#���4a8i�9O���.=�i�[�����*CsqCf��%�h4<�a4.x�J7]���&�ϟ5��V�:öV�R;jګ����s�gv�a��z�`	��A*���T3%�^t�'a`si�%���&d�[t�ϗ,�<������&ɤ�=Ǧ����5yKk�ɦ)��Ĭ��dS��,6�R�'�dP"���}`�8����������o�;"���� ��=�"{��ŃfEy}9�y�Z��2����X+iF��#��6{��Y1.��[���l�r�2k䦹�O�+tW���焙օx���i?�r��f"D��I����51�i�����9�oL�.��뗀U��� ���/ |�Q%�T�,�h�tg#�ޜd&&e�|�Ʈc�*�=����ܘkS$Ęӫ��O��v��Q��'Lt�%����IHk��A��}����D��;�S���Hk�]sû�eg��L20���5Uv�p��H��{��$�-6P@I�]x[;+|�2I���'^�\w��
����dt(r(ˤ+���X��7дF�B�ɀq-��9�v��� �52(�<�T��컃��#�6�Y�?�c���=u���"�`��zM5���0�v@ P|�v�ػ3�_��Ee�2d�N?�����U�g�8P�\�H�7�jm|��e����S�����wؔ��]m+igN�Aj�>�Qgv�*������_������P����aݸ=����,��ۿ.�v�&G���f5�YW�V�M;��e��9E/�����-pu4z����%�(�i��~����XO�Lf��:��6��wb��1K�v������C鏃\�����޽����L�*����b|�O�?������NSXz�b=A�R�dʵ�Q��Rlc�������9��9�\��&��Hh���۴jY+=�Ը
���qB'M=�=�k���x:�L|��c���Fxg��:wAtG�7������ԯ��)���^�:z(!��Q�͘c�S]��@{w���3��f~P'���\ߑׯ����hl7�S=I?Dz���.nT�1���31H���!O�jW7Gi�%,����#�{�˼��� ZZ��W�P�_q�8Xf|�y��3�?Gv�q�ɤ�12�1R+%�Ѵ�kHM2#}�F`��WP��x#b;84J����Ÿ�0�Q�������DF�������}�Ph�qPE��]��8��C�l�,��[�I�����/�Z^�Z��FV�U޷�J���Y�� �ݷp����Ru���4���v���-��{7Cl����C�+�t�)�xNg�lz�*'=�`�g�?}I���0㰬��K6KuK��1�l�n�W�,�0Y-r�{�~�f�>o�Ћk������B�L��2��7=�HϚE�Lt�d�9|`��P��+b�]2mj�f�C�cN��#	�N}���\*~)�1�<z�V�<�F0M�V�sF�a/w��{e��˺�F��t��SҠ�E��%����5B���&��$��+K�QR��*�����=`8�H���&�%�"�������u���n7'0��B��vh�������WX�9���ȑ'_s̱o6���/P��v+6X�;,Z� �g��孊��y�=7�����Qp�i�귺['���9�I��m�ֳ���;���!' ��A0���F��_!� Z�[K��S�~���/a�ۅ�}���~���,����ʓ�Ԫ�-*>�As�a ��������ޜku7`�����gr�����Z����qݘs�a@}�n5MM6f9�cm�σ���l�����*�#����ܰ�D	������P����S�LUς)�L���^�5���ʊ7��[e��He�m�ihHҧ��>��}}N��k�15w�~�d�7��p\���Qjj�%��{��P�t��Q�P=�ȱ9V'���M����4�C�9͛&V���"�I<���z������u�����k��8��#�ҊL��v��C��l�G��x�sZ�B����@���x�%�OG��W:��u9�z��BU삇���u���@fX_�9�酓�\����.�6�<U2n�y�"C�شȀPb�$'<���]ޘ"� 8��ec���������ߙ��Nq�id]��\5���͡��ղl��q���^b3��$��Y��Rw��EC�S��7(�b=�z��uMI51���;�ͧ�W�0b�V��g�,�z����0���,A����C���<�dV��\(�>|�������u%�vpŖ(�L��ӈn�&�F?L�����~/�l�~%�i��Аk�x�#)a�r�rȃkq��b�{�'��k3������C��j'L�6o1Ew�M4w2L�	��� ���hnĕ	�R�!R��B��f�a����D��^��qT!�(n���(�/\�5��1)@���.�5	��1�/�:]BYg�Ȩn��@��l�!R���ՐG��L��ݥ�H�d����z��=�. X-�*Ӝ1���x/�t��d��͈SZ����Y���|δ�3p��8��#.�\J�*eUK%���-��qd�()�a}��̚�L:�E?�H���I^��a�7�'}O)��d���iR�Tf�z��͈�BN�c�;�F���?���
���1	���2�%sμE���>G��,%���f�L�ˋj`{^�)��{<���xDW��-2�e�xxq�e������Ǻ��i��Lь�C<̍�cY��և��M�k�����b�8��w�ky�X+��hd�F�s:�}=�J��ԅ�?;��P�1k�-���~���{����V%��_���#pd��7y�j^Z�6����D��qih^�J-YyCދ��g� \/l�NI�µX`{ JyzE<�x*�TJ;ՙG��kC��+���ԜS!ƒڊ@�Ϙ��1<������C���1�7d�hV�*�ką�MԸ�k��%/��ן��j���>#-y!҉f���x�"��k��� �NBq�J�
�QF̤���ZeR�d��"iX��j�̡X�?�B� m#W�^��&p]�X�wV�6Nl�8��C_g)-��-K���Afㆰ/{~�A�����0� 7/�)c�-�ʮ,62)4�jg}��}v�1��WHro����,�׸w������<׸+�����鐝�#����i�;݊�ʱ$��/�Gl�qS*�Ld���r�N�6�b�?��n���B�3�%�˯����r���}���D4��@�'M�r����VU�F�D0:�˚��I#�#(Tä��Kn����f|tM�;�[��[��x���+]����?�����~� �7G!7Ɏ�iБ�P[*������WI��'A��sϫ�v60��=,�u���>�S�+a�j
*����a�vŬK��:�I�e����,�[�CW�O"��8y��Y��@�g��^�4����5���Д�
��!���Z�'&�ݬ�:�8^����ܿ�]����A������{*"�*��$����ˉ%�G����+��!��lz��녃x&�A���/��z	x!M�j.��6���JN�18r7�� �.��$����ٸ\cu�Y�Űr&}t_ů������(��:M���Hhd{�# �t���-� ����-�5�#^���9��2���7N~hpHoH����==kP��>���pP!2!����8��Q̮�4��;�C���X�z�3��`�����[�fѡ��cV�Tp�a��\�1�T,��Q"�Q������M�n��������m��;�d[ra�N�������3.�������͟x�at� ��V�R�VR���*~z<�q2g@�!���~^ ��z{YF�:�mz���Kpzeds�w4���>�1,��>,v�Zv|�]0�7Ŀ�j�&�����'7�ڦZd�zB����0锜w��2[�]�n4�4>�g�;��N�Pu҅7}�wRυMao�ƀX������c/ը^U=���_������&)�D�C9:���ֽg����Ɔ؁g��#4�-�uB{5v��+���!G�DY"��1�F�i��P���r�۾�Ħ4�]6Y�;������N�Ğ��*$����3J�5��Sx��~��(��c�^gN����l���[�ء5����������υ��^�;����⠒J���5
�UB�d������{uӬ��nm��/��hM��d�l�ֵ[�C�a�AqV��I΄�����yǔx��U����;�zF��ό9H�j�����z�>���������F3g35�Tr`���C��^_ϊ`���&��I�kCI���Y����-��ki*�ɞ��]��>g�M��6�c�`��V:�.yHuR[F�ܶ)3�x��{�>`�W�_?�$�+p�]����#NkPJ�V{L̶f��~���l��z_��
6 �A���\Ԏ����J��g��h��t�_��.7�8>N�r\##�A��4S�H"�Z�E�ĿXwfn
W�#5��(�K���Q�t�����ڛ��63S����l�,p��BVw�5Y�y�?ϻAn��A�\d�X;��-���*j �#�8���h}{||�S�QY[�_V�g�2|u�W����3ز#\��0
j8�i��{3i�6i"8o���8�Х��\��F5:�Į�����2�tz����1k��͢�V��xt�\Z�4�HOT�q�Fj��{@EK�W��i�V��=m_�8�no�|l.h�9�V�������pA#>���(c�L\Ψ��&�U�}��C+�N{_UU�=�����8F��Z`xI1�0�p+A,��;�I�2]�P�6��7	�9pV/XO�e��d/& ����բ�]�қ�!���zP�����0jG���mL*Ⱥ���dm�/ ��fV����8��F�l�t�k��G�XxZ|�^�����J�nr�)8}��k���Y�X5���-�{H��t����3� ���N��|�I6G���;8���b-A�Z��$52��x)Q-I\e~cc�daFmG��Q��R�*1����F���}t�=�oV&u+����LR@T�ڬƣU~ �Kڲ�0WA��]�e<N�D)��
u�:���I���|"n�Z�4�����=E��2�b6�\^  �[%�}%�;X�I��e�+�sx#��9d�o�8�PUq$L="��_>�l;H9���D��ob\�LOE~��%Tt�t�b;�а��	�'�����$������~Şϻ���O���`b<��VZC����hj$*�r�X=P�c���/����K�r��ʿ}�a�8�0�n�<�@��;�9콹9�m\��l�&8c��HVM�e:W�h�5Č�P۝�M���{�����"�wi�C@-:q�%kt���Nt#�N,wB���|��:�D>�������'�=�$K�$1$"2�XW5�r��;|  ��?�Nng���Y�d�����{d�άr6���2���nn���Z:��ٔo�d$��-�R�kz~5/CD����c�B�����T���Y�s��Wwp�@��8�	�A
�hRr)1V�V�����&�>��|,t��4%�^R����
��VM��� ��[F9��=�A�3�#�ͭE�}6Ʋ�8J���V{bun*FOp�q��TG^WȊ�mQ�a,Ȯ�1�d�\a���ZT�2[!��Ї�����9߾5�M*���1���cR8`�|�*|����*���b��3��s7�c����J~=϶�a��uU6_�!5��V9Gqu#�R��u5ӥ�+D@f���)	�)CW���2�"��IK��b���߷��]$��hҦlq�I�(5|i�Ä�+���J����QL�!a���/�CUd�
3�z�0�����0�
��B~��M����CH'w{Q�z����������7�.�%~����?�̽��+X/Q��ǵ�,39��Ob�<C��Xl�����陑
�g��)ͅ?��.%���fQF^w2�z���._N�o�����!����Ϸ��26��E��2�.��^ #�>�7��{��h׿��m�>�%<;��$B�4�l�puAn;��Q2������3ǂ�G��
,*:��XD8���C�j^հ���2d<�%���u ���U�����5�@��#Ow/���U)�� �q�>�v�N1,���Dխ]26 ��j�V�>� ��vmq��$J���}�;���<ff`�'���`{�,�i�5�
uV����U�v�<aD��ߞE�@�on��)b��F|��ny���y�}���k����/�R�Iה�TI.���s��S��w1�n3!��\4�F�c</��0W���GR����5�!���+�5%�����3��A���A�mf^��3�u�C���'1S&A��,k��:P2���F���7q�e@yV8��.u�K��]f�E���S1�)���OmF���5�67+�,l��c�`���2K��)R�gm6)����t�R���1��zqH}�{�%`l�Ab��DK��>ŔgQ&R\E�T����u�"�4K;*�?{u�X+�f"���˵p�2�Ah�����R4�4����(>n���!�� myb_��(%��W�v��uv�Đ��j״+°����$�C�X�U�M���ʹ��ar�*M
v����E����oʗ_}U����f"!�����Kcf������t�2�X��3�g�A��].6ǪER�|�{�[i>~.T��t�e�ud���ͷ�w1�Ry��TBõ?+�DpO�w�j��=�Z���Xr�!	��,�oe�T��7�1נ頱�e�i�~AS�kf���4Y[��셰z����ɘ��ʲWң��4�6�3�<�wr��}��_I՟VѸ'v;�:�CI�ڽ�b١�Y�>3R�\`�
$�]'O�Pm�\/1�6���\"(��P�T`����h>0X�t}�cr�D|I[yf�S.�i`?�n�!�N�۬�ﲴ*���O�1��Q����k�R���g����]��t�W�LN�� 6U��HTDv�k#��_�����
E�U�+��%����1�Hky�j���3��mR�w�Tα���}쎕
���42G�#����i{��1�c�XV�w]�Fd�z�����)hR�ؘ\�ѹ�Pp�6��@dC��?�<H�_~��p�.�'�`�lh���.���6f�����rCo������ ��,�r�]���'��^�q-���(���:{/1>8�j'��KEN�<��^�/.��Fp�ȫ��E �I@�p����&�"��b�
�4S���e����i�{��WG��iF���?��RD�/�b����3@�ˮ����zftrk;����EU\���ILZ�(�)n�5.ɟ(�?��`���t	��Q��j6�@#��Pu)��W��bJ�*�ոp�x{�nB5�c��[���6�3J��8�����esg�AtI~f�g��R�g�����$�E��}ۋ��2<)������Nn��_Ӕ�e�:5^Gi�h��C>"�ɱC0���!(|��Z�
�*�J���]Փ>`� l�zaQiة�!c�s�#����eá��)�㺤GLN��U ��r٥��h�Y��c�
T��_ �~�eS��'�ܝN�����Y��s�c-V��}]'}�1�e�K2��Px���ShA��鮀@�&&���cb��H����F+o��@�Z�>���^���^��w����(�4O?�r �Y=|�Pt���Iy���`:�@,��� 0Zx?A���HS� B�<�X�do��T��@Rr��t��l�@��1��P��Ϻ��)����>��a����>���2�����賙U�\�}���^��m���?�M��	�ҮN�[��n%V��J�馕�7�J3.����ԤL����Q�����F	6���	��W9^����a�9N$����T~ `A"|>)1E��@��X��$�!;��4?$	��]d9�%}�}=��^�@VR���1I���1�Z�Q����<��#���|C!8�����p ��)���y��dJ����D�a�'��SG>�"�$ ��Z�P�r�Za��'IJ\�_}�uy���?6���(Rr��nxP�T���Dd�] )�HG}G��:!��k���4��W� 3�E&q�C�Al��i�vb�̂0��$���#uW�'U
�����^�d�Oܲ�N���8T�b|��wܿ��ǐW��K:���գ��)�+3�]�W�N� J��B� Ho��5�#��X�H�T��pS��ٳ�K'�`e"������]%ܻZsu[㝼��KWW7���j����G�Χ������SoI̒|�zc���'Ƙ�z��}<R5>�m�3�?7��wv�Jxٳ$%͈"�3F3d���0S..���6(����H�FJLż��i�]�vĄ�}��j��OC�G�6���W�6��U��=`��c�-���$-�^�S(�������I��z��Sb����7&EۊظVu4��J$,�(�d��	���Z��5�Ȯ������6���R�~��uh޼y]����}�P�g⣲�� �!e.�]qI_��8�ҟ���%戓�JUW�釡��la1���"��\��)鯂Z�{B^.($���ߙ�EtV�n^i�ٸ�iX��i�s�1{�ݻ�K�=��f[��a��݉��2��4WQ�vc�|:'t�����F��Yȗ�$�A�g��lpkۙۃ
�O:ݖ��/>dYZ���c%�fs�Iy̞�O0E�р����db5J�����Uoƒ}�j�S]3Nv����$��I��{\��mZP+o�{�IU�gNC`E�y~/y���HP�e����`�1nܜ���t���w����~���3���b������ǜ
��)'��t:j�}]�ᦅU�,�k�~���n���  Y�$��UM� W�pgp��e��"1L6��@?3�DJ�Bl���la`��8QW�k�-�r\��.�.rd�]:�Ϛ~��1gy���_|Y���?�?��O�Tr3(U��%0��\q��&Z�p�օ����C�h����a�I�dp"�۵��U�����V��5�n)�գ��3�k������Tum��8~}�7�T*<��g�fF����dS�f߮��F;�p�Qѫd��t��l�D���Pzᒻݒ� y���fե{p�
�n�X���J�2ةՍ٪�asMR�Xq].&洷�	��6�R�X��t:�����4��t��}ڀ�C��,Hc#͟�H皑*史8?춱�}r���',6B$��,'�lD�v7uЇ�mt��|
���Sf�P��v���e������b��/>�r��w��%�����sp�t�r�n��_6���!p���5	/r��0�V���[���}8>^ܤ��L����M/���#1>w��Ƶ6�9'�<gl(����(�\���M������f��t>p�����++��É���v���G���e�/�b �o���M�ԴZE��JNnН�Ì��d^J��g���;7F����d!���J��`�� s��K�y��Խ�58hڪ�Dq�555
�tg�p�%�L!��(�1T�� �� ���9��%v潦�d5��>�2 ق��x���y��=	�
]�zt��I�S&�~5�P_���{�6T���k�7&����CO���3�,Ϯ�^��PQ�8ϱ��(�d��CN#d�h.��)���(a�s�����ݭ��a��ګt�}R�g!�$���:w��RiF�q��NJA�ٶ���:��+&%��͖:�kl�7b�����T�o��5;YS�ҍ7dor�,�� x� �]<�����z�d7W�L4�ʪ��vP����C��t��
ݶ\5���R�����w
�AX� ;+��>����X�*�Q�d1[L�"������`yˡ�(�>Kc �E`�>���Gy����F(�o��_~�e���Ct��d2�r����Z89Ǚ��Z��'��˂��o���&�M)]�Ъm�:щ֚qF��B��YdUx>������Kz���=��(�l��)�#V�ڭ�b�I���"��`��LG�Ԁ� Z�Eާ�tUF�1]s%�,�{�U����c�b�@7�?���}7\f��R���*/�#�]
�X̥���ZE�<�X(�b�\�Sƥ%0}�����;U���!�;fN'�v&��|�����ϧ_c�'_��T��ʵ} vI��Xfv������.��D���/p!�� ���x7��5���oI�o�wڬ⡜P���B �%I�[m(!��4Y`�����Ƨ:N���A�6HD���:�Yf��i,�Hb�S7�q݃l��61�;�Dn�#�J�ɫ0O�r(��l@
���	c�^L�,����:��ˑYd�n���w�Cd��}������hP���"�qTBȈN}~�s�9���X��P��n8ĵ��k�����p7w���%;�Y��ӎ*��Щ�� ��/��u���(�LA�F6�ݐ�7JI��#��������U2GSe<^σ+�Ę
(�-�[��y����v���Yڡ6L����x� ��`腁Q��M)9^�Q6��~UE�#�E��R3��Ś�#�� T�b|����>�]f�����R�xiYK&O�x6*�w/�6j^6�ڿ�w�i -Z\n$�x��?���c7�"�i����p�&�H_���fѤ��ؕ�-g).�[a����˙<�H}�ścS�
���Ac^2jL�zB���*lL
�:�p��3P3o���>p���o�^{�Sӕ�q4�J�X`5X�
��(�p��L�&;
6Qg~V#/ؔ���.�R�&��i_���iX���]|�8|� !��Bbd�. '�j_n���7[����X���������F�e�����V����+|�;V�Zx�w�������~r��Y��rM����t���I�]í�˛����߽�o)(g���pEљȼ�U�=p���Jc�e1)@�Ɂ.�kd龜q}�y�/l�̟�ا��Y�I@�,��q�s:(8[�dW[jv.�=���sb���?�X;sD�6���0��Z�o/��I��B�Xjѡ�l�V̲�j6�/���a������:-U��x���~WZ!�� ��K��fZ���������_|i�`�^"2QFw_�q����.��i/����t'��`-��`�c���g��Ѓ��E]=�j��z��KN M�����cu�c��S�T�l�>U�}"����#���x��!H��,K2^
Q*�8�#�M���1cJK�15�������#���y�0���bk�<���dU62I��uh#�%�:���>�����TW��88�8��|��|�����o�)���-+e��.��b�t'=Җf���ϣ�Og�47<R,F�LuS������ˬ�,'`���';K�Q��B''��Fq�l�-� W��������]�(��^!���X��KU�ծ8+�#�&M�9!p&�{vZ9wn���!nP%�ǞX�=�c�h`w(5a�#lU&�$-��0W���8y�J�t�$W�Άw�)�z��:��ý\'���W�UP�ɫU�}c��9�yD���覥��P������i@힆�� �Ͽh5���."�%��O�2zi���.���w�4x֤Ƒ��6��60d�l <$Ԧ5q!kS. �g`>��m"�M��lw��5?��շz��9u�N[���6{,��:Q4��+=e8�h�J;����E�q'�D��1��q�>(H��ӡ����2;M"��Y�8zӒ��DVv�7ؚ���X�ꏸZ@P�Jtj������W�/�,_��H���#��lo��X(�}8e��'9Z��M�e�����Xh]�V\b��5���5�+=��@y}E��gG\3>���N�Tv�#�-�����N)�7.�"��de�w,K�JO�o�����/���['�����V��A���-4⢍�f�52��0	�\�������L}�OZP�n���V46� �1�eQ�}Ⱦ��ȠI؅:Ʀ���u<o����d�p�oVezd#
�Q�k��>a-6*���+�{�Z��e@-������I6{�D� � ً������]k�fr�SŌ�3>�� �5&���o\��=�Qr�{��Y�.�L�o9_%ݖ=l�:n>��P"G�D�nܨ��	������H�8f��kh�~�)V!x;��+�vj(�B.>�3*��!Q�J��}�4�F.d�M����o�ʼ��t�Bz�����������ge�T/�H�����eL&}��oが�����&r��h���J>b�R�Q�I��#X�%��	ZWBL5k1¥~� �g|ཪ�ws�&ɵ��xU^��yL9�M��3a��ͷ�ˀ5��6��<8h�bnqN�lȞa��e�o߽�.�?���H�;4	�:i�Ƹ\����]�A`]=�.������(�h�.�`�Ǟ�>0�R���k5ՌqY2�ζپ��E?1N����-Gpc�e��Y
�s�>�zxo�ў,�m���8�{v�����9���:^�$�^�Y�
�m��$��K����0%�7J>8�G�f���_�72��aB�0>Q����)��Z��ΰ	ئ��*�q�Ş%pB�*6EH�o�qh��@?*0/�'~H����>���b�	1���r�H���r27~_�/b�D�����C�q��K�l@} �`��k'�6�OĵL/�~����Y��f1Q�C���B�j��{̝��Ed��~�m�/�KR��p�׃�w��x܆�2�un�J�?H�"�In��r%%�:g3d	�NQ�u�.����GM0am2#�TȜ�D:��^U �'���9,�HƉ�ב��),d���Ͻ������~��
�T��������;	9����C�Uc�&��;������b�V�������3o���DՓ	�jRЀ-�0���{h
l��W�Y������/��]K�����ۺ��J���^=4��Ÿ�I�ԈFs�]�j���3K���灔�88�q�r�2E�L�v�a�ՓT�̳��!}��6�dŬD�&k��䚷�Ժ*F0Q�/�p6MS-�"��{<��av�n�!&DzbNv+�f�y��:��/;����Jw��Eb�KJ���d�8�0��|�m������w���i��^k�+!p�:lg�Ц�T:-FJ5L�'�rlF�8^���'y��)��s�gqo ����#��S�3)Ll�yD��c`�h�{� � �&�\g}vO����ʔi݅UG`�UZ��뗋��� VQo��cε��1P�n��g�s' 	�'�L z�f�9x�&l�,�}��e����{�D=�_��iw��"�7lJ�H�=f�6��'�$��W�#�"�A�C{�*�Ҍ+�+��4ߙ�ui=��W�?kO�f��@ox�� &`5Nu]�-zUN����6걓��;�Z��^i'���e^�f��P�eD�'�Ԙ���[	���l�G��#�eǌ�s��dɸ� Ύ"6p�l���Ml�lH�FT/��|�X\�sl\|������Ѱ	_�+5%f)�ω��w�(B7Qe&�*��9��43�����J�Hjj�n7ʚ���q�Vå3��97%(���jZ�Օ(��H'�5��(,�kS"!Ԛ���,Ia;1�ƴ��i8RT�XU�����1'��W_Ei��3	)gٮN8�����n��`��(�þ��j��f�F����饨Jxɜ1��]�1��6���D����d)���������>�� 'R\'��P�Qk�?���=�� l��O?m��?"�����/��x��V�7џ����s���}W�pks�������5̜<3HUq�>3��Kb�e''�Eb ܃{x�B���W�yj(f��x5�Di���ke���������>�	�Á���0Ǌwנ�O�~��TN|~��jgtL]��eT��@����@ʧ�ԏr��ޤ}}ĩ{:�EFc&|�����b玞I���<�v��1�����1��n��+�n�<z-4O/����x�'��K��\ѿi��zՌn+�� �N~�Zdhp���e(�E#:o����i���򔿍������J�� �$�[nrQg�1���T.f�Cv�9#-�(�P�&�����>pb�2��G���������W_�"�-RDQ�#y�75VZ�u7�vR�w���n�aټ+� X>S��T;vd=���>Cq���	�f�rs*nYYF�/����Q�w�u��s��ױ��P�X'���w�`�������DE@���\8�`M��,�df��<����f�x�b\�u������ ��/Q�@�p�����z ϢҘ罻��{mHJB|Ʊ"�Z���Y"	�$�N);�hLo�-�)v�X�j��^����5�aX)\�8]xyP\6��D����7�&(��'�3��9y�TJN�SZ��+gZ"���El;dO�R��V�.:�A[��;C�DXȸcp.]���s�h 5d�s�X�.Iڴ��wv��M��l��qJh� cb1XX�������IE@8��.3X�ۄ�5T�e�p���}ƙ�}Z<ur{�^��U�x�?�}�0�s��X�HX�gN�`@��C���u4���6��/o)k=�	 ?޾{��CfC��+ )Ȟ�+�+o6C(�n,�[e�l�)�-�b��Y�4bcv�F-�_�Y��5G�����	3c��f�� ��?��K�e;P���6�d��pܴ���>`5O�=�cvW�actUF������$�2���k��/�IЍ�R�=k��	U��b�>�Q�OVIS�ꈷ����z0e囈d��<{�����1u#�����Y�������{͇���<������D�����_W5.#�����k�i0��cvi����Gc�C�5���:�x�UŅ`G�����9/:;�Ke ��MЏ\��TK�dL���8nx�����5ʗ���ZO����~t�ƀT�����_��x�5kX9N2�a����<��)�րot��'RJ��£�������@\�P��dH�^A�Axɉ<h�A�c*��i�@�Zt6I�;�E���\�cˮt玴)2�י�>���*�s��]
��9`8�U(��!G(}�����Ҡ(�̝�\�u��*d]�@αF��?��c������-+���^�4.M�<���g��?�e(|�Ӊ	Fe4l���:��}��[\PZ�����N[��M�&��9�Ιz6�p�pm"�H���F�����{��m�ջ̦s5� `9���e��೸���/ۨpW8m	B�ìTR�*������68����k�S�Q	5���k������L���h�!�\CZI���2,# ��Œ>ݱ����9��f�Y�:N~x��׻�2'����!�+p�@�!ށ�j�� �}�O�g�I��>�Ն�N"J�[����z��{۞��jt�/�UyM��G��~�"���1��N�����X;�����h]p�ʘ�g�U4SR�<CH���N҅���,���3i��%�R`1 �$���M"�Ɛ�K>|��>i8����ߘ�;�'����*%[�* �҇x�9�}�#]����z��2�3É�P� ��؈$�)U'�+pA��i=M�G\���;�2�N�a��Y`���O����e���E�F��|s1��.���7����B�e㎸+��1�����i{0\l�3��������hx͕,�@�u]�������/_�d��&���:����9I�ґY������a��Y!#8Q`d�ޓ��@��I�r�ќsF��R�k����EpmΨHk0��uU��"�6�4�I	�#t:#�*724tn߽���77Cv���1��	0ɔEF
Z̐�Q��5K�;�"#����iv��(���"#�e�$��I ���q�C��6+2�/>�"v=������b!E�&�[]�	�}�b��/����|�͗A{y��m8:bA}��Eཻ���z˓JM�L�9�`"#b�O[�q�,1���)u��������\�S��v�M̩���r��H���Ў��Rͥ��gB ��N&w�!��;�q7�B�(�qH�w�c�v$��c�,�5���o�)�|�m<§�l-�s���������G�@��^�%YjC~�+�d'�UpH�8 Y�<��8X(�� �pO��\�����%^��l~���o񖀓����D��=�e��Y[��MS���>�d�Q5���|NfμL�;�&��-��~�_AISƏ�#H�1Xq��E�ac�������%�|�x�c2)�:�7�Pz�\=<��ڍ����dŌ15�>qѧ��E��ׁ��������M�L�s���R��%7}M�;��A����j�n�^a��'F�"G�]�>QLt�W�e)�Ow��%��;��q3� �6sBE�X[e'<4���U⺌�>�i�6�Ȕ��9��3�P��(2(��hT@�~;X�&5�A�oS��H4t�S�R6*���&r%�^($BE*ro��/��j���;	�~'A�6�dL%�;�Lc���.��v9�)����DWׄhd.�ǝ���Cy�&���܅���A����8�8���,	����W]3oؠ�a�3l=�%d����Ę�-6��|ƴ��3N�	qݐ \؝��y�=�"C�����%n��QǺfv���Q�/k̳���3Ձ�#F���e׃ʊ� �dc�Ɇ^*���c��.1�[yM�0�]�]S�;tSwH���h���^B�pC�J%68	���ۀl�l8�:�ٍD"��b��r���խP�����x�/y��'��40���Uj][�S��h+*�z;�c�]��q2�$C�(7*��i�e��yJoo�$��]f�Vw
���f8O�{�/�&V}�%$ �)	'	�P�v>oA.2?����@L?K�<Kx�����6*�aO^���c�m�=%��(��6�����@�Rѡ'9�U�a<�gM>�0�U��a�I�Mς%���>,���D�w�G��DؙkԴ�|�����$ �g=Ŷ���1f���yC���4ixU���C����۳�����l-��
ݛ��t!hp�P;����_�ں"�B�K^��*#p�����*���P2�����>��/# ����cв7] ��d���{_X��@�Ή��O��N}�IJYUSw栆Dw|Y���W�К$�~��\8F��'ڤ,ܙt8
\��e5��$����z�����;&A�*q�8�� �Em��qφ����X=�;&#��y���E ��X���M�&vmm���7�i �i���)y�R�(li=��uɓ�4� �����MR�	n�jY�^O�^=��,��LA�R�"�g�E���wB2R�0��y�ir��5OF��wZ8(7V�����2O�YI�����):�;np�����Mx������$%��Qn����L�:GYW����ӹ�ٝ,W,\���Q_m�84�P���C�	�,���M�RK�%2R9����m�RǸ�mpFQ���h� ��-�e(*}��7D*ቩ�� 9���*��{���q�{Rs�q�������V8aW!,�$���⻾y�yr(��#p��᧟&�`�;0����a ��{`&���Q�S@���$z�j�[�2t�bϨu������:%�m=ȆI=�'	��|�a�5v$��kg<�d�q����\<G`�A��ljH�Ӻ��Hs���I����D{���5�k���P�'��C��Ω]O#B�{����]��[h�hئ����'a���8}�I��i�H�t�bS`Nк�^�(�M˱
O!f��C���a�T]��`�/	���<�T�oŋ#@�x�d�����>Ep�N��:�u�cy�����Y�|��R�*Kf�.��W���!��e`���w��p���� ��#2��^�[�g��,�ҀjΚZٍ��0��Ԟ��x�EG{-�Y��6���*w!�KK���f�����e�e��#����ct�Ew�ꡌ��a��PX���������If�1�/��ux\�k��	6���i��L�SU�"�(�r��-Cf�ʇ"�!�h������Hh��K󮛳B;K��a|��%'Q��\Y�CJ���&5����ʖ���;�p�y,��r���s�a:h8��N���E�ǆs��I�3n��p���.�gi�I-cW�N�Fp�M5Z�w�q�:��б��Z*?����^�{�{m�,���|�6#5��%�>��ul�"�v�N__�OE[e�����/�*�e,�������US�CŧS��6�ZK�T���/�!D�8��6�s��Nc��������e�!zB5��6ے%l,��T���q��,Y{��yW�M���+�4��rf,S�N�@������-)B�Px'=
��Z�9B���,ߘ�x+��[j�&�^��O�d]��ԯ�D��È��,'�h��Ӂ�C�z��p���xĕ���@���8�u��a�,=�,�ӽ�K��޼��u@�u����	����+	���-�Z���s�t�Տ�6��fS�e@���ﶬyˊ�����T\O��������q��޲$f��;( ��Y�JW��gk�����f~?|��t�5/5�hK%���p+= 5L�LLѠ6
���CY4�y7�?|��ho�X��^u���g��;[���2W���y|��O��oj�	��3E�� ��܃���[]�-V;g�p��;@ਦ�Ms�r2�.5��6��-U�OVY/C��@�]�Z�S FMXx��~'>]i����>��fe�&K���%��OC�nM���
�{�w' ���{��+��Xl.
/\���h�*U��@36GX��s^�1$��9�˴�����TeG�4�:�G�����ɻ-(�����n�}�GȂl�� �e�r{�.!p�}����0��Ha���`,:��ļ6>���%�v�&��&��b-�l(�Ӄ��I�+i��>)Ox�W[���5(J����D�Qd�Z{��(�����3l�����m\/t�����?~_ d��^�d$�W��!�6[v�kA�c���u�~4��n�n"����˯?She�8԰��q��A2��M�Q�|3��'�ظe�V�p�0ƺHD=��Γ��NZ��\�Ǩ����2��;��ǟq�$��pv�tS�j���jcٖ-\���b����t�<�:O��� �﷝�:&���U������慻9�Yk/"���A��G�O�������4�,��#�N<e�z��{�"�6�@ו�_�����T��T(
��i�?𪕸��,/�S���^.(\|4d,sM��yɌ�N�}�$�(Ё��n��o�S�L�?;�I�QG��'5nŋD�����\����P���R
��v;�����Y��s�T���n�x�F1b	�bd�_n~��WQ�Y����Y``�<�z����%*��Q��>�p�0xZx���>�|�����I���������c4��e���"�˟�����x6����θh��k���/�Ͽ�T~�������=�>����qm`��|�l10��5O�|زU�L�T�}e����W�A����57*���?������~�É%`��!�3|P۠B>W������3���٨&��"ړ���%����)�g쿸0R� ����4"F%��x��`�A��Iך���j8�,T����YL�NE�f�h�TI
��8D�ݥ��m�uEw�laPҖc~n7֘���Gkr�0��j��郒��L�ڮ��M]��?�G�@�}��wf�Q������3���2��i<P�>ޘ]=U֪uh/�*X�V�Sg"12�FJLt0��󒁗�W,�/�@�<ʼظ�/kH�m
A���%QB�U<w�h�%,9٥��C�Jg4��&=�P�������;��3�.OϮ��x����2Kټ'���T�  H�x��&���$�?�U o�C&l5�I�|���_|�Edh_m���_}8(7������dG��V0]�9uЧz6�`���m��~��ϣY����+������.\xǀ(pq8aF�6�pJ��!�,�SY���Ѕ����i�j)f�w{?*�A8(�4��xOyu6ga�3E\�q�UǬ��UQ�)�|�QT����B��v�i]�OaQ��R�b�N{�V����7V��U����
�k!�����~1`�=��AՕ�G�'�S�ޢI{Q���ā���d��>��şMݮ��_�������7Q7LK�l8�Y&6ǩ��P�]]GV����!H׀�8�|]8*׎�q����-�~&���S���ʊW��(;䃤�(.AN��{�r�g��b9��:�3!�<2�k�Eh����h.���,�� ȗ��D*��޽6�����c4���a,�����(�d�Q�5��KW��km�š��C̸:��4A4�~(3�C��^_�y� ��@I����/� ��쀋Ҏ�U|���B���wo# _p9�\2o�nd�����L���Q����c����s�1�9��;�3�-뒐�+&<�[T�<xԛ�O?q
h/�¶)�Ȥ�����b[����<T�A�B�?I�ד��MN7#1�x��CCV~�+�ݸ�ɹ�c���Zd�ۚ� �����5�jM`�E@T���/�����^�Yx��O����x~�,��&?Gmh�����hj7����n+uMG�V�	b�9��n�u����EY�45;�K}��@�����M�TǨ̫v����a(�+������
M��J���EAe�9a�p�TY�{\���R�cн���.�{�ۨ�s�|��0����.7��9l��Y]�fP.�]�0��/)���(�_o�:29,�yR']�w���w~�H-�F��)�x���5�Iu���c�r.�Ł����T+�S��=�-���Ki�7�̷=�Cku:��RK[d��(m������~��6���;�Qi��{�d�b�Q=��`���+3\��Е�{��qN��.uk!�{�	u��Z�����&��?�#&���b�~/��>�`���`0|H!�j7�"�o���C�k�u��!>/u.>}�Ďɝ�5�y���UtC_�F��#��ʹ���=}�G`��KT8&�m�jew07��z��{c�gJ�)y�u�� ��:�u�ΰ�:�Fw1X�'�<�l�3Eq��m��[� ��̬���wn�U=�5	�����FW�{'����k�h��Z�XT^�\���|n�y��e�g�kQL�ci����W���Xl�l5 y:��N���Fٱ�Y�W��;m�(�G�B��j'5g����˖������񚇄�]�J��l�������t���;9F =KWx����Z����6�|��mf���jb.{꽎�R��\o@G؎��U�@��Ӊ׿�-ց��;�c�2���6����x�g4�Pz#��?H�
����7�N�� \�nx�<f��s��cZS[�5f��k�'��X�P5�o�|���Y~}6Rq�� ��UҊ��lJ=���Ac���D኶k�!��ϳ�B��ؓg�#>�\�_B����k��L��T
c��O�ǵv�~߃�,NjRE�V8*���y��X^�����tN5��=�a���s����[/��U�c��`��m���Y���Tux�`��9�-J�|A�<(|XdO����8�iK���ԤEsQ�[y#�9��a�2��<�|p!#!aRp�7��R�ĝ�D�Ņ^���+ڌ����q��
D\�ܓ�H�HKL7��5R�Y�I�+_������p<^��J�ԡ��>m�� l�>t��C�^��Ț����;��
�?|���^�ad�UE��a�lt~u�a���g ���+���}��1 Pt���hL`�J�������&���@�/E��]�_���.dgo�3T��R���o"���ߕ���"J�z��}�R�SI�|C06�9G6H �/��!NP�)p�n���60WRs��hئ��5��;�������ot��ܻ����x�XCƌC�����:�����c|F�,���ͯ�i��t$K:�4=���?%�ӏ�	��f� 8J�gh���I'v��1�\�<�CPc���2���N�,���A�3���.�UnoN&�,h'�Yg��1=��x�`~52h�>q���"'���H���l��kD�X�x��b�cK֎L���u	1��`lNt56>�J���3��ZS��"�x�J�(/�Ag�lPۛ&��}�d��L�h�$����<	���i�,����g��G��~��������+N�л�0���+u�_�B�-�B�g�*cB#�0tK��i�M�@:*��: E������7Z��(����}���u���_#;5���lo����a@��A౏G�mSoµ��D'�X0J�%�|ڮ2�fF���z^��Hf�ȉ� ���3����������/.o>��|����g���At��
�>���_N�q�+6g`F�f�_~�EP��%A��.˫�S�NGX�q@a��7|���%�<�;�M���όJ���s����������L������o���E8 �Ò�*�"��ᅍ���$���������NN�?jk��YS{����R@��Y���4Df��z-�U2/J��X�%5��\u��@i�`���ԣ��6:ٸX+�"K2��i�B�E�X9���'�+;%mTCLիK�G�b`�xNz�h e����"ӵ��5�)Us�R$��jX�{$V�y�TbRy�r���2��XϢ���?B,�y2��[t��.#�"�'�3��x��ą����H��ڍ�g�YtӦh����씧|�rkm"�C`Y�f��;u�Bc)�y��O �]l���W׹@c�
�$�ӹf���D�o�	L��/>����F����~-�����= 5��n^<+_��P�"�2Q���=(#��� $��'�&�N�@Yʋ-��)��C�<�2�_~��@5��^����z_���������ٟL�tݮf�*��U���@
�R|�g�X�O��b��`��_�M7�弹'�zv|�Z�u�i��0f����SY�q]�˘͗�g�ЀV�g����������C@78،�#���A��޿-ϟ��%���!n���y��*�q`�'�eF]JzGE�N��(���hL���(T�����!"�h&�j ����8�ٸ�d}35�:�.������S�\q���ׂ"̤e���n6W����'m�7x��G�N��\�:�T6����[�ݶ�9�r}������Ԡk��uf��$W�}���c����N�
��o�_K뛾�-�O�:�EM�0X]����=��Q]<C7;�Ew�=K�ȴ�-z0�
��Y"���2þ�;��R�|�7���X������l��1kQ-����#C�	k��1���@!�a,xȠ���h57��FH�=j!�U�v�{ G���!c���^�޽Du���>f#mɶC<>��uy��M��}g�w3�Nx]��QG�xR����������PA�ߥ��NUK
0�����f�j}t�Xr�l�WB�+-���H��_��۵{ ��������8�^o-�^�V`:U��q�Q
i�;�O��4�!yʆ��O��x�]mB��w���	��s�k)V�
���9S�Aa8��C'LN(D��]�(�k7�K���Ȗ�H�8<�$9��(w��W��=mP=�Õ�f�����0�"XV�=���/��79��F6Fb��ͤ��I�D�����٤�S弝�ǱY��xc'���Vwo���a1*�eI4��_xF-�ƚ�g���V��#&�C�7ǋ�7T�����,�5Me<�(=�G���)r��t~��m��F&u#�b"��eiG^�sΆ�|ox�n�/n��e�[���#��*;�� �lX�[>"���g�2	w㽀���P�xI{�"���ڂbf�\�ic��1�&&�� ����A��XN���[~����>�\�
�v1�nk�}�C�˵�����h�][X�l���P��-A\O|�>���  ��IDATߋ��-�y�]��>���N�'�<�B_��W|��.�m��4�Al��LX�9�:ÿ��5�*sbT3Ͽ� �R�ڄ�^<��[��8uO�)Rw�$E06�㡤h&�����@�����YTU�k�|iN]�u���p_޽[��G�h���A��p�_>�`����%w�f����ɍ�&6�`�����:}Dd�l��e8��.6�i}��>�t�E�f4��J�e��xt8��@�ˎ��H�����ҝp�F�Ө�2-��A�o>�S}����[�Mv'.^����x5�h��bx�ȯ��>K!d6T%�Ha��8U*-<��)sg�)�,:`���Nk�eVVJ�ƃ7Ns҆)^��h/!��[���ܬh aQ��oʷ�|]޼&&
f��b �Ա�C~�Y�zw�|�w��)�|�M����M�[�_~��Ƃ!U��Z��B;�E3�6������F��})����`�vh"}��F�0 �]��e����ʇ��۠9��Fw����m��1�R(S��Y3R����)� ���$��u�x��: �딕\��PSSHdM/*f�5��k���	�ߕ���o	�t'xOɢs��t���Z� MF�u�h�U���Urx;N;��g�;�p>`���N��:^Rk�2���5��о���0\f���D~}=	���Q�)��aZ�e��cK��W������PV/���Ҧ�˚����i�]�KQ>�c�y���	J�WܳO���AJr�"����e��7X]?Ǆ�u"����}��7p��A�f(�,kb=X��7��o#a�<Q��^l7����\ѱvC��SN�-h(]�|��@Ou�g�BQi��5*HA:I���A�����*����8�iZ�S�P�F/�8T�3"p���T6I(ci<�!DD�~j�Ll(@A�߮/�]!��RV�e�?�����y�9�9�z�Ck�ٛ�R���Px���#1X�|8G�q���̑[LR_����v��Ӓ����}r.�c��lJ�e�W�X�$�&�t ���Y(KZ'E����澦fm;*슫Mh fG!��[��� =�d=����N09��r�q؅�8��X�HL��h����}=Mi49�ZW��.�MY.i"�m���i���OA�|r6��1��б.����Ac���=�D;bVY����r��8�@�"��q�>��8���+�@as�R��&���0)t|�k�2��;r�����q�E|�O���32�}�A#��������c��ǂ�� �	Y	��>���o�9&_���f��c#�X��Χ�" ���/�y������U���e�k0�F.��p�h,Ɒ��rR�H�!T��Y`��]�|�YP�����l� J�{͸��R{��f����5d�L~���*úy�(���`�� �#�ZCЍ��C�bd��R9�旆�������O�6Ξ�����y�}��2��!I��O������x�2������<y� �^��u�����?��1=O�.�*�����Y3��Cl�Tx�!�Ɗ�9DY[|v�]{J�ղ��6���K��2��F�X����1���ML0+>��L���:�Y�߽�eN)WǄ0g4l�۵&3�C˅UV�$n��9����Q#�ss@�N�OJ��:8�z�@�|�H���Iٸ��U����eqt	U�=[�l�A¶֍�ccV_�J�<1��1���@�C�����@�#���G�16gC�]�$`��i,lp��&���G'G�W����u-9�Ex�j�q�w��<�C@ WA�:_����K���J_�Z��B��^n��D�(X���
��t���v�Јrv��|Խ�H�h�BX���ͩ�	�g�l�@j�:.HN�E6�VM̀"���M���8,�>I���v�o����J}�x��3B�C�4��e�1����eqt�����Ѧz��~�Kg]��.��Dl�M�]܇���l:�ݟ=�A���r�?0=]'CP� ����I��w�+�m2)��Z���n���.��j8����2St���^\�ģc�����bp�N�S�$��K4d�<��t�{�ntʸ�5��S��j�rֈ9�p�݅~/���LFPɀ��e��
�O�1����ϋf�Em �����c�Oz/�-����ׇ��5/�.G-�r/B�$A�hh^āA�Z�iј(�AP0v
�y�5C��M��`����М YY�	������+Fʷ��jQ3S��=��v�L(�T6�������jϮ>Ns��av▢�t���)����`x�8dH�����==RX"3RfX(;�����������%���:l�b&�>����k��@D���Y���޲��^������ �Qu7�@�(#���=�*��@+���T~����e�(ȏ?�P~�(d󠌕kq����&6��|S�뛬0�8$r����;'��2����������ʅָ��$�oQ��,����n���o���S�S�����o�~��Ͽ�A0)�d�z��p����K���3��u]iK�q�u*�l)�#���$���%��J�kf����`��A��؃�cMF4,`��vأ��W���Z� -V~���[�Ł��HQ�a�hxd�S$${	�Ԅ��z�fDLEIi]��1�&N�����\޷���~�������j:�?�
�d�Υ�"t�B�d���-ܬ��b�7:�σ7HG�3튥�΍�i��i%Ǆ|s쒣:��$���ߧ&��"�-婿xT��1�zz�7J'��}�]�`9_~�6JU��0����~|��82��~��%�n�RY%2l��neI|�^�1pD�H�W���f�JzJ,���i�X�@��h��C63kS6Fq�"<qG�����QLKR�X�a�}{��ɻ�V��}6�Ɖ��2���Q���~-�%��Y�`�*�/�����w	��G�=���_��~�{;��QnS+76�̨��˲�&r$ѓ���� &����={����k�������?_�|���px�},_5A_�s���� *�����AL9WG֞�x�2�՚��`�(�+��O=�5�F�=�tK1���~-O9�ᠱV;@S�隁���J�� Kq��Z�x�u�t���nt.�@8m{��m����Թ��f�����t�6�>)�/��"|{Z\�Z�΋dy¡|��K�U�|��E+�v���#�����Re�hG��jW2+���n���X�婘"����v�Y��d�}ts��U�),r��a��6)F��0��[d?w�F"0h3}�㣰�ƍ�߁b��e-��wDC��N�Eo� �at����x�G���۳�1��<�A��n0EI�%����ܨJ�a�������TR
�;=�1������������[p�[\�\Q����qO��Q�2&dǯ_3�����+���#N��	L���.՘fѰƱ
�x�x�������3��g���ա��_�w���)��u�Ѥ5	ܚS~r��E�|_<nI:����j�'=gU������kv�Ro���&U.s�4��6_���|��=�I;�o*�1r�wÒ�E���/N|�����=�"J�=ଝk�ی�x��JZ��+�%�q�?@?tf��_Ү��H�������z��7�-'|����&A��~��N��x��t���>F�0�@m�@^@�H�ߧ�.�N�)��I��T�-pȓ_u�y17v�����.��(��+}���TP�-н�)F��Ѳ����D�bF��#�[�	-O`�hp�u.����H���xu�_W%�p�f	uu]1�=�H=������ڡ	�##=����Gs6C����\�Rz��!�lD���{��������Cu��g�A�@����������������Ͱ�U�����
��?
�-5��T�APBs@��cڇJU�?�c�z��W�7'�Na����}.@-0��a����Wo5w������BG_�Lf�/E+��;$�u:��
pO�rc�L~^9i��b�����d�w�[j7�2�"�`Fz/і��8���V�E�$����Ie�
�"Fnփ�9�*�؟8h���FV,O2[]7�x��}φ�f�A�v:�1f�U��g����'��l����?��&�*���I�����K�ɥo�0mԯI��&@Y��[�:�,�`㵽�հ��lY�(=V7F�R0�T�:X��K�9UD��X���<��/1Z�w��׻��(WW���� ��l���uJ�&�p*&����o��SJ���gP�y���M�%�h#�c4i����]d�6U,,���F�̾L%�&�̓I��������G ԰ٵ-h��V����@e�_���ypF�Ɂ�vG�1+9����(,��,��V�ml��Y�ڠ�f5'촐8���8����M_,5s�e��ξ'��8��t�2{�Il�G(�o��/�]�U���<D ��>�2�e����v���"4Q��Oe�J#򞹤J*�(��+�����������(<�x��3����.��!�(UY��eb�� 1k�ӏ�Q�$��X�3��b�Yf׼5\T%�-W�����ൟ���S��|���3e,տ�������L]Z�7�?^ ��T�9GlJ�^3ၕ=�������iv�y
�<���,�7i��<f�	������8����?�Yw=�,����?���'���A3��Vc.��Ƥ�N���,��$�S۴���ߕ�U!3 2�㣂ω�2�� G�o�5�73h��|Q:�.���޲�����g��C:��[9u��t(��7���!�l�e]Lu�%u{�Qh�zѽ����DK�W!%xw�<2�'\�y�*&��䲛dwf�>��;mY�a���,�j4]�Ze�C�1���MH��JA��g|�uU�ULg����T#Z��`%������l}!.x*�����U8�v�O�W�c�5�2���A���{�Q�p������UZ3��˔3�[��Lg9��x7��!��|�/j�ӕ�!8= ������N�׭i��s��	��]�&��贸�|B���%��IH�>Q����o�5�_�y���,��Q'>������Od.�E��{�L�]���3]�w�кa��XS��؏9��q�ܐ�I� �ȴ)�a�Tܗc���t.�w�����Pxz��u�'Q��<r� ~��3�"@"P#-G��u������y�Q!�b:׮�>�h2���0˳3K��*`�N~��3"�.z����*ȡ�A0iZ��eb�t_r��t�}v��/ބWՋ�����תV8��'�13M6�J�!lH>d�b�S�@z{'�)����vV�*�6�8������e�.|t�52i�A�'|&@R!xk�2rخ�!���b���7S5�&��8OY�[l;�G���&'�o�ZXE7��	{̒匀���!���K����]�Vλzp�q[m��B<ڬ����{v�\�vP [��gC��&�ux�bĦ>:���F����<�]��~s@+�4��b��f�-�I�k�nS�V����zp-ހ���%n@4$`�L!�ҏb$s-�!�J�A�/fE����|��ӹ����8�y�U����+� ?��j�KMe�W_}2���_ߖߐe|���UF
u�)4,��)Q�2E/r߼�T�{	i�NA4�-{z��e
<D�>�ʌ� ;�ef)֓�o;ZHk�d���!����©��fFhT8���GRW"�R����*Kr�o��!a�\U��pƋ�xY�c���N�K��X"�7yn��g��������}r#-��=�#�<��~��DZ�|+��0n<gFJ��}�}��(���>�8���p�o�鞥tU�EcEp�Z�u*�P{M�H�a!��vD�f�
��A��R!�0��F�$	��s]��a�����"�u	
��c��2΃���i��.I��P3R_/�C"��2���k��u5#M�o]R�q�,���q�T����k�/���=��]TF7�������P<���Z%��fPf�Y)'�]�b�uF��.w��?��å�񔾙�������vgr�@�Es��kk�Ic��[�|S.%���A]ʁ�͚�b����A%�&�.Ơ�ס6�V�������BlZ]��5S��\Ӄ�&q�����t��2�<�m)����Ta�uM�{hJ�I�4����w[��ߣR��w��ML��V�C���l��
� �'|��.�)g�p�>o�Dٍy�C����Ϙ���]��N����D?׃DU|p�%h]S��9�J����m�Z!;�����0u���C��&�t����^L�MբU��Y1{�m�Fs)3�&1�����MMj09� �A�WRЭ���������������E�	3tM�6���&K��֪M�S�6 ^`�Pk�ZkH3F|:����NB�=�X����r�%�L���tJ�F�I��.:��^~�}O����ғ���<>1t��X���g��V����э���ލ�!3/� ��_��KhzFp���� E�l��
.�F)�M�!Sk��`�N�.�@o��ٞ��N�#��������|9ZW�^�!�좊 K�W�x�_����7+��ch��S�@PQ�W[r����Tn�o�ci�W��JI+�暁��������������fv���m\�B�����<���
MC\̛�y��ġx�ֳ��2R�j���G�H���Uф�؀ԙFVgv��Z�f�a'����@/˚��e�ChLM]K�I�a�ks�CY���{����*�޲Wu�c-���8#D����r�贜�d�}~����I�3JR�� VS-u��=j��wc�H���R� ��Y�3,ӝ�c��~���MO77�?ٵwF�6�yZj���f���dB������#>���tb���)f����H���^�u(h�$14�6A>��Ѯ�C��P 1=bn4	gQI�����L���,�u��)@�Q>'Ή�� �E������l݂(g��S*�t�pW�iM�q��'�N�>�)��y�� ;mj{��U��t��z{
y�I�0� �o��m�F,39�tl<��
L0Q��v${����V�8Ȱ	���?��`�i������E{�������[f�h�Dvs])��G�ܜU��b��Kn�_�ɦDS�l�M�˷i�Rg�:���G� %�@�������97iCs�n���V�{gIʍ�y��6��w��3e��������ֺ�a�a���l3���`�6�A�4�e[0��q[���=xP8s���1ى5E��Ks7�}��C�oi�����kVc��t���C���'0��
�����1����E�DJ�˙S�,F���hz�؟���*�c�*�����k�굃f��R?�ʬ�i?�G��!kC�r�[唝�x-�K��X�X����Mau~�vp�ݕ��d�F��*�)�L<�+�=7���dx�#SZՀh�+�1L|�b�p����
Ii��j\y���kg��O��%��i!�\ ����r{�!��Pjڂ�*��9cbE�r�*�D�$�?�! ���q���۸V]��\n��L�����!�o�A#�0���^�0p�C���Wu����]���e|���x�".���gE���`P��Y��Vxj�tͿ�}��V?�{b��ա��7|��*j�<�6�
!����A
{n��y�����0q���J��u����3��s�k�\Q�`L0�"^�)Z�������sm����Xէ1�4TR�.��Zi���L?���i����PoN���(Z{�� S.�H�9g{�����i�����D��H ������xg橖Ķ��u	G��\����g9�ҝ�,Xl�~�rŠ���ͭa��=H�}���w�Y��~4��l��ն��L��T������V�)��h(��-��>�o+�`���i~�L�#��-ʀ���4�1���}nw_���wAm��A��:p����n��]���A_��:p�z��O����F�J�R�M[@C���g/��B�{n����v_
I�iӬ�c��n�)��h�t]�+߷�0�Ȑ'Nt�Χ�����	f�n�z��yx��@@/�Q�Nj�q�l��	j��^9c�������1GF3�j�	+X�����a���'n����^������aIf������g�6h�����9D�K�G6�յw5�I����,Q`�� <Ѐ�;�"ڷHR�g��^f��Uz�X��$ᮚ���i6��4�E�ާG>)�JF�Z���3U!f��a�}H�(H{�o]~�L�פ���z�8b��g�2���Y|u�9|�����M��/�?K�#�f���.K�LC(8������n�2VdG��F3I��R��s=_��d��l+�pp�zHy�c���cmW v�6���Ǹ쭭��o~tȯ8���� 2��B�����W*�8����꓂i��M�����һ���y'���(����fP(�Ϲ�.��5�5)�`�+]i� ��(d��S����lG(�X��@R���!��`-p)�a@�u
LT^�2O|��-D>|�n@�����jaq�kL���M�q�؛�m�Y#"�B-^����*�A���3h��-ᛑO���҄%���I�z8���vQl�ئG�92�
��ì��6������B�Qe(�_�;�V�yټ���pz���c�k��mk��&�Y�O�$���N�b�|DT��1�Ҝpܨ�������0|Ռ��J-(������p(�P	"36�s��et/A�#ձ|���0�>R�σ����97�²�Tq��L�����|���BJ.��f_�npK����g�^L�Ш1p��1��}Lė����Xٸ�c#/�U?�|/�f���:�P�<�!=�&2��xy:(v��o��t!��	�H�49��2��Ha��`j�2�9C���1�:�l��W��l�:�4'�D�������ܘ�����}H3���׌vO��b�G
�m�7&�0�QH�7��k�{iZNp���v>||�������(�L
�#t	���>���l����䁖̎�T��M��������\�a�1W|2i]gañDs��׽h��@�L������<�+�sV�7��x�!~�.cm<6��,�g�_��/����w�r�ػ�N�{ǽ�[Cym����z>m09�V����9~�_X�(��B����Wp��U$�/��� -���L,�=��Y����dB��d7A>�0��Axd]�������)��"��Cܽ_rʄ��w��:���#n4��a�g�!�{�A�3�h�Z���ʴ��{и梲�*{��n��D����{����ՃG�6>Eh�.S.J��c��5]A�&�z{�BW�(�~�_�iXO:��6�	��
�0[wӍ��Ͽ�"����B����M9e��k��繍�a����hfK�	g���>��r+���O� ��ǿ�sBx����S�Lk���n*x?(m����j>���d���U0��)x���Z7x��={�k��J\��V�xh_3�&��v�%������΁����x[�Յ��gۺ{�g�hL{��`u.���2Y+4����K�6���gńɏu/'5RM����լ� ZᲊI?���T�#�S���v�Zb�ɯ����zj��TK��8��Lc�8����9�*GO-E"�z/Z�GC�;��iY��"L�v4P{�iE	�./\�z_,ú�f�I�u�q-<7\'ZtE����28�.C�"f;���£2<�r\s����״R\���������#��h��Zet`I9�%6�����M�𓺉��Y.�4��4j�������%1B���� �G �b�8$�NI���޲��q�B���̝Lf��)N��C����z�n�UNj����(?��}������T*���FMhb<�M�譆J���|>����bB<
C4�t�Ӵ�:a.�~����V�@$\�,Ns����m��9��,�Ln��� �aai��6;Y�������j�u��	�tf/�k�,CMgM=�S�Q�=��"iXm\����:�U�w�R�M�t�Ƅ&�����2�ܶbz�S8$2RߌR��ی�6j�A3�p�xý"P�����.EL�
�G��V�h`���-�H�iF�WzX�Y� �6��^`u�����Z�)��2���A�62��_5Ia��4��^o���R�EYKSI���*c����M�=�0��< ��N�ҟ�.��&`�:MiA C�̍H�W��j堹y����D�얷�5�8�V-�潺���:��a������ut3�����c����c��pR�!����AU@,ϼ�!��6+N(��*U��_����>�ry��}f�2)]�=!�Mﮕ���Y|�`7�Y��9����Km�������:�7WwQS��X��vи�a��{$(�!��� Ty�c��&��_����/Q���HM�*����i���X�d�ܗW�(Cn�!�8�g�����}�,�]�z����2��I���nbܴ4i�o��z�8J�g�G�b����N��vX��4���b��O��C��]b!��FF�����]r$ɑ��{\���
�*���r8�v�����2�yCv7�PH��׺���Y$��9˙藝( 3w35UQQ,�����'~�<O*��S��M�t����͂w���e�m6�f%�O7>D��C�n"X���]���A�n�"3����Ŕ�a���`zʃ��Ʀsu�f�e6vai�ꀳ�̠ź(�3E���
�~
��q;Am�N�,�Հ��L<:�;+��%]ދ��Nl
n���0�,��A\\i��Y&[�SE��Y�b�{Bɿc�#� ~�� ~��r���VT�䍦�y�kŜ�W��j��}�6)M��>&�b��SVU��J�D�\���3k� +w�#�6��k>H����o�0m2/u��QY�-Y"�X���s� `�_�52�A=_�\S��U�c�]]Kg�5ȭY���k;��og�WB?�Ȭzƾt_d�W���&�V*J=S;�4̉
c�����?���v���{�;�Z��(�����Y���T�oN[�,�y��f*O�B�P�Q������C^`(]�OY>pE�`���"��f഍�e�O�"^+�{��H����u�}��hDl4����m�4�_�>U�v��j
Ȑ��	#����;�QH�8�ח)qY��@���.�1
����s
{N��B����r˚��O���/?�İ���Ҳ#�Q�_.T���/=���sP]�}���I�R�t1�d�FgA�V�/w�3PF�r3�Р4��cv���or��,
{�}&� �3u�oDo���Vl%s�f�����,�C��Uԉ��=~��М�*�\�&����f++E#t7d`��$Q;<��͑HL����5*��'~�g�=�'|�/�,K1SХ�ȴ��s�@�ڬv�s̸fk!>^~�x��<SjJ�a�ԝ�	���$�1��R�E����w9v�Pw�X��>;�(H��3�>�N/�R9����|����+�����P��"���!�~���O*�2�E�F��Y�k,�}t�Dit7K dR������m����������0dَ/�8o�������L�N��YE�����	k`40�Y@�! �|/���b�l��'L���s��1��b8`�O$��0GkX��S�o���.�k��ʪS.�C�%V�Y����I�D�� ��̟�����qA���Nѥ�쿼إR�5���$�F�g�T��u�e��T3�P:݈W��۷�۷�Rl��͏�|.4Q� ����$�e-��sc�ڤ�5��斮�s��YT?T�J�=}�Y�1+M4�N��**X�K�#��rۓ�3�|��*���`��yގ��;�O1k��]��!T]^�g�C�\]�(�׉�vo����}�N��:+N��R�tͰvW2�n��=�X�]���@%�Hkc�f�yRu�y�L4:��;�u*��~�'�Z|S���0<��ɦF�U8���jH�{��&q`x�2՟�pqȖ�0�-�o����Ϳp�/뒥I��5�T�̣J���q��@a����W6�~��G,_R��a�#(�W�s�Q���n|�7�ƅ;%�0T� ;?�y��rsL��Ԍ��Κ�����c�ۂ%����_�o⯃W�����5���Ҵ,F�1��`zX�54���֭*�p��������mU���`�8L�y�-��z��!���d���c� %�[��G���@~Q��|n��L��P���ݧ�xm�|�� {Kv�`\�M0p�h�In�U� 5L�=�q6	�t�2t�Н��m�4���15�x���2�U�3��8G&���wXJ]��w�y*�u����̤Bj�s�w+���Z��\·���`��FC�"9ʰc2�����uu|ׁ��P'��0�z�������{��9���<�*�%�g���É�����h.�$�@�i[�b�? EɄ`�E�@�����LQ�+}ɊO�QV�uqs/դ�ۮ�*�*9=K�R��r�$���*~�L�����������	&�d�%7E8b2���z�εs�1�9J�q��{J�q�;�u�$ h૯^�Nde(��x�S�FՇh@���� ��J0��ǁ�<ӲbV%�0�m�m�����kq�]UWJ{�NՃp�"����Q��#��y�0*���B�'뚕��Hp]�������m8��C|u���c�����^Q�����nQ��z�4�@�m3��Sgy�
�;��D9�a�ґz�DV�&���5&q_�;��-;�Tq�R���b��e�.���Jdanژ��L����ו���}����B��������*�KŴ�k�&c��q	��+U4�Ү�U��e�`�y����6���&����6S�oÅ[p�\f�͡��J
��a��hfou�1.�S3�.\P-��5�L�F�Qj�^��app�4P�q�e�#X(�f%L�x���a��L�P�V�u'p]k�~���i�0��[|]lB�~��w�сq����+ΰ�X)�pS������m��S{�
�����d��SO���E��O��9m��Y�������llt��Gܘ�-c�l$�1��<f�!:܋c꾣=��>߅�SnԶ	Q�+aY�Xb�ŕ�>G%�r����
JP?|�gգf��َ�I�u��v��[0�9�sz��p��(VUs�&pe@OB���,at���v)�d��ş[EGwMA8��ȴtؾ̃p���-Ȇ�-����)�°�M�C|g�`HZad�K���d�Jr�m�U ��h_�@6��Ftݷ�E����8�:##��	�̮�nD��U1L��ؕ$hr	��
i����'=�px������C��:�-ʄ�����3N�=�l����Aj�i��ZXHk��C���RͯL��&�s��Z^	S���0�o���J�o߽Uix���s�6,�i&x_]}��>3R��)�Zx���*#�Fj6�i���:4m{ܷ߼�'�?��?��a����'��'~��oۦ��ӧ '�$��=�ŀ�fVt5�i�`�2�e���w��wߕ������g�Pa����Z��c{e!|�?[���EKY�0_���%!0&�L���e���4�+<�|�8Z�"6���5�WF���)�ߐ�撟K���a���/����q���P��}Í}G;�;��]�>��6t��h-�@������|���1�k�i���챌ƩrY���}�����sY�w1��EsP�i)�?ex�A ��vH ��sb��H#˴r?^��̽hyd�\�rB����8�����9Y��ڜHE�=k)Ⱥ����r_�>�_M =�w*��^^��mP����U�?3ԦW�9�Oo��D1���R��_��?��*�*��W�hf�����|�8E�f<��S��%*��S �{	n�4 �������F m�����~@߼�E���U����"H�b$?2�͍��NT���6�\E�l�yьS���}TS���q���9�6o��9�8�0�1�S�p$��0�υ�:�8�lI��;b�k6"����}X"k0�V�����f��{&�a/�k\}����9-*w���
9��$\��Z	�s���2Mi����˟C��/巏����K�n?���G�����F�g��4��{ҾUT��\�`���~�¸��
�Y,XYe�Y������R;��X��C~�&

 �@��@�osp�mRfI�]M��Z�\�UW&�k��TkҬ���^9��l��4��_�=��gi�Ms(#D��d#0����Y�-�ݯi�`rc�����1CĮV��=�������2{�f���Y<���%6X	\�	��a��Z���.��w��w�����ђ�
�<KL���Ҝ|���u�V������XJdbKr��3}u�4^d~�	� �+k��G%CNu�Bxn�)�#H�<�d3Ɂ��#�J���8g��x��/5oN9��6'y��$�e���va�w�9�]s��<$���Ķ���H��P��>�	¤�r�����B���m.&ܗ��M<��|���M����Q	�P�z:�Z������� �Q�=6����MnX]���Qy/L�\Jd�yH�5Ƌ��E3c1���6���p�>�A��b`/p�>)��A�+?��.���\<�7�2ј�{�?Z�8A��p����e�{z���Q�2x���,TYf���)�)�e�
9�D��4<@���`��	�f�H�WZ��j���J�1�����A���Q4���j�ղ�^ex����d)�_Χ[�ߗ��ɬXG��U�1�}�@�`�}}�&��S�|�gO�ipg�-@���@�N�������Z�a��n��>V��x�<[�,(
}��5�s��/WV~��1;;�ݠAYL��(�)�1�hc}�N�m��,c�ͥ���I�d�k��bmH�}�A��ӻ*9�Ċ�Nu�_�2�\=(ܙB2{)ҟ�{b�6ⳌX�3�'����w�6ǭ��?���CI~�j\X��iPcm��x���5@P{����iul?Tzת9n0�m��?���y�]엟%N�)�7��(�RW�&���|��4�&���a���e�� x3��~��Z8.2h�]��]�aߗ���4���F�~	��1�o6B�	���<�1�UJT|9���s�.4V[�ԣ�]TE6��A�n?�,��:�0c�؃l��(����.�;/�AaӏݣDZµ��}�u "|3� �B9lB�=�����H�Q��V�����u��s�U����u(�A�jzw}���������jdm��2˒A��h�Ԍ��{���-rRG�E]ES8���:����a�(e)�N��P<�CԀYD�y\%&��/Vy�ȈQ>,d82�[�%�1�fN9;�@z8�W'����3j��l}�y.�Jji��4���u[�R�77G�kjA���k.���&*w�Dtl����&�w��x�,�����#P��P���H�Rq�Qdof��<1��uf��6�yd�B��m���b�	ҰV�(��˿������|��Q8�OY���`ĳ�w�BAp���D��9IRmb@||T3����]p��bM���4y��I��a ����)�a��ӓ �K4Q��/��n� =Ji��1���o�^���{|ޢ�D��tp�j��ʹ�E=���\�j:o����jU2��.�;5&�]�xo�'�U^�j�-M���F0�
Xe�N���u��nV����jE��$��H�_��.�#⿯����U��73R<O�����:�F��'�`	>}��rIc��]���B�������٥�5�>sT-d`�
l����y�{j��.aUw1&J<��F��Y�d�}\��,!8�M Sm���k��g~����x}�JB\�;�qL_�����Z����2%�'	b�	�&�*M�\��rtq�in*�%\�X���J�Q�\aB_�5�ΕɲY+,7����ǘdy|�ͿN�Z(YZ��Izۯ��/��*��/�J�;1<�>�a;��������m���샎�GeM^mMO�!�y�
6y�lҎ��Zƃ�b[���p ��ݻ�Y?�&��l8�;۫!���5�A����_�� DV��tf��|W��]��ޮ��/c��"�d_��͒{{MU`%'���ǡV��4s"g�]ҏ���ág���2���R��՞�[EU���kl���m�3M��|i~�k��RI�J	�xOIHD�Z7x��$���~}tW~V��7�8�^�^����&�6���a!�>�t*����i#��S��b��O4�7KS�� eQW�!S���������_���Ngv�倫�[#�`�h��o��J��S�$l�_�p���n0�c�0�S.QYV�� b�n(3�([Ks��1���86�m-���%���LY��ڔ��΃��D�eXɠ[�-��=�g& & �h#���NZ.�1Qt���ŽBP���L�������O���筤W#�xv�A�T���f���(zJz��S4w�@ uy�������b~'���S���n=p�A����*2��ۗ$���p��ÇP�*ѐ���N��H�@:���D}e����/�<�*�U�n��֜l5tG]�]'�>�T��EE ��C�Oc��ޑy.���$~��@��Z��@_�ރۛ�7K��6��X*q��	��x����g؍�y��49�Lׁ�ҴL��1PW����9Ú�C��^��
��t���8S�xq�5�e��B�k���kDF�i�{�O<Vb��ɵ{�R�H��K��ݐ�G�(��;̉��Ϯ�'p��X�w�Vz�馌iS�.3R�[<��m�
��gn&�~A����>tQ)N����@>G�9)2�������J{lLa|�E��zJ�C6[dC0I�%Iٚ]�Ӂ�V���<;�ȄrI(��k�*.YV�w<G��ؠ,�3#�F�������?�ݲ���.��4���-(���	-�'f��Z���@��O�JWz�V$����\�F6,��)�.��n'��DPΩ{������'�������}���t�H(4f�܋��i2���@!��*2WR�愸���a��jR:������xb�lF/���T��r��S�5FUoȍE/����.�!?dS�t5����eL�n�}�����������Yk-�?�p
ރ�JV����/�w�ޅt�%t[�!�T���Ͳ\�	���(����/��x��@<�0Q��:�^C,�P�c�-FZ�JPg�Y�!3X�+?v�W�/ty��	=��N!�[�u��͇]t������"5!N@]�]]� ���cF��w�������e]�kԲv��g =�n1қ[b��%��\F�'F 5V�C����9bxP	C��̓��%n��5`|#�=!{
1pY���Kg�5��]����W��n�ajT]�ՙt�������X���Ǟ��B��[&UL�E��,w����?3�y�f��ھ�u�㩻�i���n�}����9�<�Yb ��8p��2(~�	zM��Z
�Ja���
���:��\�g�X~���b��_}���^�Za@�\���7~G�����9��б�Mk��z��*q��ԇ��Jި)���Ͻ׉mOUp���\b������S�-TF�['�RMB����̨�\;�����R��?�q�ӆ��2/�0`�s3Q�����d3��PKƷ�;q�M4�Wz�]�S��d�5t�򺏓G�Y�׾U�7�~��I:���%)No͕+�00WˠSS	���s����áR���w�@�a�s�{�9��L��xt����#���tִU�y�Q4���K���$��R5��8� �SO�Y�SB��ϸ��:B��*�/����2W�-;��jW�,���l\K9�>0��xX�/��*�Hl�����<=^¡u_.5(v���m:�M:���AX��HC���o>�&���0Bl���O%6'���!D �P|�Fm�L��9����>��W�_�y���E���.ɷ��=ƙ�
h�"HB�?�^����M�k��$�� ԇ-�Z��Kt�`2�9�6q(�}�<�x�N���m�a������E����1H�?���T�|W&Kp6�>esNr�C��FJ٢&�����1�l�Dy}a��\p�����>�v�6̂�_��l�?��W�P3S�t��-�Pi������H���*.fRy���i۶_k�i]�Id��>|�'o���|߇c���.���]}�N�o�4;�$�K�\���d)Ԍ��	���5h���1�Z��8�iU��K,��m���,>�5s-F�Z�a�ټx!�%9k�q�]�=9�0��,X;�$��EF��/1��;�����-K`T(	{�AW��)f��k���� !?��^Kf>Ź��S�T҃��)@%j<�$9w��,�b4"�s��lΡ�������w���0��?�(���=+�q���Fe�1w��W[���¸��ޱ����*�:q��G:ǄW�Ȃ9c�˯œm�,�gN�!�d8ĸ��M~:�����v���'ѷ[PG@���
�{f�m �J�!���)��\�8�8D<�[{�k�˩�= p�z�6����@�πr^J��b?_����Ͳ�.�(N�H����y^��IH�c�N���K������%�a��=��	ASN< �>gbe������Á���ki� CPL�����gZ��u���gy�#]�����ȃ�g����eW�AjF�{�h�W7��C*�*�&�K6�y�E[R'ؙ�1�|�t�7��s��'���F����%ʺ��|�^������6>F/�m���{�������#mT��)F�uʌT*T���矸�+޾�}�n���Y08N	vBW����X��V͌��y���`N�))��-�9��߅t������� ��Q�q�`�̔���A/�y=q�p�_o䙆u���!�A
�9��*��#�)k}�w�3 �H͜�)��Y���w��kS��1?�d��8[[���8��Dy��W�_DP�WE0F�����Ge�����/&�N�����&O��������`��+
��:�f�Z8ݨ���b��D���d���S���^�$���4S_�yw��������,�b��)�Y�x~J>�W�a��	��'�I�H\p���)L��Q��9�x�~)V���� �-۟$t� �tb������Z��`��XӿJ���'���Qz!�*8mV�S*NOy������I�T�A���a�b����Ooys넻�}�l�"7��%���[##n�Ag�&�㔂d�g�=����H�7A�3w��ж8��NK�mG�
��%���ڞ_�"ޏj��ı'�5���nn3@Æb]�A��P��خB*���S?����k�Y��C���Þ�8��yW�/5#+a�{�����u*;�UP�J%��>����?�#34�~�����&�?�;��9�h�⿱�����IQ��DQm�Ϝ����۷Qb�x��i�}6x��y�ÎU��~N&�����x�߽{�l��\4�°�Cs���'Zd�3��ɦp�<�Εn���
�2=ixq `��ݮ'��J+x:H�����l&��qU�e�Y��@������hX%�������r�=���,LL\w��l�Y��n���Y�h]���X�vϐ��]��넱��[���σl�+<R�,��b�����'�ˋ�S-cfj.c�-!�'E��OUO'����>;i��N8'��A����HE%Ѣ��s�3���;�v���ob�ׄ+�g��B��'�;e��&ӳ�c��v,�n����=3ҋ|���|XGKX���Jɛp{����^7������C�t^�zC)_t7�U�;$&���gO��i�5�)�$O����#��,3l�GG��`������(�Ⱦ��8(��Ǉ;� �Y����]��"����/�=܏{�b�Ǹ磈��~��������-֬��oY�#CE 7����P=�(�5���.e��bM�bX\c��$���C̦+ F������ .!kc���5Ք�>���ܥ���u���A�����!�c�<º�r���gT�Դ=Z;c��k��]4��;Y�L�H���!��Ӱ��Cb�OOUO����~ga��A?��qSȰ�n�ȫ�+�H���c��j��6����M����vב�Y���fSl)��+G�h6��d�%��&���꺨�y�Jv)%ʩ.|i�7@ٸwv�������� {|��
�9M���;[�bX�m�{�u4�v�	��D�g�wp�MG�_���k|��?��?�	<�\;d��L�,�xf�C��iqSOAZn2Rw~�gzN�MQ��AT"f����n��X-0�x8��l��f��h�Ǜ<�k�?�u=�۱����_P�z,�Gr�m��.Kt��u
�\�2���`J�Z���]���ZwP2n�.88~��G�z�l=+�o�޲�o���=�3d�*E������?F(�fd��k�A��3����U��?��O���%5ǁ�E��z�e�G2�ސ�"��'�<]�L0#��L�%��Ԃ.�\3R�.��--ŵP��\��:�}�@���cc�h0���>ǐ����P��-��㣦��]϶�ց�dÅM��;n�K�.'��:��wŕ�S,%�t�m��U�q*���E0~jL��s[�����������oF�����H� Z�e���9�~A�j:�J}�RԦ����xB�"�SӐm�FbN���58eh+�ݒ7�?�M�<��Ǭ~���^R��(�J8R����g���#m����62 ��92x6G��TƂD��ݜv�����7��y�&�����~6/@Cn�`q�~%�K�Ҽnk��*�i'��@�Q:,�� Z
7�n; �}�K*�)�51�L��#���g5
Un.*�)���t���q��n���?x"e�qQu�q|���:��`4���|U���P�#�}�M,6*Hњ��!&��y/�F�m�O$:��\�:�7���8����ϗ'fy�`��������Exء����c�&����4�LO�\4��߅��3E���6j�c��6Dڧ��8JZ�wY��K\23�H2,{�5�Xdw�ߗ��������DNK���]�o7����������.&��p���R!:��+Ҷ�h�t���:���!���
���䥝�kjۻh1�/2�6�u�[�c�䳙Zp�T���>�Uc�ւ�Ԉy�%�<4�}v�G��RC��h\~��>2��cz�.x��Ң����R�Bɰ"�����c{ &��\R��e���Y&�V�����X��\� �2��ڜ�d���������Y�����_KS'{f�/ev��@�_HN�$��eu3N�1�nw�a���.lc�q�񿔌+O�5u�Р��w���_��9BX��y��gW���Zb).�/;`�><q>����������7�8d�@½�Ͱ����o޲�|p��\��JM�c4"���-��@������A�+Q��X�Ct{�l�\_H���<Q��ٵ��!E{%��9��5�Ws4�P��=�����0N��l%�w� ��b���V�/圛}Y+��,O���4ɇ���	G$)L$�J����3nՅ��\�� ���1q�qʽZ�1j %�wx��X�Ɗ��&�@&̋b�V�r����m ��d)��P�U(��tK��u ��~�]2\��iҸ��������	��i�_�-�k�{�0w���@�2b��齻�%�p4Z���!�Cl�9&5��1g�����RK4y�UӴ�g^���.�-��p���kf@����s#�A'
Eh���m,k
���tj��*o#�����O�>0K�H$6:�&ў �:mL�d��K�m�S���z
���k�`Gn�������;3�Ȇ.Y?{%t}�h��bi	�텙�2сYX��i��r��F�����Y^1��k��w��A��L�������4�/�����
m>�4��Y�;�����m=>U���&�����̵`��=f�_���l"��E5���R�������o����r۱���dY̡��� >� �� ��wwK��?�q �ґ������'��Y])Y�e�bZ�9����A��:���,S[f�z�XlȢ!��zU���z ��)x0���j���{ux0�K�=�RO$�C��vekTF�0O�>n�{"�{��.�_�?�8�hZ3R_/<���646�p�3�ps1��Tlb�����D��4�Y\_m=x*��ҴC�!�7���T���,Qm������<� ����|�L���c�`K%��O�����P7G97�"C	��~����?���/Rf������1�����=���?�q"̘�/^�����_�;�5Gb��0�U�x�Y���X�Os����:N�S4�� ��`w.e���J�!�0�`_(�EFP��J�� K�)޲�`�A��.W�E�5�?7��yAWU�n�5� p�!+7fV������ՐqUÌ��Fx������(P<]���U��`���H7�ͮLHB� �����/Yv�ٲcg�]c�fXf	�^qܻ[6��UG`W���j�Ah��I���^1��ɧiv�X���S�3\-٪��F���Y��Lr��\����C^/Q�
��g�^4�A.5���U�����`�k��Ʃ��W��j,�7U˕t�4�0ph�w�l��re,�v���>W�������]��R$����HG�bA��X"�X w�ҥ��q�� *�@�f��wƁ�T���I����0'��[yG��z�@�3�ee#��:�7��<���>>�JP���ŮK��NڟbZ��vM����[��k�ܮ�;�jb]`�A}��"���6��湌��p�KN�`����w�H�>0��j��1,��#���FԐ�/]bU��BUΣ����~_e�8	�=R<B�ͷ�M��1&*amb�8�&�7c�i��T�����HqN��[9xn�83�\{?;Xj�W/�O�>l��m��5�N�3�]�Q��r$U�1��O�������9L�.���\���J����\��D�j�!e�'M�ʹ�"���kjةkbI�E��)��9�6Y�Z���k! ����N��*>����]Q�i�I�����I��J�(t�.�{��Hi�a����n�������Z����k�Ef�,V�U�&��ϐ2�h�Q5�Z�e�v� +XI���/XG��<�;��Nx������C�� -$��B����'
�;<I�'�ҽ"Fy�g�� 
�lvU4-����ޅ�L�����:_�$�&�k<!Ȗ5G
�ѺyDrs�����[H[Qi2&"�8p=�Z\1!��K��������%^<�b*
�q3���ʄܙ�
@C�pBuH����&iDM�A�D��I��>~T�&�9��V��Ÿ�SQR�B�ㆠ6A�h�����a�� \s�r�MC�mБ��0`
x훯ި���60�C� ��?Q��#e��g2L4�Zb$Yx�'�&���et7����#��jm�Z�G�O�'�N1z#�l0"ၘ�K����O���KZgҶ���goz��l�s�g��s-��5���$�75�w�>� M.���� �am ����NA<-�Ԩ�Z��zb���.E[�������Wx�|ք��
Ho����[v1�q��gbq�ͱA4�x6����Z�4�Zn8��(�MĽ,MW�^'砣lr`#���s�x�����d��j.�x���:�D�b~:������e�@�Ȏ�[��̆��.��7 X�r�7��Q
H(���Ԍ��@
���Nie=�Hi��W3�+��xщ]�:���Y�aWr�3#-�tX��kjQ
��'�aps�s&��[��>^h�@\K�["p��BF��O<^�Щ��mc���4n�>gR��yQ�!&\�����GF���ÿQd�f�����o�|�ꛯx ��NC
2��X3�Q!T��<��*��}IȬ��<*Hh,��a�Z�k�(�Y������G6������2���w�����U�{%8}��q臄�j��N6՞��$��25Mr�AW��LנT��ǫ:�u �D5�����J_�FH_z��H�>[}�}�&ED��R�?�W#�k��Ԗg�̤68�����g���د�H�PEa{u��>Lhr@�6��c]��щ�,6�Z��I�8le���54���|B� z���9T��A~R�u��^�(�ڟ�aQދ%YW"�U���x<���e6w[��+?�224[���n+���x޲���Y��Gt�?*���u�'��q����ڂ���}��Y�y�x�%b��>�9�	xs���p�Qa����l|,�-X|���m���N��Z*��香�l��y����׻��vd铦�X�`�gV���q�Yr|֧U�K�iɔ`��tʵb�̤��~u��Rkfd��(��N���i��_�T�?o�q�NA	Z��#�ȶ��s��a���@,��_ʿ��^�y\�-c���^�ం��=�C>n7��%��!,u��ތ�*��Wt¬)���uS��Z#!����9q�I�����:e��pMq��u��[�"�B�0�P4�;P�!���!ǟ#�;Ӝ�w��X<���Ont������.��%2Y\O�������TT	�l�y?;�/�~<vy-9p��k��p���9�]}���2�8K�A��&�H|��K׽�u +�Ⱦ$6c@Z�ɒ����5,�w#�S47��n6q��H�6N�%AzƖe=n�g�$����h��dC�~x��m�R���!N���
�w[ ݽ߂aP�>�߅���)O���)����N��T���qVQ@@�������[����ɱ��R|]`��H&���ö ���X��N��@=
l.YU]9r�Z��-�Dp�t'��8)㇀���P��-uՔ���/&��a�;pS��&�d�|�C�vp� ��᧟���K�j�ڞP˸����3_	�t%Љ�5�o	���a�fo�z������	���D0�t��q,�?=�~�5iEaC
����_�l����^�|�d>}*�sj��YSm��m��2N|�*đs����e�U��C��q]BT��}B<H��k�L���2�9yv����g����qv>�<������z�!yp�����1A�Oqv��~_��T�':�GOAI���@���X�
`/(�C܈Xꨯ94t����D�2ϳҒ�+���6��	lȿt��(U��`o��>�x���R���|>޶�s���q�⍭w8�p�/,��M��H_�E� x@���k��X���-|���cQ�̞i��ʹ�`NEm�D���R��;D���莛ma@_˧�ч��,)�)��j0������Rw+A�Ң���j����(N�������������w����#x��?�5���m���I?m��@�2O5<+�u��C�XJtL5^jq�\;fp>؞�i�í#���Dռ�$�(�T8ѵ���ϳ����&׶���	��W�x�2���,����4#M7���Tl^��Rv�ʙ-��]\[T(�@z)�����0���H1�
�j���!�MŒ�#;vT�u�H�x�+�e� ��5�L��v?\g$��ll�|��DxP��2� l����C֟����2�SfMID���Su7�p�M//���"���ce��EC�ң,e c<���7������E��]c�S��p8x�	�YO�]�$�9�:Zw��tO�ߠ������J����E��9s�e��I��|L[�uI.�50�n҉6ש�>h� *Kx�H[��Bn���:6X�
57~f��[�!���	7��K���%�޿���C��1�b؇��:�L��E2��(B�3�H�er&[���TT�?`Jf*���G/ �k.��Os�ۦ�~G�Ydu)܏����ۭD<޲��������_��� �F��$ħ���I0���&�>@��9�DֺӔӶ���'fF�(�2�ǘ�Z��|<�����Ĝ�x� d�qؾ�ɒ�Ko\�����G@����>o��->Rĺ� Zm�H;�ñ&X��9�!F��ȂD��/<��[��  ��� +͇�3�]���0F�"������ן�����՛a������EԵ]^��cW>�W�ŋ�+y�77/#�^�<L�h%��2.�΂L*�х���@d��5a��x���X9=���ӂB��2���-@Mg���%)�!& z�|�f�nL���P�,�>��wC	ח�_$8�#�}xM~�3�f�@!�ZE:�%� ]V/�<�O�z�UXm���sZH��v�lܐ Y�1XSs�>�fB`� � M����"�n��M�h��t�b�5�c]3�ﭚ	?�	���_�s"(Y�v�:9e��dv�"|s�Xoד�>���@�ɩ)Z�xm0��(��Ϟb¢���=) "{?���D��b��r�t�N�gf9�4�1=�lE���E�݊�;m�i
+� NC�n?�D�?�4�p/����t^F~NO�A�L��������`zn��(+�~��M����&&��x�ߧC'�9����隳d�.O�,	]�"@ޜ���&�w�}���l�� ��=�$ӷd�C�uRݿgsO��S>�br�I�ٴ���+���N0�c�Y7�| �2s�z���%J�h<�5��bt�5V,x$�/�c��3CU�t_3�uۙ��B��9��f���5:��t�aT���KmƐ�+]�ur��W���{9̊t��nS�H��r��Օ+=�K�#�p�������?�����?���h��
d?��83=i��#8�{77����5���B=���f�r��r�֘XZ��AX�^-MѬ)���2i�(բH!�TXSu.��Z�!:�5SO�FN��Cp���d2�W��]J�����æ��EM����$'HdH���>PY�$�gP���\������(�U8��E#O��
R��6�E�q:\"��R�B��0��-4Q�cO* MXg�e��qrR��s�g�f���\�jaоo�:ݔr�M�.��d�FE��9�q	,� N��/؁G#�7_�w�9~4���Θ<�M29<q:��q��	�h���/^�{��%�ws_get%�N�~���b�HM�5TWf�h83¸�&�j���=�7�p��J@7����*y^�0�*	�5\�q��Ͷ��C��]6|,�"�ʧ���'E��i'��@z��q�_�C	�⪒̼�ꛬi;����Q�N�\�����K1�fS[���	�]�X] ������V��7�\��Z��+���e5�)�>"#�M8�i{
���h�3��3 -q���"
N�@���I�����>�A��3�)�E<�x2+�ʥd�'��Ճe��e�o�dse5�vΛ�� C�5}f}S���9�}�X�+62Jdr
{��"��1�ى�=>e =�8FE@�]6-��W���Q���i��sHd%J���9�@�#�8v1\BukM؃ԣ�hZ��?�x?��k��k����T��!�G}8��I'�- ����gd�>`�׾d�.�-�����3=��"�ӖcV��SP�����ٲ�O��X ����2E�}U����4��N][X��-s��c$遶������XQ�-s&.��b�I���lѦ<-��>wj:EO @�FCy����'e�_]�NF��ɴ�#���F�ā�
�=��5�T��03<$��~a�#c�Z�J�On6>f (�9�G����}f��iFZ�F۵X�e-V��	gz�3��:`���7m�'�\���J�X���ol�Wߡ9kjfMk ��yb��X�4'H���7=�[���?M�ȧ[ٰ*0�a�l!���L�qWҦ��ʉ��}�SbKƎ}�׸�iԗyȊa
:~���}�}V@��s�җ�}�D5s=ĽH#�Q[�0SZ�:R��l���t�w��1�K��������44��:�4��a%��u�{"fU�����-mL�$���9� �4!���sd�͖e�c��Hć=��'�)TD�f �
Vj�S��"!��k6dS��	Kb�����p��l���'�4�x8&%)��W\3@��3|��s�y���M4m�����K�y<���J�L����*.
����y�7�!���5�`b�}�s'f���4���L��ji�'u%'i3��rZ뺣�%F3Ą�i&��U�k��.�6氱�9�<�h6�X�� ���Z'O[@]�!Q7jMha�q�Z�hAz)�saFSG�9-�U�JfP�n|��s��;���)k�V�� ��Z28U {������Z�'S��M`n9��"s��K)���'��L
Ze�K�1��_rI�s\�g�JO0�F�t�C,�����E�;�6m_�x��W��ݓ�� u��r�I&	��0XC�c�k��j߰Y�I��:�dR�m��~#���T-5V��V�S�&>��2Ppr1�e+���v,�jg�bjq�Ptإ�-K���'�%j��Y���?����� ��H5�S�-����9j����縇��;������K�ks]#��f�٤E
ρ� �W��s�&v�'��vR��=�(1�'�)�X���DK}A_��z��K�8�������i�2˝�c�儀��1&��ɇ�U��'Mu�A�r[˜6�Sd��9KM4N�@A�8�����]��}R���5mhhx�mG�D��fJNZD3�MM��I`���a����Ű,~X�g����p����Q)��E��VҲL)�/p��R���g�e��rZ��i��%7��Z�!���Θ<Q?E�Z�,1��N�92��}����49��%1䔶�2F*o3�w�_J��Z��(S�z�&bm����&�Fo��c^3z<�F�8�P�b��� O(`�
�~B'���ǧ�3r��z�xmu�OU��)50L�=e��<�4�������M�l�=��g���f#-�;'�nd��$�������L�,���V8��"��Qe�تy��&��:ց�8ܽ·UU�9�W����6=��{=�*����ʤ�M�P�g �����ߤ� ���� g���Z��NF�������e~�j����`��Y�;NS�Kć �ٸPy�E�#��>���.������x:�G��%�cuB���O�3g�T��5��x�$i�ɒ�*~岕���.$���}�U�d9��.��v��5�σLbV*�sd��F�=��(���F�G<�pI3n���i��P@��i5���|�<����s�
��B�ťi6�r�����~�s��]x�nn�<dOG�:݇o7�=���%3IP�\>�%"vAW�E>�8��G�y��>�Y�D>��0�����8��ۥ��dmM�> �Q�����lin�ԇ(	N�=�í5�&Ɛ��3�լL���q�d����n�fn�����r�����1U�TB�K���P�ܼ�Qҡ��k�	����Jg�������,[�{����3_<�%��}W����f�_mE��_�塹��	TU�������@��q��ε�9J}���p�ׁ_�PGO��YYEw�*�E0�{�f��V�qP�+J�ژ�n�A�U�#:��5��O����eY8��Lh��A_�YY�{I���U�ɧ6����k3d����\����R�\Y���eA`���9��$v7�6->��Vڛ]'u����p�<�L��O�gX�Δ���3_���ǢY��ǧz >��r����P6�.#;�n:��p�G�X�}Y0�ٰ�� �;�9�!����M�{��	�5�^����{��KP�4ذfl�X	G9=��wIu�W(�ә��}��k��k��ϒQ�ĵDv���׵�0���Bɫ\ݸZ�r����6���:SK�Wَ�������Ď�W����.���$|�wS}8@���`zTl�������}���k_+�z�\$_�=A�?��J]h���Hɝ�8�K<l�Y�F$O�<�|13Y�,��Zl �;�<M/cH�B[�0�gw����ύ� YLy8�&1f6�2�����zfxnN�AwB������=��/}<?�4QIk�y��M}�jU����� ����k)�LY���5��C�=f�bgR��V��+�clof��6۵ZF�?��E�1B.����N|�)�<fH�梎��)#�H�����pfe���穝	���	��	�17�����G*3i�*���߇�m����A<�����EXvۀ��X�����f���@�uOQ�h,W';Ձ�	vəxJ��i�^jZkc-D�Ԩ�}�i��J���%�ֶ�v���i��3MO���~�ld9��a�s_��P=>t��Y�|��.��%���CQ��U���¤�����)�G[$�	GEvR�=��+���uio|��J3]�]�]�6t�`N�y��M���
�?74ok��{ ��tY���B'z������� ��1!%r�>ħ=���A�t�C �#��U>f�2<�KdȘ���,J@�,��l?�ot����k�l��*���r��%����NϸWV���!q����(���y��טl�^�v�Ye������>ph�,�)2�%8�]Y-*3����Ů�������Ԅ�ի0�������&Gm��b� Ȫ3�6zS��oYM��j�C������_��0\I����N�Dؤ6���]�.JUi������n��BhИlK4��[�I���V4��C� \b�4��?Ԅ _j-_R����A�>���@[�5��:�l9˞�P�j�WMX�}�1+V/V�#�d�X��Ka��s־��ݖ�3T�'�M0�v�M۶B����#�q���xW7��¶�+e�)��*�0� ���֫���2y���������]͂����D냇_�J2A-���,�m�[-�K��3�j���d���ǃpB�X��j��t>D�%�V:��趒/�������hq$\ �����7E����}~^ә̭�#>CR�b�RR��9S
,cZi]����R��|�ʎ������v�<Dy7g�J�M/�P�Cո�jI�efoq�'�������k�K���4�����
㸡�MD<=���p}���^
)GS9�$�0��-s��v?(��y�3޻���u��u�:�QE��>��މ��_}�-� bx�c�^U�����}��~��0���z���]r}Ծ�*%6tfYό�N!���Ῥ�G<A_ժM��9��Rg�]�@[R{�#�M���o���Ȁ[G��uļ�|����_	�>b�k�v����]���/����,I�U����!���.!/ɻ��J_r1�B��D��\��˚KW�IS*͸%-����&,�D�s�'n���'���������	Y|�SY�3d����0^��rNK�1���U/�r���!��ԃ�ŲZORAx�Ćp4d[��b��e:ܠ�̾�5M�}@�Ϗ9��Nr�@��D�K[���r��������m�/�8�u�����B���Xw�|\GAYR��g暍�׷������	}���"&���u�bYj���7��u{����E)N�aTB��ԻKd�,�k�6)K���t������ͳ��W��>���b�`B�����E�64w�������h����:I���96w1s�1_k�2�ѝb]��3�c?�g]	qo��$*�)�k������9� �áB��T'��]�d���o��m�z���5�����ia<�&��{R��\��]i�9K�dG�Tu�&��}���ܲ�OL��O�!�(;�]�V���s�3�w���RZh�A�xblj���	�X\H�����u�=-�DFl��$2 �1/S�/�w�U��>��J,a;�5}m���� �2�HoU�S��^�fzs
��'m�ؔ>L<�:E����-k8���_�	!�Zm��i��RS�T���P�����\ތTqz�r{/�1�RLZCńT�yy�Li0y��`��^�d�̴;Q����������.���(��99���uB��]�]��a���=BKȸ�%��̆��W�⽒n��Ur�����j�%0쒓b��y�f~�/޼����r�:��V�A!>�0�u[��|�,J2��K(�h�l�
XKf��{�qR��>z
�5�m�p���K�i��nxpd�Ԭ׬4��l9��j�jicbf���h��=�O��&H;Sb"��f��N0]-�q̍��5fܿ(��]Z����xӱ9�Z�d�!�ۜ̉�6$������w�T�P*��vpq��H��>��.����f�ѕ�	��U�.H�u�b�&���Q�n�&S�t��jM=Jd$K4����v�y��)p*<;�������k4{�m�)�'l�I��-~J���+�4��ih#�C�٫;�r������};G9�gp���¤`�k^)�O���tX��<�mY��8(\�\?���LR��B�ʴ�c<W��x�0De������ݾX��)�us�9,G��@�;�@@�ä�5��^�w��F]"�-���*V鵚ڿ����<8��߯߼���*�h��9�u�V}�p͊��`���VL5�]�dB���b�7]��$�,
�AKt��&dP����*FЧm/��ST��.Ka�w��/�/1u���w_���`�ą�w�N�����f��Q�57��ڻ)���)�o>a�G��Q�k�%B	_�Ǉ��ࢻ<��t�!�10���I�'�I�yM2:~�X�(ݠ�'9��2�~1S��F��A ���t͝C��l�����Ѷ,��t��#8B��WF�$���%�gջ(e�	B��MBt4�(��w	�ēG���,�!7+���z���Gv�/�bz��H�ЁF� ����G�mf��OA/k~�קXg�43v���Eb���ٗ��<��pn<_��$�9�ֵ��.���{�f�QƂn*�R�j8���i�N�����o4֦ ��kc �O�W�l��֒��	��Ӏr��9�~�����S��& W��ǚ�A��3�e��T��8x��Vy����D4}hǚ��@���cp���7Z�8R��Y6��=9��!��-��#�mf�\���IQz���Y����Ӈ����kR_�><ijI��g6�@�W����'�T�<��U�>X�2���2����;��}0�_�����ge���>�o�V/p�T�������ЂK�+_���`L&c�&����A�1�'_kOf��'Uo�J+�����;�����2�nw�Oܩ\�"H����O�����B@Ĥ�
��NZ�}t��Hh(F*�'ٶ|���@T%�箛�x�����\tW�H�1�,��u����K��9�r����6qKr;}oDn_�=q�@:Q�ڢӮ@q��g������C�ϐ�l���
l�Ֆ��֙h,� ^9G	}I|�4��,3s 9�j"�z�e5����C�[�W{�n�z�J&H<\|_�z0�����}��R	m�&0`���:�:L�Fa#����w�ԋ3��"��ր?�����}�f�4�SӮ�{��.�}Z��4�M����n�UV�V�u���cy��W?����׆x&,&�'��uA�ơ�c�ׇ�ϴ1������͢��.;���:���HCFjf6Q��>]$�[S9��B��t:���ۖ2���;20�|����R3���6��K�����܎�w��c�\�i6L�>��,T-� 㮕�"�x���Fx�]����,r��p32#��)|���s�U�EӪ����(	�-g��[3��Ȱ���=�(QUr
�R����&�Z�y����I�~7�<�i�����!02�}�s�
Pu�?%�|(G����Ll��L�ko0�D�re��CN�N�)��\��l�́5��b��Oh��E�i-��3�s�$ �N��Ժ�3�0O�쾁��'�1��fܰ�>?03X�~�9��s���(D�������-��G������Xtk�p�ɠ�l0�e����e3�Qq���20�� �%��Q��>�7Y췿s���!�/������c`�*�=?lҞ��T�I�o�-&�C�W�x��|��x�w��]��2��%KQ�WⷂW(es�}n������i��Ff'L�u��t,ns.�����k�.F_dܑ�g΍���)���Ӌ<e�B�*�88�<K�JY�c3`�~�ޟ ���;���#�����Ŀ;#��<F ES�6JS�[��-VmXk���Ă����ײeLS�m�LY�g���w ,V���,\LTV�Q��5BQg�}�� �?D�&lD��N���+�=�u�7^����ˤ�-�}���<�	G��R+���T�C��=� ܚ,U)*�*<��Ly���@��\�����1�����?���8S�O]��댴\em0��+V�ox�����t
��p������GqfZ:S�v!��4�K �s��i�( L��F7�'h:h��&<>�o�T�IK�D>�cz��OvN[�D��٠��̹��V럯&<�宱H�^�B_ת���:���d���T��-J��.!U���N0��9�%N�jג�C�䆎�&����yl��v[٭���ƽ�A�@ʏ�WJ�AP�;#�H��
��yq?�ud��W�>�6yÿS��$=K�	k�8�m<�W�X��s����Qi������Gv��������~���J
��0I��c��=Ž��WQ�H����Ȏ/ղ[�MDh�κH�s�nrŽ�{���@�� fw���;py�l����x}�Nrqh��q�h@N��z�Y����4V;�.n�}1�����y����FZ*m�)��t��#��_e���%�ƨ�N�]��]�%~~��-EV��G�#
�İ���Q�r��@AO�R� �㘤�d��"���z%���{�4�jp-Z,��Rg�e0n��#�����u3����yi������ts��،R,��Y��)u0�ވmAk8d���PM�T���ׁoh�7@)�~��o��7؁w~T�2�K�)i��-�����pC���5B���Ҵ��4������D�a�m	�%���n�>�=]5Mo���t;�ldU�F^��f"մ�ˠ�i#�S�� i�B��op�s��@���k���:�΄I�5�^�<bTW�Ō4��lt��&@�F �~�,���9�=@a�n��V��:��\��a���"����n��pi2�v�F�2��`ָ����1�qi4I�:0��*����7���9���<�ԟ�z��-i����& �������t(�򄌴�����}�<o�`���>3X+�+:���XN��h��.K�3�Pc����N�gn��}���u�L����\ũ4I���p(�P�SV��m�������k��s!�\�-�����P��k�.�B��C���V��:�Vf3%E���(s��:��v�od^�f\C�9�8.���@���<��Tb׀��'��!�Qn�`�,�S x<��r�ğ�j�xz�nK,��.G�{�����T�9�ES��r�)"��/�,��v�,<�C3J{�t���-o�>L����]o)I�M�+6>� ���%'���DԳ�jϮ���K��x�kJ���P�*K�-ģ��/V|;�X�)�#��+������{�J�'7�I�r�jn��]�٩�w�#���X���BIq�"��x �#�^�����
n�ӈu�cֱo2����H}j�bq�V�ť��0s�%)*Õ�PλG��9�,�x��;S�l'/#q�a�u�����@?�C9Y%��oޖo߾-o�~� +n��P�8p�vIO��$�Xl�ۯo����Ş��є�
� F�p<2[Sm
Qm(|N�{����l���O)��e�mS9���9��*	d�nHP�iY3�J��X��bRDYԁټ��	N���ɭ����i����NMm��w,�v��1'4������-���uEM������@�4�b|Qv��rj){^; *|��1��!�z������ꬪ� V7��J���F(�[��gw�O�-�\2�f>��������g�aa���C��gTS)�}��q2�s�n�FN�a�r�*��K<t�39����f<|L������XGD��d߶7  ����/�P�\��zpr��h7�����e��s��=�F�ɏ���V�*Rrd���k>)�&�U*�?>e ��D-�t!s��16K�Z�SK>J��;^�1"e?���%?��N���N68pY��ݻo���,��O�T~����ÿ�������J�ol���N����onI�Ɨ&�\���e������/���"����=\����~u�X�4�1%�6��6į�ICn̪XU7#J_S�hC�]w�ɺ�]td�xnO,�Bvξ�����J����.�<�Y^����>-B�����r~�����)�F��6z'��/X��U
������P��-�kM�߾O&����H��cB{y�/�v��0Y��(��gp?�'��Eը^Ǜ�-�_u��̒U�0�`r��z����ό+��9,+����e�y*�n�KN�m�܈�,ｏ�i��M��PQ[����~����В�Jc(]�awE�/�IC(~���*�'��+AWgT�_��[���<u���
s�����ׄ�6�Fz�G�_��h��e]�N�֛%3�ظِ�������Tl3R4(� ;e?Rt_������<����C�ם5�8�s�S%���~[������������|^�g��2[舾�dHw _mпE �F���o�߼�*�u=d�q�������}P6�Y��x~|N�>���s�*idfE'�a�Ms��E�xEF�4n�N�Q�8�4{�:�ZNN�_1K����� ��~�M��1�ȆFi�Յ �M"~���dvK8l��k@��5�A���jDh�]��w���� ���^m���o�����-�����;#MH)�8�y�.Qj�G���K@s`�%�\��>��3��=>�G���]SN`L!_�ʟ�ڈ�k���le<��җA0O�j�%a#>�]5��t`4;�/?o\_AB��c6�Z��"膫����gz^���/b�Dއ��o�����#�U8 ���ä�8�~���i�W�mZe6a؇��}}�b���L m:�k��2�v���qCJ�!��k*��&	{�bVVM�8�\�Z���A�G�hڟ�� �`w̎Z�E�>�ca��
��%�E|P�Qs��w�8s�9j��D����m�b�D��>��A�q����.�T�;� !���Yb�8�u~�������7�Xa�P ѱd�r����y���%�?��3��j�'L�����^C����5��n���P�����&z:?e���:��4�f�C�3�`� ���cg:�m��!f���<�������@'��2>S6�ǤU���T����I's'�j���<�u��`[h�b9�T7�jp�!a�黨�bͧ��$\v�*Q�:o�F	���2DzM��.
v� �kӹ�p=��l۰M�P�������j���b<s�f|�u�*	�����C`��j���k����������8�����~4��MgƟ�G�wqy��W����_yTt�tF=玕�;���-?r��ty��*������/:���"4�������F�I�w�h:��
Ej4�mʳF.&Y0��`�Opf��φ�ۆ��͛��W_QG3�{*��(�ǒ����j*�Ρ��,�8%���b��;'y_j�4���>}ܾ~�w��>I�>�ָ�=<����`J�	n�IӇ�KW�ǫ?�̂��\X��1��@ ���,��sL�AK�)����^���z�Ce ��½����Ӣ�%�(��
;�����;N��r�8�*ԍ���"���ƷѓS��)ֶ���q�.(3�l�D�dC�+��#�}D���^�뚴��1g���G�a{Ox��|T&s �+�p5{����t��Y�����Am�u��q&�N��P�:&>K<��������J���C���Fh4u�Ŕ�m�s\��T|�6�pM�t�{w��r��=��X�����z��T�3�v8�S��8���K��)���G���~�RJ��O��v^��k��3�R2;B����%��5� ��z�p�5����x-��#^=	�Ѩ���;�t���3W���M���1�~7r|ᐉ"����{��c����V�o�2�ZS^�x��7��%?z1ne��-�}�J<���]������PO1]�@��>j�QrW1c^��蕉`ڑ'MܱD0�8�����o�F����C����`�BN,j���������>$��N�Cn�{�q;�)A~[Θ�a/�P���=Ҋ�2f0e,*:k��뜳�����/^�~Lѽ�Fu��}���;C���%S0�h���Qih��(����U��m����u� �������)������.�L�t��Kx�1	�[����^������sׅ:��b�mZS3U��Y�b_�Ȗ�V�8-��]<��<�#E�;S�E^&@l(m�6)K�Q��(��	O㙊X�w�|7�X��6]��d��X�]Wv�Ӯf�_��ͪ�����@fGMJ�S��Q�T�J� �����p���r�񲛨��a��E߭������)ѹ�-��"h h��ق)��� ��sH�1��bs���V�2�TRpk�aC��cŔV���Q��/DC����v�댷�%�����YRŏ�O͸��ۤJ!�����!�_Ra:��].�t~���<����%��nAb��rV�_c�-���.�����z�uz��lN�S�t����sj��}Nj��U�Ÿ�h�L�9�A��"HM����fx�)��	��Q��v��1#%�T(�%�\���E�|`p�窻��KdT�[첔�]��P��"�Z��#�i��E��{Uk�f���	�i�5���]:;�c?�ڴ\��x<Z����\X?v
�t��Ӎ�!��5�^�������*��?N\�)�`�Ch�l��a��?��G#��eWϛ�<�8z��)Q����gv�%ˣ5�o$����v�����KM���ؑ�)���7p�J�UGM�!�YQ,�g�g�'|G�R)��b[���Yz<'h#h\��nu|���p��G @�v�mޭ��$7��N���ٌAg{�wT)�  �8�|�F�d��ap�rd?�Oل!�Li���4qU��v\�C6ָ�l(!X"[j �����i(O/�x�BE�큀�n9qm�_V=[�O��
z���~ `��
�����0 �^��0K����0���4���􉃑�����<��Aa���wI���A�`��C(�K��ݴ����uêr���� d��S��Ug&%,�x=2;_�9�����k�e�?+���`7�B�~gP��?�QJQ��>�j���G����I!��s`��Mx��JE���?&�;����4�8��G�`�4�>Y��
[G�4�C�v���5�ڃ���P@�zT�k ->��/jҜ�%	��P������L�����
Q�\-�m�a�J��&'�Z�Z������bQ��"��5�}t
��#����b�XPq�.y��9��x^��O/^�S#J��MⷃrOLid@��)o���Ǔ��^�1SEKN�Gooz;������_���g�fIC��|0��)O]�֪���ߡ�:Ӫ���'6N�o[vv����	��Au����ߥm��l7N舕�*d9e`���H�M���l��sy��W� �p�|����G�5���±Yiǎ�L�� C�nf��kbY��E<�ʴkH��&?������^ۑ$I��9	�Y���|�=���s�av�{���d]TD�,�Y3}�E�hdeA���TEEE�I<`"����{W�)[	�p��fe\��1>Hj:	�ȡq�7���6�&��xs[5.��ʾ0�l��6��4�*�w��I��B0��0�#e�� �EQ4�D���>���~ q�AЄ�O+���^C%�����3+�R;8��$���+W���>��(j*Ji�S�F�H[���$��i�d���&#5��&��OOt�����J�I87��f}���.Ū�t���U�O����
���	��VX��j������~�瑪���T���%.:������綉����[����g��G�s�)26H(iFpCѵ�N��c���?%O����f�a��Y�.�/��Ϣ��=�A�M�^�y����y��u��!]J�GZ�Θ�hF!�{�ρ���w�i�m2\ |����]g�is����������oݳ��#�.���(�I׊�# ���`�s���	M����Q����:�Jպ1"�<�����L���x]&S��:�kř���.;��^���j�*�p�܍�P#<6��9�L)���$�4�Yt�4�:)J�g=#Af�;ds��߬�N�P+��o߄���h�n{�!�3\362�H$�u͌o�s���Ѕ���*�Z�������~��>�m�0�(�?���9�Z=w����i�E�V־f�K�`�ʣ|3���m\D��r0mJ�8a�鶄).O��'Mκ.k�P������� i5b�8/sf
�(AAA�.�'[����_�?GG�%۾z�����Jט���NǰP޲�(b2�Z��Z��%	���>�e�mWv�3�A��^�LnE]Rak�s�Į�X��3�v����S �ۥxC��cg�$�9>�P_p�B0C�A�4��)C�]?D��f6RN�=�FdT M|߇�K��LX&��:��+��I鹣u�*�e-o׺�Kut��&ˡ��gb=5Sv/�'z�T�w��W�s��{��V4�>�*(Kǐ���0��=g �
X؝�H��r��:�ߗM�֡�%*�\���_�z�����D��������~��]�;���w���C�T��~�)��ł����d�H���7�XQ��k��C:
W�x0�2��4���?�5_C��,���bX������˷m��w��#���0��_��`��}嬕��������"�I���"�X/��J��74n��[+�3�[[�a�M��'1�}tH�-�y�(*��)/A�(QR۹��+hz/�'�a ����t�n,|<U`<��M>���dJR吶�)N��$7v=e��Fz�ṑ�r��$4R�)�"���Y�9����YZ��/������~��i��c� � (�@K����3�Ev��e�����������E�$ϵ�:sn�z���d�'ݎ̓�m纫��ns�N�*;�-�.i�?e����@A�v��E��WT�Ᏻx�����Q��=��~��(2����^#W�=�9\Ʒ��A7��2U���^�w�Ux��^��	bD�=X
����
P�2��;&�29����x~���4<U���Y"*�!3�6a��h��}�r*��]�? q>aUYL֋ l����Φ��
�5��ן6����d������	L��1f�"�˺��ҷ%��E�����:ɗ��2]��s�s?��WYs�4�HwU4�6�w��"^�i4�>&H�8����L-R���#���Iʟ�S�xGe�#�43��&f�Z~N� �T�?�]���9��3@X��j�ݼ���R�R�x�˅A�WCd������uL��v �q8?�z�l���iE��?�O:i[�	��0�~Ն�^+g�q�y�|��rQ�#K�,�7i��03cp�>w�K�T�gD�s��`�i�iu7�����0��Z!�Avǥ�ݘJ;�N���n�t��M[�g8�$'dr��쁅�'4�l�;����\o�}4tx��om6�Q�:��fo~�JGS��ÊJ�3�a���p��>�L4|����6�WV�z㸓��tZ)�Rj�i�hаy��O���ǽ|x�X���*�Is�N�
�������������ĭo�o�ݟ��5�&0�F.d��g��e�ܓQ%ox[���M�	�ߚ���+V�!�%"M�|�)�fS~��0����1�b�$U�c�,W���S>DAJz��#���|�n4��㩋 �<@��S+VX�c]כNe�g�y����g���H�>d�v��&lU��zr!��z:wWU!���4=�90�)}���EҬ��/w���w��ZI*������5�c݀���ԯ<�f���UU�J	?����1�a�ǥf���u���۔�F��^т���5\�yn6��冩\����~�L��.2?sC�l*yOz�u��,c�lDU��!>SCi��T��I#\K6g�e�Z��}D ��	�
�t�E���w}�_Mi
f���l��7$v�jx���E�;56���1m:9I����V�}���\y`�~��ݖ������/��,r�nu%c�I��4�̹�J�n�H�\�_dnFw��RT��}���Q��Yu'��\�Gz��v3�!΀��j2�����?G7?�z�<l��wt</(!.q����Yt��~>�~�/Ȍ%�wo��F��>|z���pO
��}�e��ɛ�>R��!���t[t�_8�	퀟~��|�����>mY�p�2.Cfj��I�� ��ipwO �&3;�$����v�AYB�ߟ5.�L��a<`��d�k^�	|�,�JP�
�zj�Ѫ�9/� X���N
jr���:�mo���ܓ@~a�Χ�>�4AS�>+wVG�|'\��3*�K��w��.2{\S�N��� v���V���|����t4S���� ���$[�������kx�륑b�B����f��t>�A��+�V4:�9Z*Wqr֥]
)ĝ�2�AJ�ˊR��2m���27�ێ�r�$ׯB��m��n'2�ei�˲ˇ���u��f����F�*�jb�C�� ୕6����7]�x�Ncl���	�ޕ��**�Oe���P2����Q�
�r�U3|�P`Q����u:(����C�g�I�����R�Yv�(���@�_�i8Xp�M�Aĭ5+F4��I:���U�;���������Rf���80e���ݩ�3	��Ӽ�����A���xN4�v���������~�Y*� )F<�Ɇ�/~σ��E)֌�KWՒ�p��Ț ��5@��>�:���
&�t��c��qϑ��?ż?�w���*C�Y��� �{�PL)�q;;+b�E'��8:�۽���������\��OSn�N��"bd��C�F��z,���u�h�5bZ�����>��xx%�7U��b�Y=�e1�p��H�棓���U�h6�e+�j���;������gM,U���R}�����ƭR���2�Z!|�_�W]{㤼�~!Χ ���3RO��,]�����P}�o>�_gQJ\ގ��"�̥�n}�,�+�2H��0 ���#;��]Ⱦ��r�y�;��I�S~���q����l��ö��ȱܝ������_��������-t���S̶�D�x���e�����D����a�<.����>q�9><LA�U^!���e��>q#AAW?�8���_9��,#����&n�I"& �k s��v�k^�v�$�t����fU�c]O�Fp��u/û/_�D��t�l���Q�y�8{R|�Y�nZ;x��*[��sMB6��%�w��jz�U
8�?~�����;YĦ���'������`~��4��Y��+5�����LoB�� W�*Np�IJ��߄�Q��s�f'��A5��C���6��q����&�Ki�3W�Ff�s�����z�����,÷(�~��9�yW`�Y*����	H����xb��VUk��u���$:-N�,{is��g��� �C`��u��������v^}}��t���i�����^*��g^9���`0J��b��@�@�Zm�ٽ�����qm���%��v�R��L��X#���=������
Iw[f�>(J��7��r�y����t-��?�ٿ�������q+}q�8������ز����s�r�5 ��4O��b�<�/���%��%_̾Cc@��h����������c%�&Nhl���c���;lȤ�������>��
D�I����v���x�X�O�yhFV&\oi0��dY���[�U�`�d��"2w�!Sqc����=)���2�ޝ�o?�Wٺ��
ci_�XLA��o�&�:/�m�qؘ���~�g��2�@za?�FnW٪��h���^���楸d�h��R�_$��wc���X��������$�N<lb_��V1:�f��r]p��c��d8ßL;�n�jw��B�>�M�D�X*�?�����,`9^ja$꯺7�-Zj~ږ������@�'���-�f]nL�B���SdDA��eDH�5���I3؝>�*���'�_�!Q��j�BD>�J'-��M`�M�A�ԲNc(�G���顜� 5<�z�����
#��54�@Ei�I������?�������@����	S���9߿��F>��2NRL*ɞ6�lD��T��yfs
_�8x�_>�2ﰯ�t�F9渗��A
�,��%��EI��?���*��Kf���s�N�B,����߱�F�����Q��s�C���1Q��L���h@�(׮Q��g]��ڇiov�]y�U������}&[���	U�����Wr���m�n�����1 R7���+�v�eiܔ�1�3]Ū`��c�-��0{_ҋ<1,�yN��h:��t>�b�����2y���Ƹ�{��A}����h
�{u�8�i�:�}��
=�<�g���[�{[k�LB��k��j�ۃ}l2��V��j۪ +�7�^�����zţ?ID�=}���Z���n՚��&���'{�_(;��ဠ9�oِ�����p�Y�j@](���5ښ��=7��N�K�"w��83��ih5��=Cl`��&x�S�T,� ����΅�¦aa"�B�r��?����Q~���#�3&��?���N��ӝJ�O�s;�#��I����{MNu����>]ʗ�)`�о\Y`�(^��1��턗�.z��;~��~�B���
�K`��}����|�Yq�C
��!�q�B����5>72L01�R/ ����p8�s��_,Gyj�WC��`����5r����V�G�7iM�^� �wp(9��Sn]� v\G�925'9��J���fs��[��3����y|���Ý�	T���fw֪(J"����]H�R�T�����8�v�� �����3��?<�G 
r� �`�������;�#���GN�u�c�?N]v���T�m�/��Y�$��l6c����k�k�����2��v�$1%ߎ��Q_���TiT.��o���eb��5�Mp�DM��$e�
//�lV%�d�x�������q<��K:<x��
���:V�کXz��6f��<��aBaJ0[��d��((ːaOe�扌�ܫ��uCS������"��b�x�e�wЄ�]:�t8
�!4�\����(c�|�\�-�]�_]�U�����!)���=�E�/75,�vz��%1�� /&0�-[9C�s	�'�x��|�#FN�7$��|�j#�K37zm�^����1l0l�;���n���u���ρ�Rq���lҠ�k���;e���7w�|tŢ&�e'B���V���,<� ���*�C����矻,�I._�`m�r�!N��j�a5��K���;��E9�\S�|� 5Q��Lz�ES}�/�;\^�Z��hG��g��9�MoI�I�޽
����O��R�j�[��1�#��J�-^ږ��U$� �����?SK{Kx�KJ_�S��,}�8��1N�A��y��O�I��1[�O>9kK��;��5 ��&� L�󲞢���w����UD6��u�,�����D�C�����q#��B��~x`Ge	0V3J��g)�ܔ���&��`�nz\����}ϭ|O����.�9�+]1�X��@��^D�
B=���-"3�˺ُ���AW2��x(���ii�����E���8�/k\я��iv�K��r��e*)O�0wq]@$�ߛ��k!�޲J��R{�9gq<�Կ��c�lb3_<��^e���EpQ�}��;��tȍ=�I����6�����h���I!���Y��@DJ1n��D�$^�*L�1��X�]��v��#l�)�1��u�:R�֤�x��|D�(�k�)��5}��0���:�� .q|�O���j��*f���߮�op�6�d�����u�ɝ3g>9J����Õ��@�6�g��ȟ;i��1Ƿ���(�<c��%�A�k̆Ƹ-���'���X����5�=��~��tK ޼Z�5\N�"��-*�w͘�sv�q�7ŵ!�����اǓQ� @�uX�Z;�x�uK��+��$� �'����lӞ�T�y�2���sX�O�u0gP�����a����I�'}k#�X����:�n��d�ꮿmd�Y�h:��r���i��ف�@Y�/)�LݓC�"S��w����O���V/M6�d��;���~ps��JN������8�Y�@7ub{F0��E4nD�i2-��ݐ����H~4)v�hss�͉%������CX|�PBa�.�R�{T滫Mb�x.9��r�B:)yJ�Q�+B���kb��U��>�-X�����lTe�m��v��{�=�_Mi_;e�K@�xe��Dn7�pӀ��.��D+��{��r��t?��=��au� ���n���!?P��H�U�B�ˎ��E�Y����ɑ���4/���9At���U�Hi��t&���Gzm�����o����b��CRu띑��D�ׁ5�vl�[k	��x~,~tϱ!�]��U���d��9M�X!P��^e`ڏGy�Y`m �ڰ���N�wC�8��)��Z[׍Y��8L�h!����&��۽�T���v����1�	���N�A�4Y5$�g�*,kN��������<	ϔfC����A��̒]�9,���c�O����4�Fʠ�!�k�2�{�T��~4�i�*3��+kf��i�Y�Y���B�������N�9�1Xdy}�q"���SjkT��9�6�r��f�QU�xq�����L߳jܺ�e���_�������[?�d���ԔnU)_��i��%���h�����EtG8Č���z:��ۈ7V�d+�4&`����rf�5�i�;I����7~h\w�,:��q���U�x��otI���c۱sF1���xXn0�8eE���G���^�$���3�Jf�MY͵[C�=��&v?�C/`�9���¾{���l�E���f�$L��h|uူ�g�(:�p��9��թ9��w��c}ob��4���s����q'Z�-�������1\7�T���k�Y���)3�~H��,ӋԾ��S��(�1�N�R~����s��'.e��$"���I�ρ�B(���#���hN�w:%�M���U�g;ꖵ����c����g�~)�߯�z�QF��������3�mЇ-]��Fų�X��%��	ۍ�l���zm�R1�g3�!$U��˾Jا4��ϑ���b�S�)�f��*����Ds�8i}����WN�V�Vк�ʚ2e�Vc,N����}|Rs<rigNy�ԓO!n�P ��?�:��h�&5���j �ɿ_�=jr�1���Ԣ��s�L�%g�$�9);�n�0X�I��᱄��y�;�A#�&薜 �b�UË�*C<�J�'��s���m��I����-��~���~JQ���	��Z)����Մ#����{(�ј���:�["�YS���M Q5��\�fk�u����K��,~���7�3h����d����s�^��_q3sȩ>D�˜TVH����gp��� um0�R��3��+� .�q7����ϋ���զ�&L<�Z��X�p,��0/�c�ሻ���>k9O�ܪ��yni_A=\Ki�Q�+���5�q���g�g�;��#0�pR��W��l[,���\Ҏ{M YYo���z��g_�0�5��Q��e�����#.�g����f}�ƥ�5.]�$�*ߣP���c��J�ͰWL�8mY�5&��ǐ��S�N��9�"�hC=����[�7���#0��Jn�m��yf@�˝F[���E�S���Ox��	;�|�yzƻ<������"P����e�^� `�I%[	n��0!ٹ� �Q�S%�%�������Zf�����R�"])��[ m�l�=���~��(��ձ��c��*��C�kpIn�{��^��Y��>df������9��b�3�Uv�Ywj��^����OQ{<vE�&�*�\u���RXyִ��,�s<(#��(dy_<Y�,��8#�B`��}� C\�
P�H<�		e�P�z��j��)�tzIA+�ה��
~��&����A�CP?�D�Xx5m��������ϙ,�Z�W�Z"����Ƕ[UK������0���� �Iy#�Kro�cNR_�e(W��9��]���q�As�P@u���µ%R�sTzU%k[~/�hsS�{`�#ۂb�U΢�d=����
�K|������w˜�;�sd����"����Y�f�`^��/�=��E:����2.�NU���p���%��ך�#3�Qx�;Ü���'oķŭ�d]��Lu1��Dդ\�2�v��8x2�i�-�m� ����IK�ɵ�4w���R��gUV�V5�`�u�Њ�p�G�����l�X�����k.�^3���x����s��Kg�r���`�M@�N�+��+ENju٣��)]�d)2�yN�Ӳ�G0逨\�'R�0�4#Q(f��s��Y��Sy�0[3�*�I��e����/5#��"��η	U�!v��?}+�&����m��s�~��xRlRg�~��`ĲT7|�#��8Ҫӛ����SF�|Y_5Ub���!����<E������X��yMQ�g���-���"������K���Lx_)���$�x������tn6����p�Ӳ���&��	|��jY�o5t��vF�g0#�Nk�t�Y����hF�`^{�02�P��᪦����Zf���1\ K
d�1����U�,[d���}�J�`�|G�]�6.x����bD�����qp-�9{	g�Ti�!2eWf�_v���J#���3h`v;�`�=���7�k��]�Ed��2�*^����~���R�2G����+9+;F�I�Y���.V�wr��q�e�i����#����j�Qv��H�����g��NE$T��§^ι�>��a�É�T�Ⱥ�|��f1�zOy�8�7+�zo�؛��U`4����D���ƞ���n�,��l�՗I�P�!�9�q�WJ-���kD���<�T�����Sr�4i����t&�!���� ��9�����c����Z��׿� �J�5�ٌG�PJ����)t��ۣp�o�l��M��_C�Σt�@z�pσJի��3�T���L�`�x��4�����"���T&J*�1�Y!��+������jS�2U?�w����Ỹ;q���տ�����R����sL���KY^�h�\E��|6��r�*���`z��Ń!��@�&z�l�,��}�-n���6�}TD:d��FP.�Yr��,�S1Z��G�Z��l����:Q��	��,��a/w�52I���+��.�a�� �����:}
k��-����y��0��`�3>&D��^��u�Ux�l�<x}`��F�k�S������π�l�.����<�e��Ȏ�<�k�2OH�����n?׬6GD+U�[!���\�k��}��8����m������y�b~�rS�s����`�]x��9^j�`�jv�,�ܼ�� v3i�l�_`CU�b�C�=���+���?���g�����B�m��MCΰ��o��Z�����H��熒�D
�x�oZ������zs��zyvw1+�6�YaY����lr^���7e�^��?��s��OP���?~/��;�@/ �4���UF:P�g��%Fp��|�}��o����������Y��j2 �B��������VV��N'7	H����yϗ�e��i�>�L��2�o��:D�b6X�e>Z*Ek�S�3:�b`��2����E�2�]��[e��Xr�[��PX�����Sv1A$�mdj��_2pO�9�$�F�i�H��m,�=�k� =`հ$b��5�L8c���H��#������/����1?w	M�_� �ۥ_t��y��w���:#5��b����Ig�HE�Ǫ������ϩM�8��Χd��\,�唋�V
���3�Lk��U��Dpnn\Xa�x)Z������)�i��<��� bG�=p$��4_���%-��x�]./1{��K<������TTHoE7�#d��A�u���6,dʰ�L��6�_�=�}��1g�B�˚�
���ݹ@�p�t�C��8H�U�l�Χ����i˸?��,!ܶ����_~�F�R.�w]�bZ���u�EN���>��������My�?n%p�%����9�`~�B� �	Y������C�-Hu�,���!���ch����;��C��޴��TY���Ҽ��������A7H�
�YҒd�@��f��.�1���2�^�~�6�ٴjEj&��-Q�+;[��XK�0y5�Maz���{R&��u�'�G%;l���KX`�#���T���G$��)��2���u���)��]�;��ܴ�. .(o��B+m�A��lJ��p\x�]/C��+�#�0^���I5����/<7��Fm�����-s;�V��=�*P��%�e�� b�\�_ҵ�����&n8Ɖ!�.������l9��@*�(��zg������@
�P4�5�6��@ ��P�0��)�it+w�@�����@�,��ᰋ���D�}z��|���x��c�����P
N�݀	bAl7~ �|�Hs� �Tt����Rg�c�@�Yٛ�2g�J���L	bDHQ޸���m�T�<w��9�<G0mC�]��q����u�>K\L�HF�v+^<S@��s�y�OUd�?|�v�0ᩤ�?������~;T�	�s�V�C����1�&ͱ���C���H�.1�ET!|�@�����vZ��ԭ骡�[�﬍���cC��qX�w�D�hL�#�O	T�'��I�Kxl:X���˵	�Pe]�po�F�k�p ͉�yJ�'])I�+������xO���)�E��I�N��Y�7W�h
_��}���i�����v��#���%m�9�A�r�d���ҹ6��y�"�ax�mٰM�b(�/,��f��?���0�kd���z��7W1h��k3 ��vpd�ù��7�0����Z_g���.��T=�։�f�w`q!~ S��!���ٮWEsJ�%��\�q���i�`�/6A7�QR|���ȓ���Jz�ة?D����Q���:
��?A:��q_���Hˢ@z��Yi4��]���=�xB{�3K$���ve{?�بo�Ǜf��u��=���Kd��J�|+{�E��#2>*4f#�T.P���_b�g�"��{�-�sN���������ݛ���o?�_~�%����e�J��P,O�w?lY�����e����\�,tQ����=3�`G�i�NT����ɡ��Ʀ8��hL�M���
Ń!��P�
:�JM���|��lh��e��p�ʢ�cj>*��tU��NR������I�W�Ʃ�d�!9��f��A���r������:������MG\�@�U��.�*7
|�\f���?G �����~�C5A�_� .s��1�Y��gZU̪����tFe�L�u�r��1W
��1,���K���N������
����2/�V�k�֜����fiW�&�_RN"r+���a��1�׾�!�E��Z��^��3�}9t{��Z``k M�9ۢ��O�8V��U2E$�/���B�׌�)1��0#f{�R�aVJ��52�lܲ�~.(�q���Nwߨ)7Qd#���ۅT��}n(��E	�R�����A���AGEَ)�>����v���b�=�0q�0��� ��rB�+y¸.���ٰ�#�)�ˋ��z.��3s��Ɇ�Y`*D&SzQ�(��Lf�i��wrKg�œIb�>2���R��@����IsE��Z��@�a��ö�ͅo��|����K�`#X*�t� sO1ߴ�f��p�C�U�u2W:O��S�����t��X�a6�6�+
�%���T9ᮻ�T� ��z��\^����������I�li�.m��t%7o�ʼ�ғ�n�Ĭ�i��ÈC�R2��L��y~1�YH���9�:�}��ݫ����Xitb����F mh"q=�������G�O�*�щ�'�a�r�Ɩ:���B*�G:c�\SkjN�,!���x�#��	wՄIX�vUs�+]^`��Q�~�=�Xt��XA�u)��ꋄhDG�� ���m�~ز�-#3�ֶ��M4Gc����\īj	���M���[C� �
���We�3g����N^Q�p�������|Z@d76���S]�6.z�K
;�ň#���~W<�v����I4�7�����϶rt�끳X7A���jd���SS+�m��I���1�PWXgi��Nxݕ�ƺ�94�w+6�V!hS���8k�+@`�UM�����'���*z2�)6�����u�N&����Fgw4q�i��!��|����LV3ȯ�&�Q�<��٢�p��ݨ�A�h�}"˽�� I��\Y&�]V�QJ���>zO�XhV�5������5�vm|�[��E}�E�6����B$�G�[�4��b��j'��8*�N��Ȧ�7?K����+x�m8w�cZc�B�H̕�����6A�X�)�����<
]>��	Z�[ E0�.���!�,�ycdn{?w�&w�_���� ��1�����{��	��;Z#pw���#���$>�z�\�(E�l!��e��vˊ���+
,kB�B"��]4x�����J�8��LꤞԵ��SBϪ]1?�P��I4tǭO���1��K8l��$}Nz�(^���E^�]�_�*́���[
N;��jvZ�����l��/��θ� N1ɷ��j�ʪ��fk��R�JMO�PW�ig��)cx:3�`D�F�d�%��W�=����Ƭ���w�|XG"�4_�o+�5��1L�8���J���8C��OXo�zp4�	�WN�圿iJR	{�g`A4)�w�A�1/��z5�sDc���
k6�U�n�j���&�5���������˟|ys�jX�@3����M��]'��I�6D	��ڵw�� P�m�ՙ�/���9D@��������DYLV�ܮ�0���AW7�73R
#�lt�h��ib-!)�$i=d��fM~��-�~��j��l�>���.&x���(�	�#>P����ޅ�ɞ�Y�@|X|y��ml�"C�6	^):S�mُ���y��3�}jL���A�2$_��C �+<p8a�6 x1l�����+��2�8�Tn�t���ͅ,���*��r�
�;���#-]KM���Oڮ?I�م����,���\�� 9�o���0�f�v��k�J�,�Kt�cd��?��~��?�Ϳ�����2���m�Z���@�4JcV@\c��G9=�W�_q����v�qo\e�y��t3���_~�6�ω�����x*qQ�{�‥"�Kz���A��;�WU0\�)���e�zE�G�A �)�gS�BY�ĞZwU�|�/�VFʘK�`̕�t���.[eD�$ �
�������K��BG'��,s&=��m�Zb�v��CʾA�l�EJ�1�h��K>��W��=?��̿q� �/W�c��w�52�T��>Pc�� t�S�+o\Y�geūI͐^J:� z��\���2L���#�(?&އ��-+-�1A���E�C� =JY@N���z%T�>��zK{���H�*�M�`V�j̢�s���7o�^� �.�n�e.Ehv
���(�����s����2~��46#Z�.Ӌf�`[��y(�Fv'��֠5I�)���b�jt��e|�Q�Z�۔����r1��)��`?�*X��:k�n��y���7��ؽeC!hc�Ú��G಺�ؽP�p�Y1X�&���>C�Mq��*uR�=���U��׳��rjhqe*�m˜ڧK{��3�d�5�5����i���W���IG?��Z��	���`��y� ϟ��lS�^s�XLෝϧb)��S���QX+��2s�\��i���l�9��R�Y��T�&40�G�B?n��xZ�r��l��wq�z��,�R��h������j��C@|�]r��d�ұ�|��$e��.��cjf�>�V�LO*���p��x�Yc��̎Q����O[F�Kd|o� \�1��i�|�{�U��4���NЕ  0��)P��&g��@yﲊ���NG��AΘ��!v-��)��,XDgb��x��t���¬L�fUvJ��p���;؍'P���U���zI�	��!`��5�����v���xp��=�E�!hz���}J��}x|E�U�c�j;�%)�	m�}�$�ۭY�ǜ/
�s�?~.2������+(a��P0c[v�7l��&@�=�(ziӆ��X���?���U#�[��EW|N��������6|��𙥾*�K>�SMi���(܀���}�~��������,|:�cf0|m�\c\����[������1��X�A�X��腦X�^n����D
��pнfnxt;�[��[O���zI��X�jF�S����MbOuV��$�=�c�����<����H��D�A)�	��i�OR!��l&������
�������l?�p�:#�,p{�B1���sՠ�uh�0��*���:��cl%�����^�Hyd�ߘ�57w84ws6D�Vc&(��6#u�R��,O�u]m�}�8X��նoH)�@�������ޕJk"}M��'���D��"E��]^���n��>�oX�7|��u#KPe�(���=M �&�vs��~%��r���*9�Y*`F�{�Ā���wx.��e��<���[z�U3� 1���{��FL��t��x�T�p�}�`�ç�U���k�K(����)e��VP�2Ҹ�-F�OZ����en��'v���� �R�ڣ�5/��,�T�(;�2w�L��g������ ZJ��D�g�Kӫ�6���]I^!3��|	��Ҙ���$x�6��8u�{.#0� ̅�z�]��ϫ$�z
���-�#r��Y��펢��j+��d�c>�'�l2I���nh2ɾA�x�=qo~хSW��'��%�Ʒ*�)M�&����8��"��#���M�kۘ���(�e�:�du�j<6���Q��;���+u�M��x���4�ډ�1g�}k�W	�G��i�9�tc��^��k�V��?S�}�ܜ��v�,=�f͢���A�����и�)D�9'L��(ɯ6���Ӑ6-~�kI��k�t+696�srO�P5�������y���}72������>_�Z����:���o2T<�4�j4����W��(����F���N���t�w������&>\ȬM	�{�ڮ�&5� ;i҂3�T��ԅ6�R���R�r6�SBh8}~�T%� ���&::��g�z��(�I�>�Ɉ���I���.�AC�^P#=d��fC	����2�9f����1�Ȝ�F�}�~�~+��`��0]>�� ���0"}��`2����niқt�_Euri�6��g�&NI⦏=絙� P����g��g��+�r�c�VI�{�����${����(�W���C3�)�;�7c`��'�R�}b�Weie]�˼�`p�fT?��l��t洔U��
8g8
&��z�ϟ3{���5��@���;]KŒ����S5{?P$bax����~���N���������ON�{���{+��>�7Δ#k�R������MFm�V�V�شDd���e����V۠�J��y[�4[�M"o�B�����3F~M�8]��������ec7�7ʬc����@�M�g��4ik��3�7>���2q�љ2@�,�9�PV+�W��+�6?o6Ƀ6�?� �#�����$lt��;w��r�D����kE���<R�=����i�BzpL�&ş�ՙ|���^�ԥ�E>Ձ 6V(m���/P�~����S!��}��{�]�8�	%�[G\Ϡ�|�Xln��}qx����0�s���kmcH��9������F8�>,>/"��^N��)�.���[���=�\~�����������r͌�M�
b�v�C��(���s�@��I��rƾh���P�M�Q���ߞ�*}'�0�Z��uκ\�H�b,��o��rfz��@Z�+��M�����^�,����� �Iez�x�c\�Y����I{Sr�C�{6Ogz7��p6j?0c�9N�} �c�#�,�!^�ą����4?�W�6��F�|��5lW��>��O�m�&�����Z�(L ��(�:;)�{� d���ɻ��_3Rlk~" b
�⹫�^Z�ūʒݼ�����h�t�I�=��[I� ���?�?��#�L��x7�{/�4���[q<ǻw�#3���c�72N�f���;��E �&��N�����H��(���f&Vf6���� �&�_�a@� ����X�x�UR�k����1M�O�w��E{���AY��X��H�tFc\�L�
`�|�/l�D6�����#��e�{�J� $����ֻ�V������5����#�c����Լ`�����ß'��}1F�k��x��9$�.����ɰ-v�1I��#���l	��_<>ݪ�R���5��2�D���S7� e�O���1�cik<��`zS��ͼ�Y��V��i9��y�Q}�����u����A����!�:����TJ����;X�`�`���T%*�G������2Rܨ�@qڮ+2p�h����ė��i�9(jDm���$	��z &��ɬ�N�Bo��t�Su������5קYybrt��U�c�:�i|T�+*˧�'(�o�<mCa��e���M)��4��K��D�,<�kʷiA]m���MA������<jgB��˹|��$�EߝP^
C���yxf����>o�������~8vnω�?-��B�g��Bpz����-?jы���_g�Y�w�}n$d�>��Ŋ���w���҆��o���p"��p�M6�e4�J����ް��p&����0�.�� �!6+��(�l[�,�5Fj��~�.���B;�(j�$i<�Yp�!��U<s�:Ġ��Ȑ�|��@{���(�=f��e�d����ʎ�8h(U	3�h���2�)�B|�AS�c~�M�H{`XSɸ!��ԫ�)D��,v����q?�*{��>�M��'�ph@�|�U���V6��d���C1�k��s]^��7]�t�����K�iy�����A`ۂfH}�l�AsIV�{��-�zۤ+�~[��d,^oy�������%��7�sP�E3�l�v�I��*)R�C��\lz�����&�<C�2F�w̎߼��?[jYh�jp�ԙ!:Ѝ�͠[�lΙm�/�{�N��DЬ����)4�"d���O���R�A�I�7u	��Gᰩ*#z��N`K[f6�.45X�0a�����x�����%2z�&L1�����놛�v_�|9��}���u�A	v�G�3����W~�V�$�3�44�[�]�� ���u�Mm�A!6���5>'�~�u�2��^�b=Q���;&��EJ�n !��(�q��c��`��t?�z|1X�n�U��t�<�4N⸛q�	u��-�2e��J��c �Ѹa��tE��㬾3�Vr~�O�f�X]7ϱ�^�YF[�p���c�\j ��"&dz�&����.|ä��L�?�J��@�u��sOYd��V�/�����&���"k��iT��ƫƓcnU�#�\�6�}T��7X+�7��n5=��䦄�y;�M�݋0�����$�j�ƓLݘ���'{)�1�B<�����=��O_e�s4Xp�� 7=�ٲtuD���w[���w�>�������#�g� ��ec�(_pS��=AdDc�1'�$fM?��d�Yo" 2���(j��lK�y�5��Ev''�hF���^D�:���8��.I��?=��T��Y��(pL�0�B�]� μ�W�����'/3��v0���Қ�sQ���,~��2R��&��9���(��4��[E�����?g0x����Q�0r�	��#�x�(��َ�9>R�b�^�y�M�������+krp��Yރ �/}m���}`�P��3�v�W1��gg�n&��~"������5fK��A{�\��q�}��	#��/����pd�q�b�s�����ӑ-����+��(m͗!V�%�:�XL�D�oe����w0]o�O%#��S���%�F�_[��v�}��S��h:���Uz8		6���҂�]��(nDJsb��ǔ��@<�Z�ܺЏ@��'����]�����6����-��)+]���;�?F�>t�*� ��nv'���5������Q�13��9W����#{��f)X��)P�M�R'n���Z�%�O��wH�K<g��gȡ�B�#8(�c"K����8f�Oa=��q�{\�=K�c=(4�JW�%J�#U��RWao�*4|͹x�O$���^-���g�FYflN[֖B5��4S�%���������j���ԤX��x���R�d!�P2�C;��� ��u3�{Ҹ�����C��%�E�ks��Y�g���D[T�sW)���D�b#��L��t��j�y+�R��?G\��V��?{k���qX/�8���ZI[b��?7���0�M��=�.K��{�l�Q^0N�-q5�DIe�j�� Y��J�^s��D���S#N�AΘ8��d<�}����փ,%&iO�?�����=K<!T��q� ��)��>:܀�ep�2k����������D`�u<_�jw$�u`�猦�0#���}F`3�{��b+cQ�T�D��ƪ�m;D�4���@.��9*K
{<�i9+��m|6b��j��u�)�U�U��D��,1�)N��i��y:�s��if�m�e�	�wr�)�0��ɑ�R���Ig[WPI���[+<ί��(1;rG��t�<�ʤ1�w=��>f��g�"�{]q�A�@�lg�#ѽL%bf�i1+���O}бVA�},��U�ö�x���"��]h����E�4JF�G�8���Q�&�D�rM�c4L1H���
m5�Ӻ�=`�e_
E.�Ӥ��P'O�\���76����M)[�í8�/6�l�3u�r]�Xmi�}�zj�6�+�,g�8�������5�p֚�n��Vw��CҢZ��^��|oƷ�����5d�A�lt������
����hm��W�(N��7ǜ@��)������C|��x�V��<|I��U��ڭ�y8؟���h]�D��â*����Fm�^K�XS/I:M�DǛs�g��Ĩh�3)� �x�p�:����P~`�68��p�ʪMx�cm�w޽{G�Y��˒���׫�)C���
������T�Z�":�J�t��=џ`p�ش�@K�>�G�{y�/�&��M�"�j��l�����2k�]�ʒ~(Ց��Cf~}��a"\v�븫��y�e2�V^�5i��`�ǿ?=���l�E�u��\�����V��� �aٙӄ�.>/ /04޿�7Ɵ�NZ�Cb�d+�%&�rm���}��-��L�����x'�F�`BuK�sHpc�*I����$̜X|��.�J����	�\�Wͦ�+�R�,cl&��9�T�{�]4��YVtn ��h,.��f �w��PZV/�d}���A��5�N ��ǔ���VѶڒ0*�`򶅳�@G�3�o�f�L�"L�DAiBz0��L0U��%��x�xmtÂw��H�e�4E��92\���#^�\)&	6�9��s���v��6����;��%q֮���}�um�Q�Ly�V^ e
4\�OŘ�x�_��	�� 1p�L�2�|1������g�M�M ��X�� \��/OdMi�]�����U�"��ԎY}s�ǽÅ�ld��������;L�8� ��f��Z1m�;ƚg��L�YR�U��������x���F��YP��Bf��	���y��������`I]��z�fX��STd�ځ"�!�A��=�q?2��z��9��àY���+�J�E��ۯ�T��+��� )�=G�A�K�Qp�ȸ%�"|���k�\n����S����zE����L��͊J�qiB��|ب���<�������/7�vX��d>��������w����fn`�����։὘�KU%|]eÁ���"�C ozmP9�x<�x��q��~�L�T�َQ��I�f��}����SLو�~�Rlv�=��猪C�Z�L�a��l���� ��� �k*���P�S�"���u�������%�c/.&����>�>*Z��ucJ��BWt��!���:��[��b�6�����q��]/�!)���2{�	��~����,l,�+�QEM��`����V��\�szoF��k�5M�MB���# Ws�f��C8�	B�r�xf@EjL�#)��a��������U�ͨ��`��p�p�0��'��R4n_(�XJ��1���L�� \��I����IpCi�* 1��^$\�mV�n.*���賒��u�Ʌ��+�>T"���}�D�#��۰^K��0��SZ7a4���շ���?�*,��fM��s���	a���b	���F~���>��N��]i���]���T;粖<��^�Bn!6jb�����-����tb)l	�(w��G�*m�ÉO���8����{l�]�_�ŤqB<_t��C%oG U�0���c��{������6�'ܼ\�1yt>i��}-��ذmS���Q���i�V�|U���S�)���&��jD:S25+��+E���!�V:�J��R��m�4�����F3)�OTosʌe"�5��'��4�vV�
�=L;e�+���}<al���~�C�	���"p�3-5��>h?$|��۟NɅ�ʭ���x��eפ�]������t+P ݿ�%ۃ�iנ��AA�JU�m0��J�p �p+�VȹO�P�{��[��H \c���}�;M�տ��d�?e�m*����G�V#�)�o���#c\��}�r���Ԅ�z��<06�<e2j�mN܋��wS~��@c9f���FV�$�v�ϣ�)O���\�O��1�}�H��`LC ����v[��.F�{��-!��[���d.	E��!���K<�.�C�ɰ���h)�^Ʊ��鿡?e`Rv��=��x��q���{�ciu8fi��XZE_+/���Iݜ�����2DI}U���.e��G  �N�����,*1�k���BZ�HN�&�` ���w>N����pH�典�ul�&s%����1_<0<�M��L̎�����Oze)#�ӟ��#���؈�c��a���>���t+X�����%���bkl���ݒT����;pƞiF���}��V�y���x���up}����+�~�������^���uS�n�k��Kl��س�J��������^�������N�Q����zpz"�;Sd��X�N`���������h��hS�XZ��6+]o���l��'����v���X<sݐn��R�O&���ߤ�Ku�n�3 ���k>������	��%��i��z���S}lbA�yL�G��q���ze�?1��*�����b�\���Z��7���H�u�ϦHj�~K6E��̛j-�]Ԥ��>cJ�����w����oݨ%Oxz3I�|�*d!��n�{/���~��FoW�W6<	�j�!��]�Փ��_n4Fv�W�ǇIL%�����b!�J;�D����L��ǽ�w�U���FsBTQ�`���˥w�P�Cs�y��\}ש�P��RN.�S�D�F}��	�8�4�bv��y(�	��'�	5�9�eC�O8-�$���wM�hYd��=d(ёǥ}ߛO��)��o_ߢ4k�\��U�kڃ]x>��i{>~4N�8&��S_��#�8��T�Ab�)����SG.�S��1վd7�⯵���`$���a񺝞ٵ�c����k"��3�[}=_�]���c�rO�YsP0���(N�>��3+���)���ՉY![�L|��{�c�Z ;�0K��o|lR9��T�k�μ:׽�H͍�P�!�q��|R���=�؝4�p��El����x>���C�büX��㺄p7�IL��sC�6�12#W 9�L_o���z���w���cB>��&�����F���[�6��"��z����O}�Z�b��2֋��yp7zo̮��z_�ه�P�L.�vX--J��E��@�a����3���m�s�*���5ýw��d�ě�A%��*.ܿ�=�
���jư��ʣhm��KMZ`&Zo���@g��.��}�=37��U�>sғI�)�����Yw�������^�3�֩��5���f��U�������im�'��=	�*9�B?���E�9�pM�]��_���bFAw��.@y�����ǆ���v����-4�H8�F��(�]$��xlԧ��T>���I��X��4�X��{*O"n_�^��sl2��¾�6����Z���MS,ED����ݨ`��B1�O"���QSC�KC��`�w��I-ߖf�kk�&��@5��Ȟ���X
�/�&�8r���l�x�t΃��1�7_A���s;��1S퇍�C��ȵ��F��B1q[MҸ�3����=-Ό�!I��D%�zP�}��Mڱ��w/GL����F�+'	gB�SrINE36Nو:����d��'m�&X~�?<�]z�_�lk������P� &�kA
R�?
��=�4��	���j����h����8��_Ͷ'�4�k���I��8�R����S�L�tU������kM3~�4(��d��v$������7��T�6�.�=&'P���{��E�H�@�Ы<��~�,g��A�29-.�=͑	�cX��z��]�4:0~���~+��Q���	SG�����^i|��7rU������9S�N�0S̔�45���;���.<qcQ�'r��΍�K��԰��zV�������*��Z�u�e��Mðy6w$Y�?7I'�n�A�������E�x��}p;�l�ϋ�x��Ld���� �{F� ��O�ʯ��z����G��`�� lr�{Џ�	7��K�ӎ��02������$]/t��{�֏]Ј��M�.���D3� �D�@�.�W�ŀƔ��*���{���5���Уows͜i1���ݮ�)JY~���6�)��/̸1��@2!�W;ER�hD�lՐS�ɡ�&L�j���Q*D��C�y��,�кj,���G�!XK����51m�(�(j?e��� ����W�}m���JqbJ�S٥d�R��/^�甓:a{���s��n�#d!nE�ĩ�]��B�
\/LT�cɮ������>���Y��{�H�pZ���h��f���=nA��1�v�_b�b������GPy�n����PUq���Vd�x�!tX��L/=4=���rJ~溊:ӑ�o^WY�z?Un7��z�An�K��>G����Ex;�Н�E	8�&��s��~cנ/lЃ	��k��;���=6�:xO��~/�ZX��8���m��SfTlz����$[��]�2tj���j��v(�w�^8������6�#�&��t�Q�����>.%�,"NZ��!�Ϩzt�^���\Z��K&nf�B�0ɔ㥄�(ޣ���$���"L����P��8��<t(��J0,�ܶ?��;��A�3��59�.ߣ1�����Y�$B��.qO�ڥK���Y�7�E�3V��/�N[S�ȁإy���&��Z~ ��f�{3�c��� M�pw�n���ȸ:�J���|�~q��^�װ'�PkQG7��;y���t"��q.Ҹ�p�02��  ��IDAT���~ FFX�v�Tו�N���;e3�SG�Z���cz$�B��!H�g����c�
6Ps���!D�\\��!�҇�o�,&I�ɻ�tE.*/[К̄!����	(�k��&��ǃ����H3��;݇��.�a��y,�?������"VMH�����MIT���CmԤMĶ�Tx���m����௎
��s�K
���cN���}��=���� ��C��cα3�Y��N$^Y��\c�{��`Q��9��5fs���!JT�d7|y�߂!� T���?	V"�f5�����7����"���˥����B�9��y���$�N�w{Q��4�R}x���A+*��q�s��{��1�<���R���^����9Ox��P�L>r4� Q����.��[+;3n�κ�3G�C�F�"yE�}��U�WEV	m�.�u�E�H}��:�6Ğ�^���ʭ������I�h:��H-�onr<,l3��̖%U�������ę3构q l��,��j��h%��M7_`=�W������	�Q@f����{FFzO��I�2Ә��2Q�:���s��#����h=����O:j��I���Z�z��m�����>K3S:�>8��e��G�#�
!�z7�[�o�k������P�rז�[R ��}��I��|���U�Yd�[���w������ ���6$����ӏ��[Ъ�������ߛ*"�"sX�EYG:On�E�郦�P"V�0x��5���~���}��W������C�0tQ�XY���g�������S�%���;����iԗXK����=���oNuTREfR@ΰ�����A�8��^B�L����R8��	���5����a~Z��>�8��Y�(.RI"G{[�{R�&{X�BV�=��4ޖ�E�y�];fasO��&��x�>o�<�2�ه����2�{�{�V�%�H'eA{�%��}��8�q}���=�|@��}�עnh��T/WfU�z��d]k��R���3�I�ϏN�1u���N`���I�/�$�v}�N������D�>�s�+ �&�~T�PܽA�=.��k�٘S4��jDP���.�%P��k��Ut�,q��I�ӹ��@�Q�:��	3��v'JLbq:ÇI@���xe��e����q��C�s�-o+�ʤ�[���.�N������Tӿ��������Z������n"~�*(�w�O7D�� ��{��*�%No"���=ߕ�=6�$^�E�����t��ڮc�{�m= s�񅪨nd2A��~�&]%{��l"�V����%����sm��n%]���}9���=TA���7�j���٢�O��-R���_�4p�y��d�t���0XH�S��.<3�⾆�����ہ_�e�y۠{�}Ϸ��{t�E�����}�����GZ���Q��0X���o ��A�7C{�J�]E"?�Bj��S�W{�JИVMU��Ҁ���Y`��)U�]��;Z�h,!��Nz�̢Q�# X��ٹ'u���\c/<U�;�j�A3�^b<�c��ox!�:p����C��exo,��d><��&s��q�T��<	�%c`�bF gss��Z)�زD�ObN���"�R�����������Yq?�����Ӏ޼݂�{*�G�f�M���,nB��u8�bY|/��1^g^���B�`�*F'��-����e�O�p䵛d�r���$��#��F\G)���-N4���T�9��F��t�s��u�N�ֶ�4����y,���U]��٤�8�EzH	�3�_������3��R�I�*%��"k�~�����g��n��X�����OټTCj/�6���$7rsŔ���P����uyн�i����6o�_��W_U�$�u�ɛ/�BϜȥ�x9�4�"gP�E���9�(&^�}�t�W iZ��ɴ�]�ى�dUn�=��d̘JD#(=W�%m2�Ȑ�ϋ�86�8�P�)�e�ۜ:�T~�2�ԝO4?l��v��3 �������V�q �&-eI�ҳ�����ۛ��En��PG1��F մ�ˇ-�~��r�5�(�� Ư�&e�Ĥ�!��xMd�?��c\���-�|8f�&D-�C�r�zpg����ChGqQ���Y4(�Ϗ��A��Pħϟ4Eӑ�V�214�{e-�i�Sgp�B]Kt_~��i8,�`�/�=/��ܐ�i����UE6�ʲ�'>��k�6BpY��"G�7Ҹ�J�oS��ڰ^3a�	I5���iQ.���M|�*����9q3^��7�ii�`,\�^|��s�}�7T&�z�,�j��6�v�bĚ��n�o��Ϥ�V�
���3ES�*�%gS��_ߦ?��n�Hk��^�a�8*�A<��jx���>����z�����7N�����c�1|w��g�?W�,��]3�iI�kv��s&�_�9��~؉- ��xϡ���T;/��Ӑ�� �$�ǝbd��V���<�	O�!���<R6S��GP�Pj�M^�bAc|ũ�]%�!�^�On�I~���G��)���1K F��a��A��R���:6EEH���o?�����X�K����U<�l����{�&p�J�IG� :������!��K�j�Aɕ�9ѡ+-C=T���{m����e|���@�F��2�r�\��Gubj4��M)b8-tg�C�/�e~(��]rH[��6#]$'�*#�M�gV�I���s�X*�������+�^JWkm�����=�4WP�L4�Yq|�~m���1��4�U����C�7���&!�����+�L\kp)h������H�|�_%�Miπ�㆒�ã�\�p�`����Ė��
G�J��/x�4���ο�[����2�w�⟕��4�i^�q[h�eq�X���x��58~^��T=	e�tOh�@�C�ng��Η>()y����3O0�Ud���:������e˴h�6��Q8g�Kn.�}�Ic![���p��I��t:�[Ui̱��Eb���[�;���6��� �`^��^�I� �_:v�*��r�'����M����
�p8_��V��wR�Bf��X���h6����Uv��<�,�jP۳j�I��SW]�E2u���Uk^�c�>X�x�ƽ�6�w�d/�z(��f�;�*�3�z����t���n�P������̀��4V&N2H�"q�t�-D$�^����V�y Q�/�jp̢3�}�8ܤ�`�Ι(t'"�b�A5�=Uyм.k6jo�A�[m��0�+p%��=�:��Ԡ�5�a�뫔���W�M��^��&�T�kv���BI���d�K� ��˳�O�)o���)MB��W�';��AYj�u]��.��@-���ށt]S���A�3=Ɔ@���~��c�l�@|~�8QF8dp�_�Ƃ��,�Nq���1� ��\�������9z��39Eǒg��lA�[��M�Ͽ���q�\���XRpj���N���eI<u@�#kj�PA�o诵$�:9�ީiP���tj/�"瓲l����Fr�].]]P[F��4�Ϛ����u��^�f��$/rugP�'^'XԔ���8lp$�B1�}6��3���v
�_70�&��<�r,v.g^MTc�8rdp�5��qe�,7�_X����b���@�l�(�����S+SG.nm��s�F��D|v�K�)�n/4����g��S
�X]�M�j���f����n��hN�9�Vշe�dfT㭗O�cI����J����H[�������Qݔ�]��6��+>�N�}��n��k�d�^�#�;�c��[��cS��$��f�{X,{Uhշz�o��T���H|�����_"=�-F����^�T�3R�,Ъ�>@�	�� �AJ@�� �\В%���� ���݋��� M	���ৗ��g�W���xݾ	�4�õl9y<)^B	=����H�3X�i���@�]\+o��)N�I\/��u`������膚i���j��޽��#���'��d��.Ӿ��KþډSP��Ģ��U�t��-Ɨ�����L��ɲ�F���T���mv %s���� �.P�LU�=y�]C�p�T/4��P�1!�� ���4����w��^�-�_2<f�J�p���&}�e�T��z ,��:��z�m�Z�a��/F����F���x����1�s���k���Ag���gcL1ǉZ�ދ�l^sv�o2�.$���8�5����7=�����Ϛ���Ж�U��H@w �~<.�B��V��͂䉸�\p�:~�.fQyj��O�X���t���o�z� 4�� ���ł&�@����Ʃ�U�-�1g���G�����1��t��F״�'8J>7i>�Qx|$Q�J�K��9�l�PK�0�&Jh��߹�n���Xx.˝Ӵ�&���gE B%
Y[���'2�7o��T�DiR 7U3��J<�����*�uo�'�3��qXj���)2��uv�=�rqW�b��i�X�\	%7����a�����)�˕�YA5<b�?��E>�����0b<�S�ڎ��j�QKYV;Q���(kn��X���9H�.���"�Y��kЯ�A�^2uA�C�W��
��!�f@$U	���$�x��vKY�ػkr8����鑭�<������=�o�T�J�&����u¹6��\�R��f��?��&ʋ�S��^+�pA0Zf��5������R�%��x�+4����2`䥃��&�_�6���<Ź�i�0�_wM9��7 ����b�rOy�����/�)���ܘ�5���sR��Φ��Ά�AԜ��P1,opv!r1����R��0km��(/K#d����=D	�&��&>_l��������xN+�L�|�Y�r����m5�[t`	� ������O?���xt�q�;;�I��~�F܏?�T~��/�V6�>R��|f�EY6�>������t�z��z����u��]�Oݽ�R~�2E����Z ���K�l�Qٰ�I�y�����a`��`�Rv�����:�Y#�9��_5�i>�${*�K���ƽ}�was���s�У�YMމ}�5��lYtߨ=��F��lχ×�V<�Q�=�Z�=�)�@C%L�IQ4?ڇT)�w~{ 2�f��{n.����WM~|q�켴)�_}��͎��jm����\�Γ�TVU���R{�I����2=�7���h2'E�R���eZ'�[6�v���3�K�Y��˩ ��^Ԅ��F��@��P]
����m����`����@ ş#� �n���E�n�3�<�s����vBʥ�ׯ��UZݺT�j����%������=]��>�5dSg���Ɵ��v"����O��H$~���K���#����В�8�E#EUu��@S,�����I�wI��zD�H����<"{��n���K��pannC��Q3�c�/�M��y���쭾E�j���X��書�����FLCJJ\���.�P����l؎F� Cܫ���y�ۉF�s���p9�[���dw��bMN��]��c��T�)(Z���)Y������0�{W�ik�Wһ�"��b׫*��"J�)Ӷ<U֜��d��Q�:�����'��;R{8�%g�s(�&�s{^$�s�^ԁ��:���*_8�{�:�n2sk�!���:���43*d���{-�b&�']���X�Mvz�m�h�.x�4����H'5~�Pە�0��5����}����{�,p�~�1���\/�OU�Sx[��U��#��g�#ɓq�g!p���dMuEq̅����x��q;����q�G�tU��Pz�CR<����m1"2rj��:+�ł\�j�ԩQ����ny���Ƒ�!��:kR��BMI��IVG_��^^�z3��Q��|���1.�_�����.���x�T�Rn�&-����M�B��Ïq��Ui*'b��\�������Q!�K���E�qрE��*Jk���%��c��v�Y��0w�E4y�b&�bU��¸�[�+�긝���E>��2��ܜ��
���2�����:�bFض�NGr�q���M�[$HRD���C�ȣ���q*^1
n�>�ױ),0��~Q����z.�E �L�[g߄Ae3öWz�}N菮��Ҭ iN�a)��ئ:(��AT�J��ƞSF}.%����I��1yY�l��K�(����y���V���g)-�K����>�
'u�w��C<�&�xB%���q�.�M��rC�ի��ȬHx,DC��8=&���M�M���(���2�h�,g�;�⨅��]yI���{�W?蘙F��#2Hsb
�nc�RἚX����|�b�$�D�����������C�E�.�V���#���=C��2h�OԽ�� ��!<s:��wG>�ė#mq~3��%}B5!_�D�tg����7۽��r�4�Q|SD*g��
��3�M��q����ؤ�^"¹P5��L@#�q��y4xv� u]F.����d�.n^���b�1ԩ�{��UB;a��	�U�?���@�G��!�z.<b�~;�i�-�6�L���+���b�{��g:~�#!��	��
w5W+1=�Z�Fg���	!W�K؎�I�����~)�_�zB��t7�3����]�n��Y��>:�X06�/8�Wڇ����TV5���V���&�����Z��'����5�x�F>����K�K��UEt���m �`,r������lH���t٘���G����m��eAj�Q�>S�|�1t���j8���j����t�)qG�I�~ئ^F8���8���15q�(q[U��^|���OS|Ϗ?|�.��xhhP���F�Ψt �O��=�>	F	BD��)���T�Ksh�r�8qt��6���ȧ���6׍�;Rl���8Dҏ�r��` ��A��3�F��ad`H9ǇT��.jJ��>J㔢�t*q�V[�S���a
skH��?��:݄3!A��:��קa�1f�Ӏ���f�gCٜ�72�o�{�{C��n1�b��u��QH�H��b���KNw���x�=6�ջ��h��X�5��64���p8��P��b,%�ʵu˥	�|�yb_��7�QҔ�L��i/>F�"���K��D�2�p�/]U�/I5���U,��l�دړZD���ìt�E����Z�ٻ���#_Z�O����͈ʘ�`�Cm��E�7JD�q ����EG�iΛ-�2��� y�R��[q�Fc�@�uR=%����؜��������7ٻ%m�|���4��#Jp7/��}
(ț��/��P��zu�!����~�����ϱ8!�3���nd��ėc69�=���b�$ҪgU�W�k����!��yC,���)^�ϴ�'�Ց#*��戔��F�l�؆��!���ځ�3^�+�v��xm�˯,�mQ�Ku���xG#r��ԟmOJ�ǡ*iݤq)�E+:�hKn#Ү]W\o�g��dHQ�CD
����.x�0�fv�Z���y*\C#��4'��x���H����	��ރ��#��P�Z�lA����掛 nl4��ب��,�g!w.�=j��|r��כ#����9|t˹��\��+(
(��'s��}�deT<}8"4�%��'7[X5.��E�=f���ڷ]Dj������ x��
�����TzHМt���x��:��]�u�ޘ�-ʓ�t=[��1�Ϯ�1��DǦ*�0��s�QX�چZ�m��Tg7)�4�N�T�+1ψ�o�ݽ�XY�?
���9���p�zѻ\,&,��(��9;1��x���<��B���.��:�$,\$�2Y����hWV�� �1�{&<I�3"�R�A���bӓL��l���wq!��`q*"�HS%~��yI�n�������O�o4����%뒚��G��v��Oc�0���\0XU� ���x�Ւb����#N����@������EG��Tih6n$0U�5�k)����i��#���O[\�ް_��h<�
&�䭶R|	�Z�0�\o׌�L�_f��I#T�	�wӂ�T�"�x�u��m��T�:�v�1P�=a��Ep�Z����V2i�V	�{��q�ZcZ���!]�g�@1i[EY�H�"w}��7�5أb�G��iN�+������D��?y��kg�犏YN�i��T�� �;%�peRم0H�� �"�
���aR��[����c/؈��fK]:	���N���!��~��>����\a4H��M�>���ؔ��,o���w�q)�w0��f�ӆ���Ť�Q�%�b��dt�*n����ES�[� p�,����7�J�{�60,��3=&m.R/�d�Y��e�qY<�kz����F��sMo�0�j����~ۮ�#goVw��0S�}\G\P�8η��� ��"���8�T��w����v�^�������ޒƧ�na@���x�Y����{����=v�yFu�ӡỐ�9c�u���Ң0j��P_6Q�Q��]b~M���4�tC�� �}�1M<p=�=Vj�^��2�ل��4����ޘjG1�v��m�Sk���u�T2��\�������J?0����!�/�ע�T}V���3�~|\%�z5智+4���,T\X�������W�"����JjD>����|0��O�֜�b��ԕhHQ {�N����Jx������0�2���CL�m�4n��9�������$!e��Pm��5@��;�<Wj�S�Vt�6q��QRͲ�wgQ�]�lZ�5��� =+d��<���M���Gn Ec<����Z��#����Y�A�F�rM��Y��jG�k��G�jޫ�k��v��G/Lz��xn��\`�kQ 0C�%Sv���M�U�|����c�9�����F�tϖ^;�0��{Q�lHq�WuW��1��}��Ga�l�ը���B�B�x�b'�(�f�D�U���1��@���c��=����p����+q�9qP^�UtAgY���䗛!����d�^���tO'�;V ��� f�k-�i'`A�P�Z�Y�ON�׈"Ӷ�dc�L�%��=տ�3*�1λ��|�'��ִ̍���R}b�^�]���M-�(��$�m#^/�n���t�r��C`J0Z,L�W&\�)�%��JW�G�A���D���T�P=z�&��!�������W���@�h7��X�
���v/9��������p��|n\�P
#K\w>"R�7谰E3������=�7mBwO-�ȃ�t>���Fy�S!� Z{&C���L�|�齎��i䐨/����"$U�Y����3�����xT�a�?&�� ����-�����^S/��5�@
�5�j�0dt�h�gJ�W�_���j���.w��3K�*����K�+�{�F��8b�V�"7�圆�:
����G����	5Z|u�����g�ܢZ�'�O��]��"�ahF� [�=f搆����#�'Z�o�#-Md�*��G��p��Ӎ
R\?A��iD[9I�$�"��[����eڿ<1��x�c�9�֛��2�BG�nѢ2	��&s1�r�����̋{".�~ࠍ Z�B�̂G%�ՠ�\m5�!g�����g{����4PQ���^&�	��n��{3�k=(�J�ǄoĸDUu�L�R�����#����#a/B7{���^�*�V���-k7�� t)���j�R@��O(�˛�*uI(��hV-MՕQ����2^޹/�;~Wj:�G4l��nv.�������_o�c��X/)1�h�8��`�#��;���3�i+�T��bl��?)����㘱����J�&S��yK�]9v���*�&N*����e�N�A���z��K�}�~�ߜ� #���k�߉��h}��z���m�cP�=����uk�rܲ���>+�5�Q�N'M,�`c�A=�7�훫�̖�5�f�ĝ��V�b��r9Ĺ��FѷT%)��D��[⥶��cj_�8�hY�%�np%��{QO��EE�=����QXt��Ţ>��Ӑ�ct������Ά���T��T�$Rc�{.�B�FA��q��t��
�
q�ٶE<Z~KQ�hL��HF*䉞�k�L��J#�eH�����LV��f��CO�4C��Q��.����M���Q�#GS�
Et��"1�{r����Z��x�"H���,Cڕ���p]
+���Ǜ�����O�6{�4ε�d����N�[R�zeF��T����EE��O4��!�4�����6b!^J5�{5C��#�d��3�̼�������ib&��&�$���_8읱��kD��H����:�6֟&��ʐ�]���=����vkBa�׵Tc�jM˷1i�U�hU����|��b/��Ŏ�-��k��@e*[��u�C]�D�lU='���}Y|Ԗ�?�F�����ڜw�Q�?q��L�vU!�ѠN�4�%�~ȋ��/eh�������v�P�(%��Q�"���h,E�Z�����rtH;����Z|�=���t.>����S!A��.fD�+�*�ָt
�"ƬH�;�Cr*	w�}o���Y���n��
��b�����x��Um͓R�t%�
��%�Ʀ����A����� ��RQ�:[�q�%�r��"+s��q�7�.֪��Z+5B���s�G���Ql��i�^xN"�S~U!�����k�����K�4F4i�gj��;-R}�T�Ņ��։E ffu��;�R�C�_��MF�c5��+�3S�
 �b��� ��%=���\�VS�`�DC����Y�!��Pä!t�9Y��0pVW�����?iY)!�}�����.��J�U-fQ4��۔U�n��v������o��I�����1P��>YOcZ�b��i<��[K��`){�v��/F�g�M	�O^�SGeWi��tGQ�aH���Q몍��P�=��A�k�ۭ�����+e�.+|KIɱ�iQ>׊�0Re8&ٷ���̇�@L���Mek�Z�`�t��&��-�<G��zӺuiR`S�zu��;�J�5Rfij�wu-Ɍ�`����VQ�J�6�5F�����tV��I�Ѻ�Οm)C*i�Pt�����6�!�'�?;��y��ȹ�V�E�OO��<�`�b�"ϕ�ٹ��zLc�%��Nc�[���	~���(�RA�#P���р��0
��A�]��#�^%�la���_O� �o!l�; 6uc�Q���Ɛ�<9AƲ4s���6-��.�(�,�Z\S��RP�>)��
��w���b���?��il����Y��b��hѲ2�4�ջ�S�j��6��\�Pz�=~y	��E�L��=ON�G`��?�@`92�~�tK�����`�n�B�Y�M*=đ�]5�7��t��?�g�rArc�� j�ӚOv����4a(
@o<�3�MK�xȔφ�Y^���|!P��P���f��+���Y����*�⚖���\Y�ݶ��aX%*A<0"I:�5&W#�!�����Nfe윘����HqUl�� �PU����e�d:���#K���h�=��_�vP�ԟ"J<����4Gh��󪢌��E]����A���Ǡ�qr�C����*�qO =�C	����zd 1d�w�a���`M�ym��g��4�د�<�M�K5#�}�in�QI~�I����YMɑ~�|����u�"�	�2fc��*�Lxh�D��*���{�bl?|]=6:��q�}h�#��\�[ո�^7ʘXM�=�Q�huʩ�f�E*�P�KG�?*��ڊ�t�aa��!������Z@��ϐ�i?I��`��|�8�X��\��nP?S��ȸF���W �A��h�y]�9���;�9*�9��.����5���s��^ڝ���g�%��"+���D axb]�:�u%�9�ms�<Ε����KyAҪ\�m�1���)b�[�*\����H��Q��3���kZ�_�L@*���%���*ve]��n�(9y8{�������6�] �n婳�������LS��w��A>FpfH\�(�>���M�1��~�8t���]g�_Y�[��WR��s�#r傒��.t#F��7_l�zqi|O(�mN�bڿgt�jn�ⶸ���0�j~����aL��(`V䏾}e�1\kr��}�(�ef5F��>�K��c�\~j�M{ �XF�ɚT� w�:��U�э�8��~g��{�J��ߏ�8ztd�n�&0y���S؛�ӏ���аYXؠ�A��
P���5��W�gbj���^�*�ö0̡�
��pocCG�ŞC����G����q�/T��zV�b��"�&�T����횿��ƦȢGH~ 7c-n�Ԯ�;1� b��ո!�����P��0Nq���]4I�U����:!�.q�e ԂGd4�W�a��݌�]sJI�5F���&,m�[�����*�Ltw��^(��u����>6]>��O����jjp�J%/v�����*b��BG�fEة�����̏�BT�D��F�,��c��{�"��BX��Rt��1��'���}�'����g�)�jUJF��L��I��6�X���zl�;��?ӽ�� Χg��d&mй�3�-��R���`v��$Ak������,R�^'��撲a�ZI�J7�P,6��wT�
7(�71rz����ܲ��[Kt�`;6�suT��/[�AZKQ
���$��s�7L1X_��u�����C�%r���׬���V
��>�*��c�Ɗ���j@�۟xCq��r�W�kaHQ,�1�Tp�� /O�5�O��x؎���٧K��N2��؀7��]WG��(��Tx�~�r3Bcy���b�ޓ�uM1��:O(�S����9n�rn9�$v��`}��s@�"۝	��]���m���)Y���Q�u"��&(;=�ӯ��R�?���Ջ�>�G������>~��H���5y��ً���5��C�7�o���t���9�����U`��-�~�ɶ۹=�"��r�B]�9ڬxq̈́�u��K��*����9�b`y�8/�/���ð6ƍ���b@⺿/��1�wռu�X��N�u�������'XȄ�.��
�L�(�R+�U�����G�����1��C�Ȕ�N_ �l�H��V�d�s��ZF�#gjT���_1���X��\y�����`6�ǵ��&>��L���b�z�q���%�0��H�lI���3T��|��z�x/e�թAD�Q���K�F���C�[v|CbB�Ȝ8_ø������zT���J���젇�rU��I�"���Շ��,��y�yDF���x�BC:o�eݜ��?!�s�8����0�QRܭ�X3H�����8�I��ݜ�V��T(R��00>�Rۄ�4Y�&�օ�:%e��-����.�B�"�E���g��x�+�Ό�c
��"7�Q틞=c��7G>����ǆ�
cs/E�I�h=^��ub�Զ��DGˊz_U�6Í{���\?z�Ȋ���z�X��Ѩ��|�7���E�'�]F� ���E�0$��������ߌ�*"�W�p�<�:�ѫ.R��,÷��V�d�a���s9~�1�������A#�R��I���!�~��T�MWٛ��ɬv�����Q�n_�^�����+nk5�� ���X.� 3���n� ��Y�2��M�ƇjH��[�x���D�5��'U by�޾(���>z�;F���:�[�r�:"��xzu�ġ*��s��0�l
h0�a�x��ɐ�ۿ�!�.�)RJ�l�!�Ȳ��cbD�l�\�H��Érf�3��,7B q-Ðn絎���g��?+_|�y�h
j�j/���
�������B�Y�]F���34J�'�%ƪf��*U�K�ԭ�)�*�t���:����/�3S�eɓ���*á�uL'آG�͞�񬍓��E�0�[`=�f�a������Fd#���b:H�����A��=�7fƗ���X�ZL�q�H8�/���=7�|O��U814N��Q\�!0��Q�Z�,?��$n\��������,>�1�x�*U�IDj��$�YY�1f�7��k�ݶ��gV� �ŗ�>E����8�O>�����G�E��o��v3���z���j��X��Kc��U4�#r�W��Y;�ʇ�����䨑�TcagEI��Z����V�!7=�ڛ`O�ș��ۈ|����-����.+QY�xވ�^��{�Oh�fZ�M6�8NŤ��0�FąBJ�h�B֢J�{�=�@��@��Zn(O�Ņ4��4Lg�⭳GSD'����M���[���+)�S���#���Z�H�u��WQ�����R}ިU�k��9�wM���b���F�hT�%��{c���������]J�A��Y�1��H1
Og<Τ��b�����6���;hin�m8��#�����y:"m?�}b�*r`سǌԶYv����3p��g\�C�Fj�ZE����&3T"����L��CK�3�4���&�s|I�K{�W�m;�c=B�@�N�(�_Fu��*�kA�l8N�wNѝk�m�s��y�y��~sԐA	;�Z�k#GÛ�H�&����M���������W�����џ�w���wk)���[=�񖩥/�m��!�͈Uf4�����!"N�kR�'�o!���EvD����=͎J��X,��Rq<��j���$2�hIS��0V%��e�.$��Hr��G�ؔ��e͛��Ѱ1,W�*�*��v ZI��s�"�3B
�]y�s�d�9�9�8C	��B_�~U`�G�i�cl�(�D��G`Dq��Aϧ�xWGq���.�,�x�T��X��ɧ�s�8�qG�v�P{ū���ciLh�v]D�ky����f�^�1$q��7�4��;�}T��\#ϧ���1C�x�Z���oN��#Z �hQ�vj��R���!�T:'���W���6�\�H��j\Qz��5�+�R�jV�G0K��O��1��9)��|ּ*�m�yqm���s��l���d�=��b������k�sٰsME!������S2�v���i?���DFu-��7skL�)|kҎ���sW��4�	:�����s�S����;	+��	��:t�K92���Srn���z��nN��^΅�<f�ex�����l{�c�%�v	QL�z���aC�E�E���I����F��-�F��k��쮣)'��������{f^c<����xs�F�w����9f�GFpc_+���E�����(Nݟ8n9",��14��<u�]dl�UY����	!t��ɛ{���,��an`�>�fzmdd�u�J��}n����ê�h�8Ҙ�e9��a�$\v�X;5"�۔�R��
_C�!��0�#����߶�0+bZ3[1��c��tMD�\�S@^�Ͽ�"DU(}	�Q:w8�I�-�����Sߦt�� )��V�Pf�o�%�@%�nQ���Y,��,�T)9;0���1*0��=����E1�5�#)i�tp}�e�QJ:��ݹ%4����t?zAՊ�>2u�Z#�**�)�Ǎ��&�1��'�ψ��A����7^���0}:�811�4%%�ZZ�Zշ�(��K�@Q~:3x���l}T�`��]�e��I��o
%c�#�f����~v��F�Cu6���t���f�ɑ�R�z�A`�6���6-�C���<wG�����~c*����r�Sbp�<Iͽ�F}��j���b.� �A���FʅG@���̭�5$yȪ�}q�Jӭ��M�(V0C�ǖ�]y_8O�z�SgQ��<��iM���~
C���h�Pd��$t3翳��XqlY�N��o��H��f@Sە�&�$�'_�lL[��N���X��U~��b��ߥf���L03�={��J���z�3���,�ͩ	1g�jL�X�^���������oǊ�k���F�%K�l��uf�O��ZϽ�xj��|aR��n�޽�}����e��D�W��,�0!E�6��&���l��Y,��u����p�(��FR!RZ�MF�����!��19�v�'��宖��9h�"#V,��~��NA5j΢L��{�g�u��7C�,�Y̢d��L��9���i͋��Ϟ���)���{�5מ��u�@���-�Aao]k{cF�p����l��_h�Q�¹����y ��C��وn:�L�)72�mhmB�����"�#�PF��5.uMb�\�<!�q/?��siL\�aX�/�q�~�i���(���������$ֶj��2����H�RG�G����#�#�ߌ3^y]��u�P������y��ߨ���#�*F���Q�%u�s-�{�}�Ԭ�"zҔ6b�_t>6O��^��%�k�"�����e���"/���V�r��)Ys� v�~a�Z/���-�]��6�iD]�O���u3/�]t:��=��~�)���J4��.��b1)�`��>%զ����\,1�$:�п�{:�������q-e���Jy�E�ݤ˅��^��{�1�Y��"=HvܰBʛ�^J��מY��+\WU�!�|�ѳ�4��يF^�?�A�X�&$�[U�9?�Ƶ�,�l�V-���R/+�ہ�|+&��.������ǿX_��0�f�pNW:ɘw����������䀻��!��s�n7g?�Ϗ�D��O?��gB�g�kQ��*��.|��>q:eO���!fh!b=�Ё�x�6�*rͭ���5�4��ocr@F�����crfE*�D�6��d��9�2�*�y��MD����c*��.�$�#��]~S#Ns�B��\ǻ���R�*�6~�Aָ�OL�hG�~����F�n�&n8���m�# پ��]ҨN3'�F�R(x�=�ܐ�2�-��Ze�h�fXP#�'��jPCZ#Ҷ�^1=��݅JC����r��P��?چJ�3"�C��t]�X4m��-qQ�1�S'�h��[�4�qqM��s�Q���H�ZU�����e���f�\��-�1�FT��H��l��� �*��?�k�H�v�Uo�ⰻ497X�rϐ�1���e���w)�|I��5��#f	���<k�֢~��#!c[�ٌ�?������#x�����~�*��6�Yت�/��~��7��}�)��M/_���,��������!u	*���k��ǟ�w�}W�����Q�X�0z�#蠞�n���4҆��߶�����_�X��p�@���V�h�t�S�v�sD�f��Ԉ�U��yg�h*drˈ�w	��2�D%��& 2ѹ�k�\I�����CHT?��d-iHT��P`���)���/�e��N��Y��5"e p�ʔ��H�nn-���qF�Ci�O�xV�t�گ�OQۦֈ��W����}������E"�&0�#�R�f�2A�YR��I�Ե���!�G	l��ז�����,U������]��x6���^dbbMA~��co�����-N��e������<�!fZ�ac�Zz�ƫ�=�ړ���;e�x����^~�S��Tٰ���W��%@���	�"F>3btj�����" gʔ�S)�4�q�@Ȇq��_8]Rs���?g���Xޤ��8:��H[]��u��L���L���>R_�aP��q�����w׻r�g?��ry�BS�s�;��9�-d40>��%"ݟ�I�)�JX�X�Q�ߢB�*8(1�繖.W�g�q��������lǉ����I�p��̸�V�u��	p�?#��3�*�l\��9�V�;�����y��T1�4r����*�ߨ���:�aDb���~X�UU��ΐ֌����L[d�����J���e���T���	+1B?"Zl?k�I-�i�l-�AQ�(C3�Ȣj<p$��Lk׵n*�ox�7�HYawʍ!lå���Q�R���Ðj�X�H�7�M^��KP+��s��� �]S%��W"
?�b�'�22�!���X	�R�q%8����I�x�°t`�Zf��R��=�Ǯz��pԽ��,�° E���fHM�	��3���3\+`�A{ꚬ�:Ud
G��/?����O�.�ѝ�h���)`�p�f:6�{E�B�#�hup8D����b���l��L�
cX?�p�A=px�b]!���Sh ��1��_�`ǋpQ��/!��9��c����f�.ځ�����,91���Yu^�`�<���fAA˪���,;B%���?A��+�a%�u�U�9⡝���:vP'�L��Ei���u2�֙0��ua[tpp5[���J8�#��ΠVL�v&��&����D�{`����faV)�]���'1ӎ�)+n<;fYX(Jiz�V2Q�ww���%�<k���0�b��!�ڈ40���!�Ξ=St��~��W�\Шd��y2jTD�p`���R�xđ}�_�׈T��RQ�H{���Fb�ӆ��ōj��y�E��������ѯ1<o<�;ص-�O�<���m�.�K*7yl��$�cS�(���8��-���T0R�~��t�����(j�F��8�2���E3�Uq���}��q5��Xܺ���w��}Q����-��2R;��ݴ���K; ��/?Ә"��:x���kn4ڛaH1�.�^�FJ�0�5
����.i,]d,2�Kp���82�q�j�m�p���pU|�ڜ�U���1����JF�Z?����#8��A�:�T��R�LݳBX|���������o�}U�8��]��.?�+O&��R���K���_����OF��Z�6m��{ѯ�-�j�I`>��!��lW�:Ŕ���*=�O���9�&8��0�B�?��R+�A��"N+�������=��	r,�X��F�R4���J�nr�Z7���n#x�%��6!=e�0�㚴&W���Λ���!+�,M�5��IJ���{<ߧ%`[<).�ϛ1�1x�B���Q�ڼ����Vr����0���)>�BP`F����Fט�L6GKn�L�)�:\�v�i�Ny]�lH-��@i="�(�m�.�	��%��R[$��Au�*�h���Q����J9���6G��u~|G�6���O��l�
��`_��`��W���p�l!6.��9/�)���� 9��A�|iD_�Aǡja�X5�G�����J�5�f��o��ВU�k�ƀ@m�è�]j�1���\�2%G^���0�Uk�����:�f�{L�<1ޙ��ʍ5��|�裭�si���B��-�4��je��-�U��U���z���hχ�����\܋7\]�1�d[��7�*����N,%S|SX\�J�vf�׵')cDM�g�M�ֻ��A_hU_DsQt�墬Us�4��N�ƯN��vE}���N�۹j�wѽtU�8^Հ��_�1�|���~�Ba�1�~�(�U䧼'չ`S�h����9���J�O[Z��8��T�bʉ∧���ZII+%#�Z,�(�c�V 3��u����?㘀��s�Nu�"�I��VӒ����IBK�~��mctw�~o����GQ؁����SFMД�S
� ¾��H��)��8����"K�ɕ��x�?�~��e�)�/�c3�y���'9,Ns�t@�ևJٲ����m���H�$�w<F1k��zn��ґ���,�7�E�Mg�]�e�"jդ�M8�v��<�X�6w��=�F�{q�"�&�49��KNeVl�u�U)UX]ɷ���c�|�f���3une=�iȌ�/�wY;�y��\*N��9���E��B�J�ż�~�<R*pj���9Qqo���YԚ(���<�K ��j��n�Mq�0�仆^L���;��N�Y�+Z����5Ҳ����n�,����٭
[,��8/�qτ! ���E��`R�ƭ�ś�e_df`�4F~0.x�S��f���l�M1=s�Z�N�g8�F�̎�V\��oRg��Pr|�m���嫯��w�r��謺'QY�bK�2���#5v���ǟ�:"B;D;������+�l���o׸Ơ)Eg��Qb�2�^�W�܎�6<�5�o�H������{'>s�b�y�WICj9K��vP�5�?ѣT��ȬG�	�r	︍�t�^unžOYj�� κ�z6�,;�m��,��\�UEw��9�C��;x�?1����C#{p��W>b*��!�!ጦ�վg�k/w�[�Šy��R�ة�D��I�?�"R��x���K��S	�4�98�*���Įޕ�w�aH��T�F�5ʀ{�C�L���L���R͎�I�$4c�meշ�I7@��\J��PĪ�"RG"BD��2e�u=���s�I�H��.��5PG�\q�Q 
8�w~�Rߤ�o<���*���6"��\P�/[�X�
W������(y����YE,��co�kq3:5+��Z���F��5-hK�����P��G+�v,���~�Q�lL���j%�Ћ#RЩ~�"�I]җ/C���?��vD�Q&�|���h5���f��G�3�:��L���,�7����l�uAΙQ�&_8�j!x�>������2�ttPD���3����f��mW��D�9h�_��})����1�n�n6�������mՠ������V�������4ŷ�"~P�㍴+z4���E
��f��wHc��M�~@�4�ۅ�[,E������+�Y��b��[�1�6�JI���*��3�;���������T�D��>D���t!�)��@�S��#T�J�8�kj$�˸�fH��0PQL"��*g��K|W���c�h��-��0r�<�z�v���D��Q��S��Oʖ<�#<p�F�>3Ԕ©<0�S�P�KR{��Y�����f�5����%����(C�� ���\��j���{��Zώ�c���nxꨮ ���|�(�s8\��h�s�~)��[$
c
�j#���sf"2i�,��L*��Q����D
�zU�f1�t8�SJ��]�&Vg��jƌ���cJ(���Ԙ�O��e`q�L�"��`�:/�ǵ��4s�j��⼮Yl��Hv��4V�wz9sVm}/�fI[� wm��Z�j<�:���/��XR?��;.�=tv���;�R�As3Y]E��ZS+hlܭ�@�ń�I�D��#E����m�7
,��UD�ہ^7�c�,�w%SsM�r���%��ԧ��jU��C��4ҁNE��"����-�rH��7�9�"i,BN0��>S�"E���1]�=�ʏ�����I��C���w���6��H����T�z�����!�D��;ҟv��b�K����^<�7�����Kuv2Cٷ+cX����c��l����=����A��}�E���Q��/�^����������B�C*D�hU7�V0����A�
l���'F��b$ƒ�7yDf�x)��5��j\\��RKw�~-�������o���~�`cn>�m2��Q�M�[?me�����r.�=v���"�
��gh�Z���]n����Ұ8ڡe��3�[mh�l�	wM$�ϩ��G� �ZB��7F�uO˭q'S�<�����x^�����.L
鮕Lk���+� 3R|��p˛�g����h2���nz`p1WF_É�U�M��N��C���>f+��؍��M�<��@-`]�����6bGT�"	6��;��b�<��Q(�L�Xo~܊�_.�0�G�I��p�TuĵŦ��OU_O�ާ��sxn+��{ދ�^'�aH�����E�C�f� C)l��oK�6�R*v���&~ٌ���=Ry��CΟ"�|3f�)>��\�^�C�	F�J��V�R���>�~B+���__�����g��_~���l�i���kyP�N�����Z8�s��i�tq����Q��y�����'�.}�2~�1�H�7b�$"s��-;����$�J��~�z���]ُ~�9e#A��q>r��.�k�A^�X��{���<׌�]V��;#�G�y�b�>��{���q�/�;(gj`且�H��aulC�3�'�ߪ�Юf�c�Ac���GF�^�<�򇏮��!m�T̓F�߁�����ɔj�Y��8��V�(�Hznn�E�M��Ж�T�:~׭�����GsgЪ��M~S��g�u������R�"�]X�q�7t��u푯�|8�!!��ל�c��c�'�܁*���b���6)� �,�h#���M�o� ����"�E	�W8��������cEC���ﭰ�o�2WxL	haB�����p�u)�L~��8��@����a/�BY6vB�~��w�~[���W�O?)�~�Iy���a�ax�	��޽[�ea���|�}F���<Ρ�tٮ�� �}\��Q����~��1k�ш�e�k��g�30p�0�)3��bOrD\wz�yJSR�JWS[ޫ}T��u]��M��xL����gqe�9f����F���#�#EVM����(��+�j@0)2���$����2���Ň[#���Dv6��1B�("]��8�/� ��w�A��6Þ���49��|X�%�_��,5����3)˅4��M'�50��EV��"=�Y8�Cj�q��/_��"����Q�!�O=^��f��WE�D��b�g� z�w#�ñA.���X�$����@��i��(Ea��G��ǏH�x`�ww�D�m�RLU~RRlHG`�6<���͸|��7[���f�87<�l��S���rj��ӺVt�C�`H�7SfDh���KtH+z��5�:[��~�ڛ���)���+G憌(��et[W�����z]�w���w�bT�q�P��)�B�n�}'um��9*{&���v��~��wq�Xk��ʛ��d3���pA��������:�)�?k�Fu�ն�5��f��s�����<�$V��,Jj*�
Q�ҽV/�G��Y}6�[��1]<%1�N�!5vV]�!�P�C:�	�۱Z.)��7S,������2�E{��E���Zc�=<�5v�R���� m�q�b%���Э�w]Y�aµ|�0���/cs�Z�
�����n���XtMG_=_\� ���B@e���ZT��ٖjw�B�
����ia o"�������`�KV�=���P� ��[� �!��[c�*j����h���nf ZB�%|~��X�a�tn��g��uI����mH��v�h
��+�(��?ޫ�g�Xa���BV1���F������-��.!�c�m�AYC��*h%e�i�]��>�y�O��6�5���G�ڃ�^p;��G ��h�I�r*x��͈�M���$Ļ��)���{�D4��﴾���F�����~�Eekc����g5�QlSAqgH-�oԁ�ŸٴP�I�a��rf��_��h�05��
���N�u����.j"�)�4�v܃2*g�C_U�n�*p=}��W	�6��k�B�b^��J8��d�P�b��|�\q�t�]kEL[8@V�F�MTZ?w�dH��Qh���jL��K���Un��H]�"�A�1<2>�#. .N��
O\�EUwa$g��2-{T�'g;�E1���56<��04�C�.Q�6I�Q�%��$�E�璚���;E��=;�@��H��=�3E��j�D�|���)SO��;U��E�����Y���l�r���k5����j٬V�_C��믿N��)f�+"�!ϱ�������f�	�)
.��@b��!N�6���3�Ӄ��^Ʃ����q��6"5(�F}�NF��eu���T?�Yѯ�������)Y8�c\?�8kEP2Z�{���HD��}_�Y�yH��Aw�we�h��((�Q��'c���(��p�y�ax�n�����Ѱz��m
#�᎒����U�8**5��Ա�(���A��"��� ϐ��.p]���G�I��x.X��cX�d�0��^GWᯑ���S���30˥�u��J#�iH�$���hC;V#�bOO�S�`�c ��i4ԡx���Յ35)���,n!��W�����}8GUn��E`�
�\���J4�Z��=�|�ߣ�Y�������HU���Ű�Z�-��nu����HK�W�H�7=��a�(�E;�5�|�;F��V��Fv�?/1DMv��%(���?#�}��Щ|�I?� "�
#�s3�������(.�}�
��� pX�#,ցf|Ϥ.�Y�����ҍ��y����6�ǽB;�� �������I r�p����^m�����]F�2�V ��燓�!P�������oU\�(�ir������+�;�)�ݳg���)��fd:�Y���-�]i�&2�g���H�׼?�����'���ܰo��])�}����.�5�y��ٜܺn����v�������kd���;��h���}Z�b6�Z��0*mO���ȥ婢�7�"b�q=̅��I�޽��Z8��g9�x�p6Y��4 �?g�%�i���� GDq`t�s�Ũ�N$TĹ�������0=nț:~�'=�15x�����pA;Q�"�3N���K�<d�psUU􍶘��:���~�N���/���*��Y5�;�bRt�(>�$[䅈�_~+��y�m�g!:��?}Q>�����g��1���]֥D}Rj�i��`oOd8���T��������1�ch/�j���g�ך�~Uƭ�-��Xa�pJ�?�T�9��+D���r��I�0��0���sQ�p�/23���i\$�H�f�[^��	t�g���I�ݵ�Aj�����*���#G��NC��fԦO3C�� F��\(#�@�_����Ogk�2D=��	~��z�7(Ԩs�&ѳ�Z��FN�۱6�Êך/O�{��њj�5rP��]����хQ�.u�@[|�b}M�ۂU[ds�Ŧ����Laj#R����\��'�l�1Ń#%.ۉ�'='7q�۸كZ��%���
�I��c~�ma=f�y��hm߿1=\|`��B$�6�!)S�w�g�釒��{]�3�]�����S���ļ�ۂ�9r��@ŊyJ�uRw�H�U��2��ϊ�%�(�)`L�h���;��k�#�kQ�䩙�[��z��Aq��_�-� <E"�fSM\ģ��p.�-�f+�G$�_D1J{��{�yu�̄�J�8����1��ᜧ[�*X��WC
����}h�C	��}���O~��g�p��)�
0Fo?��PdY���}��8W\�y��^���W�b�A����Ґ&才��ms��������q���u,�-��:���F�BJm�.�?}Z�X
�,K�d�K,eB���>#�Z�b�GQM��i��କ5����P��ݎ%�Rg$'��}�z��U�S�̼w��a�#ڲv��0~a��m���}S�Z��Q���h-�����(�M�u�,
)��=ᵀCa޽���WQ)�ᩔ���mh~k�BZ�Eަ��*g8U9�:���ߞ� Y��o��z�����cl��*gB͹`�b �c�I�2�e���W]CCO����^lIu�����b	xaL�|�ȅ�tv3��������y'�8<�fvJ���a�@��~|>8�0.��>ތ�ˏ^��mE���3qa���,Z�h��[����	r�s�MF&�o焨�$<�x]�_���9����C��W��?DA���p�V���y���KS0�9��rt�}� �gk6�ZgcX�7~g��ؓ��k>�5��)�]�Y���8V	M~x8V=�
��Ұ��͛ ����mw��N��ɤ1)�:��*��0ɦZ�]ک�4'6��9�V9*/[~���������~�X	�>�NrIj�M$|��,�,�1jŐ���Y$lb�=�������:F!6�sQ�t�s�C�*Z� 
7dL+Lqu�:ra�(婎�����(���K��M��Ɉ`�s�.��-��B��IF��鄽�{�ݝ��k�%'g����(61JY����Nf��=��bn>'DIP��1�5*ˈp��ӗ��-�E
jL�aloM��[C
m�P�~�q-o��]Ch1Ez�h����E~����+��4��=�
op�f�P���{�p+rAvS7�\t/A&0n���8����7ߊ�L��~G�y��9��6�|]�؎����p0�_o�	�'84���(,m��NG��<;�j���nǪLt��
�YFq���4�=~j$٬@Z��Oc�7�ǞSe��F���Ŵ�[�Mf�XZ�v֠���<���u�T�5Z��
��p����4Y�Zo�u4�����<q�	�Q���oXF,rd�����Q��nY3nl���!���rj��۝Rt.�~�,�ʂ��V�S���q�47�-A���;ElY��lH1�BF�M)�,2p�MQ&�����_�UR�s2%ޤBQYӐ�cd�~?�B�>QfayQ�ע�nW1��tÈ.�:�+n�2�=�R(��16�5oy-)��+�eE݄�,	*w%ǳx\oܗy�E
�+�NH�q��n����2�6#�oa(����,b�M�Gډ����_��Fq�Π�[$����-`�����9@.�CP]�������F
�����\)����z%�0�?G���m�����o��pR{c�p�,؍ZC5j�I��v{�t`������8o�m��'����"A�)��J� �DjL��x���,kٍ�� �O-CQ�Swvڝ���A�;H�?� v>������
�����0���l|�گ�h{��#[�+V�r��mr��i1�>�5��4��]��1V%q�?2��E���h�Nw$U�NC�	��C�3��8zUF�4cφ���şm[��4KZ��ݲW����93�ѹ4e(�^4QӋ'���d��R䈮�0�3�i��#�,i5�N�Fb?�\E[�<�5�>wW�������$(�k洖�֚��Mx���QR��3u�fα!�s�63"B,�����sbఒ�|�RGp46^p5�Y�*��B
�]�Aw��Et��)����>	�g%/�%]U+*h8Z�w�p�p�	-��Àa�w�H���ϿG���P� �t����w-S�(�)p:�;i>W8ZEWpވ>��~����V�����$� �kP��.ڤ�a.�{�(�F�z�T�u������m��L��~�yD���֠�Y�׮����>8bme'Yp��DO�KN�u�ü�Q���)���l��{R:�1a&�/j;��3�d��vk��$�ڳE�����},jIe��r�����Ol�fs��*V���T��G�	Y���)k/s��#�t�+5��҈f/�M��]�9��"Z�=�O&��5����%c]:�%�e �Ɇ�!�:�a�z<4���E�?�MC:�M>hV���FZ~��bʅ��-��u�%k�e�"�6j�ƈ��Ն�3��W�:U�يo��`ҔX|� �uX����	NsUgg�A�cA��(�=��K�ԙ6��R�k��*T�_}DJ����M�޲��d
\�U��Gr��!:B�;�Y ���y�r��]���{��q���RC���F�H�9��oX@�Z��'|�駟�?��O����ߢ�t�Us:	bՇ4<���0��M��ѭ�k:*C����/��	��}ܯ����q&LP/�����:�<z�˺/X\[�
�O����B=����Zh���d�m�� m��)���UЌu�����p��9M%+܆�ܮ�����Ų�xM�Z_<�&ܼ��l�@��^Ly.�X�=��ir��u��|;� ۜ�zl���`�۸�c�����<��?�K���v�!m�����Βa'А|���W��x���&<܂����.������{����F����Z������Ѩ7�uM���^��~�U���80��B�w]m�6C�����ٳ�R���Jg��Q�gMk(H�̌Z�ʫ�#�͢�+v����w��	�����L���:b/��V��*���:��m��0�䍲�m��A�ĺ�9��Ȣ�҈��3i�D��A��zyK�!:�%�򀽻t��X�)�=��E���_����d�RBT�9��Y��J�����vD�塚c�7��;�5�
�<�� xZgw:��b�W>5��X���u�,^kc�[�=Ũ�f��t�*W%N�/0�9�Y9�B T�$���;��=�u������e���5%�B�`,yE����ȸl4�����:���!�tۂH.�m�^;�����z�If�m�NMqs�:��\U��}�#���R��s|q���������4ྯ��o�Eԡw���w�F�W��h!�A�ޒ'5v�4*�E�u���=��7�s������֙L��Q�NY��8�����C���{��n��D�FZ2v���X���NllG]X4G]2�"�[ve�!QSz��#�80���ֿ��aЂ<�Q���A��W��Ғj�.Ϥ��~"r�{�V֗"��s��|T$���+<8�jt�����)���J���F����8�G�̓]�k�(��>ݢ�?o�(i�}��^��wa����0~�M�]�� �c���"���!����t�m��Y?�:�8\�����~P�����k�߯���b�u�wY�΂ ~8<�#��Τ|o��x�B3�5a
���k�~����%s�f���6M�Wërxq�(޴3\c��j����a� �ܨ�w�/�)ǚ�cp�F�i�U_u��o\�;�t���t^�'F�N��c�L�KkPK�s[2BuJY�����額A.�\��y,@���>�{7��RqJ�\v'G����}��fE�璋��e\��w;.�"�o��I�#l��I�G�1�$���x��O~P�.�M$b��:M��Β���&\ґ9��+#��Ė�%�Q,���%�@�dBZ��Hk��?d���+UJ���/������Q�gn��3��J��iR���/u,�"�x���+��뺃(��6��®S]qn���ۺ�X&�)=��o��-��X5.k�R��$U�A4�;�k^R��m����hG�$�m&���δ�K\WXd����6^�Q�t�#�;Q{l$KW�_����ډF7��c�����/Ű���-�����JZ�
ծ�X���jT�0�g�]M��{�U�>��3��2Z�>,q����C�
�.��d�L��������z�����t�Ր�A$�q�`5��@�<�T?���h5!��!����2�6���J{yA/l� 8͸��\���Vꗁ��Kꔍ��+�FaQ��.�Q�uO3����x
L��Ȗ�\k��U �Ŧ6)��Qo��q{_햺��ޅ��۵�E��G9��~]�R9E?8�����1VZ���@_�D�+�_V�S���T_�y
��@�P���\+�+|\>���0\�Hm@�T��*B�u(��z4���a�W��*����,@K�ߨ�Nv�Q̈�>��s������崻IgV���Q��������va�q��bJà��hi�|��wuV"�_S�
߇H:&�n�8F���(�QU�2�9��fu��a�%��'r��u�m��|.��8L�pc���%N��;�"b�^������!�ac��3�!���g����!u����9rV�3{#��yN��=$;�T.�	�������Ycs���i�;�4�M��vȸ@`���.5��xK�;	h��nS�|�ۅ���Q���%

�4�У?���Qh�5�!�hy���]��H��E1���R�7	O+��)$��<:�����ңN�t���!��`���"B�N�:mOA��0>.�#�ш�ψ������.���?S	݆O��g�}��@�1�:���"��)�!sc�3`\���?�?m�.�� �s�.)MŤ�2h4���ӭ27�V�Ҭs�ݶL��Zz��v%��sD�������
B0�X?�/�T��X;�/0eD����K!%�EL���g�!F:>���17�4	�X�4�m�FF�
�0ϐO;[K��g%����7;砗0~L�����@��3�\��Qo�ڣ>Z���F�������p8�u.ָ>}��X���լ��!��p}�ɾ��CR3tP\�1+9��މ��ة'&���I�k��F��9S�]��U�j z��T��E�9�֌���e4ZJ�6��!����S��r־� ]q)]S�Q�)�_��C`���hVM7��Kc�ܜ�ٺ0�o���~z�������X6���n���n�G%�l(�s�9����)o�jS�C�,�6
aH�������^����w��/�����c��1x�Q~wL�i2���hFx��an/�v0 ��ҿ��/Q�7��s6�7��נ�E���X����mV�,��J9��c�����E�1tn3DW5e���>x�72��H�h��t��i
��gwv���tO}�03=���)~���èk��<Bpb�p��,D���ʑ��Y?"ړWj8���.����E�tI��4��$�<��ru6��P��p����z�b��,b��o�uDCzK�8 ���D�0�_|�����V��gʐ��Y)�1�5l�#8ړ��(K͝��}���Zkt]+�Q3xm������F�������m��ɢ�	�K�T��M�s*�,�R�I�"+U��SϿ.�+��T��:�t
h垵iGe�ʒ��nw�����j�2���]6(�$��k�s�[�5��cG4�݃�t��nt��G��*�3��l��4
ÕS��V�5�s�l�Jc�}t����`��gI���R��5k��tJ���GN�|��]��Gt/�.�s\���8�b��3#�y��mW$�Nɏ�`]w����I�hs�~V�I�>�I��v٭�l��9���]��،(�\K�:���H{U���G߭�r��Q��F�*�I��R�ȹ���q���2�*���Q�t�k~�<F���%�D�;LB$׆v�OoѦlu�U��M�R?L��P��{\��`�����|/�����x�Á��̵�`������ZS�r�ܖ�N���5����K�����\ܡf65��ĪQ�*s�Ͷ�A����=U�{W�z���2�/�]D#v�H`��;t*���86����(�4"�4���ÐD|O���n�]j�L�5�����97?6��U3Ut��)kױ�Pp��ʵ��hI�x��	g���X%�.�N,�����Cj��0��������y��_��fI g�e�TD����e�M�$���9��>Ȉ:�+k��(��MU��Xx�͘[�(Q������?��d&���01��\����ET��k��񘥦��ӳ���h	�H���B;mН����ls��%��^�����k�[:&;W�!�;������b0ju��Xv�'�H��B�!�/�9�4Z�Y�C��]�c�&I\����>�!rV7*�<XTAJ[�E�(P�	L�A��z\<V��^�r��%�B���"�J����F������}$�z�/����x}�ٔ��<�'f�W��N,Θw<q~6�}l^c}�����.�� �jA�'}D�x��VcY|���
�n���ے�tA���0�N�p<���5h�R�xh�ȡ�Lה�s
R�~��0=X�Y�e��v5�_Oݞ�#"SA�1�3?�zJ��#�"�5hvT���T�
�VP|��˟���)�G����?]I���ގ�=9����7#��' ;ߦYƠTgx��(�{�9��
̈��z66�L�ɱ���!ź�J=)�Eݹ��T���,�hk
�;.ˠ숑:>�tj����3��h�����be�WN��H�5��U�9Z�I$�W�M��-D��s}��t5+@&@�F���p۱��}���퉨�ڶ�c����͕\ٵ�$��J����`Q��)��j�'�������y/Z�*#�NbG<W��q��	��l���:���}�e~bH�DX<u��d�[T�>܊Hk�i���̋i���Z���U���	-*��p�"u�y�i{[��'OAcPuӂN��k�J昆����;FFE.刦��07��T�,����{1o�otzϓYw��J<����J�T��˟7X-iAk*����B��,yE���O5��0~'�,J�FcĒW���L.��Q ��B|J��lpd�`)Rj��55�Y��yi*"6d�n(g!�q誂�e�~��(䬔�����rS��k���/��(4���x�~��>5��ˣ�vh)�H�J���Zi)�_��q�Rg;-�0N���A����Zm��1)���k%��q=K�� :O��Yb�oGqa���cmj����y?�7� x�h^��V���t���|&������~�I�v 1]�8�^�*/�]�o�J#M�c�w�������iIE(z��6Ga�S���J��b�(PSMk�|/�Ջ�d,������ǻ.M�3H��s��o}K�H�����~7Ym�ۅ�5m��Q��꠮{E^-�LX��I5t�O}Wv*�2���+�ۧ�C�F��1$�ȁ�pd&�tgʈ�c�1-��NQ����/C�������[�9h(J���/��R�ԩ-���ߡ ��H�_b2'����g����[���uI��}��t
���B�8�����R���v~�y*�c-�hBa3NbuT+�@�NLqCs�l�W�GN%^m��F�W�i�}j��u���i�G7WZ\��Qc��(j}�>>�(�ПP�F�R������U�@���T��p5&\�{.p��~��7G�<֡�x.W�$"�Y�:�1v[����^Ȅ�O-��\[c� �]��s��DDG��U����wh��I�3�Wu�2ݗ`<r1?��;{o3��)�{l�#���w_c=1�J���� ���Na���R��E���蜹v�=&Q�0�Uu��i�q�v8��N�ya�m�g��a��	���d���ت�o:�n���)�?��,�ZT�	w[%ѽԈ
\�"Bx�HQ�q9�8q��a�葑��=�ד�h|����e3WnC#ԝ���Wl�ܾ��K�{B���U��;ӈ_/��hBw���!��ڦ�}x�M�Z���?ǽ�����r�!��*m��yW��k-4F�*�t=#�ܫ]�g��F���/����o�OY`r���͚ɸg�pL0�6�������W�\�`H�V�8�5�M��c纇:���A���Ru�K�'�n�s�{~<O	�$�#����b�0�j<:ʖ[fgf~�8o�e�ƃ�:�ҨK����d�,��eۦۯwV�T����ڐV��ũiQ?��R]<B<fy��������!m�`��_���I����d���$C�����x���HQl�c�8�C�Ԉ��R�|ʈ�T"�.��o���,�h|00�Rv'eٽ{�E�p��4 bV�Ų��A��[��7�V�a%�=���>�C��$�"Z]aV���X>�;�,��97,���r��F|7�5���1��t(��r՛��/2���_�ߏ��ׯ?ۢQV�?�{��-�P���������:��[\꣨��/�3;{Ta�J_E0����Xv/��t�<2{�(V0Cv�dD*#6P� kz������#M^oM
��F�G���x���T�b�S��>!'!����ӑ���Fx�;v�5C�]Ȋ�k(����*ϔ�������%�r�(�6h��*�`g�����2�+��{����ω�{���E<�x]o��_a_��O�y�>��l���^؄�z��R5�35_��PZ	ZM9ǵ���X!�]j.��	|�.��.��P����_D�t�b4��Ԑ�A��!n�u)�Z�A��WsJ�
'2��E.���"��fQՑ�1��9ӳ�b�����y{]Ǌ�e�ےF�8Y{1S��@ ܑN��w]v�DBE!V�ORf*�K�϶��(���H���{n&8%��0ڦ�v��a@`</Ѳ9��"F������4-<}j��p�2��C���[u�C����a�=�x�j�:x�0h:���a���/�����Y���5H�PA5
D九CU�Z�Da	�Q���,)���\��Uųz��N��8vDs8�A?c�H>6v�3W29�i�U���f�L("��"��oa�~F�>�Q��ШRtܭ�S�rJ�!�J:��d���,�u��X�IYՐ�xy!C-�]*��X/�0�p���LH�65�֘�C��M�[2^�	�c��q�ޚ4�m��#��T�="B��O�̟�V�>qU�;��n�,45Xl�*�"]à�����v�Q�\����ESDI�i9M��u Į�j^����?$�}�F��	x9��\TI=t������h��-�<Cp��NB��9�d�ZS�X�w��1d��k�91Ǽ��W���d8��D`lB��x,?x3J:$�5Ƽ��.��t�������bRxg,��#�h�(
E�����QFJ*1�|�V<��9�6��˚�����I[���,)"��c�mH-���榉�}O�:#O��Y���3'<p���ypG�����E��D[lz�qF�iD�px8��3�<�a���9��\�EE��)�O.�\�q��UǱ1	s�1�H������OֆM�J��8����G�A3�I57��&��z4f6��T�6HW�A$��L8{�W��g_����Q��	�RL��~l���ר��JV�N8���ħl*������*,
T���T�rڽL�k��!E�-����!�U<I+��3U�c�=��⁛���"��iG��`�ys7�+pו�ô�Ò����@=�(�b���2�K����T����&Fz,��"b���{��Ҧ��XFW�|�ICz͡y����zS���k[Ȝtz ��D J�z��<RD�5�3�s�t^a�bX�VC���v]����#�<q�0��P�b�[��Ɛ5K�ف�g&��s��'eNYxd���\Ӗ�����������q��-������ÐZ��$��7"Rd;6�7�Z�kK�DT��=�/\�Y�r�юV�f�WE��]�Zz��e�<4$�?F4���4[��ɐ���+�x�~���\c���͠���Q�|\�s�-��pB�CR�'�r���4�Jb�}�tp�@CBQ�Ђ��q<ƽ��5���^��׼v�,m�<"�JSG��Cl8����Gۛ��q$IW �%�<=���?l�ݙn�$�@U�infQ$u�ՃEudFx�����{i��$���sׯ�@�.��COX�Ar��$���_��
��_e�]��ᒅ�n���Yz<4�7qQ���)+	9+�Y/K�TK������7���w7�\��fٞ����Ξ�Ln�1i���b��U��n7ǖu�"�)>#wA&;���-�,_I�6��ⶄU���*f�5A����D�L��=˙��$�����=Đ/�|����4T���ĜA;X�#~~��`�U��盤���c6{ч�TkrKOSU�7_�YpFಡ�?ݱ#�꺇�{fa,%#C���'TP������St���F�B݆ڟ��c�^����U�z�;`�y�*�>�;jOV)���<}!t_[I7��m�:S��r)ל�1Eύ;�ќ4�_���=E�G�O�nz��!���)�{j=�$M�=׫3��z���>��Z�~W�Q��� �ܾ�:7��hwz��^b�ۍ�7�����_�w�k_�t05�:�MF7PO�f��LE"�
�5Q�8V���e�����+��H�E���� [A��<����t�m������Ae?�h@U@�?S�98����N���7�|ZA��K�����cF��Z��p9�[�v���ߐ^�
�t"��zY�Jڧ�$�5�2��1��z��?���R�Q��R�.6̓#��^�
���]�+�/m���;���i�{�Ԗ�kv���k�i-����R�(��Z��,L5��"ؿD�j>/��sՑ�tU�>�A\r����:U(��Kzv٨ժDE�1���}���Z�7���I�K�Nl�jc��^����E9v�]~2ஂ�d_o���W�����ӧAw�(J�8�p��!�Xw'�N:�P��}�n�\Is�Ţ2{:�brp�CԦ�)�Mܳ�Z�c;n���$ǁ/� vƜ�p�I1�VtH���5�&w�	��7����kM�w�I�m�Ѓ���'Q�Vaa�Y������8�YN!��1nJ4�����!J��*�j��+SMR��3A�:�9pyy����K\h˩#��a�ün��G�V�]g�����rw��*��i-R-�n�7�=�X�*�I��i~�7	��Ԟ�#���$M��l����r�F&���.���G l��9��;y��0��2��2j�<�!��%D?���YS]�mv/�=1]�Q�F���h�!8B���鲳`W(�4�B�������S`��^6/d����ŚƵ�e�>O���M*��%�Z�pbhM^��+����sM'98|Y�ĺ�hs4��'��&�=LQ9��^������E�������*ؤ� �� �� �ɥ�z�����1�W��� �v�#f���@���ҐO���^Ģ��V'O+�V��t�m�=���,�tCg��m��!�'�]����h�}���o�Fr��}r��s�|\���L�n8͓�#dCX�������������o�dF����x�;ix`�I���ʎ�������ÿ��K\���F�����-�S��SE:�<{u��B�K�Y��u������I����f-��yR}6v�OќB)�(�uI6�f ?�L�jy�k@�O�!�k�n��-�t�*@{���
��l��a(^=�{h�(G��3#��G��C��3!Cw!�&q@=9-4d�G��$�`H�;���gZ�|f���b�[���f'v����"e*MJ�^//�)@mKd���'�d�]Ng�`f���P{8�rP�
�2�Yn���� ��|B�QS]�T{m'DD�����堄�d��Z��.K�k��	d��fCC������������a�����7��;��%�
�t@E�set� Ȫ��s��|b��'Ɗ�$��������2u��'
�7�)gk�l?&��,r߾��J��&���2��Ϳ�����+����[���-cq	vp�Ml<i��>�R�"�u���wఠ��������3�ƠjQɃ��2��֘ePbp�bb�������g�Pcv}\�f\��F�W݅v�N3PK��S9�j����@Yj��X�Y��7KG�&s� ����#�"me��`bv�57�-�Ɲ�#���yF/�ezA��B��ћ�d78���V9҃^�Ճ�r4���rZ�3C9iZ-Wc��16*J?�ǍƤ�*8õ���(��N�"(���:=��I8 ���/���N.����@�sS�[�o�'b��Ab,�x�ֿ�&#��2�}�z�������C.�6��O|~�����I��#�V�t�}{NћC�z�������Z���0�):��Ԥ���]��\��舲�!�����p�Pu5)����XݽrV�}�:�h�*fCZA�4m.M$[��.�j�xʟ��3Jv_`��κ��<����[��.�BC<&Q��=���:�!�;Jz�zn�0���6:�o��y�vdM�xP&�I�\B�$��؄Ѕl8h����ufP9$��R�9�i��;i�����C|G�(3Y�m-�6��GM� ���L4Up��uks��YF�"�����$J#�~�̏�)�Y(� �\¿I5�)6�Sl�
C�Y@\�p�<������Qaʟ᪬sTv�����A)��Z��)���,8������h�5���BU��7>�ǒX3�*h1�P�8m�u�jz�v�fp�(	F�����O��},���5��{~��h���D'S���uh�P�S��r5�g�E#�d ��{�w�_��!SĎ
��"��	�������
�]��k�X�ȫxn)u:��N����i+JN����sw 'm��Ϧ��]��k��N\\)׆�iV���7+Q�ǣ�ߐ����W��:��Az�vus�k��"�?<�wCI�쩠�r�F�R1G=SL@�;�I��\HY>���-�6�GTL��ׅ	j��\h�D&��T��猍���X/>w%�.�$�H8�ZE�y��K�@�����{��8�{�Μ�>�x�d�^��~�46&Kύf譵YR%����?�Z�&�#���c���E����C�øn޿o��G� ����0I��$([%�8���P�����p>~��(�0����%�7?EC�Sy��w"������_����*�5����~����im�J ߼?>��qGU$���<�Lz�C<�C�0W%#0�	Av�	�Q�9�m{�r��;x_����ϟc�j�	A�f���G9�:I|�����X�
$R�j�1�n���>�}�uP�8т�ҟ>=��xo8�pXұ��`Ҡ�5�0^/�Go���F�^瘘�0a�=�}��碵�S�0��[l4��ju>Mk���l;#�$�MY��ɫ�^�x�ke����w)/��
�8^eñ�z�H:�c�W������Q�i/*M:��@ܳ(-k���I�\b2���K�[��qҌ�׈���Kx�<�^U�����Wf�F�DE��k-���v�1�`M�'c����5؊�u�ȼ �ahW�K�3E͓P����\��#�k=�ѯ��Җ�N99Уt�Jt�\].N�a/��1샑M!���	����Qvɸ.�PT] @�u��X#�{�z*�Ѐ���h����Fc�Âd�x��P�w]8�rg�?b�J�O�M�u���:�����?
Yt����90�y���}P��}��9�i"�5�W�
rm1 �,��@��w����M"�>Ή�r"���������Qd��y��O������9އ\"�o���I��?�(2a������KH?š��A���f�M�����}ܶ1���A��䃄Vnӵ���W��*�i���0���
H�T�����G�`W��+K��k-�/'*�ʦ�#ַ,�R��6f��|������m̮��4x��ã���@�A��b���o�5�}��B����EA���ZCЃ��,���7�v���"B6��g��V��ܗ�0�lQ:z��"�<�΁x�S��t".�.8���� ��6r�,�l�]��s�QS"H�r�� 1�¹�{~�A�v{��e�nI��\@�����MA�Q�]#��ks YB)Q^�xsd�����9>J���q��(��u���T.�1��^�����R����#�b����M��Ƿ���G'��Z(���&���G�VO�J�2h8����>���,?��kc@���[�W�e�	Ki7/���P^V���>V<��L�C�e�0����X~��;�ϟ^i�c����8��m���Ĳs��Ʊ��:����.�~�6�H�>{v�cp"���<$������q\���qd�x\d�q�1�z.ဨ�x���ஜ/MϢ�_G��&Lr�dlg)v����z����3�k���҆��)q�_�?�l���DT���7�+u��&5��.
��6*g�ݾ�#�f����<�Ήz��d�5�i%w�����N��Pl�Aafr����t��M�$(^G��}��F9-��R��jx͛�uIk)
���6i{��)+
�"p�s(���s"��i4�LD�z�Öt"���¨�T��ކ|�U�O1�ݕ8<^� q[.�T�G ��U��׽U��Ɔ��4�X����N�)�2Q�������t���,�oH_?F0����3�&���h3|�h������E�1�V�����Lm���A�]���^"�}]��E �H�P"C �k�Z>��%��g��X�� ��� ZĽ��w�����a����JTS�I�Gq/������1_��ܷ�AΚj�3i�3�8�=JR;��J8M�b�E�Z�k0O��8��tן��9�n�u61�zyu�\��s+��f�����q8a�]�& ��/���@�ʱ�7�dwL�hY;���9W u�� s�I�^��gB*�@ϻ�~e��6YR��J��[42��;N���m8����Y�^4	7�\���frt��D]e�]d]���;/2��"�F1%t�EH�Љ�M��s��{��뚳���`(�_�I�A�ڳK@����|�G�6�ͳ�ЀO���͗�ٳ��N+��*>��W���5����c�|w|�3�!��CK����-$�@�ڢL��A�!X��#3zz<EF4��g���4�YjH�P�6�f�(9�m�p0$pH]`>}
�A����gpoH�zzzZ���Ncઠ�m�ff��4�T��'�7����/�	�ϟ�˻�~����4�2���5������xo;`�ȑ�a��������~(03BFZ�C�����=�@LӞ�ȅ/ܛ�;�Jg]oǚ����t���XC�g���M/Yu(s�D��FjV��X�rTz���l��N�])��X� ��}ߘ�ڀT�'.u_b�����Y�E�1�!�g���Ω����zY���4�N��N�ά׍w��j!fKm�֌��%v������5�Ly����{!2@a�������<����F�]�8���C���qȔH2*���D�.#���.��i���ZF�.�
ϰb�F�L��=�i���D�P���'u�%���E��ڙ3�cgg.bdQ��cr�(,��-���+�	�^��W�ϛT��Ӎ�#�\\�l��fA�9{�Y-�����A�E�?�|Ytd�ȓ� �m��lݪ�!�R��'e��I�O�t�y����Yu�	���&XP{?2Øk7���z�oR'�2c�'���*����h�@D΢vE`����/X�`8s�Pƶ]���s=�������sw�<��9b����[��቗P*�4Fv�l���1֋3y�q�I�
�1&����Ou��� Iȝ�߱6@g{~f�fyʃ���M�̓�b����AL��Ǟ��^z��E�-���vS���+v 㾭�ڴٴ.k�4u�`k��d��Kh7��EV���qm�(�lu�� �L���|��!�N�V�Q�� ��[�@b(�֨֊����7����dvϠe�p�<�;�&�O3������N: N}ʾ�l �K	�r��N8 M�2�cw�����SC�h�$�CM���S��u�v��[���6������{��[�6���f*11�o]�[���
��ѭ�MG��YJ���Q�l�����q�:`��B��48�륈�9�%�?��Oy�c<1�"eL9�t<��f�82�z�`�yB���)�Z�g��Ee����^�
	!-L�I��l����ŭ�E��D�9�f�]�)����׌���L	x9\X�w�38:f���ؤ��I�}/%OYŁrҰAY��O�
��a '
�#x��VѴ��D��!5�?�R�nFl���f��(�W�V]�m3���M!��F��Y}����y�������Z�>�߇��'/ٱ$�TдH�J&9�V�|���G�{���?�[����ԋvc�h[�Y�	ߜ�s΋�bw��47(�����B�˼
nZ��!#m�Ѹ�lt;�c�.Q��L �:�(qv�C�9,��:��Z�0���,��!PY�|���>��q�'g��5�K^h/�b&�e�p�#hE��j £�\�ө��i�.阞Y�2R`y��u�(wH�-
�2R�U-�=~��1I:�T�I4�S<�cp\��x!���ۏ�!�@���~����u\W��m�m�ue���@J��W��{�P1ե	�5���ag���Y�f����˨ό���C���,�d�葝O·�~{e�$�[�7o�i����\]��P���އ%�����mHL;�A�+!���z�`�)��ک罸�@sוR���kC�o�F#;bʟw��U��E�Ӏ5@�^�p}N�Ep(���$V��vB��cÖ�C�����?��A�>��Q�GG���s�w�E�RS�=Pݧ(p~��U�Ө~%-*�g	~t2��������HsZ�� ���)�2+,�1�G���EK�?'U�����]JB&ʏ'l©�"��z��/�v#+�N�(^�R��S;��5H�A.��x����&jZ[r5�f��,Ѕ.��+I��,b� �Mg����B�Sf�=�j�<@Mu�F��4��C
���M4��ؕ�F�3��妃U��ڠ.�m���XJ����pd�H��e�u��H4������5�;XV>3�Q��E�A����kN�W+p�Lԝjg�س��}5c�k�m톅�����@�e�Y�$�֫��^���#56��N�%R��o�@�����;��ٱ���-�b����<j?@����y튣-p�|؅�^�5�SOy"�k���~�K���Z1��l6�@���b\�ӆʠ���7(�gG���g#�i��oc��u�"Et�y $�T6���YV6�"��}��i�D`e�{ٚM*Ŧ��d{S*E�� ն�iVԬbu`��C2e�)�/�S<;��^�Ag�r]���P����@�g ��"��ɩ���Q<�v��)+�D�-��PI�C'�G	��Y{��G���:�2��|zJ򼗨qPܓ���u -f`qz���fxC��K]�J��U���d���ꉁ���Gُ��<���%�r������򗫺��T���$y�t��j��dO�)��vZ���!qH��Uƹ�W�e�IRZ�0��<�	�a�����W�w@Q�۞�d�h��Zn������(�V>q`k�ٍg��9�}���At�x����*���/��Y4������u����Z
��x�rs�Y���͘J:}�VGPA�~�<1��βXG���yNT�@����+��=y�\7�n�
:[��Ak�3��Rf�x(p�eS����Le�S��4t�%q�:�ϸ4�閥�3� ����)�*ŵ��̦��3S���Ag�L�&�����sy>�'8��z�E�b�e��H/1�s8&��2�&g�P��|�@�=?Jo��1��A��x/�J��ׯ�����D�}��9p��Z���)s6�\Γ�>�ߡ�8��r��2����`�x����p=qDl�ęnM&��D�EA���_����ս�oyy�,����Pl�TI�#�)�u�v<��QA<̗gk�.�[���&��L��6�$~�A-�N�E}�T���*�܅M����IX�*F�C��-� ��b��� ���Ӎ��Kǆs&'}�rG�|?��O1���-(��L�?����0���:Q2����tk����w:�}/ޤR(T�vnD�xx�}�H��ٳܳz_{��vF:@����c�M��]���(�}8@:����ܺYT���M��K��"��Yw�/w�tSFjm�^��m��@fO�������x�d!����M0�)2��כ&ep�%/����c��ڙ�Rc�1Y����2�~�����E��w��V�"40�?����X/(��;�ie�a���n|t]fQ�?��~��j������g��T�JT1v�{��拌��Z^8ʫ,ބ�<Ħ1��K����E ��XN�H��Ǣ&!}w�����)����?�/:D.z���� ���ݓub�q��JQw���:X�ڥ�gJ�i��j��JJ1{&�:�O���A��R{��Ą@��k�5�?���m�-��F��"��z�MNc��_Gį��� ��Գ�1gt֔��iW;�E4�Q�ZX�I�-��&뛆�S ڠ(� ��) �E��>7���k�qRZKf���dBD��v�TWf �tƯ���?���1OS�Lv$i|>Kpa������:�gv�դ�@��_��)��U�#����#F�48�\�]��?��l~��H"�^)׆�2���U��1ˍ�zzb@l癱�0�
n���~F����X!��w>H�ً={���{#��b��.&+��h>a�}�v)�SWXx,�.B�A���+���w�0H& 6�����:��P¿}���{+�����uVy���[����8i�b?ZfQA.��:�/�=�/��N9�΁���l:d-�iv����kH|�b�����=�P�g���c���@8�4�[c��]/�t�T��{�԰�ޜod	���"��Tc��=a�[�w�L��ke���� `�58��E�G�����{��ߍ��;$���{7�콦ٝ>�f���&�7�l<�	��}���Cn���\�q�^��o�(`��]���F@�SY� �˸�����b�:0����x�v-��73
�9�<ˣ��%>��A�`AK{e˶���l��%�X�F#p]լ��9�1�[��Y��*�8�j|�Q�hp ��cZX�1,>h�A�f(uC���%Ki�.�+�������� M ��qm0s��?�ԟI4;�^���_�J���b�G�X��9�����}C���������=�c��|&���q�,����I~���di�2kF>iGRײ�B45	~_�`�`��cTdNڢ�dt��f�³|��D�(��/̽n�K�\]
����M�[7Gs���t�t��Vj�/u:r�(��Ȱ���H�{��4�>�f���b��V���%����X�+Q-��I8i�i
��B�����%����X��K�m�>�d3��)�S֪m	6LMׯ�2#�� �U��e��JXx��G��x���
)�|J�Z,wO�M�9��M��6f�4U&��i�A�<vC�Wף��YQ�����Bdիl�䅮�;Q�wkx�[�x�tVĶ�4(��iu�  !��o�������'�4��tV�Gf1X���p�7<��+�;����1��?���as���߄;���V������Z�1=q>~Y��jV���	��93(�}�>Є�
V�8$ı��� (�i�w��k���ӎ�{��)���y��90@`[�ەk��������fN�5)����*�#^/��cr�)����SB6uϲ�������p��"�[��UMKq2��0�4�Q�H�Cp����T�2�#<ΐ�T��CvQ��MUK7��y�X���d�o����/]���>�BAu�%��%�48���ڹ�KzH�/��[�����;��=�[S��}(� e�4��O�ւ	�����5��:�U�)i5�TU�M�pY�7���t�[<����H��S;�M�����}�p�j]���'v1Mb�S���i7�Ry�6��P9�p��"�{��l�
����Q�`�*}~~as�~[�w�8�!nR��s�ĩb�\�ul6H{��_�o�mN�0!:;��q����.D�q���Ø~`���ld��\e4dN��ŦH@C����3�|�D�0�>���Mc�^31n(̝�2���U��V��1(�|z�u"����o7lOE�|oN*M�Zi�b8fO�t�,3�:�V�#yP� ���b�w{���oѕjC�ƌ/g�I�� ^�2�4=�4��	��mKHq���
������^̓�w�y�i��T�Z�����S������_��^�m�:��u��	�ߒ�]37(ğ3�jbx0:�~=!���)J�SLEt9�L�^�i7���o���B���<�a�{�h$��Jadv������ )�>Ȑm9ι���5�N,-��Pv{͸	��	�W�=b荻����x�uEP��`�������X��Մ�?<=
Ҙ3�<�#�,n/����8=��o� �v�q���9�u���hx �GV��v6���J@J6K��-%�kB��9P����i��;��A�J& z_+�u�"�?�߹�<^k���y&�T�7�d�+�v��T�Ǝ��k{��!x3��^�Ǯ8�����s�M~��b
�>�0�K^<�Aέ�g�=o)GB��Ps�|S%E�ʸ��3f��M�/ga�� �aί�F
��8��ޜ�G�i��?�9�{.�X�t�����F�"�ޕ���&�6�Ѷ�7��[�֓����ds�䲰9T2���^¢d�M�2d�����o�����>	�\7I�ֳ�u
9��\Oݦ�o7)3
`'��}vm�Ɨ��V�H�ͅ����nI��x��3�c���k��4'�z6�u ݄)35���ծ�%u)Wa�fT���!���~�v~<�n�U���9����\�߾��Wo*��ש�IXup��L�)����qN�<C9��8W��X��w���9�g�������pQ��nuܷ�@�D���R�z)[M�E8��)�~� ��[��?����� �
�l�1�@�j�M�A��]���̫�#p�~xT�q���mP���U��QJSn�ڕ�^W���;�y�G@��$�}��л�^m��t#�!� [N\��-��)0r%���=ǟO		���R��u�i�U��P#���9��������x|�#m�h�rs�48gt
u��PX�C^,�ͳ��������a'�L$�Q�|�]��L`le���-q�%����d��'d��j��V�F�Ӱ��qk��'H���JQOzK��e��ϧ30wC���A��D�����Y� �i'�5M�����.��\�_��$�6����D;��d��!K�E�����gI�]�^��I��a�������l�8h���x�Ȫ������-y'�k~/�24����X\^��?���O+��>_kC�nV
c6��u�O�q����A�F��J����Y����.G�V�=u�4��|1�
���fp���)���G�u����2{��㯒�NL���ł9��cO�*5ĵ�|��ʰ9�B�o���pH"�l�cvO*��¸���'���Wٞ#p�6�Ȟp��\W��)!�1���C��ڑ��EAT��lp�&�C��v��o�2��mjN͍:Ԡ� /�3G���T�����������a�SK^P���I�.`�
��B��\T2+����LRC�`0�Z�=\�����9N��T��Y��jC<����H�H�ͻ�!�j�l������B�r��tv�;��Ҷe�V��G���T�L���z̊��ޑ	�>P�>�	�\5F��N�̳�~ȞVM\��_/��[���X)��*�7�+�ݕ�˪XνuD������|�߻zp������M��_��څ�W:���Z�`��h0AC �5�����J��vCf���T����8��hm�|_���T�e<���`@FMqh��w�K[��-/%�E:!�RR���:½�=O���?V?C����^[Bk�<��^��1���k���.z9{&�/����u��'��E�ON5AR����C���)O��M�ʕv�1*&"�)x�)�S���IrA��6v���<e��`C��Ħ��ER����s��GM&���"�������fT��R�GׁԓV>4��٢2�U���j@���q���	Xg �U�zu>q��^)U�^�qx�\)��������M�Xg�x���J �Q��]����%V�+Ǜ?��1/	����5�Q(�G6H��i�̌��Db<O�{�Hm��뷪���vS٧��v�@35x�}�V*�t��(?W'���qi�5/T�����+-aH)���a�M6	�{�F���s�NU�o�4`0�kɷ���m�lD2�0މ0�8�,�=k#hE�{ӠΞ��6�����HF��މ�'�t7���pz�d���Ғ��j�1�I
�����v�#����	�������\3Ҍ�y�kǯ�f�f�ܰU����c���B�l�A&N���~�D�CNk�B�`G<jZ
4�.�A=)���h�\q/�Q����(AcE*�]��tgW�c@^�sm0���Jڔ�I�y����G��
��u���USP%��a� �i���J �Ҧԍ�l�p�\M5�7������T�������>׀	�Z��:�)����� o:��>�lF��u��GPb}�"�x�')�b�uW�~�����%a�P��B>D���b7-���.�<�^BԼ���3����%�T��##�J�*���3�|fL�a���A��:.�g������h@���9+����eAZx.POJ`pHU�j���k����M\��㘦�̲.BI>d���}:S����O����d �0A�a]-C��Z��F�����F���O��/m����i�u�a�W��,�\D^H��Dƹ�m�;)�HE�I��i'��<i֜���TP O�Jpv��cg��ݙ�����rn�����kL	3�7v���<�BMĀd���(%he;(&&Z����ߋ�����"�����`s�.2�ۜ�Vˇ~�e���������'MѾ��K��	_��q�T��p�2��iL�P>�RL2��:�����r9�st&�����bdM�����9d�.):����Y����`�!���'w��9��<_4���q՛h�I3��).O�h[��g~��w�	��-e���{���וz��!��k�M8p�^/}�mVڮC߫d�d�(�>zQ׼�|�C��:�ͭ\�Y��<�����uO���S)�7�ЍF�gK��xc�{����s�<����&�&�%l�+� �'wi�O���[�?����W�)�ea�|��9qb#<pAѨ	L6�.��d�[���QB�_,��K�F������Tm�>���X��V*G��m#&��}�_�s�{sF�Ƿ����g���~w�z�&��ޤ9��W�97�)-��O���e2;09�.`�9H�����<j2{4TRJ'�@��^���� ���������wm(��P��@����]2{�}��l;��ْ�p���~�(��!��Nn���� �S��/�l�L8I;7�Y�I�4��O���kD�+zз{6�½ ���5��t��Ra��HKi	'�Ze|�N��Jm��C^j��{�f rd�щ�-Я�q��ٙ~f�Seܰ�h ��!Ý���C��U��A��0/��P�B�:#��=�ŝ�z4������� w���$7�J�u	�@�0��k��Km_�9	��
���;,�n�56����;t���GS#��$죄�x�;� ��5�ۮ�&�ŧ���7k)*@(C��	�HM���ZD��*�X=AUr\�!�go�H�!��W�D���Ec�k9�?��S�6>��s� ���M�|�x(W�KJ���|jp�oU��S�=΋h`�1��������9��+��zaS.������������n�L� �0������*d�󭔦�C+�*=�����M���l4ua�\9�X,g����0ډ�����h>-�~������$�]���<W�H�6���Ī�J�wgہ!����C&�GM�AWT�����\���j�#�}���ة+������:��Ӽ'Q8p_o����[�s�w��N�rruR����|.�8���_�Q���j��o���=/蠓��h�����h�#��{���[�$u��NYbn�#(ޮ�$����0�S.<�#uOM{�t�k�1���2@�d�Ň���X��2S)%
��]����&+5�a��6��,�IB�{e���eOy�q�uH�j�� �q���(����K]\�Y'���yT*�CG����NM�.��7Mm�eQE�םe����A�5��;��>]��=u�k������6����<[e*ᭁ���M��d ��ds�\�q��J\;��Yk5醟le��A&8b� �ö�$�:����+�*a�h���o���2ŗ���~{#�'��Z��v/�N����E-Av���������W�^R[�������u�� RZ{ߔ|�;�z��8�9xQ����	�y��J00�5|�)<�H�rCsJV���V�r���sXPO䚢J=MY�x&�����+����o��m���1���8fM��u�9ȘTo�cU��p�t�~Z��R9�Wv�ŗ+���>|��y`^$4dG1.��r�Ml8�Ү��:���%q*y�|�������o3�Mݓ�6�pc���%�3��ږ:yG�{��lD50�8�Ao��M�좻�`�pZ�Yf���,��9:�ƣZ/(3�Tz�R�8�2��6��Z�|?��f���4���{��{M��� {�	'�L�0��.�T�-vMk��*N������b`َ��nnW� �C�e2�C�����[
߻z�&ݯ(�����4�v17PE�y�Qz� ���p�T�y���= �	�Q��#��w\��"̤F����~gC	2��N-�^���d�v`�Ӄԟ��z�u�V(~����x�������@ho&���Õb���*��6�(�&��c�݅,��aO�7��_<�	���͵�n��vRP�xv7�F�$&H��q��b?�;�dsȪQ�q�/��T	<�عIrNߛk��u�C��W��I��6%��G32c��5�ˇC�qA�G^�恾�A�)&N�v��M��D�B��o��+�,j2!xDV"�l^�,�	�����c����%=��r��NW��uW��fGW7�DʍԛmK�z̸oc�w\o7��ۏjȬ���P`r����:�d�^���� �၁����-;�7�w��Ip23�WZJ�Z�d �@�Z	�83�mIu0h�td�6�ǀ���X�-�l�L\g��@�I��n�����*�b��`��Kj;`;�s��V���nj?|H)-�'��
fPߛcB�R!���	Wv�\�ig� {��d�b���ס��ņ�5�e��&i��]��X̹�FK�G���.�X�.�Ya���MU��*�x���4J��'��Rl�FG���q�8�2�v#�&�� �
��#��{��%D� �̋v s#��1St�Gv��� �-N��t'.Z���{���Z���Y�0�3��v�V�K�%�$�ȗ�E�&���)K�Ȟ��R��.�IN�&�GF�X6 -���*x�q�#��4���9�\���8=u��C�b�YsN��e��n��Z�|�>"[���H*�ҁ��`�����rd!o��fɛ��]��ΰn�9�,Jͬ��kP;�΂�~�m`��56�q���(��U"�eD�ٲf�lZ���!�
��f��������8�v�@��6�U�bL�F�p*��؍�2�i�0�������z`�7%I[⪮ڒ(��]���6m��)���ăx�q}fNW�gӚI�s�bV���[4��� &��|<Q��ja4�+j�Ep]��.�;��zC'�	��/�Ocs�w-�\���tk�v(\$_ܢ��l��[���ݞ%U���lB��Д"{��p(�C��6g�'����R�Kل3�$�ki����ԩ��*(ߺ�J
r���>��˞��`��|�:r��j�˵�N񾆻��ϒ]y�}�yv���0)݃\eP���(*�W�t�4^LӞ���6wWL���ߔE����ݑ=_�{�s���@pg��2��*XUC6���2��1[7�JWED2�뛀m������RU�9��2������D����yL���S��0��nB�$�"vVw|}a�ى���8�aF�q������c^O��H`X�w{)v��{��U�j٫ÃY8��|��;7T[m�]a��׺l��^��`���,���FU���w7��d���M�j[�D�C/w��jjc~&���H·���4eU�K =l�a
�9K�*uv�TS\H]d�}��$�%��A�������PX����|�G���ARFi�믿1��ܕ-
_��G6�B�/��;<�z��&�n�W͋ǍBgz���5G�˅x�Ό�I��f���l��, �K]�D�4��%k�Iޮp:c�}Gs86\?���Y.��>9�g�� Q������A��T�Oy}Z �AqU� �˛�2,�+�6���|Px��z���a�=zH��oӁo;q7�z���nE&>�=��!��6}����	@�;���{k�"4��H���;o\7�Z�c�ӉV y�"�T)��PN��'G��xJi��y�0êe*�{嶎�4wݻ��d 1u�ϓL����fx$�Ьqg����y�:�2�0�xx߳I�tb�1��N�0q��M�U=�{o�-�������Ҿ���l����.d~5?��=%����ӧ���|�M����`GfLM��xS/<f�N����,c5 m��w/�>O�|�P)'	-�RÓ�A?S��=�?���T=y[�^�6�H:K��������@��C�O���g��ncf��"ٓ_�剬wM�u�Y�.)�@����p��=�F01<����"��g�w����m"�&F�<�T�yV�����q�`�����)=��F��e�����4eҍV�=�
O��'��Toj0yw��P3Dp�R�̒���ؠ��8V�	|ѹc�|:�0��XDzqݬM ��Y4}��;�қ�������A3�W�����Ca.�߿�5��#����`������k�9��cI�*$t�j��-k��*�M~��u0ދ'(1����Tŵ������>�_R��+�3A_4�8F5Z��[]��Q�r�8^��:%%�_:�c7��s�̀pK�i^A�9O�S�N0�:n��A���`���8�w�^��w����4�04�y��z��;�7��������C,��, R;��O<�����8~I�7��=�0H`��C�R���i$FH,�Y2n$�AэS�~Cvf��Ւ��&|qxu�DWk�v�H��u�B�X�D�����"��t����R�}��XX"�>Dx�yܪ�gسt�(Rk೓  TևtC,Y ��Kb���	��=O�9���С������x��fu���s�w������ij�7��CND�Z�sl��_#�Q��ȕ�͆.�6���J_E�q��p��V�e?�p�����������@��d9�i8�d���������v��GB!_���y�^�F'�����.�J��t�-�&��H�z0��n��%c����u6NH�D��f|xIz�=w�2�\�8;NFJ���O�A�y�#�Fs��&`�l��e�טj�ƻ��\ڗ?y0]_Se��P<.���2fi~.;��/������eJ�E���4>q��y�Lm��ׄn�P�ڻ2x�T���F�9�k��e3L��6��Y�V�n�k)�4��|�hSX�a`v��'��fv��^�ZQ�P�r� /VKj9j�@��
xa�Cc�~}b_��B�5lC�{�}�M'��l�q'ecK��<�4D`}L��I�Ђ<!�8�%{`�lѳҊu�,p9��G/��m�����T[�2T:�6���݆(���A�BҼS4�	��G%1��ާ�ot���K%,w�IO:]3��ĩ,'��~�k��)� ��Y�[[ ��dG�����1��]@�G6���+��Bc�r�sLY�t0v,��!��l�Ԣl��{ ��6�.�ec�VD��z�O�"�6���e�Q�v����u]��8m���FE��Ѯ���b���7��%6��?���f�VO�U�`ΐ��&K���U�{�������^<�͋���ub�Z�����*��ZvoV��tYFw�אS���"�����j.i��;R|_�y����f�H�3����{ʛ~ϗ@��5}���At5��{P܍\�(���m��jɟ��U�j�?�纃<~d0���40߶����#a�x�%'�ꤔ�i<�ͩ�MSa�kLY��@ځ�׮EY�z��Z�Bb�]�0�,���b�\�(m�w�D.��T���r-V��m�0����MP�%��dbn�Y5Fi=�U<��_:�4
9)��N���lP!�tox :��F\���ǭfל�@�(9���J�{�Pk"klpXw�݄�>AHW9��ő&P�mW'^�Y���2��E ��އ�g�A�a����~��'��u�b��n����������d�5 ͳ�V�u9Ŗ
M��`Piq�i�m����� ��cy���n�yѐExa{�Ėƞ�"=��o2���>��~���{�<y#P�A]�oL�c��6ܼ�,,��r�l����D�:sDF5*&H�&/4b����
�����QS[W�{y<�������.�������
�.�P��½AF
#86�^�Y�����"q���tw��^����ڢ޴�r�@s�՜�:�[�=�J���,)��v[�����Sq�~�m�^Wm�q�!Hڌ�У&��>�<�G���X�t4W��Op����
{��)�y���JR�~ۛ)_48�.��r�\����>r����~���F�����.�����[I��y�lJ�5�~n�ƺ�>�ҽdF�,=���S�Y�k�O�Ij�5\	���_��RS�/Z@_��6x~'�$�z�q�]j)hG�P qf��eZ1׈�]�v�7��g��z��91�d`�����Y_���ḩ?i4nf��n
`�tJBv1���x]u7���%�	۫�Z��%R�.���Ϝ�gad�},���`�Nb�z(cߧ�%��$M,����#�nKR���wZ�������sٴ$Y9	�%��t�c[�um6����o�=�M��n�����`b��J�o�g��Y��7Q�[ı.f���Fl7�5�`C������x�u�]Z�!��}���n��Pu�xK�=�W�L	٘+�^��>��z���F���׍�%��ɍ�v�t.'9�..��z}.KQ�ݒ��,���0�8��O���mm��u,���u4�m��]Y)t(>?��=��YY6���{���{ߙe��Nr�+��a��N��o��c����a ����B7Л�a���jRJh�0*��6z!�s�����@�]�Ɍs`Q}7�w�.(�r�PO�o.�7�Ln�鲲1��5��1[�AR۷�5��Y�����I��FJP{�o��d4����8n%��i*��i8�M��d�x�}���g[,�a�E?ц��?~:�
7vUU�"W�k�ƺع�`��K�A��#ػ,��m�V�#���U���x�X�֔k����K4^;�6�ei��0�Lq��4Ռ�np��������`�����鋽ݭK��?�2�n��*����FS���MN�t��J)Y�sj?)�;8����.A���:�l�((b?0��E�7e��.�{Ů�+�)�#K��^Z3�:�o��&D��Z� �����1�wf��9��� ]c����M��E1��j�o��~�0R��?��΢"$�ZxdV�vG���	��T,8q���� � �R֪1�2_�ų�8j89�js�>ﹸ��\�c)�ŁB�%�2܀h�j3L��$Rl蝍"p�(#H�۶	*`w<4Ew_���ٝ��pm�[�y�r�-5Ե����I�A��"��IM$���.��m_�13�a����=�W�>΢�E����Ȥbn���x�l��a����X�#(tZ�&��⮮ ��"o5���Y�~�ᴵ�otf�\7�V��{��XC��8X���q�c�|������'x�F��9��4	��m����^�9��"�yO\%�r�ޘ����%f�5�"���>�1[�1�$���^P�֜x�qτ�Tq��:������&�ld$`d���SR4�^!�8�J��5�������,-��y�-��Ɖ���\�C��F~�LQ��C6�����T�8����X�We���OK{\dd����b5�[n;"���Ơ,���Sg��V�{�w<�D�Fwt�t�ŵ q�.�
r�H�{��j��&;w�������1���Y�\Yf��=���x�Z��;��߽1���`�L��q����In��q����j����������84(f���������u(�@Τ�E)�f�kT1P��^HG����|��m�}�tࠡ�*އM�B�ے�5,3epۅ���|�Vy�=Ƥ�A<:/�����)�qOZ͞�g���4�!=ծϟ�0C�9> pX�� ��]���/Z���e��w�T�g u�#���ΌY׾C]ۤ��׏C[���{f�Ūe%L3p<����ة)d�a��U�� ��~�jZf�T�_'D[�E�),��)��@s#.+�I��"�:��)�Jʖ����Oү�z��O�O�#j�a��=�`B�i�T��C��8���]�l��r2�������EP�MxF7�]3��2���P�b�p� �o�W��z��]E���Ke̙3�����P��4�����I�(�Q��n��a�ު�5���0�7⠊�e�G	u>O��G$�^��Y
�*�6�Yn���iw�k�E6K��cP��Vv�C	�0���¶��\;f��Ԡ��+�_���C#�1fS)Mkڸ��ۘ�ff���b��HT�l����ˋ3
��UwЍ&�nN4k$ޫ��)\L��JΔ����t��-�X����_�_��L�*�FC�+:)w������Ө�m������$� �hk�u�&h0_�N;1�ܟ�S�&���8s����Q��l�*�£e8 c���/��䜽G��������*�@�������N��?���ฌ��5�jb�:K�6�B$d�)�y[�Ӛl�`� ��.5�*3���z���|*{�\�1%P �Kj����Y4y�@�b~5�۲��zU���|��S��z1U�x�l�;���Y��3~�kT�����?�L�]J4�8�0��c��S6���}�ƴ�K!M�\Śp�$&��+8�q<��)��XR,�ɂ�x<�#�����Z�KS�VL��wU~��b�球��'��vg��(TR������U����{U3�ǒ<� �ע� �j�źC���-�q/O���J�K�Q��%	��x���҇���L]�w�TMD^C���Cl"���zkϞ�_-�m��EW�\���SO1�9�{�S5���)1H�/��s���H;�/�hT��Q-��4H�xWf�8��;C��<��uM�r���*��{�k�5ww��}X�"���_7����bF
�����L�A�B~��L�4ѣ>�HԹ�%6=���g,� =���&��a���EQm,U��������������o�9y��7�*��H����!`GU۱tw��04p�l�1��XG5C�X������4{d��3S���W&�#�"軙�\��I�A��:c*�����:��~�H!����{ٞ���$,9�>��><$��
�
mYӟ$�+�3ҾvT=�y�6�i`��w��g���Z����Q���u���r:8��%:�vj��j���0�:�~#��a|�0�?�89��
�{f9l�ؚ�6�<F�u3�:�L:LjQ\.lB���SVd���Q��\&���40K-�6\��������8�1l<�_��
>�8��G�\�;��	Vx��s���A����T���)�E�&��D�Cq�=&���4��5_��Dl.�LW�c�Wӷ�u����Oi`4��'�ZS�ƶ
̙Z�)�.�J�vL�8E��uSe�	1���R�˒~;7)�{��٥q�{��eP��2'q&���� �\�!�B�?;f6��^�]�0D��{�%�rH��bsS�c��f��v��F�xʳ��x,�EM�Mx˷�n�I
��p�8�4a�o�%�+�VPM��~��U������s\Y�C�זj2�3ՋzUfm8�}byZ�%u���XY��(P{{l�o�ynW+�|so��ڱ�pI��nb�	��D��u^8=,��~)��?`pN���^]�꜑�0�J�.��w��4$�M��ʌ���l
m}�T��A�%��8wދ��\�=����s�HLʣ)e]��|*�z����/]l^�W��w|P^1KHN�̲S<S���5�D&+���}E&�U8H��.Nfϡ���^<:��/Һ :�R�}��s�4&Cv��8ɞ5�����FJ���&><>�WC�s��B0����bP��g����|֩�$���-` 7̐eq<q�fu(���b6ҩ�>�۷���K�/ov
R���į�̑Fg>L���h\�.H#q��,8�T~<�P�D�1�w��B��^?�N��G)�����!��՘%��~3�!���Q��t��,�ƪnn�Q����lf���[s<дQ����4]}��@��{���Swl�4�]�hSh8\R�������/����5�Oݡ<�k�2K�.�H������:u�����qF�n.1��j7Z{�T���k�(��Ln�3��:����h(šmp;����]L����D�'�e��\�ʬ�2m�V,ٵ�5�3_�v4��/Pq��<>�vG�N�{8	.�T��3EE��M�����I��Uf���R+8���O��|]�57Rq9"ƅ����M��ᕒMw���f�M�5�N�^��_d�k<'���e�AC�Hʇ�L�V&lƀrBm��������o��x?�I���(�_4��(���Ǹy��L�N�9Vo�����~�&�îN�k�N&~��}`q��{t����|>��D	C,`�:��;�3%��-b �p.tۙ��y[xx"P�>~���͝]��p��,��"�lU\�muG����RI]zc�^��;o�N�oɡ���X�,����`G��jJ8|� ����9��`wOAў�&��M*����"վ�1Q����(׃�8W[��	y� ���4p���u5[����m<�,�����ǚ��<Q�;Jz$A:����^��3QO�U!�[|&���?�{
���X�3J�d �U@����U��/^�E��F%�I�m�t+6x����<�bO��S-�s �:������.���y�\�F݋@���Wݤ8�F�����^"��=ǉ5�V���`11�61[>�	����4�v���莯�L�YdW��s��@�`l����IZFD���O?�F��!��Qc>/��-��d�|/Cn�4�Y��~�����ު�%����ܹk��\��qAꘗk�wy�����g���&���҈�p�]�l&=�u~��ww��Xxϟ_��ʒL��G0���4o^	��4a�1\��c/Z�R���@�I�m����2�ڏc�p�l$z�����*�<��zS�c��Z�ۥ��*c��x�6+�VA�������]$Ɉ@�je��?�������a�#��`s�Hc4T�b�`P�vK��h��p����b0��A�cŲ�<�C�g ��tw�*�E'Vk5Y脥\`��N�H{�S$?�����P�G#�����u�Mw��#㉅v�/r���x}>��)�$/;Ħ}
a��nJ��41�ߋ�5�:;��\��6!/���k擟��]v����$^7�K�k`Gp�^K�����ī#�w�|��z�f�<��4��Q� ����t�h��K������뱝�mv-����O�[����J\֦j�qe�W4��=*Ni|����M4?�L\t� �F@�S7EM+��]�=1-"?+�>p( ��V)�h`��|d"��-��t��p�������/�^nV����R�<�r���3�I���cv����3T�f�f�jj��7��/9�K	5�ㄱ��i�~cd�t9?�5:��=S�� ���ˍ����=�b��"���3��$���)�l/:�)KM�w��6�*��hś�W�E������q�����̊�a��GPK1\K��j������+���@�%���}��ŮP��*l�,SG��_o�rT��xFO&�e�k>M1�������$#���x� ��irK�i��:%ǉ��(P��"�E%,�=�ׯ"�~���du�w��<ܝ����b}�^�=�$���SU���yQ��w�¡�����Yt^k��@ng�O�n�K����b���/�������)V�F�h�L�wqm>?��L�A{�e�����:4��P_v�/a���f�����b����?|�X~����M�>~�ݻ��������ԍ��I��0+T����fyX3̞�U
�T���3���� �羞�0Y֪��9��ɐe�fծ!�	�6�|���6��ж��u*N6�cIK��hhk9�8��ם��Ǌm,�m�R1�AnM3��A�C�K�D��&���?8c͇��]M=⒬�����@	�`�z�����j��n�k��]V"���f�.7N�����t�(گ���[�H�.fu�\n�}�&�������}w�~3���W`�_�H��\7�Y�y�����7�6���pKqx@�V �}�"�	"v�)Ze���?�x��=.�X;�Y��f�r��b4/�����U��:�[u�Blq]YNL����{PHƪN�tO �}��G����^T,ݰ������{+����C`ԁ�{P���_5�>e��f|�;�Ί��)u��Ty�����ٷ5��@zd�0WQjdT�����H;������������im�~����M�.YC�����u� H��<-t��#,��{�UN�!��ou�o�N��h���i�b���>Ӂ0��>��-Hd�X���!4�σCy��Yk�r����#�Z!��ּ�4�S�&�c�{�;@���е������T�gK��JtTbx���ɒ*�e�����!�%��鳚���,v�;���𹑑6��w���j@�Y�j��*��V��d���d�۹��EЯ׎����%��7ގU�\,_�)xG�4T�A�>nH`:��J3h�Ϙe��\�I�_n)p�S���Ţzg��N����͘�x`մ�EC���q!g�����h����A��c|d.�kӠ��*�̚f��)-�ۙ4�ٓ#����st!�e�O��0� j"�KņS��7����E�Π����7e�j;�כ�0�#F���&b�!���:�p8+����O�M��B+��[�+{M��L�Q%�u6���7a}��53�,\ra�2yS!w��w�d��b���n�Q�_��u��3�롯���A+�Ը��=��6�L�z��H�7���-L\��~��OA�rύΩ2c̃��\���-t~��[�?/�����o�u&�	���[l�t�〴ݲ>ST/C�D��rvܰM�D��K��)~���ߧީ!��ڬ�_�Y��?�?�ROC;�������\�a�M�\���_���ߊr�.�Gi��-F�8U�;՛���E�8&K�Y�)T�i�{�4Yƾ���Y3髀j�B`�s��j����bsX����#��\���΢�+�'?�^�s�DVWH�Y�׷W��:Z Aw���������:�Nm��44S�-� A��ry.z�@��;�����AX� �|<G�*m+�/I���Olq�o�5��G�H�$[�tvsD��_^r�r���+��@AZ�����#X<P(�Q��i'�)�����kN��{v��(s!\.�6��(�ͱE&�������ǉ���ʦ�y�4L���G5�o+"j\��CC�V;���5|��������{}�+i��l��I�ޒ-�k ̡e�~/x�%`�G*�������p��u)ֲkBM�/���Z9��!��:ߥ����YK�R�������S�'��`�E(�pl~uƸ菛���H�!�C�t�}W��V,6�	3��C ���}�(�n�ΕH���S�ʓ�;ǒ�sFQ�_�W�Y��Sd��B��'2�����Y�Ƞ_xn�8�K�4섿RG��3�5_�y�1�����T)����ܫ0�-��Q`�L�]�{4�.���{� $0�@���>x���-:�8Hx �
�]ⵝ�����j��cp��{�F���:!(,1Yrk2�i/�~<B:�&�?��Lenǒי݉�Q��+�:>��Ǻ<S�
%-9��<��Fut��Ŋ�K�+)Kl���GY��\NҫJ��'�Z�����6:��ߢ{�2v�s�b��L��B��3��W6�S�����T�z��B��%1��]���oB�B��h ��U��YuH-�_��A,?�uͪ����#��`m�:%XǨ�e�?�k�av	Z�q�n�Y�-N��um���{g�O]�GbD�AH�:c��L-e���%���FP�A��`Zt����N �X-|"n�yDc*R�wC�$���q�r���t��i��R��*6���cMч>?e�N�Ys�z�jW�MS;�^�!.g5�c�ח� 4	cG���M�1��wlڟ�����\��	����Q�?����5n0��#���^���������x�Re�|�y�y�r��1��L�^7/l�km֔�YX~m
���kԶi
��pP��&�*J�-�[�[�a��(S�*V\�k�Ӧb �
�>Ȃ�#CD��z�{�R�e��t4�ǲT�Xf6+gޓ���F�2��&�w�ѿ�\M�'T?�Wa>k��P��8כ�� "2ʸ��!���[y\�L��5�����.�� �X����/�� @��<q>}��;��y����jθ�5,��Z�������'/)g��U:�U���WF ��51@���z��$���{O7}	�v���KQ��}ի�M���'���_v��&.��6"�;2����K�z�jHO�N7'\h2n{�\x]N��TZ4�ƒ�6����6�`�gF�f�ϱx�i�#�^@����w�蘃���������#�{��mQ�4�>k>_0 ���L'�h��
���V,��	���D��F_����/�����?�Y~����`�=��?�9���v��>=��S��'��15������q.��m� ���g~����#3#����SN{%�c��5c�|�8�V��ٷ'6�T������c�`�?�)��*m�����r�疘K̇{|�{�s�R��p=p�����5��~�k���1��!��1��u���G's�z�*�8��N~��yM����X�ޣ���x_�sֆ�PvN%�q\;`�ͬ;˫H|-d���(����",�A�m���X�s��0����s~x�U�b�0l���jm\V]԰�^m\ԍ��o=���Wu)�=�E��)�kIa�
Z�M�":]ca�1:K��w��+�Y��]bq�@�8�:�<�izƆ0�Z�I�� :�I�E��|��<�aO�; ($�������w��(������~*���=���'6,��	�����X0�$��.V����m+vR�B$���)�'��}� ��SN�,3�g�od$��Ս�,�v�Ɠr�׭�T��w�E�~QG]%����8��%�0|&���uu*�J�溘)��˫J�؈�:M�T1׮#��VEur�v�|^�*a�%�㯏�5���]mg���zg�7�0Q�&_�=X���9�C: bMvv��P_2�zϱ�G7�+8�
 �f�m�cf��6�0�`�瑱��q�r�%k�����,�G�9���	���d�:*���4�Y�R^����@m�'�}��H_4�*��h��-rͪY��٬<�[���G�ϛK�7�פ����ڶ{op�ٵ��������E���KM<�P��p��7x�:�jw���8�E�-*]��H��9�l��cࡲpF@���I�S�_�I�ۿ�[|v4���U�7�A����l������_��n��7�|�Iq\����*5ԣ�~����������8'�u���fH��>��1ex�)��x���ه̢Ln��R�R��^>�����葝]��.�*M�n"��P�E������\^OY��A"+����|���h~%S���f��M8+�[�y�y�~�,iLݴ��%;����!�4E`	]TK���!<=N���������R�U��9|T6K�b�!59�m�
Ǭ�|Q)��e- ��^K:y*�wי�!����n��Gwj���((�r�Y��Gr���4Y%J&���%|?T����k��k�VA4��ac-1��WϲR���X5��A�3��Wm�1�Z�2����m��X.r��D���{�*,;ݸ��z\o≙I���ԓ���	��H�u�B"S�s-j@�ۺ$%���Y��ɹ,W�@I+�^��eO���-�~�:W�L��?&@~,�!��OG�_O�I�S��eׂ�$�˯���z�R8�۬Idſ��ׇ���)/R�)��u���E�bdsX��6�lU܇^gH�	�����P�A��� �&`�cs�@C�<�'�e��[�e�������>:�H�g��;�V2�i�հ7�����(�c|��msbvQv��+mQn�1U�r��R�u�=��iu-~2�E��>�����*�	x�ڕSfq�����:p�جQQT���,!kU����+=_s��0���^��L�x��.�A	j݄�>����ۮƝ��zQ��|~���u��)�>�D�K�D|Vi�>\����6X��wod���"#�Z��S����7pxM �|�7^�_UFT;����n�]�f�V7&O�V=]1(`�������M��h[Qt��񧼁 ��OkRglMRDU�RR
<�_ڑ#���q��'�<t
8�@�s	������w�>=�����G���"�������|�m�w2=z�o�MB �t�*S�G�ʇ�<��c���ߒ��@Z�G��\޽{_>��$�G��i<EP\%��MP�(�3`�.0p-�Hp�L��awq��~���-��s< k
!���%���d�wg  ��IDAT_Ш�k�i�C.R]�.��;�lz��h���Buy~V|����$�Fx]��n�k�O?�����=:�/���3\ҳ�=��Y�\�!�[��ά�P�(��KK=~(Q����߹���z"=�1���0���ܪ�3G:HW���cu�p_��K@�[�Y��&��>���e���>��E�'��vi��({�69��I�ڌ�]XzR'������W��(�  ̚�i�vDddՀ��j��bLw������ps:����Y��� ��f�2�+k��JX�)��1\�3��,�*?�2��Z�f�TÿSPe{�1��l-Q5��jZ���ؗ�h��X#m�W���r9\����0Ͼ� j�wY�ه��:����0��[+��>)aF�R�mB��5�����������4�ꥩu�B�*U��A��E��5�u���纋s��Lӕ!,�ACz�ѷQ�qS���;^#i�a�r�=i8�U��Oz��^��m^�i3���X~��O<����Z9�E(:�h�u�y[��s��AOCva�7�s����<4�`8aDϸV��@}?�S����VZ߮��d^�,GT�l���p |�w!t�X.�F�N[�S�!�Nk\cqw���z����r`l�Ez�<�qhO�~*��	���׏���}�~R<8y�cb�P�ق�Z���8�������B�J��'\es|x�[�aq�t�O�����i`�-Q��4��;"B����ҁ��o9�5��j5j}�_$�D/3�c��㐑�_O��3�x0_�	5��'z�{J/V}ZG�UF��Hv):�0/�P��5��%
M.����
k�v���ѻM�|�v�c�pbWic���ڈ<�RJ[�����k��T�Jb��s#��~5|��TW|��M��V���^�C˚a��l���l,�r\�a !����Q�=��hk��U�8D9�)�X	Pm|]��w���1D/���^
������=1Ϸo��t��mhѪ�Hp��P-ߞ�c>��:�����"�.��w�6�?]�A;�Y��<G@҇Ioj`V��c���Z������eh����B��N�ϛ�ɀ�n^��ݳm��J�ghO�B�쐾8L��Z(s@C��)}|������z���=Z��3�(�%X]CK�D�7�J��q��c����WZ�{3͵����[�8�-��l(ׂw��Wm�L���1�R#C�D�>z"]m����bRtQ�����$��m�
>"�a'�sG�.i_���޴Ϋ�s�!�]s,эb-�T6�qA��N�sF[�5j05R	�d�d����ݜ�Z�/�&�%����B��*B�X��`!�~��ۇ�Q?������V�|K����0���k>МŲ��,���O�&Bf�Ui <S�<3A�]`o}��d!��N@R���秒���l��0wiۂ���]ވ�"����NŜQ����@��Bch�V~��c�05�?��c��!��u�>�� ��Kr�3���"Qu(u��k�������"N���,�{�|����e�Ӌ�gHTUR8�/�Abm8�'?��>�������F���� RQ�F�eh�띥����-�q�����1�H Y���мL�Ơ�*=ku�x���R\A�{9��ɋ�flL�U�S�J�D�Ё��""gЪ��=��9�E'o��}
# ��һ<�XsH���P:Jr�D�W�ċ��&S��0�bոw�k�o���� e��5��|�1ͬN��	%+�1j؏�j�.�^�B���je����2����߂M#��K�}�u��X�<�-@�^\�U��<s��:���G`���u���ΐ��o�]��9	�-V��U�W�`۰�4�,5NƩ��>K!�@�z3 ���kp!�Pp�.��ʎ^��ɖ�����^℣!1[�T��8t90�9�$s�p����}L�;^#���=�z��X��E��pX����T�Z��=��gR���HZ��zp�:P��%�3d>��8~�ˌ���駔;��O+g�s[��q��Z&�c_�yh"Q��`/ң�$��$�7o�D;�}(��~Bj�mi;���)g�un5vG����i���lr�Q��JUw�-�K������T�ϓG����a]�tVc�9�aHo�9���Rn2$݂F=�������z�\S	�]�~%#���l�51m7�62]�5L��Y�o�#"��䪟V�6�<ٖH�{t��v�k=���9.	�<0Bs��0Ta��Nh�����H�9��<C��#X��cZ���ђ<�4��Sf)Z�4CY-p�Y�tu��3�Ԧ�72�R��J��cyh"Xl0��lt
!]���;"�K���a��Pa�G
�pa�O�S
�ڐ�#%x����ft�G���P�ϫ��t��8����d��Io�Y�J[�15+��6����Ɇ�;�#���D�
Fߏ��_ߔ7o�2a�k���4�ǌK�1���%؍ ����m��u[�2�&ч�o �_��h�������},o߼�C6��_hH�وZ�׉�%��9J���==���p�ҵv4�E8��KB<(w]�g�7r4��X)j�H�X�S�L,ѻjI߅��^Y�`R��.E�/瞆\s������c�j�lޯ�����lc���в�Y�Sb�ɛ�^(�[��|��L#��(���e�/p�.���ե��G���ɋ�6b%�Ĳ�����Y�����^,��AY��d^G����0�kӮyA�������i�K�d�q��\ȇ�acʠB4�bPV��rs:UHL_B��2G5ԅߤS���N�X�㶧��>E�׳3ͧk��⠰Z}��k{MUa�q�|��ey��=�(`���N%�%C�2_�w�Sx�"�[)~�ČX�
+�!�œ�g��-<TP��0l� سRk�-v��P�]�N�����w$�[�B�5�Z#�Φ��Q�Ϻw�QBwme��~L~�zA�R�MxV+6QKF�Tq�\a24���Kf��L���\Yk�li������v�MIl���G���碽Ū*�l�]�2K�W�J����&i-�O�Y[o_� P������2��~��Wrc�>�hZ��f�@��u=G��!:q��2�K*�m��V��8e�9z�9Z��}.#�{*���n���՞Xr�S�ut΢����)�I�D��%W��d�&1�J�xw�8��i9tŦ�ʘڀ������#�Va��c��`+e�@�~a��XG�9#�z����_�b�Ν3�V��������8+i���5�-��	(����Wϑf�Z�8
��&�o���^���k��I���9���	�����<D4?1�r�b�GXD��jD�4K�ɺ�,��G8)���}� �Ђ(K[�1�7 ����>�p��=��҉B/'~��ç ��)����(�}��q���Ko%ޡ���a0���A��yd�(��\EW,Z3���2lK�Z������ e(��_l��B7�eSC?q��]���(t^�w��&ץv�mK�f��s���z��2�䎒��(����224�e�K6����x�+�B�e���wFJ��j��y�l
�3��*N�/��c�����_��^�#�C���~`/��p�z:?Fbv��}n����Y%����1���^���RNY�4�W�ZHs�G�~-��ڂ�����w�k�zg��2v�c�,<�-�<���u�P+:G	aU3W�UI��9n0���C���[m��-��Id�1���F�L�,V#-I�͕&�F����ҔJf�?�-���S�y���'d�6�MY����J��)/��1q��<��"�ڦ9����2��õ�:d����)�t��/E���.�%��j� �~Qo�%��0C�*ŉ��g�O4��Q��6�{�٨����b-Xm�>1�5� L}�ف/$pQ%E��i���u!�:�1����{��C�!z_ݤ'���?(*�tű��A�	��H��OJP���3vAV��p>��ċ��LSRo�uY������g\[󐌔L"��B[w��{�@?	ۭ�p^B ���ST=�`��"�ɸN1vMx�59���H�������c��A����q�>f�11�$�*���w'��ݗ�f���	���k�n�Ҙ.���&���1�+�������V׶��������͘�O�XXy3(	�N�U�xj2�F/�Tu�2ɄL��+uc%�a��Y���BV�KϠ��������^<	u.��O�՘�JC��� އ��H��O�$��һYU6���ƶe�|\zf��J���h2꩘<����̔��W؏��z�U�بv���۵�����_)��.�pUתr���W�~�p�*�[��Mܖ�z�,Xm�iB��nf�)`�ǺR5L!�(O�!�|,�~[�ʱX]n��D��P�%��mMFAS�_�\�ɳns�H����� ��:/E�B�5��]�$7$���X��~�]a���K'�(V��q�A
���)J)MΗ�V�K��61�6��S���5�3�4T�
Y�^Eg�r��l�2WHep �8o�K<��a�pЁ�W�V
&�Ǯ��~��ג�y����ʈ���<��_gHWc�/M�a1f�k�}Ye>|�P�qs�ͅe�
"���m����)Ú9�jN����pg�%���dh�W5o�"�X��0Rߍš�z_�*.��<�VR��+���m�z<��!�fL�	�gS�}��������%z��ɝ�4PVvghop>�t1D/r4�rz�,�;Ѹ"q��%GQ��cSx��3��k�9�җ:LNJ`�o��>&<��1�wl8�e����݇��um��㰁��K(��=����]�]���Ŀ�mRoe�=Œ��2�1�u1����ܖ�} >-�O����B��2�X��	�G����f4���6��6������u:uU�:�3�w?��������ݽ�O�At�ct��Eb�@x|�]i%��t�:���h���&~�;sn-�]?F��4�5ۺ��U@�@��h��>�wR��ۮk���h 9F�1E����!�
ߏ������S�tLΨ���^P��<m7��	�LU{ DŘ�ܜV�4���H?��E#��;l�nh=G}��!���z�5Sr�������o<)wͬnu^~���o�-����l<$%�ݹ�5���K����tzg.�.�� q��Ȉ��3'�NLюRHc�'�������Ǣr�fեx
=�aȓ��0)S�Ds������C.����4���V�tzJ���ȭP���!^Jk��Q����횝�Ŝ�۪9��LE�#��=��f9�}��x��d�qm5���{yՀP�]0�7���f��4�ZIj�'�X����������0�}]oݪ���9�c�}΢"oF�qC@ᕺ�����1m�H�V_޼���ٌ!k`0n��
{�R�O���J"�'��a2֭\T�|z�QX#�n��*��O�mU��rr�
��j�:���8��t,�џY<Ğ����X����r�2憮���8���@LP1!*�ҺZ���!mK���X#������1mCb..A�������s����B�l����1�p",����ɫ_w�4�����H�x����ρޝ) ���ՙ�IτiO<����u��K,�p�b�t�ߎ�CPO��f��S�2�2��Gڐ^.ǀ'f^g�
���.Vx����2,!Q�h���Ю�f�(2��G?| ������c�4����V��w"��:�yyBw3=���]������:��q,q��Zg�G�''�PFr�9���2W^0��݌�{��kߪ<�	��sz,b���2rAU�A2��e�����X�sr�}����gS7>w�H�<Re��������`�Ix���421���n0"Ps�o|�Bmp�=m��Q�MJ=b�݇�����1�w�w�R�P��
J�j��Y~��Hh��+x�������( �/��yI�W��԰6�H�?�5��[�<���������mmC��8�ܒƆT��!���>l��{���'a���Q�Lkn[�l�I��������z�w��29cL��t��S��n�����1m�Yu��5�n���zV���k�DM�YKm�����`eǝ�L���qc��n�M���w�0sU�,G�ml���8_js/���9jȷ�eس�jj�[��P��+=OʥV���~�S�G]ʰ��7�C.��=��B�?0��k��V3P^7�����x�����4a������q���g�uP�(0�y�����Z]���U����t�\�V����(�Q�f�K 'by��l��܄��rׂR$�b耇c\�i96�)�8Q$P�}���p�ǥ���w{�ڠ�^�`��5'��,��C�3���b3đ��zꃱ}z�oxBo�W�e�o�s��7�����5�~�%9���C3�����ƻ�5j�wN��U�I�os#��5re����G�%g��O���Z]iʝ�JͶqLW!�Lvt�A�b��Q�a� ��c�8��L�b{.��[�T"b���OYI�����t��_.j���'&���]��k��6)U����po�!�hq��XO/�P�9@�����[�8פG�h��hLˇG������q�5z،��HI���NGʔ���R��h~V�E\�S&��{���{;�@�[��J%tk,N�M�,/��u)kz�N�8Ӌ��|�j8�s������](�|R��50ג�K������Nԡ���Z�^�*��)��2�=;������;���r�����B ���	"��R'���������=۸���y�,�&���iYU����L�؋�Γ�}����!>U,��<�)��Ω%
�*{��X��^�U���:�܂���F�ڙ�i[�"�+�٩��&�����:0K@a��'Lk�)>7�y�����9eb$��?���)�O�"�d���լ�9��Z�A5���0,����;p�JQ�76���,f c�0�������� k9� ��3{��úm�����%���%���{���57#��0��OO!<�D%�H�����1����.<.��Z�!=~g/X$���h����ח]w���w����!�f����\�-���bv�C�C ݡ��]a��9fcRcz�s���bdY�^^����Z��!�+������bq=*�84Do�����"K��J��2_?_�\ǁ���=�'óF��B��J��V_�꿎u�IM��W��5�IɡO��NF���ܮY^i	��#Iz��k�]�.�s'A3����5Ԉ�Q<̉�w�k��tH�b�ϣ�����Kp�������:P��1�]�N_�;���P�P��w� �AX�io��ZD���V�^�(��!l����	�6�Za��bH�|�OY_�� 08۟�jh0�ZI�5eB+�,��z��ga�
�t�&5�]2�b�5�/i�$66E������Yi1\�g��-��'�!|�:���j�γ����
�X��dc6	��Ճn=QWx�K�.6��aq�񘇉�������	ä�x�Ww]+�Sj}t�P�Gc�U1��iѝ�sP}���L��U0��r^��rD��G���j�n(�!#��8M���y�P	�B�M�y��ɨy����^��"�GI�"�� 5��`Ms����r7���R=�n��~!�?uC@#ԒX����z��4e�Z�B�]JK-��ژ����s�r�+j@5]Iυ'J����u8��L�
U��J8j��q@8%��n�Ʉet�<t]� �߶n>�W
N�����z���Ҿw����D�����t�rm��f���^�ǟП��y��!͖a�<W0;ܩDMD�K���%[�Nzx������/(pq�%��U}�m��F���8Gݲt	�w��1���$�D����(��Ĥ��"$r�W&������(�[���Y:�?�uL�����ˮ�o3ε��U��"~'Nɖͻ�}�ډ�ΦV!�Oz�U��Ɋ���B&W|�3f����:0���cؗ9��;�A{�9���	8z񥊱��UG�N-6���Fu��|/_�q�_�	A���1'W��C����ǽO���'ەz�.�'+@-тZ��DǭJeϹD�ob��~��T�@��'�C���'m�Q|�4�+�Bs�{�D��*��9�����ݻ�����D�g3�`T�*ϗ��]*��7uo�*��U�}��cG�f0t�&������e����9����,��.]�FѤ�R�]��5�i�O�걷��jC�?[wt��1�1�����d�»�Ø
��!���7*�0��'�;,���ݧY�/��2{��uG���P
��H����8��zm�ſ�"I���\L�$
׼do{]>4Fw9M�q�Z=G8=dr��,��ܰc���X��k���t<{2�Ui�͸squn�ّ���#i�h 3ҿ�nT����$��MWңv��U@G��`1��/(\�S]P���G�>8�T�%#��$BT�������&�	O���{K�9����EMťU�G�땺PW��^M�iH�=��w���}d7�	���B���k�R&C�z�`��S��� y��n��ZC�������t��z��>aER���?ʎH�ͪCa��#0xV|����u^�׆ԥ�6��)`�<۞(��{@y�(KK�#n|�]�+��(i64U�k�o��@��a�D����K-��t��׮4F�όi�	�k�=��BF�dh�厣Hףկ���Ah��_��D,��֚�9��0�_lO�o`p��r0E���t�E����6qw0Mj�p������d�&���o�F�@mA����Yױ����0�%��*�0\a��O���#��.@n�(o�>�b��x��J�_�,s��w�E��O���(kJ�����T�(H������^U@x/[
s��������a���$�3��"���%E���Q�z���BQ�!���8��P�Q?�~�.y�^쵕wŏ+��U7�+�w5��;缃!�rBc�UnΆt�����ϥ&I��lBK�}���x�s��a��3���yx��2>MkpX��!2�P�"��/<@�Ѣ::�ؓpl^F���W���J��Өu��R$aH_��"qm���K�z����)���.�Ϯ��9�lR�e��=�-qb�b!zXDao-WӶ_�����'jjȯ:�Zٔ�=��$�^^��6%��x�zb�7�<���6�<��$���0A���qی���8�. �Jf�5hCV�M�����@���*��	RO�7�k�ͽk)3ƛ������:�̓c�kRk��U]|�s��ѳC+���g��DSN75�H�BS�c��D[;l�k�5��YO���0v����R{���7�Cra$�������W+�׎y{��9�[�2�L�Ҷ�le�w���/�B�Ob����Cm�k�l��*�����_���^I�5:Td"�rn<�� ��4���t�9����x:���˗/��>�����.�S��#�]�t	��EF}J-Q~|׳��"�ƹ��Yg�a0N�gL`>| n�!"�����UF�o?q'5ҘJmU>GnE^5�6L��]��[wQ��h7�$ݚ�Ve����ǅh�M�&�mV	��L��I�r�jﲕsTҕ<$��uؒK��ޓ}t^ך��J��n������{#���x�:����k�ȑTu�*��O/".g-��Z�j�{Jqe����B@�O�qAnT��Ss]����I��J1b�@��ϥ]�MqfZJ��9�9���83�	���|I��������ʧ��vw�����y��H�ϧ�\�]�iHc,��]��q��=#%�'�(n�=P�)z�K��OC!��WM��~a.$�H\;�H�/�� P�P�{���w �B�/<|���a�n���g�q�P�������x�?�}��J]�}*-�(�h��)�xBj!})�����ﶟx@�}� ��J��i�5�Iu�s&��?N�؎�/�W_}ɍGm�O��[�Ic��ׯ^����|��W���k?�'����e�eR�ٽ)��Cm���u�����.��To�
�"��}ˬ9*!�dX�)o���W��h#��*�u�ϑ���u�)�
ׅRS9���6��=�܂��Ҥ���5�6+�;D�3|�8�I4I]W��ikT'z���*����=Ww�p1�"�h��N|��a\4����reL��Ue��1Ғ�hkH�&�8�R5�s=��wt	2�1��q�}[x_}�u�*44�]M��\�����	��a����m���ꟺu�5��}p��r�նa���C��-�=7!�N�����Q���W0�w��ײ�a'��3$u��}���<�Ż$�l|+�]e�]�s�J�xw"[c���-j�c����]�ɪ�H栖���7L�`��~m�%�hxP���R$������?��C�����c��-==�5�ȗ/��Y���_��	�����m�|�'�bl��#[P�t(�`���`����7R��q c�E�~�X�~���������ͷ�n�T�i:�p��хa�G*����J?vP��4髰�f����p�g�`�Aa�h�Ib��ZZ�����s���������*����[��Z�����X#�t)�|�� ��ƅ�~sA 0t�h��Q����Ɯ�!��z(gY����8��:�NnEa9�*�x�EC3h�p��%��hXG촓�헵�R������#m���H[�SM�T��{wz�UQ`1�*
�`vO;e��mqCe�� � `r9eE�I�fX>���x|�a��w���x
��'�0hC���=�B1��){0�t��D!/����}/��mzk���lP��z���0����ؼ�W�!�a��AV_|>\e�aX�㐋J��$"���P4�ڟ�_�
��T
۴�&C1gn����Eu[ASwA���W�%;��q�Yg�U�f�Wqp�0�	,�F=��p�].�|��a�JDI�A�e'գ'
Z��1�	hi��st���z�"��q���2��P]�z���/ʷ�~S�zyY�R8��!g; k��^��"�b�c\;�lF��J6� �^�ܡʧ'�GIk/Q=��a��%�X~�1�ΐ<.�p�D�o?F�]p��e>�������f0��8fՒ�E\�[����m�ђ�K�:�5�Gf;�jw|?}���u�ϕl^$��NU��5����{���o����gF�?��!5-��T��>}\k���'D]�>)9�l�IG��-<p(����`���؀���*�<+�f�&�s�$���"�%�{R�N�FJ�m$�/7�Em�2�<�ȅ�V�ۂ�f��R�}���nO��x��ó*z7�b�R�����&=;z�x�p��������O>D���`?ܑ�l��4(������|LӋ���-n�
�p��%ۊ`�[?�i�����kq�OO�Hor�s,/mB��۞�|�Uy�
$�G�d<�	�A����z����67����KW��'�~~������'�#�u��e��'�b���;#Q�B(*�Ǖ�f�N=�����:-����c>��~��.��rŘ��>qP�6C4X�T�ڌ>��iN��⋢���������#�051H�J/wc��F�R���)o�'5F���>e�ɂ�(C5G����n�����[���
L��ҳ���]U��r��m���3v���i2����j��1:
Ko��\��V�k�1fw۠?��k议�?39թ�s���0��_�!OfǢO^��f���=	+Y\_;��B���ә�"�G������I�V(qCC8�S���5����6��L�w(�c�L��=qx	u�L��C�x=�������y��-%���O`x�����C�F������X�\�0���$O6��leN"���L��Q�Sxg8�C0�;9!u	��j90�`C�s��5�]%��m1��!D~��{��ڋ��.��g4��5�	�Ib^�����_���mPU&f���n�b"������������s��"e�5[ ��a��`����.��g�ox��ާ�u1#Fg�7�4U��H��>S��D��,���5ƾ����oޕ��OYb���7���1_���R_���б��3�'��w���-��_��8�L@)�d��ԏ��ʓd���EG�Btao��񖒆k���98<n��0�����#����b�W��z�:4�<4���������0�CCO�xf�""`�L�~N���ձ�r[�;�F�RѠ�����,bM|�����<R���?�[&|����3܃�6�JH'�UN� ��0_��摾(?��3�?��s`Kj*G�8��Sd�JcDC`7jr�km~��a�����E��n����%��6���L��[G ���/�Bd(��<Y$#�PN����=�`�x���J~D�v�cC��Ʃ/�
?��MP�W���N	�ɚ�2�$��3�����c���������n߉q���#��?��C��+(�+wm=�U�q�g��v���[����曯�����{;l���T�6f�8��"��z�ۘ���w�����ۡ�[��`���o���-�Ex���w����c�jlH����]]���5|+A�w6����&��X��`H�G
CzwI�1������5�g��Q!�-��������ٯ��e�|�T��<�`������ �?��Ss���a����T5X%������P���j�^�8<r?z\��]C�N�xb�=~z"�	�] ��tD?3��՞j���􎸌A��>��I��8�]�$��I3?�� OQKBb�lo)��R��*�Mll^�+�6��+m-�X��TX��K�k<���Ҿ!5ϲ>�u"��X�lU�.�CK�8W�{�h���M��;���������O����Y�iW�I�QXNp������������[.ns���a�J,d�7���81<�!`b��йD�B��RxxJ [�%\33���cL���SP�;����=�܅��L/Ix~��İ����n!���=���RO+`�7I�Q��MO�x�3a� �j���T�_m�A�T�N!}&Y�B&�#�x����������eL!�|�������W�y;�9�=�m�$�o�v�)�2�s�D<<�c񓚧��J��m^8�>�dl^��*����l%8�4:����Ŀ�#����q�$�3mX��3���k�,��?(��蕱�r�V��ϫ��I*eE��F��I��%.
��:%����Ն�ɶF�U`څ.q
��c8-s�0�����G���!Q�ͣ+jS\"��=�>�a��}͸��ۯ����liS��_X��W�xCB�;X?�����CgfhCz
Bl	�ƈ}s�!~�7�E"U��l[Acל�|؅Qjq�.��tڻ�1�nCߧ0�]�J)3DH_�R1� ���&{)E���*p=dT�$���"�vOh��O���'��(N���&b��fdDeP`x��Hw��Ϸ���u�'��t�=��q�����?H(e�K�<��~��M�0������g�7Y.�y��p{;0���`P�w�L&�#���f�%\l�%a����~*����f�ߒ��7���J���ű�(�I.�뱹�Y��"R�sJ��f3�KV�� ]��������)�m�١w�ד�}6�;�B���!r��pTDL���!Ն��^x�(��ݷ�rnp����?	�`>�lp3��5- 3�ASO,������N4�ǧh�3$s	�~���yO�$.%�2�O�<3����(����qfS+\�Gy��Q�{�����X��y홧=D;pU/^2��Dqe�V5�s���}'����[v����:����ꚗm*C�Gԧ�w���Q���/�?O�s�j�^֔wC��P�ޱ�o	��
X�ǃ���Co��BZR�Kʈ����ݲ���+2-H텅=���^R+S,+W"ܳ!�6��@���8���/��ɐ�l���Ķ��&���0X����Ɗ�[^��D)x�Ґ�F�a�fD]���Fx������1Ï���矣��nbsQM��w�&���維�ٷ��[mҳ��慝�O�)�c�~C�=�.�l�8�0����e�;�Q�7
oM<�[Q*�/jA���j�����S7���:�&��"Arz��`�����<�o"���p"�]m�a�����]%[ԓ]�(zW�3q�/7C��������s���'��lb��t��1�p�w���Ɯ�E�Ѷ�t����t�жȁZ����=�2Bez��n��	��K8$�N?��N�� I�zH�Ť�SP�B#A��6jj* �?+j`��,�,T�ȑ"��<P\��H�uW�b��|�.%�ҹ�=��ӧ9����xCȇW�b����M�\��#���s#*�o=�L35o��Mڪ����P�«p%S����v�&s
�ݴ*W$���F�5�����LцbYݭ4����U���E��y�Hr�C�ñ�:d��gy
j�2h�v۾���9��C(�/)ʂE�:�{�yz��D��4�k�*�w�� *H�jt����Q�y�������JZn�Њ�����8��WW)c+��I���cS����ƌL9���N	���W5�T�!���~N^������R���U��eZ����	��E0�h'�V/�������1Ϣq����7�D�uM]\+��Ç]�B؁��g4�싵����x�9���ڄ��L�������'�Q�ծjO;&QJ)�g��5��e���\�}{�4E]QYEX�Ɓ�����������(J���58,�]���l�:F!�iU�RJ\�Tқ2�-a�z������ΠC�r�+�sm����"kae�` �B��|iJ����n�p�M�}-�S��Q��l�5��pMFNk`�L!���=s�]I%�]Ы�.p����ث�Q�I��c$~W׽�Њy�0�}����7Uo�s.J�kE�ffp4�.z�8��d��wݛ>#�0��A���Ccdq�1Ĳ�!�R��K�^��*����f`��_�R����+b`��CӘ�{�=WrO�!��k���ay�L��,�Q)��������XC	�Cc�X�����_���G����`(��bN��<��g�u��¸�;zL��M�;6�8�wi@��f���Y_t̶��,����!6�ˏ�u�]��aX�	Ǟ{|RKo[0��pI'�N���[>�e�Ȥ׭_�3��pm���{]*������1Λ!c����l��M�>�6,tԻz+.��=���+�^y��zi9�u�}���Gg�)<��ôL���,���"ؚ���K���ܘ�����[�NY�p�/SXp]A߻��:rJ�?R�@�$n3��!d���A����X�Ŋ�0\��h'�ܜ�bϸf����sY�΢�x�D"4�j�_��{k#�V����ӦRS3
Ta��]P�`�0>���n����9����7'�*���G)2�!Kq�������H�� ��u���Ƣ������ߕ��C��_���B�ɐ���Q2ȇ|.|������������x�ΙG��9����5���D��W'LM��plHa��>����f������=	���!u��������w齐�vW%ۖX����%�Yb�P�Sԋ�PF�)hi��0BC��\_���vL$a�2��pv�"��u����=�ۛbؿ����m��`�@y?yo*�>�%"�Y���v#�]����
�i��6v�z���4ϭuj"L���Vf�`��J�ĥ��=�v�}�8g��j62�S��叠��oՈ�����?��e�9g�-a��	�����V&�'�v�Ľ8|J�t����D3���x���ǣ���a�%,�)q,��y3$�~���ڕM��� *�{I��)�����IKe�����N�i��0b��}O��v����,�g��..��a��2����1�x��/�>���mM�2�������z����1$��������葂�
����Sļ���bx� ��X�3��?mzR1�xP���)p�����j�"��t*|<K���<�&��ȚF�&��6cx]lo\��$���
�witi_!���HK�Zd&�]��6�i����9Go$W�����鲂�R�(�{�.n{�Q��zy����a.B�,�kۉ#����7^�^*]XQ��dr	��1��
�?#�y�qpT�׸��;�o8HSO8���v�I����k�(�:�����J��D���6�����g��`S��B>*1���K�d,mD9�}Md$�� �x��Z*N�������y	�>����(O����\��D��ءfq�1�JWZ�i�k���B%���$?D�^���,a�Ƕ�Ϟ��.�崮)��l3C�X�.�3~U�/Y���^���nv�R2�=�%��B��k�&���z�6��H���DԻ��-�uFs�l�׭$�j�Q�OCu��t�f56i��>��u`��d����k�ؠ�5>>�>���>V�6���[z�dE!A
���:ĤIqR���`�j���q�y��1�-Aj��%��V%�ΧS:UKbI'�/�y}oQ��j��b�BPs�C�d�h��P�&��W[�j%�`����_�f�s>K�كdn8�*#6��O���(��h�G{�X�.-U[�c0'�
2{�
>$�dSqw��b�|η��oG�Հ�����m>��o�Zsl֮v���$Y�<�]3	��:P� k�����3pa����˸���Ioyf}-�Y}ډx�E�er������\b��x���6Bć����X`Y����5��Z@�%�_���C�{H��dR+�,R_8�)6������<�Xý�!/"\OlVx0x��@�z��%��,��m��#�Q�!\��E�G���AI3OTf�����,��ō5@,��o0ڡ1�2�cx�k�^>03��F�s���R.��>��P,�톘]���Y]*�*e�FI'�� ����~�	�60O�;�|=��}$Pv����Œ�u��6B��Ma������p�z(Zs�X=���L��v0~���9�,<��Z��ԥ#����9<Y]C�
YW?Tn5Ǧ[��H�ܒ�!`*s3d$���5�ԙ��@v�`���fdk]�ӕ��y���}�mDM��=�zTt؍�/1�Hp�<u"Cf�,E�WlQ?3�����a۞�����6"���I}Hb�ru�t�i�1L�\�&�7���|��^}�6b��������N\��t 9�I3��v��9�d���#v�'�M3��I�>�{��5|NW��Ӗ}���z�!��I!����J��5��?���p���d��]�����!�)-Q�e��b� a������7����k
i� ⾔9�D�(�Nﶟ�e�XJ�t��� x/���oh���ص�/c���Ӏv��	C,k�4r7���{6���c�B���������)EHv�Α�]Y��q��f��07��m
d@�نC��.��X�׫4^����`��L��է�Lq���	�l���o���?����,g�3��1�E���wsť��]�1����cO9B�#~��~������� ��ʩ��%��o#�~܅�VeY�ç��+�a]"�dxNFTv}$���������w�`Y7��^�`^&�ߪi�}��~����G�?vnߨ�U��76��1Ro2sX��Fy���␥+]/�B�L���h�)4cS�}:�uF���ym��$����P�]�Fn}�2!�&���L���R�y�0��L���c�FscuR�b��IP���J����gE��q��;��%�Dɩv�� �������|����xU<pS����j�9Ƶ��I�)�/|P����F��&ۊɈ�ϡ6!��ÛS�(f2@]&%Z����9��:����<vg����c��.��I�wƗ�)�����I�"K�cJ��w�>9����[� v�|P˔+�K��0�_�\�7�|C���1�:;N�.��[@�0W��C:?I��E���J���.X	C����]�&]{war��'6<G䱬��>;�|9g$�Xi�s0`N��R5��՚|V�N��K�;�B����[����ϵ��b#���=Ғאa}pK��#���=�e6
��ye�&�r�|��	/8���=�.���'yFE��YmL��%�R��q�{���{�+D���4�/��P+IL�Q���:i$V�`�eeR��$���=�4�ۢaF��Kb���j��Z����l��q�ws��J�<lR�s�I揽���,��5���$<��Ÿ~���̼J9��w^%�G���3^��#�ܢ$��9I��5�q�P0���xd���jD��ܮ��F��2.4� �5�4�݇��^�!:#A�g�h%��:E��[%a��a"��RJW�<�CKB�0�qX8W�l�Y�����]&O�������S;vY)DJ0�/���	Z�Z��	Q�S1�a,�p;�nFiZaǰ��� ��o`y���� ��b�u�ys�WQY�)����
��qﲶ"��ۧ��m�"�K2|ҋ�h7�O&���J�duD5cY�xxo�Sx���ж��g	��2��hKK���w��]�x���$�*y����(C�ΚcV��Iƨ<��F���@�V�.���J�+����~�"g�B#��DI�1�������Ğ0/�y�sH!|LRxv2��I9y��X(��z��\���?Gi$ƚ��,�������G��?��+iX�ٞ�q�h�gx:��K�߷\�
�V`8\��@u���0�~F��%v���(��ږ;�@�탄�ק5C���+�9Q�q�8��+�}�֐�8Vr}���m.��?�rI�v���5<�6�y�lOT3}� ��Ƈ�m���A���^�!�:�r��2�Q����3R��F:�4�'�'��Ȑ>�z�u�Q�N��Z	d��%��Ү��SY(=�&����9�l8Cl��Vg�X[�I���>ց���ݫl%�a�̒���X��^|���zZ����N�,c؁r�����#+�6�Jnm���kK���}nN���о�@;��p���sT��iO�ւ=yNn�R���x�҄^��>_��(��� ���gumo�6�!5�1�@q�N�d�C�85J��Tr��~Hc
� �G�>�ZҐR�g0���p��s��")"�_R��=�³���a\������4��t2Ieq�t���ު���_}�q�1�UE�1�����=�'��Ht8�>E).���'T`�8@���J�z;�!������,1�0��@.p��-K�WLf	�y|����t~9�Z~��M��]�����c���[��B\D�K��6�n	`��/�܅�Yĸn���0�<saA3Ú'v=�G��u
����]��*����SV�����֩�{���p��˸���?��ch�v%�	��TU�X�k���Y�=�ġb���X��Ú�Q��sHoO��L���2N:��j%��}&�����I�]|�y��'���?{4��C���&w��s��鰎�sc�(� �`u�>J����U�ҥ������F�F|I'
�P�9D�)��_�,��޾5�.�d�uR�YW�z�X��k�%�������M܈(�,ۺ2�G��>��2¬�a]�G��2��&;fV�8|��\A�q8Qj�ݻ��~(���/��'����@U�%�������n�u�)Y����>�C	���oB�D8��eM�#n[f���1ď(=�^����7�-4O����JOV8��V����%�v�d���O�����K��E�7;u^8Ň��S�y�.��O�S$ N<h~�<�����xQo#uT���$��R�x�p}�:[�
���N�.�!�S,VY]{�����Y�#ˋ'	q�;ȁ���D��qX��柆���y�C�]xhd�@�_�*���c�҉��&I��)���Y9n��?~M�[KV��A�s��{�'������zϗ��լY�e��P�%��ژ%ıd�!���uŽ��9
/��TB%�u��v����8���=������g���df�G�y
{<'�BZ�վ{�aux��\�[t��9BQs�$v�1đ�ĉ��%��,j�:���QU}�^�U8�R3�����<�a^`�c`�a�y��g�hv,��RXt�g�7oB�|=�2-F�0��GS�7�v��/����Z�O�+f2Bq�)�Cp��M��a�=�B(�/��j�ܴ�׺P�Z���������	E�j����c�ш��o�oyM���&�l^�/0 ��,=���W�����c@u��`!��"��͟���)Y0��`;$=�Ɓ�5
��i[C�%b��6f0�0D?��Oz�7��T����kU��~d(���k�&OT�S�6� � ե�c�ŶWXauCz�gI���׉93-l<�2����3�x�k�p
�ou׻<zU��uȮ�̶/�Z��0�1�X3��¿�r�R�O]�(%�Q�G�ޟ��b���$~���0T�tP�A��wGm;���w���SG.��ƹd�j+y�\Zz�v�?��?�a^�Ol�=��5��
黰D�eRykDI����M��.�H�>j�w� �z��a3�E���=Hb�0Vؤ΄2D?�i��%h�22���x�s����$x��d({||�x���]~7�3Y�I#����������t<,f\76�K.�ĵ���*���3	^��e���������R�5�`��Q��~~�p�}o ���8�0����C&=�{e͟�>�B��X�#���a.%�b�#�YǇm�u0l�ǵ� ���e�M�ۻ@a�w̃����-�As'�������'	Ct�,:�v�w������/��F��O���w��Z�!�Ѣ!���k0��!uj�Z�R�vM��z�pw{a��I�b+�����~;���P������'e��i��V�F�6�=�|��7X�R�'�qs#ąn�.�6�8�q�1��MA��E-Ä\k�O�T�7k|�Kէ��NF�KC���j;{N�Nc�!;��c�UEߪ셅1����,��,�Mc���?2��G���2<���#-W�K<ؑs�Oe���(�*)�+�	� ��'g4��E��J�5/L#���c�{���E�"s3Ǧ��']E5Q%3�}�,->��lT�Q�Ix�O�'nc�Τ�5����f(�o���#S�'F�*��JX���$)�
���^���X�6�����
��}I0[��9��=�v
���Z��2F�Q�6ju����P��-�N�oW����{�-�A�c �O�t�S��=$p��t%�$܂���?L�F��݆�4mJxaJP��v˰�I�0DNRY��M�{�:��6Ը�K� ���ǀ�`DѠQ��.��U9aI�飸���@^��HԍplB�#G�LCr�k� 4�@9j{=e+�@�b�+M�oE�X�4��T�+��ō���*Th��}��Q��2}�X+�*:�)�mDI��P�%�_�F;ӱ���}�K��P�7{�J[UK9����`��y	' ��������������3um�����Cõ����e�L��{�K%k��%^m%�q.c,
��{�%iH���4��s�]�P~~j����l�R �FV=��  �����;�2�v�w^�1�	��租~REKp34}�g�!��)��c��!0����i���=�C����U[���x��\5�@�Z>G����ڿIc֙�Q��Cȓ��K̽�9�m��D7�!�(��g6[�B��$�l��WBD����e2��_T�b����>hX�f�អ����#�q�xF"3n�{����Z`�7��<�]庁�] /�~�R�����?D�s����D�H�d)97�<�@��v�.��*���ό�p8���OC�l碄g��F�����B�YPK�y�Y������k��Q&��lBMz��!��8]�mX�|�����d��CeCIOѢ�L�"��,
믩sm��V%�l�!ʥx��On�'-ђ�5�l��0��V�ħ
�E��Z�[4�.�?�ssFN��6���t���հ7�8�į��}Z0V�J-p����>���gM���$�O曣`AY2`�
a+�\CK�Ǡ�z���Ln�0�
�?e���/qx\�,��s���-�)<§�6�;&�Jf��!�Ӑv�Aݲ�?�ޏl���S�>FI)QR��>�z���������t}���}|b)���
W�t�WB��:�0,s�w�5�6�3�.I�_���J^��y��n���$0�,�UA�O^�"����7�}���N!��"�i9�p�irI�|EO��0��d���a�GK-"3G����� ���v:�M	9G�O_�B�#�o/s҇�pq��4W"��zL��Ԯ1s&�������&3�Dy��G%5D�+��*����Z!5���(&��ó�I��Z���;�0'�fO¸�q��A��w?�[U<��pV�T�#��'�L�j��¯�
Lcz(�ɉ�� �:���$Dr��Ё��3V�sa�����%��T������@/�fy��c��ܰ5�x���r
5�'��St�<� �t^t�||b���<���X������䰆 ����1Z�I\wɝAu#JH�܌��44"Ӭ��!�����w��γ{�wN���!��=�w	��a�tHKu�8�NO���9���E�e� d����cp;�[7�&.ġ'�AU��7�A~�"�yZҘ�!�ü:zN��C�8�]���X���;$�v��8с�?�݇S��kܟ�	�7�I���P�f�����(��((0>�a�k�k�]�����1qыү(S�F��{hNUz��C��X7����qb�1��9�^K��[5������3����#�-�m�X�s}^+
��qm�mT}�Hd֎u=\x�R�Suc�
�q1VV�k"�V"��g��ז�?��9ѩ0���d����7,.Nf�T��
����h,��^I�>H{��^�٫'٪8y�g����Y�
I'�l�:�u��<�x�pY�3�Q�?k� ��6'��7F\�L�Y^({�r�v�>nV�t�3#���
��VŦ	�*��ƅ��*YfW�0q��{d�
4u���F���TK	sE������tʺh%��c,%��t����fh>���}5�����üϾ��-�rp�}�n!4�z��LkV.ל�%
G��u��za�<:c�8�%��5�������9���r<"A��l։�b����s+J[M	�t�+iT��m2�\y�}-:!�3�,K4��C�i,$d���eaO�1�	��!�Z�U�"����x?�	�g�q��1��.f���]����H3@��k�p����L�I�J�W2�gz��t�
�퍖���&�Jz��^����O.�BHm�{h�#U(`umf��t����.��,1^4SS��!��c>[2�����H�X�Ș��Ϋ��W���=��*�ӻxۭJ�<����D`a��=S�ݵ2��6Y�m��a��J��ҷ����R�Qj��ł��VVhD�A�+Iկ1��e��.�l�I2���K���x}�v�{��k^Y�m>\�#�C)��<	F�F���Bn�1c�,�N���E+�I�$�W��Uo�#f��$��w�'~D���I�:��^��E�H"��E-?���{�z�H;�mN��z��[�Dey�fP����t��1i<��x��k/�9��G /�e���n��,p�==Ȼ�o��k�j����cDe��jRY��Կ��_�p��
	1�\R<�<�W98���i��ڝ�n��̕\.�	���M��;镆�6�Ø)�tLQhu���ɦ���1�W�����[������4�!CƓ�	�����,j�a�A]zs�4��@[��E�B�����F@<m�l^hP��xd?�W�j�ҫt��}�j޵p�|j'}�0�A�Ϙ�y�0_��������=�uۃ�x�6�'��sx����ī��`����4���� tPȃR�i��YJ-�5m�_;qE��$���ڠ�^'��{X�7kt@�I��S���8�2�E�CO#�J�ٙfv�l�1���0�sxS]gOt��mm�3{��DSf���>�u�GY㲖L\�hԎ< Q��ǒڦ>��BU�a���cw ���qx<��C&�����F>"�%�����0�����>4��0�i���������h�=6�]�t&Q�(%�p4�z�w\�r�g�������H�u"��OAӺ/��}��<����`�T���`B����G���In4�F-ib�����S@H�
r$j�ЙB��1��6�^+�e��a���ц�1�W?���1�DYf�׶�=�к.�P��L$�c_d��;t2��<�����v�-����q������x΁u�"a`�K<t]�{���]����*��G74^P�[5-�d�*L�ז�;Wq1�圸�At�~U�	���BBor���m:���'��K�dH�Q�xv},�9k��Q�v���+�X���UX��6`_��H����7w�=灰DM�#�W�j�!��ջ��?
^�3�c�z�oc�����j��3æ��u����c�]�K�{S��,��ac�J^�0V�
�hbUVR7��X/N
9����Q�h�w��aw�CF�g��ֺs�-��O��iI��Y�͹g�Ɋ���t�@�-}�+���j�� �A����lX����5R�s����]&��HVK��i<�{z����!��#i������ 7�x�cj��� ���2!0SU�P��3,_hXݳ��*:���Z;?0�"Xa
�B�g�nYq��mei�P4���Aa2 �M��pE�*V���>C�0�d�슉C��u���1&�ba�j��=��tE�a�� �{.V3�Tl��L�nk%d|#��Ơ�^%��r�L�Hx"Ad愠��2���q�=�4��E�0V�n�׸"1#]��e��`o�5mp&j��m@i֜�cH�Z�yQƾ�Nڹ;CP�lԆ���t��o8+���֐�)�D���'*V�(�Duޅ#R�+��:s�>6:�}��Jvy���<�[c{L�6K�{w"���`��z�}zo��?�ۭ��5t&� �]���^R�RG�����3���N�.�>����*Ʉx�!!�>Q� �"��|���Ԭ��ظx��4�G��&z�~gL���'�%5{op�UM�N��uZ�6q>���9���`��W��]���u�R���<������rKj{���B)�(���Զ$�7�g�&���.�_O&�?X^S���9#Q�}���Zoץ����QJz�]��2�5Y`~.=>�	$Ew�D�����cH?W�cSH����r�yS�U�C��d�Gh|c�<QWr!�B�+
8�X�
���)����ީ�t�]�;������2^�����W�^r�]� �ld����R>�m��n��v��������Km-�sqCps��YK�Hm^��1�وWY����:��~8}��?,�p�vS9d1K#����e��q�^����BK�6����DG�&<��MAK|1BjT�Z��k�.Y�VnK;z�8��;���*���r>?~ʜ�x��=�NQ�r��Z�)n�)�L���Y:`��y���`�3�h���s�uu�W@�ځ+K���2�lL��v��:So\��5�t�ך5�i[y�Gzݣ�m��ӹ?��`9���F�E?��8��3���z01Ԥ�Jh[��ۆ�N��A��I咧���%0$	���ԗ�{	�����~CR.�r�U��jYZ4�pc�l�8-a���l�ݺ$�d�6��$�ӑ�l/O��	�W�;�\/_��^Ay���%,��
!Ђ1�f�|WW�&{���K$È��c�*Ԧ| ��i�*c{�bo(<&Z�����v��n�`�LCY*=jH:��U�>O�I�3�p �������k��Y��mwA�P�m���;\��CrNbC�֐�}3�QaS���5 %W��h���@�����$v�Cqa�UU\�gnťH��=��z�"������41�,��	��@6マ�t!�к��À��}B�7��|(g�TӇ�Pey����bB�^�~�_?#�-�l���s�����<�!����U	!����
I�W����2r�w#W�V��z]�
��_���~ICtg�����7�E(L��wo��l�hlk���O%��$����C�}r��_LEA�U��C�D���\b�ج��d�o������~��O� �!#���V�I�X��k��C��"�\*���?�Vx3+��Okx�%�4��9�� �PP����f���Ik[d��}~^�d֎F��]&~���A���R8���t���f��q�<x��Yyq'��T�^�k�����=��8�a O5�M����q[g7�����]_�2Cޅ�R�{��x]��m:
h�|'y��.��e��|�����C��P�1v|��%�f��^�SߥPP��&��b�쬄���v[���*��#�:�7g�4)26C�nkf������{ᰬM	ys�`ɠ#�:���v�J�Qc?��\�m�v�f���d*�Ms��7�����z�������_;$��P�l K]�f T�M{V9�)�D�}�d4hG��w��~����̶���Px����Ր�Cu`�����ET!1��Nl�n���#.x_8 �O��m~�fL��l�S��?�")y�k.(q��������5=������m���qϐ�`?��%k�UB�*
U�&����$��D<_��4eB}_Ss�Ԇ'єzZ��8�D;hh�kdPZv��nܚ���(��M��$��ɭ��8����!	'CZf�Z�4%\���=Q����p4eK��� JOOe�~7$������u�[YE��{�<nƒun�3� x6+��C��@���9��9&�n�!`H���iL(/m�tڜx�����s����Oi��v36Z��bW���޾|��Wعs�30*�
���ژ�� %���A�"=i$[��-��YF(|`�>>\��,��׫�}����}��c�t�����\�X?=sVۖ�w�B��"؍V�
|��!��S���1��N��d����ڤ�����vaC����jn�Qx�_s�kF�3;��?�2�5��Ꭵ�#�w��Șdy�~F���q�33p��L�Ȣ	.��&oF~'.;v>'N�v��4U,L�6DdG7�ӓ�'w�C`�ڗ�RЧ��䅒-kV�H�t����	����¢϶a6�2�5Hֵ���cc�Xx,w�X��C�����l�q�<7o�yP�.i4�`��rF���y���kQ����M����(�mM��(WE���/K�Q�G*Y��f�|c� 4�۾�6<����C�6��q�7��-8h�߾����Ǉ{�ԕ}v[^�|V�������QZ���G�����0��ț��'��ֆ�V���ё��*5�����/�S���Ǐh�������O۵QUڲ#�͈�#�Ð���<R55���Q���,�r���L�h�]��<��=�$��n׾���N���{�<ExCx���i�!�CLC�dֺy�=U������$I�b�̌.]��y���,�C�G�I؎�S����W�%U�P�]I-Vm���[Ѯ��>������Ë"�wI�0r��7McM����?0��V�������V�z�7\�_�4�WV��]��O�
h�2AG1�ݒ����%��H��ϖ�Rkla��/�
=X>�޾s�V��x�x�떍�bJu�,;}�:�%��Lc)�����$�E���LZ��XI����jf��'vt!]_������3a?�p���c=� .v �ɫ��B�W"��s���]�����:��8�Y��$J��YR���$������w�p��!�1Re�W6��w&/w�o�B��8?�_�ܞ���_ыe�9��`gHV��w��Q��ܨQ��P�T�gw���YTm�b�^j����	KE�.BZ���3,URt.�%7����[9�g���@��ah}�񐸭�z�����:R��k-� k�(�=q�����L����~:J�H	cS"��1��1C�����Ո6��]��\������Ⴞ2I�H��!�x�VE�����#���m���ui�j�s���g���x�`���Da`�����t�K�l����ߘ_U58���	�xZ��)]d���47�1g�d`;mߠ=M�ū|;�ָJ�k�ey���ܯ��`��KL��jt���t*��Z��"�Դ��<~�V�08x#G�?��f۠��a�������~��W�s��j1[{Y�N]a�@��M��:��Vf�a�u*�|̆m-��MRrQx��9�P��vy� ��Ð���w+<�5�,����y�.tZ����)��<��� �m�σ��%?|(�͈�e�u_�e����>1�_l�ź���u�a�
l����K��fK
�������B����ݭ:hx��>��P��a�ޖ}�)�w
��]�V�NC��0ڨ�W���~Z�zD��.��<EDW\�;�7D���!y����d�j.	��Q,`�1�B��m��F�՘&�����ϠV��ަ�>��{���=�b��0p|a�1	��y�V���ۡ8ӋUe�%D���������?K��v��/��jd���Gʯ���7�+�����C���\����wR4�Y�*0`W��Bw#e}u�����x�I�I��FU�ifЇ��/���c�0���|�&v�<���"c#|��������<�c3���2�m��:A�2��m.��+.�'��*���y�MN�B޳�MtX|b��������D���+gI�A�����VϥU�u�P����D���I�q�D�VY_N:��gx�bF�K���NzK���fr��Y����!�pϐ��a۸_~�U����JzT�8*�|�����^����>]���=����<��N!���,_m��:�xBQ��9:��$.�#ؐ�`�H�h���z�����q%�lxN�� x���ޤǆ�o���=�S�e;����,}4�� �������?�R�V��Z%�[o���n?6%.��:�)�HoRe��h%��k�B��*C*�^�=%����g)T��w`�@��ի�������.#پ7�`��]���~f[�Q_��V����Q�?1��Ɔ�CZ7���:�� �[��5�ChNeJ�B�H-]e>�Z���1�B�m���u� �q�Z���	��ZE(��>��,Թ��Y5�k@2�0nh6�������n`Ha�ݠ�3��P���o�����v��!�َ��<�1�'I#��`����>H�Jmƥ����(�%��p��υ��C�2�9��`��6ـ*"� �j,�n⾸��J����.�zI��ң-�Llv��/�������2��#���*���5������s����_��C���������
����q�L��_��(S��,�:�����=ҋ�}�/^��������?ŵ�܊���ٳ8�#2��ݻ$޳|v�^Ԙ���[���a��1e",(D��*�ּz��?co��q$FfV�t7I��fg����}����I"�7�:��473�(��TT	h�P������9>{���~��r@�Tΰ�'��]��웈�:^�7���B�����;P߰��3�!am���K���f�l������{�߃�̲ҧ��ǈ��s�+ƞ1�#
V�{���Y�a6�{GG��,}�% �(P��,��q8�߳��7z��^�w�ڻ�[]�)��(���s����E����۝��]bb�]V'E���\�6��#T�i��Is"1w������+R��H�+���a��Q�O�H����O?�(�����}_;�fF����L�Er5��]�/�F9���g�_�V�4��g��=9ApaGE\׷�����%�����d�`ɋ+��6�K#%�=�ɕ��%�uH�f,l�s1��l�;W�md[؋C�m̑Y��Z��4�_�� �?����K�2�!�|������0�2��gR�>F+�V�������D��zۈx?x�NJa��i��b$�������p��?|����횎L��'���=� ���5)~�e3�WC�Y������5�+�5X	�Ԏ�U���׮���U�9G�l@ a(�Ȏ-�٪�Q]a�c�0��Ӷ���#7��^�`�QQ�5��	���j�b>�(�"0勞lh���V�p$�K�} �X��!s�]iݎ9���ꝲ�ik+��N�����/��4�i2'-�u�摶ofC갳��2����YVd�#�pu]�ϔ�h����>�g������B2�ť_�P���$���4��6�:�`�1!*����@4GL�8�R$K��NȾ�0`�K��X#�:.�G($A0<�sdP?�
>�X����
p7E�t:����D�c�c
_���:P�����I,by�)}7L7�׬F�v�8N'yħT���}Q����t7�AQ�t��ԣ�I��J�ge��MNm��P	���
�? y�M��s��>G8��CM?	���əY��К,����߻�xL)��M�y�h�)��! D�^��.ƚj�L6�JyT��!�^#�ެ;��=b�~1ָW<L�k5f�ی�]py/gbӅ����]�Y��(�1����%�(�0�C���W/q��o�8�4��+[���#�_�@���NIOt�s*����Ÿ�ÁѨ�MCr�t����:E�S8n7����4���~e�~I{�e����W�}{��J[�wԟ���y1xm�"%��e�q&�0`��j3�]sq>9jQWL9�ލ:�X@��)��V!���>2����2aR�#}���������O����y+�X���i[�0���q���+,J��Y���ҕ5Ðv!x{��S|>��+gb1��2xćX008�a�z0v�ې�c�E#��H�����';�fѱ�!��G�I7��o�zN��2DU���,o������R�Q��Y_�"�))U�v��'�������x�?��>Z��!\fa�'�M��#x�3�=��9���$��G�Y�������F港�R�$��Hw:l:U��H��=RWŽ���jZ������H.UڰK~����!�ǔr>֨��юǽ!������sQ�U�߈lP�W_��BΘ+F#�J���-�|?��z������sxPdUY&j�N]�C�{~PKq��w1v\K��1BĴ`F�E-�Tw/s(o�ƴ�m��u��qH�M�>q���:�L!E	�ǆN�o��l�j� ��.���]$. �gYL}PP����� x �D���tL�m��u�X�z���-ۥ'C���vǘ$`F�@�4!Ģ��!Dq��/q�D�Yv�Y^9*�]�l��q���y@�R�^�8��;����`���e��c�n}$+^^N�5�$/�v�~@�i/l�ka��p
	�$E��p���B�	�.��y_��*�p(j9ž�0�vo/�UyQ�x����M<ewem�*��Rw]V��a{`gؐ����1������e��nG����;uJ�w�	�b:�R�%���Fu����1i=6�*XG{E��kz����I���N�#�z
�C��&� s&+_�$��I.�+��b�`��I�Y4/�=-��7�h�AR~&�7��7J#�h���VBA�dS���4�NV��� u��޲��:�E�YM�$Hzg ����ImR��ldY����2*���"��dΪLԽd�1O�bü@'4Z#����7�,�7������:��&�K�}y��6�����Nde���D��܉q�(�9
��>/B�Yc;�-a�c���(�����[B��B�Hn��3k�q�/��-kme͖�l����]y�V�b���[�����g����d�/�����J���ڮg�a�>��E٥��P�R�[�O0,�|�@(ĭ��0�����Qq�&E*0ե��Z�c�J&����ފ�6��//'2ҋ���]���ʨ
G3�r��}�\�xUr�M�e�9Z�.�g��T���e`H�糄V��;#&8fXLn5��CVEb�M�7�j�J�"ӘY~$5��u��,(M�����0��o��o���£��`������-J<�mªr����x8$�g e]n����K�Wj����-xbJ�,}�ྑH���P�Β��=�N̒�.�g��Y��2_㞿4����'=;�kIX /���J�	Q�4�i�]�h����|Wa`I���S�"���>\��w�����@���M9�	u�˧U�����80K��D���hNG�H�w�����q���1�["L2���$V�q
�{z�*+1iD���~E.ݗ�����X,%w���I0�O�6��%��/��B.$UT���-%�`D����$P��f������%�~�XK��g?tpf���Fq���;���/c<.���.�R���#4�!f�M�6��������0>V=�5��c�wC�	�kQ���8�[m��ۑ���t2�
q��ؕ�_S"��wd�EP��4�pquT��<�s�]!����!�W��z�71�RZC ���*��k�j��(���|���t�)i=��x3��d����5GF�1�6��%8��~���p�z� >I�kʪ�h^:8���P�6���a��P��T�Ev&2��������n�ID��ꃼT�5�6�6��rIWu����Hm��kT'%���������׶�L�nMյ_��f�a�B���n�����X`/�7{����&'��G��%�媖�+%�T,g�Ӎ����n�k���֒H��H�t���CQQ3n�2�p�I��"Ga�,<�)��1<R&S��O���a����&p���/ݮ���FZ�}�	�؛�F%/�m♗�-���Ң2@4�Ʌ�7d@�jQ�6l;$%s���Hx��0���T��^��U"�ӵZ��� ��vip��y��
O�<�亳?�f��\�X��]�Gb���E!�0�b{��׷���"���4�b'g�We��]��:���6?�oh2���X�Y�{!c!Zq���4�M扞�������՗L6/sM*g(�ђz0�8���"�j���Zp�^)��(���Y��zN����	��I�[���*; 0�טA�S}~��לc��|�{�gOr5����k�R�GҚ���ԕ��5'���Y��=7�Q�T����rRVSt���v �wE`v%��9��,[mt�̠���F���AE��@�QTT%�(OnH!�S��,kz��ĭ&yaK-a����"h����U�E�L�����^C�|�����wa�������Xy+��"C�T�a��)k��9���}�� b�����)��q�{5ɢ3���ܜI�bxgv[	:��I���;	�����o~�5ᳱ��P¼�$N�Ćղ�7�~AȞ#�Ì?���|�F)����`I�{�|O�T���ͥ�.9
8���ciY�,u/��k��5��n����-��r����0�8��#�Xr�j�:��b�5Ǝs�&����9y�~RM�,�H�c�8��ry�{y#�fq�|[~�`�Ũˌ9����_#R����/�H�sV�,��6pǵb= �2�۽���� ��;сx*n����� cK臒��G%\�,4�k&�m�ر��7���T%[~�mb������lP�+�|�� ����J�㼈��b�h��]�OC��BL�
-n\�FZV�%Ɛe�ͩC<�a�CCaHA㘩�c"s�:?>H�O��P�.V)km���۝|WM@8䞍�5�j����odn��𧠺 �YCteR�]�Э�C�S"��#{�!u8�E���]����aXq�.5�[��4�]z��/w���s���1�$��րDv4<�;�2#���°�-���܌ij9�('}Ì��-��[����S�� C\1�-5P�lM����2�Ɖ� ��p���N<�z[,����Klb$�X�t
.��l�����`������:��u�K��rz��a���t� ����S���b���];p0CN'e��Kzڟ�B&�0�DV�&1��w�#0�H8a�`�p����)�ۏM)%M���g�*�=�����*�ދU��}�[��馤V�6�F�E�W� �7�m�#JC��!�6�<�i/�%�)��a��{�5�B&br�Ւ.-�����kc}�n��)�,��*�G�S���-���dp�3�P���Ъ�<��P���{3Y����"&�r=�a;�Cf0$a�M�cM�*�-�xH�4y�ܐɩ�^�{A��4l��a'�)l�����_���>�0��Ҟ!�}����<Ix���J���3Ԯt�G��s�jQ��u�T'ϐ�u�s���W��{���hM��5��7u�WI&�'{�q����;)4�-������0\�\
Q�� =�ș]#S_ˁ/�4�C�v<��,��M������p�G��\�kNTfg�N��(��(wz	x�����:L੝�"���E��8�	��#���?
��A�ͺ?�#���}�� �@� �5��4�>��A[{<�#)�h�6"*E�0�x����?EH�z������n��-��fd�u�����dl��Uv�+Φ��Y�{���Р���E��P���Эq�� ~���f�V����-ڮ���e��$���:�\��H��g}�a������I�1wT���(��|3#�V�(9����z+mm��=@bUL��17�[~��7n``	�U��.km�S���T\��&��T�=��޹K%�j9���~����JS�z���!�Uh{S�� ��\ƝD����I�Հ�4b+3��=�IS�E	?��h�b��o|NNo�Ezv7 ]F
��!��x��G�H��Ø�yIl�=vjoq˨� h=wT�a���Ab����~���M`^X@q�}�w�|*+�T��MlN��`��s*lB�37$��`S��&z kA^����G	����˜�x�T��iQS�H����JH&/�+EE�?Zh��;߈��v��,���o�w��>�O���)�?| ��|I�����w�s�<O5I���X��I$'sW�;6;�u����e��9�a ��=j�`�XD�kE�]���W9>-NZ�+��4i&� 2fX�ޅ�k5���Az��v��t�QhM�|<��;���}�^3�gq�!����Ƴ2��b�f�ݣ)W�� ���̧̒��paޔ��R�jl�������$=�Z���ͤ�MJX)�'�����'6(K/Q"������*����f  �WB�����З`8���9�ZO�?�han` �E�!Ø|���lw�m����~g:����˛����`1����QɵP%Z��1����#ta�g��*�{���b
D�&������C���P���<`�B�k
ܠ��Y���#w }����k�S2��A#���X5?�c����a(B���O���ew���"o�����#�����(�9��hk�o�&�+w;��Hu0��c/���k M>7*���������������Cw2�NSڮ�w
�i�Ae{�H+���UѮW7qH	���vm��I��&�ZZ����#v�kV�"�w ���|�yOyj��ΗKPW��#�1�W�ʐ
#5UTz�꯭N�V��B�4Z"s�DJ~x��z��Xn�aR��@%Pv(1�](�@n����O65SM��*6�T'���rN�r��
x�-ԉb��,N���\�
�9���\P��ק/Q�!�h!�D{wW�+6ڶ���������N�N�z��E�:V�X�vM��B�-<�K�
P�`n��S7��L�'��m�Yj�Ȩ$ͨ��I��0�0
n<X��C�����(�T:�/�z&��훸w$��w�OOa`�6����!�Q8�,1z>�~Kա܀:���G�c��j{S0H,Y�����Ps� J?~�nC������}�h\�蹗;2�K�dG5��,}�_m�ʐ�i��n�C�Q>z�>� 0<(��ケ�������������fB4�ߔ������h��D��]��*E\��ą���+pB�0+�ُ�V�yRe�޶��M/\�}����A5iͣ��8[o��&��=�Ѵ��x��k���~c���b�t_}C�:;�����j��	���$�"æ�̰z~��X��`�v4.���J�:���y�;v�a�i�/V�
�`��Hè��,b+�9��\5���v�P&:DZ���S\UxG�㟢~z����&���{z��=�lc�F�=�=�D4 `���?n!��X��9ل�yM�PI�6�SD䇁B(�(L�^Z/c6KH�X#d���Q�V�t4������䦦oJz�˚!�H�1��o��TB;��a��À8h�����g�(��M1�`:���L�������S�͔��#�dF��DYl�mgk���L�oL�{�#������r<�4'�"�1�m�ktx,�9��I���4 �b�6�LH]�#�ヮc;�q}(�E���	����X^�ϗ������������ט7JlBbW�#��.Tۆ�%t�v1���X>�s?Pkk�c���	�r���w_��i=��m��������ޒ^gM0�J�S;��ǵ���Ȗ���LAkMK�\������%b	^�H(����?�J�ۼ�������������!H�Wf�k	����H��]�t+q
����V)�O8�m�^���XlP䁌¢(!ݮT'��Zx�%qXj ད�L�v=����������˗����5�*����EaA��L�y�SOq��
7_�I�q(���E����lX��Sx��C���%�����:HB��L}���캤*M���6��۸-oi������_���?��Oq��!0�sA�	O�ġB�<�����_�k���a=Z:o����D��Uh]U��7:	��px`����ت{��l3z�6�{��p�ᷳ�0���Ѳ��Qz�>,���ӟ���kzbu�_��桥�W*ck1���3ߛ�a��p��QūX��y�|Yc��#��������)
�7�J���-��{���N��D3?�I;\~p<�w؇����^�P����I-��/���RigQ�AO8ztO�����ř�������=43�Oc]���>�����&#�ũlٻImj^F�Y�ɀ�u�� wmYS�:�E�$77Jwu��L����d��V���c$�2H�b��_�*][�>ܝT�z:��F��^��pJ��7���F�R�SfI)6QrX�JEull�*&�ӧ�[��a3����&�A}mhH�ğ*�j�X�����,LL=�b��d��@b�=
�õ^B-�`�O������5��j�=΃��df<�67Gxx�kcEۍe��1��PI���|�xT]�zg�8��z ~���aH!�����a���H��	��2;��ڸy݄�X�ġDCJX��3��{Jhڞ?�C�=PU!����;te6�+� �x^����9�Ž��4�he�׿�5�Ƹ_J��Q5�D-��Du��H���ʻfS3��44�9�ۯhF1"�h����y��Or^���bMR�Io��ivg�Y�s62�)DιO��ƹ�|/˗�w�7�.R��U}L�A�?��XF��PT©��^�z�a��f����F�	���۲�Δ�%�m6��E�ȩ�!<��Q��E��ܲi��ȉ$r�/1H�=�3�Ђ9���t��v�m��[PP�%8`�����mH��{��B�k�߮o%�vH�Td5�0ٞظ�$P��D��|mH��P��@�ݻ?���������O����#�*�4��	�)D�jJ�-��7�R,�����?'���~/C�-C�҇q��|x�1���X
�b��1��?΃�*ċa$�{<��J�9�B��n�dx���[��s-a�xl�58łb�#�X���D�&�3�p��u�=��_�e$�c��G,E-Gܶ�t9x�_`D�>�p����ݔ*�!+x�A��i$$f*���9`,����Fi��(�(�Q-�%�	����B����N�!�"Nl�G��u��Z�F������k�G������-.JF@�ݏ��ZK�=�*�\��:|S��e̤%bM�0��H�U���6���R|� ����k>,���<���e��T��g�8w���e�jn�:��<�ր6����u��_U�����K���d����E�j���z�'��ߌ����s��:y`)�ܳ#ט��J�g���N.�rw¤�
�CҔp��q�ԋ8���{��Dۀ^��B�t�Z������;���-���v{�k� Y�-ŵ������q�jX�@#J���/� ��pK���rg	y�kx2T!��-u�_�x���>�t9���.]��`��fYj����IB��O��;�z)���o��@���YcxyC �]352��{���u:%7�H�!��Ir|m�Y�����7�4v#���|�A�C`˘'7p����7SSg�K��O�t/R�Bb��������� �P�kj�D��b�/��\�v���*L�y��+���6���}��UHY��y� ��\A-�,���悮)�n�LJ/58*�a�Z)��
A�ߵ�����Y�ƈ���M�6I�(��IJYBo�����|=w�pg'S���Yi�O����K�Xq�8���˼ġ6P�>�{bb� ��^�	���`�L�v��w�қ�o����R��S��~��!��cp��l+�\4֏Qq���m����h���zZX ecӘ�����I�	8��0��5W��hA�m�',�%��������������I�0N�P����k�wެ�5��!�e��UA�T�ҎMo �"=�1�j� ��N��$���HÆ3<7�
���W�d|��n�X�4;a�����$����&��)#�^o�#�F&�޳G
�8���e��b��B
���d3¨ņg�=|�MmN��J�c��������o^=��y�W����q8Q�e�{�a����-�5�w�tf�ۏ?�J�҉�8;�0&؆H4�:	�����WX�k	�����db�%�Л��C�n�L\�@d���S���|��Z���j��^0ڣ�I@g�����a��:/q4.�d]�j]�����>���|����12vK�h����,�|��+y���^S�h���'e����0wo	�u�B�[�n�fu1}�U7�S�%�v����m�0�A�]�����h&�y�ġ�I��~����m8���́41a��#i��Kdv8T|z�Mj�ς�����D������q'���`l�3�oC��]�3Q��v]�̆TViq
x��=�20��Ы���H� ��п���5����5	� ��w�ƁЊ�`Ȣ��2�a,7C�v�^��r#�ʐ>=똡646?<D�N�3t (���yV)�˹�;�(�k�i~��=�<�O�_��J��)q�g}���cs���P�)��A0ScرM���Y�\����I�7^c�n�(�D/
���M��{R�\�����)"iɲ�s�4=�Z�%�L
�ĺ
���E�t;�
i��n��S�sF�@W#�d0"�5�\K:;p0p-L�����ihP7M��S���8�x�����>���B�p�9�`�
IW�	&�9�=�$^Ӄ.�����B���Y�I��4Ȯ���b_'�k�ii�����f�������i\_�H�_|_�u��{�]q=y�$�
��F�̜�^v�v���X�Z�pE�qB�rb�P2�
�e�+�P�xy![�&����~�s�h$."[�*���f��y���?��B�m��bivYed�$~'���X�?B�0�d	 �{��L�n3�X��((!e��>��B�
/���9�uӓ;8�J<�V�k�g^ۅ���3<�)�N�dƈ�*��ł�̡��O'�Iz�k�N �e���"�þT���}�����O�В���"����AqM�M��m�}��B���h��a�	���� �6a���vzHZ^s�P)��S�`��7��!��퉯0�g��A&���cC���q �v�������d��^�6��Ř1^L,.J����懶�3�x���Y����{�μ��A�{�Aq~��6�r���L�iNN�e�J'MgteU����%?'�1��e0�-�(�Z[�{��p�%��������]W�+�V~D�L��wu���˴�iD��O�T��o�T;����Ѳ_s�-��dj��n���M�f�6keG�N�D��o7������1�Oj���.�+VQ���![� <F�F�j� Y�Y�L�/}$
�������&�h1��]���s�Q��b�IH�⾭D �j��o�ah�nބ�3�F��wؾ?l_/{������<�q���C,�;póp�$9[8{J���y�:�%hf���
�|A�Fk ��{��fab����/5"�X�x�n�\�U�&d��;j�Ѻ��ց��Y�k�HP|a�-��篟Ch�k`׷䃚k���snLd�*q,Y�vQo0"x/�0�0b�����
�M���X�o�$����0S��\H�m^����/f�5�N;�.G�l�hٌ��`���c9������z�[���h�Z*#g;L
 68���pjӉέ:u6�$�7�M�2Y��QUێ�6>U�S{NC�ίA�ݏ�-��Hܪh;���C%�Os�p����]�Y>L!;��g]g�җ;h`W^ҊE�η;���p�u�������J�
{)�k���Cd��L��(�c���k���Ϻdb��nj[{��^��Y�N�aa|��>2�l-��N����u�+��z��Q_�x-�欮��E��ɨ({�*�ݥ��HG%Ix`\s�Gk�b�{�=��s!Ro�ޤ�R?8�&Qc�o\tOq(�f[��I23ܟ��^�>�{�U���,t��\S�R[|�;�+�j����p��3o~���&0f^�����#�9z��U�$�Bu3(^��:�t�S�a�@��{�S����zM;��dX�YG+�Q���)\��s	#��˩��0h��C�8=�RC�+�U�Qq8�������	#�P�|odn�j�5)1�`���Xv��)<����xS�ҔE 0潔�Kw��������\��믌$/ّ��H@'�IG��E��K}\OW=R�ש��/�JjĖ5�O�*�d	E'ɛb������$�	����o=Rf���ҹ��N�T�G��JE�Fsf8�!����3ae�Gʒ�蕔��U"�0h3�S��h�-7�U�!N��W����}-����p(#���%�A�m�GƆgi��m3>��(�̉�B/?{ܐ�\,D\�w���a,������/�q�SrSN�H�c���(qoT�	\p�̥�';aֵٞ)b���+������)�ŚI�B�Mp;��,�[���82��*���F�f��p�pHQ�BUubџ?}�>D4�%��3�dx9�!u�H��}u��ݮ���k�g��-�7;$�T�����8*4�ݐ��=$��=���R�u �h6D��B���ꖬ��m�݈Ra���8̖�	�wT�r����GB5h�ѓ[�'��5�#a�c����b��M�JO�G�_��vۚ�*g����o$�MO7=��i_,#�ݢ�*8��<��M8K�>Q�А�2�� A�5c�l7��&2���J�V��I8�OG�k�.�[j�Z2U���j�>�v
q��kM���I5�1�ᥭ)v���8h����D�Ԕo,W!��/���1+E��׀G�+zq,�����Q}�v�����|�U��uc�$Ai���L2�� o�C�򮾯��B����[y�EgU҈�h~�����OM��$�^a:���k{n4��9��z/�v��M�:dw�|Vg�}�:Z�ؤ6�+��:��v��-��=��5��M��ϙ\��5�y����c���Ϝ��V���T�n'&2ݓ��2�t���}�bzH��>!�eC<V��^�ưԱ׆$��Uf\W���ι�Y1�a^q�BWQyz�[V-���L( b`Ik�F�	x��vE��y�=8�D\�X?1���2OR��ʒW��Ki�@[ϒ�]�vơ�9�I�����e[xS�\{�=�2Jͯ�J��[���msO�����y��>��>*���MM�!>>����j�x��(�8�K�,�2����J���>P�xk]�7�u C�l�(���֪��x 9�k�D���(�f'�|���L��*^&��2����q䱭Jp��pC�ә�X8��7fNy\�XݔĳQ�gu���^a�9�{�Ck�^��f��<Kc�<I���6�r'mWc9���Zۤ8�]db�������&|��!�R����M�k߉�ʓ����74F�DI!N��ajV�d;+X��GC��{�S?n���
Y��X8C�&qZZ��K����`t�_&;G%a�I^$�㹧G:�Tq_Ŀ����=������cHF:R��׾���)�Ö���q�)�o�A*Mq�l{��Z,zF
$I���*i����S$����JϾ�c�����;�a�#�{�3�C&5���א@t�eb�,��Co���R��E{is`�j���e�~M��>2S_��|���Y�]��un	 u��)1�7%�m�N�O����*�lF( 	8
ps{q ���Tg���1x�I�a�@6������B<��;�|p�ZE4fƿ��.J\��S��T<%~~K��4�X$
wbiw����S�Nɫ��ha@㹰/Tv��hn��N/Wz�{�z?�<x6#p~���w$������d6۫��2�뚑D�Yxa��ڧ`�R�r�uS[�P�U&���ˬE'�U���]u�p�wl�֢3��90��tr1色�pMDuؙ:0�K$p�&vC�x|6�<0�s?#S �IH�d��z!6�$x3�ö&$�0p��q$�:`���?�����Zד�5Ԡ=���M�Bl1.��yf���(��a���7[}������w�V�����r��ն�O���]4Fڐb�̓��o��à�����%���I.�������<����{�kb�s�����<��l�i���e�1x�G��a�LcZ]e��"���o�]��:�^T2F,��EaYf�4�>��H�w]#3���o��..��M��� [�̵���p8�� G,ȵ����P�p�Mg��<DSYz��__^;.=�/&����R�zOxYK}J�x�^4��o+�B�k����J|�2�c�"brgm~O%uWXE��[w� Bv��H��5��n)`�y�D[������"���3Y���оq!4ELO!�x����<|{�_{�f��늉�U*-T�#ݪX*`m��A���o�AP�����ǲ-t�gG��%�9�kt�Sݰ�Q�ipA����Ε����X�{B2��j�5��*���{�6���,,���G���4��'��c�ӗ�o�ڎeP� ���C�;ڬ�������a�v%�GT�	�ar�h=�i�{m�''�*!w�oA<&��<�.=wG���C8�~ʱ[h
	�7�1�w6�J���g��kN&[�R��f�~�j˷�}[3���N�Q{|�v ߑYb�z�>� ��Za��4PL&����7�yδM�,�!��N�IwcNT*N���Ɩܰ��Tc���<��&�{_+�G�#D�W�v1�5���Z���/�S1��f�z��x�˚�=���
Q;�w�J���L���k4�QQ
�@�}�o��d ��������	(�*�]��e���ȯ����Z�*a�Z�v��8�ם	��� ��	;��,���uE�39��	�c7��ҊxO�h"��t��*K�q'��q�>�{��E�2����mvr:꺪ɍ0⥲h`�.���pXGL���V����#M�k�N,^���6h�&���l�֢k�5:��k ���;& �Ŕ�x�J���]�kz��!��&v.����t#<�;�ͷ		X���y�9������g��t��F��NX��]-u^��ҙLZ����iQv�&
�$��a͞m1��|�P��'��=~��Z�ۄ�=���u��AV^\ԻfV��k�c��/Sn:׊����c�+<�RuM�yQ�t����ڠ�=���m��4�����X������-$����q(��L,��g����=�R{4r��Pc��wj�G���/��1Q�3��&%|`��*_���Yd��:��N�a�'���b�D��J
Rr�U*�U������y��EF�V�WY�-�e��ΐ.����lb<�B��F��q����6���]8:}2�[��5���k��^M����W�tM�G]g�>aL�>��zLq��5��O'���%qX���D��{|���
����/����v6^������5�19���K,2ƾT��Д�����*5ئ���
A#`�'HQ�_է4֥��{�]����!����?�h����q��=^�א򄭓��k�I�v@õo���%|_�!N�x≁G)�+��{e[ {�5\�ă�R�?�$B�;�u��]��z���������=����T�X}�����̺����>F� fe{�u��#�������f{^L�p,�[�P	�h6&���x�J��{��N��h-�J�5?��^�Պ�!,��'$d�ZvyPZ9��Ƀ͵p�]8��,w�1���I��O���`��yP��q=6�L%�"qٻE���x�'���>��M8�ݍ)54/:���:p��Pv]��6�yPX��n#v]5�;�e���Ν�p����x�u��;k���FĆ�E*�*ʞc_��hbWrAGv
�(�Y+/�Y����ԡ�Ȧ�LX,[��{��"Wt�8�c����p�H�C� X��,������_�����p#D;e� ��f|VN�z�y�A�������i�M,]�^O��7��1n����͝��R����Hj]~,"R=�5k#L�4D5|�wxj�A1��:#ۉ��s'#$]�>x�!R�Vq���d#j��bC�W/i�<��_�t3����_����qa���;y�ʊ��5g1:�x��^^g>E���o�hӌ<G-i]׻��r�K�V��k��=���J�]��]z`�3�L��^�1O	Dy���Ax�`���:%��"��݌�ݦTkzMY��8+u��
싸q.���oӔ�37�q�n���	:WdD	�l���/Un����F������C}|PD<�d"*�*K��hM#y�P3bՕ��(!��Z(��X;�v�e3s<�Q�]
W-���`�/Z�M�u��Y�C��\��M�)s��3�� Q�cѯǍ
V/w����X�7�R���v���4Ѻ��u�����N����o{�2J�$p��eć��bB������Z8&�>����<��R��^����LU8]���,��J��k�C�:yэh�L�]��٢���k��G��BlF�m,��zR��ކ����V�>F%M�x�p�\SݑW�	Wy.�{D%˲�w�����x��=�c��:ݱ �L��UZ���V��o��8 ��/��gQ�,j;rI�� pq[�"�}��d���s�qm�]$���[&@��UOϭ(��:Fu�z�]��w]BH6r��X�p4�A%�s����1�mcFf�	��å5z�W����G�}�@D��������0�K%���>���ޡ�p#:���pPұ֡����n<���c�0P�)�%��xs"�s�C ���LNE{i1jܘ�纬�3��'	�D��f)ECb/7���)�ɪ������������6�ڊv�x����Ա�O�s@��!}y��Q�à^N稚�tr�juF+v�G�i���s9�3t����|����=�-OV/�rvQ�D�4�R���z�
M�+
�Nǣ4<��I���U�\�9��n)>�9hY�&��N�x%���Y�
�ǂ�6*�~(V�!��eS���ZRd��8�.�ܐ��wi�,'�eץ��^jIa��l�{�־�z���$�}fuǬ�2~�V��i���RNnQ��%3�֑���>*�X��].�	�8�X.<:m��|�ڣ�'@�����㲨���YO�.bWV{��v�{ݼ�]1����Sx�oh�u]���lFW��sB"/�&|N=�(�܌�K��C>�a�)�6V���2�+���*i[J�ب1�S�4�� ��A�Epz�9���W��䱚Wno�k��ʗlJ؜x;���.�B��'R���Xv�/����L<��'���1�MCZ�xLK n�*#�B:�ol'����z�D���y�����l�qr�PY4%���
/.]t=1VNK��P^5ܫ»���ny�j_��M�o���
��bO��s�Cz�Wm��ٍ��������Q�kUon%��O�n}�䅈D��`�{��H=�b�됯�Ē���6�C�0���X�~O��d���s��a&5��fzPc�R�+Ԓ�RK*ãɹZ� n-�I���^�}�QLk�Q�a���c��c�k��U�@F���H��5��Ns�#����H
m�'v�u�ڲW	+^�T�^���ȯKdC7d8kc֮
��C�.>d����oE���f���'�;cr<C`�Y&���*<H�7v<� �T���V��4��a�`D���tR�$Ɗ}JW-�ݲ�W�d1�I2�U��|�=�Dv�x��m_�!_��;ϴsh���דM�]3�tK`��N0�4/�	���!��#N�4h�K�/lA��=hĂB�����������RccaVK
��C���d,���b�l�[���g���	K��i7�̸��FE����QmS(g������A���97P�2*jTu��)c��H��H|>^��M)��DL�H���u&��uU;�[⢫�yW�������u��a���r�.*���?��U	_1�z���eY���cq�������O5��ʳݩH-kf��e-�W�z��������,��J�pZ�*^�$^x���]'N�`ϰ^�o�����יִW���x\�����3E�U�A9���������(a��wQTIUb(��{�um����hC,O��������&f���w�%�<Z��/ۊ�|l}2�՝~}�V}��
F��/@OJ*�>�IM.��=v�E5d�����O��\�ᑋ�����4�u�Q2*��a�גX�iN/�]$�G�b����eᬀ��|?�ȼy2Q�%Nil��
M$- w��SY��rR��m�� �sd�a@v��V�����{�YӮb�� I�s%�nTqBu�z\��6��w%�vm6�&jfU�C�%B�m�a���5ծ����llx�7�[F� ��-�?���X�X1�Us�^O�`��\-ڲ�ڶ�e���.N
���ľO��Mw��U�Ȣ�-T�w��o2�J�p�rl��N�:���;d޲��v{J��^�䯖��v��E�\L2�9(^�z�)4f�[G���S���:]!b�\w9��{��.��?g�1x�Kh�^�Ě"�mL,��s��#�X�{���E�#{j�&L���8�4�P0>ꮤ\��6f�q���Z��lp1pYM8W�0�ˠh�&����%婵���w�����i�;/�%Cu��|%���wq�_g���r�"�db(�ǩ�剕�!Y9�)��>H�ԩL�T<�H�왘Xw�p�kS�V=&f)��5���&yb؀�2���C����{�?��I�*K��9�Lu+��5��R���I�&���<�R=��*��Eet��4�0wY\eZ�̅�ǽ�}GZQ�d��1S�g��V�xA������a������9��)�:�L�)�s2g�J�(��^��<����4�Ri�cޗ�f�E�h��:7�z��-*�̵۩rN�n���W��R<��X���1�Ӎ�!D�1�HbfDf8��~'Ϟ�e'����]���N�PP�g>=})?��S@](|	�-���-pO1��-_6㈯62lB��y�QU�����U>��J��HyVcj�t�@eN��	N(��-���1%�����R!�bj׼��z	f��Z���z�mZG���U8��j,�C����z���[��l~W���3����5���"�޸��*<RO�9��r�2IE9���|�<�úg�-gp�Re�lH����:��u�Q.�����$�	�#}s�E�M/�y��fQj�p�5���{fZ���@wI�Q���cV�"��=1���/�ѳZKT���&�H������:�Hx\�����{�n	�A/�ӎ5����v;|�1�HAW��ޔ�R����`Α�|��x��G�;��d�����2D^��u�z�j�=D~e��" x���%�����k�N�a����(��|�kQk%W�6����$�̛�7b1��K�E�:������,>�,��ƾ��~(���b6bP��厞��"ܥ�\2�/���:#Y�.��⸖���qL˭mK_-fRiHb'�G��z�)�e�nkYwe�3=�&����֚��gz69s�`$3�!q�HD��^d�'�f3̣�������&#On�@p��{�f�XE�,�kk3���`eҦ��;��}��p��1�>�o�`-2�פ_i��&kWT�,���;g�&�tà
����
��WKV
!�����cTN��/O�<^�)��������!D�Yy�x�S�c�ba��M+ӣ�S
3�M� �5'��ʫBpư����>���'�9e���{��[�=y�5�1(1�z��]�~X�O�"!�j��6�����u��f[(p�CD��F ��u���V{��H���P��p��|G�1��	=��S4Un��?"R��<�獱��;&|�����բ�QXk��{eK8��(ʜjR覆o�g����I:�WF�r�c_
;&����N>{��7tÃ�9kW?v]��5��k���AM������k~�x�Y�лo<'������͓�Mr3=���3�h��0*+,*P�%���D�T�f�(=���l}�d��SE����V
O�7����!��^C���OT'���y��}����S�L$<Z'l���{QYtZ��6����7a���N�������P}�6���]v�]�,�"�|C^��{�X�_gO�jD��ט�ǽ�/+�w�^��#��yR+�t������PM��� �e����t��a�Gv�k���u���N=��!0Jnr�!�Ƙ��̗m,��s��0�ͪ'\@�J��������)Y�!��J�b�0^ļ���L�i��RĂ���Um�FE��<�kI�a?���!a Fe�����y��w{V�BIOKvC�UC�C�8�ҹ6~�~�!���J�anΈ��&lF�© �أ��k��ߔw�.���E�~MZC��O����6?m����ln3&¯����6i(B:O�DTU�u��j��Zj��N7�4(��oY�k�4�z,KU#ϧ�݄�.ٌ�d]�dc�,�!�p���ܼ�o~W!�^�>wG��|���� wN,5"֋�s�a�V����.K.�ҁk"���Fqz�f�K[6�w�D����+U��4��}V��[3�Ъa���K(�������k��=�p�S�l�a�uJ�플�e[c��{��ʟ����F���^�u5m��c1f,�}�.����RT��#1����<�t,���K.pX��rhN�y�/݋�
�W]�!/�VO�EG�h�R��B��p'ެ�*�&Ml��'�]��`7�$���O��6�N���x��H���,�P�cq%��65Th ��V�֧H���Ed��䆯v��4�����7�bm�4���������1m=S���#�����yu՘ti\pC��g�,X�e��du(�r�>��j��H:B����C5���m��9�W7]���е�ӛ��2jS��r�u��F�EQ�p�!r�T�c����J�N��
sU�hW,��&0�8u�O#1Mt(��c��� s�@w��'�pN9y�Y��!x�8�nW�-����	��΋��a�J 8�/��}�����9U���8iA�4ٻ�G$��v"��k\�}W�Fd���ø�jZ�q�2
�X8���C|�b��J��,�i;���B�Qx��Û�����b�5Z�`�,W�.�!/�n�x���y�0�h�8M)���j��lc�Wj���P���q5s�K��-ڍ�k^K��'v��N�b]b�E����,k�*��h�* ���:�F��TL�����>�
����K�o�W��4�t��H����j(CW��S��J,uPwԙ��W��K��׏zf����ߵ��?ڛ<lCj:AhQ�)��ȯܫ6-�g�?p�CD8���A�.''��J��E�����~f�R��6᷺�kaC8��pmWU�����W�˩�OMF��.!m��C�Q�˪�IFuJ8�%}���Ȱ���y��B���M#�0�ُg����B��rn��}��x+)^P������Ҙ,/h��L���A����A��a�E��n�:�1h�2��V��uM���x��Am-�ā����� �2�J1���TFɲL�u\.0�E%����{�b́d"���k
�Rq\�22�7&�F����6�)�����d 7���Yz��ż阌�A�P�e\E\��k'"�o�j��
tb���M�C1
:Y��YT��	$mG�jH��^@C���)Ա���a��U��*��cF���]Ib-G�n)		�g��Кmd�p)�����ְ�W-_��_�[���-i�-{��%�k���=��1��⃢�qx���&=��n�� ����n���E��y���f�نT���ر�g�C�Gڋ�%�8-ѕRl�uYű���y��)k�@�b��N�v~k��f�=)6`0>���:��瀿PCp�Ka3���>�(=%��3��f�Ӆ����5̵�q�ILS���h�Ø�@�1���>�_�����X`��4�_�Iq�>�
����U��e�x��8�f]k��V��:��-5��e;�m[W�o��}����5��k�I'п��Z�y��01���rUy�"���%%oy0'.W��V�(��[ɚ�5���F��$&z����g���N-�6e�g���$f�N�揓v�9m�
tW��P�ڌ�5��/�{v"O|v[�(��~���Ȅ�@��Q�Z=�Ю5$�����3V8���i�n�>�o�����cӷ	�jn��GZ�@����v�Hca	����=r�����Y%��aEx�
�%�$l���cO��r0&���=�@�o�`dFu���'��d���%��j�96��k?�4���z:��V��O����:��Px-a$�&��l�f4nC��ޥ6[�*&Z��أ�%����)E8�B�CK����ZT-b��\�����،�.@�CׄR^G�Ҫ�M��]$,��l���L�y�h`�����Wa���4Yf�-���&M�5�H�H����T���X�sɫ�ѡ{c��}���=�{i�rkuŭbp-�,�/��PT%���A�ҳ3�)(i*, Z�D��/����WW�i8[����*-ks :�s/�I�2��pT�Jv,��uU��W�������)D ��wa*ٙ�ὶF�WM^~�&3_߼G�gB{ߴ'�$6����7�S��F(�bRE������<�I�GX�� b*/�-TH�`IO����µ��|����|�og�VNJ�"�_�밢�Z�y2����qo����d�{�oV�M�'{�^��]�	O~����jVK^މ>,�$�0<p�|����!N�c������Zk���	��ϊ�v�c��`��Rhܝ�ˑ�YM�Y���H�Q���(�ۉ�*���ZLt՚��_Q̔8sSFo�Q�����j���IJR��
S�Xq���c�(��rwh�=�L�s&9ZCw��W�۲�`�:ו��u��ap�0�>�Ӊ����6'���4Y���)$�6��F��r��[�ŞpzÅ�Z���ƿ��$[(��9VyUf��	2�5��Ŀݣɏ�4὆�%cVn5����z�I�E��q�ZX���HKNX�������O/ϕv�p׋� ���]X굗D\�xG�+mHټ���K@o�Bod{�L`=J��I�V,�R��A����N.���^�x�2s�Ϊ���7cr�|XуXR����~�������B�k���uS�k���$�D3�,�ѳ���DX�_>��:d�߽}������n���g�)=?�z�@f����$���cj�6��!]��'ʚ}F���W���g��:��:l�5��Đ��j%[T_��0����_��&F�A�k�������n��p_&�#|��R[�_����Eq����(H|X����F��1}*{��M�	#7O-L��A<�5��*�}�����\���=>4����߯w���I����I�A��u���[�)YZ�]�m۞ؐ&�D�C���/�m/ڞ��c��?}�֤���ʐ֬�-zK٩�E��^���2��h���ɛ.V	�����$��ca� p��zz��W}��d�J��;6�E4$���=���(�K<ɓ�*�`��A�v���7i��ITx�#-@l`���W� �څ�e �]0ۓ.sS�RSU���]ӫ�CN��4W���,�|O��*OМ�v�2�.�����s��
��oa��1a��&<�ɧ��+^g�Rk7�޷>ܳ}F��^��J"��{j vE�G]�m�5��:�p�H�!�Y�t`�2���ϱ!(�<�QÚN��|��Q��Yһ�BQ.ZH
�b(h�JJk���"g��]I���3¢��tĭ������azc�k��#�ӣ���E�����ޢ�`�I_v%-j)�2�Z��۩�K8W4ص�i��u��Yts�c���_-�	�i��_vk��WƳ4xWJ�@��Q]j��J�PV��T�?���±�rg�M��tx%ʞ�(�67�{�g�A��>��,J�_�����L��~��&��<~�m|���D'��J��9�cj9_%���%�>&e��Z�W�'�-ԛ ��ϗ:ָW�~w��N�K��kT���W!h<��١ .�;�Y�b���O�ɳ)��v�alġ��lQ�)H��1yj�.�$U ���B*��B���b�쨹_�o&�H��MY�� z&����4 P��A�>n9�ɬ�xɇ��b�Q_���%��ji7�A��Aǵ8#��h�]$��R�/
��@:ņ�t����'*������O�c%��]�?q+%a��#��,����کo�r�F�ڙp�i�=�t�@=rb
���ӧd~�3#O��(�|TH���O�FC�C��������R�����ب�k"{�R���kRv{=�ad�P���5�MN5���mwG����ҙ8�buF.i}5�6���^e��W���F�I���W �2�^��{w���P?�֯	�����y3�Q�=��DX��G���ߔ~�!�"]�.�[P�6�O�2�Y�����>����� �UZ�;Ȑ�HSV�B���A�y9�*3���1�>�]�n4�U��Exd-�;K�[K���Hӱ&�����2f�lƲ�Å�UjBJx!{����AӁ���8s	�Un��nA/�	�c�WV��6��]W�|R2:({X����v��Z0C0�Qʌ�vi[�&JO�@�� �#�i�1�Wg�����*�q��:���;[�&�>���#"ϫ��?*�(&�&q8L�6o�rԡ�KU,c�&ޯ��P�B%�U��Huߵ�m�u�Dy2���&��J'Ls(.[���*87�}�Fg�Vޔ��.�V��Z���eؖ�t*�Y�5k�R��;g�>��߱�u瓱�Qz���qI5��H}�Ixd�|��WjR2�[[�2LiN%v�>C�e��劒!��`�]�+�����YU>��|&Y�5���+U��M����a�k�o� �#�͌j�a�������nI.�q@��t,��'N}f�Oi
'G&�#���m#��_�ەr7G({\#�����>W�Rm�.���_���̿�՚#�U���A�5��&��;s�GpTw ��~��.��%s�a�<��Sb*l��Q��[{h���G�w4up�?�ˌ{�������> N����c���Tq������L(�`�}����k��1��Yk��~޻���vdL��zN�ߝ��`<{�]T��Y`��c�����}FC��!9��3�;/���0���]��X��O�iD
\��P4��н��ߗ��`f�f���~�TC졖�RF���Ң�&-.��!bN.�C'��d�mB��
wJuA��9�,������X�;E$^b��f�
Nv7���z�]gע����N@����ow��x#�����$V��T�/��u��ș[�WKW)�X���G�B\�a���YJH��lP-'F��]l�����_����x�2�����}\��vVoX�zK�x��
��kv��0�W��ɧ��:B'̾�=��	Zp�"���D��=�j�m�t]f��S~MV��y��ૌ+>J��T�p!��C�v�]x�"�TY���(|�Gʱ��P+X��.�I�$vk�[f�W~6���1^�É��5qVg�]\	��H��\v��K��b�L]�A�O<q�X�6���pw4��d�W�L]��d�4E�%�ׯ�ၗu�3�{k(�p׵F)�h��|��<<I��\�^��{��o�x�L:�#��R/��nc�'1�eN�cO�X46���e-�!���J-��0?�#����!�[���=��J
X�)�+@Y��X�g}�<^Y�W�_���s��i�=��P8�v�� T�Tn/p'tR�II��a�l�)1�(=,P��� ��Z�!��D����7��L&��o?��'|���}uH�A��rr��T��Ξ3�!�����eb/2�s
yX~m��1�u���`�OYpb����$���=��T�W�*t������^�`�r1�W�pMzT���1�Ga���yʄ����'Z[THlWL7����5�Z���=Fٮ�9չV�ti�)L�r.Ge�5KlT�����h_k��^�"�(7��б9�����u/�2���3���L�H���ʊ�X�"�I��N�α�Ux������h�c�u?ġ\J��u��2����hc~���>���Qګ.m��:>��_'�Vҧ�������rQ@�!���^�4��]�@Hp����j){�֡�g��cm��bm2*���������Y}�H���y�ʂi3��}3pMY� J°W�N���;�Ђ�;�@:�q��7e�[��5��6+���k9���vV�F`�+z�WT�yLT�Q��`9����le
^ʚ׽�g��ݡ�dW��Iz����El�(�KO��J���lf��Q����ccٴ�)�bp�,��+g��,�J������b^�\*��ZoaJ<�uO�C�n�hWҳ��/湫(���+�r�5���h`�VN�sOOĒ�^߮���-��/���<�a�0�Az~*������;b��;@M�lFN���\�SVRU#�1�����q�غ�U��zZ����H*�R�vv�QT�I���hWvE����ʳȠv��w�B�gu�8W�0�/�ad�6����׀Ȩ�&�����%�v�u��`ɚz����L�~8
LN]v�u5ު�C����7��t�����:�g[��U�����r�����~����z����WU8��q�XǕ�A�G%�����r�$�Eq�MV���ր����r20x.�+�e�"�(���.��n|f��n������6�P�Eg{O��3� ���qW���-�V�R�x�N�B�j�j�t(MJ[�
a^�;�F�uX�!h@7ʆ9�����"�b��� k.&:D�|��һ�r�y��Z1�"��a}l\%�\Aey2�w��-ϐ0�1�NQ���խ�ſ[���3�Ɲ�ɝ4AyȄ"��k�e��ϯQZ��\�`b�@����jed�]��k*�ʬ��ޙ�[x��wmw��2K�����4-�$���u��	����*#{�UȈ��jL��~ތכ�S'm�(M�����.�/[�������"E}f�}�y��U��5����oa��ر����7���x'��)�s��V��2�w)�R1P%?=/������#���G��s���;�Z�Sw�z��#�]������ꂉ�\�r�a9�>�k����ˀ�69heB���u��}�.I:g�@}��Noyn����%�̤���]I����T�-,����΅���@��̃�ix�xN�<; Ng$�JI�0f���DBeύ��֒F��	zi}aȖ�Q���>.����Iw���ғ�����XފJ����!��Ɵ��T+*��SV ��g'�M�Ë�ܪ�Uz��]Զ8��%������`h0��y�l��y���G��a�o��S�~a�`jԪ1톒n4�7F��K�͎���ǌ]_��<w��c�S$��zd��h�)A:��;�{���W������*c��rۀ�u���ǜ��������8�=�JeH�O�;Ц�\��
]���h�`��9�a�M�����n`��0���V�i�5��4�4������P�<���V$���&�w�v�2��u{�[����(�"��������҉\7���MhR�W*��XC��v�r(&|w�bp�W
[y�TI5��Sߥq�ڃ�B�-��k��.E�9��Q��64؈c��w։ff��ϝT�FR�8M��5��P�;��A^(�.czc�`ovS�X�Z�$qm�U����MWI�����|�!�� o�vf��T����|!�c^خ�6��C<�=K@)/�a����Vb���l�L���smS����U��k���a��`�H:�X�W�Z��+�w�q�g���;+���T�ٱwה�D�*-ؐ���hZW�{�r�e��өn��;U�R�x����7���|��!�EP��ۜ��4Gq}_�X�]g�� <���,�X�M���/�^��:�O*�މU�z���O����3.�1�u���1�꣒U�U�K���ժ���b�4�.��Na�t�!u� ��s���Z}����=����$?�W��"����Lы���DI6���GTl����/p�_�n-�}�T�I9dg�Y�u�!*���ֱ��$�H�M	���6�-��>fe�Y�r�GJC
lu��{_�NMۘ�FI�P/Ah�K�z+�/�{ZtJ�#*C�^�q���I�H�!y讓�XzP>��p\��Y��0lw������EU����ݗ0��z�g����{L��ue9�׶��>p\��_��ܳ�;wI^�Y��Qҝ0s�!<�E�NF���:�7F�	����WľP4Ќ��J��6肊�"�6PWm�}^��~� �p��3����)!*�NVmYx�o7C�����|��L?��S���ۛ��n�����	����9��g?'n#���`���A�{R�G%�;o�W0�_������z��<��x��5�Ӱs[��lh���2�Є��1�d���(�t8�|���4j�^�ڵ�h�\m��������Wu~cP)���0ŧ/U��Τ���N�8d����x]/5qBos*G)��|���f޾y����R{���?$>\�g���V��}�ކW�\�<�
�'���p��r�ȐJ$�
��0/�O1�0j�-N������~���a3d��fj-PrP��}����N!�Zq> Qb�ڗ���Q���岴�Ɲ7�s^�P�to��iv7��D�!������j׀U�1��sh�&EK\����xL\2*�8bp�#�h+�o���W���Պ}��U��Ry�v@-����x�1[-פW�8�0�n?NFE�'޾�uτ�SR������GBzO�_y/�E��%���c�哆1�I�4��?���ۯi��9���7T��t�z��I�i�ik��͵F�N4��<E�Y��vuOmM2f	+��7��WiFV*�Ҵ�v���n'�Vo`��᳼�Evy	ٚ�lOq%*v4U��Pib ��Q�]�B�5�Nt,hj@r�Gk���9��x���u��5!��D�1^>��iJ	-���u�lI�N�x�yI��K|�b���(������0S;g�"9�z描��ݷ�E���qd��D����^e���/5�p�P)bnҤ}��J���UICL]QW1���g�e�Ϟ�AX?�:�3kG�bm���~	��0�1�`N\K�зrX�	��t_I�!���m�Z�qa���A����gy�c(vUϓI-�=YSC���"n�\���y��9$��B���r�VC������r�����DR����o�h��K-�#a�`�H�w�-k��Ŷװ�0�Ad�U�F�5���_�Sݐ��7���I�I5r�Mo�}I�!����o�H��r�.i$6��wF%�B���� !d�W��J�XP�F�P�����x������C�����Bk��x_>��P>~�(���~����`�<���w��o�-�����trN�y'��YO���!T���*i���fm~���9*N&�V����ph=�K�e~�¾������]D�0�x�W�c.�m��������O������5��>~�@C0I� Lč���+��o����p�DT'>|?��q�I:F�U�0ø*������S������l3)pGa��ˇ�C�Ł���p���Z�!�A�A�������"o�^Q�-�2�~�n��T�O
����ݽ���j��|Q�5���I�I�G;�ų[�pZ]&�H�׆�Ѫ�!8��u�'S��r6�5�kCK��r�0�6l��X�&�/�H���`����������������oY&������{e ��oZ�_7�~��(%=�4����U�����Jj8$���gu_fZ���{N�Y�Qڀs9��5�qwҭ�?io�帑,n�Y�v��˻s���?�ͼso�%�T[.\@��[D0�����lfe� ��p777/�je��e���UOo`5�Y�,��Ř���y�(5��a�nb&�;7'KL�w����n�~��݈ޣJ�!�I�bJ�_�zI�F냒�ݵEg��5зw/������<FC0�x�d�e���׮⼏��6�&�_���T*��?E�80=��yO"��0ϼ�q�wS��{��MNn8��>`m��Չ�� X���Y����1O		�������<y	87�;trU�0��z�]U���\,�l,蜐��g���C���;�֕7�.�����ʅ򼷷�^^���v�f��%IL� �t���J�V��@
]��� &V�E�K��4DS�V�~��q^���>�CFo��x��e`�;��S.K���]��(,Թݵ�
�D�ƶ��ҕ�WlE�ڎ~��V��Ԧ��XH����wK���x��ϓ����ؙ�DλG$0l$�]7����
��fc��j��I�gJ&���#>��]�1��R�`�vY�x�#�������W���^z!�|��ۤ�o^+	�{��E�EY�DOlOa��$���#k����y-hKq�(�\<ZzzOG��^B����onI#�cѵ�eT�]Ȱ\G�bO1��"|��O��2��H1|?I9
�ߑw+�&�����X��z��=e�o��l�(-p�g�wi.=�$�'�B�&i�n
�޸���c��\�1C~�Q�I/QN��w3��O�Tg)�"�a�7$C��A��<���cn��B����&�^/N'�%��L"��:�� J`�--ўa�Ǡ�B�z^����B�s�D�k��m��Ebv����r��1��|a.���8E�-Q?Ye��ps�.P̬�Q�n���Ι��B���{�ŶF��xJ�>/)�-�i� �l#���9Y�ϫ��kv�nW?��Klԕ�ƞ�)�|��C�#Z%S�1�ֱ��|���s��;�;:1P�u-:�?��}���b�.1��r(�&{��}���X�����]���%��������J�Q�&��>|�A�7�n�_�|�L"�U�^��7<�.�X&h�_M�=Cg�?�{)��׺�9x���M���	��ŋ[rH��@z��PD�Xũ�f���������F�'eT� ����`nj� �-=T(*9��y	}?||�>��{��&^ב�ZGS6\��F�U�GM}^&�)z'9�c�;m����a,p�`|qm���J��qz<_,���y��m�S�p���b�l�wN^K�������uЮ�`�R�Dv��+VD��@CH���������SRiK,�:��=�:	f��a
����QYk9"Sx�؜aH�Q����=U-��pJ���Q��!'��{R\e:fC���S���~�]�%�a��p�D�� 1Ίs�����^�d�+���9i
T��E��	<i�x�T���Y�^�-�']m����5:ӐV;��M�l�]�`Xw�܉�-��� ��x�[��!2�S�G*x@��-�gL����#V���SH���ǔ�iڎ}�1�d��ݨ���M����/���M�>e@!j��#���o<Gx����+B��8��n,Jߞh,��?��=�����~/�*���}QB��h@��c�G
e"\���=>V��rC/�~lw�v����,�	^��~�Ţ	!>�s\������o����n۱D �c���M���w&�p�?���'lD!����-�|E)�]�U��*�2�9�<�����#�ae�}�H��	:"�����bQb��@d@�Ї԰n�>|L���W���74·	�s�U��zcvȶ�F�����1Ģ�{����miC�4���A�ݹ#k�tR~T8�~LA����(X04UwЊ]�v=�܎c>�~�N�M�%\��=6�}�[��;&os��/+�e��9�i%B�&g�M۲�7<�� �>ĺ�g�w�r�X��-�'l�7���f F�w�;�99�k��.*�9�:?�y��0?C%���<կ?��SJ%{{���n�x�2��T;�ɑ��"�w��)ė����8���U(� �]*e�s:��Z��C�"����(	�{�����BNx�x��������D�u?�����;>0";�T�םq���ijڂ��+ZZd$zi���?�g����W���d��cū�嚰)�v����.�GD��O?-����IK����!e�7���m﹡2`N+�l7˫��+�*���>2{b���1�_�1%�S�G�X�⏏bJ�C'�-���cA>>�>1����ȧT�A�[��
�7���נp1�E�\�����{�J�jYV�ʉ�����2�Wq��n����pe��8i�xzZg���_�{;;ic�k�5�B� fCk�O��$];Q��	{�L�G�q�%�����wW'	}4A�D5_"�\��3a'���1��,-��l�y���E;3�*��D��l�y|�q�V��B�)'��J��-�X�\v0���o���6[�s?�~s��J��.�֢��~4��B��T73�S(�7*C�wm�1أ*0� �W�ccq1|_����_��z����aL `wL�8�8�F�=m�A��&g, ��Y[s����d�g��q�bl'�1f|-D~OC�ب�tՂb#3�D/
�Ft�Sb1�}v��1)�^��x�{�͖s`Rky#�f�&y�H�L��Ѝ2�0\�7�2��x¦���^�:r}���%�X�G��~Z·��i�F��"�!�EE���hl:8>5����M�Yo>+q2�ksFXk�� �����y�]�xo�?y3�|M/C����Y�;�1�w*�#x��B5s��7��u�y/��:X!B
�˙a�6� ��5D���{�C���ыж!�=��xraE�(i2�p�po�4MIf+Y-�.�"��T�"��!�u�"RD��xy���:[_+��F����e,��/�Ϥ*��_�;��Z{c�uf�Ύ��w���`Rt��~uU��^+Nv��`�_��l2o/��Ljxv`(wg��2E�,_#��f�ey�K�i<rM��7��_:p@y�eAX����;��y섛�����L*OOr~�r��mf{��J�um�3�aHʈg	G�݋.�� 煨�bD?S6����cj̫�"䑞X��ǻw�;�K8�٬s)��$/��KдC��F�&�� �o<Gb-=/<؋�<�kLṹ.z����y	M��y�.x���=���4�i2��k���8����n).S�԰�F�X&�f��5a<��☙x��mDfYZ2��cz)�R�+�[ݓ� xa�xi�J�z��2xrH6��WQ��S�LNFS�
�B��gr-c���2��U��GZ�\���#��NRTV�.eCz}M)'�T������	�����T��si�.H�,kВ*�l��nV�_��7��������=��h��8�?<�B��Dty_x��n,gv�s]�o��1�&'�����GQ�Ty˓��pܘ���7�2K�b#K�)佨C���B_�ÌZ����X0"�u!ϋ�7d.�0��Ы�~�P�q���<��z��sm7��Ԙ�t�=4=�K�7N�F���*�ι�f�,b׵�E�e���$2*�_��7����EL!�헋�UE�E�^yLMQ�r�Vx_�>Ĝ)�ӻ̲�'�w���r��L���dZ�9��A�r�<n�ϕc� ���.��!�����E��?��k=Mj��j�*R���M�w�^�g����ѹ�1�xN+4O9��b�Xm�}Ӛ&��F��_Z�#	馀hi�4�L��|��1^u0��|s�6m�i�N�R02l:�U^W�t����S`�K�����쉖��i���K;�Ͳ�;�������{M&��w��.��09�AF8��M"N�����!]#�O�OM�XG+%s|�P�#ͦU��E��SЖ��!isI'��u��P�"�'P;㚝�%����i]����*_.�A��""�4n�5E�������=j�#��Q�Ѭd
զI��U^�|�.X/� ƄP�z��H��
!*iR�J�c*�p$�e�ƺx6Zt+��]c��n��Z&���a�?�����_���{����{z��5y�H����d�Ԋ�c���<-�� ���a����
s7ߟ1�Ѵڨd(�.�Kѩ���;����iP��GF>�Qr�z���<����������$���-��)�,R	ׂ��t�!A�k�9wI8��KqJ�~�\�܈Q�	M����/A).wI�z�[�SV͊�t�x�!&ݏ�X;�<I��.��g�ꂻ�� �S�.�a
WX�z�;�Yq�}³�8IJR�"5�$��F�{�Q��E(��}�/l��m$����5MW����gc����B�-���1��a����v�^�D���� C�
$%乖֨nP�kL�nY8���ь�s�lK1L���F�x��` �%�p�4P����}��t�<)ک��[A�gM�$���N6�5gj1��!킃��&=!��4�Ԣ,u�g�h��0�'N*2
F�$!��0<,=]�yw����FS�1P��uC4M��@X�����I�Y	���:K�����7DR
�������_�i����p8�-���B��$�1]2N4R��Y������?��H����].�w�Ȭ2އ�p� ���>�cj��9�3$����� ��p�����&ϑڸy�0O��r+碞�� E$�Y1��̶��R!�He�EoL�18��\ٷ�Á{ Y繶nn-�<��@c��X�Ѐ7��\Z��^��Q5$ش�1�m�3�uQ��t���K�F���Bt�ק�V:����P�:2������]����6��o0�/=��p�@%%a���nc�3xͤ;���	/�\J$<���=��Q�͡1�F��e֏"Ja�h,�p�2;��q�����ͳoS�Aۅ�!�ζ"�z)C�0��`����D����I}��1Z��Z�6�͍s���4aD�!�A1�Hq��m��D!p�Cx�����E�ۻ܏�c���ӕ-�8@�z|�s0�i*���ď<�˘�4Y�h�n��JeAEB	�o���x�2����i�x�;����Hu]��t�^<ʮ#i$B0A�}
�(�t�c��'])�F�*C]|GT��﮷�t'+�S�S�Im����;�����F����*��+��S�%�D�/�Br�O}Mycè�[[�S���  ��IDATPYe��h��(;1L>����� j Mlw�ˢ�c�
8?P��i�P��>VGU�U��1T��WٺK6��IY|9l�i�b�k#aZ�;��R���Ą1�<R�'9��LĆ����
����S5��l�$�s���C�ɆT�+)����R��\e!�����`pQ�O��U���z��J�[B�.>�Lm>�%Qg���h�E��7r�����6T�����{�8��Q*R}�<do��.��&U+�QB�H�4�������+s�rc��n����+��C���Ix��1�mh�<!h�/�7�Os;g��CC�-w���i�����Cђ���@"������s8./�H"�l�e�A�ܯ��8L� vL~�7Lz_KA,WG�a�yN6�l �5"��JMܤ.����g��ңmb���عbsC#���r�y5���)a�pV�a�jf��9�?)�L�@���K��Q���*�)'�\����<4NY&/�h";�ceg&�R, Ǌ-r�_p�\UUY<�<В���񼦚��\]y���Q@��t��UrA�RdQ�7è�NX�#���\~n(���~��=��Տ>=3�_!����_3�ƭ8.��*�,��5��h�4,7�B%���e�:��ء��1ӂ�KS��j�I�T%̬~�0�c�cp^ �Ls���[0h�2����F<D�RS7��N���2�n�^�e �Cy��2Kn�����e��FoM��y�<E,����\�&V_���$��>H��l0ɽ��Y"M��%�x&���!��2�����h�����C!����j�2E-{���)A�Wu ��y{sԝ�Bd5�&h=8vo�d�%�a�T%d�ם8/A�K���Cήt�uRr�)�*�����̕]pIY�f��eq�)Z��#h>��4bZ��
��C�����Q��%������cN�D�h�OA�p�P"7*Ҕup�	y���f0�_�����yj����aqx0W�~*Q�γ��s0c�Ic�� �E`�e���ju(^�`-�]�/ �#3dR.]m�ҏ͑H��[��ײ�_V.=���{@��D�3rM��4Iy�4	�^�=�s!b�h�	��!�X��vp	f��c޻���r)����:��>F��Ꮼ��*��ց��.o
���X��OcU3�(/d�b�뙮i���l�H�mB�t�F�'���Q��l��>�0��ȕ�-��J�c��X�zS$�0�0p����:)[�!#	zh�f��,C����TBAD�aB^P!�c��j���BCm�%�6�V�9�t�]�O�t�u��G:���:xR�����KR�Bų�u)���|�U����������S�iˌ��j"q%�PT��[{�1��pO�㮚j�҅��^e���H����"�@�
a�ŧ���6!w��4#a�D�Ou��,�s|�b�s�����]y�}@l�g&�wxٗ(�H3ƁT�h�q	��y����D�C��Y1(��lt}���x1&P}�z�!uCL'�0?��i�y��Ќx�)R�e�g���{4M����C{�S�*>A��	�H�x
��|�OX���/�Z�o�ʕ@�020�o,��KN&�Γ��N�v����YgC_�@0�����L���sL4z�{�L���w�sD����e�m�<�<>A��Y&"����B���Jэ�^"5=�>iLa��H�� j� CD̩����kc*P'��|���d=fa6�^?���1��	���af	�"J�`Ԕ�$��~�w�oB�c�н_�S<E��0�i�^,�BS��2yPG߭���|�N���x�00>���E�בOc#�d���&�Z'��k�͉�)6�>BV��8���x�S=���
%���7��|�??���it�����=�(�;&h�I��X�#˹4��ײ8�c�^�����)��󹌻���	eVMEx����d�x��[֭�t��]$�����׃ǣjXE�%ʙ�F�+Ӿx8�W~S�Oבy=z�oz����3��69;��A;]��^X/Z�n���@�'�j�M٧�ꬌg���̬i̝�R�\�D�Վ��x\�i'G�F���\V�����	Yw��7����5�����8�q����Lc�p'K_c��+��[NkVbWF=;�c����&&#��6�Mn�V���r4k�`ln��{���>��2�i����֑H�a�4���[m��R|f���(�����> �3H���G1�i,1�������K��^A�qoY�~����L����N�����)B7�{w�|A9DWRs	��ep���7�T�L��箊���56�ɂȎ���"9�8o(�xV?(���:�6��q���r8P�����Lرtr��,|�A��������R����e]
W�̈+,5���{{mug�����&Z��R���qiOm2�LF���&�Md�\L�w�����zw;{���K�38�)ڀX���w{����pw
{�a�c|.�z��^�Q�8Z��([��Ӹ��i�d6�F?�������8�ӕ!�������m�x��%+����U;ߵ��m��3E�e:-7'��I�\�C��"�]��4������_�_��b��u�0���ls�=o�A"��8�2!`��OU��>?��+{�\ΜH����B`g=4���2�P�R��Ezё���x��s�XtQ�G�q`��JT� ����a�~��0,��I��"�B��,)�O�/�%��U�2zq�0��p�3Ce{��̩u��y��p+�����ł�y"C
/_�u�lH�4��(�u)�G��U}���[.2(����y�P�8��>)ǿ--6�����0G$��ݍhW�Qv��L��d�`8Pi+��j�"�#̇��cA�����~3�w�$CNY;u����9����p�b�Tk�-<NC#��ǵ����
�w�tn&�%C_E�ϩ`��s^J97��.��8.�+�dEG��$�2K`��M��C߅�9�s�J���9�a�ٕ���SXy�_rb�3������<R�dʡG��P�QKa�KX^���b�V�̸�B�C��R��Gw���u��U�����	c2�uj�jX>�x�w5���I/�!�7�YO��`���׭<'R(�������CVW��T����CJ��PEb<6|?�x�@c�a���dC����V��^Z���.�7��L�d��Z��g!H�5���nh�`��3<��������{XD�w72�n�B�c�� �t��3tP�R%���>��ݝ���x�!�b0���E�H��d�ժ2�߈OyD/���孳�l����ȱY�J$3<.�#=lR�[��<�)�����U�N�,���65E�[�1�!*�MTx�0�R�zAhO;M�zMS���Mꜙ�Z���A���E��9a%��"0��0*�e�+�OB4*�<��������i� �Q��ې�aV���٨;
�\x���4�ٌ'�/��{�W3)j��\��s4�d��9o�H8f ��n�4��Ɛ���E6��RTd�z`�ƵJ��f�pF��0R1:��o.*S���ւ�4����rU�˽\꧳v� H^�e~��p���K��]��UY�%9��#�<�c���a���̽���*`����g�_����Q��91g�1�\��5�$�^�]��?ޥ�>.���2���q�-�4��<��A�Lx�sN���u�9D� vn�;��̃�B-;ڠ�F�#��\RM>#,<#�{�5�?�MC�ȋb�eW�`Q���㑑E����4l)Zu#I!&�Q����q�g§x�G%�\���bPV���1Z��>��I��UpsN�\Y�
8��g,^UI�W���ߩ����&�A��`b�U�J���>8Ņ�g��ھ�c��QZ�iZӠ*���0��̥�Q��sc���c�.���=�!��[.ǝ��yV���`��R��U���y��<g��{�F���}�h�n\M�*���q��_�����WZ����<�v�yҫu��-�Q`1Ñ��դ�S��P` $�fS��
����:�)���a��hC�:&�0��.,�o���Z!��0�0�W�މ���U.G�Am"���>zѻ?�To�?���%������5������bpc
"�)����*���O�6�f4%D`���oC?3�R���Ӂ	�!J-ɑ$��z�&��$���>�M���v��bi���%�י�ۜÐZ|��G'-K�ɋPR\^wauƞ�ߐ�{x����_����)�u%#�s����Py��a9�{W	nq�iT9�Ӽ�}��chx�Q�s{��8�J��� y�G�NP�'c$xԗ�<�Z������K?�]�E�����D�AY�s��X|�B����K��_⾫
̎�+��ؤ]԰�뷦Ja�\(����*�#^z�J�Z�.L�̛�%����N���Wخ��X�^�(���X�,��I��.����*��i������ў< _��]�K��	����,��%g3�����C���}��c�bOq�=� Q�=�߇p�<x"�'؆We����b�1e���v	�_�o�v��+�e�n�r�epD�j��ۢ����!O�,�?JC���.��X����+/�\���X�������>!�a5˿��	,�3���J����gE���IՎ����XC\ML^�]l,cL�K�6ɭ$�q�}��bs����h.JD���OJ�IG��J����P����4.#t���S����P�s�MGx�e��D&l.��c3>h����YO۔;4�i�(��oZ�)�ٳ����q\�B�4�Q�����Bvo�]v�9!��%�ߚ�,�,8��;���m$^�����U����1oǱ4�:�ο��(�E�-���t�5�Xz����`����$[]e��Y�c�{l�.Ӫ��4]j���Q����O�؎0� �`�VT+���t�(rF����M�����.�uhoRrex��+{�2��6R���Q�kL!a�ɜI�jBx�m�&C#�&N^�����97A�QT]t�mצ)��Vb�x[��r��ᖎ�:ވm���I����ي�<��V��x�������
�R�!��?�	���{�yb��q]sg%�A�H�*���/o�^)p�U���h̭� Ɓ�<ga�j�r�Ha�mw*Br�A�����#�7uE�L�_�+4�E�t-ˇes���-��"ه��k���n��,��D>qL>}����ӠO+�}V�
)>-�s>�����te4�mw�+x�z&��!���x~�j�Om�S诺�\��}�TIVV�r�Q��Dx/d
u�50��<u���FW�F��� sa
݁N��S�5ݪ�kz#��鄖�:�`]'�JQ�H����B;�\����0M=y���4?�4��>�{��I�MS��S���9������ƛ��s���I�%S(�H�]���.(N���y�P���8N:����ν�q"������jǻ�&pdH-���q�����W�>Ϲ��jF�����z��tYwc�^위1����%:`n���:g�6udh~���RA��S���{��-E$��q���5������C���O;���&}����}o{���s^��h�*hx��r�~�9W"ΏS6��U%�S���u�僙>�P��$Oq�po�\l�+�6�ʀ?�?����1�pG�+E8��-e �r��k�_��K���.�/��Nm�QE,n���J�޳0��z/b��%��M��T8k��������z%O�x��X���ɵ����-\�.=�pJF�Px3��S�Rj�ioiHk�w1~W��I��ǣa��lW�,*�v���*ڥ�N��M��Ѵ��wb��#��1�wu�9vWu�(���o�i������Ƴ��<�aL���đ��&��� �k�ŋ}�o��ֳ�d��ܲ��-C�c��`�L�c,tL,�ﮌ`�C��ϱs��M�@�&�q�x���� 퉕%��`Տƥ���\S�N�R�*�m�~���s$B�M���t�s�����-.<�U�t�Nkn�� ����6�+E��&�W�bN���1��s`K�g<�D+Q��	^5�!��E�K�@�xȘ3�迅�ۋ͛�)qxJ�H�C]��@�(]'wh�v�N����H��P�?e�-��Qrj�7y��zOǌ�q�-�#�s�,���S����<��m���C�����=���2�0��N��I����r{�Ґ�'e឵�Ѷ�ڷl)CXp���Zy��C���(
�C?BUfk�sa^J���6���+�ި�&���$���7��4�]��C�omʌ�&�_ӳH��(�((�d�d��9�%�RN`{|�6�ŘV1ͯ'�j�EO쑆�i�������)�5�!�4W�����G	�L�,<Ҩ�c��0f�4Z8I�=�"w�L�r�>�D�H����JS��L�m!TYGIh H���92��tc�T8ڊ�k�T'E�w~
����xۍ&�.M�͑�-B��-��>5A�A��]FѲ����LVcf)cg&E+k{ɉ#����a��-A9�v��GnX¬.U�Wi/�_�s�#�~Y����D�8�fv��<n��\�dkJI
쮄u��Q�O);m�V[�wӯ�N�C�Q��DT�����"�e> B���XL����k��VM�$,�y���?��ۉ�9���Բ�]p>*)�X�c�ZP����;U��8A34��jf���h��Sf���<�F2��D�L�f���$3�Ҏ�� �2�`�^�S�E�zHQ���!���zu%�E��E
c������c���a���R�v9Mynφ�lc����+����.0���ޣ^O�!�Ě�,n��]�w��"�!`C ��6Ё[� �N��Cd�Ι����H��@_��^B�b ���XJ��'.�I��{�}�*�p���qno��ciQ��YVO�;X 0�02�(cܚ(�LA�bM��vx��!�ҩ�N�+�ğ�wJQ�\�
�F��p�ƃ����ƈ�u�i*��<ct��""�8!�va]{y�YuW�>M�FXS07'?��!�W��w�D�OA���:,�x�	>g��0sq'ݙ2�ax����H&�ޭ+*�*�FB.N:q�jC��}s!���J���Q,�?ERF��"�����x��z 06��U"��9r	1gm4ovQX�}���ǜ"��=�K�S���Ӛ\�m���_��rTR�)�
�1w�����>�{qݻ�8s�#Ā�Ԃ'r,��S��ں��(A��C�W3��x.$#IĎBA����UEh��
��k���l�G��Gې�߬�5��1[��6�.��]��.�]��-#Z���"��А�dH1p��C�%=?T�DX��hCQ��M�ݴ�0Ȅd��W��E�3�à�$(���;���w̾��3�y�g/Q]t��]������2˸������e78�]܍+���������V�g鉎F`6ؙ�R��O�����
���a2*��f�9:��t����j%��+}W�����l�Jxh}Ty��	�˘��)��-�h�G�C�����)��Հ�_&='$-og�G��	R�tZ$A��1ۘ5�ԇ`��$7���Աm�eU��S��1k���.�N!�܍y��%�;��c(��Qv9�F�l������^ZES�!{��(ヾHF�I��El�۶�p�3lP������lG�S��W*��<����%���L9���=J�����؟�'��#�Y;��r>.+55j@⊘k���	}�6�Բ�G.4J�5!�9u���U��X��}�~.8�1H��1���7��j��Q&����f�������b(�ĂG�`��q	��A���$ٷ���T�<��z�y���D�>t�:5F�A��Zp�.���7�~�ԛ	�Z�����ڻ68�dkN
�y.+��&ZY��-������&T���m\W<���RL�6x}���Y}#f���K�wT��7���snr�!ƞO��-,�n+��������s]����fڎu]	I��]L噊�q>�+��w���&�O�9� {)�Der�*n9�\y��'�eG���#�A����Vx}�ы����H���ܠo���͐G?i��gvy�MO��Hs��/C�����*��Sb󒶩� ĭC"�d�K������͌�	7���b+�/�;���b�_T��`pAm�駟����Ɉ����[k��1]6��@7��_�.Ag4WYc;��V���YI�ψ� s&�A��=������6��f�U� Rrɕ�Im"������k�����cri�@���c/�	�I�[۵Z����ҩ���v��`��v"���1�H�\i(5�B��Zє_��H�p`2�c�%y�Mϛ��x'��(t�j�kgWr��]�ͺoU7ѠEuap�՜�ؐ�ĢE�:��N5�E��sS�4qLMS����uZعWV�G3��6�Km��Ԅz|5��89y��Eg��,�.3\J\����>f�i<\���
";3�R�'�����1O���M�I]��d�8�56w�F�DjVD;�&YR�j՜J�����]�����c�x��G�#�@��jm[�0��5-V,���aC�d�\��	g��ɛ����E����Κ�N������]E�_5�ϭ蜾�h���/<�"Ag]AS�ܒ��i;����񯺎5y���n����q� ��C���.x�ێ�Aл�������d��ذ'�D�55�/ш��=��ۈk ��������Ń�ڵ-�xƸ�q�F�q�Š�)p?	�����H���D�U�d����7V�a%���X��~��#�߯Cp��J�����3A�����a������k!(a.e҄6�����U���ݠ#>��4
�a���x�nn\����|�}��e�Z՜r"m�7<0Y���>���a��2-J���]=Y�@�@�t�r�l\������Tĵ�%1Ŧ�W�K��=���n�E=�sn�33kL�����C_3U���f��s$��l�8�!^2�ĸ�a[�E�5k؞�&w� m�1�]n�"�2��Yb>�ʯA����!�\ѩ���]Ń"�i�N��N���x�Ϟ�v�G��+��kƔT��x` �����Aw���lXQ�ʒON�[���җ,F�&2C���τ�,	g"Ivg�t}���>�� ���vI��dx~��I)e}�r~�
�N5�h���<���R-�k���FX]�*{�����/�B��xٓG/��0E�ᄽ-�7�bFQ�[a�ؐ�������!w_mKF�<H"��7@�ݶ��Q2����������	����ڥ�%Qg$�.ޣ����\��������� ̩qױ+��^���><`c���~P���xF8d������1zw�o�&�Q�1)x�NܳKE%qe-�92���W9�"w"f�K�$��M�'^c����p��v$��Xc<f�k���6�H�vc(�[ fb��.Z9CC0{r?�g�k]k�+�j��N����L�gf	=�i%��0��.�9a�-�c��~�1[���o�C�6"�E	$$Z����ÑaC�n��z�l��T��\IԹIW٭��]�^@c�O&��x˲˔�̟𨰁��[���6yq�D[ʘKJ��c�X-I���a�-~5�OQ�}���8Gd//�>�(]\�!���h$�})�zr�^�>�FuCW���"�Ι�秫R֡8t���<)��H����5�	��/�Ƣ�PJI�3����Yb3'#DV=��J���Dω	��<���#`���x�!�3n�ίg��iL�x?�`�E%��	�q<�E.w�+�c�s��3�0�L:�e�~#�~^�!gx
������H_Ef�FS��&��V��`��jYG�F+� y���S'{���K�����1n�}1�p��T8���(q-�f��]{%���F��K$�앚cZ�%23V� jP9�n�##��Umflw�ƙ��N�`�'��g�V?Ex���髏9ciM����:g�bfE��26�%������f������5��Emrn�>X�N��6�5�W�켟�����Rp����}��榺����B�zƃ�	��VDo�K�[���n��Kf�+~���W�����X����c�x���y����1�6D9m�N�8��g���&O�K�g��&���}`���NA��=c��������H@A�xp���C]�>�C;����8WX��fM���B��w��n�*��� ��oB�%�=�u������X.+� H�f��Pk�!���~/���b���!O�9��	:a嚣}�U�6�@��C����2JB���<wBQ]��y��w[�:I�p����lQ��F��KKn�v$=)���ׂq�8��$G{�Ӝ�T�-ojF���������&��6t�+�S$�Y�����(��Xx��K��jK�?������9xN�G�*��q*��BR���&���5�����H�}Q�PL���ڐ������n�V��S_0'�R1������l	&S�d�Px��`�Quò!����U�h	��Dٻ')���ل7�C������^����Ի��g$fOS�"�>�hbh։�9�D�¹K��;�j��F3g�YN���]^�2������uv�����d���)�9�ǁ^cD%A�P�K�%5Xӵ���YGey|�D�#�p����m���H��a�=^�sj��T���̖"ژ;y�h�����:0�&��C�ҜY�*Rj��S�>o�K�������۪��gET�����X#�Z��V��U�_M�������\9B�H�1h^M�rv��&*�v����+���>�k�u$}�/����ӥ��l��S������� ��[q]`�Aߪ˽sR�+��rKDX^��}n\+K��i��~)ü��Y�IB0�!��:qh����-Cߝ;"��g�	�=ɶ�H��5Ì}����N��V���9��0�]���n�j#����$]�X���\D�E��<�x.?���+�6��A0�7��OgC'aܾ�*@���x�7o�r� *��,mă�XM�JR-X�Dr,��Pܙ��Sag�0��e�V9�M� O���iO��dvAln+D$L8�S�n���7�~�Gc{�Cqs��8�1����H|hvƽ�8�C�ŷ������H�f�3�h������~FU+���׼Y�sl��O�{�H�Z��<�ې���p�E�xP.a�*;T���j�f�-|����p\SzJ��#�t��Bg ��k��8��J�[%��}��-Q���6�.wP�XQ�7���bH���1��M��%�"톈j��~M�p\]��4���L���hx<�`wr4���*�>�/���}֯%}w��ژ����@��y��l2%*B�|�eeꨋ��2E�O�|�u���9�}����&y���$m�%"��+P�re��̞&B]ݤ&9	bH��%�W���I�,	��U"�U޸d�j���M#TQ\ͷ��b&����v&)g��Ʀn��<��s(��`�3��Ha
�!k���)��U�5a��ish��,T���nB�x^󜮼Br������(=T)��0pq	�T��>ۖ���R<���7��O��*2��H �wVfB'(;T�jRM��XƗI<Ѷ�`a��)������;ww7���S�=��8�J's��:pe��HV�P����KV�z���J �kC�(�!�4孉r'���F��v�2�&0w�+\�s�)UWT����!$����N���M��^_D���K�r�g��!h��z��)�zI�����]����[�o���㻹a�A6n�.��H��{��1��������"��U5�<8q�{���1�Z�#4܊������w+$n�]!�w�C��V�!(t-ܻ�+\��)b�2,��y�İ^�� �EQVG���6㐙>��U�L�`4I�C	�mӔ>rw�B�LPŐ�,�ۖ�hO��"ߓ�/f��}`����y����yr�>�36������Ԇm���G�?�o�"��¯��Ǽ��C��vT�VA�W�>C\m+%|���h�7C�%�`�=��FmP|�y,d�CZ5]u�]�C���%��V�06�HN�{����͖������z��WB�(:�ΰs��T�����!�]�ެg{8ກ�tY{�1��x���~��ni0ב�f���O'��Ԙ�[W�6�%
��ę�h�<����%��5��E��-a/�`r�7'�,�}E�J)(]�\��D�e{�T"�(�T�jDdng���Md�o�K��ό�@\�sV�n0��ۚXz{	'�����5�4l�37�:B���^)�Yk�/�����I)y�hu���̮����jr�I��B��d1#�$t�t��q�;Q�d��|u�x��P*�/�C�L�mԕsw%���%,1xOؠW�pN�Ñ�ܱ��kNr�;��7�R��S/�Cl0/�^�k��[u#M�N1V�r��1�"fS#��0�?l���Tb�fo��Ʉ�%`����7V��:C5��Mz,�m�]W�S�#D���}{�?=E�M��I�+�7��]�v�9!�ǜ�8��a, +��f�jbc���P���4O����q�)7S`ԋ�r����b��2uY�p�&�t�M̑d��~�aĿ�!]��]tW8`�X�R
�������0�>��h�4 �Nv����<n�=����mx���KT�T��m�zl�\���W�M������Y���q�;EC�/f���x<0G\>�Vα�9���Q��$e�.ӛ����l��f�-C��ک������9l� 3X#�T%�W��z-fu�2���������4�6 ��P��I���������8��8�>v��>ǍxZ<�6��P�aHD|������յS�$(���å��R8��	����E����R�a��zHw'a��A͸<�@��͆�Aoj,�)L:�ډ�P�	���#�����o7�Øܓ����fW��7�M�,X.�l�\�Ŧ}w�93	9�P�Hno@���)&.�G�)p�.2���w�T�j];b�nZ&��2�諒��]�ʫ����-�0�l�r��.����t���@���K������5؟�չO���H2"<��|�jJ��i�$�x��;qbI]XsS-$���훷�j@��
CJ���c��mN��������Q�-����j�����Ԥ�%��Nz�f$����_��-�S�7b':sk�H��#5��v�Ϙ�b�L��zM�_nC�"�#C^!H�x�!0فg�Z)j�"�ms����yNn�Ҷ
�aH��g�q����̌��!3��� U�deE��_�u_㡳�|��/���!\З�K����l�r'`$����^<!l!%�G��
��/�!/6y�&�G�ʈ�NIv�o�h�9L�6�+��i6�H�r�u���B#�	�j঺��ۻZ�N�������Z�QgsK���E�4�:�xOH �,(ã��%����ڶ���6�x���88y˄��v�LB{�Wl��8���ڸ�Ɏ�\@Q\���%��:o�C%�p�ʺ#tfk��Õ�;��pC5Z�����D��;���6,�j���?�tSDT�m�>"�p���v�/2�(?V��h{�CUrd/��c$T���n�4����v�>Z���Ŏ�Z[���li�1�E�0@�C��0�b�,�b�Đw�r;7��(ڿ�������A�2t3Ny�?�K�]@s�>8�a�nK�*ZS��)g͕�*��5Dk���z�Q��d]�	p��*��1:����ʭ���8���=7��u������J�#��ԔJ��c��iﺴk��dNaf
���!���<D�0��=�7���;���V�Wig��2U��9H�[�r�+�RC]��_sQ�0n�%�r)d�����k�ׁcm�˅�W�h�����n��b��?�����)�=S~����m�/!w����K/o�to����T��K�
�.��|F��������}�.�+1+��M�To#���J,(��]"���ϼwmNr�59�B�ɭ��jD(0����e,�jV0�����+;v�c�YBN1eڊ��P�W��\�"TBC��������@�Æ�^�yI�0z*�����͎E�{��àc>L���ެKrs�̉��3��1��RlL��Օ=M{�b�
���2�R�K�V���!�D�%A��p8�y��T�����K�z�\#���n/�T��g�ț�߷U.��rn_�Sj.Y}�y�*�^�MW�9Z>t�����~��lSR��PW��0\O�Su���{�1dC�e�|iy;=- �0.�Z;Ĵ� ��u��r
N|�S6���esά {�;N�m6��@�>�d6�颤U^�1*,��lc��<�*�QdZ]RGjɬn�۝zr�Ӑ���\#��Ř��x���U�,���e-ry��L?]�Ncľ5˸���lu'g������zu��`���z��҈�_��62�T���2޷�/���������8E�\S��s_&S�Q��gx�cb�������!<�B��|����g%�#Gt��\ "�$~$�����|3��%�&��я<ɿ��s�I��,�#�!uG�1".i���]�w{��	�s����z���n2}�1�.��)Fw]�������K�ٍ2���M�,�!E1Fx���͜rI�;ǣ^�`���p[�2�`U�wj�8_R;?x0��XG�S��Wt+p�ϼW�d2�������霍mz��lG�lb1��=�~��U����}@���Mh�9'������Be��#��;ע&A➛���
�%$�p�L/��V��'�����x+n���Ԏ��SZiW��s�Xvu5QFX�q~�
�{�X���P`�W�7��v	�N��m4�p�/��9���x=Rzp1�ct��VJ��e�����ĕ�*a��<�����y���W	7���4�QE��6��N˸��.s|e0T5��nk����=���P��9G��[>�nJ-�Z�9���ޔ�8�t� L����y���ٚ�:�
/W���%��h1��@��1���T��I���^�z��k��[OL2��`_��=�3ÀJ�f��%��
����=��n�n�#Y���XK�K9��+��x�/��
�5�I@�mЋ��rDF�!�c�K�� :���ec�e1GO��:ڲz��Y9��+UkS��p����YU��"�UG��ҝ���::j�'��[M���4rs�%1����Ѹ��<_������3�$�zcn�����e�t�v�N�c�����}�u�M̹��g�Đ[���%lq�{�j�p\J3�h�ǰl���!3�c?������q@����m���Iҍ�!��L���U�,��m��D�������e2=�9�X�h� ���A���F�7���ݤW���:����@��y� h!�;��Z�F�u�dL�,�x���wm<�ɖ_��+�t��*�/�1ƔKy�X����}�w�M����O���۸�{�ܓ4��+�!U��zA�nu5����+�fl1b�Ô>}�ϡW�`k�@.��	��"qq?�-�������?���I�����=���ś<��#�H�lE7О`�h<}�~��46����zا�4
3��0I���7o���}������xhK�Ԏsǁ�����a|���F����������e��::W���B��K�Q�]�y���x�b��uj�6�n���u�ڂgN�D}໊Xq���=+������+m��,~�hP\��p�y��
�sl�EeQ�e½�;#��s	ӝHz�;G�n�Ve�W�J� f�fD�y�W�ȉ�d�z�J����[�|X������m}�o
p�)J��a�0)��9{/������m��n�]|�g�0��'�jҕ��V��ZR}�8�9��4��&��dVWO$������{�����;,��͊���c��h�a������&�k�L��vd"M�2�!ii4�(" ft�����;�L��k�h	!�
�Yh}f�,Y;c��
��3o���6�Qw��y��MX�Ȩ#�D:σ�t�E�^�x
�������9��O˩)�����Bgv�2�,����znsd)|���!+�K0f1>���!��ǟ�O��-���i�s����ç�p<-��,�ܔv�l�6��|��m����Ć��z�����o��r�S԰ҊpEd�œE<%�%�߿��OB`4�T::��z�VT�����K	p�� :T
̐D���I��t<��v�s�T\E�s��"�8V�I;�1i�>J�G:�=H�_�C)�&W�1a�P:8ݝ�/���E��7�0��\���S����]8���l9�E6�஻���q��Y?�kW�Y><L?EWhgeI]80^i�P8�-���)X �#ue����G:��u��u�L$Q�4��g�"הJ�8\�}�oA���9bR�B�*�T����}����v(&ҧ�md�&e�������<��wT�?g�-���i,����~ym�s��u��D��=����j�/����bDOT臤�n1�/_�`����B�?��K-��H��mt���ky	Lh�VzJ�
^���O�u�C���%d=�I"̫U�(��T� u'=�a�+��ό ^����+&A�m�X.�&y�����%�~w/�J�|nX��͔���l,�N�<\���}����2�(���u���P�m�J��p��(�Uŏ�~Z6�?ӧ������x!	�~>�I��C�0�0�^�y�~���?���`����������/���+F��w�|�FБ�&�	|��o�r�)?3鈱��G
���	M�9����	�w�r�j܏�Ζ9���~0��A�h,�f0��{%l�k�ޤ�v͹��i�"�9-�U:�Q��TրP⩋�Et>P[�
�{��Ex��i�ᢡ����\�l�Io�o��@ö�ŋX*L���336[��"��*�Ԩ�0QA��$�S^���$��.k��XX&�~A����k��~�;��o>��X�,��ɕm?���~E��ؓB9�e�<@X�x�ъC8�6cdH������V�Cb��g�ڹ�|2QFMё�	O�G�[���=�6����D��~ܬp��@|��Q���|�	ju����냐�LJ���K7�;�����f;y��g�q���0[8G�\Q�V�޾���U�7RJu�@�X�?+05����g�c83tSc�đ ��ɠ)�#���7�1CV���XN1����WA�W�!�r�"��	���7��X��	����Z��_����_����Y�.��6�1f˛����%0L/pm*�6^5����.F��׸`�Y#������74h�3G.�z��Ⰶ�+���P%�po(2-ĵ	�#��݄�ng�:(���ؚ�B�t���pQ��{�� ���I���o�NT�#n6��e.����3Mp����IT�I�a�s^+9ǒ܏J�����t��F4��Pj?{�%2�}��k��=
��Ե��V[y���hq6P�,���*5��y��1@$FT�'�[��jڐ��fK��^^�ƀ9�J�hC����\�<�a��}�����r�G�g�>D���g��i���2�{������d�����|�(�ؕ�N�(X�R��ǳ{�br�0�O^�T�*:��R���7�z�ԕD�h8�R�K�jwV�U��Z.�:���A�P�[4h�y�]I�9JW��e� &�=Q��cU�H�i�b�/�X._���^�,�����o��.}��w4b�Nܫ����￥�������8f��fk���������՝t�2J�W���*�]E�w�;`Pً,�7�s�{�����׋ф�y"?:�:O1�$�2j�j�'*B׼m�_s���qB5�ؤ�2+�9��6ox�7J:͜�Y��,��Ê�������Ms�(������in�ۼ�Ԙ/��/�|1��!�S��{S��`�h^.�|��[s�E�%��ls�^���=�P�����aH��u��4�~���!,��H��i/���M�+�ΉOy�~]������1��`���vhkB�1�#�i�1�	ə�)0��*W�ecó �/߁���k������)H1Р �A>P��z��XT�q�����d�Ɓ��\��-f]״[�ߴ%�Q��8���� ��7K��-ѓ�b��n���!x�nG�Rי�E��p*���x�G���w` ��ɤnJ0.��Kg��Hs��l��jX���au9�o��7G� �X-F��6(D	�?��<�g���_	�������^�����O	���[15L��:�31fC��jh'�d�)T�@�#�̞ߨ�c�j �6�D�_����s	����@��M�{+�{�#�d���+�fe��]���˜���]��Zs}���<�9��������n��=+!:DiÍ~�2Ow�d^c�g����y��HM��X8p���}�^�i��0�)��.'p�y�G�ϳ~�ިy'�/��־�H�U�)��N�Ōa����
Ƭr�c�ջ�PF��-��V�C�`C!t�6w�Ӡ$E�c�l2N��Jd�=�8�n{���&��D�m�i"�ާ��^;�%$[Srm��C�:�<��?�w��C*dE���h<Wa����n/V���G�o0�K�Z�ω�ϡ���Q�)1�<5�,��s�H�.���j;�ˢG8E���ZQ ;��@B<I�j50Y�ٔ���QPTc��ǜ�x?��4���ᔩtSH2�4y��!æ�ӏ?��o���8o@X�����@O�UA�h�E�c5�����-���jEDG��D��q��[<�r#bBF��(1�x���_hȥ�����9��b]E;�L��f�LC�j���?�9���ܯe��q�����A{E��"��W�ywںUۿ��m������=�Й���%��Ys��a��:ڑ�h�3��A1���ʓ4�2��/�����L	}Ơ�cP~N�nU���A���ĩz�x�]��J�ꎜ>��&�S��2�0{��C�H|t���� >c<EU6MrC0�ש�p5/�~o��؊��^D���w�ty 2w��ar>�i�,*�Zww|l(�L�s��a1�x��t�B&��I���d�>5e���;���l'��D�����e��MT�zEX7<g,Vp���Ar��V#�hEb5�6�0l*�4Q�|X��6l<��rb�C3�>,Mxw�=h'��~5rj�4=�(��#�2]Ox�?��st�L�F���Q���>���kF
������M������e<1_F�U��h]�1hEl���镼Ub:v��w�r������x̠�=U�Z�$�Tb���+�������NZ�AA�w�1ccAD"1Ϊ����0��_Rƞ!�)���|F�����{�'���D�Z��$��	K�'Ut�OWx��H`_��T�х�<�bD��m*R�*��q����)�o|�&���|��>����hyvaH]Q!���!Mj߻5|[�9n�T��  �v�]h�Ӝ��"4ڸ�{�	�{8 ߐ�ƚ^{s�-I�������0��k!��E{�d�G	�T�=�|��ux�=��x�B$z9����/���\�&w�?O��>����!�Cq�U@�V0eO����\�<�.g7��U!ԘG��
�`:DM8&�&o�wR�xY�jHW���K]�\�q�5��7�]�܆"3(X6�%��8�i c�l��v��׺׸V<r"2��8d��g�}�2�y�6}����}g��0L�_d����{�ws�������y�d�}��)�����Qe7D�K�V-Ԁ��DT&F#���o�����G�޽��>%ť���Ue߫Wo��m⸂�J��1�Y���æa�
y��@�*�C��nal���u`�q�9�L�N�*��O���&�
L��H��
�:����$�Wc�.P��7_x�^+�1,�)1�⸺i.t6:)YP|L�Y,-�k�(/g����v�7!�ڀe�6���R�����-B]��<K�g:gж�@��3i��N���6↍<R-��H'y��)��q�D��a�&(�kVBϳUh�rN{'}XL\5��ۧ}��1�v��=!D�
���?|\<�O�V�`(|�Lh�}x`7NH�a3px��pߝ)g�ex�:ҡ���9���Iʤ8.��H'4*d�.^S��������X���O�,��"%8nr^���0gN���U���S9.h-�ˈq�kK{%ЦHxΐJR��G�뒾����J!
�kÆ���q:[U��3�ىs������sot�ϟ�`��J��e�6o�8��U_{z���s����I��p$v�����ת���H ^hϬ�(K�7�4��+p���cF��M�Q��F��@�[޽^�9�*!��r��j����_獎%���i��a!�GCW5�I��y"��UC�*W��T��M9R!{`񜛱4 ��Yzh�����9U3Xd�
L���HSع�wϟ)º��c�u����R����Ӌ��R����X�m��\r&�]$�����h�4��U
ÊQ�*à���}N
�抩��-=�M�W�QGޯ�
+\q��ߗ���Ű������V��S��٪_g>���x<e>��J]�e��)q�Pk�����ד	!y�
��Á�		���;��� �#<h^Έ+thtp��ܣɚ�� �Km����~�*	�a�~�fy��,��RʃJF�,�՘��^+����p� ϡu���	��D�����ԃ��|����n��5�{ 0�*E�d�T�-��+V.�����t�/��̐~���<�:T���0���LnaX<\�\��D"���=�3x��k��H�k-$*��14q�3�s����͡�:��X���ղQmyk�j���p� 6�M��4���{��HD�ϔ$j�,k!dv��~�1ob��9c�8wќ��?e�Z#5;>��R�W�+�!a�d#��(�cR��vJ��kH�p���$�ֶ��7hO�L�YS.r,C�^@=냃{�{��gā\���Y���\�R䀹�md��zC�*Φw�3�R��p�$�a����r��T[��#����P���}�Zv�4�U�}�}�ʐ�x��"�F�E5C�D�w�MMk�������|�>Y�<�.!_hal���QыtZ��� `����C�h�h-N} e�����Ta�k0ygO��?/c�*��/"4��Q�"�c�)ƃ����^=zRr��^sI��f�1�!�r��s��T�P�e�C�%�Mt�-e�H�`LXu�d�}�~Hj�	�Q�f@A�r���4�#BoF$��� �똏�By,s�&6{lr���?}�!}|���ɱ�mw] �x���V�/��hvK�&s>�X�$`䍧��R�L9�Q"G9H�/ב�d�<燊��t��[�Ug
X���׻*@{��T�h<�q����X��B�չ�*�d���'GƵ!��Sd,����\g��3٘6
)Mՙ��h�dI��}���$���Y55᧔����r%�$�$�N��$,�H�X�͜�}�6)�[¢�/�M�v
!;�=ڻ�F����lı����D(#HC:�#qq�'JoT��F4�YLSeH�\Dzn�x��@o��v�2��٨�$%%k`̇h�P�3���;��O�5��F�ڧ?P��tgZ����L.��Q�=T��n'�Mn^.�EY΁qN�W��?0��&	pjQ��Ǖ�]L
�l��cx_$��9��5�����͹	�=Rx��,��T� _��c�ґ~�1g�?}��͎b�Q�&d���3�8.�����R�o�~C�:0B#5i�u<-ǖG�t���%.h��F�$lfxR�g^�M5��6���n]^�:��lE`�xЈ�8����e�=ۮ�����l$OM�������	hm�q]���)����>�?F0P�
-j/O{�ִ��4=TQ�;)sqL���S�m_پ��h�ƪIW;�W����w¼&�_ь�9�p殄5���B�R�a޵���2�Xp��|c�Τ��Т����hʓ�������v�����@X�(��g�v/u�u��n�';�dd�Q�V��h�"��c�F���*�qTP��m�"E
|�Z��g���'��mt>�՜ͯ���)ZN����t��8&�]"�p,L�t��;BR�����}�޲jG�4�V��iʊ,ƠD^����Us�PN^Pm!{�Ә��%5.ᥱ\���3u5;�J�O��B����	Z��q<ED#e�5�2B���u�#7l��D��l��������2�q�ߜ"Id��ןKu)s7E��e�織x���+p��]]!���Ű����'}�h���a�M%�=��S�/�Y��Ҕ���M&W3V҉�3{�M)jP��AFxtr�>�au�@�f`��K�Ũ�_�7_��&�\�����dIm�+u����Y�_�������x�o�ض9A2��%)�&u <CG4��nEޗ���P���3S6��E�z��`,�������EB���ˇz,���t7[a����9 �dq�ݻ?*���� �,}E݁]rU�b�p_@O��MD=���ˤ���l񻻹ͤ{֛cG�B�96�c4�c��[*�x"�ӂzfQ�)��%�I�����K���V���4��wO2`�qbROك�!Z�J�:ȺCl�Ǝ����R�tΟoA�j��S6kCT;b�(tn������Im�72���[Sr�R�M���bq��v�GJЍ�C��3�4�I7A@?e);��VK�X�8^�!�qkW٘�>E�!�Oz: }�O�(qNY��h��n����a
(`H�=OQ����
����J����"<�ip�����RT�5$��"����el xnO�h�UaiS^<���D�%�m�f��܍�i��$�X��b�����y!�dJ��uŒ4��ޕ��˧�i�̘r~�z��h��4�2a��i=�bb���%vqV��0�O�!A�;��?/5y""��E�rQ�SV��y��(�iG��X�d�������\�rmOO��}�A��J��F����=�-�ت^(�q	C�9}:]h����Z���b��Z\Ӭ�ވ�K��u�Y�]���SS�(�[�?{}6�
�ֹ=2��1<3d��:c����Ĭ�J�����U߿�ԭ��=!'u!P햛�SH�ɻR?��X۫��.͙�P��!]�Zg�3�I�;���aՓo�:x���TȞ(������Y߻�B�i�"C�ce�4�4�c`�dy,� �p�$�`Y��>xYC��b⓰�%W��[����c�춱R���^�q�Ȝ%B#U�UD�����5���#,������ �?���9���r�-�QѨ�n�vyn�*���<�s�����^�:��ht�I�3�ڔ%�q�u�L�͍Z�Q����5@����<���fj�0��b�w}eC����X�Da�<�ݪ���-$D�9��5�z��lmC�JU:��&o���3MA��8S'"Q�w�t�`���a���ĉ~�E;zz�G�󪖖��&x'X��ʹܵ�l�֑pi#��%�`X�7�w�{Qկ7�z�=�"�#x�kqt	���<.A7��ا�k�A�Q��m��:%���7?�qs�1�T����<M`��d$��,3�c&%n���0oTQY}K�c��ğdHy��/��ʨ}uT���<Nt/}���!��K(�b9P��U���C�Z���AlH|b񁆆369�s��o޾Y����#�-<I��eLnwڠ]Y'q��3�PfIY�p�P����Hś��Rجq��c��� �#�6hv�1��U�m\I���Κ^�pu�Ӝ�>,����X�3�{�!�/TΆC��zf�M4E4<DGi��@&���W)_��3e��<�>I;��u��T�l�Ӟ�7D|'�uL��[�QK`喛�|\��钡&z�mg����*su�������C}󟔈�p�J��{k�D�Z�up�t2x�R�ìE�$�K2W�]BJxiY85�C�n'��Oו72�4�:�BY�^��i�-�5�� ?^�?��?s�#Y��S��9���ܭT4����]O��d��ޓeOjL��Л�(���ٛvG�$Ib�G 򨫻w摻��������73�]]����pw�\f����Yb6�	 w35UQQ�b��F� JVȔ�j[��*�Rj7v��[<��=��x;s��'~9YP������f�Bֆ��B�8Nfq�ee-\ے-���BkiE:�JD4�p��P
��̵m�%'�tД<��ZZu]JM�!� ��X>W��U��ͫ�*w���*�#+_|�܃V1]��\$�#ۗR�)t5D��le�,�=a���l=z �T��|�p_���F�Cm����]��$%�T;i2ֆ7fZm�}IVB5Xo�rl�ڔG�N�l��!���~���ӣ`=����g�p�p������s`ct�O՜r��2�u��η��c���se�����*���k�)��GBײO�jg��a�.w�v��s�-�Yꆦ�ͱ-�4<��lޜL.᯶2` �`�;�����cv�N�W%$+�Wl��Ģ��kB���ܪ}��T��AEguSI�$
*��ԩڻ$g�ͩ�T3����ИHXf9��!q�+�M0r�^^*�<^I�R�(�Pn2ۍ#|o���$	�	^�!e��0�P��f�; ��b�� N�x�w�q�U�Jj?S�/o�'�*8�Pw��m�Xa����$����$����i�M-"��pM^_�\����gW��|��8�.kÄ�!�}n�����T��^ȭv)]�g�acj�:WCa��:s��C8�!^��?~���}zW��L�T9J� ���y�6�Mn�b�]�ԖvZ�]/	
�<a�//��f�2�3��x0��a�@KNj����x���R�ʠ���7ۖ@IL�� ���߮y�q5���}�(;� _��dZ��.�֤p���_V���k��a����4���R-���e�����`�B�P�9%h5/R������t'`�()�u�ϕD��b�z͂*; ����
��أ���*�w�C�$���"Bt���gss�I�����>7%�A�F׿�Hqf�]���կVw��Q�L]�$+�63�[ن�hTu]���C� t�F� r/��z�y/��:2Ql�w^�g7���.�7HF�*���f�6���Bޘ5��Ha���kWtM���J�
N9Z�J���C�h�Z���K\-�Ji� �2�~�L&Ͱ�f����m���a5#�ԬF]�c՝=O��zY#�'O�2#�k�R�VA4���*�lq ��5;	��X�{�bU�o}������q<�� |����ӱ��R�h�R(x�������"�˻�qO?|��ғ�ܿs�� *3,&c��osBc�L�iC��)��Wր�3����A�aZ(R��E��u��j��9�tew�c}=<�<�t?����]
�.�7V@�H��˄e��v�=�n��Q�	��Rs����_C}���䲰W,��ڼq6g}��\&� e�Ud3�����jF/̀H��l�٩�k8&��J���s�]P����d �2>
F���ke���-�$68�U�ЦؤZ9��������9��,k���.*�����kp��<q(�l"�dTqmSb���Y�\��AY���̓`�����&�{.���-�ͪg�|����ԎF��\A/A4�^>'U�X�f���-�]�י}�����x�FZv���մ�(�5�{��+Gi�R51�qʹ9��9���� �
�����P����yM �]�c�������o�e���5ʲ�&W-�����$cػ��JL��Z�j�6��>�QT�)U�M!,\��p�2����_�ıyD���϶�#���	ߊ/ueO�W ]��Tȥo�誠GA \��7����vo�5�����Um	\�NemJ� ���_�=���|��-k	�b�����]�<W���&誹��?3s9����H�N9�mW���.c�C�楖�����F(����'ˌs�jQ�RD�r����C�k��Vg>��+�/�+��*>�uo�oiC?�϶�+�v��R)TyT������A��@�\���.��YVO�(3�N(��T�����J�=��@T�+���dY͈R��Vz��1t�1[���F����KyM��q=��V��W�T��v�Q5�K;�]%d��P����a�Mf�W� �<$�rYls�;�2���p�^G�>�N��o�fk���<]*EI��R'�8����E��P1Y�(ax�(�xY�ocC��#�wU�svCs���j���T]1�F��eׇ��;tt����(Mu�rn���s�'؉��*�&�������I�`�L?�3�
��1+M����w*��E���$D�Q��lú�4�K� �H�Qq�^�.~��2/�ґ#���ə�����X�[M�:7��n� Y6i�vn�	�efr�윳�Y�x&a�K��t���8$��PZ"C{�6>���}��]��D�yb�z#�	#Nnh_���������q*�ɲ �B�7z�	E����K���2�*��F3�
#AL_� 81k9�K�v[+���?7�N&�����a����Lt{���F�yWޫ��# FK@^�\���@:֡�L��N9$L��A�M�@��?e��`���ؑ<앵�����6\U��b�=lK��>\(i��n��)GF�'�OQ�R�Ҫk��Zs�_^5�|y�Ը�a0e�\�}.�w���A����/�#��ݽ����u�M8&��=�@j:��XY8��/�.��컈�OT��Ņ��W�����g+:����P���š��̓�V4P�Ĵ��:5���o'����U�;X�H��ݻn�O��5��| X�4M�`6�G��
`h���¢V�:m�L͞`u� !=
J�����e��N�m��=�7���eM�\*l��d2V�v������b��f&����q�jfL�<�Y%�����֧� Wfj����|;�õ���J�����?���j�{Rr�Y>��ù�0F ڊ^�,e�wQn�W8D�;75<>��_�x��vM)%$`e����Lg���|��#�k�=(�\�B�l\M��q�	W����ў��K�y�u�o��v�VX!YQ���:��ܦZ�����d��D��#�����iZ�}�Ɵ�ftv���-q��ȡ���o�[�c�YU��g�u��3~:I�>f�i��������$x�Y+�]�kD���_K��뮊J6_ת�a�K��2�J������+^�JN��xjKPJ5����oƃ)�q�)f�}���V�����?f�-��+C�@+��!�e3p�7�M{3��R*��њ�^�i��*�^1�t�͒yk��<1AOB7�)3wT�Ѱ�N]P�{�mr�e�Hq�^R�������O���X�ݓ4��l�4ͳʙ���`>�Ue6KE-X�"k{��H��W
�h�f2k`�AY2�C�����׻�ֻ+�:�T�D��z907���V��~o�~~wh#v\Ȫ�'7c�:�H,���ȱ]��TBm��@}:ߠH�x�un��Ɋ��6YSi荄�$��xr����܍�X��\"����3�G�ܥ�|7>gLUi��x�v�Б����ŪW������p~?o3,%0Ԛ,��gM�<ص@6�[ �C� �7��1`~�~G�Jg�	X�\��N���Vԙ�Ǒ�Zګ
��"�:�!�62��6�����T �����YdQr!W�s�	����E�S���;������z-���+����{��J��w�S��ѕݪ���[%JJ�5�n-����g���k��]J�)����ͬosm�EzHM7����$VGm_�-�$�T��n/<P�\��XXE(��������/n�C�c{�w]�B��HU�o/f���ظ�q�cF*��h�*lyl8�%��lN"�����D�����Pr�sY�/����%��󽙋��v��R���9�tU�`r�i�ќ�<! K}xp��o�^:��������S���0`L̼R�3��,�Y���L06�d[MԱQ�f[�s��c5|����g�l�o&�
s���a1gWΚ{��	�i���hK���_ه~�JJ��L���R�����L�ԭ�To�9\�R�(��c�����8̳:������S+��Zt�0�H�!���� k���u��=��֨k�N��L30�`$'?����2�� ������d�-[�~	�ے���)�?&��Z���+1q��haݯ叁4L�}7����$����\C�r��ΐ���ܵ�3R�ͺ�O?��&���g�E����ހt�[��V��m����i���_�k�������s 똡6��a|�SMĿ��^|RNv�81V�����QF�G�z̾�Vݩg�l�73�K�W���X�X3,���TO��ṫ;���Ӵ0���V@v��6�p��59����)��0�q�QB5j��zeԢ`u%)�y��:��k� NKd��3�t+�/|wN��=j�����$w�'� z X��7zr�<x��l����bLB ����8?h1A6�����٢�S����r����lH&�g���|h�0�v��w�4?���wC�K//Y�F+&X�փw�����kz��hG��

���Xu���{g�ſ��/u�L���&AY�0���Ǌwʉv@_W��ACu_��I�O���Ҳ�L�-p�����>3}D[v�9n�Gj<'�p\���(C}1�d�]۹0����+��TD��������e�Pl���fJ"bL���r�h��0;���;a��IfcO�Ƣ�xz؞����:���.�Ɏ��������l�g�c_��x�?�]�|�Wc���I��ga\)';7�NG���y�PuEx [���yq�{��gk�t��F���ݼ��I�:��I�k�����#�_d���qJ2,:ȿ}��~f�:�I����Ar7gq1{F���|4��#�\�{��S���
����矊\p�3��.��*Y�<�Xg�7��v�#i��WY��<	�r�n,YC(�A4��\3�Ҳ�uP���Edh0	\׫���#�b���I9�]o��,��X3�Q�*p>]+_l�+��w�]ۃ�oa�'9Pt�x]��VoZj%��s>���d%��믲��DҏЎ2��s"6��I$�V|t5a�M�T�=�Qn�2�g�ð��R�}/ݽX��*V��P�y���蝶c�2 �޵nT��m�;���Q���f���&\1��K�"a2u�6��ѳT'Y��R��=��!G�����K|+?N�?;��<��z)����K�5�2d8�J�))H�9+c���E4}�����I ��S׫�x��=���)b���������|�O���Aԡ�_H�8U�l/�4��x���0�0�e���P�����1���ʵ��?���U�,�7�$��g��9�P6xwV�ɱ[fw�$ie��
s������+�-2��M��t��Ρ��]Wn�2냃e�=�-m�vXK#V��R��ɲp�o����*��uW�0����(��L�e��S��?�<����`�E��Q�K�D��^Nl�j�4��4ʰ����%�~k����m��e�oqS/L��������{��*zQ�7�6V��\���J��g�'<>D}�����MW��k���g�Zj�v|nj�FMj1�p5o{���g�Y?�}��fb���}�B�J`�N�X��f�����Ev��� 뉿֎��lIܬ���J^.�uss��*F���řc����减Xf {�9�ۍ�������Aj��Z��9����;��~�!^"��gbKT:�SwRp�a	���q
#{��_\dRx?�_���,3�NA����Dǆ5�/����u������H���|��Y0�,�O���&���<��F��))��9�!=�A�=���]����R0��� �u������\�A0�����v͓��î5ڢ7������Z�.�K������=�~Cx���t���J���F;ԃ~�8]׆󆸞\$��wX���x��d�� D1��`��XPM��3��Z��v8���#1��(.Su��iWG|�Q��ҩRC�h�I��-�IW��/�\��ޥL��XGG���
�?�W{v:�K��O��x-�G�V��o����^.�l�����u��\'&Z�[m�L6ܧ*��S�c��]�Jl�M�9�V�hwU���ٰ�i�������7t�4���lj��{���&CU�^dYuLKK�~w��_*Ƒ�����٥L�'��M�v6��D
k�"<y(�kq�t�����������D�;O}
+P)]����� t����ba�Bs��,����U`�0��3�/��s04���=�_7#�X�"��ڼ�-}��a��M�w`��L/�_~�I>�)<O�g~����!�}&�T2w��=�F!��f�X�
��?m��x';�x�Q�����"��(��8�4�|l	ޞ��R�K�1(���<��t��D\t��޵ݷB��k��Jq��\�����}��;�RQ��Ww��k�8�<�&����o�X/go�V�
�^7'�OG��3Cm
���_�p�Fu?�e�&�$$�D#�C�4���&8j��a?��[-�� �v�t�����'3��@���l6(+e96���I����x&��>,�XqX�+��VV���e����i�y']Zu!d���p��Z�S�>�Q
�"�<��X�g���3�:k���ɻ��.���b�g��6�3��Q�t��]0�]@hI �E�p-���r�����MiV�I�9i�U�h1�zD���"���GM.�&O�3�dw���b����ww4�� ܳ�����V�u"|�����I� �f5��2#=q��\��=�>5�\FƇ�p�� �37Ȳ]���M���������x�����v�#�e�ˤL�}y�20F8�	��u��^�bΠD�ٲ�&bA���%6^�e���\e�]�鯩������<��T�җ�_�
bFur�%�����~���"uU�#��X��Vĭ�ays�hVۂ��t�d�|0���_��.w����E�w��'% �N*�:q�_�AO-��T��F���;�	��A�uUsK�ߍ��/l���x�p�ӟ����_~����վV���]�3�k%��L�m{���H�{~B.6�ý@S���SN_��@q�Mq0UU�����T��ˤ�=tn�6u^�6�'ׄp�Em�w�wб�:j[j��-:ޗ��zmk\t��*���|E.��3�c��w�i���v@��x�gnV:��ӽbP�p/6@�B��R��X���<�]~��9�������ֹ��Uy��X(Ͽl����3�6e���*���SƄ�b��t�o���w�/�e)1�j��(�ДO�*FMe�9�с��Yc�(`�=
�6�-(R��F��;��"���|�A�@�,Rg�O�i�uz7UɿX���F_����w��3ʭ)�Cm�-������_^>WFƃ���6�tlX�u>i"8sC��:���8������ٛ-�4w��ݪY	�\�����|��L��ޙ�W��~�87��_-�+�#o���<�/yz!����i���[�)]8�� ���]�T|�W[����WHY�졁���
&:���X�0j��Py�Z {�(����:H6`u���c4:#��w�I$d�x_"x�����T�o��s%�DqZ8{�a}w�}�-LX��\i�f�z#�w��H_gus�b�j�A�Y�����O!Ϸ?1mmA�M0ݳvj�5���s2��a�HuM��W>�&��k�@zs �[�[�E�ND��>K�����e��`���q�y�\Ɲ\��{h�O��W���x��~f`̜-�#����e�{�,qv��ij.=3�Ʃ����������Z<X:z����`˲���y������L0Fu�ZH��52w����L��?Y�X�Ќ��1��l�������5�/�tI�M'����L�B��qo��l���VN8�x <h��� �u��w�-��������n���PB���JHp����x����T�8H�:�zr�=������
��34b�V�	j�3��Liny])-�,����^���] �}���c���p��z�~C�ה��[Q���ָ�n���5�����R��` ����o�<�~!�����pSn��:|4��H-�K�j��u�**pE?o�)�y��Z�O[M�{�����	��9\T���0�:C��>N%c�I�/}�����oƠ�7�/��kEa����ochp�?ӮQ�G���.������Ͷ�#���ke��E],��b��f�'���l�4�>q�ܧF���Ha-�Sr���X;�6�f�L�q�O�N�/����pN�s�q$��_=Ut:);�=���l$m�c-Ii�(���C���-�<�{=Uy��0���Miz2ܑ�Zf�9�I(-;>��Ł!^o��"n��oNR)?�/����4VjH�Պ"c�׫n���4�����8��6���ٱpclt��__� �~ ��AWQ�&36N/�*���t���i+�>y��8y�'L�ݕ�md1e�>�2�GZy�cP&w%��؄^�ρ�F
|�q0>�Ú�R�8����N���U��Ҩ���F G�������ߥ�o��K�u�k)�'3��c�9��* ֆ�Q	of�a�0�h����ꤘ�+�k��}(P��4ݍ�P_���5Ga����gW#�[6�;������|�nf�,x��\2��$����Di��#�v���l�m��zk��"n6@����\ꌬ������H�yW`��~})�W������7��H!����b��"�XS\u�W�ǥ�'��y=�cz2ٸ�k��c����S]e8�����<3�-+����r��mdc�������:x$5�1<|@�ꤘ�X�S�ĵ�?2�S�}s���s:K->8Ny�c�
糲����uց�Nx�pҜ�W:d~�@Chb�dUS|�n�չ�ar9��k��݄��n�ʯ���N�),Ȕ 6��?~-�x��՘*4�n�K���3����d���	19�6��ަ����.����J���u�1{�������A%|�?��2PT_�}fV&��VL���[8LSQ"�ܮ�to",+���#�;�Wa�i�������{��8��G�w��U����+���Ӥ
�	{��%�F��x������.��D�
�냃���?G2�*k�1�����-@�z�WJ��Jw?�#��{�4*�n�fQ}����`�&�V�s�ҵ2�%����Q3��S㦮X���ț��/w5�"���L�����e���1ݲ=FY=:����Q��A;���%��Z��͖���G��_�dͣT��T�c��� ��;��Kw��~-ͧ��x��4��XF]ѡ|�J0�������Bc���V;ͫ1�⒝��E_��oZ�|}�=�sIԜG�C��vB�¿�J#�}w���K;\�Ԉ�O��y�ZU|h�O]u����ܙ�����N��|��߷����ݫ�<�\o4>;HDd߈B���;z�_O�2^�7��d����Vc���^1�I,�{m0N�����(�˟�K�l�R�0�AFH�{W����YhAY����M�HO��p��Z,����:|���%���IR�^g��:`���`{d{��u(����o� '��"qe��KU��%��Kl�����|y5Q~�"C�A�P�,2��L��~f����!�E�XW
��E��=JIw���6L�����_��mSfށ��K=�Sv0��[٨o�X�����#�v�Ics���ˋ�1�U��uWG�h��9��/Δ�~�:��b��n�
�r�3,�3�ȏ�Z�c�q)b|�&�v8=����MC���@������r=��.l
�E@�BK#�'��`R;�I�(K�XX�m��)�4��ɨ4�H�^t���r���y,QM�(J	��
\���,�� �^����3�x_�__�o)��,��Q������z�	M
d���ū���N���]�!?��N��������Q�"���'��u��*AG��
��!fO�dn�'��	��*�n��&�C@ȔP*���扜��V��A��w!����$"A�(��  �N�6�]W�@ F�(�.R�l��:�;���^����D��U�4�W��'r���ך����8���\M������6�����t-�J���b���:���[O"���+���^�����A���Hk׾��oS�҉~0�Q���|:qZA���N&K^�Cx�%����'OiL$��F0��d�Bn�,���/�9m�)��e���)K�i��/n��<,���J���O�}s�>J�H�N�#p�}�d�&�GjBn�8��z�)K'�e�Ց�V������?_oM̫��ص=���`Q��O[&���r�{m��x�~֚NZq��ػ<�kT��%~zd�q�.��912��()������=�TO��K��a����x�QNϮ*������տ�q:2�����6[��V	��E�MR*`�l���M���b.�γ�F��u2m�0
���k��OKl�A�F�R�����������~%M68��
-<��C��ÊǬ�Ш]ڡ�ks�A��N^���q��Jە͠��-%���n���ވG�VI��D�Z�� %xO���T�$vȲ���믿�#�4��d	1�Ɂ��Ң����(����:��i;pN�:�]�7�1.o�B��B�׾v�}�݇�Q���_��i\��6 ����6��`����H,�M2Ǉ�g�����#�2��"�uo/� �}��4a�:�l�PԠ`!�*K�}�n��1Έ � 穉PZVs
���p�5���4�U�8�z��'@޸{A���s��f>\%p}����K^���0'}le�|�����(��G�>����+�1��u�|�)G���6�bU-�
�p��O|I��n��)�e =���yRQ�d۰�ZWY	����Hu����韬.?�R�5���Rim����N� S���D#�U��P�ƥ�e�8_~�u_\!����� �H�d�@���3q�����
�����u>���l;
V�e/�@�ʵC����S���@
~�G�����|WqteM�~7b)�q\�/��2����U�����K���P�8���������p�X�n��
1I��3�=�A+k='c!�����5b��̿�"�Tl~-�4���Q&�t;�[�,���{j��v���@���ߕ?�d!�v����}.�2�k��2�.5�q�J��]#[�� ��i>�A���i!�_a��)הJ�b��l�7Մ��o)���R�|n�Tb��,@��.j����3#]��'e���jZ��z���}��md��u�a�T�����J��b���lG-�BF6�,�c�]$E	��-E�����q���c�:*g�8�S"K:X��s�o1D�@���#2Rtg nTDw�Y���><�] �|r!~j��P������w�:���B��������A��i9����33=9��q6׬�SC����@z^�u�/���-P?�Cű��.�V}WF�Ȯ<�%��A����@�������r2�k��t�c��De%���y���X���x�
N�w`�}u�������o�Q����?����O8�̀�PC�F�>�uw��2������=j��G��w&�ͧ���x�N$Q�ik?L.籞��;�bڔ�ܖX�ⅰR:J��-�׹��x�7�j�59�M6�i�oDQ�&��d�yC{�v�s�#`�-S7�qe�:�p"�W��D���s%R��_�j��E���p�����e
g��x�-
�/a�~�;������`qE������Q0���̒
�����.R��K)��k@��,r���9L��~b�s��I����P�����R�����K��2ƶ�3�p�8�g���L;S:t��$ʿ���xq��V�|��3-�cvS �Q����"��������ȉ��Ã��ޱ�����Me������{^���h�b�}�x�o����!܌�_�9apj>0��B�j�oޤx�7W4�w���L�
w7%�(Ac�܋��*˹��m�QX���
:>�t�ޟ�Q�[q��P%��=��g��5P���%��V/�^ko�,_��v�.y��7VL���<���IMd�m���&�k�C!�we_��m1S�k�'���g�z��^i���OU�����i�QL��&���Z���pG���>z�R�� 1?O^��P~�
��gdU���X�|~e��p6�'bB�IP��2)�?��h"��8%�k	i�(����<Iu�]��DAɉ��V{B�}f�S&���S�
�,z4�r �2�d��r��|׆�ٴ�r��_����BJ̕핛�ݳ������ ��A80����X"ne���^�޲�=��dD�~�ޔ:�Ƙ&��_ܡŃ��4RӤ����7b��Ͽ�S����ؒHɩAH�jy�)[މ�/x}|����ߘ�r��_������sB��y�N��M(6��D��ɴ��ަm�"�3����`��3���kq���}�=#@��δP�͖�����ֱd鮄o��� ޛF��>����r5�q�_P	�wMR�K���`~��'s�����1R~�A8d)�k���ؠ��u7��Y��t�	��66�'�
��ʰ�o��r�`K�h���v������y�����Qal��^*�jZV4$��S�լ����nݗ�|����]�P���~��{u�+\�u�-��3�t�	r�D6�����nv2^��_��P��`ꁛ�x�M�I��R�T�Jp�vS�6��!#��^0s_.hi�!���D��M+[@�G� �|��cU��U
6N:�̎M�_��(�CS�8���b�̏[`}��7P��,z}}��ݗ/�L/�T
��zy�a�,��R�	Jb��-(;-�QlZ(#Ǯ/7�s9���5�g�};L҅����?�@�L��`@$.V*��H���=�T����ȿ���/��_8�y:K�`5W�����:̈́��h�\��b��ץ�+-<N��zJ����9|PpvY��rsE��;�gB'�����'pY�u1�:C�-�ܾH_�`x�sr����@%1W��Ls�\�3�A����յ��\jU�@�C�9M( ]^��~�$�u�vW�������c���Z�����uTyL��Ca��ą8qh�{�����N�鋟]�B�8z��9'9g�K�͵/+�η�e�6bv���	��ث�Q�M�Q���,�ר{�q�6��z1�����'=2'N_u�Q�gw���C:{�] 7��2�[}��=���%ݩ��w'����@#A
J�������eL ��m�OO� =���Y�T�z/���[��e��i"wm�ApUiL�>��R<��q�l�a�<��M��n8em���;����q�����#�-E�R��~�r|�|��������3t��G�+�o_�0�'v�E��@3چH�Ye篼�T�v٧Z#x"�g�������Ϭ�d7����+�~v���8<�9��
5���8j���N���J�pf��i��?�	��\[/�t�')Y��M\�O�a3w�eأm�T��&��n�@C��yTwL.F� �V���j����k��T�ȫڶp���͇���$���=+�.t5B0۵��w~Q�΀K\F#�)��!䫛U��?�U�sk$��P���Ĳ�A�lo}�Ӯf�����7���;��v��R)%L}�E\�œ7���2��@U���NX��(*��PkuUL	��m� 8�h�La߱&��qZ�z��^��n�!��N��C����n�Zn���=�����U#����Lժ��U��4\��v�t��ה��q� ��2�
xVp����Fc�=f��P�zS�.�l��g��e�қM:��"���R�l4>kD&R�����C��2l�S���5��GvWTb�w:�^��]�7
����nK�˳����e�:I)>!k�2uЈ�>���`a�����M��0�P��6-ٵAz����_�cv��mt:v�M�Z<}���65�46��,���F67���_ .|kSX�_%��nx����,���dū�B��	\i�;n
QϤ~وK�)4'40�R�K)	���_�M�𑯅��Dq�j��R����tʚIG;�y0�}�u�O�+�@3�}w��~e���)ֽ���~�����w����Z��\�y�0�����N��9l��%�
(��Փ%X
)Ur��g�޼�uN㙔!N�� �hv�$���8�b"�������*�s��`lm��b��`���q�l�pT�A0~���ȆR�}^~⟾\�T�Q���4�@��&e�������D��Y���\7�u^�͗�A����+�HP��EY�n7<����En;K��efh�eQ�nf��l?3�xsH���K�*�3��+�6Ov����]Y�,�ss�~{/h�����l����d���s��<���-P v@Ɯ������ �kf&n ͞]D�/�a������'X!9�Ek��-^K(gG�Ƌy1�ܽ� �@6�)�z!.\��6�c]k�t���*�H�u��R��,�V���`���G�t��c��-Y��撁��+#&{.�x���d��\�Xv/Ǘ�w�2:��|:�+���Zi:�#[��(��[��k0c���v}6�([I_�s��i}��/&�"�=�|��dl��yї�-,�&S��e�T���Ԥ1���m U�X�B+�F�����x�����Y���"��a$f�N7��J��E�)�e�I���H�I������4Ը:oA0Z�P���3/]��K���~'���@�LP ���
�	��H�m�NlW<[?W�P���m�����,-#�٨��`b�{e"{�M��=��)�˫4���!*�B�}��2�q�nvrӽv���*�CT̏��)#e�	��C6m�,a��&�L��u��(lr�ؐp�3�"���f<�x�ceW71�|�{�b��?�t*�k�X(n�:�"�?8 R�u�����<�����/�Zۍ@��^���y���ێ�!�xTAk���µ�����MwN��sH�iPV}�=�a���ܰہU��*`�J�F�}Wa����M�rF�ᓢDJ�SL��N��o�x��p�e9� `���c�1�l�������R�7��@���w���{�\^b�������F%1�:؍�y�I!�ry���N&�&��1rP-��fX�@����@d��tR��3��p?0kC<�f�&3J�D��X�}�]�-덇�x8q�b�"�I
HT"_��C� ?��z�<�_��Y���q�#�}^��	�}}7�6�՛����昺�ť���@��3���Y�����zD\��m�H;������5��<
��z��>֬c��&Sp��B�ƙ�����ͫ�нR:���ᰄY��5�m��0���ck3T8�n~�����{R�ah�AM��-���C!}x��
�(K���{�RjC���X�!����^���zt���GCU<���A�@��X�Gi7sV+I\%౽� �5��kyD2my���G��Wke�,9��Z������vϣ��|�˰[��f�
Gޯ�7ӓn��b����}�H��]��� ��I�H������܀���_�|�aA�p�D�q�Mz���&\n̓��B���eX|S���V�z�t7�f�I�5Màϧ�t�b��M���C��/��CU!�wȒ֚����vR������W/�����@��-��H���:ƫ&r2_o�7�q>�R���b³T�|�#��֎di�����R�{��U�R�p����d��tb�����y}\M���c�&��󼡰Q}jU�k���xr��l����3����^�D�8�S�0/�Ц�`��e�n�b��~��rQa�����P!�o� ���bX�0����!FnG�>�D��z��ǒ�0Qfy�ŷ�������O.WS�p0�ƚ��6B�%}�g�a����t�PTOH�[�ڸI�ƥFq�����̓!f��`���񺧳�2�*�>���j��|�t��ܬ}������e�u���3��SK�#Ҩk̥���E�7ͦl��+�Ԕ�� �͕�8�}��:mq��#�����⩳�F�y������SE�=��[�̦�����@ ��1�/��D�����Ӷ��9�S�u�Au�|2��i�X���$�1�M����&�K�~�woN��c�������o�/u��(<M�K��q<Y+���r	.~vz�*d\ۮ.g:�#D`�@s�4S	*���T^K�]+��%
����V���/�ŝ�⍮�Z�8v����C��s�I""a�K^�>X���_������\�T&��I��V>��Xz� Yq�Sޥ�,�S68�>&X���N�#'w�ϕ2U��3���� s1G�f�u����j�p�հ�����}�&u`/�^�_NVC�P:�Bx�����h��1L ��]C�e�oゖH� �x�3� l��V�I||�>�z�[*��nh�A�AVN���ҴhT6��8��*x���+��a�r6�vL���h�i���7��n�#1�>}�?F������T;W�3����O��KM����Aʕ�)\g6:q�C�^�B^k�d���lj�'Ns��E��AJ�d��9v6[,;�$>�R""�;M�Lu��dů�<O\K�zAc!�DF�E�M>�Ub�����I���WMA���LgX�o
��LG7qn�C��e6d�e/��W�N.����U������
�g�߳�:x�N+M�|�k_9�����5�l>�|���[���SS/�2a�g]�X����ϞL<t��f��?�1�C��C�"�Q[jCZ�<"4k�W�[5|��Q!�~�T���*��4�����p:���:�">�w�޶m�
����U^0��u���z%������̭F��g�㞢TD�t��H�7�FP��hhTά��`V�����$>5Ϧ�I�ppj��4��z�Ϧ\�!��͕G��hyOk�;����0s�>���X��Mi�cD}�#l�_y�lj�sx���j+'o���D�(h�m��k�<&������p뢶��2��~V�y��F��9ܖ�?|t��f�*���bA"������[M��)�:9�,���;X=`v�n�˥��a$, <������⫛)�7��ȃi�ś{���*��Sv�XiS"߯U�*���]�q��Iq���r�s��J&�_��Va�A}�olNN�s�������;1_���L̙�>��_�����~E��x����9�C��o���%�Wg~b��MƱ���)#�iv�����첓(��K�bVs47V��^�q	���.Kq��>|���[�X�4Q`F��M��tXw����q���jE��2�s�p�J)Q�=���%6��-+��������'��]���?����%� ����y0�������o�+�G�2q��?X�4:	3�+�Gуo��KZ!�^���Y4�:L{&6k�cխv�I)��>n�oBg�Vw��m ��+ѹ��ͬ������FE�A�o2���Cqd/Q�>��H��*P%~�����O_�m	3�� n�>UA���� Xvvr�?�F?Y�Iֱ"ccS��t2ɷi�1�"FD�8�l�v)˩QfX�Zo�J����ѯ�����vs�H�����&��|��5l�?wIPO��8ؠO��x~d8_=�q��#��F���B���x���\���]�w�쀠�b�qf��O+�<!3����8
)Lt�7�0ZXe�<Hj�ԷH�3�����6���L�c�>d�y�>��I�r��\���AM��`��j)�c��0��bq���Im&�h��~������#����}���{LVlSsb�� ��\�m���5����<��R��`�- "�'q�U�K���$:D�c���p\��J�K'��_��_�P�ۿ�+?�vx�6SS�B�I�+���ĺ���~�u���d�2>��;�-NL��1/�_�?��:wc9�&������7wy���_�e�� "b�T�hn�l�q8b1>Äu(��2���}�?0�b�����d�asKmG|���T�� Y�tg~��ؗ��4Â��!
;ڱ�t.w�kc,��F	�$��Ju��uI�Z�,5�j�t� �F����W׻*U�k�;_�S��tu�5xD~N���L�`ۇoŋ���]*��RT��I�f�Y:�P��/[ �Z<��8�:k~ܘ2F�]��u���ɫ�v_�;P����R��ܽ��'s�_�἖p>{�KӇ|�>����'�׋�6��]}������7�"�F�5�22�qG`ӓ����.�4\u=�A��ڎ���@$e���++�4X�bSÆ�˟�ˠr}fy��uR�"?�􋼙�p�͖�3lCh�J�/�ٚ�f2�+��OR��_h�n� �oO߫����hG�'���fó�q�c��Ï?2���˿����X���ȥ%1����owilA=�G���/���֪k?Ն����I�Ib�h��O��߼��v�����H]���yc�n�Ӎ[ �->�.|��^�z��=�Z{:��3)��(+�����D|�(��+D����'�c��_-t2�j�� ~R�y+Ǯۆ ߭�@s���~	�mB`�){�xc
�ݜ�GԺg�$E�fJ*�\�$�E�D�(=�<�\�W
�`���9u�w[�����x/�W\"��Û\�*X]�.U����PR�hf�0(m�w�i��ͫ�X�����m����������J�NO!t�,|+[��)��9�����=����^�u�kt�NƱ���>Y\�	��&EUO*�P��S��l��
�A�C>�5�L��� ���\͓T�ū�j8�w�1��n8`A۟#Ix��o��2SBsi�T���>C/d��Ǟ��p�H[���Spq�}�]�>Ø��7[f� B���{���*\!c�]�Pf����5E�e��׻&�"L�)�+5	�j?�� ��O<Jbڸ����3b�:��U�`��ާ]�V��)Ş�W��j��=�KR7[Ì���%K���5�?u])m��}�޴�ޘ�0`�bܩ�'�v��"<K��RJ��Sj��^f��àE��)?��;	7�n�We'wz�?9k�ƣ��Ǒڥl�1���E�F�&:Y�2.�Ƞ<�;���3tw)n�����9�_�1k�/+G��|��;���:	LO���#�[�O����J�I��ڶ�m��8F��Z��YpUl�N2^�M����c�M�y�wlNj��F�y�-���d��13,��O��	GdBPw?nY%2�m3�c�`�ejU_�����~|B%���<�~bP����`���9�j�ƹvg����Ayג�a�[uv�ԥ��Y��3\5cN��`�o��]�!r�v��)_1�;M�]5�ò_���l��b����8�z3����b���&�M4�Dy+���-����Llbw^{�x����S���v�!������\�-Pa/�w`�H����\zޱ�/`t������t��ζ��${���n=<=�_��33n�@��~�~w���!�ö7�z�l���,η4�Xt�OAU3�c���D��O|�W�����P��d�]Wꁮq�H�BUV<v�4���Z�<9��H1-a4�y�O�N�R���9r|p�"�~>J�^_��t��;��q���R~����]y,��㲝�0�Cq�����v�x�l�Rfa����g���_[�Cj��Wj7�;\��Tʫ��N�X.nH�9�7Սn�`��Ձ��&3,x8�(������/�y8�KU��c͖��.�"R�,��m��(��X�=Q �/T��+�8����m�˭gPE�,���;~_�������>��{�9�b�B:Yٗ��������Gn�����O΢���L�`��P�rJ����
<����L��̩�x���ޏ���M��ܤ
z�G�ͅu���;O�
8sⵝi���+���
��>Ax[t=��H/����0���t�;�HlP����̴pH_�{�2�sM@�蠐͖��^U����=&�\��~��O�iYp0#���N�S�:�;�n��"�k��gLUa��� 
ϳ-"�=l���?�"�ʠu�zy���H�q�u <<�y}���7mkH
^{����80�QԵ��1n}�C��A�&�v{fО���b�}i@��N�{�~Hy.X���y��������w��&�� uv����|��C�8
������E_]*0����tw��ϓ�$�>Z���)�2d�7�}�s��U�/�����D��x���_I�|w�}H%�`F8Cs͡�J;vX��\���D�p��Nd/����޳n*�#��8	���L$����Ҋ%`���}aɉ��0��~"���,.�e><������
3 ���@���T��7�xxdjG@�0����6���>MņE��ּ#�� �O�	-'�;A�%�El�m�4gW$ڬ@ g�	�����o�+��+��sTy���8��J����<�x�Q%=z�������^�o�$�7Ԉ�atƟ �Q��2�1����$%��� �"ZU߂gۙ~F>��px���.�Pa
H��SρQ��%jO���N�F;��0^��6�pe��B����Kc��o`����5��`��GN�/���N!��.T��k#&��c�.��J���#�"�_�\3�t�������q�,`-�8��ũ�E7g2e�7" g����?����,�UvEv�]��&�g�4˄�	���-�����fѺ�$)?<ý�7'�W�V�Yj�⏦W0;?���|FgW���T|�G���6~S��ɺ_ ��.mZ��㺊�}I�Je�N���~)�2�ژV�����f��l�-͡�Z�g�)QL����r��B�Ɵ!p��P8"Y*��j[����Ar��Zù�Y	3yt�7Բ�g��&�lg7P�fݛəd2��o��<��������A��]/|�:��� ��p�QE���{�%`
��<HyhR
��(��wσ��Gv�3%��!�]�.)�f�
��!M�YW=�8�q�<մ�(���Jp���&�vnU�Mp^��ݺ��23F�ٸ����,�c�-���ƤٕY�{�X�;k�Koa�������@��6f��O	@]=���˷����)����`�2�eY�/��z�l��X�0��	i��F�hp���^��쁪v��Q��Ʊ\��hτᔇJ.�a�)S���)�g���g8@�\�uo���b �R�����ukJ�n�) l����_��M��T��T\f(��s��,�ۼsF��ܾ6l�wyn���K��I�J.6_4y�`*��2E���>n�BL/�,;H�;��b�e��?�䡇�S�뻲���04(��v��y ��<g�y��V�PP��+�Xwq啃j1͏�-C_I��<���櫍��h=`�\�K=�r�f=���&��GWrً��|ئ��CmY��y��>�~&�β���=����6$P��"�#h(��xp���>y�M�i�
��7ʛ3X3kHF�X�Zik�f������U��vBQ�y6ѦY��y<]���2�R�}�M��Y�i�:X�M�{o��o�f��(��xg,K�'c}c;Y���+Vɛ�@��Pyv�f��C������I�����7��rA|��0� ��@!�S��:�l�����1�6�L���7�,U�4��m���Ԫ�*�q�D��ݱ�F����q&�B\6e���pi�t�Cv�&��!�؝Ovf�d*(W�D!OBE�\�J-���H���ښ��ڔ`g�Ŷכa�W��.:]�f$��yV>?m���x?n��[�iF=J��#��뾽�'�m�����(;���Y%�z�;�>�Z�p֕�ԍZwI*�Y%�/�h�d��(���@WX��wQ��4�Nk�|��z��'ixĳ����u�\M}��i�i��}<5�3|����l��|'!�p�F4����Z��"B+qϲ�	���DK^&���PM�^fB���Ì�MH�g���H{��/�V{���Q�����Atט��h��u���[vJ3H��ĉ��S4��xS6�ѸL�d��D�S�̞��x��MK��;��R�&���x}i'hW�d��o�`�.����	T@������� 9�^T���b���q��kཡ���JÙ5��F��P����k!�CX�����ҩ�J>�<�nW7]n�����)�}�2İ:#��P����Wu.g��$�6��9��>,����0SU,��1�S����_�q��r�Ag(��O ��ֵ�C��e�|����`�1I����*=M�v�k�C����J����ƾZ�>ȁ�{7w���A����n�L�kȬ������揶+a��Vq]DZ"S�`D�c��y=�z�>E��l}V��:�?]ūU��k�%a"�I�e�恃�9WM��k���$ל9��J�P.ŰY�=M����ap�v � ��Ե��.h�Q���v�u�Vǁd�f5��h�d��xN��j��`�I�e���)��������ʰe���Q�&�@�((f�>�l��%�Hz�~}	�~�HX�x���e��\��]zrଈ�2J�^�c¤P����q���I���Rx�������"r�����ط��Nl��
 �jz��`�����Uz(\q��{�����T��Jf�]�����ܥg�@
��f㽸`����0�����;�"c�F:��[m�f�H���`O-��8H��Au�����3;�2�^+���4)[kFaFJ�ZJ@���������Z+v����y���z&/�����$/�Gf���z����q/�>�v�v�2WJa:�U� �p�+���8���,����ڸ3;�d�Ս���?:	�1�az��`�w*��>M5I�g	�����Ǐ<��Hb��s�O�c�1F����FBw�/�:����pk6��ܡ�Sj��>���-,�o�8�Ǌ��V*�sϦnלI6:��7e�#�&1�C�vIX�J]>gG T�7��i��D��7�2��Ycݸ}�Y���վ�
�s|oj0�FJUQ"�|���DGm09v>p�j5U�i��=Uӷ�˒l2y(q����د�'}f�!>�Ƙ�������tP�O��1�E!N\�]�Z��j�bC�;���Ql �e����en�����oϠ����չm��٨,�o�0M�k���}�Dϵ�~�5V��0�a�Ƨ;¶l�����~X��2xť�~2���7MMt-С��5�p���j��L�gZ��G�z��3�󶻻#��N���t������G=1��3�<���w�꣉wH��ٽD߂@�v�&�=.���{�h����Բo<�jF�%0q b�I�M_x��4�[�����Up_k��K���?�r��jW�����_�M���,{��P������oF�y��� �ՕO��=���Ѹ�;��o1Oƍ5n!;��?���tLCQH��:��(���29��Ep �����(��#5�����7�Yh�k��p%p�N���.+m���|̨X(�4�	ZK4%}��t����?��792k�>�å^3�N1�xQ���<�g:��!�d��B;�,��K@��7�+R��c짛;e����s-��a)�,��7��N�+㓭1֔��l�e�[�D&�2���y0�p?�f�%������ژ��,Q�᠁��Ws#�N|{;�U�w�)3�mY.�����Q\^��v�W���G)����V�PS5�OSWKmD�z�X(��tiUÕk�7\��3���J[B̮ջ��:��M���&l�t�]���9M�V����Yw�(a>��C���b;`��Y�m?�A�C�
�;���5�Ρ���>{��z7Z��Q�#�c��6�����=>-o����Þ���� �承���"Cw2Tz�܏e:M,7ɖ-&X3�A�i����S�\И��[�v�J��9x��d��)�Rk�c�c�swA/�ucF�Z�3k9Z?�f��0Zj��l�ɾB<��R�ڞ�q�@q#!�q�M���A�H����M#O��)3Vԩ��k\'o�Z��u���/m�a� F?=Jq��f�ʨ���m`y��*�_�s�\�4#�8%gDsqk������(�ǡ���R) EÊT�Z"�6�!A�gG���Z�3B`^J���+]*>�ϣ����b�c��M�"v�]��d�(��	q3eC{H���T��^��\$��Za����PY�HP�{mf��PX���h� ܗ��⦨�}v�V�c6����� �a�j��J	�[쑗�����Ҙ�^UU��J��.1R`E
�|�����C�q�%*t�b)�K�l�Y80�u�dS$+��+�	�Xc��QK�#_�hC�`���P�]��v���k2����Hs3�-��t���q@�4��f�y�H�lu�U=�[��
��(|�4lPث��Q7��%��0Հ*W��MY�.��v[����,2����4�5� 9���JJ���KiM���٣6�"ST�cv2�����`��4uᢽ^�8������?VL�U]�8jx������L��U����])q����q��۶Ŋ�~�[��p>��O[i�$�e����:�q�d���]l9���Z1-q>��������/�c� /i����˼f�ֶ��ut�)ϚW��g�h$m�W7I���16&Qr�cѪ�z(�ĕB��.1㛛/Θ��[�l���Y�&�G'��Mi����>/T���I7�wj��Ln����X���F^���qۗ��"�K]Cԛ��k��z5\���%>#�ĕ�@�?lz�De�tlJpL�HW7�?S��ӛDN�p��P)����kb��\qiʾ�qe�˛N�Z�����O���H�F�`�;J��_<m���ғ�[�,�#����J��	�\8R�K
-0^��mR��N�(��V��hl\Es��`�%�X��
��I��؈��h���J�Ֆ�������;�>Y(燥�oj)���m���F�(�f���7�@��H�� ���\!���FA*M��ĎA/���B<����:�.��K)Aa���p��TQ?HE}�[�ƌt;x�- ��������ޒok����1��>��tw@%>���Q��V�db�V�(�nܶqZ05i1���v��4��v�H��G|��ZaFxO�߂�ӻG�;�o��7�
��؟ �\=f�{X�%�*�_c�J��hm��r2��p ��2k�γ������B!��Z�b �Ǚ�$Ě)7y���:���x��(��;�NI�����e�'�`h��U��.�6��@�
Y�(A��ˊ��52�]��L2鸴�\��e�f�-����������O�<Y�@\�6F���D�٧�FEO��� H��v�3�Ȍ�D�㖑��IڱM	��!�*L)����8��4��LQB�V���ɢ�Ň���6��f�k����mŅG�M�yn��բ,��]}��$��a�_����~����N#������Wwt�T¾�������z��-�V��u<�*��/�~/����e��3��#R�9����~�:f~��� ����Hl�e�4,L �L�[����[�Z��o]FM�����`0_Լ�&��@��6���>�ֆe������6�V#E�7����H&�G�%ّ�@��������^���`U��s�s�ք������*�q��U;ƚ���(D�_^����+	�rc��'��r^*<�DTy88�@w��J �b���>�b�&����ul�2�ci�/#_#���ۋ���Y�ʬ7M:	W��D�Mu��|;ҾP/ .�����k5��o!V��s���W�)	c���?H+�� �{N��1c�O�`^
"{B�8KOQt�fO��ˏ?��e[9zF�HL�*�fj��"��jA�?~�/�����5_o"	��{7�H�򔱣��UV�&�+h( �\����ߡN�F�k��W�wS�z�4��vn��-t�����6�a7D��	)�'똲���2��J���H�E���h=>l9S��7�O<�y��TX��d}��5�M�.#�:4��1w�y|.�*!`uc�&I'Y�e�Yvv�+�+�'���//�<AJ(����>���	�D�����?���b=�d���������l�����J�@�5�Ġ�sp�����u��A�V,g1	�������]>R�ִ9�Sq��:�Y֚]���^��/^S�{`�A��������9R��u��O��������C}��G7������)�Qdb10	��L^9{@��2��e3>?��p�}�OSRd��{��K��:�ݦ��@�+����>Wa7�Z0-j,v-����4�����5�5�l�"R��7k}��DP�2�C�A�%.r8Q�s��l��J�����- �mlwϘ�M�u�Jp�rz6܊)�ѣh�(���v&�_ܘ���l�S�(J�8%�j��nڌ-e}��ف�&%��I�`�ؗ�Uk��P��3���I��P������� ,��[��]bhףJ��vX�X|X�q$͂�������G�Z=�"��Q����]J��-�L~��\}�WW�Φ��q��d��?W7�}ȺA��wV5�K��^T�@4I����Œ��j���d�{��E_�����M�P��F9�L'������Ⲽ9��@zoͬ��5#--S;�g��i�����E����	'���C���~}u� ��0`D��Vb�耱+�~�q_GTs
�_`alR:ǚ6�O������Bg�K��)a��!7��#�{��[��w\�_����W!4�j�-}�Zv�=�)ȷM$�Y1��A��^��{2ֲ;��Ƭ�O��k-�Ӏ�-P�L:�k��h��IXq�)p>��R��� 0R=�JF�ũ��u?��Z�C(/� �r�{��^C���� �5�K|t�W�&o�縴F�G�R��5����u�E��+E@0���^a:�<k%�<�8�L`0[v�r�>��/��
9J�K�&�M�d_�T4��7�]%pH�RR|�I�7f��J,��:Ү�I��
�;nWu��yv�|�%�1��/���W�Qg�eo��0D�Rez);1K�%X,c+K�$�eԳ~:<0�Q�	�˶9����<]��6��ٝ�4㣀OT"���T�R�h�ŌDM���q��@f�?�mD�a����+�L��b Ȍ��^��Xb�=z�cs]X�$����>�Z�*=��Y�n5Mn��+�O��Zc���[�
(���T)����ҾI�V�LO�z�3ۂܮ�,�{�Mi����p���O5~���)؜�Q��o�Ӑ����i�1�H9�r@�%JD&pjqn�l�J,s��#�͑ԣ7I�F�)�'O�W�Ndc����l���$�zq@L�xm|Ԕ]��)��X)�p)�r�9�Be�J��x a��J�n���τ��(�yv7V������'@5r�Q�~1w]��b�K��(�a׺�{�﵅�p�����l�4-#�,Vp���p�ƃ5�q�s���V~�;��s��~�3��zN-�(� �<6�8�Q�B�� �UӍ]'s�0X�g�(��h�ㆉ�����k}�gԋm��\;>~�ڕ�6
ތ-8e=������9/�|�רӘ4�������qY��������l�6�z���} ����-�Ë5��ɖ�iu�Ѹ���A1�gC8����vϣ����\b�����s�h��{U��UY�Bs�؜]����5�N�5�0����{=���X~�Q����~��v�`ޕ=ސ���s�Z���і"S.��,�A�S\��q��x�]E�EWn<�C���w�UZ$��1����o�Ի2-4_�3  �o��fg��=W���%i
aaH���'��L'	'�9XU�O&�Y���t�t�M&^�x���W黳����χ�w�s^Ԑ���7N|��cĳ��k��,�/���S�U�:�6�*Ӛk��䮙y0qRjP
*SG9�C�� ;h� �YA�5���i٦�T�\v����c-��,������B��`U"ken�j�
�L6U�P�H?������A%(_'��t;Rz|�䀺�w�ٺ�Gn�B��ų��y�����G�IoT��W5����,����u�i��6�i���=�������,�/�%ؔ�x�On�.�@38?=�~�7�`
�e]�v+5k_�;�T �Xʩ��t�hL��Li��~l:�vG\h�_NW!���=R0K��m�&�`)�:J�	�Y�$��ђ���}����T�^\������,���L>�nwp�(�t�������b��=��r�Zi�Jԑ°d�t�x6Q7'�Ͼ�ť˙�t!6.�{�Nz�O*a!<��n���2���~1�q�ϟ?��>Y�\*7y�^�i+\�?��~��°���zBX��)%A��jY�&�q��V!#�'�d>H��7!z�?�2�v訂^���h��d�ir�	^��r@�iN�	�RQ�Nѱ{�\�(�M�N�Y]�KQ+�z��K{�����Y�9�u�Cpe���z���^��n�]D˱F��2]i�����r{�H.~��8��,�����oAs�:3<�#&�`-~e���q��(�]j��a!��U?:+�%2�D�A9�Aj�&�����3��#�j�����@�� ����2j~>>�ii>�b��¹�
�Zzѭ��#ˏ�'>�1��^�{�EĽ�g:cm�u�Ī�n���m��-߬6�Y'�q�>*i��uܠ��t��7Ѯ��$��T�����.��{W����Y�D��qGv������NZ����F�eyA�U� �%�ɲ����0�ə^��0*�Wn�K����/m��ȑMU���gfw����a{����v���d>���7�jW��T*�y �@ ���#��1���3��<)`-�3U���_����V�������޿|A)*��us��c��QU35�G-<��^��1,U޶3�͹�����+�Ed�7�0�aHc؏.�=�l(�����JH ��qR���CM�4^�m�m��m����~�����?�I�)��F�ʽ���ȸ��3�[kk��v��̂�9��A��H`�R�l�gޏ"��]��y�ρ��LD-�����X[�j�ٍ���'_�!EJ�؍Iy�P޲����ʵg�wo�Z�l8����u���^��٘�:!��y��r�i���֟�<t�g�����V�KA'������6�2�G��K��<Q%Wm�}ޟ�x�ϻ�~�=w�$)7[���I�%Ze�}��Zd�C#��g��Q����C�!B������0���X=(h��Ҩ�V�"�Zuk��$®�)嘭�'��Ʌ�X��<Aq3���?��,u��)�Yg�vnj�v#�	!��x}��X4�Zyb���Bzy��^�S.<��BY1`�߿b#Fk�ی�ׯ�^��:�b}������{�����z&}��&}R��0�4(e#�5Ee�p@�����V�S�n��d�;�[��dي
c����ۯ�q����/���`"�����EB>ѓ?/k�*U���z���i
�ڙ|Y_)X<*T4H����`\.Y�4���S�,4wJ�g(y���SW���Qĸo1�0����}�^;54y��s��� @����&wO�4'�;���E�<c�*C�qq&V�е�������(���&��3#�����rm���d�`�j="9�vD>6�r�M/A]�Np��cܗڔxa����t��]n*� �+���["�Lt�X<?a�iB��C��Rق�d��MiW���?7��} v�
U����� ��q��d�j,([����C��K�PpU�@��W��B4�ͬ��f� ������}%�z�|co�%�-7w�3�����z�)|#���z%��{ŏ��n~�W>�*��Ȁ״9��[��%k�i���a<%�熀I�r����Kp�p"�y�:=*h��d�oKg�w9-̻g���ˎ��lz��s���l��fHW�\n��?�؍�o~���w#���?��)n���n�-O�:uyn,v���NؚtU!
>6����`p�ޗ����2�N���!:����(�=����,<�=+��yzF1�uw�}=��٘S�_�pftn7D�T�[Iv��v{�Oj�U�����ɤ�����0�1i�g��G	�W/,�!�|�M�lݛ����{�a؞q�qw�����m�#�vW������r��Wt�Z���¢�*��ȁ?��OQ��a�k(������Rr�����|��ND�3�����Ϫ������T�Y%�RHr�`��-��ƃ�����`Fˆ��%��	$��i96� �`|bA�g�fD W8�4�$���{d�'��΅�'b�k��b�U����[kX��,+��-6��������Ðz�Ӱ�siA�N�����e�� zf&��ؿ 3Z�`(
N�T��m�1mL��Bt_dY��6��ǁ}^�g�1q!��F��0o�Hq������/|v��2���+�ӈI�(��5P�j������yp��=C��qſ��Ĥ����G���7:t�%�`�9�x��.h�q��>�*�Р0'4b`� ��#*!�%y�77^7
4;�v��<X�h<��C1��gJ�|s��8s��r�>����G�ucJ`7F��AC���Ǻ\�h�>Q|�p�F���=i���m_��?w�P�E�h����W5:��0�4e�Y�v7F6�E��'����SM&�ϼ�0��^�ǅz��	;��-�Wȑ�'�I���Z.��� �wt眨`�����f������޽}j������mC_�>�}p-����N=县��;5�e���As���$����v�$�����UF�����*UZ�B5�7.y�+5@����,��,.E �I��ps�G�έ#7��.��mv���a�ipq������BݟWX���!fщ�N8P�Ѡ���c�i�>���>��������� ��o�����?���*�����G����'�왑,�ah}�m�Xh7����{dF�?C��@����:���D²��D��y�=�L6�g���V��ye��w����X�}��#L7o��4���+�����6�N�za�ݕb7sp6��Le�7>����)[}�[o�-�W*M��`��{��
�����<B0G����a�r>N���#��ןC&���e�3��-�,l_��ܸ�u�Jο^ d��Φ����b�׏�(���^������m�21�I�98-T0T��߰�:�$���7:~gH3�υ_hQJH�Ӭ�NU�X��%�m�ZӐ�f����&pdIW���-|��1#:y��7��t��[�(��B�ejx瞱y9nH������n�vb��6�������Y�+ۥ�@��9q���4�>����|�	|,�7�7�lV�Qy
��V�f|�_�O�|�M[_�d!+��I��ֿ2����+�k�)��i5
�%�i�H�B��p��<Sn��&��{cڴ>���}@�fgb��@��B�H���z+yR���cK	i�/�W���%ʐO��{��3�6^f������s���F���!��P��3�K�Y��8#�	1x��/��=Cq��&=����P��C�(B#�EW��
f6�vc�A�����9f�S��ʂ�l}�<��ȺXٵ����9����Ma�o��
ÃPO�u��!eg	�}"�Ƣ�;N�	!%h_�
8�<���̲a�+�|���Ys<l-���dZ{�8���m�M�Ġ�F�Ml��ATы��w��-������%�W���e�ģk�}z��C�M{�a8÷�J&P�#=�"ch���Ic1L0�x!��O}#����/ho��:�(&��H�)js	#J���/��ed!r<9^��"\�:k���>�6��D��]�O�-�g��q:m�R`}��gv1��� C�N�A�oj�n�Z�B ޥ���Y}$嬌o���ɕ� �c2w×���R�*�U^��/��nՐ��*#�<�N^���<:MI��8'���o�~{�[��������ް��ܓ���s:�c7`��C�	������+��|����sҘ�H։�kt1Z)f8�pb[/5~|����u����*���[`~�4��=� �y��mjWf�}�X����B��4Ҵa'|p���M�"�1���S���9)7�I|��F���^R�x���"����5�����W�Y��>��=���p�z@������u_�����i��,#5
f�=�����߽Ay���O�}t�u�ߛ���P4iM��<Fg
S�
�����e��oN�{y�*���h�H[Q�o%��[Ң��)0�!3���FR�V6��K�����-�����Ҭ�-�'VmL���ې!��yz��1]�	�}oh�<ٗ3w�����4��S�� ��ܫ5��pƆ�#3���0X8�������%m�	$d�آ���@�uԈ��3��к���T��N�f��ȞV�9��Y��ɍ�Qm`栭}`��A��q��!��3��=�Ep'���&P��>3�w��O�O�G��G��[��po!���p6nf�:Y���0���T�4d����޿{�m��c��û}�~�:���.�
Z�׺�:�u�9�k�q8Y�0[�&h���(�ܰ^�Y�P(a$v[^%7q̣��Ek!�����vO<I>�	E��ѷul��%j��9�������.D��6&���!Ltu�)2��Ǐ����}��}H�gWQ	Rgqʣ����>�ٲ���`����޿������޹�C���ݾ�9�\2Ac�i�x:E��Cx��7y���<���P̎/%gz3J���T��0Q�D'����%7;�wѵ`J�,�D��k��p�<�"��q7�9�aj�_Yx��$O�ps�s���a�RGy�g�%g���28�<���2�O����.�lz�o�B�"�T�缩F8�Gц�33j;d�����{��#ՂΩ�/L�� ����I�U	@�,�C-:�y�L��ϖ����y�D\zεt���۔<�#ܱ��ƭ�zg0P	;����^��p�F�vQ���:�ujFTl$8�"�k�pgE3n|m-M�o֟~��x]m���\�9�\}�0al̀{����%6ͧ&�^�T`c7�� j�[�����
��6Cݷ7$��&�8{c�{v�>�����j�ɓE#X%��^�qA�G?`m�^/�<q�90��mt�h4�N�ʪ�-N�X�9���t������NH��8�NT����c z�Q������Ă8�_�'����_=�����E��
*�4���5g�
(xݓ��T��^H�H	By���aP��h�Z�lG�Ոv����L�!�X=˩���t��5�l�h�����?�*�Dv����{�`xRo�-Ly����4p7��Ƶ�t�Q��ۂ�3:�jA����}�Ήu��s���I�=E��|�/�2hG�N�+�/Gf����
[]���@g��-�9{xk�=< �r����o]s��i�yb:`{ �m�Ĝ��\<�(�I���H��0������p�qlA1:o3�3�X+bDR0B�����I�w���0��Ȍ��Ó{aKp��;U��%���(����D�WEж7�HY`"������ZԿ&b#�>��)�-�2ڞ8gxui�y~`}�l1#T��^��^u����������0B�.7jFG|���G4���sim�}-�ky�=pR�i{�7��J�#��߯�؈��H��$��A8`�ܡ?�H��DoU	#D�b���[���@~��J ���e7�����g�Kpv^$�ɦʢ)V4�c������z���+��+y�n(Ƽ
:}�7����yF�v-��=B�����;�n���p�ݛ���π?4e��C#{ 8i1���:�i��c��#Q��M{=dq�@�[�&(N|�`a"w����96�NՑ��#[A?==��2#j���M�~�U�J*US�ΐ���x���T���\^pY	|Y	��xr�2���9��;��:GP[��� �-~{�'bkW����VϬ��L�������p��`%D־$�(Z3�s>�x��,�̵yТt�+��[c� r���Kx�H>9V�V*E��d���ب}c"�%J��|��y)X�r=Z2��?;����zW�[�]������ G�R�ݐ���{�0#z��0FҦ�x�)�*x�5�:���]�-q_a�g� #�d�p�hl�e!5��P��6%�i��4y��{���σ�#w(ͬ�Z���DuG�����<M��Qc{#�H2�SdWiw��a!�����l��ϤQ<PՈ��S��{��É!C�M_���0t��鑊� oQ�BKCz˲V0�2��L���	�V'?� F2G�8Hԗ��<�d�E��C43|� \0��Jm�:�[CM%#�dU τ7,����)��MyI�����j�Zq��mSgʱ��m��w�W5A��mK����:��ptA�Ul�k�]Fo���H:i92�'��(���>Oy��M�T�s���q�+��`�<x��@��IQ*;�<��!�!�v�i$���z�᧤�I�F[='�
���u(���9�������M���'g����̻g�-�o��x��"6�$�^[�L�	����g 6��+�������o�����^���eY�V�]"*�i�=�C���x_$�r��ॗ�h�ύH�#��K�b���3�b4<#�u.f�N�uh"i��D���mH�^�@�y����=d`=zΣ}	*�.厪�=��@'�2�ټk
�����]p�N�4Sx7G�8Wax��I�q���V�U��3X�\E%�l�-hpQ��6�
c���X~�s&#�Eb���	��N79	wD�F�u#�d���U/s�Ԩ
�W�5���Lj^\&�f���]�Kc���
�ӌ��n���T��;R&�n�Խ��x�H��!�N�1)F��R�#�Bh͵ḭ�%�P���8�[��#���4ȳR;(;�I���HN-
B�|������?0x�V&J�e/?�G��@�	��)@����h�������X����9X�yv���Jc�1�����i����2J��:�ʖ1ef~+)6�ؤG(/�v�����gc����/�i�4t�D2#}�R�<R�-�4Gخ��]�w^�i���M�SQ����7�g�yIj�jo�J����0�j�!u'�<�s�qH�C��\a�s����C�7��Ux.O������
*���7&b����3��l`wn߽��%�����Ql>-r�\A��~��S�}�(c�ߥ�g�d�S���u2a�-<����G����K�9��U	֜���-�*b	O�Y�$)���7�*d,P��DàmM訵R�y
�B��3��s�BR�mޤ�a�7�qg;�)	�Ф���(��	X4�-5��w���5Mم�x�HT�C��>�{3%)��>8�IQ�*�&�[A$1'�F�ĭޣ��7�Se����~`	��_��3C
���zr'�Ƴt���3�?���7/9c6������!+���2;��k�xW�R�h��]؝{A"�2숯-�<Ƣ��!	���$�FId�4ʲ1T��	�V�#��$��w�Jq���~D��ϖA��VO���S�>�<�2���4�@�|��]Ѧ��ww ��N3��R�1~Y��$ޤ-�f������C�I�L i��3����{xP�X)6p�fh�I#��܂���p��P�e���u%�[Tȵy �cԺ5�;�m���5��U])�k�=@	r�iD�xOS���$�3� ��S�4�C��hz�qǹ�o&��������P�^�?��(���qO�8�c���-�8T^	m�(b��?���b5^.jUn=C{�/����h�dr'���@t�x83*���: 4/���@+BF�8��	 լl�c$�!%�|��c-hR{O�Ak%9�'�39��!���}7�xː�4@�!���N��� �E8�(A�/�a��.��^ANsn�֎�Qy��[����;�p���B�����m��Y���J�<�%��ͳ�}�m����� �Q58սt�1�1Kg���8�����8�Q��2���)��$��r�vY����z�۩b��b�g)��yM*Q�����#�3c]tz�8l�^��)�����KƱZ���E4N�Vw�H2�a){%�+86��Ǎ������W�N�����B}�v�\�Z��DBx�~�IP�FM��Z���A��{�K������@� ���$�:NX����{C�&���9ZIU�^a�?�au��h/��cՂt`V
V{З
[*�$XMkU��A�z���}�� ճ�������?thB��@@Z�DNʁ����?��b7�J�"B��.$��x�4@���U,�!7����(9�qJ�%<��'u����I�ޗ�4�M�'{���n��ԾV,z��
�:JJ�jǁM����6�f��զ�yf�IoC$�tb&��l6[E�������&~'.����D&_�(�;��q7�,ȮdH�$�Ҙ
OU���^�u�0e�5��������5#I�dc�J����OO���׵�1!E��v0"Cs����n��#��4<�&C��:zE߷ɆCv��r#:�G�`�F¿6���~��`��Q����%R΄��d==��ޖ�)�=N����EY���>��|�>�?��!���v�lgL(a�M��J��x�+'`���քl�HeK�a2�A;02�+�H���Ƽ
`&���\.�L��q+���6Bq�C3�FR�t��j5�q��\�)����ݝ1�F5��*Y�Cq�&+�!��WC��B�c࢏�TV�#��z��^<
���Rq%�J́�i�<��E(Ӭ����rS����[�ҹ+�RcM*Y�O��<�<ĸ�@��6��'U�V�����k��������O<S��ږ�m�$B`H�Z��,����H�5d�����aY���;-�O�7�uO�^�����6��Q}��%
?4�0h��m�;��TK�̤o��%Ӣ3m:�{� ��C���Բ r��(��(@ˍ�G+�4�h��F V��=$���=ĎO���#T��a��3(A3�Cv-,�%J�[���%nM	N9@�ޑpF��i����n�� h�[�̼���GF��U-}����-��j&e�� �A�����0�����xH�8fì�T��ȸzB�8Q�AB�[��9S�t����T�觔?:E{���~��{�!��̆*a��"�- �,䏚73O�"g_^�d;,�X���v�Kȃ*>^�H>�JxGy>=�<S~K�=�6����Zp|s��<B/ �� �9�fԷԝ��������c�)��6FK��^�F5��A�2�%1��6��,T2��! ���b���&r�k8��vzc4���yX��TEKx��2yqv�� nA�=��k� ��(D�ׯ��?��B��@'�E���/1�G�֞�=#	�C��9F�D��	F�� (��l��L��Q4�SOf�'��|o�5���MWi8��rⳑ�Dɹ+��:YE�{��δ�׍�ajJ��nL2i�jj�{���5�1�����ݰ����Gvf�S�n(ڷ������{w=�$�Z�bH��Id�<��tC�N�(�|
C*��]Va��	*������}G�.�ą���F\��k���S��=1R��!A0�<����d�����P#Gr!w�ŧ�f�Sd�'ǝ6$�DAѤ"���l��Z4�ؤ��^�������X�v#�(#�F��U^u'�B����$��"c*O��j�8�:���C�� ���ѝ�ɮ����S%��^��%ճũg�a����~��D�I�sxB�<���sьi��k��`-��XDa�]�ЁG��&j��P� ƺ����V��v��|hNk�}evx�Ŕ*W�hS�herb�-*������h�&����բy2�ǘ�W=�����?�P�*�ݸ=c^"z[�⠇���ᗘ���W1�5$���Fz�7�G�a5xZ�Z��PJ�F�Ⱥ�p��df�B+��3lP�����恙껌�7�s�9�012�O@�>E+ZK�l���8��$�:�)^�� ��~��; jo��,A �B(��l{�t.����k�[f|��sy�6.�^�Dc
A���z��tW���k���d�:�^��v��|�Hn��	;G��c��l��5��WHә9�����E�$��Qk:��0FX/�L�򴭝�{k�/����GO�̱���� ('U���	��lTg!f���P��Ȧv^eա9��.n�!J
���,h �<��њ��DʖXC�ڿ����b��T���}��'����}��([�H���CKy�q�m�pf�Y�ʵ��	CzU'��B����R�f��
Iއ����h�� jeltR`������[��]s�X�A�;&��P��+U�A��W�BA?Ո�Af-H��Ha߄�:K���KO,�O��M@c;4M>�(�C3/.��Cg�	�5u�����������{����6y��p�Ka4��T��B��b�Y�į[�?.�s|�)��������k�x�(��感�ћBW���_���mI�1o�_u�_�$���͛�5[�Ki'2�!��7��p>��?�Ȏ4\K��Ʒ���-el#O$�7z�"�CUI�Y�X{��V�14�5�Fy,��EXG��2z���}�hG��=�k��� ��4�0x��ؕQG��W�20���6Щ��a�b��ځh���4���#y�à&}		Uj�C&6�v�l��(�PQ��	&h�"#(OZ���RS�B�>'����38��w�lBle��u����fQ8�2fs6�T��u��E�7�K`��9�U"?F�#�v�f�0�V��9K��f̈́��m%<�\jϮo����OȊda�?sQ�@����2���Y&�,��-�"U�s����ނ��Ʃ}ٝ��7�������v�L��?�P>���d��<M�`�~]=Awc����	��c-��� ,0M�NC�Tw�m�IS�f`��!6dx���� {��1��eKOk��B�qP�U6vi�~�}�PI�aǢoI��gE(>���kv�@�'�Z<Bu\G�|{!�֛B2�����3;(B�	�����zʋ��"�[`����A&�R��vm��V�s��7��Y���; *3�żj�����a�H�+�у�H/�B�Eo��|��*E�o�*[�'!+��ښ��Ւ0����*�.�fߟ}�3d�q��AL�8�q�!mgޫg�aD�`�5��s텈ak:x��l�;��8�m�z�u��~��~N#�Kl1w��I�<�v��ү0�ޙbY"
UN'�jFz�J��:�H#c�;��IB���m��E�U)8iU�ɕ����������]�u[�z�X�*̨�bx2麷&_�ᬩ�Xn�B��n�cxEZ�G�ֆ�X�Kt�;��&�B�ӳ��'m�ǽ ��\ST��ЈK�崧��HU�Dٺm�s��E1�	������hv*�IOlm�񬮁��+�sTC?�X��诬o��CZ��_�H�ܸP}�͓�N`[���1�FT�-���I��8������PÄ�AQ(�b�]ЉJ��Q�4�6$m�7|Ll�s¨c~|���!G��(��*�zk8��!�l����5x�4vu�n��L�Wf��1�Ps?�X]윆�|"�^�y�tj�n���9�{���HmM�Sb�2��\��}�l����'*S��ӲF��y���Lc�"y��Z��������0�7z�*���ƴE@t�:x��r�Tᗰ�Ȅ�@�:e�+��M#��j�<��h.8=+m.�O�)��N:n3͘`'Z/�����D���D� ��0�0$��I�$�F��da��ĳ�0��������|b#�=��R�����Z1]>6�� �+s��!զ(�- <*<� !�\ѫV�E��
��I�����uȠ ��KUіI7  ��IDATX�i���;l�y[l*y'�Pfpe$u�o�O0/f�Ϭ��}����M~z�c���e���,!���9ɩk�d d��"/�.$���qZeL�x:�I�5��~�t&֚k71D��A��	�')��u�t���Xɦk�b]HR9��E]�h��a
�^�=hs	OW����w��\D 4[L��֚����|��I&�o�y0�W���� q8S+֌�B~o-�U������=b3T�4,�`���zgZ�G��6e�E�PF�ɐ�W�c>y�w{wsj��+�Ѹ)ԑ'dX��m1�h�Cɾ;9ز�&��:��%�:��	��O� Rưr�6p�H`��-�s�t��g���,�qÚ:Ͷ]<��x��������M��&8A����&�`���!�P{���k۾=���%��Q�n��Ђճtze�٦��Au𾬋��񄐴�3����ɉ1�i"�'�D���G�1JhQ�|����;�q������1�u����$�qh���E$|�5R�*ML�T����HN��e?�.U4��B��yE1DJǵ���y�뚇?!�c�����S>/��+<5Js	?�']��^_�s��l`d4J�����u-rv����µ�9��lln��[���6*"���T���S�ǯ������s����5 ������䡆*��o@0�Ř��� ���֛����3V�.��%?S�\�����Ҳ��e�`�A&ë؅��Y��C�ϡ8h>PG��K��V>&ʓ���~�����C��ֲ�x��"co�R��� V�h\�2���C��Q(��?m�OJM�Wԛ�bÐ1� '��$2�s�;ٗ��J0d%�+�=ȳ��`OC�l6��-��F�&����I�B�s<S���ᴔ�����Fe��Y�����C�~��>��IG7v���zx�� @�p�9G3<;~ַ5����-_�7##i�#����Y��K��kp:O��v4��H�����o-�xKg��z�.��C�߾,�+�)�mM�
^,a�
7z]c��'�Ea�t�kX���@22�P�O��DDF�L}��m���������?����-O0�.�s�t�G���g����u�$1���<ٱ������P�F�s拶��b�{�ͤ/)��RTw�-�	}�a�����[���0ɶ1�O%�k�����Iy-��a�� �u���D�U�,��6S9j>��*�����fl�!�K���~������%F����sXn7z�p�2�)C�5�
w
%Hƻ|��2gC�0�g*�?;�ll�Z�����+ժTaT������E<���k8�Ґ.(��0q��8gba-��iH��J���%U�IF},ܭE�U,1����sx�)�T�F�")0�#�9����oL��?J
�%z=Ӡq��p��I*�t���c���q=*y��# �\� {4����2d.�m4��#Y��5�[�y��!lk�~����8yUC�Z�VB�W���ҷ0uc���`H��Bo��oƇ��6u������ZVǁ�#�����?h���@з�5z����68�H4y����.�ۭE@�p�<�HHi��_Z�<Ҟ*�p��"i��U6�ήI����5���}�/�a +��r�r>*1�	�]��� O�W��̓5����Ž�Oz3�/���U��u��0�`]/�gP���L�P���tM�PO>���-�pķW`ZBn��A ���M�a�杊� �]o�$k+��s�*7d���w\�-C\�p��1E�[a���֚������6��¿=d���e��~� ��
�ڈM%�+�,�0��$p��7��=���ū��B��O��Ao�煂�9D�;���s���-��_}L�0�}�γf�\k��;�u��qy8]��n�	���}RԾ;4�ԍ�9ᎎhf� c�m�N�2��u�>	˛G/�ņ^��K�7i�����H�	UG�2�m�*�v�S�y�7"�&��KV���n@�g�k��|�G�	3������ߧ}M]�����O?�N��^z�_�pb�<R���L̓�Õ�ɐ1�O�7�Bk����S��R�M^���q�k��=���D�_;�/��c����j܇�u�=�(��}T�����钺��~�hW*���g)ۍ�*�*`�|a��M�J+e�E� 5��~�]dH�4��8 )����YhZ�>4�p��	l�XJt�F�t�O��_�_�	}ޑImA#1��󔑓�r	�w�М���u�����S�2�gs�^y<\�؀2� RϨ�qxa4��r�C�q	CT��l�ǚڿW�=+�ҋ-OR�	�G����@=W������|]/t�j���(
�A�;��,�_)0����v���4�{~�\����Ό���~~��T��ӛG��"3�u.g��k�#������P��wnU{���5�k�;�f�D}fR����@x���;�i�XX��C���?��=������݉z�����),�m�ZfK�ݘB�BЏ�9����2_��1Ѥ9,`iz�����u��F�#�zuԳ�TB�xI�q��^���	�#T)�7-��v*w�:�N�$�駟=�8xu�]m��4�6֗�����׿��)W�"��F�:�������\e��)T�R�Ěf�>f��� XJm36�����"|� �V�#�4��>��w�F�*�\`��o�*��D� �
�v}��^�-.y ^3�Β�O��dz+m�GfX�gQ���p�*���uԈ�%44�Gz�`L�a����T�ދ����R�*��
#�O,���5덉R\H�����I�o��nkC����PZ�F�qh*�5�}}���ZJ$� �sp�ʻ.^����I����~{i�wO���Ș��12Cw{�	E�5�c��r�_+{-�5�j�������w��`1�2��7��Օ��F�0L��#�5և`����_����Ç��/n���/fK�pްQ�;�����������C���Z�$�x.�-7躙�����/y�Phnc�yl����y���}h�R��d@˟��^��K�a��X��	�^IC��yi.���ވ�9F�y
R���ׯ�a���z^��0C��<J3��e�C��OU�l�7��X�]x���M�3R�N�� ��^����܀���9��/7����]�,c�p��e%P��'����B�?)\-��K�]�~�Q��oYg=�1����eM����Rz�|+�LM�Qna@S��v�d�JIK����j򽷃�*c�Lxm�mG�/�'Qx���(�Ƃo=<�
�Zpd�[L_��A	n�XR�04�4J��>��'{6-�&e_"Yu��G��}�<{2����{=��(/UuYT>�C� A����*͸�8|��L��9;3��'j����;u&z��ռ�5�x7�c�x��}l��=��ĩ9L��~���K]�g�ӛ���a1!P�b��5�]DF��%��Ci��@�{�����P��U�҈�����GZ~,�u�����Z�zn����zߣ�xf��{��믿��Yϗ���/�/�y��_b�fVk ��99���~����Jr��a�����waM�L6������`'9U�D��l1�^#8a|��XsFï����w�֢0�Sh�<Ю�P�$�њ�g��]�����ſ�߆n�|J�ŦvbȍF���zl+�]/'�F�Z�������U����r�"�%~c8Z˔�Qm@�&%%}ٳ����>3��s-o��ꞡHT���\"lUqȫ>�HBs���0�K������j���z3�v���w����j$7S%��ئ�ac��q�c�i�&ܰE�N������D��,9N�ϕ�S~��-P[Ϗ�<�2�`N���P���k�-d�����kTP��I�G��u{����G++W����ٲ�\��a���k3�|U���0m~��Qdq�қ�н⺃(4��0�=�M�Rm�Lx�XU��H�SPVx��	~c�&�^����;;]^����^=%/]���F3lϰ����g7&V}d�����C�8v}����������w����F���mc�P=J���0>I�8$��pH֬�`d)����	�8�a��kT�}ߤXH��z�^�7�x�fc`��\l|�hH�G��&}�h���T�l��ӧO����ϝi|��э)B3`px�$ԛ�:����<+4DR���������?�I�+E�+װR�����K��MKt��p��e�g(��F��`7�-ɛ�\�?���G5��0���@l��q����~�:����?��%-Դ�s��kH��7��@M�"���K��"b�鑣*i	O��±T�M0G⠕;kk�<Q�u_��q�	�R������5���u�|�("�p�H��֋㵞Trk+X5�[������������e�SVӍ��yD�!�G���!SH6��GZ!p���;���.B
�?��Y�j��9���O��=�D-�f�4�=Rm���	��O���������o� �bt����]_v�?�6z�jG!��hS޿k>��D:5�`ߓ� �c�\5��Mrj�Ka�=��G���q��y��w3Z��ԖLPr�6�_��78Fy2�b!ݗ�����fs�H��j�6i1�Ka|;�G;&$������)�ky����W���PRN^�LOf���¸ps�!E���z9#��]�Bo����i&� ���G=��x
~&��%�ٟ��H�6t
�QR��\,�6B�'?�bnm�?=��6���(&����}���������d/K�(J8�QucQ�5-���нF�}�d��z���1} ����5hp6f�/��ze�9E�asCEC�?�W6>���԰��v��e{6;�?�Ǻ��ʵ)#)#�i�#�:�2R��?S�:���ϗ�.�v��1��2�U�rp��c@I����ռ{�#M���_={6I�z��î����mHi��*�7a������Ÿ�g��%�B��W
n���뿹�[`�^�9e�E_,܈�E�EUI������~>�r��(�˵$�m_D��ϕS5��i!�K�D� �lk� ��&c0�H@�QU�*�L�h f'�iM¨a���>���0��H�m#:������'=zMvm��|���>v�싿���/�^���+������x�dH�^�(��Ңe3��4�g����1��ȼ�� �	�k�2Tz��S�^jYݗ+=��d=����8E�s$���!<-
-�f0ͥ������땉�[%��~{+��^��u��(Eϯл���xE��`{�׷��y�O�����k���{sL��Vѧ&M�L�&��=������m|��Lv�i���:���N�5�~-Ga������� bm�Vig_�!�a	"x�ͯ���r0����`T��}�(/t[	�3����ڊ�ꆷ���^.t����M]��$��r9}utT}М��C�<�e�0�K�$|� yHCTGܖV�d���L����@��:�z0�D�����6ڀdr�Q�3H��B!��3���{�q�xo?.=�-��֘p���-T�ά�u��}j�݈Z+c��jr�H=����3� �Оg��&��D9RWό�~�ʡ3ͯ��Q�}Q�D��M�ߖ�{xs/�|�Y��+*p)l�^׆��g�0�;�t��%t��ل5�����a��D�V����F�VOgMRJ$��n�W��"�%� ���Q�\cy��.��J����n���˯�4H{5�@{4�J�g}�Y"���8���Q�7M��f�:g��-^��rhu�E�� ]��j�l^��Q{�ʧ���y.9.�dg���86F��U�﵃�����W�L�ފjx���7 *��{ ���Di�k@�J�����;b<с���3�����yH���P51y�N��>�!�	>�d�3��F�z7dcJ�-�HiFq�����;x���%�`�GzѼNYK��WL�M�1��&E�6l�~f���9Z?� K���oϬ<7Ǔ����*���<���fp�v��g������$~��O�{V�^<#M/��M��f�����/����'ь^e� �c���:�gay����:ƼO��_��/�+��g��&�!z#f��f�(�Vx�ߞ!�}y}�'o�����Ȣ���-�7��w����%�4�`(Rq�_�D�_y@���Zn�4���/~(��g�9h>nh�]���,���J1{$<q���Yy��0���K�A�ͮ[ʊפ��
����xeh������x�v�@L��<��m�Gm�)ǸO��k�A1J��phݘ1��[�.�A��):���3��%�?����^�B��������:_��߽�"l"��ipC���#[���`�M	�em^u�n��M告:h���rISw��#���=����Z�iu��]x>��k�d�غ����@�q��\��V���� �hQR^���]�,~?$�������"�ᚼ
UH��B�ֻz%���[HB��f*ʈ:#���#���U솰E��C�Ps%ff������B���l��R�kF�J�f�R���Je!�ί���;Q�⋝���y���gFv��+K�+��v���M��)��%.����no�}���EHףc*�k֍�#D�rTu�J
����^x���~��eU���y�9 �W�"�EGC�}�̯�53�J��>7W�A�	q��kO�0K� P�A��i�������Bs�x����y%�P��P5��mu���{֚ծg�{�)���D�a�E�E4j�\ғ��󢌗[V*0U���l��-��2��Ψ~���]�[��G/��H`�SW��?FB���bu8��������ҠNA�Z���=�\��sE_��\�����)f��=��RT��^S��ڔ�<�y�£�x+޶�N�d;�?���OM�<̓�K ���S��5���� a�虡��ױ��2����\�%��ၭ����b�F%N�pf)���"����i|��!��Ub)(�}p������1��{m�AM��[�������#-�G֢II���@O�젇	����tf�
�a�,��c$�������@!�g��a]f�	���8H�~
�����Z!5o�ڲk��K����%VJF��h�w^��*�9�%0�tK�J�9�nG*�	r9����%��@�q|�_L���(!��u,��,`��nٜ��O�(��>sf����(=���p�k������NB�i�o:�8�v��o��D�U}����⤩�8�R��sO��Pw��b�ѕ2��h����
��)k�O�\�2�[ܾo����ԝt�frJG���A~`O(�|�����qnC�w�a�a5F�V��hk�s�B(� Q̄��{)��j�lۖ���8M@�^�9��8�|�Bi�w[�
���.�Ր�[��T,����ܠ�ْ�^2�RwOc�Y�Z�ը��Sփ?��8�%�GC��gS)fXb���B�+�V㒅
��9��U��Ͼm�e��"��Yj�HS��{&�	%�	9[�/>9�f�،93��p�1�(K[39���[��4O�Dt�����6�ڸ�Xu��#�^vF�U� �i�g;M���V���+��9sb\ ]��4$�K�Ģz�o��k��Z1�=Ӕ�p��Z��A4��Ϝ^e����H�a���@^E͠��X�q�K'�,�2���QB(�����:�J�vC�ғ��������Ə���q Ӌ��k�R�H&x����y���iM�mv]��-��M�� ]*�Vd����u�j3���}�H�k��� LvZ?>2��jMQ
��Ή[�jt���Voy�(�&#�%�'��9�I��O�u_]~ϵ�ke�4��vǊ����K�	�FG�͟�Θ�v��W��&D��밐�
�k��eQd7OYJ�_�c<Q!輨ĒA�E� �$z�	�V}>{�C���~��Vf�{z���'�w��;<�G�*S��[��i��ѷ���S쯚?�s�%�j�z94�kG��� L[�8��;3s�R:�L�����/ѝ"<qFsF�b�NI1Wv�5��
(~�~�%M�&%��^K�����rE����^��m�v�1H�L��X'�H�4?����<ȉ��v����}�XB���6�clȊ��{��7��Ĥ����~>^���^s��p��!�¼�Fib�1�4�<�&�`&�����癉H����n	�>j��#X��t��:�Nćט�m�U:7���������<;�Nl�W�w=�d��Kcv����id��F,V�@�z)���HF��DWQzt34b`�+�E�����{Y�H��m�G2"l>�aa �����a��\I�fе���TIǳf��xk����I\���A�G�-�kK��]RnP�}�p\�>Q@&���5��������Q��:;:pu�I#a�U�M���ɨ�mm:���y��������
�1�)�7&r-
s�Cd�%A�Mp�][�����X�V\iv��ɱ/��g�z(��[4زMm!��CM���̪F����d�i CC�����nz.i8�ؚ���G�?K؎�{��G*�سm�_��X%�G՞�x�wϬ�>%~Dϲ*�(�o��񊗷��Og�������Y�8���3�	%��[�O��`����.K,kX��t�u�L�n\Nx����N�Ff
�bl]c�(<Jݣ_��\�Lu}m���� ����)ȡzy��J����N�ߝk� 	�d$����J�f�b��r<���|E����z�����)������D����Ycoz��
�i���՘�NY�G�q}
��E<�9���R!�g�i t�ߧ
܅�ԓ��R����DM�3�Z�u�q
���Y{�*���L����� 
��H�NG��o��йx||�Cv@�<��Z/��ER=�;���)�ڨ_>�}��������UDl��A�yx~H��G�L�����2߲�5� %_�m��n'��yT<L���Gc9�	���Pt��b����\��Sb��v� ^����W���S������"2��3e��N%X�.G� I쁈����c0=V��&X�y��Ku"���n����E(�]WK(%� N�}s�u�0L�k�y�<�J75]��tְ/���wWrŗ=z��F=�e�#���6�0���B�Հo[?&?��s��g|�{��ʒ�:_�o�9������ׇ����w~��g�\3n�%�>�/���q�8؄҃i�%�����)����X'eJ��[z�����`ֿ���u������F�p�������r��z�6��4�������gBQ�S�pc�}�m�}"d�P �w�g�tv�ѭ�����G7+ѵ��k9�'������"㋃�Sge=1�$+oA�pp����p��T4B��%:b�Sn`?y�,|șUD��d2K�pz�'�����dx����:��w*N�rё�~��V���������g�����}��'�PO�m��n�$ʾ[�n)������O���4�����:z`m�X�8p2t�xVz�Bu�Z�ў9�>�ث!���	+��Y�b�2˙���c���ʘf��L��`�3m��QB!p�4�����Cf��I>E_�{%���n	u#�ε *_�����Gf�o�>���1ƭiT�T�o��Ӊ��I���#t�L���?h�������G�r���� v��ri[��-��N���ƫr����!Ґ��ф�&UPϣv!�� �j�b����h�3��"��p��L��/��ɲ1Oh�-�"XF�*Ғ�r�y
�N�`hk��'�����Қ���B�����tcy�N���=y\��d�MC����*��0���%/!m�c	⟀u5%yZ�B1��� �2'&�.A(�M�kA0��B(+'���yv!�o��YG�µ{|̦hØ�=�+�����X�dA���-�M��e󨓼-��tHZz?�1���72���%��b�������px�Ej+B ��~�g�D��<Kz���g�n�q��{�����"1ha��̓Jx��G6�4��D0ڀ��|#�V{��s+I�i�}Vq�a����4E�DF�&|}��R� 8󠓟<��G-zC%8O����	����٘�uU�ގ��W�Ƒ��z�P�X
A"�P�d�{`�W�^��vO��y��{8^���y�n_,�`u��;�Eg��d6C��1eN�+�I�!��d˚Yx�0mJ�ʾ�^^�7�,4N�ĭB>���� ȕ7C��m#�b��L��4��Չ�M(��Q5S��(�[8YcTH�x*�'8�i�2#�p�+��D� ��D��� �Ao��Nb�L�W>M �[X�NI���iOz0�?Dj�8 nx���"�L�@R���(-�\�5�(0��{�&W�1Q9��Z;,؍ắ [?��D*�e��_��՚��'��uINȀ��m��ck��"9E����a��Q*����4J��FQ��z0P:���9��Q�]in<#�[��Fz�T1�3��d��=�Z��-9���T����@R�o�b�ʪa=�~���]
�����U�Ȳ<���n����
r�#�n�E�X�)��q(���v�R
3����?
��+}�6�۽I����gci��=�8�e�Cz��H�A�ˤ/I��u�`�p�v��@��0�cd�e*OpݶX�
��@FĿ�\�7s���	T�NWK��{�9�~o�Ǧ`�/�*��&e�;6��q<��	E���&)Wʑ�yZ�6�f����]��p��I�F�O��X��gT�",ϭwC�y��5=�X?v�=Jj�N���P��.
]�Ů�Қ4���צ�S7h=$e���y� ��H�� ���]ԧLؑ28�k+��V���\�5$`��Ud��h2�|eBi�k>n���l&L~W�\�?E����^��B;�ʻ"�DkpE[W��E�=�w���x�5 ���6F+ј��e���m��w��y���
��nأ��j�m�G�Y����a���x��Zmas����U�#+2Z�yMYs��}�ó��pT�Q�a�ڽ��H�A^���G1�ū��]�Ji���o}榋�~���g!�yzO�B��	?��'� ��<tk�e���H���np=���r�k�D�I��w��*.���=�,8�+Ac�&{�\������
����,�K#W��� �Ry�f�
 �޼?O}x�SRV�}϶�#+EfNl�@��>29D(�Q|�&�*�}��������$�
K�r%g&�G��{㵼O%��� �b(UQX��z_HL*�0��r0�v���8^;kK�yB#=J%�4g$3�}���^0�����w�W�PPcZ�������������t��VEj�5�Ͼ�o��&����U����R�"��z����Q��Ǻ�ٿZp�g��G?�F��[eõ	�/��G�oٳ�O��F{�U�\b�Xw_0��He_�����dx�ln�PQQ�O�62�epʦ4,eh'���
o�V_ؤJ�׾OlKb����BJ7�� C�F��J\ś�:�-�(*��(+F�ڽ7ڪ7:7NXTSRO�f��+~�>�B�H���$���Q##�k
�D(�{��f���I�Q�c!��c-�
z�2��s=���rO�AW	�Ŀ��g�CR��)ֈ�>g�����`Հ�Ƭ�+�H�d��W�47�dD
�5>ֈc��с�з�I=8T�%o����J���!�-i�[�����Z���=�sd�3V
RY��f�jFH��^^��:��5^46�W`Wn���#;p8'����{C:�ŕFT�?�u[|7�mWV/A�U�Mb�q�K�])�B���Y�P�YU�,���ޘ� P7|:�eZ;d�����]�T�B�W��
+ܟL� �F-��6�-'�o�rt��AAG2�f���5c�$�/��U���+j,���J�Na�Ě���<���k����m��7*���1*�&��J$d��/��#�{=���M^<�C�.�^�����s9)D?��m��jR�
�b�ci}r�#�t�\�S�0E������KF.�ےc��%�Gz���}�{��{=;P�A�JN0�1�{��[[��Ҏ'�T�T�Heü�˓E�B0J�ײv*OɳB��!"�nWBz��BgxJ��ʊ-	�g��!mMsro\��������N�!���z<�+6r����!�&R,=ڠ0-���K�J��?��IZ��k�2r��V°hLඖ$��56�}y�(7�D�V�0(٤���b6�A�\�F�[aP>�.��$�ɘ��|�%�6��
3uǶF9��W	��t����w�������Q�1��;
��;�,q��͝��L�lM�Sz�%�tZ�m�e�������Z[��Gn�|V{�U=�d�x���2������BG$�Svo|�1�Keg� ��T+��K�
�|�v��_��?��ڢ�iO��[����2�����L9Ӏ�~V26��S_�~V�h[5�!���H��16c�.f3@��r��&�+T�3�9�IkI� �qJ��Rѧ�0tS�y+ޟ����Pe��5���?�!6��	���	\ɛh>��8D�i�j�4���6&l6f5I��A��c\/)[�=[ve����vO���K�CL���-��ʲ6b��ۿ�T���^[����8\���6DS�����W9����0#��y���q���jk�|>���� ��O���L8%wQ�p�~'����t�9'��Y��dUG�	_[t���m/ܿ�N��n)8y��s��@�!���%+H�
��4��,<��T� �?	�c���=�w�KMؕ�մ�/7��ϕ�x�㛏U��]�1��\+n��VA��s%#����y�EJ�c*���yJX��$mD�U󥹚X5&ÿ4�<�C�VM�o(K��FaH3�;�������+O�,Fҹ�Z�~*��|1t���Z�׹E��D��$t-~�͘�3�>�{)����2�20��̀��[ԏ��X{[�m0��BZ��T?<
>[�W� %Ɛ͇R9�~�n8uu��u=�d�mOz�,};SD�=<��@������ocs�ʦ��q/�3UC��7̌�\��@����>���X���Z+/Q85���J��D�G�Y�Wx[�Ű�nJ�}|���<�շ~�{&�Z1�Ca4����ш�0҈�w���W�Z:���[w~埱<Q�x����c썭 ���p���������.�/�A$s�
�]�F��y���g֭�[�	%���Ys�T� j�����?�QXm-m��M�+�ȯ?	�7�������t�w�R��x��FeH�������xc��0���{�)����9yV�v�Z\>�ŐЁ<�Ɠ8-�a��)����{�%aW �X���hl�e�P+��|��9���=�D�?�c��·�D=�1u#�O����VH����p^�{��*��)�#{�Yb�eL-�{=����W#�G����Hc,�2��%Z��p&O&��:XQ:�yP�PHj[�!������h�^��gT;�AQ;��a��H��Z҃�i���Q��c�W1��h�RR�9��+?gb_��!�nI��\~�uam�5{��RyoJ���M=v���ɾF��	,��JD4j�[�YN��, D�T!o)=� ҅O�P/�M��h�Г����iz�%���^'.J����5��sEH~�N�or��X���Ky��=�,�*[�����J��<��縁8)���U�#�v�rduT��%���㖷�wo��H��X�v�Mkഩ���4b� �d.��שM}���8��/V������l�޲��/���/�ևxh�e�?V}v|��Q́�aS�[x��q�%�kO�䦸?�����(�?�_�"t�P6<�e�씚������Ȍ�` 4Q��Č���Z���G�P�ʁL<��'����"�����#
A���;��5������d��<@$]�:�ש#�5�U`]I���Ű�������4����o5��{[��.�?w�1/�~�܅�p(��K�#��S���AL�����Z�O�\�s��們fH��x UYHj�%F| Nh"kO��P����c�w-�s�n��v��m�E������y�s)Գ���M�S�ZJ�	:�,fW��8(�1È�g��]/�i{��%0�m:`*:��kD�*�)N��f�%�a�����B}]�B� ���V�hn�=L����Y�j��|P[@�b���9�c��T�i���z���^۰��m��l��fK��PQ�����dٖR�ڷ�mM��s�jM	g��g��w̏_�*�`>*C��C�ND�&v�[�62L�;{�q�1�z/���#���y��IN<Ķ��h�3"!��	�5��֩_�!�jwT9"�!�G�V!�*�T:��G�v0����oV���Y�R9&��$�'�>��E�fj����<p-*��g��[��+���9)��w:UD�͌��*�%ޮ��:ΧbH/Njwל�峲�]��ĄZ;jX��0���,�[��3L9`��.��k���<�8k)a�'��@�-F�qÑ�d��[�90��Dg7CH����Λw7fkR�&��*������zi'.����/O�~�=7��ǌ�8��uid��p���j2�-���]�fs�ݐ��J�x��Z���-��*���V�#�`y�7���V��=�%���R�l�ֽ�95�kNQQۀ��.fn��`�jV���59��%L�V6S�	�6�=E�ys��fz�����	�Zz�G"���XK��Ęסx�CJ�+hF��v��Ġ�[�f�3�ͻ�;���,A�Sb�M���BJ�^JI�;�q�#��l�)!�`��X��O��������5�.�	g<�%��`e������Nʃ3�'.����7��!���Ki��,��!6��@�GY;��r��-��'\�yp�$f*����6b,�[���]K;[�*�a��eɊ�~TfOC���OLS�_x�%�����I�W�<� 6y��s�ic�����mE�QW?x�a�$�+nz�c(� �3��/��$����s�x<(���z�7�ÍS��B7e^}-Y����a�y?PU���5�|��h�3�v��R�ul xˌ��4���l�e�QNzu��z�)�����j��V~�(uuouagw4\�T��ҹe�x��iD�labɹQ���}|h+3���v���s'�S����x\�n��������L�̑p��u
�O�ȼ�J��	%���	���CP1�.�?�EA[�bZ�מWa���u�By|@��j,����hd���ᾮ�>�*a<�K��l���9c��]ɧ����g_�6(ޘ�m��k�ɓ�6�?�p�p���)�=���Z�#mxy���+�SW�b��0|�Yn���gW���p��S���ٮ/5���6��a!�p.jnȃ|S��W�߳)՘@���u�TE�Q��ͤ�����bHÓ�ސ!Sh|���+���M��(�hdZ��]�ߪQs.����0�1؏d&���NkLR��Pޛ���Z���O�R`��S}L��hZi%R+2���D\ч�V#1����<M�˓6��&	"[�gF�g�pJ�˼��l��g��s�L}��cd}� 鱬�P+�A�f�C�-+�����!	5O�9[2�0�������j�+���ď�֖�ze6x�SQ^NJQ�'x�-V$�VЄ`_�Z�լ{?{cD�<od��T5-J�����E�+�1H������I[J3�6u,U�0@�r�HU�Y��3��b�Ʀ��C#
u	MF��K?l̑���f�%F�;���Wb<����Rh��k�7��$n���2����Xɫ��QRJNX��IC-.י��ƃA��Z=$������Y��LJ���Ǿ,\o���co��-1�]�9m,����-�v���H�J^���fFPՕ�¼��Io���o�JR�=u9,a�YN����w���n�Z����{�D�d�_uy"Ai圧��F�2�je�I�R�q\�r�����&l���1��u�Vi�s��0�O�a��Z6׼!���h�W�*��'�4���!����FU�oj���їB��ͅ���	A`��K~a�3R�P6Oy��UY�ۺm>���?Hhl��;�����x���d�Y�U'�xP��2*ԩڶ�1��w�A�%~YD [�ыW�h"[Y	��EkYi��}wy��*a}g�j�Z@O��f9+Jh�\8ĩ��{n��{#� ����T��:���C��,IY�������	L�U�
��L�Ł2NGY׮�[r�"��{�/��2���X)Ό|�a�A�\وǽ�!Z�܋9�r���qC��R��.�Z�ɃG��d����l������ܨ���-�}_�1�P�)K���
����!E)��n��U����p��[\�Q�� �[N��(Ƒ�e���cl��%���I����\���)Љ56V�N'�hT[�F�;sA��.jA�
�zʓ�,`���]=Pvu0�+�w��2p:H�	8��`ȗ�A/�`�y�jn�����KY�U�njl��x�z�
��n���Nb�W���/nEP�E����3h�vMo�^�D-�{8x�����!���t�OF��2ێF�!��#B�����в��݆�a�Vv�Uģ�Ud�{t޽F�.�s�ͤs�ۘ��"�ۺXC\F0K�F!�?��$��n�oES�Ác�<����j�TlT�K���C����DZE�-���g`%��[���7W���K[gf�#�Z5p��x&ws�����u��Mc �$�2A��M�����F�w���n�rS�DϒZ�����0�y���?�7a���O-�<�v1��_u=���������u5L��wLjddP�L�	�j���4���!�/��*~����/�E�Wk���񹃒;iH3��a�8���OZ���F������~�����X{�����z1��N���V�/����G��/o��)x�UW��yL���!\mb�"g����p@��d҅��Z��	>��n���\ә��u"Ｓ.Q���o�jW�T�!۳�S]ac��A�l}sJO����FBF1�~Y=��k�WC
�
k��Q��b��O�yl\�Am�ӗ��r���A���D	�(P�V^{-;�����5m�U�;�B� �u���ǅ��m�_Ƕ�k��'�����%=��H&PLX�	m��].K��Q�T�e�
�{Q�[&���U��s��,И�g^:[Ġl�1��cN���V����7�u�Uꖌ�P��@W"p�ҋ�F%:Q��T7p��Aj:��Hw�G|H�4
Ð��X�0���RZ��܌�z�3�y�Y��)>���#��CQ�훸�\��Lw 6�}��A�5���;��%B�I8�i�=u>�r�Ciɽܢ�G�tF��a�����m���|��ѐPJ��B�;�P)G�$������sG�����|N��?2RG�?�ߊGş��`+I�zў���VfW���A������6҉'m=�e�8"�r�)��a,i���~ҙ�x2�Sn��B�T����Z+�C�c6���n���4��������A�D޿p˲��0���Q�q��� ��=<����*���r��f�|?6����-�ؚ�Ҥ�e�����h2t�2*8 >8������X����P+k?�_���Ua�\�e�5zC��s�4��@����k�U�5�w��[+��tB�pL&��mwi@hM����|::��m�o:f�q��>pZ����ɛ-{6��h'�q+y����'����!������u%&�
��* �)�'Ӗ�`�E��n[��)$ת҂��~>��|�ѵ��>�.�AR2*|7�I��b-Ƴ\*2'�0
e!�^���j��o��;J�ޓpc�|O2��k�i�I���Ɔo�:�X�,�x�5f�HB!���6$f�&��0N�ʩ�b/u�9P���¬��L��`�������Wd��Z.�b u���	ȉ�)��vwM��H��A�,����ǁ�ʿ�!��9��y���<����C��1�L<�8w��`���0��6t�H!����ض���I�8�T�Y��C�	�-?:"�!���:0���+y�	rY���#~��a�!�{o�6�k�������:t�aԛ�7B�#y��0��*��� ի�=	+Ȱrb�O}1�&ߥ6Q�|��߭�79z��a�O{8�n%^�we�OzD)d�gik� �:8�[����7�{n�$�䡈z� I&# �8no�e��P�����}T5��[��PC4Пr-t%�������e� ��]��eN���������쿟O��!>ϝ�e���!��mˆl߽�{��xώu���5���������w���ǘ��A� ?[��2-p�ko8~8G�����ݱ$7��{Dfr�K��F��>����y���nI���B2��xa0�H�J�3!e����;0 ��}6���s#�g��If�A`JsSC2	D���o�W�8�?0G���������������#��:H�.����T�N�8)Y-��]i�y6����DL�ս����lύ�O=A�E�=�@��*��t	EzeD���VP��#��#���	�e��MKM0"s.�!� ���[V�={��	0�e-���T1�e�*�����k���T��$8F��Ze��ʫ�]��y�$3�]ɓ�I��M�X�K��K�3Ct,��;[%R$-���&Q�v����@��[ey�آ継�3�D����tx�ͼ���E1�Ϻ����o�i�oBg�"t%<��Z��M�`�3w#ބSdP���C�?��KR�.k����6�=�����(��O�<�r��^0���&�0�q���,�JB��6�Z�h�Z�^VK|f����*��X�q"Vb#�E��0�}��zX�2�.�5s(׏��$Bu�زY1�q��0�P�U�И���Y^E-K���󭊵/q>=o��c�oV�߸V���d�9D�3��,����P5�|��rtj�̾UJ*vuX�r!3%�b�}�L��l����T��A�E�����2�!~���eֵ��C���|��Ϧ{M�ϤK\���`�s՝S=�d����ƞ��y	٨5���Q_$�KI'��Q��f-�?h�0e�U����G[��U�{��<_��[�����?�g��4��]O�բ�ruE����ݖ���e)�6y�ZM���,)LR�����^AQ�N#U�f�XU2�W�4��;�IQ^*Ҟ�R�#��CR ��RΗ���Ÿ���<K̍��Zhn��be��4�!;-B*��|*}%"�&v�W�A�N��d�%>��\�q������O�^��V��������-
F�"dRF��d7Q��]L:�-�u�"���F�(�r�k�F��p"��T%�}�+���4����{�������S��;�w4��q4���US��,�eȹ	�R�rl�M�tk%.���Z*c�EȮ��<�3��5�hX*l=e�*Ӎ|9$��^ݎ9>X�LL%Z�.W�{(�@�a�ge�R�&u��!�XJukd����f>��.��
�O���&�����Gv�R�1fI�c���ׇ��%:�l�(�z���m�h�[wC��ZD�=������Dy܅��V�؞w쑜3D��@d����,�F��u1N�I���҆;؋�9?�V;eii�h�xo�eI�8d�J��"�2�L�+�����]�཭�-�:Z���sYE�Z3�{(8 ��0U�ԳL���|�ޒ;[�RWK/t�+ġ�n~�X_��*$T]�P����BU-�|��/#�ò'�P=��2�Q���j��#n��y�ʲ��K7��F*6*sc��%��B��v/���ܽ��<���_#�+Y�������WE��{�ZA5�h���C	X�]� �(�\���T⾠����6c�O�y+.��Ń��q���L/����i�X��%3�Sco��o�DV�W�����c��͑hWLV}I�=n��Ҹ��!�a�%����H�m���$7�n4�V����d��*�?�U���b��:��qR�֔�c��i��	��Z��ZG>� ](D�� ����8�U�p���	@���Kσ�wy�Ճ5�h�l3yY����y/�Z[��*����:�ׄjK���7P.z{4�Q��G2C���Zl����H��y��ǫa�]4�2|޴�J�nN��]bq�+
5��+�y~Hڪzy�e��g�)s��Z.�]¥�%b��z���m,[��7c�]J鬺ڸ�E���{8f�D�S�_O7}�b�lPT�c��ŎE��rO�ɺ ��D(g��Ʃ��B"�K�m��?Zt��A�ne���|ΡW#��F��D1\�����P|ٻ��R���M������J�ֿ��$�=��#/m��_+)U�E)d�Z���W�-��p�U.�� ]��>?�P������N@�7kx^6 `�2�ZPӸEL�ҍ2]6��4�3� �*��Eq��v_Ch(o�DpϾ5���9��銪�+�x��9	4U�eCo-�f���H+Р���%u*N�|.��	����9���ڕ5�֏��v.��~Y�Y|O� �3D��$�朝�[��&%t����T��בi*�HP����ޔ�]��"��oj�"����Kר��
�p�-V���O����Z�R͡���h�8g����iΡ�>F���b�Ҟ��2E_њ<�&�R�]�Wʮһ�$�e(��]S���h�D�9�j�Qkb��k���UO���x�2�آ���|u�7�$�J10t-k��MM�x��E���F��s��@��	���ƺ��wB��VV�qh���d=A�?o�g�*��Ik���dGPC/���!j�U�u���֘����"=�c�ɗkT�ӶU)�}��k���[�h�~��ʲm�^��Q�k�h��)%P8a����#7@���2^4�ə�k�Ak�\����2��ӵ����Jݚ���~RZ//�U��n}���aN%;gV_�]�a5WT~�2u��v �!�y�b��L%�
Z���-�J.�gm�s�E��U�dU4Cue�
F���狢k�|^���_����ĳt?�1�i�shM�zU�EE�g�}�b����М�D�e>�N4%��"�4"Ul H��Х���C~8c��$n�ҰҘ��H��4XBY�L�*��˸l��񔆽����k�$�w���I)fٖ�UԄ>Z�Ֆ������n����ַ�AP���z�!�����u&|�Z�,��MZ��OO�Ae*W���������v^�N�Xc� M�y�*�m=y��\�^�B^�gK�lE����������7�H�ˮ=�
�޴ٚZ&JF����U�Rs�U,99�Uiuz��HA\��,2{�]�D��7X��,��g)r�y^��q�^����؋�A+�N2y���u��+�OV��X2�4�b��_dP+J,�2�Gu�ɲ�-����רwݯք<��dJEl��(�f�=ǹK68�&Os�|��zn�<q�zN�2��H�e�� X^e��$��Mx��>OR���,[��e�*� NT+h��'򊂰C�%Kd��l䃪�hy�:��.~��m�
��׋�M��ed���FGuS����Vo��[n	�$%:�,Ua}j�_}�9+Q��5GA�)
��F)й��2�>��(6%��K�a�Yv$�3dU_ם���D3��Z���d���"��N���_޻X�ӥ��~���KgG3��6�<��F��R�Ȧ�Q�*��F��Nz&^�VW���_�hYkFH��0!��;���ͽo�M-e܌R�Lq�ԫs\N�{��\��^�x�)_�`v_W�KI�����^̓��ǋ�}��J�ni�"�W�����ō�U���Hx
�7�)����h�j�^3�}���1�����~z���k��ŭ�F%�f3?��YP}gG���﷔���_6ISj��%�%��EFe��u�=8�M;�T�<��w�ie� qn_ ������kb�m�1�]�ޣVjqȍ��yTM�My�B�1�K����V��~�z�R��t}C��P�j=U�J�(����ͽ\�W�/�!�4d*��#JW���e�
$�2�K����z��ac��fy92z�L���U#A�:��G��k-�q��?k���4�������ȉֵ����FS�������.-���I7d�cp��Ja�X^�������R�U��}�x�%�YZq��ma1�0��/I�I7��|~{�t�+���x�j+���AB~מ@xEq���sҷ���NOw0�z^1׎{ma��u�U^^��ҥ�ʽ�Q�#�Š���_W�yi�QK$��ߠ�Q���ҽ祐Li �2FGɥZjۄ������[��eL�Ja�w�9x�=�ߋ�2�/:Y^��W��}ͱ] &y��׫�K��7?_S@5�?,�yލH����{���q�˺
����y������cq�;�MۋUr��oJ|1UU��q�H+�7�n�	(>��=�$F=��ܻ4m�xM&2��6e�eN�(Ѯ\2�Q���+���@�Y�F�u�l�c��
��C�Pq���~gޚ�+گ�ՖP�*�K�$#ueP7ϵE��t��#z�N�r�pRn��j��-ׯ�|�i�N��iI�q�DC���,��(��j
Wu��gmk��OJ��t�K_��
|�o��17ܺ��O�?U��ԕ�ac�c����JW[��hʆ�ى-���{���gv;3��ɋ+��d�Ĩ���t)=��y#��/�����d��4�NyZ��w��������l�~�W�V�*6���c����xy��:�.��MG��c�"��������|�DC��� �nĽl�(8��K��H��i��
q���D��B������eLk�ZrNe47���S���V<�3iu��p�[�v؜�P�i�\y/)�9�Tf�-����1���[t�ɷ���鳾��<-B�C��cJ����H����J}�	a"b3Wc=pcn�����N�5��y�Ϸ�^<��]�U)\�b��� ��I��7���l4$�L��eZ|���lF+鲼x���ӓ�Y�E�ͤ�0'��qU�/c��ZkL�3]iI@Eh�"Һ��@H��kG���G��e��*U�w�u|�D����Mn\�Q��u����CvX����F��[�]�Z����7eu��|���{j�G��{p�0K���ϒ��Y�"�%%�7�Z�*䋹I�L��m�޺��$6��e!���9�=�>B�[R�$O2��������_
w���_!@G����8�NK��6덲īQ���V��3ͭ�Y�Xk����m����0gX"VDx-[S,á���V�=~��/�%�4�~����"�0����2��y��V�pe�hD����gS"ͺ��x���j߅7�{�> K���W���Ÿ��|&i��Zk����X�kh��r�
����BX[Sg��1�����6)t�t�U�ǧ���� a^R���Z,�n�����g�1�c_3 �J�8\�J�͞�o�S��YQM�1ֺ�z,q�ih5���D4�O�K��l���^�I��ۍ�ܳ�lpe�~u}^��)�K�s����)m���~�jk[�������"���ꦾ;	T��E��>��ؑ��wfۓ�YL�:��egh�^5�)^�R��F����)����*�M׫kP�`�ѫ�)�S��=�{%})y�T�l��#� &����g
���żS��޷��໗�~YJq��d`	���>��L*�2�o&��������R����Шȸ`e��o:��29�Ks��� ѥ�jv7�|ټѯ	op�b�]XiԆy�\7����&m�9�$x�}�rz�q�f~�����b�`;�x��),ukŵ"��F���h�ёP�!c��n����P*K!����fl���;ۚ�^)L)�n o��M�ι����4S����H����֍F0�t��w_�!ϋ̡2�y��-�:����N�d�#iY�9�^1$6ڸdb��M�W��՚��l���3Ou���}�|����Q�\�g��L��E��Jt��hc$r�ܮx�&�;�(s��0�����XW��\�a	���=�#TGh��jP�=����k�ҥ�oelrx��Ht�Hc�y���.����Wz�6�Y�mLV��8
ٜ�,($��f8S��"j��7������fzĝR�jw��Ԟ�-�Ԣ�j]���p�iY\+� �R�U�$��n����4�����Y"�l[ht��� W�۰GVݲzSRk������
a��Om�!R��?��Ӝ=?'�cK��J6�e�]�Z1�QRY]���H�������67�f{M^Vc�[���!������(�4��)Hc�
�Kk�ϩJ-(A����>iE�5F�\/��˒������g*_�^�Ȱ��EN%�,�����;� 2�w�S`��}y;s�-�6�7�΄N�����󳿑l�Gj1��r�ʒ��ut]�I�<�l��Պ$Z�퍡�bc��EHx���M�e��v�ï]t�����y+��:v��u�n�/g�pB������E�{a�g,i�=�7�Xk�s��I��A��u��ى��,��s���^%_R���spZ$4��X�� �d�X��Ms����ׅ��bT��k(���l�]{�l\7������$<�RW'�M!�%��[ěƀ�VB>C۸��>�R[<����4��\J��4"�"A�^8���X�^�)o_���`q��>�K��m��]`�|� ]nj��zl�zA�0�hf"e;y�� ��r�1�����ID��i]�u�U�5����s��Kl�V/4G�/�vM�����y�CC�SQu�+]�<F.x�@�o_���A٘��%�1�� L�w6�5D�z:wݒ�s���"e��e����NA^w�c=M[���2v���Tq��s����s
��]�f*��5�4{6�3�l�������x����"�d3��^Ќ[뗈�_ULR[��s&zL%�0��{ܠ�������Jt��;��OW��<�qɹ�^2��&������,��r����M��Ұ�{S_[Wzj�3������z{(^�Hw Q���b�X6/�����kkmn��8�K��X�Vf�r�b�� �M�7]��j���a����0������o��{����9ц�,{�.�@Ԗu�-6AC��
�U��qI�ƆAHt�.�<G�0[Z��+��5n�����{;s��	�!J�RP�xG�X����"�}���F�Y^Ύ�;Qْ
���rWEZ�iU����oY��'u��!B��N��Kkr:(�\��K҃i�B�W!�r^���pO�*�HS���bo�a��ѧ�H4/����+(՝sܫ�.J��yM_ob�.Qcx@c X뭻l������t5�m�'ä9y�ş�,�ٔ	P�*�S!�M8�����cL_�����<�<˖�t��M��r�IY�Ɖd>��M�kd^�B<�������**ݪ}ICA�U�.۟��Y��j��B(I��H@of�U���3{�m�̅��Ѽ����=3�*��r�t�òE�2/Ky�pGˀ� cRx��p<�'�P�c�H6�pnK�����oj�]��sf�s6����o[J�Lu�8�K�I^�+?|=���B֢�S���8�.0�"��kڛ*>�6�x�z�[]\a��µ�0)c�q��=��ܦ�fQ�b1H��8���!��K��$Y�򨞓<�h��s;kz*X��fhua���|����a����z hݍ:Q)�ch�x���"���'�'e-��1���1Y��*{R��#S�6�ە���\jL�ݥl�|����U�_�Zu��dMԲ�
�(�M����a�l=�C���%��z���{�LI�SG�=2SYR(Hۖai���._]�9ؕ��/��'@|�t-JQyZ�i�����H�9%̒P�����b��BƜLD�.��Z�Ǭp&�~xbWsrl�.��#z�}���q��mtť��"�+��1����E����m�\K�䐂��v�&�j�vyHbp��o�Cʑ	$m��"�j�(��P����.�6nC(=?K��+�*�dˠb�\`[/ ��5����aРuʡ/p+j(ni�ۓq�$P[�,�k�}	ۢ����$σ�m��v����x.����l�]��`����\xs���ʐ���� ��ǹ43e���%�&nm�����@H�[�F��>�j,l����%�Y���=ۙaG��s��lɧH�IN�vE�Xc����w����Λ���"��䝊F�~�0?�.V��_���w�nh���Ҋ"uڊa�Y
&����s���ΡdC�.B�� b�R��DϧS[l3,�v�����}����y�ʥ��ue٩]9C;�d<r����TZ�i��M��r0*�3n<�y��y���f�b����\X�x/l�q��ST��,R:�[�7@�n��;�R�z-�Y5-6H����!B�F���q��2��J,K��F!��p]��u!��"<�t��,�'?w�j�����	��ZE �)���E�=Y������MTN�	p�M!��\W��LzGQ�z�k+ `�"=��t�4���ihh��fw,!Q���b���)r�{Dz x*�[�hhy1����Ev�꞉'�\�s�k�ze��`R�G���{F��{Yd�=&�U�#V1� ���mR$�,�n�H���c�*"U�G"ѪL[KD�!���i�̨�\Qָ��ue�J{���T�n����%��n�xX�m���m��j{��P��0#?/�ҍ�}`!"p����K5W8c.H�R�g
��v�s���=���I�-=��O�B�RM~R_t��ќ+�u,��ļ\��Ukq4��ثMtu�:���H)"40
���I����L�3�A����!�C�yD�~���;G2K�?��ۏ��F�*��r9["�rvis|��g�-;3�� I475�'�����LK6�г]s,76i�Z{6���/�U!�  ��t�es�?u/

㾟��X� 4_�3;t"R�06J��b��@�mٔO+� �75�s����)T�!�s�1�x��5Kl��RH��f��R�p�І�5�ܓ��� H�����r4g�	f��8�X'"=�썮ȹ/C^	�^U�5�I&e͖�ߴ��ٺ�[2�U+����Q��=�v+t�V_�9Jњ��s@��TA��n@s{_2��=1kw>Q������n�M��^B�7\C���;C�qi")tL��{���+n���J�����θ�}���e�_W�&w��V�;��LYs�Lp�2Ae�9�ݍ�WI ȯ����]c��'�P�OɆ�\B6ۢ��F�����@�C"Cs�BZ�t�S�1�-�]�'���uDS��8FC�Uxm2�d꿇@�t�x�i��1�����74�i|:�:.Mͷ�^��o˘��|n���p�\&w�^�]5���'��s����L�#��v�=A�h�j����њ�5��K��(���3�L1n0��+c�s�P��Aw�_ho)���sE������V>�,���vI�r����K�:�SO����5���o%l��*�(U)�.���0�+NSV�^U���y>[SC�1J��~W!�s�B�F6�X|�����5š�}\��GB���:�� ����Ն����� �����D�}.	J���B���k�+��ɓ��rщ�%�&�m*̃9b��w���~�,d9��M�c|���G�z��x���存[�a�J���$w!͐C�2f�<�!��R�mn�I[c@o�&�M=��j�MM���!�#y����P�JU\��̙��3_.��%�-jޒk�(�0����Los䘎Cd�w��V�2�)��:���e���3Tp�5��=����etw�o �e�(�����������N[�]_�4P��*�\��	��	���HԳĢ������H)�✂j�V^:<;-����v��Xh�Ui�����}��l�3k"�mK��?��T�)�e�UA���c#t�h�T�/*y6͞S�� ���Ꝝ/�0MFky���759�ͅhLɅ�c���:n�xKE���{�AT�XmT�h������ln%����{����$eLJ��X&�ڹ��ؼ����]��^Y�.���إ���J�6�)r�5rG�z���~]�9��m=B��{�k'�z�s���Aw�f���,)Rq��{Y��R�dF���dR�A�v!xR覕��tĵw�����^Jh�_h��ο����p�fA^[ܺP���W���96��
�z����ѝ�𪫵�\�^��,W,T3B�(�N��%�P�Ew��{\x��,�W�IlK �8��|���:])�XǷ\��=n�j.����x��eN�Q G�w��@z=����=d�z��'󱇂�z4���T�R<)�.)��=�1�Ƕ��O�cp�c����;"u��a]۞���o�D���8T�$�8�kH�5�i��k�`�c��Y���%qj�FQ��}�����~���yW���άCTy���Y�L�#��z���	���m�"ou�$G�P����<l���y�'_(RCI���I����dx	�*�W�^/�bE<WV*�qY���S�{�JCq���=����)Ф�k�Du������Nܧ�H��f��^��8.�3�?f#�ڹ�|��|�	0��̩������1��߫F�n�g��F��Q9��D}�Is��fL�c��=�z�%ⷘ���
�!JR]�@����ҫ�F�qm����1b��D71]qO�V��l�j����Wg���d���#K�4�c�m�5&Z+���>,t!i�¬qBmK�x|��1����Y��%�ϫ�4��ɝ�z�5S�m����bgr^�)��N�*���^a]���佗�<�s�����D�%<�<�<�r>>��=Q�!��Uq��xA��y���}��W�z0֌<�3~5FJ��owww����~B;C���pյ�k�H�V�Hu�k�B/%�E]��D�r��K(�����Ӫ�P�6; ��u�4�G�Zn� �B7������z��ƌ_ή �Hp]+@C��3��qQ+�+�(C#�����(��l�Ce�{U6C&�,�]hZ�=9��9ϜS���l��'^�{��D�`��v%���W���}� SҐ�M_�ێX��C'4t�I�1�5x�K��t��e8K��23���*����}�?��U�q-�.+�(E>���tU1؃����&��׬��q]��=��5u��&�>[����ZY�o&]��3�g�qoX�݌a\Na��.T��F�绹��kd�y�Ǔ)Q\w�}��]T�܀�U�{���51���q/�rQhs�Ǩ����TcU��Eϔ����z���o߆"��/�Hщ������H�G(ͻ�T�0�T��נ�&MV���-��B�븄�!Re�*�
��$��ה͝U�}�m�Ly &y�T�(f�l&%;����j���x��*O���̮�[͂.>aBE�kیA��8��=I���n��a�!j���׬�(U��4L�Ŧ;Me�8Ű���܎����O1�.w�\��N��Ѕ)����[,Ȍ#v3^�w��(/�aɰ�-a2���>P�ސ��Hz�m�T�ol^�lw.JJ���)U_����o�Q���t�p�%�Ft7$��F�jO�c��5>�쨡�}���o�r9� �(ZKMdF��*lE���/���W����"��^1_x���%;���T6%Sj�@����P)A��H.OPn�&�lc�� ϧMx����� �S����y�1Q�1����eW�:��4�W1�+!ү��zU��HG������*�|�T��2��|�po����Ѭ��l�]��N
�:ȭ���n�H$HJ�)�pY�G©ʇD;YŲx����`� 9��F�;�Y� !T��0a�վ���/����s���Q	W�ǹJ���`|�1�6��
�O	�B9��kݳZ��ω+ڝcۘ5�"�;;:�v=�x��ۛt�"���K7�簄�-o���XkQI�n��ڦ���B |����K�&�nE������?P��B��0$�O�͓��������=@í}
�|~�qu��gO��I@����C������O.����)� Kz:�R�Z1"�\5��nW��V��דL�qo��^�tVR)� Ej4,$#��=�k	c�5��óL�?]~�+Ƈ�^��Fp(6Q�4F���Ӣ��``�n����Ye�dp��㊌��G��T����(N'�B���kD���2:�����Si5��Mr�l��7%h�GE�%�v�(krJG�.n)�(�j�04b���qL���x��PY:���j��'޷��m.D�V�E�`^��r�k��f\���$Q���y(�>���:�#���M����%��j�+������Lj$J����竲#@tg�)D���M���S|6��R]����@a[
�CYt�!��~?G�M
R���aۖP�����Ɛ�]Q4cx�r���Ux_��b���	��S!���?������(����qdX�Lxx������C�^�*�+��/h?�}�|�w|����c%��/��@a�}[�odX�2i�}�+�j-�P�����q(�B B�|�A}
G�pWZe�V�L���c� %���ֽf<+���3�5��s���@�J^�<ͱM����?�����+��9�]ʺ{�޺+`1��Uf|7i�т@u#��d�>����p��!�`8��Z�K�`S��9��1Ez���u����Y֧u@�J�������u�OP��V���sK!�>o�6�@����v8h1��~p~�Nm[��i��{G�TV$�Y��T��s��M	_D��6�o�D��<)�F�;�:�9�R�����Z�����:�X�xAyZՐ��&a�qѲ'O�&G<��MO����;��W=vd����,���0k���`��h� <�C��+D_��}�k��3(Fk��"g؋e�T�DA�H|4?��W�,E�p��a���fl�������O�!\o<;�H
�
�������d�C�2\w��$�}Ng_�K̞�KYO/=��v��-ۍ�%�o-�|�3�٠κ��&�U ]�H���T�^oV.�����w�T�Z{'���э��u�`H������(�!�)��JK��!�#
��U.XZ�}�D���lbpbL��ͧ��
��YdW/h3,�M�����m��,�fc�m����f�Bg�f�֑�hV<Ks��8�g "�*����2�ٝ�@!���}_?�/�g�ޞ=���Z��N��\_�K�i�3K��su��nf���I���*�(���>~����8�K'
�.��~K�yrJ(H�E\��ӎ��ŸK7R�GgF�O1�H��M��n�uE,�%���C.����>/`x�(ҡd��kk�5B�"�k,�a�ǻ0�;SJ�Xxl�������Xo�O�S?G�ʞ���p���9���aP��H��7�<��-F���
���9v�7�QB%��֩9�Ԃ�4#��IB��I{ck�ϐƧ��l�c��d���2����o�1Y2����<"Ż�ץ��Ɗ�b&�Vy� 7�;��mK��P��֤-��Q��ʳ#����l7S���~$�"8�EKcq�7o͊���/�Ç�� �! L���ú���u �ie����-f�>.N8.� �	eZ���72��8�ֳ5O��CQɝ�畕U�a*YF\삟g��,m�B�7���C�mm��P�_�8��*N�%>�]Y�u�M�>w���ڻ�6��8���Ap�3�������H<��Gs��Ї�7eb@�C���z2�~�����qëJ���m5ȎE�2�Lp�r�^z��/Śm����ؒ�'W�N�ꕃ8�������z>����yK7�d��̦˃!
$�0d��1���OxU5���dU.���`�����������N��a�k������c�/�fgc���b�8� %@��}��ݭ��$O�a��B��/	�L���0�x�W E���>⭶V�g��A�`�ݛ�!����G�� �9����h�����
��� e$�2]bB7�c��!d�E��\�K(RQ+4xh@������&��Ӌ-@e��^E�������;���������O?��aU�o�e���⋙�/W��>z&�q2�"����׊
�:��4�B��g+��ȑ*��PR������z|�R��(�`A�Į��U�U���x�/�VxV�Ʃ�%�"�٭�[����	��(Ct{�r	�3�(�#�Z�0`.1�_}�U(Q"���z���.����)�sO�����ɲ�9f��yȤژ�NX���=�JXA1z�nq��+�j�?;��U���ܖbZ1�Ȓ�*�]��ݻw�8ܵ�����==�s0��oq�+�����u��B�����۷�L�`�t@�1�R��)y�2���䝡�J��.(�O�?۽���9`}f��0oQa8��*�;�0�b���gH�����c��axA�W�Ŵ�aݽ����->��a� �Hq�Cҝ �"���m��5�>����_���҉q��1?��<$�ب�N[
��R�z��@ִ)��+Þ�0T�	<&�eL7�����Í�����}�bj��"iqCh!X�����}�ȸ��?��~���U����:�m��Y�T���?��zC�#�	����}�����r��ŬiA�������f��ȖYu�٠�!�N��`��ΐ����u��ݝŸX�ؑ�\I� p�0,���(�����X�oL�qNSP��N1��ި�()��1@�7���7��u������Psko޾1񹽿I��hڊU��@�٨M%���� �wͶ�н)>j-�J��>����גަ��uL�"F\�iUr�;��#���R��`,a�/��~�~0y�}��dTن��V%�*b&�pN(�Z�Fo�{��a]g��=RZ�9q����?������w�f�>����O��fw����\� b��,�
�3�B�\���<=��)f�;���B��sךԪ]d�eH�H������C"��B6�|tgi\�Ǉ��K�p�<����� E�gȀ��q˴�}�"w��T��_*�Ɠ#>=�-��%�+�آ��1& (D��~����cRޯH ��& �t,��@�*`���5�B�z3�+
������kQ_Y%�d�\z��ص.�㰉äU=D#c�?�*�A���4���.��!㞮�`��-�.XkYE��ňq2tW�M*�P�&fWVo^����U�~5��sB��\�)�Y�	�\-CӗP(X���/#��
(��=V�!�`c"�ǖjO>_��~Θ鲄��Y�Z==>��y
�����BNl�q�}�,t�h;�9!o?���B�����*@q@[�y�e&;�qQ(c���c��V@����_���8�5���e���ƓR���JJp�Q��Z��}(XR劜	>�d}ǳ?����w �{Ý/b�Q�F�� ��1'��ޮ����2T2�8�J���u2�S�Y���$Ӣ�;��c_"��&ܕ��_���+����"�[)R�0�䉩�\ɬ���b!�_~��·�;����_�$�3h��h�,Ѓ��:���^�����tr������O�����D�Τ|Q�N��Hҟ��)K�!��{��e���\���L�nDD��@]�p>XnX��*#:y�c((.�Y��`���U�]q+{�C#��+:��v?�����f��/��b����=��Y2k��^@xP���Y��"D��)b�ճxa���S�	M��Uqb3	V�A6��ע�=vW�B�{��������x�XJLW�6@COD�0^S0f{6�H�ҭ���dn��H�����^^:����$�Z��E^d��ԕ4$*{܋2�_���3��p �Sb��IԻ"�=e�����/�����㺗�\�lМ�%�)�Q9S�0����'e��(;U!,� �CZ7f ��*(}�-&+�x�i:o�Z2V��-M+Y&u���4,��Ev��FN�'-�V5��H�>;�>���oG%�P�ל�>�B9�_���0��Z\jU�O+�� �e���Dd�po�(L�ϨD:y���*P��x/��a�(����Ǘ��?!���!N"�[��f@_��]i���bx��ɔ���NP>.�'�.�D���l͓v����VK��X�h9BpS1F�ɡA0b�pOE��k9"4�s?8�i�1�\���}�[��5~⚘�_?��I�3㭗S�$j��ӟ�������2Er��UiT&�x�������:�ό/����qFk�$�EF�rV|�P�}^���7_[�U+J�a,q~��-~?M.sR��-VO�x��w����b������c�]�ڳA��2���ra��`��E~�uv}�A͈�;���[����x���ft��޽�sclqN��Q��'w�l���ΏO����0��bxG2>�(n�0ח_2��@%��ט7��Ֆ�%	*���R��֝3L������4�8���P��e���[-DԲ��t��
��㺴S��f�'��&GJUu����K�,.�ɂ����O�?�Ы�$�2�l�ᦉ/)�عP��s�H�͒3�-���N��U��i�ЛE$IX|��T>,i�!�0/,��.�=\��YH�>;�D4���r�ĉ$��K�O�z�}(1���d¤$����|q�'^#���{�gWlcS)#P'��-�@�X��o�ǧ���̅"Z��[^	k�v_Gk��p�$mjQS����������q�~?�_�r>�5���J�$s.���q��:���nYcs�QJg�b�����mF�1g��4R�GM�Ϙ��Fơ`�[��a��bA�2�<Df�	pL�L�&�wβ����=V�?D�&�R�Ԣ�nF�����P�%E�g���Z�����K��8�;c�-in�ښ�t�
�\!nz���� ���(�B�Cܧ�қjʍn�W?K!����o���o�ұ�p�����y6�X�z�ÇP8�Bt=n�}+;E�熙^�Z���9�l�19۹p�Ϫ��0����7���_�/�6�z涮��	4ג�X�rQ��W0��U�}�d�6�e��㧾��n��@���/���EĹT�1zW"�_�ɛ��� ����E�R�_�J�/&�ޘ�5OǷ��zk"�����)N%���U�S)|t'�����a\��B�??�4?N����a}�>�}"�� �D����,s}�.5b�G�ĵ,��x�]��-t4�w���++�U�CC@�?�����&Vٱ"3�'�!|VqE+-������(����!}�?x!���d��X>�<���@�h�U>���y��J$}����L���ɾ�q?�ThG�n�M�2ݬ�QZ6}&�E^����u�$އƩ�I7�d���N�¸4/!d��h����&b,l}������E�].5~V���&�6&�+�T֚��v+����s[|n�W�b��TRQ��57�¿q��R`�k��!�'���<0㈸��$�){��!�$f/��� ����AA�-���ظ�Ȟkﮈ)R�p/�qYk��=,c�5�G���%�0w������?��?V�D+[��,r��']F`[����;�t���&� a	e!�Y��q�[|4��Dɖ=8�_Q50R�~���=���Od5|��l_�n>�A�ӳ+u�ÆDuw��`0VV��9�8[�u�����z����c�{"�m{�Nɘl�Ȯe��1����@ō���F'2��Po�CR$)UY'�ϡP�%㼃�JHE�V�^�)J�UNL�|狖�U�^��!I�ǋqM���\���1"�#�?���a��g����M[޸�PHt�W�@�̙�Fw���Ժ����
�����(��¨W���J�J���l�R�{r	庶W����БYt���JU���z�v������(�m��Z��BTQ�X?OCS̧�#�f�{/%�b=�<`�pb���&��!+q<d ^�-e�H��4^�/��dUѝ�%�P1�������4
����;xv����qa(��S���p���Ѹ� ����/vN�O�A�B�H~�b���Ѕ���;RCF�w�F������PƔ��)�8�=�K4O.� ��RoW��X(�����n���7\w�Kܻ�ʍ�o�>b�1�k�BZ���]�4�;�A� n6?<��~��_}n���sɤ3��?�����;G�^=�F��crO� ˅n���GK��E}0�D/������|ë�X�1��s��x|^߿u����.�1K(D<��t�iwWy�Rj"�l�W����]����gCų�8��í#��� ����x�i�<_���*�*���_�2�����ӯT��|�Z����{[����I�W����z:U)r߸��6��o�=�y@�5BrB�f��� ֊�h�~d��Wq�8�z������K�����^��'i��� �L7ۚo�����A��h�H�sܜ2�p��#ӣH���/�;���5����u�.�E,<罻�8�n.H�ѳ����ӝ�K`(,���!�q�/�Z@%��|������X5�OO>��%�K�4ј�9�#֌�f�b6Z���p�T�\t��;�v��@�
��.��<�J����I���Qߠ#���b`���Z,�m�'Ɗ�E
c(�L�?�6�￰��0Ηܱ����5�ŀ�;�;��<�G�ޟ�Cx5�^b� s�q)�:}7R<�(F�ųܘK�9�����-d�l,[��0:�R��Ce�����O&�޷&˻�bޛ�	o
��=�հ%�3׷��)���UER��5�u�M���=��k�i�2Z�P����µ�aD1366Jo�k�g���P�t��\܇���R5k_u[(ّF#��Ͷ�^�������׌U[��+�7���XE�Y�Le(�8[����[۰Յ{{��
�	��n�ܯ��u��h�CZ~|F.&GM(�U��;/����b�X<AYq�kX�����?9O�C�)N��d��a,���3����,���ǟ��M�-�r����o8f�`q>a<�����L|p��vz(R�8�Tԗ)b����|�8����}祧�JX�tq��������w.�%�<>�4U�]� =�1�
k@f�[x�x_.w�0bE��yX��\��q�#|D~{($ݷ5M�g-�h��k��`���.�'w�ob�����#	�d1�=r�d��b��TǑ(h �Ǩg!�M$��2Wfh�N.�S�|��Iw6�"��qB<�Ь.e�ay3j�S]W��ɥE�X��m5_p�P�d@�t��#�W����.0���9n�W��BJdg�^��ւn՛�fX��ǿ�����3\����78�����]7^��h�=g�䩹��0�${�`KT�s퉨��l�6fBp��q�~�7���-�ƞ�B��g6�I4>�7������ x��g>쐈t5��.��z�J�� N���Q����$Q������ZRN�!z@��om�￶���ovO�|�M��߶/��2j���^X����F�R'%� <�0����-h��f����H´�n�8��{���)Qܳ�9]*U���CW��O?�+��=�iݭ�:,�/V"()k�] �A<�{w�(�ÝO*�B��b���r����Q����φ�n{�c�M&9.2l/<�[���yrw���S�N��u�q�莻S{�?9.�Oœ�G��'ƣ��\#ɉD����M�W������sd�3�Z�S�_��o��e�"����T�j��ܑ��F����8�4�zw��Fz�ɴq��':O�}�0�^֌y�(�)ۄT4�$ܹ��&Ej���J}�q}�R�����mA��� O'�K�AW�Gj�����|���"-٤���-S���+Z��Tk�a�ٶ n<l��N���#�-l�*�C��	 Z�F���P�Bj��)���8��7��3n��Eh�5lv�Q���M@��j��cq��Y	T�xR����.�:�Db����>3��v9��7`Q��,��r�������z0d&/沙�u��๕>���˷7�����Dm��deеg��ήO��4#/N�qҹ��aάф�8����l�c������'��2cG����2w0d�}#�|WE��?Ի�;*�Q�_�,2&��s�)�y�|�Pu��D�/xc��0�}G-N��&&� ;���"o�vc��G�X�'� �6�B"@@ٳ��nrS���W	Y�}�FB��B	�]�K�j�U���L O�������;���ͳ�6� q��*A�6��x啌Lm�r�<u<�RURsm����I�I+�擇�����H7�'����3��J`Z�%MN��1 ��{� "�n�*D$���I�V���������d�ѫ_p?IE��frHI�WuI��)w+ȘX
��3�����YՅ����n�:v@�����i
��w�sq�\4 P��L���u��ۼ���S�p�����1n�S�쁬��W%(�V�8N��aR�[裓�w{�b�'���t��T0�\Gۣʹ��-��j!���ͳ�֚�%��?������O?�x��\ͺ�xp]�U�=*qZ����%l1�[�>�ʠ�!���ҍ<d��<8'��x����U���a*Ҩ�h\����aI�dN.kU�2DH�⹕������-�g9�6�S���L�>��ZW��W��{�� ��17�ߋ���%/R�L�ђ�5���*o�yBV��Œ8�|=��γ����"��Wyj�ㅱ�a�=��S
��!C�,�?a���u�����5�4������g������&Nq���أ5����}Z�#Ăb36׊!��-w�dFRM�] }��C�$��M����U����4��v���^	�0h˒ƶ|��A�R�j�JU'Y��gO>d�]���4��N,�V�1#Q���Y�g|H��X��a�3���?������	b���|3w��ث�njj��K���4�ME�Ɔ��Ο�1�;e޽���cg�R�����K��뼖$Y�Ż��_��T#o(0>zl�}�]`����@lϬd����ў�|~::0IԠ��N�y��%9	�����z�=o,��t{��^����2�09��w��2]X~VJ����;{숌��'�5妑��T���:5�b{V_m7�����(�g�;*4UF�����M����8�}�`ct�a!R)]�c��a�����`�P�ry{���QT�E4��'B�0��Rk��cc-������?Y�<��zz��T�+�z(dﵲ%��=��4���������ɃЁH/9a�X����(9�w�&,p�q��0| pVYuv!JƮ�ޭ:(W�7�������ˋň{#!y���5G�S<+���gM��i�*	���ؓu�Iޞ,���C���{���Ǫ����5��gvɹ��l�i+l�H�w�kp�����j���m\��%{����)�⻉^"֊��D<m�(�%����ԃU-���&җ��ϐ�{�x���H�v�
�#)D\|0~�7���?�bW9*��_}eJ]����#x� ��$�->��-�&����(HGn ����m,������|cq�/�� i_Cd���k��3�qk�Y�Cdtq����#�"Z�!�er�L��yt���ݳo�A~um�&D������-5���gӴXǸg�2vIER�d�|2�Q#n�>�"U�}��?��"��8�O��",�)��m�Ⰻ����?c��+��"��������1;�yM��"��q`�KR[�'<RG��[AsYz��j~7�(��J���ܵaZ& v�s衆��Y��W9��ذ���a�����vAL�߾��<Z�f���m8�Ư��s�.�/^��^h�;?jk�1�x
����'�1p���;�֒]�G��8��1�jP58��j�������
���H��t��i��m|Zw��q�j�k�](s2�[� �J(������5�}R�D�!GQ��T���N[hfU�@�
����s�S���DCOA�"+� ȇ���s�}��,�����Vu���]��Ũ����K�I&d���}(`�-n��l�U�L���~�bƌٗT-�Ы���ØՂ
��QUD7��>E������<�\�"c�bO�2���F��Ѝ{b�O<�m�Ε������s\_� �E
IK�h������R�ݷ�{�~lbOZ��=���{���s�RhT%���.���K�|��E�������X��
�Nd�2���-�z|�"�B7�?o_�Ba�)�j�W(N�����Nŧ�E�+R�]�����_عH������+L�8 .�sxVeNVH� �9�hIIT@�5)s��Ʌ"���{�P�+�vp5���jy�ث>=>:!�%�f�NL�(�����ʀ4�[�����؆xOTH^ Q-��'G����w�/Z��H\$WS�����He��VE
��T�yTB}r%�geOT��=���"�g����zlA�m5���bq��g�?������HَRк���5�d���66�BIȷ���Ǫ���L�X��i*L��o���O9'R���]po���̿5����s&r������T��<\��L�O쎛��fU69�f�c��*�OM{!�+Jz�'��h�^��[M�.S(:��Crn��5h|Kq���t{씱��#�T�W�JC/�����Cª��	�-p&��~~t�p�&�'�"ǝ*:Xc�N��j�V/�G
�����s�b>XsƇX�C�K(;�C��h�����sW����t�Ϧ���	h"�^��ݞ���!/ >����`qP�����wW�(q�l~¹ =��	���߿��ד�]�e}�~�w�}�!�7�cB��	��Ǭ)���Q�σNN�����wZ�e��^K(�RA ��!]k=�������������g����P�k�7ǵU1d{�Y�"�C��A5�wN�BÂe/�m(F�(�ڄ� t��� &�D7��ʤ��˄�y�Pj� ]
�V6�`Ƶ����A��?����?�Lַ
6C��m�E�S(,�{8I��M(�~\��o�Ka�JV���"�``��7� �H�׃��5��ό�����4pڠS'�9��  �vN�ސl�n���]���{���hz���)
)6G���D�2յ�A�W��Fl�#�='��Y�F�\���KK�jY��iN�ڻ�����Ҵq	J�-��@{.��=�Xoqͳ[E}E�Z�E�]i�g�E`=�����B(�R`P+ƭ���'������V�)�e�C�j*��1�5�HX¹��˟-�޽p��._������S gܯzEVt"!�g �#���Z��q`I��ʬ;�cqw.d�Q/c��@Y��⮐��	��{��45ߖ[�0���U�M�}������+��"����&[�E�Ě�\)*{,φ[��T�Z =׏^�k��ֈ<���C2{m}��u֖�ֿ�6�U�]$�{$�$i�]d=�9OsY۪p�^'�@a�)���P w;e�S'I^�%��#7?�,��h2.h|..��ȴuL��^e�C�����V��<�ZH�q���潗�k�F��H��Ԥ�<�y��������G��('���}{��	�{����n �	�:��uڅ��{�/�ϵ��>糺m�2BC\����	�����X�FT%�H�ݵ���'*����G��1y������b ���^U%�J�.R[T"R�ڜ���n/�k���j�T��������w^4�[�MZ�sR|�����6�~5R���ف��ڳ�f�Zm��?�2�uѪ��dfR��9���Zat�\�}�_�80Q>w�?���v��L˵��T^��r\�==*g��'L�AZ��W14$��J�1��֤��9��-����O0.��!7�H!㪤���8"kE+N��y�jZ��,.��*��H +�=��=���`�6���i�LŊ&�ٶ����y��r�Ϟ2*�J�U�ܝ+Mzd�J����X��ݓ����+ � m�'��J��k%�Z�t�T�?	������'z��'��r1�$��J�$�'��|!^&�X��=�ҶRM_�t����)��g���r�-���}����@����|���
:D��	�QPO|y�n����Hd�JAYB(����*�Z
|K��9�dA���BS������51��{�c1���,��P����-��`
Jt'�%*/M����@d����N���}��ح��bc�ڹ�����qKCesnu��R'�o����سqLl?��S��BruC��a�8V�әat�TSe��8�_z	�nv]G�\�+dB�f��V=���0оS�N�]�Ձ��K���0�J����N�U<��#2�7^֊Ј�ܠ�_����xm7_�� M�4b����{��ِ��!��㆕)������NM޲GK\� '7^�$�2�]��?�Ǐ,�Ѧ�*)_Zҿ*\^�|�@_K4m~�(�Х��*m���	�T����bp{Q�Bc�Ȋ���g{���pa���C}�7N��y� �H>��0�
�b����q�����2ˌ����[�ekNoai�ު���@�����v�ɰ��S�n��w�r�1���
��i�� �Jj��e˺�{�l4����wn�+� �]�n�l�.�ώ=��nn��T��uj��]'�]^����=�.�� $����+�	]ԕ�K�ݾ-W.��}��L����4�
��}{���'n��h��s(Ѥ���n��#���}|fS�;�j�'C[�R(���9�-$�b��H���FƵz�~���j[����6���{K��2gm��x/4��%b��LGW��)����8i����)�S}ie�d���j��Y���1~�<��S��G�q*�)�)Dz:=�:�U���6�1�ρ~�ǣE�m�\�XS`��dU[�HCq��_D�5,���Yd�8!�ɗԾ�j�M��b�u�ܓ/(5�9̒C�A����n�*��"p��oCv����l���j�E� W3���6B�3�%���O�l�yu�0Hn�Y��(��N�i�a�R-����%�h_���" �s��.<`$52t���F-��� .�{��)'KRA��V#O�	�XUKM�HW�=�#v%E�k����{d��5 �9D�
D:����y�f�էS�'� ���7��?����K
�:&�L:�#�[&~��'����>DR���x����ܳ���D��|��/�\y*c)�F4,���$��tk�X߈9��8���mv&g�+ �h[O��<�W��S�C*�ը��]6��{���۷I�R�P��0�PҊ����D�*��M)y�:����pQ]Ĭ������"���i�F1[=����jK#{&o���>�i���{J������ ����4㣆|<�i�<)��߹������jYm��n/*%����QZ��{�+�s�
�����3�e|��d�IǸs�򥡺G��l ��g�EH�j�P�v�e����5~U�b�¥=F��g*��+Ɠ3��=G/�gS����w�{����~�IƗ�D�w�ΓY��I{8Y����
NYnm-����u�d(�'oF��BJ.��o��Y�8ȅ���	���:�iC��pҞR�'wpXA�/B��L��W��ʘ�$�ԗ%WKha��$r�u#��IݤQͮa��R�������
�eb�� *�98��s�=`\l���q��W���Y��Do���'���D��:.��(([_���QZ[A��{�
���Iq́ܩ\� 3�<�nb/��	@������ѥ,{���(g�*���Ԏq�{�-S����g��Sŀ.	z�h�-���<�3DD�s$�ΗdU��/e裄���z�t�_|�����ض��"Rf�TO�O����<�{v�����9��V&MJR������b;/sRu#��m |��@1�P����)��&�{����@�r5ɰph���ѧ+ў[1Hq�b�2��
����γ]�W�L��ۃ]R��� �������G�.F8� �ݶaq�|��l�|�#R�Z0\��׃#��Qaa�U+X��ַ�\� P�bU��6�I��ӈ���V����UH�11%�|Yj��?��A��R��b^���/M��]_q�Gߙ�6����h���q˗��A����z����������پ�
9\��3�a �"VW "�k>ll���}���#KZ!H� &l��>&�*�J�� �����a�����>�.hj�Y�:*K?�T�R���4vv��U�_X��F\�!��/�#�X�l�$Y5��ۺ4��Ge!3���f}��U'��������
��K6��ի������Uw��>�8N�M{d\E�]
�h�JxH�rO�n5��:�	�\?�͔���ל�
S �˩�ߙb) ���g�7�>d狄�yur��\�l[6[�$��BoR¤*x�s���j�x� �z3ܘ�1��^t��i�P���^s�nqځ;��(�����-[d�Η���|�>�*ە��-w�\5Q�<q7��9����	�y͋E(BP��w����	�w�|�R��������Yq0�MZ�y>���y���B�9�g5�8E�����qÝ��]p�Iyr�~
�h
e*9���xY;>6�:K�q��5h>x¤mb�эi69���n8i��IQU�	E�Eݎr�81�Ѯ���� �v�G��.�వ�xd�r�����)��<��%�!w��=�d���M��.��BN=�szfY�IN���ʧ\/���:��]��?6d�*p%@���D!R,�h��S�pO^�� ��]�"���g�x��P���8�Bʾ5�x]|�7�F�H�"�J�[���ܴ�Z�ظ���@X�5��-�RI�6�{�4�%�;\���7��Ƚ~�W당"�7��$� ��Zu1��]�U�C=h�o�o͞���TՊ��}����g����0+L�mev�i�<�W�xR�B����W��dwܒb=-��ޥ��w��u�0\����z|T��y��[Pdܛ��PZIR���D�\�0��ה�����#]�bE&�ٷ|&�<�@� M�L��S��ڸi*'e���Z�A�ùŕ���*�N]�Ll�f�V ��)1�Z���竚M�j��ŸY����'c��Ԏ9�u�K�UW(�%&��`;G��ϩP:?��wＤ����hZ4@b-n$$;��f����b��W��e9���O;�׌��o8���Go�|�&��D�T�J��^z�K��dm�����%m�=b����Y��A6��$xs�#��`�H�b	P��S�5�����!>�~�ۤ�''�ʲ��~.{o+&�d��8V��
\�����2�
�3ÙƤ�"7Q�Ce���(YP�߬J�޾��}X]Y	s�VntT��Nʕ7��^��ۣ�F�p+�]~2�/���������n��J���h���$q:R��?��3����D�"5>+*����(Q�yts��W�~~���~�k��G���㻦u��]r�+kB��Ç�gH�iPM��8uo���W�Mff��2f��f�0ؒ_�Tx�����}�si�YV�A������Θ,�l��ی;+���~�9�⦪2N������U��}-�1T�F[؟��8��̃ws��z�nĨ5�	���܂=���k�6n<���՗X�Qy�HO�ܽ�Q#�H��?����/ވ��)Zұ�F�TS?���_=~�־_!�q�mH�^L�77��~��%����95E���g��ҍI�WqX��L���ɮY��}�mr�e!]�}��=:���$w�[�~0tc� KoM-�_�h�Z�Zf�r"���ӟ�d�tn���u���EcB"��qS7z,j���÷�rq�S�*$?��C�n�>�0�g��C��/��x���c[�����s"CR��{��-ka�	JV16.b�Sj�}�h��@�b���u��Vp�R]KD�$��%���A�B��������%c��ۏ?N�̈os{��T�y����=��^�l���e��0nvHn(� [;�D7�d������%�J7�j��%K�� 0T�{@�0C��=C�����o��u�0c����9��7ߌ�/��j��'O4���)�+�v�9��E�����,����� !~p�g̞�,��Ay��l��[���%x��/��;ǵ��N�``���������o�7[�?$b� �B�o19���o�F��ʔJ�w�朊����t��>gB��q��p�� �Ɓ3���GGi��`i��S_��~>��]�={v���Rz�������8�X�� �`�:�/J�g��h�>&R�� Bc�VёVNn'�d�M٠�C��+�"� kQ��<zB#��aW�O���1ceJP�[��R��'�vu�fŨ'Kk�!� e���#$ג�烳�L� e!a�՗�*���%����@Y��+��˿�����{n���s�'t��|�|�-�|O���B۲h+	.T���6��n>y;�v�jȣ�]7���v���e��+T$z3���,��[�(qn0x4���õ����]Bi�H9�������
�Ϧ�w���θaRV!�������Y���c>�Jp�N*�V�G�A�Xz���z�#�!����q}Əv�`�b����"�1<���<iǈ,M�-=�Z|�[��k��?��>�L����Dh��wr"��♗�ƙ�"KHɝ�����Q�'��a_��R���`�G��k^�J���[�V1)���"��sdH���)�@,�\���b��?H�$5İ$Ѫ|��p�����pr4�T��\!����b��:J��P$8��K@��zA��>�q>� ���s�KxȽ����b|��ch{����d�D>�5�W_~e�Ol	ۖ���8�6�����{R�*J��F���a�^N���������c,���:�JV��I���=����*��R�K���bIhW�q�Ap:�{���T��yWiq�m=��֛[��]��/I���u����)^��]�����8�*�Xi%Y8�A��x��;o;�|��L�g��_�k�q���EIRS����nY(P)׀8�
�T}�~�d2x��ų����	kGr���1ҪP������mE�l�QWqQO�]���"��L�v�-�yX�K�؏i/���pqe:9R�L��1A��)`�"*Ū���Q���UҶ �)Rc����6s�=t��cr����������^}�)�Z.8{�Ԓg>��U��@�����.>����&g��0j�bX���;���1�=Q�:$1S:�1���}�?'������`���*-$6�^�.��?X#�'�!9c���kـˎ�����JV'a쭦�_�U�O|��Q��V�"��T�K	-*�l�A%�{��k8��������b藡�7��[��ۦ�)f����Z�����8B[P�7^j��v��v�KŮ�Q��L=y�喸WŢ1��E�3�@�)c��Å���8���+Cow��<��>;<������GשOG�pA>(��x�R>C9�32��]鷰���U��h�*�w��K��Z�9b�b������F������Wh����te(�W�����i��;1y+�i��+�����[�O�J�ҥT�BE�*�&q�98�`E��ܨG��+s/0M����@��T��~ٗ2K��E��O5����K��n�E�ͬ�[` fY3HO��'�?�X��!�2�2��9>�7�5W)��C[��Sr��ңR�:�{]��Ѳ�H�=#�j|�U�Ɲ��؍���ֲ�B����;:�1�O�R�9<���͹Yq4��`Ht��Ð�n.��<���jՙ�-ʋE�Y��,��P�Ns���k��c8G(5�?�Gۢ��P���ߣѼ��m��O������*��e��[�#O���]�)e��E>nr���q���# Ej
?Ш���^�6O��u�v+�a�\�U�"	՗�~g9�a�V79%K(�*�<dH�{^��w|���h��P���������:|���W1��Q����@�R�ኈ͙�Lڟ�Af��-A���q��)X�9�~��R�r��*p�L��p���C;�;m��U JV�^�%�Q���%������MĻ�Yz5f>���z�/� ~�(���P���u�4")s�u�|{(a�  T�8�����a�ϛUa��>�+	Ξ]����}��nV��#V���5���?��ܬ��̕���'�\-�d3폎Ȳ�E���NO(fp�����[�����
�P��bØ!��P@�8��K�\����JF�KW&8��њ0�^��]�Γ��<��Uf*A�k�v���)Yy���s6�|}��Ɓ�6������5�A>>�����Z�b�����B�{��tt�0�
�p>�;˖q����j2��Z�d	��~�������	���	F �x!ݰA�vC����H��c����N���6_���{-I��X4R�h10P��������9���.䈞��n���{d@y��+��-��"#\����CVބd�ucC�y,��"���
�~	�T;8l�ʭP�@���n���7�wU���s������;Rr��*�j���q��G��T��ʽcHJ뭺^Ê�ѣG��PĠ�*�����4F����J�q����!�� p��m�*�Q���<6;��xԠ>:qj�ٍ�62�7���smVR��)C�X�1,��n(��<ݾ��n!�LG��P�w��<���s=b���0��/����ĺ��+5���̆{�f�uB�vu&}�x��59W��:��YP���4�) K�+}��e���vE�g�e^�,���?�-�w���y�ggZ.f ~"���\A(6�-�p���m���k���I+b�(Mڧ&��T�4 �5ıu�1l..���dbmHպ-N����9�̴>���u���9M��Z���Vq{q���|�8v�L���ƀ��pQ��K���z�:��}��0œ1��ºN��"�k�Y�d�9�S�4���UE��`�3%�'�`�J���:j� �C�C<���O#�U1V
���MI��hʨ�HiZ���������_y^U0�U�6��=��=�h�`�oN���p0��H��} ��hs��>hkEu*�0Ћ��ƵPt�4�9*���MJҖ�U����
t^ܢB��E C�ej�=S���?+�<�FR��#��p����A�6��Mq�ap�_�n���)ֆ{HJEX�y��Cj��&��6e`5�0���z+.��/o���=4:��@�^��,�.�
=�1M�|L���g��;��i��Z ΒP�Gp�Tjb%]s��w�K��1�o@1X3��z��jU�a�m~�n���-��BP˧}��К+���@8�k��� �t�8��{@�HƔ����A�zE6A	ni+c&'f�If����ڟ?�ؠ.�ݍ5ej���j�{��xO�Q��M��G����h�MA�x=�T[�J�������C��)('W��0\�#�QDki�J�O�ll��h}L@m� f�gN��a�B�5��cn����߃�l��@|u�
�c���_��mӖ�+xh��`E��i�^�ާw�Ao�>G�4^���9q����-�mU��J���~�ņ��FuV��qzcNTb,�L8����?cx^�Kt��}ZK��Na�tu��
KbY BP1����
A�:�T]5�"/�.NS!��Z�z�8�d�c�r"�Y-����k^�z'<��w�;�)`�0D�T�G}�N�.?��|≭�Q�3zԝh0�I��Y���ĵԓ T=�!�uX�#�G� �Ǣ�1*LB���ɣG�n&�F�E�/�G���S��Q����C�TY+� l������4��+���g���`3~�7���=�,�L���iU��0ҍ��_�����Ya���T�����U�u#o�d�v�jդY���� C]޹��j�v�a����Ӏ9���͡���-�9�`>��W� ^\m\�<��W`�vpgbauT����-�� ��[q\�Z���ɉ�x���������]D��˜��WB�o�k�ޑ�t�b�Q�<P�g]C^,�6�E]f�4�[��*����_
U�WWջ��H(FF��S9$ba�}I)6F&R�ד�5�|I*7�W'��8�m9I�m��}�a��CM��zN�->��h��&��*Zu��a���W����:4�)����]~�	��D��afW!"1s�%՝�$��}���^���k�ixG_mXl���5�oyF�P�4L��_~a�x0"��o=K�C0��̏i��Y��d�CFU:�xd1��k�qC���a�^$T����1d'$�~���{��Y\J�<R�%�b��Ҕ�?4��`��R0��fS������7�8I���$GRI�\�L�,D���vE;p{�/���:g��L���4oyb�{�ݨ�I<���ͨ	}��\���dl����k�\mH�UO�t7�=��js}\�.[��q4����F��OKl^9��ذ&g�R�Ѥ� �g?��$�1#��z��w��0����R\�*�#�^����w�s�#�8�^���8��tn��
�����6	�����ӏ?��C!��([F]:8�voס�}�
���9�W�m}`�t�,�D�h��TvU�Z_S�4Y{H�^㚳�2��Q%G��ϗTZ�]�pxi�P�f��Q����H
��pASC�&�J�����^G���������j�<K�ZعK�q����������8p�.�>���M$�ڴ���d�(Sb-�f�ܚ�^��~�)���/��Ž��Έ��1�*$ݖ�����K��U�����zU`���Uk'�*]�`����&BE"E}9��#I�>���=<OUٍA\��#b��=�bb(n�R��[�jP;�~�	5�a ���<.��t���0�{�)�2ڼ���u"�,/�6Z�3!�*���\0cZD�� �R�������{��*P���ȩ7�\	g8T ~+~�V�_+J4��&��8�Z�6���k��gvms�鲑��gN
T��46���6��˲`(zW��j���-�>��1(r:���v�S��D>2�$��&f�4~[�LC�8�E��K�ӤHuڅ%�X҃��P��9�<������g��x�%'\��WӦ��Rc�T�*̓$�����Ȗ�l�
�D�+�k��F�T�)���f����s����s�Q��e�5����j�K\CP>���~i<��,l�q�ya�7��b�8Z���"�ش�!�q���ru��X�乥A0�B_�I�P��w�ͨ
�TbGj:=���#e헟�t��я��S)�j�������k���	�"�wE��?��Z�%Z[O�Γd���;��yZi*:H]O9�^�!�;+���y�L@�aH.�qrq������gp�p��yx�0��)/� Js|�r$G��1#�ya�M�'�)��DID�������sL�,Muj/.��M�7mD4���:~ľ���M�3@���6���R`�˳�XSv�D�(�54��*�hZ*�r�&V�L���,(�sV�+*��j��:��"o���#%\1Gڟ�z��%��a�Kk$zsD%gk)b'�����χ��|<�H��,�&��'��Uc�T;=���6���`v�C;|�қS>{*�����t�}���>ֽ,J�(nں�,r�#̨�Ћ7�)#REWaPeL�FH�������û�$ȫ`��eC�7a���Ts�\�ү�������u�o<I��#�`̔ɣ!}i��ژ��C'e�Ee/�}�3�n��x�p5�)��#�!m9qxaX�@� �:��$�3�=Z&~)��1��9�at��0g�n�5�>{�!i�*R����{�*�]��V��������Xd�-����4d�ԊYҐ.7s����r��s��M������߼yW޽{���n�v;�1����U`����d�ؤc����o�]2s�c�PBЃQ�a��G���M��P�}���U�KU�sy��^�2��R8��9=9��&��ޏ�M���u����n�=�r�4�D�7=���!՞Qg�0S�O�{�1O�!"�B!iq�YP���������{
��2x8O`��ɑ��l��g��=�E!�z�M�~������fF��!T3�m���)�B-���<�1�T���)<g�S{Yc�Ve�n%ߐؘS:QMS�G�uӴE��w0��YSc s�D��OEP,��ż#�$��	��Q,��`��X|rk򆬚#
#�*2z����ݤ�8�wX� l���׍�bj�GD <k?&�'�	u�P��7��d�.H�D�Ti�*ir>�<x}I���ZiI��;L�{
�pѠ��x����j�e�&D�@݈�Є����n�Z�Jnn|��S�1a���4�F���"����fJI8��,��g���Sm����u�I�i�����b��k�Rv�H�)G�(�Dѷ�(�Hڮ�W6��#�-i�0f2�08�b��j���aL��G�j^�(֬4NS�Y�n��N��m��KqKm�ܓ�����V�fJ����",)]h�@���`��sS��,������O��3�an��2���>j�,�7 ە,?+�l��Mx��h���TH�ӣU��.���!�.�A�v;���hW��G��lB�P<7#�׏(H5F�Ɖ�^�����"���W_H��5�(����j�6�>���Ԋ��ʭϷ����z�� IPWU]��e#�ֹ���>��╊2�(}^��=o@#���R��A$d �`X�y�ɕ�x�C���u�zY�~��7���FZ�,�t���/^�V���ܥ/�����(��8�"��.n��j�kH���v�9�W�Ţ�MD�tt�Fi�&���F�?)�S��"��:��cv�]#����%��m��>,�S˶mR�`��	eS'@�4�us��ɩ�:�ɉ*#?xD��D%>?5wy��w�gP�0��a/`_��^H���ui��y�Kd��r�;YHӓ� hR���E]��~��B~�c����oֿ㐼i��2qm+�l��Ş	��*l�a�+e��.�E�r��\E/̐rF�(B2�����3���ߒi��[����>��GX��~F�)��䆰���#�4X��\���s>y�>�E-�u:�~ly�&�����n}���7ߚ`�w�}g�
*���zy`�֟1"�l�_|��Arc�[b+��'q��7��ESt���W.i�E��>�4C�ԍ��u2<��~��#Efs.��$C���YB�����ɉ��V(5	E*��Bup��i�������D�9��h)�FW�`�+��\C��Z�c���*c���R7(�%/�/R?S!���,&� �_;ۧ�ŦN$�{�8-Re���&���eIU l<��v�i�p��t��$ں�<y=��?C�4�a�����ԍًG'��й3��x(�z���(�SSW ︁��U�蠒3[<B3�p>[�I���ûw��T*8w�8�}���@C�s7t�����Լnj��=�W=m&Q*�����:��V	��H==�*_�rtu90Eh�8k}�vX��iܤe �8��6�F��^��������jE�}x��5&���*,t&������z�HQ��6QΖGF�/���juX_����ܐ��C'Ux��*�s��ѐR����(�J��j~����F	�!C��(|^�Ф4'm��N���.�5���)wj��g:��A����iDo�w
$����ِ�xc���{��Rہ]O�Ȳ����[���(W#sXP%.[���u-"���7����"�\2+e�*f �����9FD�3g��NMΊ)9��6�x��\�2</
�R6N�b���=�Ԑ���ċ�tV��I�rfxD5���V���j��o�:��Q���� I��_.�H)C���J�h�&��*���	�Tl�JQ�O��Ε�����Nޮ��3.E��z-R+/M%��t��ڸ��<�u����n���.-`�;� KX�$��6ý~��.�5�H#��H��֍��&��ޱ[��,�a�R׵�P�g�Y5/κ�i�)fŽs��U[1�|b�j�J�� q�6hC���60*�-T]]�wk:�Ť�9��k2D��J�p��X�̬�k(�]S�#>O�ugN�|�<]�<��K��d��·�PL��0�����mp�`!�U��I�	,E��eq�2>s^�=��H�'ߧF��u��5�;����5�Kma[�X������z��̩~�O[���4|���5E�Y���h=�ͷ����K�t�
�����9��c�*�9~�^�]�j�T���F
�oJB��.{�J'?`�c��E7���5.�k���k��uL�Zw�~��Ee��9�FVv~��ܥ�(�Yr�th�y�C���:�{}�2����kae���W�`�م�ŏCtß�}m�;�Fѭ+���*����X#�w1����n��yCJ�O�A�kt��(�0٦�['@'�E����6����M���2�Qt�(4�scQ�q=���#z[���G�fOC*��������B�,]�r&Z�t��8�I�h]���T=� ��Gfsj�AU���`FfG71_��(	n�0Mda��2o|v6�� C����>9�����7��5aM��u/�Lf>V��9��iۀpp�m�4�v��D0~�j�3k��it���Iy�U�	����U@�&���>3�ɚo����_\6���?5"ޤPXŐroz����w���]I��m��}Sy����/Ν���b��\a��t���v���;W�ñv,�;�C:9�>� $�4l�,I�K��ܨe!��qyXS��t�n��ϑ�*���q�$�9a��!�����F�+�	��v �I3���͠��w��w��?���������h��At&fD���6�f�#"0C�ۯģ�RJNc3�w`���Å!��?��	OXQ�h���^B��`R���vTP����g�	0p=ۂMD���2������Ed��<���ÐJ|EІ����߫7O("�g8XW�v�0��L�¯S�T|UF�]��beh4	0{QA*����o�P�Q���,�����tV���\�E*��O������
�짳���8�%G?�\�>`]-
Kd-���0C:Q��9��^��mH�N�YٙhH</�g��P<S��V���Z6���wCU9�g��	��:і""������e��l���tM5}�>�sC��i$(a�����x�K�V�cDL��ؠ��T�T�¹���#�>�����x*=�t'���IC������vw&�l�-��:��\�NG�GS�_S�k����u)E@=������&�L����f��Tv��}���%�T[A��bbQ<ĵ�����&� ~G�����ɝgm=:�KE{�C�.+�=�Kr��GQM��8��mOO��8�߯��5*�����{	n++���������z.\���Ɯ��T�.c���MZU�3��8G�5X1���ZMoo���I�G*�a�OKy?�F����k�8�U��z�qΚkh�j��w�%��)�`��JQ�c��ДAm)L5�Є
�Hgj�sxP��H�ƿk�2*-�kDj
(W���IŦ��|�C8���ۼ�J���:���؆/`�v,��Z�r�Ar���w5dK" ��D<j��z�"n<i=�F�W���8�]xU��H�T����+-sN�䠹�oa����hm�
ޅx�4&�{�OPT�_�v�7���9Q����SdL��&�֩�K�|�9�:T��r��Q�\%Hѓ�kFUK�K49����%�&��v�a�^I9_�-Q�O��[X��f��˚�L#�F�m�sV�y�m%�V:�4t#x���'&~^1��Q-H�97���r ���l�{�])J{F�<��۷A3�uύԕ�H�A8�gkrr!y����\޼}kFgS�7J�P'�y�c��ɀ�T��0�x����Љ+�)f}T�~Op^_�������ޠډ�u`v@��߯����˥s����s�r6֧ع���܈F�:&]>a����!��y��F��>u�I]ʍ��ϼr�ɟ��H#����5EH<�">�.Լ�`���.�f�D�z{ĉ�G&�� B��!��6܇�gG��I�P�����[��4OQt�������QJs�n�X�zG׍��߫�՚���U�������J8d��v)Mᐁ��k�a-V���>(=u5����d�c9�)ءt6���F����`-H�i(N;�2C�}����יS_��jOԺ	�����Ë�R{�ʬT��lƴ������'�����l�����=�SoE�38E�6%��2�$���`*d�����C�M��+�K�jB�u���i�lL]X-�=���Q�u0�oo?2���#MJSt��e��n�T�:��M��&E��i*D������Mx�R$̞�����>6�u(�����L�unң+�o�܄�HY蘣�&#R�p6K�Fb�H��yp�Sr_�ۍc��.�Rb��E�`�pY�H�a\�A���7B"��Hka
���0k��}���-�W��W��Qh<�v�"�:�ͬ(T����:��`I�n��m�x&"YTt�����������훷A��\]A����﬏�9�F��"�I�K�\Έ�*��ˇ��_ߛ�Tt��a����������.�\��;��=e��%���d9�ַ�{fN������eLy 	e4%G_�}��>�;ƸǠ�;�r=$����Bm��~�9Q �^{��믿�b><Q�����mo�>���z�J�sAD���u�W�g+�s���8M��z�xI	��#l��o�L��j)q6�x��jr?�uKo"�E$�k{�fE���zw�{S�P�d+�2���gt�қ�k��^}?��Lj�i&.����hty�_5V�,�����7m��%�ϩyi�n��;&Q��%������j�E���'��k�`�\E�C�>�JO�=�H�q�@����v1ي;'�	$�u{�C�բ�yd�qOoh�M��S/��hT�K����U�p=$3�`>���1�N�?ygx���&r���.�I�M�n]#��u�P�3��iZ�N-KC�(�"'<��<p���,�Y�����~�������60���5q@Ιm�HǓ7�
{ݠÒ�B�~�c�Rt�<��V����.����(=����ڥ�����{��h�y�u���Vө�>b$f[6�I������Xk�3��0x+wN5���v�5?*X	�l�z4�SM;��j���a���B����(~9~��'�4�����?%鏀�(Z	#���=Baz�0�nlJ�8���n�,%�tK� ��a|��h��ru�Z��aQ�Q��� ��� {)��76�ҵ-ʘSM(NC4v��dj��}��i==i�H�\FV����զr\Dvn��C����E@v>��B�D`@Es�5 j��q\��HӤ8%j�����/0�����՚�,���ѽ�R�_u�\�#F͡g,�"����^t��O���q�ށ�u��������+�"g=F0d8�QzM�j���S;m!�9�YB�W�o?TX�p\���o�����z�zF�2��A�����N�VU���[�9��T2����Sݟz��o�����|L����}�j��O� dJY@M���f`z����Y�Lg�p�D1.�wTJ����G��H��,�E%�
Ye)�y���K�W�����o5�o����ٟ������Q=#�s��rY�����<r�u���$���!�GO!��Մ���`%� C%`�D��u��E*��M��SʞɳQ�f�/�4��w��S4qPt�ON2�~���ߣ �۽��0}xC���,2�ϑ�xo��� ��E��&;[��Dn��tY�9�ay�*�&�02|�,�US<a���6Jt�Þ�j�틗�i�:Dw��`�\^�o7v��wQPI�.>�*��>�k�9��!���K���E��u�{YG�E{Ƣ_��lz���8F��C8]v9�X:�}L3�N�GFቧ-Q]�<s��2���*~j��E�h���)�&�j����Q���:���VD*��Kij�*���~?�:���ו��$5h�p[F�h-�ߡ�V���c9�5J7CC"���3�b��R7;��������N�ąz��g�i�!����Ϫ�Yy����|�@ߨf�^�&͋/I�(���� z�zIW.�W�#��&�9Q�����G���q�'7����D�D�Y��Z����n��Ɯj�T�^��q�[��hX�^S��}��b��MQ�H]�wRJ�H��z{[$����h.P�G%��ɚ��ڄ�ňj�NC��06"��l����ײO��"�R�4@A[�����i��5�X�_�*�ީUT�G����o�%ǖ�g1����{�L�<<O���,����<JE����)i55M)�,x��l��\��:��q��4��,�s�ZXfaH}�� k��v�x�XO�&�g�s�68ǳm��r��NٴQ<2S���DtM]w�:]��q��X�3�63{�u�?e����F��垭���\�-��B��M/�d9�Y�s�t)��]SqƖe+��')C5a�M4Z�'�Ƃ������M��%~���h��� ��%�9���C$���BUY4�)1��铞��[�x��MDjyӺ�Gc2��:���=G	K�
���^��W�-_7@㇞���n��uD�@��OܹRmNimf�~����!(F0�8t8p"�S=��n@���m��}V��6��\�"#M�4cǽ��w��K_$���!���,1G�.�Rd�Q}��'�N��x։R�}�����Q�Rؙ��|�)FO(��i�@߬#%u��3c�"k<�N_�uu�4�ù�����Z�d��8�f֬#/R�r(�^K,��P�gp��� wL��J�b��}�ڂ�i?�1���9�M6h<6��&�53���v�;�7SZdnuV8�T� �EMdQ�yƵ�k&�±�Q�����H:���٭���>�-w������)L������?y�%�4��c(���s��9"U�[{7HGp��%�g��Q8�a'�ǖнύ�h�cڃ�Gm}g|��A+8����Rlo(�?�R�nLU�Tj"7�lz�t�ٍ��!z�h�<;��bw>K�|P��6 ��E��Ř�ym	� ���nh�N׀dw�%D��^���wvXLKz�t
����Xt4�(�ag���g���]��Ro\����XO8Q��9G\��EN��&R=��a�x
N���SVz���..N�G]��7:g������5� �Q����\�W�V>���'iڀ����Y\��j��޳���l���oo�ѡ���S����-��4%pu�ۄכ�Fr�y��~4�ޭ �ܺ��<��B���ޓ4�t�e�4�ʻ
eH�Qк��H�U���[����jC��B������T�4܈�^�ʘ*������"����M�K��ً*0(�b��@�!"�k,�@q}&W��Aw��mnYq��u5�� ��Â��8���<}C8
��VEJ�F��ܘR]h������G?���&��'p{�kC�8՛�m���$��p0VF�3�!�5�@��`�aP�T��ϱ���)�����$�"@�` 8����iNִ)�7���B�HB�k=����-^,�s]�v�g��'���~{���d�ɌB�	�	Eӑ�6�{���Ģ���=�j�8o�f�F�Z� �K��Z"��]�W�QG��X�f8�1ǌ0ҿq��G!�E�J�ܫ;6�8i 2����V����u�ǜj{�QM�1Ѡ�i�:�9Px�Lk�ۇA�����dkT3Ar�_�X(�$%���9�0���~�H������_�2J�
f�����L�M�wM6�|�F�xf:�l�_�@U�k��	�t�n��������H�$�1W���2�R,�rI�_�eĚ�����-�6�����WKl���Sy0��i��o�ug��F��^�i��bG�<`-{Ӂ�qн�l��K�Z�VP� ��OA���o0F;E�s�'g��5 L�BQ�H���G)��"-a��'(���-��{���9��g�*�o���68L�Y��&�1q�o�yw# �,�㜪p>/C��-:���u����$ڽ���_8Ċ������p9�.�$�����d�
b�6�WG�ZO�#(	G�SG#���!����;p�e����ं��5�����#)y�s����L��7ERM �{i,���_�^�j���C{.�U����Ft~�����3Q�v	��ȤaI�ß��kŷZ�7�vG�{Q)?g2�W��ƶ���_�v����m�\��`��P�G�w�q�h��.�[X�� �%��HE�xE��e���b���M���B���x�����ݾ��
h�OlU�z�x��Q� G
AD�SF#��q�}��;;h�?,ת2�Mf��B�/�
/C�7�r��~K����]�'Fp5��I��<��r!����)�]	��ީ��SY9��
%������&x���wC�ʽz�Ma�#�������ڇ�>���ѡ
sϮ��l���Q\��V�vJv�L#��$�ڐ�@� 6���	��0����~��fwއ��g!lp�q�ǴS����n����lE�Keh�Cʂ���F�h�L�� �1�V���J��֣Ud]?��c�l+����k2ٯ6 �a~�������#��%���O��MR�y���O]ǈB/��F'�"���%��t~��.
�9|�Q!������f¤�����$�3�t.�ն� �5��JX��{w����UC��-����))>��cH[z_�Η͍6��J�KvO��%���{��X���hz`��z�;/�ᰙƦ3%x-��y(U�����L�l�w7'����ZL�ٮ#��:"a�/���Kͥ4�ML�$����d�/įս��O}p�˾hb)�s��ud���.��a�u�S��.�&�#�·��{��F˴<�^zZ�S����]"�bRYک���%�%������ A��׫N�� 7����ԝ����L�p��.��Qg@4%8g\+֛i�.����K�1���5@��3�I���N�u��}�3�~F0<��X?��i��I�1z,�2�4�G��j���#�GƮN�e�j�>��T�tY>��T�풜8�K��K�^�����|z�ҵ0~���W������H%j�8[	���n+UQf�8I�5%�s(A�֖_�}�%�L2哃��}���������߲���^j�M)�:Q(��I:l���i�TJF����w���Q���m2g#�i�Z7f��8F>�<a����ůA�ۜ�o�_��D���c�f��)Uw���(@�V��Oc��n���:EI���������3�?�#�>�=��Z<�t��D��?5��|~0��$��QG�7�ԴA?£��Y��>O�<ԑT�i�g��r�����QpSS��Q[H���d�y��T���K"PЇpe�"��:U<aer5u�뻈�Ek��:y��H$�<g\�g�������o��jޭ�LJ�4M# ��R��h3Ϟ����Q��u<�A�Q<�T�tC���P��0��,g���@��CFimt��B��vpp�]�z����`�l}e�ǋ�r��(��)�cxwp�TT���%�&��z����H���������b��� ���ާ'�8��UU��Q�]p�$d<�)�����o?��E�~إ�ZD��c(�_.�s���T��"�NDp�H��j�%q������j�7qΝ���]lQ�*J����>�='��`KPx�}���	?�����c-�n��	9�������.+<�v�4r9-����������?
J���Yޝ���Ϯ����G����`��u�!�c��⣵��3��vf����l���Ƥ	�V�Z���4E�\���պϛ����$=9)��	��\��Z�uO`��;����f���І��'���O<j#��'�I�s�	��Z��g]�Q����)�I%n\�L͑�M���F3�iDJT����B�mkH�Aj�л5��uU%�x/�s�66W�6OD�0��!�,��)�lE<YzϹP�0�����5�8c��D�y�i�J��ڄz�
���0Gf���[� kPo�+1"�.7�B�O�&#�E-��j�� �ZFΪ0�)���e3l�H��$�b-5,u*���%�Ȱ/&6$7�� �!�7R��=ͳ��6USy��9�1{|/���M��y?�9
���q^°��&(kj�|=eH� r��ۃ�Ꮟ��o��7v�9{�~}]Mvǿ^Vߒ�l�7��m+�~��_S�z�����<;C*To�u23��a���n�(Q������ʜ�N�s�s�F՛�n���Ҁ���3�Ty�>u��R-R�	��a�^���q��Z�c[)����nw��9�8����Kߴ0�x� Ȱ71�%�,<����܄7Q��a5���N)�N�\�hK�Ϳu�O����z��3o�|0�O��������!r�3�F��pF�+�H�]$��������Ǐtalp��Y>d�J#	�-�k�}���C�/#��;�Qp�%��9Ei�FS���v�k����T�h8��8��4���(���!�9}R�Ӊ�-�K�7�(0��O%�gb��R]��~��4�&��ۯ����T��ȏ�?QyB�sۦaf��o�n��J���9ʊ��6�3����&���6��0�Qh3�~�z���K�L��+���>% �~y˶����1"�q�ǽ���c�����y1�͛K��}^�^"@��"�t�qj/���J�P�MA��ee��O�w�����g��Ŀ�*�@U�gWO5��O���;ǒm�%#�q��w)>���s}T��{]E�Qׇ0�%���9�	�*3}uq��fT�-�Ґ�MV���ʏ�.��L��C���<�ɣ��*�"�7i�"9���p�
9s�g�7�8��WE�*�ܔJ��ٙ*�TϚ���q<K���g2��A�ѝ�爵�`+��Z�P%Ew���	C��\w��#&�xj(Ǡb�al'���.�zȂ��<`Xe��T���>tK�,��~�Iےv�M�-ɳ���Mq}LU���0�\�-�g'N]g(�:u��.�`�0� T����_����N��J\=P� ^�z�"��d3����#�/Q����OL[82� ;���Y�F�	a��T���	��;if&����-���3�Xp�����4�`���,�2<k.S������)�*�b�{FTPmxEK�U{u)L^�Z��%��=|D��W�qP|�'^6�z͆��e
�*���d���PK7)�T�kէ4���H�0���o.�ei��UZ�Y7!��|��3{���P�d�DR�_U�W�D�-�M����[lVK����>'"�2Z�s��B ��J�i�Zoٓ�}�6�qW�-�N��H^��Ud�T�9�;{��5M��b��9>�0`
ҩjI}��E�A��z6�!���]t[�
�C#qev[�I;��_�εcw�p��=U�l�\԰A|�$��O����:ͮ�����瀭x?���3�F�p?��K���u(�۬!����R>ru�^$��j�����8@v��j�d�TZ���h,���Wg|�̯���{~B���	'%,��麇��Y���R-�[F��������޴��h�?2>��
:��:��A��hF&��s{���A3�1��ʐZ��EҼpy���Fc��t�v�`�#e��C¤rJ�VQ]GJO:��T%�oɶ��{}T��J�(u��'9�M�J>��ݷ�Y:����?��MC�<FE����պ^J�<�s���q5��y��KF���:h@r�:RCNI=���j%��ؼ%��,�4��11�n�,H)�Q"��g�����H�U���i܄$	3
�Ѽl����É�ˁg��wx�h���S��&� !L5]�i\�ͱm�Z�_jE͙c�{g�,�Y��:���ј�����KM���¡T���M��ދ�"��:7���:�k�F�uWזĎ�TZ/����k�kшX=O����󽋀{��=�M�,��s��z���OG!���ɮyy�dޓw}�=�+j�գv:�t�/��ܝ%T��z0�?����z'�@)#�%��C�G0����2��R���P4�B��.��9�����9f5{J0N�M�Q&�^u+���;K�I�
P��d�H%j����m��I���Eё�$�n��#/�8���ީ ��N���I���0Ҹ���_��^~n��,��a4�����3z��]"r�F�9�˿����8x�{�6�w<A�!�w������>X{�ٮ��q�5D":J��l��� ��WF��' tmU�-/�aQ�ܸMj�hZ5T��b��  ��IDAT4��mk�ŮJ���k�7BP����A�Ǝ;ͪnFׂ;����6-����0a_-��j%���.iM(����*8�Q!��>�8�b%�L��"u���H}�-���'��q�q��]W��#�T0��y��ѯ�랍aO�;>�%�������k߅��1$
jd�Ց$�2��鰧�^�s�T��0TA]K�8�Q\b �T�(|�� ���Wm�%�����.��ܲ��i,%
0��b�{�s�;�P2pl��k��f���|�dۙp�z�M �.�a���H�N� �韪�}��<��~~X~z�8^�y��(E?vm�@������?�`���~��A��ң��7}�b�"m�n?O�-!��:�X~������ǋ|0\�O��[s�'���ӈW���[�p\u��Iő!R�\Rw2�pp������6�%�7��}ui�R���
rⵊƣ�B������n#��,8�bŏ��3���d�w0��W��&�2��,�iGW��T�C�]�߸�J}QɗcA��#�4hN�62�Z�}����|�s(�*�)5X�s��I���}����E��@j�RĆ�}��.��*<��&>����}H�'���1a���`oj*��*d�����|z���2�Ri=5I!m�c�B��A�x��!�-�Z�B�ߣ��|6�9:�8���0OG,�m��cr"qs`LΧ��A4.:��x����-߸	6��)�r�n��0�go���33��ݠ 7�s#�|��Jd /;�:�0� D-�����?	z���I�U&��H����!y�����p/�R2�)Q^ߛ�'���f;@`�%�-�5)sq��F]����hb�-�^�R��fs���*�/^ܹV����qP��♍�z�%m�Ѥiq:ǵy�k�iF��Jw�d�3��?�S��L�zq���w�H;I�[A`쯓G�Z����\�qC���'�~Xm�R��W�t�X>A�hu.�7�7b�hm�4jd�����~ľ �6T�q�^0��c5�2��T8R����x�1�*�\�ݰ=�!��:�T��EZ�~9�"E���S8[��a_����-N'=ͦl`_�64���E��R�;7������!�V�RD��o3p`�900��8�V��q.y︙[�7o�2s�A{�6�6�`ja�7zt�,�`�ĈdP�9�8��B
��`'�m ��I������Ui:���s��3U�<]�ݙ��~��T�JQ�ka�����T�b��"�3��}�2��Q����޺!�3#)�)��gg+Up��q��FV$y���?Dz�ͅ�U���sBYp;�=���P��w�W"Vqi�4V�j�K�fR:]rb1�!h욵��Qvkɭ+Q	��B3�[;��B�ukFO�S\E�u�pJe0�˸�Oe���Z��l=+B�tZM�Z�ި!J>v�}�d{��+*Z7�"eFԴFO4Tl]M�c�o7G���c�gm���~��:G���E�wqI%U��^�~�L���KL@�5G�)*T�S�~�o�N�kj1��umH���
ֺ*:b�q>���6��)"њ�V� ��* �'���1�G��D���S-�*\<�G��uYс�m�����{��=�1Uꖔ����y
�N�<�ͫ��L�	�:� �`�'�x��G���8T뾼~�:7��f.)h���'�!�X��O:E�`*���=��S���n]��j���<�ڳ2�,8!a3,�H)}�T�x����&�>���Rt��0�	{Rt���p�g:��(d`�
���4m`�l�uE-�#|}�Ā訚(:c�*|^�_����n����=c\�=�#���7{I���xK�GNn=X��{��z9�yt^wA1���E�iT�K�����NjVEZKY��S$T���CP����߸��XO����v��Q�tcϧ(N����P5���{5�(�Wǔ�6;����N�Κx���K5���J�?�1��cp[GQ$ڼ��j�:�LҽJ�_]��F�"�ʺZ��o�)���h�Y-���[����2� եs�]�a�nXM�O���=p���׸����w��h��!�ya��Gћ�0�φC&buM�a[<��'���)'�yL`0�H��X"@P�4<b���Z�\L�e�}�ͳ"#�v��S)g�$a�d-������օ�лX����F�C�>DǗw$Ie���ޮ���?�bUo#W߈v���3��f��/�Msblո
�'}�Aբ��m��M�t�6�-.������e'�E9�>�����y�G��֜(�T���)̢�"A�&���1�[r@``��W��!C
c�lAJaj�Etٵ��L��`_�-*���`H��jjt��0��U7Q��7;��/6��Sb�yA!i��x�j��}�2�]=�WVC�r܇�\�}�{������[�]��^����*e�I�4�Uw\��N�����L��ij_{�0�S՟-2��@��"�lϼi{¥ψ�>K=��ԜeM�EUl, �L��M���J!�X'ۨn���'�����o7�rRuو�YS��R����7�PЁQB��f��NO���&A��?���z����=R<���)6��\5�Ŧ\N�X�4{i̹8�G%}P��4uE$``���?�aF��_~*��߽y�3��'�w�u�"�Sj���k�L�:�����/_���ֺ�@�
�R_S��៓����7��4�D��,�A�U�,��%d�}ں��E)N�3�q76�*j�LN���c���"�Dr��NG�f���C��{i�T�p4�PE��[�}tlT�*:1��
ĘQr55�[�q�3�u�����O?�lq�hf�Y��$�W7'��W���&�p��i�v�w��a�D�/&:R9!�TZs�X45U�'�^�vA����3���8$����+�����c��+&R���r�:�O#�����4�ؐ��z���o��䇗��&��!�Ȃ���}T�=�fZ�~�QR_��m��'�.9o��<e�g�'���,�&�������ތ�Gg�x���H��ro�?��QY(^��4
/��Gd|�'&�x����ޗ\��Y,%�u�%:5���N���Uiۮ��Z��o�S���-u6�ߤ���S���r\�(.�~�P�`a�4F4�-�6�Y!mn�]�G��ꞌC�~�]�%�,H��yэ�QՖ�,k�O�9]�К�Ve�0�����}-~_���+��Ql�jR�5���s�!��ZWMw�τ����{f۶��ĳ^{�&C��*AթR�X�$�+T�([k�`*��7Z3F���?,>��+�3�5^L�Ԟ�;�V�:���M�^�&�7o��a?���Q73��K�Ö�����C��2D@p^D�m�|��Tڿ�G���-�E}�i�%���:�➀�@/��F3��Ci�����<e�E�-5 _Mx��zm
	��+��S'1�=Ǌ
Cw��.�4q��mQ�R<]Lu���J��)oj3mn��!2/�ƩH�xC�GڈF`�j}T��)�n,z�3m5��
���v<�?�(ڍ"��;Í���[��	�k�w���#*�Rv)'>�H���4�(��oQh{�^�)4C�L�5���POؔ@Fk�#�<,�'.ȑ's6��"{��cО�,9�f��G�YzK�ib������W�}Qp�
Ք��a�#�P����T�u���A�V���g��S�k�6c5�P��['��Q("��4�k�}�u�>��V���>�s(���e����x���:�5�3�`�nn���>��0�^Nݠ��˚U�Q����ӏ?�
�"[U��EN�����#ҚF�����
����	'��'͵�G��Uj��# ��պ
�����&�P����kX6����)��asӐJ˓�MS�0o|.6���\���@�x����t״���P�,���v�cQ���T7	6DfA�u��EQ�KL#��ŭ/_�LT\�|&�Zq`M�V�T�T���aM�ؚ@�z=Q�8q�z����o����򹴡�Ak�l�%��F!i;�X����c�oMcN���74��
#��]I�l�	]�5iђ���q5��My����
���w�}�^ue+�	8���ׯm/=X�gp�y��=�;���gJJ�Z��~�����(d�E���������\��3.N�K�vY��������ER��U"m����s��4�Sg�D���u���� �ޑØ�v8��O���u���΋�3[��E�M8H܇ś��u�<ؗ�;�޺�-v~qn���{]��"���Ծi�Ѵ�u4�{y|���7�sCZa>5�<xW�B��8{I��i�3�ɰ��f����PK gO�D]+2y����I8QV�Ii����}vW<8�/yi�6~O���=+�鯻gi_v����b(4b��0�-
��_�:RHI��1�m�~���������x�Y������)K"�)�I�P�F���$��߿{�j�N�Z���o�[��X����Pn��4Z��U�-��:�X2}Ed��)/˛�~-�Z�D�0F4���AiFw�0�LGiԳ�w���鶺|`D������3kX_ԕqJ\�"���dxd#���%[�������g9D�3��|��Df�U��_?Z4*�[׾ꖺ���i��${W��E6N�/�ۇ���uu��(W�NJ��(��mHVJ���1�nHA?���n��Җ,���X��	�8C�|h41:��|m��U�W�%ɹG�H�S̓����4-rp��2Z��cF�����Z���z�i:�2̈K�9D�>+�FL��̱NS��k.3��B
I|\�����H��񟷈�鍷F4j�����_J TSQ)�]�&T �� o�兄�T]�X��AF���Jŋ�w��b�`a#3���H�X �)�o�FIr�)
?���#�յ�Z_��r���(T��� �C6L}ˍ�J<M�Z��R�Q���
_6��B�a�G�+.���n5l��am��i��������Ѡu�;���y`�b�t!h��� ��a����f�����:�n2��6�O�%@W׮4^a)����}�t�ڟڣf���I\:�e�UsV.H��E��Z��������\�9i@J��1rX�GZ��ҬN+��ZJ�;����Y/e����~�)�	���Wb���cI:"#4:]�K0	po�yΩ@��@�4O>�j}]�7��BD�Oe7�l� �O�Y`dQ3]/�{�]��7�8F��w���	��7�U��W8+���X��>�ɵ)��8wW6K���3�[�+���1ϭ��#�X��'T��M*#��e󅅃�@4&A�q��6��ӣ����<&1��(��c-����r`/�j*� k�-Gm����:ڇ�)�'j����/3�5���h��>�m�ׯEc3$a�vΫᓌ�h�q`Y����kQqS6�)c �~����E8�!v.���R$�lֿQ���ه��/�ص�h�D�j������iR�6J�̚꾸�su�OJ�!����y��A��gZ��nQ�X�{\�SB�#>�����q�n�c��g7vX��9��߸����+!���E��{Ҁ�O��I������������M�H��jL�������SJ���F(:����17p\ѩ#6@`���>�n	Q���\{~�Y�ѵv�cipM`Ɯ�%�[�BX�����
��?���0�k�X�c��&~�d8�9� �9���!H�ɢ|��H_���I49�thA=C4,gn�l��A����{rt���=ˌ�J�?��I�O�6M��+P�y��+p�Fx�&�a���t�ibEX�j=kZ�M�J�R��Q�ޢx^��>�3�b���95{���B4�ǈ&`H5�M�;纏q���~�hk�2��� �I׉�@T�߿_�������5H�%T�����B|�p�tɣ�����`J6#
#��%/KИQ<��K,��a=>��#�Y���o�ѨMsN�-�B���n3�߅C:�$��Do=�ų�&��&���'�Rk�Q	G�2;Dg�Q�|�:�h���� y��p5�	g?���oY��L-��	W���áVXb{7��I���=�zX�g�֢S�;�棋oc=�5H���0^T?�b��X
W�����'�ґ;y��č�����5�(�l���58f�����3���Raλ�j�%	�a���XI�fc��X�x��,>��ihx�}LQ9F�;d�|}�*q�#�gE&�I?ɔ6��~~�\�m$A#�D�i#���Ȉ���ȨV)5��H�T���,�գ,��%��"κx�'v��"n~7�N�nð�FǄQo5U��B���Z쳶����M��(4^A��S7�	s8W��W��o���HE�	_S�u�����`�l�VVl8lr(��5�^�C�jd�ihV��&���л����
�m���	�"��m����8p-U43B���[���,��A��x�	��dWX$��ɱ"���j�l]�@�%�0��)[M���p���~��ƻ����֕���:;�T�J%�.";cq� Vc���}X��V�C5KDB)
Dd���<�u?Κ�K�N�f`���1�Y*NĘ���9������UT9�Q�}UѸ%�'�a�Ԧ�"����
��M�g���.�2�(~`�C�m��v�9+u7�-$�����X�%nov,�>����z|"�)��&Q��Ƀ_c�!G0k��~'I�5-�kI�0��0}|��|��󶍍y�,� `U6�r�wC,gP���h�����y�$2�DT�J�m�Ź����cP*�Z{f+����'��x� r�vFHU���C���C���9q�MZ�=���,�]ʛ�o"W��u�������[Q�Us�{Y3Z���`ׄ��uB� ��y�"�����841ѱ�X��Z��a�H���V8r����i�wY����`�k9��) ��5µJ���{�#��7��������?��\)������LC��j`��f ������%|����pv�:��s�UTC��בbӲMV�XW�Y�)������U�P�3|�;ز�MC������Xp�S �CSJ۰`��G�����`��͡�)�Q���,�Q(<W��+�X�M��(�8�*�(���xh'b������})��nY���!UT!��FԖ�j��7�\�w��pPb������ ���C�ޑA�����´KRs��K�@Tĉ����1U���Ｐג!�Za1�~��y1^�<�C ��ǟ~J�^�8Z��6n�@.��(`���V���߈{aN��>Z�]_��SCy>��}R��GB狫�_9n��!{��הs|K6Y�I��{��*���:�\HCSWvζO���a�MU�J[��#�K��	�I����g�}�����&۸��ԩ�fܟl�Y�����G��$�i �EPU���m�󶰏`�O�S�]���w��)������eb��d3�j�;PR�ޕ_��k�5QT59?	��|\]���J�C���p��cm7��W$��lJko�-R����8O|�lJN���
�Y��?�������b�ܖ�h2<vޝ�I'��yӶ��a���j��p�W:�Y�E�1sY�*b�XƠ�yI����+��c*��<"%olr�x���r1��K\Dm���$���Z
�����|r�nQy��!:��E��X�Kfٸ��<�ج�+��:�V��'a�) [��7_S���F7	I+UV5?�;!����Zı��W�Q�!����ȞK��]��_]3@"(l��i��	+"�X���,l׳� "R�3#.TWmmY�ױ�OXMh�5j~o��x�!���>��M�&�>l��T�����iמ1I��|�6k��t�z�m���lI�B�a|PZ>^�3ۻ�>c��|�"%�a����#�*0��b6 PI
Դl?�f�mVp0z{�`�~���2�)�8�k������iB�V#��c~m����*����e��]��qT���4���<4;gU\k��f%�%����0������ �3k�X������Hq���#0�g�FVc�Z#�3�$�*�#�3��Wr[ M�S���(�qJ�8������{g�>��MSo�%�z�o7�<o�I��︑-�G���-F�	�MmeHe�j�U[y�l!L�G��v0ݰ�.A*����@��mC�K���w����`��t�G�+j�61,�AK-wqȰ�~�����'\�x���(���l���'�*u�S���I�\K���I�Wꖠ��sr�wȤ§G��p:�]ﺱ�o)]�ma�Ǌ�G�8���#�Cw����{K���8�5���� I?����S�5E�Q`jRR��;��N�H���g��W�DHm�6�����M�����M�^�ɲ����z�2�d4K��r�(:N���x�7G(��v��*�
����Z#�_�{��*%|�sV�u�9�� ��!�����9i�������Qݡ�"�Q�b�6�{�6d�V�B1ZRC��ep�=�#v��z�P�z.�t��h|�����u �4.�h�(_|��s�W��?zH��l�����KV�'P��bS���m�ҷY�hsC"�%��sc�ti����y�YC�ćƈ�ŇT�����ͺDa����GU�gF����bL��1*����H��j��!��C�����~��M��1R
)�@39�9�,*׾-*��S��%�}:�uȯ.5�9����m�d�ם���`�|V0�ѣ�ǆY<rE�Ml�p~�4� �꣪��!
�x�!	�����7? �ً�2�Ͷ3��[������7�����
S�uFf�S�7V|B�\����m��ʐ`��,U `dwWh�=K@G[0�hu��^f� 8���6=R;3Dhx��'c@�	��]2Ua��� E�N�� ����@�)�<*��x=
G��ĩ�(��@Ӕ0l�o_��^ߔ�8��3��B,�	ң��t�Ā�_��.�TI]��U��AR0���isȈ��6��c�գ���?�|n���󈴭#�6�"d0բe�[�h�����Ы�&�/J�p��f���hc�����1��4��}i�0�q������A�(̬�7������TĪg<aS�ۈ^O���z�*6���;�Do\����6��=;1l&���,%�!��W����ɢv/*Q����7Y��\>n}��!��DFa��^�z��1B�b ��} �q5���6g�9w]\�郭���0�Z�����Rl���?'wxS�]��\������5\�9�u]oonܐR	�k���v@�_x!d�(��}�'�ˎ<�xu��L�d��
u�X'c?�i�0S��VE?1�RPPCF�݉�FOb�������~�߇s�����s�����{rA�!�)E޽gy�\IÊϧ�2���ZDH��4����vސ����4���c�qc��u�ڦ:8�8��~]q�uV�nP���aːj
)���#v�=��o�F�3�p�# ��.Y�% эIUOJeL�f���ː�EL��R�>jn?��4���X�?���ǻ�p7�.F@�P��&0�F��B�*T�ߚ���`���W����xs����Ӎ�,)��y"'`
7���-XBl�BɽGcχ�e�$emX<,]s8i��߿�Ap27���ԓK��*��˘
��H�['�g*e�D��T�6����]� �iJy�B�;�*tKF�˜\�R��w\��6:����$�v�ǭ4.�׽�Q��7�&��DKC$�ȟ}�W�1����	1꒩�g��ӝW=�fwh\
ۆ[7�ZΡ��k��V<Gq�ٚ��G��	���k3���D��Ϥ���y$�"%��/Bip;7�9v��;��H���㝮�wx��t�=6�����w(���=ԋ��%��
��9�٦uc��Z�� �Q-��N����>_�������N�3�EB.�%����M�"����߿cM?��f:X�P��"�J�5Q�H��&��jOTTx{C��6�bB��� �^8��=hc^�i=�O	��sԶ�WmD� �]�q��L}4uR�R�'Uc�)ܮ�z�y�����0(����`1�s}/D#�$�ñ��,����Ԫ�r����Abˈ�S�Č��X>F���9��A�� �[a�U�OF�gK���H�9�������Z%�R�f[�M�5q��Z��O�h�m��ڽ��0�6��Z�zا$�W���T�
;��u���
XE��%��auS���c��燑B6(�a��h�a `#��!껢���@:��d�N�q�������~oYC �A]q���E��k��/����OA�E슋�:��mlLe4��������&}\���=�>f�s��"o\�YjP�P�U��SbO8�M�h�����G̜ A"AK���iJ����Pz�>�D��M칥=���?��7��c�����9tCQ�=��%�dQD֛�)3��/,%���=<�q�&�%s�"�[�̔o2���N�$�,���t*Z�9��9:����i�y3�q�y��~x8�CG��D���b;�yg���]�M���i5�[]'����~�.t���$���^}����1as=.�1!g��Dڐ��_�`E?+��	q_�=�_F� ��Q~\�z�I����P���FE�٢ \��M���zM�홌��_�Ck��N��K7��/�����$��Έؼ��sv�ᵎׁ��'��y]�ជݸҥ�q\���4>��q)���&葺����*{�v�&w����k{8BY��s�2�bWw��^�W�BBA�2&s�r,No�y�D&�P0dF�O��,\Q��^�'\�u�{
�c��Xq��*�;Up`�F�Y�t���PJ�0_vN����{���b�\Wֳ�MPYա��'[���)��|Ύu��ba[F��s>103K�a�Xt�6���1��$օ;'%�#	�PN�ϣ)�\.'Sg���&�7�s�pBmH�0	�S!�6��Re����
7���/M5�.6+�	�A�
ԖhH�����7��f��>fL�av��t���u��u2�aUǛ�X�\:y�t*3����������~o<QPJ�ۈv�#|D��o�;U�|��'"R�Q�P�hkxb ��羿���~i�����9e)�4�8P��/���Y x�S�3�h�0̈JŨ`�Qֲ�9ED�e""}�^r�0JV�p�9B��S0�|����s&������[ߏ�&�|�@�$��8#
c������+�JfM	�$��r���TR���4n}4M�TT:��0w�(�%�6��pWP�P�������v������;��>�=}tMb�y��;��GJ��^~��֣iސ==�k�	���5FZŢ�ʧ��Վ��_�Bը��8�R)D��ܥ��E.�Ns���"EHIX��2GX�y=�Cu�
���j���UŴ�H�6;�u8��b�i����ʠ+2� ˻+
%D*:��a�/67�uy��D-F1A��J|աg���N���ɡ��9Mq�¹���cgѪ��^ฅ�E�j�
Jͧ��-�V�Xa/q1�RlB.�{��_��X���ͩ@��5jl��ã�
��������$غ�j�Cg��q��)�|��(��!.��#*���8��2���ǲ�Hk�>,����E��b:-�/w�Ւ]��,gjx4"i?�g:h<���p��9��1ޤ9A�?X'���8����|O�6��4"P�c�Hgfs���X�3�P�a�����
��?J�SQ��s������{��|<D}�j�}:�P��r�6�$���Zim1A�� �h�Y����LJ���0�n�}C�	ָ_m�ܓ;�ٙ$J�&k>�:$x2���󣖥��U-���S��Wx�[�z�wXUf!��)	n���"��/v�C�1���4__g24�.�|��1Bp)�Pp�EhyJ��n�b��-�c.����&�uq��v��)�g�A;� ��:M8��}y�F�H�8�䃍�Ib("�ӣ����>'iO�u�a㷾�,Es�D)���t�'OUL��Y�Pr�=�}ai�m���X����oo�FrcR2|�`� ��(b)��;a��w������B��k�磳���R��"���]'^v��X�0.�����\/�x��K?�1\7 ��iH��3f�]@<Ț��Q� P�W֔�)����gqȫ�ۀ��ڥ�YcY ��O�A7�~��,1f&o�I8���pu9F�׾U���0��X��C�:�R7�� �p�ܮ��=�ِ���1t83F~�o����Dۯ�x���ch3�WD�H7�B3��f��:np�n�b7]|��]���jS^��M�g;�=*'�8��oKH�Q�:\K�bэ=���.�QJ���ztC)i���F[is��h(�H�V�w���ȓ�2�SP4k-0����֣��V����W嫯��4Y�6"�GO�mF9�8����3R^lVu=1U��,h�b=F_�>.59_XdE�����0��.3��fX_�x�<��Χ�R����zK�pm��,�W��Ӝ������Nmj%0�z(9���:�n��]'RS�Y_��qE�9$���e����=�ɢ!��hWT�ii� e\��۞�M���6�/�u�T-��=���gá�EU��"ņ��+b#J��ڻ!xFT{VԵibuX�_M{�$J��� ���\o�m}�Ѡ�!����_F����ώs#x�f�?a�a|2,�x���$�c?c?iԈ�>U��پ�!�N�ә�����������_�`���ć#'w�S
����zݵ�hd�)"�:�櫔�(�"k�Yt8!��&)k��j@�T�Dzҽ��xX�[�Q��!�F� ��?d�Do�h�@c�s�U�m��ۊmD�GMo��ɿ��FF�{�ٹ�DJ�0�\}߆h+>�QFaY.�zY�hn���l��S�M8�&'�;W�O��
͖�q1�>��p$�J��UOŜ�MN��
�u5\�w5�����;�X �dMS/r���R�٣V���xtm\ҶMϾ0�5ޣ�-->�m��.�wo���D��3��/� C�
7�戀�3��*�~PL���x4��J�QVi�^����mF6����y��Ce�65?��y۾�rx��� 9nO��3��9�0�T[�^s-3�3�	-U��""��6�ϤHI*��Y�f��Á8��ό�~�]��s���
��<[}�䐁��\��)�;-�����3�)nT�1ҕ��|�p'cJq�'�,�Nq��v�̻fs�dHe��O����͙��	>Q��m"�Ń��!��eʠ�m�)�Ti�-�q����nM^QM(��A_d���4i&������ņ����7��l�����3Vh7�����sZL���)����֙��}�bS��|����uF�z%UJ0��Wz���s��B�NU�,��ܣ�HPBX��֩单Q��j�������-�Ьl�}�����읾�qƇ��Ba�:�/6��zk��6��@e�V&:D�R���y̡.��*ǀBLJm��3��S�px������x�5�+�7��=Wx�R#eT�&�7�wEeë�w��B7n^DoF�[,:"���I���*��Fs|kd�~�u�~g�[���J���,-��֛7�>9-[e)�v�3lTWz'Ƕ1(D{�Eܱ��2��Ǹ�u�B���z�>�ds~�Ս��ѓ�fz�m�C�����_��"�1��z����(*U^��uY�!���t}�j6�p)�M4��^����T���-!�e������^��9�sKx��\]�TMv}n/�^���;'�F�W�$���T�u#��BI��M�]�==�v�
5�VUHPt8.��:e��f\���+C%�#�I�]����w���!I�ΑE���%�O��_|����W��OjҐf�����4�H*X��s]E�#" D¯����/�o^ݼ0j�����X�E䅆�!�񔔩�Qb��xf�������S�y�&��:o�;�S#31UT�
?��`}�����{�Z䆩���LD��c(������}�z��ʴ,���ept��T�Y%�Rx�lK�ሓw׭�Nc͡W������d�W�x��X�� Ԣ����w ���*���Y+T�j�;��������S#[4FE�D�q-һ2�S<a�t>Ť� ���y�q���ZM�h$����2Z5cA������5;LR���@���(�j�v�z]��:�Q�d���"�MD�ܘV�PvI�u:�N=�T������S�a/^U��]��PO�Dd��mR�X"В��i2��yY2��>p����\Вv52E\7��)6��7�~kt���֮ׅJ�/��HZ�$�w�."Q��de��C���P�WO�|�-~�����=�I�#��L$P�ը��R=�����ܷ�w\1Ӳ
@�7���#P3�偬���* 32���?�Ǩ��i<v��F��b!ߒ�Z��c���M�*x�ar1�I���)��m�
���1�s��[�Hݳ��K�p�O�L�����*X��'m�tu0bbk4vT|_`�@�K� T���g��$�p8���}��=����㗨����wl=��?��<>]AA�C?��qo���qqc�Yj�1�h����eCt�]�0"�U燤=�j�f�h����l�`M�E£��D���nӜ-�mg��W����~>��!�#rP���R)�������r>�T'� �눴�����[T�yn�]'������3�8E�zw\V��ղ0��4_��Q~��H�C���#��#9h^�iA���c���8e"�L�Qiske�-�1����:z��$*�*���v�.�IbU�!?��3��f�ty(�{OE�aX�̂P�v��v�}��F���m��wv�W�U׀0�eUs��n��xx�i��|\��@d����i��u(�B>�7ǈ�GNj�y�ff2v��Eu�)�� �o�Q�!hd>�Ǖ�[������YZ�-�-T2(؋d>$�JA4�k,J�c�G$!�9&S�RAH�������	9�CrI���1�WP^�R#1����|���?N�ёCl{��-dU�����FFo_�����RH�p�W��8e�������hum��#G�����U�!�8:�X$�Y9� lsj�<Ys�q�)���Q!�g�ɇ�4��uH諗��>sϫߍH��Y��T���T�?s�����i��a�����UuwYU���}���5����#R?�lB�V��^��\���V���V����M ��T,���È�����Q��ǈ����%��%��U���8��jT�H�a#�r��u>=�$ڏ7�r���>/Af7u��hׁt�\Q��>Lɨ�D��,�w��晕ToxE����~иvT��)�?u �Z4�/Tп~�hc�����LL���}b�>@��C���/�\G �껁� iF9%�: ����<�h�]E����~�xh�*J�ǲ�4O6�"�e+�Z�ʦƲ$O4(E�L��d �/)h<��N��pL��YY�S���_��R�-��mXpf�fn�\q@���|���(�s�$�(Z]@a��D�C�����[����U~N��b�~nE�m�]5�XL-��h�4�B;S�ք�1���a���5:����1���S�5�k�(nWѓA���F��}1E�tY��������e���-M7���j��������Q�_����hP����E���G��z5��n뻽%IނN��gF�x��)G�z����
8hU�ӧω]R�L��sv\��]��F�>�C(.�@8��	�+RT��T������wR���9�	0J�g�������z�~���v�cRV@Q436�� �����>1����x<�q���?伣7aX�����SUܡ���q�A�v�V"�9M��4}w����v���	���z`��F&������,zJ�8 �0�������&mE]Y��9��VT#��j{��扊�]_c�f���"o�RCa�sk$y��{��H
Vb�^\a�2�H�7��:R\�H![�]�F�5bw�J5�c|��X�Ε_��֚�s���y���$V�,�g�;�Q5S�hlD�Iu��r��	�mw$.���;�o�:�c�0O.<-q��]�طǏ�jYDwzmH_㺿1}�1��ڭ���!�[�7.���]2.X�E<�8�Z��.��>�-<l���v���z9o��~���|��.@��h�P���xy���ltN2�?d�u<�o}���r
��Ym�QQ����
�)��m�Q['`��}���F=ޥ��Dt�*r�,;"'�����>)�����UU>#L|�6X<�>���x1�V#��.�3#��`{�i�M��p8v��9(�+���|](�%Lxw�DV����1�!j>`q��]�Mv<5��|n���~��{=�2Xm��{w��=4��	�EN�Q�x�q�	�NSCxY���&�����fi"�,�6\Z��-����]c�~������Bvhx���&�sp1���|���b�زn*��Q],�og�Dy��6O�75f�T��ɐ.M�!�xv;i��L��+9z��,C���P����r����*�����x�+�WH�ݪg�#
�|�ɿ�|{Dn!��;4z�.��9mc�M5�յ����G��O���{�_Do�bW��X���N��������X/ߟ����pJ�
��S�)<?62�X=�s�mre��Y8 S�=��t��8�����;bL�.[%�H�6�9/|63`��@������9x�0KG��*����Yl�%6�vд�b�܀14���if���a�	�	�)��������y�]qX��b��Z�_ "W��
qq�m�k�4
Ǽ���ߍ�_ݥ��Z)����ف�E�&tネÍȭipY5�G�� �K��R��n��0�2�oVt��>r�q���3V#r�	����Ρx���o�b?ڡn�a�6(�I�8g�kպ;skY3�] �G����Q���u�K�,ΕQ���3��?�0I_2�v����X�L�ʃX��н�u@�u�m��ZԐ~��n���g$M�W{l�ǆ>�b~�s��j'���1n9��3Z0��)6I㕶e�/���% }�F�&Fa�į��$�����FI����੩Pyҥf�Ħ��s8����)����#�r4�U�$B���!�.W8��W|���m�{-I����)�F2&lk��/�w�Jf�b\0�W�OnTr���Et���������o��a*;�)�f��r�d��d^��}]�����[}��/�jj��(�Z�jH��sJ׭o�(z�kv�c����p��LM���hU�O������
���^�;Ӝ4)�y��#Hj;G���eyz��@���Χs�l���t �λ�<�S�����Mp�{'��Jk�.��s�J	��'ơ梅�) 9c_F��
E9N���_YB_X�����X���������w�?v���@�����ҙ�9;��j'4&�Τ�NO�Vc�P��V�p�l��<����]V|m�L�rO>�.�����J���Ѧ��p��>�J���s:j&�S_K���R��6�~.��X�)R� ��~v^��O��yR�2.9��V*�B�����:�ބr<"j|���Q�n7&-�YEG�Ƙc���dѨ$�5K��P�v�v��90*
x@cVއ�=�ѝ:�.�B�h���J�`=̈T|H�z�z(߬�]d9�&%
�ٶ�)\Q*Ν΁�Ӝ����i�~��l7{�w����4�=���/��Ic�`�#R��߾{�Њ#�V?�i5-�uQ��QV�#16��}�N�^3�e:�`�[F��BdƎ�|!E���g!S\����l|�p�PC�(.����,��B�:�YQ�M{� [ř�ې΂�Ᾱ�V�
�f�_^Ā��n.&�W�I�U�V�e�^E�՘Vkx]�����!k��b�v�ՉQ1a*-�ߤ�J��>M���IX����Ӽ�p�!n�X���7�I
��n�G9�B<��;�Ǯx�Bp2U���3��Y|��3��}�Z��]����i��Yj;�;
��C��S*s��ta��XN�H�US3(EG*�;b�Cr[�@q�)��6�]S,1�oۦi��s;F����a��i`>��ؘ�/ˉ�ա��f��>U�n��Ͼ�-V�����i8���=y����u������Ģ�Ѻ��6J^a�U��c��/��f|��h//x��|�p7�@�S��J֊&y�2���PS�0��b2q�OO҉u���eM��3��k�*j"ts ��5�9IU���^3�"��v�d&Uz��w��a�y^�������s݉r��h�ZT���oݍ�,%6fh�.ၼ#��{��Al�E��'�Anc��l��φX
 �,�̤����u���^S�5�]���@�����P�y)k�[e�_ť8h���`}fOxwƎ�9r����IL	�;�}���P_I7Y�����c��q�e�ϯ�ε��r��G�G�Y��dX b×�����XZl�Q�ݝZ�u��8�0��H}���5&:IH!$����	�� ��������*��:�����>n�*)��w��4i�.��]'cU~�
���˄�\������0�"a��WD�l�M���he���0��-1>���H�4&n Qt��t���Fƛ��uӰ��s�����rО��(%.|�����85ː�A��J�S�lp���Ug��f���N�	N�&j���*;PwO�I�T�w�F��fw؍2)�� �����_��vт���Ye<�!x-V�y��۞=��l<���_�1n��Ykt4��p�X�l��.�����̍P�:#j'dPa�v] ��rM���֠* ujo��U��UqR�]Y��n&w�r�c�y����RT�Wva<<�������!
���������FI�ƭ�&Up���fFq'�&�^~��p;��}V;gr�UCU�}Fۤ�\8e��0����e*��U��3��c�۶�"Ӂn�2��(O8�û��É?�=�#|���>��5��a�(��sF�~����+�:h����x�g�Lp��ºĢ���>�s����U���O]�T�*��޸����(gE�OyOQ��U%&쟣& DƤ�J��%�f7�xp���Z���4[�F�V���&y�!e�e�u�A���#0ȱ5����c]c����}�`�m������sG��D��g6�Cm�6v.��L���&
�`���x���嶜�����4��kE�/��{:��a��56�J�0ǳ �۠�A�
�E�o����Л�7���^81�����1�����`@ciJ]�����NI�v(��I�w�=W�������ujoS�w0�5M���������6"n�j��k`��̘�_.$���zӑ�з�B�S�� 9��)]7�bwi`�bn��I�d��k^_�s���V�������9 �'id�Ԟ@{_��k�撞�S١Q��nْ���:up�Yq�X��g�&�OK�X��P�{�eԍ�h޴b?�U9��l�0�����갔�z��9t��}���P��lN�4zU�T�������F��8W���p�x�Ð��A���Fذւ���eո^b�3�_��4��V4U��;�G�2��`�q�*���N����Ya�����r����{ŷ�,�*Wt1����(��o���(�I�#1"2%E����i�X����q��>�s#~�s�fv�l��f��`>w�EČs؏�~���k�YhS���V.�1�L�jZC|�r����Mͺ�V��J8_����e�
��%0�����3�2���LgGG
"���89+-px+?1j|j��U�������{��v�+�1�_E�a[*�5G� J���/��� ����ۨ��e�=��
)�`���!D���aq;�7+����2O�Gd�X��F{��?,��/�{;ѓ�J|P�����d4r�M��oR�z��w��7���E����n�\gqCa>4i隅����ne�~V!���%��|7ϝG$���y��ޏ��]���zz��,��a{΅���T�r�, �P�z�Q���� ��ᔾ/�"s�Ύ,t�0uQ�k�2��J�oqT��+�����Ο>�b�<ާ�@����L͌��X�b-�3�0���23��Lu_��N8�ԵM�Y�ۋ�����8�DE���	�>�j��"*m�?�q��|��_�:����E4H����:�������G�#B��t�,oc`��l�����1�|x�!�B�P�Ez���u�Ϲ�X���.n�����rX�'�J��ʡ��5|w��k���loC��6Sl��I�"��0���q�nh�a�����RT����3�+���__S��cbf6n�z���p<v �v{�5���.��	��%ػ�z�0���>K�b3������u�Yo�4[k/L��`�Vq�X`p�[�m���%�Q���}��@A�pY�Fe�
N�}�i~|�f.i/|���9-n6�%�)`/D�ls��&�o��
o�ڠ����wa$?}�T>m{��ki��������'I����=�S��:�RQ8�~(��ܧX�)+��	t`]|�ϥ��w{r��_ԣ�Fo������p�
�1�Q�8���o�7a@�//n��]G������I�����) O��e��F�i=s�|Q�Z�)��X�kB�+���G��z�W�dKf��3��P�~:,7��X�䩟���C�����a���ka^>�&��K���iH6ֽR�v�3၊�;��L����8�dE�7�~�X9�]w� �h�`�!�����]�8C_g%�bΟ�.E��kr����#�QY�@��E�H�Y��� ;s�DQd��`�)>��`"R�}��)�g����!��2#.�X��a]I5{HC�C�,��/�(0�:�&��Ո̾n���f��`�R�r�p�`|>qO8���)�K�j��/�K�hg�xK�H�u9_Ȅzg&_�u���J@C\�^mЦ�����n����������6��E��l�z�ܕ��.?��c����?�g<��PB8SлD���ě/U�$x��̶/}�0�!GK��7�Vjb;40Q���Q|�r������� N���&?s���5&+|��sf�9%��ׁ����P~���X��X�����]�N�g41)�E�t���uߗ����"l�������KZ��i�U��X�&"����]���T�;WK�n�G�8ͬ��2�22%æ���GFQ	�8h��E}���؄�-�$�����H��>����T����)������I������^J;҃�7��� |��t�TBG��
<N=<%�Ņ���ValA'��O�:�)��uF!M�P�:�U�����03;�� 
�FH�A<��fQr�Ŗg�]չ��#E�È"����+|����
����((i#�����T2����H��Ut��ɐ<FR]%Kv���{�����wUǲ�#	J�cW��&`�\XC=I _�����x�F!΃뾗��e"����cjCD�E!)�흨%l6O�@���i��b����=����v;�(&ng�$�~��b��!q9+���3���q�]�3�M:�5���FnX�����id����#�^�B�z|րlЌ�}�q/�zM� �Ѯ2d��,��`޿kd+��P����?�w��������Q�����ĕ�0�Pj�QC:z���q"(�� i�;���=�>�L���x^�qXp����ύ*�-E^�8����+9I����i�<�I6��V�%��)��s������	�;n�8�C�̩�ʡ\j��x}Q��l+�Y�of��#�+_��㔅�.�r��x�n�+Hۭ�c}�l���?IpeR'���UA���O���Kd�f�3�(REA����0��M�`T,��͈o�֕p��ƂEP���/�l�y&���k�������Ȼ.g��{�Í渏L�/lB�����_��r�RD��hH�E�1��Ǔ�Mx��y֥��4���S�:0`=�9�f��wfY��Q�<"�h*��!�s9*0�4;��� ��5���/g���N�`C�.��Ҙb��o���Y�������^{�.��Q�Qj!3�D��h7�l��Z �8�p�����Ok���1�W/=נ|�w��m�i� �IU���lF�:Ԩ4�N�E{��S"n���@s������HE~ݾ��A�G܄[�������q��4�K���D/~'��P�׬�ë��E� �Kz��}j���SL�L}UG8��-��I�|�ᨊ���j���_�K��_D�A��C�����?Ʀ�
�f(��l�+e������Et�Ӊ�g�����	���4�ќ�q	0�<l��m���8|_>���?�%�����]n�ٸ2�k��q��	��RG���Ѿf�x�C��)B�"��ʉ�6���!V6�XV�wF�KK�r��^�ws*a��c�
���pDN)?��s���?G ���oL���nBo����Q|b\�ˉ�XOo�t 6D$-
��I��G��n8��	#�$:��Ӿ�����@)�Ѣ�Gq{�P�{�S���sCW������sF�4�k|��� ^���B؋�r!����?l�{NF�y��k0c��� fW�z^ӛ^����M�jO�"�uW�����SU�Tp��o�EjSXY#vG�z72��8ȰEeK9oF��t�����n��cv$��7�s=�`Hl��$��b��U���B�w]ġ����+� ���	�'.<{i��z�JŃ�Kx��ݠ��T�!ժ>$�G�Ѐ{>�7�i'c�|S⫋�V�"(
l�M���>���n����>X�1p�QuE� �x�yI�N���� �y�V+�@�R�3��EX/�.sM�c���'���#k|(b
�v��ḚJ�UZK�k<�]]V&
��w$�� �zS��a�7�+U�T��J���p��g�u�e-�V!)�׹F�cFSYz?��ݴrY�"݀�R�v��g��v.R�H�\Ea����W�c�ָ_*=�g�0r>�G�X��m�0E�cdE����Z�+:����\�$�W��?g�m�K4���ځ�k�5����7/�<Ґ�m��b�ki�����	�'��1�6-à���V�1��`�_n^�R �EL��xJl�7��)��$�����&�u �������E������>���8�� On^��D�oZ�_��9B��Ak�_�e����!���|6""��d���g|�{�	��@�>��D��%��xE�~x�Plڢ%T�]���*������=����}~�EW����D��.�˔stb/�3��e���GyB�a6���Q�̠�.{�Tv��k��Q�Y��%ӮM�h�&��]I�67��v(�C�;��Z�(����ݩ ����mYa~1l\�N���\��E��a/Z�]Ϋ2���ꭃws����0l�����\ؽh#b�`�5��[�Ȇ��#D��b�F���M�M�/� Fa�A8��ѻ�F��?�vlN� ��J��O��0�����w׆����#lGͥ7�0[�i����M�o�%���-��Q���/�9����,���FzG����&v�t��oԆԞ���F?y���M�:�(��z��6��öؓ�z;N\���u�C	#v������?�����א�c�TM<�1f���pU*��;�O�|�<�@���ys��IA�Ɛ�#u�j�f�G�o�L@��xH�.���;���S���Q������ɝ�x>~����XGT�q/HGQh�!6�4"7:�ϱo\�u���k�k����J�P#A��E����m� �-����]�}��{�5ۜ@��\K[���J��{�^c��sT�)*�n>d5��M�Bլ^��c^R�����)eͬ�s�Q9�#�y�£����RY�2�q�LTݫ�3��V��  �s�>��F'���;�1&�*ru��L�4;rP��J���H��"|�48J� �b[�k�	�Q�|g�m���Z�PȄ��1�,5K�!�SDe<�[��ԃ�*xk��Q�2-��牎No"*U;gz��]�Op ����A͠BQ��U%>��y���pJ���o��X��$x{�2��a9G�Dt��C�E�WАަ6�F_���_�%x���o��?���
%`S|��q�� !{����ZӞ��pЁk�(�j&�ć͐���Р���+)L�*
xN;
{6��dq?��_
ǳ|�h2|4����Ѕv����O?��d\�v�!B7r3t�!�������4��r���3�qG����;��k�f*2<1{��y����`i[4�b��V�
�G�{�(�t�޲EU�5�,��ro�T�j4�b!���	��4��`i#Rub!�2}��|N6��||���ޡh��Jt��b2��"o�蠣���T*�����!Ea�T�=W��`���h����j
�^D�O���x��<�>G��p潮��r{�:%��yZ���k����� �F����H-v䂓4G�m���s�*�������'g� �B�.i�&Z���2��r��渉H�/����ɘb3,ul2^�I���V!{%D�` ���9{�M�N�^�Ȅ)!�)�?\Uཐ�춛�� ���q��s#�؀��eꆈ�#�EtD���)�+�"��*��o@4�Q �1G1�aՑ���d�Q��Rm��C�z�9�_���(<�ȳC�����!�@�"`��#ٷ�$�ً�S;R.S`�������$�q'^�slDA_��f�>�3�X��3u��?��|�E�4�L���xVq����0 x��R�NfY�����4��|f��Z�՗)4;��<�@��1#�q�h�>=1"1���ﮰ�0�F�ј��,>�H78�����.��Ql�m�����u����J=�aa�8��.3\r�i��2����b��j֔�a��e�6l3�(�|..�������(�y�4A��U�g���;2�m��ʾ���i1mH_KEU0@6��^̳�5ђ�
!��Ε�˙)ґe�^)۸f��T\F��#E�2��/�����9cm�͕�����?dDk~�!�i�w�P��}�/Yr�R	���0$���t�%6r�QnlP�9��e7��F:m��_J#����F�Bz�50�l�a�I��:��*J�G��B�}}�#��n,�ǉ�_a䤤ONfm�ͷl� l��(����f�c�O|��JLǞ��C����mT亸��5�����
,���(8����aHmX���Y���s:죰a8��L�\�&�{#�[��P�ʽ3�p����<) �h�q��.�h���{����N8��(��(8���M졯�ti���kvR��QIV�*��ݠ�u]���D@t"�}g�"Y�!2l��q��2(Ws��B7�he��!��m�`k�Q�%�����Gп4z��S���dH�ڽ��d�����fa�.�Iy�]kD[>Z�S�I)�GCU�A2=����tV�������g�dc����?����?���9ӀPOza�!Da��D}���JoI��=��;j��;��^9$�\�Ke\9z�Cј=6���1���C�5�
:�V.��^���ǿ!\AR�s�.N�=����x���H=s�$�����-f�G��;9�!�KAad��ܫ[�>Ԫ�0��?��׍�F�T4"����ȢY�I=�v�ϭ�״�N��#�����ݶ�����_��_�l:9��6�|�ݐ��!�֡��\�E�ֳ�FBN�2��Y������
G!��q���JY�]�P�^�7=뀛�ݫ��4�2'*g�i���R�y����(C���BQ!���c�yD;9��B��eI��Vڟc�gD�H�5�.��>G62��������5��rD�ۭYl㵘�?+@��]I����E��%���Q|�}F�-��m�.Q�����OGCZ~׈:��W0s�7�-,�-x�5#d�[Z�����$�k���]{!S/~Kϸ��uN�������h���D�G��TՐ�'��,K�ZS�I��}���S��KL�ޯ�e���a��a����(\G+��tDl��h�z 8�bWT=�R�Z�����z���r�����Ǝ�h���#��&��H����F���[j��$CȗSزK�W�*���l�_�F���D�%��F��F��ؕFM(��cT�}�.���ؓ���U�'6���t�
��}K��\�H'Y�m���k*k����Z�m��m��{�|iy���ಋ4/�Yc/�.&LU�X����l�y^��&+y�17E,���ܘa=���m�#D�C�jB8��LxW���\x��Z��I�������<:�m�>���H�2\�D���	�M�Emb���:尵��| ��'\���D�g�j�s�ܞ�3MU�ؑ�EI��3"�����9��ѣ!Y���AV���Ї�.�_��n�^.�Z�(v)]F����u�sSv�X�
�<�T���u}|�Ȗ!��[͚:)��zEv T2j</u�O}ya���х����Rq<�+*���P)�&�Gl��{%�U�T�-7~IC�H��Ydp�����q��+oo1��#P9Nd�1I�X�RGQA+��l��=�9T)@.p`� Z�y�=]�q�u퓦gV��f��QxP��jpDI��������s���`n�nC0>����t�.�}�WDʤh�l�3��窮�=�K�$��5�35��L(�Tv(V�2s�M�kH-����ڶ�h����>�g�pʄ�I��p����𷆴���Ɨ4�5��)jm���B��A�-��<Nh���;�f�Ζ�xc��N"s���m�wN9��@9�גl�F�!���Z�׸DJ�
,�uF��-�.2���$�Y��r�iܛ�s]C_<�#��$v�b�,���A�1� F���,������'��G*�
�w1����6�BX���|DY;���0�W��/5
�^?Iy���RU����h<*4�f�9`��JI>7j��_.z�q�D������P�=�ѽ�&����Y�#[l��|�w_���l�"z� kd�s\q�h�=5��Ҹ�)E�fRn��PN�@JU���J:��C0ӼK��(����8�Թ��(>�1�����>k�}�.<�۶�r~���mG�Ps�6Ai8�_�J���]��`UU6>Ϯ��_۲��������`��WJ�g5��\��������!U8�5��:�ۘ�*��Ԅ�Jq:Q�R���8�U*���8�A��7dcg��N���R����mק.$C	�t����)5�6��Vc]$�b>�rC����B'��r�h��H�>_�15|6+��J�n��Wg�gv���(���(��a��I��/�K�-���F�F?���"�F�0��U��W=�S1/�x�#���(�L��?��ާ����}*�?<k�'���t6�v�+c�,�B6C��2%u	X7�����"#E��ų�j�	{֙^}��"Rv��<0<>_���G�x�(7t��	�0F�{@����c�.'I2Ml3�����ԩ��8*����ݩ�Mdq�C	~�1��T�uU!�t�v��xiJm���,�͛>�J?n��s�L�oM�q%��~�n*�.��S4���p��|o�+�sF�/8��r����6�`q�R�������,:�Q��,b����~-����G�i�f}E��w��\����پ~��u+�, �]�c.,�����Z�"՝��H�Ý�f��g�n l�N��7n�n�~a�z��:Z)nx>DSa������kf�=��U�)��L��*��_��ѡ��va��;���M*��uP�@L�Z�7�n��������wQ%�^Rx���9B�t1|.�V0��Y������׿�sj,���$�=m�� ��8�(��:)�UQ�.3e��22u�meV�Cd��95Gk���E�t-�rR1�J�@b=�^�d�CR�z997*B�����`>���l��S�oR�5����7%�l�r���.�a�1.T�Z�Jbfs���8�Y��ng���T�^>��{�}{�/�{��g�kF��zz����0	GG'��y�g�V��萙�T�E�Z�2QڥZ#q�l��\����:�w�ŽN�sOS3�Z�mj�%g�����t65mM�b�������B�4�j�����=i"���'��d��cl>0����w��6��bg�>ϊ(f����{����I�*��9��mDt�����}@\�o��ݪ��`��_�dɿ<���뇁.Ɣ�x1F��4X].H�o9>i#*�!T�=����᧟��<P�}CΆ��7Cz�ro$�Wv��O����9�_��"�p����q��kC�M���z�9��Fx&S���t��o�$�
���c!n�:jzh��x��SU�P̜�u�����1GQtzԆ��c,ʶU�igDM�H�먔5SZ߻���N�~/��MS��8�,��敓9�hHG�6�\��)�(ڒO����:���9pp0�v'5,X�"��%�]0]xm5�L�!�w
�H1چ���������c�׫Z	4M�cQօ�אeT�^�`�׆s-�АVc�0�z[C����n�q[K��ʘ�)�uX��F�Ge���a�":���%�bPҮ�H�Y��;�qur�(�����g?���StP��SW��?��gu1Q���D��nݽ\=��V��(�T�H�� �9ђ�ަ�='��ip�H�(�!X�5���-8�n�� ��"��P��aK�1X�N��%6:���	�T���Ǐ[4�׈� �1�ʎ.�acA�	'��wW�5b�<�"n�EE�����0� �}sb8����@��y�5W-5舴a:b��!���������R1�ڡ����8"vZ '��J���GE--�t^�#t3f���}UQ3D��"�5F�_�U�4A� 	�s�cCm$�`0��:,o�>�s��l?�ʀH��a�=L�Ħ
������#��:nu�bC��m��v�5�;�65l�4��J�A��Ym���PV�`�)�Fu׆ϵ�ֹp**�!�
���ZC��������kXiS]z]h��-�T�ƫ["��T}����h����r�0����WX�s��Q�@��W�Es
'*����� >����K>W�	�"�SO/SO�a(	�Yxj$ �nȞa㱌���4�m��G���*��W��kN���Ew���^��zK��T��ZɿC�6ܛ�h]��r���ܣ�k�ty�4��:�;��bR����3�)P�q���J�x�߅!�/2�K�/v�?�le�z]����wKK
��h��mD�Pe@DG�XE�����`��E}�1��P�=��DL�o���f
An��Hs��@��AM��rM\��ǿ����|�@'�m 6yT��d.Ἆ��uy~� K�kz����+#Y���Jڒ�f���)jKhB9�u8ڭ��ud��o�G�<��5���-�vm�Ԭv�qi��b��K�����H�1ص* 9�����L�\*��"�O���D��"n�!:�F�a���}�#�;�]o�h��qxa��~��7.�k���ߍ��X���T�5�H��q{ߧ� P�t>˾�\?EJ���"���@1Lµ���9O�e�脱FS����r���EW|5���=J�7��!"Q��������Jjւ9�A�A�S���I��F{a�n�����Í�w	(Qj�f� ��0�\��Ҳ(W�
32C��E���27>�`A	��H�zpA�R�p��h��ܸ�C�u�$�q�����Fq	�����i�rN9t�����o$�wT��!�xk�m\Lgb��.�z>����p���n��,�L	�\"cq�4
|GR������<vb�1�P|�$x�A�km���e������:J�'��Jj)Q�,�������P5�Kc�+絭�8�
�`��X�V��y8��3W��q�Պ�:c��ν�j�����9���>�8�B��>��m;$�W�Ҁ��W	��ϔ,�HZ��8>kx�S��%*~�]0:m�(*Ǔ�ɹ|��Cy����)�=ƁG�Z��!Ҁ��J4c�%
PV%ꕶ�bָ�Q���%���bHL�#)���b�����<�s����n�^hJ�9��}:�P1�N��oQD
��CP��U���h5u������L*7�t���/�h�kYׄ[!9������Sa���E����70���P�%��S�Wi2%c�1IT���>;�@<���9;�n'}�N���p�1����[�f�3Z��c����%����z�s��[�ä|�0hr�O8'}W������Yc߰p�|-��Il�H黔��5�5�����¡���Q�Z����Լsb�����a7R~�Q��q��3LC���\���{���]U�ƈVVɫ��s���aLCCuI�^�%p"U�cFN/�f�J����;�<��m,Q��ν�:�Wx���)i�R��-=f<����h�k�K����|�%~��	#,,�~������0�:EdgC�CjH��?��vc��8��"/�匋�5����oN���f-a����a
6>"/bV�F�C�a8���O��U��lH�6�JS�ś@$���>���0<�n5�i"Q�l�Z�=0�g��*�2t8G�����)#�w\G�>i`�(N��cԼ��1&��5��Dq�T�#����(��
�d��ǰ�"��J��xg8���0J��L~]Ŭ����Nb/-�A�
�����V�˵5�a#ص:�x����ا��B't�4CY�Cn>�����3۷�g�=CcE���|�5�j��lyJvm1#����s%���*5��Z���z�r��w��s��m3�kb�SlT�yKV�甇:j��r���1�:��.	���<]1�qPtQ�X��p���c�ǥ�����Q�rS�UӬ�B�9j�����EЉ��b/�1<�W`�2�{)�*�$��d�5����5}�WD����Ƙe�
����������mh�z���ύ����P�f��ʄ�\4�ё�e���e���'����և��C\�1ו��"�Hgȳ���z�~�6IO~��o�a��L���EMF$\4��ҍEy����Θ��5'e
+��p�H�w,ʌ��<�N��᠊��^G�}�u)������!�+��E��k�a���Y����G �0��(�e��3��<2�u��
g��aB~�g�M����q<Qt���0�T�z��g{�N��V�X6����3떵 d\����(OL��{ ���PE�wwb��湫�x���N�*Q� �5� F�7���H�B���U��32βc1Ѷ7َ��7Bg���Y �_Ү�$#���e4H�`�=[?��a^.M�_XEc�Y��;
3�%��}]�6/L���t�P����샧!%�yP�y�1���k�t��������KM+q�P����c#�2hM��Ҷ�E�H#t��cY���0�Xj�*]�~�t�4 _oղՊx�)�\�#e�(}Ƶ�X:Z�l�����4n��|nq�S \�s6l�Q?ߎ����a_2��?���TK�)�(��%c��Q�~��[��^Όt<�.��ƴ��$��=8����bةӈ�o���q�Sd]_�7߈n�3�Z�X�ZᎽx��q�����C-��߉V�}n�~��r�<�B�`�|ID�떽��w��
��m��� �'�y�~S�6�X*�����%��ض\Q|vR;t]����˒[o-n�����^����E.\�1��������Դ����BMU��!�NېN���Ey����a2'�*��m�����9B|v�H�p݄�e9_=c*�Ē�ŔJ��'Q8AJ��%+���YS�Å�1��ƈV�j[P�:X�rT����.�;�T�K=�X2�R�IڇH�Xǃģ Dm�K�T͘.�#��K���*}�d�"=t�j��~f�ib���9�������e���K�Y8���^l��������������&����w͹-W�=���r�b��9�Yd{ v��8�ʴ���	�]��y�ǐ$�)zF�`�9�UD������N�����$�M	ju�PLs?>��������&���Ü���n%�|�0Ͷ����Zq~�E����\�#��w�J�m��.M���(��6���o�?����Ra�Ɛf�.pV��n:T�4�um��i��Kf��i G���������ʐ.�������&~��aeQ�[�|E�����{+�e*o��5��`�Li��T؁.�vx�w��0Hla���Z���������)&-;Z�"�4��
��m���Ez���O����#�&��L�_��s�: u�W2�Y^����.G3�����؝8�,����9"s52=|צ�pv02�ҫ��%[wW�u}�<|P�qc�l&���3��Ԍ�0e�B.�M����tɴ���£^h�k����&#�a��9�~��lһB��5�p��F�D�0:���y�ׄ�%��OZ�܃`�㨝Ӵ��v9$�Φ�x�;Ȱ�ӫ7>Z�߿w��,��9z*�.��M]�FѪ��P��0^���4R�`���Q��G7�T��s�r�kg���:(z��BSƱ�=��@`P��5Y�g�����`\��Fwl�6"�ޣ�`���T+CJ�����lL�N���Nݼ�7m�^)wi�Z�Rww��]�b�8G2�b�K)�*��w٘�na�/�����K��8��8��a]���%��ُ�>n�|���=E���i\
b���
Sq��?��������8Ɵ4];4��j�*V����nΪ��Q�,�ʄ����կZ@�+hFόrMq4Ƕ<�`���H�$7ϼ>d�8��~z��I�`-ZQ��X��Aw�Fqzk��+׃�#��eD�x?�?�!�/�G��t��
�7�7�f�{�eUA�K����]�$/�1����EY�݆-�eJ�.���1P��.��������4����\ڗ;v�X#t��3ɸ�'l%��U;�:q"Ý�u�/<����>T�+�y9�$x�j�&����{�h�Y��{��U�梳��Y�o�0�k��V��Χ����x&-��i"��)�bФ�i<S��������+S�J��K[-+�d��^�� ��6�� ���3�gZ�T��+��I�0�vZ	�莉�k7τ0[���?�T��+��mX����?�1��ɀ������Aaq��W�'�B�JX�$��3u����"�/���S�ꮁ5-�*]J��}z��4e��&]k���؏Y����Kx.�o#z���u�:���`�S�o��T��V�S%���P)P�o��>3�o��5���\&RW<Kl�S̉���B��H�$F��!����ÏL}!��h���ې�����k�[���ܸ++-�&��JIL��x�1±-��@c
��V�8�)_D%�����mo�e
cHq�E���v���7Ulb�Q�#�UN��1�I�;C:p�F�F\�����=�R������������K�{��Z���s[�~�����=ᔝT0��2��h`r�,例V�!*�>C�Wl��/�k]9�Q�a�N���H���!߼b��u^��aԆ�j~_`IA+��%�OG$�̇��xP"r�b�aېbct����b���}u��*IO�q�/p��N�yD��]PS)�!�r�]1=�	����t�CM��M��"Z�,U4*݇l���'�R����?d�NX�u��ȓ�a�HPn�V#}:P��|���TԎC��w|foB���������H_w�v�((�WA��L*6��.h+m眿����T�	Ro>��C�����M�m����g�S:(8���.��1Ac^�'G�h@����}��"�v�������E���Kj�"��P�RC�(��OI�0��~�9& �!aV���d��ΧT�
]XQ��ap�{�>)2�|�8{��߿�.����%��Cf*q�t�~V<7���
��}���:s�Qʣ����}�
��َ���y��o(rȺ�hp�gv��Hw��
��O�`�)"M�yeP[���!�
���0�h�bb�!ں��E3
 e̶+/��EqhY�sF���Q�
3-<$�go܊�� � �/�i��ӵ�$�m���ϰj�b���,��97��c�͚*F&Rc��+m�i���vEE�~>G��Q�����߳�c�Ջ���ܞ�Z�9ύޟ�\���Y���g1rW��Ey�)������Q��C� ll����:{#���^�!�����������g~.j���$�b!�p�p�۟�4��s:9��X	\������P2�3�/-�q�J�g/��If�`6K<f���u{�{�DS8,��(Dy-�9ܩc3������l��A�d��)'@�Ό�y��0d��킂U�2b��~���Qd���-��Դ�g X���&G2�M��Z��׶fd�`	�Fm�OO��4�3�g:�V��>I���+���ؿ��ʘ����*C��q2�����(��k�6�N_��0�!Ҍ��o�Cl�/�=�vLEU@J+�0�fK䔅���/ײ!P[<@�8.����BU��Bd��h�"_����`H���S�)~���)6����,c���#a]L�{����%�d��Y84PE��ǈbD�6�V�
����A����N�YxF�ka	8��(�P�����5�k�t�9�o���82����J���
�G��J[]5�޴}����+-�#l����,�jc��~[������6�Wl�.�͘2��BY%h���X�T2<Lآ�q��J��Nb�i�x3Z�QsИ6��|#������W��+f��k�jQ��]HE��ߚE�EQ�|���x�������W��~G
U����1��N�*%�<sg��&gO���+A;b�KuK�T�5�/\��Qo���Ҽ�kkgۉ8�0�cL�~:?��TzU�����׌EK�䓐����k�Y�Y���U��:+ƩL[Y�f��~��-���&�
� ��x�yJ��+�1#o^�c�w"������/�ׯx�=�؊M�L�u��5q�)g/`<�[�?���k�q`^H��t�5��R��!��)�gX ���-��JSD�������.GS1Vcp�ךl�`'\�Y�G���'�͈��z���@�\FWq���w||��CJ���R�$�_W=+��|�����qa|���o��}㮹V%�ڜ:p4��o�^T)��*co=I�_Q@Ѩ�4<����ϟ/q�0~�&آtD�h���_���{�S� �=�7�nnoum���aH��Xs@p�X&����+!��Cb�a���:*r�\���pMk��Itl���nc���10�2�o�O���ˈF7��TI"�=_2��Z\�{�g�P[0�i&��cv'����/�p
[�������t�qdT�_b���̰�ƠS�=���f`��]`���Ѷ��i��:o�r�g�o[^���u]W�j$Q�W�au�``��o�;3��(<��0f���Dj��SG�z�����X�>7&�(6?Z6�{�ZҎ/����2���F���#����Q+�6>Q���L�`n��rC���v�QTI>��e��}�x腧y�Cd��
�'�o�Se���۷S���=z�G"g׏��)AHѼ?�F�b��0�P�K����u�A��<U�����*>�W����� �-e��s��l�5�c�7Ñ�"zrKY���(���4����8	�ܤczU_�B��6��aD��3�/_ޤ�h�tQX{g�؝bf��q�:�IB*�G��YY5Ez��O�Cꞇ2o�tzǮ#�5on�e����r�fe��;�q�nG�85Vp��{5
l��ܥ5�jᳲO��9��}	���q�>vҢX������G;�F�=�iHj吴��j����������U��hP*6����z���v\��fm��+R��v��g�]gw�,TO� �'[�YP >�����1	oT�e��Y{l�������XI������|<*��l>�);R2V�y�JGZ�K���3�Iv5r(N���j�
�ot�*)���ذPN��DD�p$��pz��������Yx���UX\�-H��	��r�Z�I���i]q�Qx{�bG��I�:#V�ki[l��DpU��t[:~������Sg���ٙfHf1`O��X�7p�9���1Q��5�������=��a?�r�^�|��}���V�z�kA8�;>踺[_�c�e�Z�FWw�He�=��]-�1B��y\�?��V?,���Ԩ(ΖN�C���������g38pga9��[�+N�.��>�ښ�N�C$`�P��	Y#
{/�#�fM�n-�����Z^�F}�L�:��l�R��Y(��U�4��D6����'4���4���oCꉄV:g��1Lc�ʐ:��C8�����p^���öpH_�jm��VT�����}���\�W���DO�,�͛}<\OD��q.���N��Q�{&"��^iڭ�57����|��)9���w���&�G~	��(a�ۜ�m�⢖7� ���>[U��r&����S$���/�Q��r��"t�)����÷��׿���m��c�P����!՘�o��IU��Un+��0z��W��ḏaGD��te��Ց���<���U�o�A��6�:� 9s�6�"���^�I�B��j��v*�KF��|�t��Ǐ��o%����,�d=ԨlM��=j���a�!iV���lY$'���q��3攺�A��U���3�����X��y��[e���[ɴ}. t�a��yP�7�g�)W8e����1佖�6͸�,t����C�_��m�gTy�|���=�`�Rk�cw�P�c[�%|�\9]g3m�i�vMD���lH�hc*K{���� �a�`�ݾ7���jn��vW5}�qhD/¿�0��.r�u��i��}QD�N/��m[�W�q8L��{��`Q-���f{����5"���ϑ�y�����P����hq$���.vo�pDц�| ��~���x��G\_T';�0A�M�*�}=�%y.�X^(�oF�0��_E���A�O��x���өR�V�^�.��m]a�at�~�	�l*�#g����<(�h�Z�H��@cxNV�U���u�G�A�e8.,�uP���%��yxV����Z��C;D���{�&�d�{�&��=�m���~'%�7��G��Zo��81f.���
��W��bW2���X���";6����ߢL��NB��7�����������3i3ћ����i�k�fs-�Z'�:�m�:Z��Z����K48j�B����N#x��uknq6���ڐ"�Ҍ�*���߷α:�ׯ|�]��F���kx�*5��nE�f:0���}�_ѕU˿��/�=�h�T񬓢�I"kfX���x)x~+��z��rPy�+���m��������2�q�cV��� �RD�@4���!|���aR:����´(��d���a��)���9�'��p��B��u1�����:iL��^���m��Mό.�lP�^�[
��4���V�R
����!��`�J-��B@:�7T�w��a����Q� �?F-�e���>|H��g�ɑ�SJc���,nr�f_����u�D�x�r���xv��˶�,�}��)X���5S"�� �wq�`�#��R�pQ������	����h�8>�g���|�=�B!�a��"/��tvq��YHњц�@µ�rڬ@d]�L�����)���gB�i�?��x(�*��Z��%Y\��fc�L���|��5��2W!�g�3�{���s��&Ӽ�P�z,�-�-�\`��=;�\��-;��g����&o���R�^�{�7���,����$��:̗��������t���E��\��4�ƐZ?󠢏�ۃ6�cx����Z�:��^�9�ɒc{)图�$���X�m&b6�Sd�(�5�/��- ���n#FZx��xy �:&�=�ENN�S8��tqAo���#��"�
je{υ��"���3�)IG�İ�kO�(�F4��u¸X��a;4]�$�Vi!+��<Q(�{詛@ne	'�n�)�dO���׬��|}:�dI�&�����IǊ� ��!b�2܃��I�YP�0�œD�Q��sG���xO�f���&����k�����dG��XDߊ���?���B������m�c�5���P�J=>�>���uMO��vԅ $���9`p7S���p��?������������	��)���e��(�m�ÞY8/���\ �h���C%��p&�\�fH���0j��$�n�c����U!(�����>K�"��4w�ǳ@JO��2���ߔ����n����������!��$d�P���Rw1b{�ϝR�Xh=���6*��ۛ>S!�$C�kϼ��
���i��|���Z8��d���N��O�x ��M�`��zj/\#R
�Vc���H�MC��t3ZOY�;>��_��9(}QU��ӛ����}�Q%"RPn���6j�W�� C��3�Ut6%@����%���ME�����L}nr5_4DcFw��(FFԩP�!�c�z:q��t̌w�6����혃��x/��~�X>n߱��"��1t���fd롥b�eb��F���6�*���áS]gdD��������%�����!�Nx�h�`�����ֻ�Ю��N��b�TD���]���y;�CD���}C gRz��PCFo��_�P�:T� 3�,��p ���g�PO��w<[���f<�ƠQa�H��p��9U���Y�OR��5�p�`��U{2^�"�_qJ�;�z���gOT)F��N�QD�8���=v���j�3�NȦ?���:�)�[����{���������j����ٶ0���p���!�� C���
1i�3�6G�$N)�ߥ(�(/<��0^���V���|�h8H5����,��ssӦ0����c<=�ʢ��N��/�`z.�3w��7Ґ>�τP�p�Y�7{����3��ɰ��{C�%��?��]��O��s.�=j@*�G��}��k����Qtj=�S0�Lw�(��q�MP���n����t�>c��`�ņCH�������͌��'�_��.@�� B&�M�{�R�IŦ0 7��z�����.OrJO�.ra�b$��$�����P'cZ��B.���>k
A���)�`��6�
���=�o$<h��$�{M��Ɨ`���b�zZ �jd]�G��g8x_��(�E�Q���R��#����e��nʳm��[�<��Gz�>���X�s�Q=��~_2����U�M
��+���H�F�=0 ���E�ޭ�Ě�4��%�َ�[�] �����~U����!�?����������ar�Z�H�xE_�g�ϵ��bŖ��ag�
��T�}�C���kx��������U�=�|�F*3�2^�,%�06Gͮ�!��K��Lq�,�=9��z؂O$�u����gUBe1�MnVu�uX�H�P@��E<'�/��a3�4D�p�f�7��gB���o �X=�R�������|ԍuk.7u`���#�9�"�nN)d8Jt#���|��))Y04���}�r��ī��X�(�B6�g�5���F������K�Q���6r0ñH������s��1�A�Ն/;^�O�&��8X煎紭/���11�m�� @D�1|n�����[��h�x|�s��
a�M�)�����SMad=��E����͈����hT�����a�ʎ8\.���b�I���)&�iL�����PѾ�ʺVA��{|s'�_��?�|X�@��!��[�/��+!�����a&-�
��Ws�[H��7���6��� ��!�hL���^wJ�����D� m���|�L�X�*X��6$��`QiE\��UԆ��X�*
V�؋3i��j�F=>�	�G����3##zkB�oxﮈ��H�_�c�*⻟�E*��Pf�o����{g�v�j�)���`'�:�.���ھO3)p�Q�L�4��Tz��gu��JM|Y�ԶQ�a�.�O�b�q/�쑽<GV25{`I
U]c���m���O�i��r'N2��c� Gnx_�ge �n;�̈�����눭�6ď�~��&�`r��B�i3��x�����)���HV��34�b���*��?�J����Y���?�n�n��Jg�[�W���E�ׂE���cvΠ�٦;�AsZ��0��gwR��t�̕�m��5#�H�\�(���bR��B��u���J�la�r�ºG}��W���|����«)�X4jw֑��|���!��;y�^�4�
O���:�p�^��7;��}KqW�iL��zᪧ����E°�]�`�zHgR��KVxp[u���,��%��.�zH{]��ȜE��e;1�VMTI��w��d�`a�6X�Z&��t��4�Yh�h��� �0�`��^�����oj��� k�rVЇڈq��E:x��>1��QM�F]���,Mfõn�Gv̽�r�d���`uw,�R��{�VZ�,�p�օ�3J,f�ڨ᜻�
�	8a3�!)�7��Ե\��5���L��=��+h˸�,)��$#�3�N!�����`���H�� ya!�m^��s�0/^�fʰ�jo�F.��/1U��mqyR�S|m���~�M4��]�د���8;�2�XG���eh(��k�W�Tȋ��A��>6�E)}Ua]��I�!-���.,#�N!.UϏ>#b{�*��w���Pa�ޫ���]w������$��W
�6c��ڰ����0l��M�H�������R��(�C×�T�b�&�:uyW8����*��i�T�Pp6ǠU�~��`&j�IX䋠	��{4��c��:Q|VpJ���W����HX#�U�Tald�Z�F%eb�H��<H�Cq�:���u��`���J�7��FS5�S���Aܠ��N��=�*o�{���r\��p0�i�C��#��ߦRQN�Tm>�"* �׺T�ʮk,C���:��PÜe���C�L�N�H���g�hI���t=�0�3��̈g#��6���i?�yҨ��)���g��<'��j[뢬?���e׿�}�\b���tT��v���1R�<0G���>�g�lT���
�A�_Ԥ�@��ʨ�^���p�y^����R!I��gD9��CE��D�I��Ln��Z;�" ���$���t�(�d��d1�*�}�=��:{�����,���֮��]��j��C\	�,B���o"/
�,(L��Z��56x;���� ��M��DF���r���F��Hv���Dqx�`�®������ ��r5n���SD����{n��=�Q��\�%��)�*�k�Z��ǁ����p�E.,�ݾGwu�+O��L� �z���cD��}��u��D�^ p�|
?l��Q�3����K�1��R�t�1�V���@E-*Z'�SV�mTa8�@���"���g���]*,٨�����UZ����Ru^�	�&�����O[��*�� Қ��Y��`A�Y��M0~�k>�_�b&���ohL��<v;q����ғ��d��ض��-�tr|A�E]>nZG�/g�Ԙd��),���?_G���h���eY�)n �|W��-��Ϡ4�勶�V0 ?��$�>hD8���;��Z�6�v�J����g�/Yg���g�H�q��;��_��C��������P��⁓b����a�Ԝ�q8̫�	��F� :��Z3ӰIe*P�^�Q���Φ��&I�o@[��Rj/���̒J�^�%���#�a$�h���+5�,���h�y��|��C�3��_����P�Gѵ��9���8�������u�6Ɲ��48��P�����ٹ�PS%\�s	���Y4���>�c��"4�|,����u���������� b,���B'�&'����黽����Yi��9�f uI�S�(���U4�l]�l��+��}��K2=�o���Ad1Ǘ�h��2ژ���e��0�s��>><&3��t<!�~�|e�QPTÀ[X]�`��ʲ�\�cD���,�7e��~w{.��i x�b��ߍw+���,�y�R��ciM������̕x��d
1	W\�8�Jb-R��~�i��ڧnWuz�����~�S��\IxD+�V�j�u���r�ݏ�$�wHո��,}�gʴ��0���ƮꝢ���'H��*�T6���3	4��6��ZuIE��٢�\�7�V�T��^s�$
%�y�eW��W.�"����i�5���#�7G#��Wb�h���1��܍d�h�Lvn����Ү�Y��.�l]��ਣ��g6uQ�`�[�Y�I�84B�9A��2[	����٦���#5Ӥ*&��2/�qn���:�X\�m�'�5��K@\h�(�ptF]O�4�\��(���_5��f5h�@v%)�������A��0���0˨V�)N�>pj�uW��1�Rd��y�J���}m@kP�}��;ӟ��}U��C��DJ�y@���Q#-*��e/��l�6~@N]��!.l�N-$�i�8,��]·�b���U������,"�{Epm~[��o����V�*ks>I���������D��$��е
�8����=�p,�zϵ(��)��+�ު1d1�tG�^7b�y��^��%�ܥ�9ش0v�S���*k��Y=][Ȝ鹐�y�H
�9���Qs�p_�U�R?E�?O2�����DǶ�Q���.C��,��J�M��3/�ERJ��z�^;�fUosys�,g��Eσ�7m��i�^w�`]�Ί��ϙL���9��nG�A��Q�c�%�*��ɧ�Lxl_�b����瀱͍��j&���n!o�uP�h�g���ʛ-Pfٌ��s�H�>F9eቒwt`7��� V�̵�w��ۛ�9..�lN��^Ic��7>)�sU�k�!�!����K����O��ّ~PA�?�"��*�ϣa+�Ur��4�	�q0gW�fzd)����h#��T�_��I-02�����fɂ1B��o-}��V��@9���"6�1?4
+��|�I���)������H5��H�A��掂��\�B��k���~�(�?�{�0ɪ��VM����:��E��	�LeKnzٗ��7�؈-_r�4��Af�ScHo5G�k~z��L�}#EEo3���R�� �q*��R�HэtG��!Z7a�M�����X���	dj	�s\��_�hS�d�Ds�v_w�SR�(!W1C|���D�=�>�lx�:B��n�eD�Z���O;�6�\��ρӆC3�ϭ��#���cm�Ta�l�#�V�!����-�S�g)�=%����ۚQ��>2O��=�%���,^F�x�f���nD��0
���d�D=�w��,��(�jR�i�	W#�
�,u�c��C#�}���\D^G!�F��i��h8'a�-�o����Z��{�.6���/�{�ƽ��U
A^����z�ￓ��$B���=7�j����j��L]m���Z��{�#�������헿sV�����u�u� 1����MwȔ�r`�8O���s���:~���)R�w�mh���`uޝ�}Y,hR�/�q�hO<��y��p=q��ϟ�7:M��^�1���S�(�#\c��� �w�4�5�N
�i>�$��y�gOu��ta}��f�13�H��b4��3�MЦّ�j���r`��4|%��q-��5FQ�2B�՝�
�����w��B����.��֢C�*��9}fPQ���L�o2Ev!���`O���^���x�蹡F�!c�#ڻ.�]na��N��h<>����N�t�1B/�(H.�:3�\T:���	aͭ@gչ�s��26�r%3jK��Φ�+��?�-A�g���7Q\�,���ΐ���	��!�Ñ�K2�)�4�rVG���<{�~c�DP+���O�p\�C+^K��T94ǎ���`����5��m㌯oRdG����>��{a�cα�sJ�L���Do��K[�9;���h:O���Qɸ����V�Y><�I��Na���z?O7�B���x[��U㑓_���ϙm�P�މ���1�]U��?�ӡ�cB��D��I�b(��=�����?�9.�9Ee<Z�wWb1xQ[������*X)�xb�|��f��8)�����(��l�҅�>}��&t�������$Ir$�A���!�X�{'w��E9�[��ú�IU� /�T�ܳ�g	�%P���UI"�����T;u�M^7ͧT͝��S�v6�!
W$ ��K^'�[���0��x!�ol�m�F�-����ٺ伆6�T�h���n��{WY"���Y���L��Ч]WI�	�Ĵ��S��6{�Z�z�5]��?R�n5�oGW[�f�m��e��j���?D�XW7;�m��|:s��D�f)����0��I��Y�� �����Q���t���o�U$Y�A��r�����\`����T"jU�=���uLA��ٜ�Z�StR1X���+�-V�u�����7\J�$�s�PO_��I��sv�]L����ٙ|m�)�{��%ϗk2)<R��."�[���ok�E��@�~���l��K	p���K�K(����D��Y�P���kl(�����o~0J�oA�R��Z����+I���ԓuO]�Xx'\f��;꽡�o��q9�,�m*9�I��ä����A'ԒX�1t�旬�"�?���	�����c��`s�m�5��I����Nt�%7<�ȸcp�z�Ъfr4v��tM�q"�1^W�X�0����gz�0I❂]����C�77���N^QRR������4��U������|6R�aa���Aa>��߼fSg�;��M9k�����\R�d��0������?q�(�v'�O-[�"��Ւh�x�!�a��`@�"�}��hd���}�s�t��n�����R��93H`�P����.��#3�s����r��b00ëzJp��Y�r��둄xIZ%�YT��Y�/��+qY
�fY������O(\nY<%��P���v)��|�5��E���^#kEV����[�A8�v������г\�{C ���3��������?����� �@ښ,����Q���)C��:�\9��� ����E�����B��|;��I�q@[��h��X*��;�׊�jh���)c?wÛ�T���p k=?Q��u�2�C
���]��\g�R���d4��ލ+�d�Y��
}��>Őz�F�)B�Hp���?K���/�������5����s_�h,�d�L�{{]������6#�n�0��y��=�χ�ڥk���R'>N�N�Y:�}��C<��3�Ň*(��Q�$�q;�[)���`@��H��E��N���������suX�B7����z�:-M/4z�f���NCe���.��3�Iy����{��Vٛ,��0J����"=���̒):����f�{�N�m�p4���Մ�~��0~m���ZC,-��Ž?q�>�φn�kf���,J�^�q�=L�[ēu���u� ν<�,;SeJt1�������:]���bzѸ�y` Tx')w��c�㐊��*�vez˼�i��#�O�>l�Ǯ��j8��r��38()���4~_;��>�"���{OK�[}��W9*�Qn�W?���!�U��eҳjH	{dW<O�f�1�B�z-~��Zu���������jA�[2����6{���6zv��6I-��4���������Anu��� ,q:��k�/d��dwFy�#�k�\JInT�75o�	���oj��
�Qr��f��d�[b��;��m	^6qڬnP���7d5fI����h���UO�.ac�xNf���@\E�)g�)yt/O�`�ωa�=�9{�aC�σ`bkl��c� P�ȩ�l���Ǹ� �c-܎�������j�ۍ��a�k�#N�^��{:�)8J�g�wg�$VAq�Bț��5�T�\P�c� ,��5:Jڸ"��:���3iY�JL�RE@x��u���M��T8dƳ����΍{X�JG1d"�� �m����R� ��盰�>�Hg\G���*��\\P�
1��!�l��Af���|�70]̕����p�萯Z��L��[kS�+Q¡�����g��A��p6[_���M�d*��F%h�_��z������:.�1y��t5����$��T�ә�#�7]Ҙ8I�@�gJJU%��%��u7�Et��l�e��r���@i�����p,un}Vv�n�/wH]�Ō����xA
]ɽ'���
<V8dC��OĿ���L�:�������j�_ؤQ*k��~���4�{�U�dd/k�Âl��h�? ��e��]��ͤ�P����?�6���w�^�ǟ����g?����a�R�+�l'�܀upD��>�;�#�|I�m��z�v���Ի$�� ��4����'*�y4q�T���	�����9�aiH6a�V'u��]��PL��B���M�q�΍��(����*8g�nd�����q�=}/���B&�2ؗww8(���[�^�(���~[޽}{�_��1����K��J�ВpʲL����1#��*h��bY����e�_	������������l�v��O�/sf��=}@_���m�q�s�Ѡ~J_��I��J^��^�
4�`[��y�n{2��A-r;��QP?|A������(�_�.͜�"����]RJ���vWӣlU���v�}Ԓ�A	��0џ�����8	�]��8���|-�E�L���۲P�|��>����pk��.���)H��9�k����b��@�z>���c�x��m�F�/3ue"G
��W�)�k9�h2��f�/���!3��6��	~��L� ߌA��d�YpG�� �Z][���/MSeT���2m	����7�5�eU}ӹ�s�Ʉ�F����ymtU���&�M�R�E��bu-��GPe��9-��!L뗎���-���a a�p���ļĵƇ��ۯ����q;�?]��v;�/	����y����4��8W�y�
�=�N��e��0�I㩋��T^�����y�#m��R�if��'T��3�~6��7ֵAo!VڄX�(B5~f	`���;��a��A��&d���plb���i���ٜ?��+/�^t��qZ����1S���X��c��[]@���Sm�7�^R�E�#�#5XvM���P�l�x��t"W�2m�ʷ��I}�b����~4&Λ��28BY�G)����.���36�2�'�k��,qLS���	�c�����Sl����{֤�����`Q�ȅ0��@�>K�Ž��%~Qg���y�sjW�g�n ��NB<X�$�۷�$*���g5A�����E�ƀ�q��3I��	�X��vx�"�6�˵wD�m�
��a��n�� �S�O��P�o��8�'�Lw)�X� �yY�{��p��l|Ο��T��kHEU�0fՁ���G?�0]"�;�����[�1
�O�@+Z���&\p���p{h���_�r̬��cm�O���뷱�k��O���	o0�1��x�I��@��:�q$�))3(g�.���%�e+ZGV�'Zk4�P�X�ռLE��L�d�.�L��}��[[j�MZ��7�z�8��<�k����:]?�؛����=�\�:h�� �-Ⴌ�c����X=o���
�n\8�� v�h�Z�z�I��:����9A�߭-Р��PUC6��]뫔�����@9~���9�-=*��;6--��~v�=>�PY�&	��B����c�x����F" �-Q��^��*���m�g�����O>~�����-ZKfgTII>1;�Q~v@>�q-�����>�#��:y~��������WƈL�q	x?
��#�H�O�)+.R7<���?�esp�S�Z�;�{��� �P��o�>Ӓ�ن��6��X��sR[��#��/�0C�x���e༭�M�o晘�l���ky����œ���~?;��^	#���%���N��D:��M�����#���$?1s��j����YiPḱ��A�����T�K��Ms�r� ʇweN ��y�bë��\�9�̝�6d)� ���9�����a��i�P��_��Jf��u�AT�#-K\�Էg�'��_C�� ~8شm|c~��?�{�X�,Ec�Ȼ��Fn��02��/�C��z!�����pc�Z�2���P1�-U�ą��ZW3y����ohM�Jpo�^�=>�ԦD�����!�?O��4q�$iG�P�E�	�E>P�~�����s�[ЄGE�\�e !�zRs�9yӥT�	H��B~̊M_�ږ�s��Z��� �i����$|We}��)s
gџ�/��*l�I�G��I(�3�_�(��=�`�'��蹾�ᱝ0�\*��u�XK�g�ݲ'��yk1����Wk�<:Fj�uK�Q+F��;L�p���d{����D)���C,��L��L�]���*��4��,��rM�RN�5���M��t���Ձ�<Ek��c�U`�S.n,�����P<�m/�K<�'I��C����{�bv ���(�C��Ƶs�i��M'4��;f��C�&kɿ�V]%�;w���r�y���!��/I/2�%(T*�=gtp!5}�y��O�'{ꬮ7"/���� �=n�.��)�(�E�����Fz=�#�inX��]q��>is�ڒ]p�I>���O��x �r�j�k�qU�n�8���Vý^����m�A,���ג��7���qh ��,^�ߺ�h���Xy�x�dR�a&�
�H�@�!a��j=�J{rS��K��2�:9Q5��S�Ow���Ԁ�eD8V��V{����f�-�؋��R�����������ޔ���c�Y��V���	�褍�T����
&7E��������;��2�Ð�]����/ ���@Q�6�r�J�^��Z4�2�y�ve�ؘ�d6�
��A�ƭ��+5=�n@n���79Yn��wO[J@��*J�ꉠ-e����mZ,+xIs?�s���'҄>I����G͆[k��4��������Jn�)�2�Y'�
gi��j�A�����k..,mw������Pm�ς9J eR<<���L]�eS�V	���s�69���I�E0���2�Ku}\����j��^�a`++Jq�����<�q�;H��A�b���-�:��-5�z�,��G�E�	��O���t�4֘���F&���6&�SP�EC���	����&���w?H�:mu�C� �Ȧ��c���������\8}�`ڐ���}.��q^�H�k��i/�
��k�|+_�HM�#�jM��8%���]��&�n�s�T����;Y��#h��#��߸!�6��v��i9�X���@let���^�r:�hM��=��c�����H����k)7>�.qPB!�>�bH��2^������f@#d'ZQQ6�e��b���f��/ZQ�f��G������97+~���c,�m�&��uv�F�ۙ���	Q~�Í�k�m���=�q;+�IGԎ�4�벌K|:��5�؇}l	y�M�8ȥ�K��A�Y���i�0����W���l/��C�S�-�md�� �%T���Nk��Q6���I$aW}�bS�`W������'�*�a�����~�I8|�����`�� �2M���Ym��A��������Y�1���Ӷ�y�$Tu~�ֻiG��}Z�CDVp�1v:��fhki��[�U�K��s�G��N�HW�|�0����O�BU�����O(��W��γ�uq�?4�7������I�.?��7�[m@X���3F`[2��"/���F#+l/����^��X�`*+�,�??*�np�Ť�z�n��kaY��v���xp�G�NȠ����~T.!���߳� ���kd̕����=��wmwu��#����nz\��s�ln\e��F�3?]<G��;a���Γ;��aK�к����(��(+���~f��,�k��i����H��A�E�Ym�Sq��,l�s�=�j�5����F���;��r��능&�p��t�'�f`�%vj"��D/�vo�Х�f>~)�F�{��%�SL:��nR�*���qf_�8\��E�Y��=	�x�x/5�j���(G�3FTdUS��*� O;���2�4ͦ����y��iҵ&n\����}�#��Dw$U�o����[2U�΢�d�x��`�1u+ii:,���i��U��Wo4N���4ټ��0$�6[N�i��z�`V���S��:9��Q����ʸ��$*_4�*�}A�Y��;���k�_��49ۯ��L�ভ|_��ή5��kd�|�u�?A�]\f4��msW���EVˠ]�Lq?��ӟ�J
LB�疜ݧ����7_�ow������n`\R���4~��"���*�����`����l�%�aw��y�eߣ��ꊬ�9A��a�?�����?d��2��b%��*�5յ��<�f)�Ag�I���:�~We�@R����N<�����O�5���>��[mq��e�� Z:�G�R_l��y�uf[6��W��44�N�|��Sb��uQ���9�j�x��o�f�C$Q��Z�E���(b�� ~p0Y�[-�R5��/Q#j\*���s�-�^��֌��GR{�MSW�}$�j��KJSQ*ZSR��2���$�0��y�⦫�Z�j��۳d�iɑ>r�v�ʍ�9�^�\pm��%�������m�ݝ�}�FC�y8$���7㘣��X8�?}�����`j"2�f�n$q����h`DG�0 �j�A��t$���Z܍v����|�������̼.�s��g �۲��{�j�B����|�X��Jm0��P�<�v\��;~u� 辣3�w�;�
U��y��`XI(��{(�b��R��cs��>���. c}AiE��B��3��Է��o��6>$��&Rd7eε�[ۿR����CN�=���=lCMYF\���K��A����N�T�9�-w�F@�����̮y���Ἵ��{�Za�"ۚU6���2�;�6����a�n������߾}c������BIJNu�0='��K%��^ڈ����4�c\f�Z�!~T��t6�������]O��1��Q7�7��b}b����m�zvE�S��h/���:�h���5fޖ�+m3�N୳RaQziZ��l�J�Gg<aU�u��3�M�E��ˠ�!�z���q���3�4���b*Ь��>�=����h�f��	S�������tkv�4Վ�(F뢌��c���V��!I�v�|��+d���C�zۀ(�p��
��Y�(��:�V���[Eɹ�l��۷R:s<s]�o�㡰F���W���*N~l����O���ʟ��O�@L>���ˏ���l`�`A��o��n����?�g�����EϋD��]a����
Z�L;��M��s�(�C�R��Sh�V)0���(~���/ߔ?���D:���h����{���(���ߔ���o��sP���kQ)l�C	��dӫ�ϛ�o�]���c���M���
t���t�sn-'�gu=f�h���u�x�	��nI��G�fF
g���7���s�d�!�Q���q����^ӂ}�ئ3I�!U@y��HH�l��|H;f�e�ػ�p�)x��T)U��f�]@h��?����`f�5�u.��gn�`�~�Sͦ���6�f�K\���^G�Pߑ�n�r-�,��i4��B�\j>A˙�]�p����D�6�R�����z/6�r�o�u��/�>fsq�}8v�\U��gk�F�s���vS���-���1%q���G����g�PZ�j�ӣ�AI�.���'�v7��{�ga�94:�����W�%N�`#�����YSk��=�s�zr�Ũk_\��g����l1m���!���}�����AV��-�w���5Ij�5��&D�2�D�>�N~ס��D���.����u�542ͷ��~�кW���9i�~UU�
R������{@#�p�<Z'K1Z=�S���q`�wׄͰ� 	�@j,c��Or��A�o�r���>�U��N�k�h|����NA��"-3ᚵ8\�[<\�k����i��?�jw?;�/���Y�|D�w�Kٙ�g���.�<�	����hk	��K���Lɹ�.�e}.�Pv������w� qY��9��!b���۞2>q� *`Ƚ��?>q+dZ(OQR�=#�����L���) �0�V��>���H-�L��C6�b��4���&�<��M-�Gɉ������,n�.�AM�k~N�[�eс��AX��[����o2�w*��9��?�;RX����?O��	b)Ӕs����e'�� �3d��|H�I`��k�g�����-cň�뵏�������� &��3"�>��poI@�uz>��ú9�Hfc\/�R�?s�\FzﴢSdǲى[|/��Z��[F�dv�G���Ͻm�;����0ѣ�Yj��mu��� ���=DV��'�`L�5F�b~��!����a��57��-��c��WcGZ��v#n�ц���>�J�v����+G�5D�r>����~�>�l��2�y�}���}>��|r;��x������`'��n�����J�+?�"��[0:_2�8*���Q�I�-1�_7��N�E>
����U��&f�T�*53
��k�������7qs�*`�8:�Ӕ^1�@8�v��Yw�������n���6ʼ(1��GX�`<��#�"����<�v�>�7]�쬊R��l/�9��Tqke��o��&���dS֎Ĉ����V�C�*&^�cB~_�����<6'��c�,�f2����gÑ�#Mq "���k���ꈘ5��7x��u��5�����x�H����%?dJ#^�
�l��^��T�&����_�����{���u�f�tJ"��֩��{>s������X3�p<�ն���?���M��_����_��"$ _�~7L�R̲��K���Q5z�&0�}ϳ�W>Л�V<���Q��a+��ƚ%$����c�ˠi��������ʌ��	�/3Re1+�޼���� �G��ʹ����6̋��.v�;�j�hv�=���"�q.����T���a�� ��Lʌ4������96�S��c�� �Q�]ˏł�q�&�Y��TY�"�2	�*�
��(�U�Ԅ��h�5	�;�<uu6��v@�{��ԫb�H�?c>k�����z>�OH����x!���ݼ��ز�7������M��7ހ|2�<�>L�d8`�Iӳ�a[fp挾X gAE摺��^Uz�!j����l^)�z]��؃�����u��WuQ�E���2'T��\/b�h�Y�9x�j��k�]r�^�kr��Ư�{�/5��q���g�ӻ��U����@�x�9����C�P��.�>kC���ӭhrp1#@uJ\�@z�h�c��Fh�K��dУ��׻�\/��a�P�o���⢿��s��L�z1L?H�'��4{�*)��޶�x`6�F�Hؐ��鴉�����S#�d˒[W��[X�c�Cr�$\��D�Ϝ#���c�{��i�eP[�k�4�w��@I��9ի�X�v1�0�n G(�r���=2D�6�������V�ϑƠSMW��%57�i�m�dzd|fp)ׅ�u%'����R���uU��S#�:4T�D���*�#�3����8�H��UgF&Xg��������c�?���'H�x�N�!n���U<KOVY�o�W�a\4ۆe���U�].׫pOR|����b��\��p����{pqh�p�C {������!�G+�8�\�����	׽�I�}b䰔�������xH�+9�k�6d�������Ջ�YTC��ۆ�!��B�iRv�5Yj������E��aLڛ���p���1�{�� �8pE�s/m��5����vkN��������>�����q9�_�D6��&��N�P�1���d�HKwu�o�2\��qS���#x����x���!�`��"���Pv��WY�J��	׹����Ό3rUI���c/����T��@P�ˋ�P/��faA�`���j���m�� x�B�x�)�R`�y^�~��xKIƁt'�ؼ���y��k{Ǜ��CCg[�8ݖ�,������*�%���F*-S��%䶵�~�BƗ�)��yJ�Gݫ�cjZ�.�bUX��MNE��h7,hxh���_n�Sq��a=��h�l�"ή�yt�ٽ�(�u��b�&�b�K6��<�zцFӇ�R�����tֺ�ڧ�h�G�]]3�N���������}po�`���yr�EE��/_��τu�Aՙ���� 62pV%?��	%�xI{i�b_�ps��=m�X�`����=py�.�Dvf"�����6�����/����eоi&�4�\�'���Ɩy����e������3����	��5}߹��1N*�>6OGM�SJi0�ύ�0��`��� �<ƇbMS\�7=�O��9�0v+1�ikF��s�E��zŠ�Ec��=;�X��	-������ ?Ԓ���I�7�z�ʉ��q;<7��%�I姽��-E
�wY6b�b�yءf�
���`w���6˟�N�:Q��DQ'�BS�r~\�Ai�l�`��n�2�����x���(��7:�f��c����M�<�*����%��Q|�R�c����_���B}����דw�{A:3m��A|`@F�N�䇃n�>��1H�gF�r4�G/au_�Բ���/�jw �~�P�S3�5},�u�������׿��|���X��	��ٔ�t���HF�'.���ze2�%�(�/3R�[
߻�@����HnY5�2���C��A��l�ob܋���&S�Yr�Z��$YWnd�ܥnK��r�򔖳���]�%/ ��8���R'�}���Ɖ���tKzo��Β����	ߍ),~\<S&�Md�5��� ��]��<[l�^�L�,���Y�q�A�LA�,NLt�-�RD���'��(Oo�i=Yt�����y:�~��͔]Y4����"2�٢ȝU�x����&�p_.�Qt�dA�ZYW�/ǉ��H��\6�]�:����R� ΌG�����+!&�ڳSnT$@�>ꐆ��fN���]����3~��~��c�D��l$�:b�u���ڋ\0���P����$$�~�s����u�[�Ã�t��cjMe5��NN�U�'��C��	SL�'�\Ϣ�~�V:�Y���e�P�Np�1�L\�בW�`j_�����}�)?+�y]��O�Z^C��)X���{q��ÿ)������柚s�$�7Wүb����5���V�p� ������-M�����B	1��(iwj�Ĭx �E��P���Q�a��A�9�j1�Sjs������s_4������I����5�<r,��Vc�BΚ��$�u�$���f�;³��ÐT%c1x��y�h<ܱ逮7ԗ��Oo^��:>��Z,�C�J���6\[u�=E�Qؖ6�Ӗ�m�&�Il�:�s.�96�/�e|>l�!���,�}��=��0⼇��3$�n�]nJc�$�ӛi�F����VOs�^�+�s�R6�F|t�B؍;�2�D^�Ce����Lա�qNe�����s�9sPe���k��]	>�+ye����ӳ��!�;��1�.n�ik7=�C����G��x'���h/�)8�Ac����dp�*2য়.珧��Y�߶�N�)�,���;�bϵ:��χL�)D¹�#a!c�A�92{�m�������Gb��Uk�d��\�z��K�����(K6�;dl���."U|�� ��$����"� 	0wZG��q�x*���ޚ��Sȟ���� p���y,�bj���D�M5{�#d(ۄ?_j�M�
������8D�)�	��Z�uɓ�vΚ7���Oi������	�P`?Y�^M�F��c��90�[���w�@����.|d#[�.�IS�~Φ����!5��%q	�,'W��} �,)��w�����z���aga[�0�k�M��Q눙]!�bf��Vk�#o+K�x�l�V�����x���k	��-�D[B�>FDe4hoyg����j�1hw�����_
XL���&�r\{�In-�"�!T��"��0�v$#���31 ��m����Op>���uܮpT\L~q]�@�^s?[�1��V��+)iN�8\��9��q��Q��ىM��H�>��<"S��gs�j䶬o)PM ����T��h��oڈ��@�]i<�-/�	�t�����b6N�FT�i�F���b��XHn�8����M%nS���T�4k.S."��^�:PR�R��=�t�E*;�e�5�1��TWͲ۱F3�������('tP�c���&H���:gVϑ�����P����J�d�v'}G|h��چF�/(����U�6�����}��D�*1v9���s��T�5&��q�uu��~��q���k��#�3q�W~f�́���\�����
�@���8 �ɓ��hU�:�g�3Y.ѴقFW�y�)���:��U���d#x���eR��m�p�ʵt�#��ԔM�k��AC*�
�:�!�S~�W���y��_��^���M���+I����� �/�"�$*["^z��n e��gm��Ҿ��Ϧ�Ң~sQ�/�:�>��Y~�YR���^+��E��UcVervus�.��u~�⢴nm�_�lWo�^��|C��Fv���N"��̓���XMP�ix*ܭ��}�Lc�)d�4��F����=�>��"������^���Y��8��:U�n�[0=�̒&�"	|ɃA3,������UK��=�l\�9߫�N�5k>��}x��Wu����ὤn�����pΒ��}蚆� %��MV���Q�wQ.>QzM��J�MG� e*�?�ZQ������'N�����E	U�2J���k��6�~�M2�,Bَ���Ʃ��'���J|��Zs|{������ ۬ؖǪe-t�φ�����5�8C��c��E&Y�-�Oۑi�K����F�X�������3s|\B���]|��F��h eW�p�<��d��їA�������	��<�M�?�,2��{FrfX�F<귈�̕�^@�q��Y�mDy�:0<��C'p�|c���=[O��t��l��a׍�PY|@�E�2D��Q;���̞����ݾ�����	��ĸ��V���\<��DX�����WF���CbL"�� 8DP��
[��C-%e�]���/'
��cv�c�|�%�z�y̯�b�����1M�)a3D����7qt�yk���rY{�U�g��[�xz�p�,�}������Ɵ-L��F)1궲������Y4� {,{9�j&��[�E�.�Ӓ|H��}ec��V!S���ύ��/���Q���t@n4L�Fa�6�+���.��;}�x��ľ��J�!����'wy8:!۫R!���ʪ�=UC�Ӈmu�+֭�5U�v���� N�rH?7*�2v�-����s���H+ �m�ܴs3D�y�?J��WY�X�0�N)�!Ԓ9�o)@���!�4F�IBO��Q����r�����o���D������-6���P��`�\��͡�T���f��U>������-���)���A��'r��
28� ��d���b�c{Ƭ����
"C�kFF
ag�{e����� �U�$��츒括.��J�l�a��C��e%&���`s�T1��}_K�c�%���/�����q*�ݷq�m��9��������f���v�x�X��.�F��g�qO��q]^�E8�D�7lF����e�`0��5�7݉-A��Լ�O�a�T*��5��3�[麪�w�l��֚�ޯ�[p�B�O�&䚛ܒ}H�p����З����������@s';�g"k�Dۛ�nJ{g��3�8�G��KV��ңu�)��������z��?Ta�'�ط��s��6]K�qm�>g����oJ���oI�QY��T�r~���v�$�|ǡ��v�ÅGm>J�yN� �i�,I������Z:S �Lb�J�/�~Q[����8bY�+��tC]������g9�,yr"�5D�R{�I����0��:��ZzF��j��R�,�����4�U��}_;��=�Y��kEO"��)�mQ���)�{7D��)���N����]t�,����ce�j�F��>�=3@l�*�a^�ks�" K��n�Dè����e�7�!9�Kfz� g�/>��s[g�q�.��XJg5����R��qW%��vl�Z�x]�̓|����K�a�������Ɔ�xcS�$�|H�_r �<�-�gc���=V5*�	���!3	���Ȁc0�'�#����m+u-v�5G4՗�}�k>i$�=�~n�(����Cl,7|P��eɪ��oB�ON �ጴ	���9�t��������� ڈ=�-dp�7]/��������ù�1J#|��c�V��'��7��� �l�̅��}�	�߉��12�h߸3v��t�92Hi��('G50��Is�9����m�2#�gƵ����oLq]*(��Ye��}����e�9v`�G3�)�l����:��&G�QHƙ�*e���=%��K)���-t�03�13Ho��da��%����pM�?1x^�3p��(T���gW�4��M��5 RY�E�Bf��[?�X.���0��X�p��w��sZ#�����
���LєS���,�?Nὢ��ݕ�Bcj!�]]����c�'MM���5N�=;T>x�f��Te��5���,���I�в��&���o�q�s,�=�^jh�Z{%�U��^�jk�duT���h�L8���up���]M��o�z���YN��-�Q~"��.�f֐+�������H����G�0�>�I�0�g�h��72�*GDY�y$��{*��"�؜#��>���ByV�e���p�a����F�<熻���O��b��t��L��]L¨�Z� ��� ~�%<���g�Gb�����ӹڞ\�ªkӍ�,Kynbb�?�u��'���_~��	6��6N���Gl�e��2/y�[W`=
ЗسG��W�?�9��ӧ��#7^Ã55&�ƒ��%Y�ED���(��XC��gMU6C)]67|��<9~���&�����ǽgY�^�q�<��	�i�q�	�)�����~����L��mu�wǼ��*w%=�^�y�?T�g�+E~P�\^	��aa��D:S`�#S��Y_7�P�y��0g��HMs��oh��� ���;9���y#��6zd�����4�O�An���2Qn�kvν���n�".��C���u��"+M��gzT��/՟��8����݅�6&S�2s@#�(<Y���3�����(���(�n2Ŋ��F�X'YڇŔiJ6��(�z7%��P�萴|�k,�-���e��w�WQM�=s(�p��>��,��yROqY�Q���;�qb�`|nd-ԫ �x�����\Ж��Wx����ʴ���Y��0=�
*�ƴ�V�������Bة��/���$�hA@�P���z/)I�R}���U��q�R�Y�)j�4��Xi�q�|�%zW�lx�1���r���^��5Gfs3r�C�r,	{�o���`��[6��:����:�w;�� ��VV{�ά]<�:����k�t֧-�yg���X�3 �]�L��(P���-�]Gd]�$Ωr��J4��IB�!��L�yg4K(Y.k��6�m_��o/,�S���Wc��W-���������}��Mv�q�(�z*�co<��'9D�3�c7��I�����y����J�-�S᤬��JH�WLQڅ1���9q��YĻ�*�j�&r���^z�~]�7U#����9����6�3\�E��Ӊ�.<Hc����?������}Pq �Cٓ	��ϧoy�uх=�X�21by,���u�:S��_Z2fb1;�ߛ�o�LS�(�qݮ?�� �˝�Z;�suq�l����0�29�<5͆�b���%u��lv�3�w!J���{/�����1�Wxϯ�Y���L���h\��y��e)�!���HJ���|�
7m�'}o�2r��b3P��T�K:��g�Z���2 ���C���� ��Z]��0���1�Y=�(����a@�D�'Lr+���FQ@z�S�G}����kPX��G�����!�m�b�'�]m�l���)Ɖ�\nIퟎk�: �Y��'V���}�Oi頛��X�gP�f�N¡Y ��]0�2Ͳ��?,Ynn�tь��}����{宒�����%�{qR�B}��K*�������^�cnZ�eC���%���T�]�M���#0�lg�Z�vIA`��xo_~�e�0���N*N�Y��?�7bӂ���Oc`��J`�y̿K����~����'�IԀ-��t����:={.������17�`_�$�>��ǟ" >Kَx�n������k�Uy��?�xt�*���!9��
�	��4Js�F�Ǩ-U�������4��-��C�_Y�^I��c���!8�C��:�&_�<p;4������x���g鿺*�[���Ycd6�\�lH��ĩ�nq8���&��ϵR܍
�����yω:*[���!�c~,t%�[}��H�2��Q�0�b����Z�F�ߊqMm��LӞ�6��F�)c�ZR�Y�z���D��u�î�}��cbòwMѸsH�g�(nx��=}\NV��K^���u���8��r�#Tm�x�f�$u�era��n(x}� �)�P�FwU�'7��j���Np���^�{[�WK�d�����Z����W�aPf�&�gz�����im�1�`ab�<>�iDpD0@���ߗ�[��y���L�#������� �,L<�{*���Ȫ�EF�k��As�������]%�_�?Y�ib4қo���Ȧ�}I��00�ޔ(��̄2��G`�_ƿ�I����w�[%p����#�`Z@�@%�ydb9�R�LL�����ԫ��w?���ى�@Jؒs�\��3-:����H֚E+���W��b�V��X�p��D�3�C�Q���{��o �~/3;KL���
�l�AL?���o}�E�]����P�4��G`[~���S�%��/W�;�llkb�M m��~���ڷ���UFu���l�f���=�ۧ�7	���~(
h�JիK�ε�]g��F8ES%]W,����7?w�i�k�N��IO
Q������
�.���0�+�k���"�# �Fb�Qd�<E�,Y����6�_��_�d�2M��,q͆A��Y0ÚЀ�yv�Ǫ]���cp:�����l��������%w�,�������lrR�9d�y�ƋKq$^��ƃ���y���m�a��B����]�kn�p�a�Ԁr[�����!�k�*���W6�D>/��z���U���ۉB���<LT��@v���J[���w��c���<�F��2�d��y'��n�=5�]a.k)i)~�X�i�W�L�;�����e؎�"�1"^������X��QP&�k ��U��Ϝ$�l[l\V/{%Ss��z%�^����ے�s�_�&�&�?����x��ET��FvW�����I�8�A*N)�*a���$�
���Y���8cf-o�e�U���&��Ӣ~Z2kI�ځ#�E�I�a�f ]Ǫ��Eq���,\���%x�ʥ��l�V�:�q2�ê��O�ɱ��<�-��������i�x�z5���J�4�s��Vx�;ǊF�!��
,���>�MOʯ�1=(��`zT��mF��)w瓟��u�\~�J���C�R�$�KIj�%)l�	t��Nc�2�R2���D�id����vݤ���?��+'��Cx�X{b�kH�R��u�ܰ������N�a�2�����U�U�,���5�~�S�'�oШ��e�r̖��b~tW�(�"�N}���(���d�7��� �����O�̴���V.4��N�.������:Nlyr�h�a�C���'ao��5�ԥ���U7�ڊǐ&/_�s'�&W+#m�������T�{�)���C�������]j��p�H�9�t<��XMI?�sR3f�@6�l]�8��"��HW�|��]ROܶb�G�Y]Q��J�sjA���p���JN_Df	|�
>ۿ���.m4������qXH��P����b"�ڡP�|V�aHVC\c�xS��Ј(�l��)J���#7���?��C�*fe�U�k�@jb��-wh�D ��@j��e�9��tv���s��#��p��>>ׇ����)߇�}��G���S�I��]׶��Yk1Gr�~�N^�I�#]]�!��Q]�bQ�s8���U8C���{��>�]eM^���8���"7�AR��.p�<�`����B�<̍}�5ͺ.�d�j��E�����'���YҘ��zb�M��X�
����_�V�ŔKqԳ��8��\������ό+������~���?�w��R,�ٰK�5��7�g����t�M�w�./�o~�'mY���8K\�d���
�z*�:�bP��'��s-��U^X��K#b�`�ճ���t[��M�x1>�fO�l1��i�`������/)A�yʉ�T��1����u�����i[����*/����Z#�봮O�a"����gH�w)u�5�x*�eN�HӸ������8��pw?��t(��UA��L�����d�k ����j�����lӿPj���ee3�
\2h1O	?P��,C�|'w��M��J��R�#Pm��t~.�xnܿ9h�8}��q�)�m��]�K�������f���xm47'N{��!���jXԱXWNn`�k��b�e��FW��:�˲}��&ovi�*��U��&�sQ*,牧ć�Q�ha�o��&���	�D��7Yc�,��tlD�fF������S�j+R�jE��-$S=TsĹ����Z��"46��Z����)�����k����0dh����h�ΐ�)V�oEO�Cc/�t���j�y��]r4:bzC[����TR�ԇ���dg�A��UV�t&R��(a�{��̲ٛ��>{�*�ߋ�*��Z��/���E}�Nr<���m�X�&q �(��:��X�Sx��D����쬥�\�ɽ\D�fFG��1�8k'6�>��cs���(0jX	>�! ��ĕ;�}~�T���C���}X�D�T�q��@�A��ns������|���^�/�4PP���Ú�&2<�ږu�W`���^Z�.?�f�������� ��]��-�rW�g`�θ���w%2�k>h��2�a�`�l$����`��qC��2Q1E�WF{e_^}�*��u88���Xo�{۔"�m.)u��)YJt8�v'N�9лX���������Y�Mwc��}��X쇏O��e�y�Uq��t$9��o;���EE����Eж)`4���ܳt#��%�y��Z!���5WAN�v�xe3��E�R���hU��ߥJ�nO�V����Y�M5pƢ�^��1�c��ʢ�()�HǓ��5��>��H��Y:��s�~z��3(���(D�Z��}��q�����ݗ[�$k�!:�8�&�`U���LW���9�����e�Oz^��k<�O�q�ef��S�!ba��9i������ԫ�;��4��x-v�<���&��@:���� ��r��ޗ������z�5��$�'���0#E�����/�����:�0!<n�퍦�������qz�e�8&lT{5�h#�����5�Lt�T�������Q�ӝ���CE�A�\`po�P�!��Ə��!-L�`-��t�ꉍ>�E8>ዧ8���D����7��OMD0މ������`X�`������ډ�=%o�R3�z����[�j#Jr�Hh@�����`^V1�ԅ��Q"q��`�m�߷���x�1����}�}��۷��{X픊sR��^m�d�е���O�ʙ-5u��R�\���l|�^�oRӵ�V쵴��~�|V�	�V+�꥾�71���')�#�a�C��Ol�ڢ�7B��ISLL�O�Q������� ��)�mh����G� 5  ��IDAT	^Sd���F�M �Y\He��6��I���-'��1!�R_�\��S<���R�r��ט��A��+NHϥ�4�Eg�*�k|����:�4G�e�1��L�ϊlP�AI'�5,�JB��M9F�́�q;�t`=wqm�����z����- �������=J=dJ���C�,6���H�(�	�\Dy+HCa�0�L�x����d�>3��f߱y�M���-y����]/���`p
=�s_���~��.�i����G��Vb�Zi� ��1��A$24��b+�*����?��m|a�ʥ)����Ǟ��ڴi ���E�A\'��Q;a����i�m>�����ѕ?s ��ڼ�ɫ�Hp	2��I*\?��KE]��V_��?Pa�aKt���m��Sy����*Û�<j�ǌ��
��ګ�޿��s�>m^��m���x�-�F�����s6��:�Ns�0�����e_GILi����H�h��_�[�?����@c�I�-ʗO����٢	R;]#��/��fJ����^�	���+�G�+�%�Q:~�q�[��ĉ����xi_5%�6���Y�N�˙����]], �;��o��6��(�K�i�>	��2��D�x���d:F&�H�Sb��-��2���TEo�p>q�N�!1Y�g�)�14������0�l�t���(o8�8M�j�p��%��.�|�F��Lq�LL>S���X��|��>%��<k��Xօ����I��E;��ê`@����.��9����E��^�����DzT6$����t����Lb$wj�-�Mۢ��++%�J�/����d�;a/r%e��^�mr�l��������L8��E��F��:����`HЩD�d�5G[����T���qLq��p/=�E��������q�Gx|ٱ�oŴ��r)^�m�/p�_�ڋ)p�P�jl��%��R�� ��R8���j�Zd�7H`w�����JH<<_k=Ã�΍{����iG��Y�����h����$,u��u�����\Q>7�`���HM�5�M��N/��>�M�����:��3�[���>?���C�IZrz��0率Es����.ͨecu��Hl�����3�{�,]zL��K�MJ�kSw���a���CvAd�;
N�Y#K�i��r�DO� �l����(--Z_����q��*��~�1X�+�e���HOaZؘ��o�5Ґ ��4�C&�;I_A::&�XL<q��<�GE���U��k�O�W/�
kV�R�$�"!���k��<o���"XU��Ś����R�=��,����T<8�Pa%
O�J����޽$)/a.�XJ#x�^�l��\�X��ٶo^w��_DÊp��g0]�;�M�+���)s�Y\����*�A���BV$jtDC�H�	�(j �͜���%j'n��頎	s���dZ⦂f�O�)G�tc��}N?�A����^�/ys���7���Ep��7��[sY�=�F�Z��s�|�m����])=�s'g�5pa����g�">#-"�7��%�\��>��=��J6Ѱ�������'�"�}���کn)[��4�]Uq���E�-6c�ٿ&��A��C6(Hў�H1��C�!��agmh
2s�u{ߏ�����A,���S'`Vއg���]��G ��gk�Ȇ�t�v�fmd���[�9 lf�ގ�֬�Q��!�9#��l�K�ci����&&��� u��Ab�(zē�y�C/}�k� �~�,~)�St�������`Gׇ��q�����'T�W������ �F6��t�i��=s�ڪ�NZ���՚0v�lB�mH}��'�O�P_k��]y��S0AO¤�v�M��RC�y��.��$�������u�q�`S��g�X5I�'x>W�x<�Si|��'[sAr���#�*�ʖC�Z�f��cs<.�����)�!]Nu���|O}�m�W9���l��z���7ӕܵ�'�j�.�7a�K(�LoGs/�0"(7��"3��1_#��m��,�ρ�⑬�ރU�>(AӮ�ǋ��a�Z�k=���2�t�j��@<���m1	���;&�]y���XZ�YC"� �*{@�k�k�3�7�x�q�f�*�f�U=]VD�F��	�??���[������`K��霊����ݼa����7T�f]r�ɴQ�Y�` W1���9j�H\����0�ڳ�y�V�Z�L����{!����57�+�����ӛG�A\�_�(�������`j�%P-�'���aS�!�o����]k�� ެ\ܖֳ琝��k�g!t{�w�qp�eR-s��|J��6��u��J@��sww���Tw��pUL����.9��r��4������ڭ�"���V!���i������U�RZX���р��m��K�MO����,���SZ������&��d�¡<��kX�����	6V��8^/wJ��Q���q�M�_�
��ŋ�j%=�"���)pT��=]Yj_��C�"�F�GRK��Jd��ķty�gt�CZ9Q��9�����
g�]���˿j��[s_}��$�������Q��#@]��7�HI�qow����5�X�`�$���I�������:S.�/_�G�ş�n�'ۉ~[B����p���?7��.4#qmrXik�y�����&`:1��m~���u�p���6�������]�J6wv��w*]�A�oE��+	���fVZ�fv��T`b�B�o�<�Z�-��ɥQ�m��>�ΰ7	��^gެ�����luLӺ���%��?�`�T�J)�����i��*л�,(��+Ŗ)z�u�nndZ��l�V��Y';a����(Hm<3�~��g����{�oF0ؾ��tv
��X�ȱ��'��F~�Lai��p�D_+(�
��yӣVm���X+�<��G�[յ�'_ه]`�=7`��t	 ��p�D��*Y�'�a�N �7�0Q	����I��R15�G7�܀�RW�1�0h�cА�S)��s�YbIݣy�k�uy|k>?���T�5��1ڄQ�
�#K��XFYu�9���$��ꃲq7&��ڍ٠�m��1�/���t�F��ʪ�z����xc�x%�5���ᜐ�ݘ\����9���r��$�ȣ������TF��v�l�V1.�,���*94��te�74���J��������^��s9w��t����W'��A����z>��6�|7�P��(3����P;��1o.��8�!��Y���^�*�d6���N�}yj%���BG@�ٷ��	������m
������'q��]��sQ�Y[ܼ2���`�eł�<[a��swS��
���*9b{w(�Hw��>�
R�}�;�g�w�}�J�v�p�9⹦���	�u9�ɘT������-uD��U\�yݾ\�.iHǁ?Uy|����#�R�.�a8�IUת�׈�,�Y�S�@�k-��jXثѺ�yz�3���Um��;��!�?w��w4�f��yNۏǇ���|E��ӾIF.�}SԦSt
]�=�}�;Á.F����)!�Q�~c��X^{�S(�km}�H^�y=i DM����H}M��q�`ɉ
N��~�m$�amgt^� �K�D��P I���-Z+��Sץ[�������Q�������/�pnbg�}�6��QJ)!�i� e�xMa��d5�>_dB�[V��U'���(KZ[��V���f�Vu�yqm��]䎚���Ȓ,�#��]�{M�8�a�3Ŷ�m��n��=qPA� ��"� ƍ�[Ux�)[)J�
����c1gXI�Wf��[�y�"�^�o�A�
������u��׊�z�; B3����%��/[Y��?��C�x ��d���*rb?����'���A�G�B2�p_��[ ,�5�F������Wb�%�X�b$���Q� ��b7��z?d�Up�J�{W�d���O�R�/\W�w0�u�8�� {`�>�i���,?��Lj�]��D�l
[ʜ��I;د`>��Vގ�_���н�#/��}:�q ۵�������0P<)�}&a�!�rܒ��>�~�]~�q���?,E��.�;��D�"u��0�e�*Y9I���p��r4������>�e�M�]�6�fl-c��_���&Z�hJx>w�)�f�)𬡿��A�`Q�+�j0���Z�Ɲ��͙�婸�'�ɹ}a�n����9u*�i6����N����������st�n�.�\�x�x�j+k+[XN��!i&�5�:ϵ̟ĵ���7uU0^8���ڭ�nO �}����6�o˻�]V�p�8Y�J�Rljt�@�Q9�|���-0�\���T�m���O?FF���p���^X������s����&!�B�P��k�D_����O�7�f����b�Ŝ�MHn���� z>�����JC�mnl�Xo��s����b�n�1i��
�P��S�Ӌt
�')�6��a�Ǜ�M��%�?����㚮N8@�y��6�Sd��>~J?,�����
E~�ݧV/1 �/QN��Z��}���~/���EAu�W�����'�8FK��,J!~�z��.�Տ�fS�W.&�T)�hjO�����
�u��Y�ˌ�-z��Xe�~>-*�FM}36��{��fZ].�1��>yr��k�	,��E �\Hӫ��݈����>ˎᄾ�&�z`O�4uEϘ�Խ�<�&�sc�,23�̀l6Tp�`E�<��]������M���{�m��u?cwK;����i���	QU��x�)�����u�^bSQ5�$��.&@�x�{��n�O�yx��<d_#��o��~��~_|~���!s�����M�Ʉv*^�I��*��ľ�����35��b`|�5���o��\�&͊����@�,>!���n<�����3���#&{`���2U\˷o����TXz��Y�k��ÞSZ��m��)(;8�4�瓦Ӱ��7XcȲP�L0G���n�0�lf�����a��E���D6y2�������a�,�|Tew�:�Q��@1����i�K�®�ʎ�h$>߳rz�5q�fAO�%��z̓��.5s/��И�\�jm�����6��ܟn1uM�%|���������GПn"q)�/��V�hF-�B�tSd�^*��x� �T_{=�ʟu���S�x�{\,f�]_��3���m��e�,_���#�)�3�":�/�RO`�E�!'�,K	7�,J[�ܐ����@�B� �cO�)��Ź}R�P:���L1Ϣ�U�I�ua�g%ot��a�w?�9����/[v�6:��;'���ӗ��Fr����*���ڟ5]��<1����ǂ�츯JE��K	6&�N�n?1����{���"5�"j�7iR��]4��"7C������H�Z����
ig�O���z�������J̞�7d7<��������'�E;�����[~$��]6ȴO;7<�z�h(�ؠ^���?�i��a=��0��-��J�.�����"\9'��p=�	`�׊UcPв��ġ'!��f1z%�o!�u�>�F���ե�]���3��&�2��^Mm6uk�d닧k���,j2�f_�/��N�d*nTi�ɦ��=e��P'�i8�+�����^䦌1C�����@
��G
Q�Q�#nW-̢�g?����\2��-���3&7�,eJަ'JL�vy�bR�|�����uRC�J�r����fѥH'����)'��^p�~�2Od����lY�w�G�hm�^b6����"�� ��π����ӖA��e���a���6�����%�^)��Xcl&|6yQ�f����s�����ރ����n��.�q{����fc�iCB<��u�:Y�<s��lBxw���	�p�wm3��f�+�%�5�O�/xN��}��`-,U����E�pW�x��	����x/�X�����~��Q�@�b�7ؠ5�t��r�l.}�w��Ĕv({�[���������l����{�j^>�]���R9n�#�{�`��U!�]�MתlFiF�����|�Yέ��YX]���/�ￌz7�$�B�ڶ�?۵ߩ[�ܯϩ�khG�T'Tz���Hh�p�[E��m��O[��_`$
�]g�P�]��R�Z+	7��,w9�rUV�At���q�o��J1��e̐Ap�q����n��(����,�8���U��Ͳ�16�Z���lnL���\No��0�B�m��+c`˜��i'R`���}���{L�(K
`{���ͷ�_~�;��?�xf&�X/vJB������@*�
oW(�qw�4틦�0�P�W�!h��-d�߼�ύ��Γ���Aim�*���`�]�>�uұ,Z�/��U��Ն�>x
�*a���*�����?�@���x���Qe)uvEÁ���92�����w���=����tR�.�sL���������Il���	���[��C"5w�믾�����Qڢ#�E��V3�[O�S܀q�|�z��ob?5j�^?��C�,�	;�׋�dM79բ3v�2Z����ٻ܍m��_���z�W�F��qõ�t}Ѯ*�	�E��Q�^2W������c���0�2f�j��^��K�ِ.�J/�z����Ew�d`���U�X�OR����.,8��l����	��5��No_�,d,��"��̪H�#J��(�հ�8�7�F;�-���U5��q�<Q�x��
6�n��)��.T�a_�^���?�#.�k=����o[����_q���[��t�9@�~�6۫mc�wU�8J��:�����|�!����|�Y`��j1���M�nZ4�ο�Md�x��<�(O�E
��]b6��.�A�{��ꫯc#c�;$��8�������zl���b]�?�R��_�5��-����)2((ɿ�2�����L�5��k��w����ۧ�I��z�a��!A��t.�8(��:2q��ή��)��&�(Q�q{��"[�5�z�H�N���]V�=�P[l���5�kb�j��"�w����aOS!��OмA�mQ��̙,�E�=hdMw��XsQÉ@��v_�i4��Ϧ{wP_ƾ��* Lsf�)р�����Í闻�]ߗJ���ӑu�j�n`���;a%�P=qH�K��dR�-�N�xl��a|-R��_E@�3e�3�V�1%�ジ�����X��C?gwݣ��i�baFᙶ�-�#���U\�*(;7�c`�w�T�!efMz�$�<Oq_�B�e �Q�W<�Ο߿���6���xV����#2����|z��#}��J���x~Fऊ=՗Ne�5B@C)�k�$K
NBu�^���Np��k���t)_lb�Mɹ��E�W�/)}]�d����j���(��c��d�i3�h`^N�\����|���=l)+�g�HMX�S#��z��^���}�h'��vYk��pN�`#�pܫx�ۡx�2ЀKcWf���7����L���}a��C��ￋ���UQ/��k	�z��7�07=!���}� S�I�S;�p��Ly����VIڟ�����[vѱ)�����d�	r�L0���6��4�Y��_wg���x�~����� ̆JrY^T!h������R
���b3��e���Sj=�\\D�GK��b�=E	q���~'�5�p���<�<�1�Z6A�@���Ӯx��oP�N� �62Y({��נx3N�sNjy.�ﰫ�D��u�A�Rg��w,/m(f���l&��>||��ݲ#v�?
���|M�"6��A"���2X¿�Cv��{U��&.8O[6����p|f`��`�~ձ����3�ٳ�:�p�m�L�@�����Dbp.UbF�NtW;ĤwA��m��u]��X�r��"h6@���B�Tk�A�*=�):�o�w[�AV�a5|�; ��Hm�v���h���!��������Y�a�^�D[��{�0̼�z�a5���D Fј�� "@聆�Y�^q�~��|��)��Coù)��A�l�3���>M�q�p݂
6ŶP�>�R������ �� .k5����1�`۶SA-�?���1�k	��OR���w*N�����ڑ=g��X*���P8����ӣ�蚓�4��r�j_.RohX���)��Q�`�6
6��\(�_F���������2#e&cJw��)�X=i��2�cv�俍��",��C]�mV;
|.�aR�n�˭�3ϝ�Jc=}p|.��i�;DV�L	e��ۿ���r	e��X���:�����E��.=�)�Q���D߲�k|�����T��LB@�1�Y]PT)����<����	��.
�,	^��$|��7�o����r��n/�Fb�'��N��|X�zT�x�*�N��wB�8�8W�Ԁ�&����������m�\�k�(%��c��~�z��m������` %���5<���c`�j[�d�����x0�0�n�s��8 0O�*�q=�1�yA	��{{>H㿷l4���U���N��%F}��p��Ʒd`�վ���E�9�l��lR���RӕU{$x��$N������Ju���}��|[/M��30�����f���㒳WL�#��X]��Km�1T���rYʈ1��:ҕ�������Uc�&"⢮jRQ�T7W���Y�F�j|`q,���]0��sGv2HA���k&Y)ksP�e�.���]�T[�Uԑn�%S���?���ߛ/�����+���ۻ��R�%�_\[�v�8�vsF06Nk�P��+�2p����r�2�̗@G�ཱhd>�n��K��Zm-'��)�WB�����<<�.�ؠ47zh?lPuy�өD�Ͷ(+�	{A������,�ל�_T��`����١�I��ڮ�!�V��t�Yz,_H�k� ���w�Q�f��z�_"��p�9{�MơK�cP���؜��2�iIkp��i���h"p��X�n�����iX�s6ׅ+��x��:����g�J+�e͉HŢ�T�\�2���jx�Zm6��M�|���"֟��V�cMN�^�-U�,��q�q��L���h�{��j�sN7���ܔ(�/�8�x�g��6���5&ya�nj���|�%�{u��n��tΟ娤����[L���@5�벋K"8a��I�]�����#����e�k!X� �ed��6=�6��^vc�F%����5t�����K���6�,͝��]�cC�(+ab�U"�bN�@}ZUle������'2�!�����\� /��&���(�l�5��k�X�/���Ы�#�f,l�����#1�=�{O>dۋ��Ş�C���E�2r���Z��l�H�S\h�E��}j�_�f�E���6ꟺ�]��X�rL���^:���Ս�OŴY�ly�B�K*�]�`���S���љ��D6�6�qJ�>�*qx�(�r�حu6������r�솲��T��p�(�X�nn_�٬nGu=�W���5K����7׼��������u�n:B�{X��xϨC8!� '*� �`���A�V�0��ӧ���Y�2�_0���s�i��(b��Aa�=�씁Ya!<iƅ�7�K~cCbZQ���4��Ih����7ю$9�E#3k�{O���CJ��wλ��9W�<Q��z�7 ������<�0=$������%3�����L߱ #�>�w<�B�S����d����NDK�ÀGv�d7ު[��(dX��P�Xhr �C&����$�c�Nоk����W4�۳��谡�� 8��9\O��ht�6�X �J���C�KN�PN�<�1�.w돇��b��ذZ���8Y~�����EƎO
�5�3��Ø���|�1����|��؉����z��vbw����T��	��:��DUB]Tf[��K����f�����iy�h�����8hl�eiOtV��!�@�=u�sm��$�q`R�gO�ym�j
+�C5�;�
�n����3��r6�v#�6G�T�fuФ��&�⋲Y7�fą{2nv��MU(n�!"WY�?�L1��ǛH��@����`�����E|Avϐ�?�P�?j�����.8k�M���P_ҁt�>̱h�z䍴C���a��
]vR�A�:���o��?|ҬnH��[*��6�b��R/�es��ڶ�F �ȭ�f�{s8~҄�j'�M�x^Q�Dt2�Gd�UB�R�5\�)����ԛ�k��Y�����?��%9�QHZ4�����p8V)V�>�+�oKd�;�.tW��ͫ�Ff�(�� �h8İ16y�1��㬌%~�y�M"d&G���Ģ�<�#��>��͇���q�{T��CJ�J��ðո�a]���\B�*��!(2��Ngf�񾩠u,��H���^M�C[���A��Fad�de��۞����o�C.|b���v��Mu�C2�Rk`g�j�w8�=��ڧmTV1ew)w9���5�N���:^3���Q����Qb�$�A��7�6�.5#�Vq��gU��=j�ڕχ�_��o���Ɏ�J�Ƙ4�|=n$2P�a�	!z�Vb��4Y���XbQ���=�8�R�l.*$��.F��领������������&ZB_�4��l՚b�����gYJXޫ�l-�R�c�AM'c���u��5��>�B!0�y�V����:lrlp�����X]<������R��G�td馋��X4��f��(.���#��`"F^�)���]?�Sp'�/���u��j̹���M��eנZ��w4Sb�(���QNs�F�
���fW����F�7ŭ-s(K���������c�gk ��g-�{�/r/�(9�;k]��6}/qg��r���%9���X�?��l�c\ҜKVg⃚�2�\�ݸ	Z��%�h��kZ��'�s�	�j<z_�t�����Ic�]�WafM�7�pC������^������ߖ�7��9��nU�z,�r�V0d��Hz(/�gW��M#s4©q�Ձ4n�^&���c�8���T����}��c�F'�P.k/�m�rմ=߷�X��L�7[(�x�0 ��6��w�'�:�J3)s�C�$����U���S����F��]�ߛ���c��G�C8C���*��3� �C��oR�d+p��9v��60o\�,c��R��ﾥ�݇��s�c��� �g6�� ��$��M(�S�h�/��uw/\s��Z��*�ۊ�wS�z�%�~���r�4��'��>����ȵ��-J�p��47��S-�"��@�m`n��=��cm��������H�5B��-��.��)�*��~�<e\�,I�lhv9gm8���xT�h��(���w_S欁Wh�e�z�s� ��oO_�}�&1�V�~=2Ƒ���e�L-�~���2?[�ڨ��\�w;5w�`N�B6	o���|������ÒSCn������9E�e��{H�Wd(t�
��}��x˦�w\����h()�6����_H7a����Y_Y*��iX�B�K9K��Q6�e���'��;�usOLg+������	�M�&�Κ�~�,�e��*�X1� ����ÚA�Sey�'�1�>R�!}Ĳ�'kX�X��Y��s����h !As��_]˹�{��)>[��O?��֌�6p�;M��WJY�V�tN�/2t\L��$�U%0���"3��AH���[`�a6�@�d�O�<*Ϟ>-���M��������3�A���~����π��F��&�s�w��|�}h&X.��/��%��@%��>>��{��A�+X�杂���q�b��vǻnІ\�!�Ɖ���X�Ҕ�U=�،,:ܢ����m\[�W_��������睆���3���@������YD����yZ��2g�N	%`�Ą����p�sɕ��7K�����A�SO�4��ݡ�<#�\o��g��˽Q�E��n��Y�y)3��B�����,�Stq0Y��*l����&|>�C�!���`j������?i����(�R��ϧ�X"�Z	_��Џ��y�.�Dʹn�,���xe����Fą|�_/@)h4�ɡ�XĿ����{)��<��v�et�n���>%�9��l*.X'���7���?V�aY��`��b��2��Y�H�G����	���C6ъl���FZ)��B�&1�N��^B��ll-q?}�{ALmmD}	O����l��gO���E�$�6�IuX޽�	� �k6<n�a�!NǊX�Zij�E�7�1��͖<�	�������/��v8D���(�Ŀ'����c�y�IC?����Ա	u�g�|&��)�m��K���t<7��`:)W�I��7���>]�׫�_�#hg�z麰h"K�S����*~I����Rg������ù�?��[�3�+�cվ �����~���"�B�J�]�hJT1Ux��R����H♋���%�D�K-��n��E��Yg>U�����b�F�m$�HU],�p�u��d)�v���z�u� �����>��V���qf�2O���b�*���F��g,��E᱐��-�E|�-躼�g� �H&-e�$<A��{[;l�Re�Ɉ��{���}p��$Tsv���)өx�')t=o��=�Y��k��G�m���ML
�6���	%=�(�G��麰��v��-�����v׌�~�O�3��[v�����>ǎ/Sm�13�K�4���}����1$W*��X�g���a��1;~��gF�����Ԯ�+�ހ�4Z�lf�Z?K�n��(��Z�;$���u��&�mjq�.%Thd�|�Y8�r4佮����V����B1J��vw%���8���?����L��hr!���a��3������;��y���w�{M{Q)i�E��s�g�"`�:�t� ��a�����b���J�䶻ٕP�?P\z�v�Kw��g=��?���!D�R��b�@��7�Tļ�QĦ�hsd֎؟��N������p���kz���G� 3���HUM����d`��m�D^ه%�\��Py�.$�̙�R�w/1b��\8sb�f����8!��Ky.�������i�����I4v_�ad}�p�ߒc��	ܰ�G�BMPY^ pK�h<�shd����HѵݪQ������D���e2�=�HnEa�/��,�}���0Y�vn�D��Z%>#^Rp�n�BG�:s�JA��=��~���0�=-�vni��N|�L�:��B��Ӈhsؽ�4���\0Zږ�KO�9]�s�Sv��=w>�PD���;+(I���n����piX��k��k��'v�q���5l�6���B��Z[��n�Q!���/2r��b�������_��G�����e(�c�^��������!~_�v�i��s��Md�����P�f<M�Wؕ���S̷wwj����ǠL	�G;�)�c�;��\�pЙ�=(���Um�����:5c����<�0l�Tk�>ۨ�[ԅ�8��N���*T����}�4`�Ue�ӹ��I'h���:9L�wY�.�F��`����/^����g0%�l��:j9��k��MR<�u�,�JݻP�	%`�&��>���l��{�WY��և]��Ԭt�RŀxP����}��-��	����������&��M_���YVx��M(0 ��<)>"{�$�9�_�SlX����wi͸33`Sd�MW��������zp�9:e��	Zo��p}�P�qg�Nt����!xS ��.5
̷�1�m�m�|���tW���1�d6�%�6I�Sf������GXM�< '��x��,��s���K=O��R#�K�5S���g�d渎��?�@�=9�g)���i�Ǡ��x���)�^�l�^���+: �b�ؕ6&���%�����g6c�	B��uo8v}�f���'��7q�=�)��"x� ��W������/^�(1hpu��.�MQ���*^Nh�Q�c����6!ei���HC?�c�]�}o9�~��� �g�45rI��W�:6f����,�ur�� ���&5+���(�X��(w�47����3���/_ds+�����R�+��Rxc4�i��E7~�QjQ]�T(�ww,c�\�ww���U*�7�Xh\�`&��6G,����꤉[�x�	��g��[�5g|��^�%�]c���L�b���W���^W�om9d7Urx���H����3��k�t���h{��F>赳���HP�ر�?!SY���J{��c�n&��]�hVp8a<�ɸ�\��$b��]V+�0o3 �����f�4-�:�*�+Wpz'�Ų�F�m}B��Pz2�g&֏&�u(�o�xS���-n<+Q���|�*`Ff��^6�P����J!3�����`d�\�}�O�eC~��s��k���̻�Ae��rKxL�o�344�!���C�5����R��*̎V��Ϝ���:`�~���z]줳0H��s�6�.�qU�jB8`Uéݯ��{!�ll%~�y���(�q$�l�&g?�JZd����|BA���L���d+9@:�� B��(����8k�T���Rl_�vspc�_9��t4���|�HR~�9Wou��Ʋ}u��.��.}32WR�$:�S�~o�a =K	����Pa��.�MOR8���4�(p�f΀\,���G7������QY@�w�[7Y6/uY A�~�f�xc�d��,�4�	b��c<�f]���#˾��d9�Zt U�z���^��%���a9�VSI^g�7�s;Kt���(��ʔֳ(�(�}�9d������pד�QyD�����NA�_�i�u�
hx<y�a���<[��ω1�9gґ�W��T<2"�F�ac���	`'컠Z�M�����JW�NT����۸߸�'�y�n+��C��D���b��Rg��\q,j��M�Pe�*4�Խ�,5;]�b�a>���T���Hu��(܋��S�vRL	��:5Mw�%�N�ࢮB�Į��(�������1.^�yB���M�v�,�=B���=����5M�����l���C���M�2�� ۊ����ڜ��ח��X���!�Z%f1HGI��}�m(N����*��o�r�� ��%e}�w��#@�x�Ic��3);C"�H�BQR�y���^fv�1~x�y��h����������85��[Q�(���݊wh�9y���p��}��]����e��C% ��jpѼ]dn�y �� l/��
�F��V/\�̈́M���FMf�&�/<��n#�RO��c`7z��u���U�c����
�	K����C��7ڡEם�ߓƅ�?���i�_8짳�n�����r���^��� L��G�5D��Z�8XE5 �>��{��)��5�͈�+�n���t#��Ŭ�gQ���H�g�L���A@��R��|��Wc�u�Ր*�g��t�����z�Χ|5��}��r
qW<6�4�P�C�bbsb �v��nI�ߙ2��꨹�����K�rf���S�(�6�)ox{�`!ͱ�lK˃B��i�ԣ.w_����M��h3ITy�3M�þ��,_O	�6�w`H��ρ&'y�!�V&�/\i���G&#{����'�ի��A��p���m���P^፦�n]��ۻ�Qڨm<�T BWl/�U���3��!>�b�Ae#&0�u3�����m���9N�,ߙ��I]�K2�.��rWt]�8ƽ�^���N�D����*�Z��Z����m�g�� *!�!=��Z�R@�k�M�e�,/����6�9���%6XS�g77�ym��9�]��68�>4��OЮ6�R�~b��2��S@v��E��^C1�2���@X�K%�{u9�{}���"�hL�-D�Ў�me�
�AF���.�b����ܴ�3]���YĪO�yh���YЕ%��(K�H�3�C��f�U�ߔS��%�����NQ��Xv��jJa}Se��ϐZ�.�p9c��,V�mCa9=�}�$��ӔN�'3��/���)��d�E��bj�T2���\S��Y{L
K6/VâL�����Ds�]�wG鞁�/v�?����͵tfO�u5���j݈��Az}}�g�I��)-����������w4æ�"'�M�&�څ�!�f_~��m�@7��:o�f�����6�:;5\c�a�6g��:H�8�K�7�ᖓ\}4~>���qL��>⳾y�[��qu5bb|r#�{�8��?�:l4���r���J�����B�O����X��>|���I���As�7�ٓ�Gu��F�-�	c�8��䣧4�]�7�r*`�����^�&����C�'��/g�Kf���))KV|@�^��/T��R�9��� <���.#�΢-���2��w0�	�E`�Qf�S�R��{�]~<B]���?-
�]��@��j�f���S��n����e��L�0��'<Sq������fϕ�˰>�#��S�����`����HK5�S��2��A�%-'��M	8Z���r��R ���Gj��8Mvs��'�n���7�������tNz���;��Ca���{c����"��j�K��%�L`ӝkL�B����\��֌�w=�/�����b,����̒ڸ����[�LJ4B'�x��,�*Q�;���~TOذ}��9�^�~!�?��/囿�����i�ɣ���p������t߃���Ǖ@������{��2t =���Jg��8�9Q%/3�ޟ[�qg;p䰏��F�9V]�O&�\�dD��h޵��o��v�`Y.��5(w�/���b]�+ي)=�H{(1�βL��M5��bx��y��nZ�K.Y��U�,`�]LS�"8-��j>U0vٸ���٨9��n��є�Y�o�UF�;
���}��7�^u��9�Ug��-P�}8\��V�y����5pg�hbB�g�{�)}�%���5W�ì��f����aϧ-���1�v�̀�,��O��M|��q��W�^�R�����Ϋ&Y��D���Y�؅���b�e�*��s�Tj���%p녝�+}�����e����_�9��u;��?7��Z�8�`z�_+�6���*�_g�
�#�#�Ӓ������`�}h<���~�e���_�Z��7�Y������'�'���cܛKV>�$��4G|؈�Bh��u�����|x���Pw�k4,�܌�S��9`2$���j�S$1c2]�خƲUV�m�͗N0��i�6����T�.�e����^}X�����]{���\�I�n�@��]�Ml�5� ���4�"�&y�Ys��[�s�k{v�%48l.�-j����i07�qHuO>8�59�z���T!���%��=y���"�kP�%q��4��<Ņ�Qhӫ�b�,�>�|b��C�$W�<���ܙ���!7��Ce��I�T��C*�Ҿx����sgM�HՈ�����8*�o��#)R�&E�!�ls�!4*����8�1�J3�T�yiǏ��Qz��� 泇L�w�]�p^Nw���J֕��D�r_��뻒S}ь�T��G�ݒ��xF�{'�Q������7>:
�e�i+^i�R��'�t'd|�ʗ	���o��a�~�͟yݠ��� ���͎A)o�(��sG5r�.�Ȉ8�ޡ�Ϻ.0m���O�hl6�3�������pfR�u��aY4�s]�>�u�kI %Ľ������� ���ڔ`���U_<;ۢ��P�3�濐���P�YQ��n����\����]�t�$.�L2p�%��2��O��mb}!��w���m%�jb9����y�/������&��R�?gg��O(=�|Hl22B`R]�8��a�?��}��;�����D}�$1S��Rms��1s]�q�\ͪ��m+̲D�U�T���f����Ec�t%�M/5�א��o� ��a8�S�^\_�0*�]���hT�rR�'�{`��:S�:�m�+iX$"(4��I���n�θ��c�9�.�;�6s ups��o$�k��h�o|F����ld���`,��5�h$%�ˈ�3�E���C�~������R����@L8t�˗_~������4�"��S}-٢��ؔ��@zT���� ������勗���/ʣ�O��n���gR9\�/��V�����p?��B����ϼ�e�����錴�-�PT����k0������h����l�T�J�D��_f��T̨�����0A�_�Li��XpΜ�X/"���挟 x߬������{����Qx�=ţI�x�q�)T�?�z�)$3��]t�,PHǅ��qf��lsdh5#��jg:���9("�.��B
�׆Ї�.?�9�uJ%*o�!̬b"]<��b?�>KEV�'�'%�Ɨ���j�&��h�񉮘��F�S�L)�7.^i2�R����3�E�n��5r�������
b'�BLnͲȰ��6�.J>褶�67��f(El�
+x�K�W����{PE��&K�m3����ʢ�7Y�t	1x��H/��f��1�m/x��<z8͡&O���P��! e��/w�i?^�5Ƥ���'y���g���c�Vm��lF�t�����,�ǆ 
� �[`'J��%{�}n2�h/~]��P!������}R�l4����Tw���3�_d�bL�*i�m����_Iȯj��6`9:�����.}�g�L��X��Ew���B��
��$K�,�{l�&��T� 	��&�z�,���(��qM�
��_]O�Ti�K�MDl���y�q��~��.n[�����xN�V�G��t.�۝/Ev lWQ��!k*��M.�>t:���\��fS�l�z��(Ê�#38��^�Ao����'��Ԭ��˭��B��FUY����m�p��~�����̞��f	8HP�6j)�>�x��Vh,u��rP�������1����M�^/���)�C%�k���`�^��gyo-*�Q��,�a��yԤ����~��|l�nc.� TS�d����
Hh~���������U��@=���:��]i�����'0���~���Q�;��k�U��Cl�����Q����:�1�RM6��Y����jΚ���o�l�(�k	կ���s#a�c�Kf�=�[�@���qb[?�;�5SSi$���$^a2<-;�c�c�D���S��x7j/��9 �qG�������<�8'�r2t�D���J��R�!�ʲ������E�ϒ�<ϒ����� i̗__��q�N')�ܒ�b��ˣ�kBl +��u��e X�|��*<�y�tp;�)CQ�3�����Z����R�f� �����i��Q��	���1�6E��(9��Q��H|�[3�]	a�"c�M4�'�RJ�Q���j��Is��&�*h� ��v�2q�7R�u>���������Y��ZAs���J��)/���M�z���ܿ�aJ�'���d|�K�0��~]��g�V��φz��5@�f�	���۷l.=���m�Co�	 X�-��ޱ�艳��YM�PI�C�4�[�D�$̀b!W�S���Y�Փ�����<(y���ѵ_D;��`��"�L<\	FFKZ����<L�q����_����@j|����T��T����6�H�Klf�6�x�n#۬�(��Xﺰ>�$�'N�Md	x};g��,�M�}��������f���5*Q�8#�8��Sן��d����k��ݐ���@Q�Ǳ=5g��ܐT�J�n�g+��ؤa{A³(K�_�eI�mp�c��׽����A:��o^_�#MM����W�����:�GRrpo���.����<߀4��$[3&� [Z3�kQc�<]���f���#�>"+��ב����$JZ,0)?%n�N��%� ��*��Ǵ�U��9�m����?� ��__��ZȲ��p# F�P�<��w�/�:�vq8�b_o��t�v�
����(�C���k���Uy��>�A�'R��C�o=t�ѥ@��_��_tpt��4��i���1�T�`P�hZsQiG8k�	I3�R-�&;��7�n�e����^���)|bӾY<⒳���o<����������w`�%�HFj��I�/K^$/�(�TڍuF��7�X�U�y�sT.�������(��	�c/�Q]͘ư���Mg0� ���G����o�q�@��m�������0P�� #��(cn�򴩴���Ƹ�8p���,�����v����g����,�<__2�f X*��aX��O�١	�1M�I�s8-2�̶G���������W_1���p�!��`0�\��e��t�����!d���b��fE�A�ޢA6'��bfe���P{�$�Tt6!�Q�IYL��NT��TN��'J|+�Vq�O�	 tT�g�a�yz��B��J�Ð
[`\��H��:����n��:e� �P���De���~����Nl�]�DŅ���ߕ�?�T��O*_|�"�t��@/���˗Ϲ�p���:ʜ�Xd������퀣J��&kV��uV0���nӇ�~稵6K�jIVG!4H1��0x1l���cV�K�5�jcƾ���RfM��3��y,��?g�;[��f�Os]vG�@]r�i'���f�40��M�(:��&̚��@'u*��e`�cJ�cHs���$<��{G'������I�f�m5�H�v�B
��S��=d�J4�I��1��!����u��t��zV �]4AS:dF
[i��w�ҕ�9�eZjCd����t� \�=݊���!v#M���f���<�I�G������P����=�s�_��k���oZ����`���$��Y�aר"uY���+�sw�F9���k����L���6�"��Y�.��Vܶ&I�G��F�a��;��.��:J~�Zv�E���KG�g��{�dR|VV<WU��U ��!�f�9��Gj��,�ϲs�d�Z��ͷY~���Dd'�:���������?�R�3X�����%���&�B�<l҃���� ��m}�Q���?SO�_pN%i�Y�0��J��д(�B��ov��P�v$��J]^��hV/�s�e{�->�m?�&��T���<RO5Y�jR���S�e�ZՄ�/x�I�fq�3��1
�%8k#
�#�qc���$o��I�&Q�ȒX'���P�����/n�Q�ˢiJ�"F3�oe����	@� 4 Z�!T����Ff�����$�X��H2>_��ߤm2���w
b�އ*�)�c�@Z�l��Z��N�4��ʦ>���q�`�o�����x�u�d��������� ��s�ϟ>�pP>�cY��u�Q%��J�a܋���sS�;>��'���C7C���ǖ��!��������~���uX�\��->�` �E�7�$
jʋ��lN�Q!ߡh�Tr|������1(v	���0C�`{�w���tF1�I���I�	�k�Y4��CI��������������tWEtD� ��jGK嫫�`���9t(��=����CWԤ��q�&��N���D(�Ue:> �b�J���d�P\��+vl`9?��PɊ��yeD��V��B�^��ح榳x�x�����Z\,��&`lٷy��M��\Pu�����\-��.�ۛH�!�o��聉h����]�n�˼������4����,;c1u�ZQ��Z����I�nd m3����G��P4��)'|���Of����lP���O�D9�Qٹ��9="ˆ�?�ݬ����=�D'�{Xb�k{n�/�|�a�zٗ�5��=���r<?�I 6��o��A����ޔ��U9����3��_�_�.���o�����J��=����|ï������v#�dx��l1��Ϋ�H�`z����c��0d���7�	�K�/is�A�,`�{x�A[*�!��{��P�l�z���r 6ɽ��)J��NCW</[)���������7�P�z5a!FB�,$h=)��?��
��x)���5���t����C��S�O��w�>�#	��X��|�H��ʺ?�Y���2�'7Ot�~��E��ށ����9�to����E`^��}���3$?�ٟF��M�i�]�4���:WJe �J��=���]w�����׃��������j��GK8�#q���b%M��q\P��4�T[f�^u2�2�+K�j#�,���fLS\pf\�$S��+��D���mLa�
D2ҫ�7k�P��_U���ØD��R#�s��yR2��Jz� 9Dw�n��4iќs�۷(J;)ȫyR28��o�Y�2�4�ayK-��$�>�'M�B�ew��3���)��g1#q�?_�|��!�"��V����C�QH��SŸ�/�B�8���Gтf9����e��<�����������A�i��y;�[ȕ���TKF7n!�#z����[e�O!n����uMK6��>{��\��g����r����t�����0M�qm;�S�H&nu�U^�C����wT[S�;��V��� ��ɗ�LH�8)�L*�,p}ʺ:'�:�,�r*'�}���(3>3,6J�r?u�[|>�e)A벹�ț�kd�����g~�hI���RZn����@)"�s6�aA�w���)�0���t�Eb%|^�d7ӯW�ϕ�K����SY|DOAY���"�OPvVS��%������c�я�V��3�1��RQ�W��a�fB�瘩�I\�(u�=�XJ*f�6eՒM���w:�B�eZ��̼Wa������6����v�F�aޯχ���OW�AaS�^nmX?�<:��%m.�ޔEE)���a���c���o˟��g\{cdop(e�43�b�p9&yw��^[sv�B�Y����Xr�qHz҈�,�I�{�ξ����!�ክ�U1T0�䔇�R2����!z��7��`��af����k��#��j|�/߼���r�&W@(�?X	j?��`p���T߿���^{������~&�OX�G����>0@���æ��g8"v�+�����7Mn�" ;k��T������	���!�M����Yzo�3h��O���P�p�k��ek����H��y��@�e�����eWU��[��rN�x�¶��
$��!A�N�At��<�NJ��0F��7��]���r�w�N�*VbB��VW�� :  6*S,'��H8��x/�s�;�ŧ�ʣ��ga��fD=�+���pF-��茔��"��	xв	�����B���!�\jq���I˧����~\�u��k��I��پ���*P�@
��}@+��(��V%�Z)� ���/2��t�}��b�GyFկ��:�W���s���u�~L���ambew7�|]e�^{^��{pyq��)~3�}Vu��O
@��Ï?��u3�6a���l��q�j/�?���_����/��PڋS��Iv�v'Nx�	�u� �Ǒ���߽�P޽��̖��~��[VT�r�=	(A�&����(���/��=�]tg�!�4�d�Ӑ2S"F���&\Z?~ИiF���m3���8�A)�h���3��ϣbl.��ϕH[�\M)��y0�a8&�h<�. n�xn�U�2u ��֨&O�Y�Vt�hQKB	MgϘ��V�lr��f�/ޠ)nR��2�M�:�T2�&�ˉ����W4�{,o&X���X��ns�PrZ��mJxqrJ�Up��
��f�8�Z7Պ\W�{m�SC���y@SD9~>�O�^=7g��4�����!/+�R�>CC��D�ppM~z�;�������7���9R�Z��E�Spc�ɀFi�f@R�?Kڍ�Me�M�;�s�˸^J��Y�E22z.	{g�z�0�;��hR=�5֟���46w�����˥=)P�^�0Ĵ��P��l�*����~����y� ��	�q>��G�l�n�6�sQ��`�m�F�fӁ����}y��ܬ�2�?��M��c�m���w��r4�pս�B�K�*��{-]	�H�����s'�)CE	�{)��,T:���GL�&��}E������l�潥�x�,�=6�`���]�v�Z��v$�oG��>����s:�Gk@FB��>��V�g����ѯk�3U�?4'�!ʇ�2��F��rҁ���3��s��`�6�|8�F`g�ZAR߆ �Vvִ�ݳ�83�]C�1⃚v�sa�E��T�`D��4n��4�2?s%����Y*��e7��M*|f���Wh�K? �7���z��xԟʻ��qB�Sn���fC��^e9�q�h:blL4CAhR�ӚA���*���-Az��sO*�l�X����|ٿ'���Q�̂���0�3�i"��pswσ܊dW�Q���$j�'\��g��j*����@O���v���c��_�����y����^�� p��~�l���ՔjY�Y��v���Bb<4��1g��z�k-��x.҂m�h\�f���JVV��[����Y���Ɵ���j{6+ι;D�:�Bd���i�X�g��#��.13���aSO�x%���n��3�4N��m�B�CU��p���=eY�ʒ~�������$6�%�X���`���Y)�l�o;�nrK��i����Ũh6T�nˋ�K��P������}��ά��E�/R�@Vfp���G�geYH/����\B�c���ۋ���3��'>�tT�3J��)���~�6 ��J�_hW:�e�v<��Jz��(?���~i��8:�e�ؐ��t�H�~-c�3�ނ	��#�Hdk����UFw�̚�oY��f\X�ō#/�6��f�9�*B(����Ca��S �	�����)T������UzC���|�����GZ�N�Zsz뱂gX�Z:�;>�s�:���W����G^�o��.D�!Q�r,��j��{������q�xآ�@Ѹ<��Lٷ��C'}a$	M �M���P��:��ڥj��8Y�eChї1�t��3��m���|������ ]��ˈ�e���5_��r҇e��y�97�D�{�ʯS7+�R�8$n����6�'&�gG���K�»e	�)���^Ä���Q� �LE��1�h��Q6;�>�AT���0���Tp9�MxQ�D3�+�[ݶ/���N�2RRg�K,8�b����K����#�C��?��rd�ܯ�l�G�����'�4wv}A�B)�{��N1Jo�N��KS�5��KJ�d5��՟Ε����J���1�����'��a��.h=��@
�&J/i�rsc�b���h� Zj�ou�#���Lg�y���4�7wA�ꎙ����}��Wr� �y���~��O|߸N���(]�h!��y�|��oH��-�8�gP�w��b(����jO$�㾜8�o������	6x�q�q(aR��_�z���ua�04U�S��	"��,�.-�yr ՐSf�O� jrWҝ!����b���]���z���P/;�\>�8�6M5��l��q��<�џ���X�,~�c������Fi<�[�	(3��ɀz>�o?_���N"��\~6�Ɉx�	C�*z#��Z!���/��3Wـ��Aؽ� �B�9��6e;n�C�I�u�x�l�M���\��=�)hҕ�w������X�L,w�m����^S���[�ku8�����.�-[#�LϦ� �\�,�`o��V�-x����`��X���H/�˞�։8��t[n��<Շ�~�ݔk��K�O#)>$���__����%r� ���gϢ�\��ׯ�O}��%;��}t�1G��� ��<���5`��gӴS��T5�Ƶ��\\�usuK�`�9��c%2��u��ր�ۋ���ʂ���6F^7�������"p��U�2=�8����u7��I��zŠ#��j���K�L0{�B+8iy���d�ڝ����0pB�*T�b�$F�}}�taL���ĥS�a��Yk�l��j�ۍ;���}7�6K[�W���� �M����\%�;��җ�ҳ�fP9}��!U�b���	���C���%��3�����vI�r4$��گʌv{!�&��9�Ϸ�8G���w���^�} އG`(��}�����R��#}���9t<n�"���mG��"P��ȱ�<!�DOz��	q�f��<<T�P��*i��N|O�D B����q�~��SD�F�#�5~n䆞����Ԥ��nI}��	�e�4K��V�]�뿣�͉�CYM��@:޲\����=�;�#�]�<���؀�&�s�ݩ|Z_���X�{�#�+Ϟ<-�4+��!#�QI_���01�����oI��D��F�i�M�Ӓ�sm�<p���Ȱc$pf� �#����V�B�<At��3��뿠��
�T37G�e�a�Wql�����J���;8�	��X�t"8X������O�Z�@��Νx������(�}���6{v!�m��^xNf�࣮k�4&�s�G�֞<eՀ�;�`�Y8�LD@�n��נ���S�,0_g�JTO���{
]� �Q����;��t#G�C��{��%;�K�l���+�ge�m���=�v�Ӎ���H���p,�T��p� ��N����~� z�9ԬL�7�#q�le�j	�Y�)n��S�eT��RO$�"\H��9:��C���n)�#��F�3H��x:��x�Y<cÃtN���X�?��%f��{�7��Ԣ"r���fp,�:tB�o�� N|p�DVq8�r�i+�[����T1c�$��;Jm�y�.k37�e���=�C�����rW(��?���h>h:�Tfb }���~Q���"����>��Ȳ�ZK������bW�"����!��DB�}?���|�-E��e� '*�J�i^��� ��ei���x���Dk�
�Ŭ�k �/�t8��C���Kwpc��Ox����.�"��$䝃0K�&}`�}[��)f�'�g��0x���D���d)<�9>��l
�W#!��m��^3dH�a1f~�=���h,:���?d@���+R�zjZD3��k��#��m@^�>�!��p}���>/FbI$��Vs4��,�9���w�>���t��e�Ϊ%͎V�!?���:Mj�Z�hɲ��?>�Vܨ��*:�#g��'��{#���8{��(�v+��#�x镲3ɧ���r{Y��ip(˯�}��өb���[�iU&/�w�$���\�%�P��q1�U��c	������=?3��NQ�ز���|.�1�w��@��J~��\\��33�ȼ7Y��;>3��t#��")��V�_��0]�Y�a��@�,<��0Y������eѧu1�%?J{7�n0B
�e���(�w�-��p� � ��Z7�T�}��3 ��Wgk���8ޭ���7ߕGk;��ײp=8���z�M��Ĭ�Ns���������m(d��'i�6'���s��g�5)�����3��ʏ󫈣+]�2t���p c�ܮ��6�`���2�����e�����q���N�u�~�D��Y��=���I������~=01��E���3 �Pv�(�Az&}ӏo��ϧ����X=i��-��W̊��ɫ5��t�~��qu/0�J�_N�����0{�+�8W��vX��fu�ج��2��5��|��N
�e�}�h�Vg�_�lʥt�Wq#��+E)���.���X���+��ԑV��x�&��'H��$�)��8�-��<k����_Z�')<��7Ew22�>1K,� ���OE0D����3�!�V���?��,W��9�d�\�N�x��K{����\ҶX�+���r>+�-���P��W�*O�~���R�ϺRx8p�j�M9���Y&"P�Hh 0K]����r�0?���+L6�P
b� ��)��8�0��a�1���<D&���r�JE)M���FJ�x�!�"�"���Db�߱	�Te�p��ʺ>J]46�m��%_�M/�/��V�. =�����,?%����:��|��N�l5e�E��,
Cpx�~z[���ӣ��E�N~L*�
�ڇ�2���X�L?S�l�W0ޢ�����J�X�ptC�l���D�k�5��!��
	��&�jk�j5�_��f*Ta��v��kU��5�$�K�� ���ա����#��AZƅ4�Ds:�嶛b!rO��> ��P�@�����xJ�_�fx�F��F �Nx������t��@(?�0�t&��)��L�"l���L#x����>2��w9^	�x��/��2ũ[Q�X����`6��%)b]���� �@�TF�Ξif��:uM�I��u	��K�ސNl��ح4�(�A��Ե� YbV=Z;(s��ofI�s}�����͗l,2���!�l<Ċ$%=�h��?}�Ƃ��q�76�	�pw]4A5��Tf��?�85/z�F.~z�jW?K�v/8@�O��!r�C��o8��Ӷ��4S&n�.)W2xW�"�0�/�X��/(y�5��;>�ӷ��cX�@�p*� ޯ��ǈ����>��]�%s.�c^� �J���J����� ��M�9���.�UL"5�9Y,��[���sò)L���M:���S
�<r�Ջ@*��3� �����%���R�����X�������%˩v���#��4m,��.R��_�ݥ�0́D)%tx�<_X���(ZL���HV6��`��ӧO�b�OI�
1<W��V�@Z}*���|;N��j� i﫡�b%�Ab�k�i��{Q����5T do����g3�jܟs�?7D�<s�U�WD�/X�"'uS�75]߰����
��J��/�L�`�C�h�|�O�E]�z`��֠:-�3 Y��`��ki���e� 2u]隣���ƳJF����^`�Iߑ*�F"�nsM��.�%��-}����j�,�G5�+�IW�L
ƈ���R��~��5�SWt��W��Ϟ���7���X����L�v�]VbY��ەTTG�̤f�C4g���^Jp!������|J�̼�ρό�@e����Xf���W��}0���ۘ�:It�M)�J���ҽjY>�-xY��7�����T�п��\~��bs*��Ɍ�t?3�ӇQV��ܥ�T�G��w�������rt뱩ݍ[�8�"�*�i����io��\�%R4����Yw�W�(b�l<_@hb�/2�F��ZZ��Ȣ�č�f]ko���c����F6��[��XJ�����dKwy���s}S��=��\6�����.�.,���~/'H8!�t⼣���s͒ݑ]e0�肩�k.�a d�o|Ko!d�����Zֿ
*������`G���OL+>e����~l����{7j����
�,�ݷ�G����)�9��%�%6��ᥤ.����2�^�1L� A9l9|��Ff'�"�����L���v��)��(eia�SU���)R}���J���K��VL��!�J����8)��H��j��f�7Q�	��iwAO���m��ƭ�:}��6���{�s1���7x\l<ov��!�g�ߛl�;g`��1���K�Y/N�ǛG�|��jR�u�b�1Es]��M_���������m��dƅχ��5*NXX^��LX4�fA�6Ȕ�*dY҆���ڮ�U��e�N�KK��Ǔd�,ivY|$*�(R��N?嵰�@�.F���@�[GP�� ��rs�D��Y���ƞ�����g���t'x�� {���[Q�~�Gf0����}��0*{�Vo�n��8h�%�U��Uɼ���d��\�n�o�s���a=�&�S��2��ϩ���lb8�&ɩ�]�v��x�o`�!Z)L��- T���3�%�|�09�/k�R~��P,H�頳�_�f:`�T�m�2�x����rv�����Ϻ��E4���,80�H(>~����NR��y�sB�7}$N��#�ָ���@�X=�R4����v��ei�����E�0�F���_�	o�܁#1�i̩'җv
\%��"�Rr7�*����[7֤�NI��8�Yj�<J���/a2��bx7F�$�[�i�vV������ä˛�]J����/y�T�:�<7@7���k@'�1"Ld����pee��l߁�N�L� MkR]4g�oAi3O~Y	+X��%:��LF��pB�U���L����c��)~��pPM� `��E�㚁�;�;�Q����pH7�MDt/h^�s⥋^��%��z�a���f.��"���|`�]m0i,4���`�HmG������>Xsh�aW��*�;l������}��S@��tnR ��+�J�X�H%�#)�A)~}+�kh�b����������'1�]&=�ׁ�"�i��My���#�}V�����-a*Q��Y�89�b8��A6Ⱦ�	��'�H���KC��Q�
X��h*����s��/E�ei#q��=�r��m�ƛ�%�˺:ƣ
�7W�\w��鐚�xFs�\o�\0NR��Y���i�ޝ�:fS-��l��X��^��V�y�0s<6"тZ�ϖ��p��A��8%��
V�W�,��rf����5������U��R�@��SH,��.���sN�.%H�$���/�@�� �/h5�f��XXeL[4)f5�B�w#H%���9�N�#~�?�� ���v��0C	�����FV�����?���Ebm|�y��xFjtL��vM	����½�Gy�r��_-,0��Ti��K���?�JŽ�3ŊG��I�.��<��mGضD5�go$��~���19�Gf��{a��������zj�j���>����ә�k�j�n���@�ဓ�6[�����Wt�#��sy�KWߚA�{k��zԡ�
��:���T�pQ�"��uwY�7Yͻ�w���q��?�ڷ�����C���ҽi2�������� 9/�������^�uQy�R<	��%&b斋�+��){��м/2�e��½�W�]=����'~L%�9ic���=��),R�I�Z6㳗R�	}]� �@���b��q��7:րK��3�C|����j�@G��7���Z ���8����:ʢ#ӈ�0D,�~����FY��E��x��������C���x�,��G�n�������o&y��`s+#`���9�q�T�ɚ����_|Ů�N|0[�����y�����j�2���#�8T랛u����ǝ���Yf�%.`̡����c^��9�_?HD���N�pә�!���U���L� (&A����6|���<�f^o[��/1�Y1�3�l��.����;0��fh?4��*���}#ڵ��B]���\,����ӟ���i�I����}�iz�����G/)S�y���:�`N"�k,�"1q`��>��^����w{t�'��)ˇ�t���υL�,<\o��Y�0FC�n�����Ɇ�'���6��|xS��¬c��Xi��ʂ��v�� �ˇݧ2cl�ѩ�FP�Z*�����A����Ä�Ⱦ����+�1���,�Q���gg��ٽ��������i��x:V�� {lP��FA���d(�ݶ�Y�ǉ�41��������ݭ�ҹ9�fw�V�uo��뺚�}%ㇿ�Pǃ6�(��o�a<��բf��T�|w�'��ѐ���(�%�|ntؑ�o�����t4�qa�:�{�q�`�	er�7�CY9�qAl6&����i�{�P*�kzT%F�|%vF6l�'Ա�)�}H��m(��:���ji�rM]�\�P��|w��n�dW�m��0����݌t�L�(���&pȋ���)fW�{H��!����(E1��(�Gԃ��˅�����ٺ^/T��Am�~F�zv�Ǹ�8y��g��N�C(�/��:e����e �����j:�s� w�(��H�E��f|A��z,��٢������׻�x�3���]W��J��`9��:G4ů"�I�������ẩG��_K��u��Z	�Ӂ��m���ch��psh�˃�">-�cn�v�xx��nF�����h=]i�K{}��k�]Rg|�JH\k&���ذndCI5#]�ac��3��z���#)��A���*^;�붼-�^.1���D(��R0�{�B�\W�!U�<���2�SN٘��:�P	t@��>���x�����"�NM �X�H�(�:35��"�Ɋ������H/������g}�K�@0&�u�oxv�7IY�9Z/�^Y�U}����E��73��-)�r�^��'�RqQ����o_�����).�qӒ�>�"�R�wu�jiJ1e��-)XL�
����,�l�&Y6d0�$e6M�������L��q��z����b,M&����Y�#�+�J`\s�ŚL�A�ڮ(-&ޑ>��b�$"{��!�s"�'�a��sp1nz��Ō��S[�"]������]]tf���Q!�G��oK��?c���R�`'��qH8@�����VD�w]�Z��
%��p���0���	f:��H��h(�)��<th�&fH˕�63�C>��@�~�$T	��+�S@��xh�U�Y�RG�ƙ8�<�����I�nQ�����3���x��-��h׃��)o�gM~�J��T�JR��[��'�m�!?p[�%F)L)�e��(0��}�]�	��D&�Ũ|��P�S'm?�^�W'lƜ�>�V&l|]-����˧�F�� Z��(�2%�/��أAv[/�)����4v)R�?�2�s{T{��M�Z��F��W��q�ċ{P����e��!�����m�[m�ϽdV�4�*��3�"�7��e*4W�ጃ�or�D|�f���x�@�MpD��q�0|s���pY�}��^_�	&齎����� �z��������J�pă�Y�r~�+�w*��|�Ek�辎]�߼���Myj���FW��)i(��4]b�5����$�������Iy��%����p��նߡ��ʲ�*U��O(����P����x����͢M&B�P��CǮ�SRZ����A������t�M�K��G��.*'hc�@�Sj�,�$c*\s�"���f�S����X��Z�+�)]s���%S�o&�/�.�G܂�4&���L��V�q��FsF�`�ٷ���R"�s�b\?7�6��i͋s���@�f�,�&x·;�x//��d �葴��xt|ޥ�ƌ�� ��x�8I+�5�-�ğiC!��<�ys.��dш�4�F6�]-9�βvA��.3>��R3�6�a$�s�g�u�������,?��M���D�~�i6b�U���0.�������x;Ѿd܅HI,�6���"��<�$p��Hn6����N��7E��z�u�j�.�1��0�w�dY�8n2@���z%@h\K�Շ���
���I匠5P�e��g/J�"Ll���a���7,�}a��C�r��n�B� ����Z�Y���x�]������^������aF�5ծ/<�ߣC��ɼ&�f쏎�jO�I�����:Y�r�L�"��soO�) �-
��
�E�>��cC��C�����ư��,u�8�Z�'<<��Y{P{VՑξ�r��E�7k՛ ���vsw��u �`H�yM7���Bo�>W>$<O.��Hh&�z8���{�~}��F �vD2�(M(�񳽰�R4�����w�����l�l��/�L����\E-�ک��㸡��E&�s)�SK��C!OЬ�����?�KQs�	��`��K����v�y�K����d����g�k9�o�Ȣ����A����l�\�Ϛ��s�9	8׊�9З��Ǵ�����l��i�U��X��'C���,�zǤ:���}�>�I|��x}Oi����O�r�?k�!
���)X��d��d�_������?��P�k�4�"�/ƿ�e����f����InvL�xw1�)��]t�z���̇d�s����S�=�0��=�� ��P�W���t�i�V���@0 o��cq�wblT�֙b���s��o�Z��� ��=�������E?�( M7�m?R�U{���f���bi�������F��$��0�{��e)"�sl����^�/�q�� kl*��μ��6Z�1�Y+6�I�O^�,����7�'��%�gF�$��T��'�ܪ�i�
e(�s-e�e�?߈�WЫ�i�#����Rjf
�^-T�ϩS�E��6�k3c7?�)�C�)�" k����[B,{n&s�	8��-�)X�2��s -��-.�ES�Ą�"�js���գ1���G��C����QQ/4x�K�B7(�[�s�:��d��`˩�7�g�l��=��4q���kɿ+�I#�����
�G�|6����/� ����e��<�e��[/�A`OQ�ܮ��xw�cҦ=�Qچ�׎�����f�T}����l�1�K���_���tNH��;��eG|;]��W�t+ ����	��l�Gp	#@�z���R�Ė�\�-ϳ������8Z��g���7�b�?�����_S��/�s��?�'3�5��=��T�<r��?�*����� ��Ȉ ���+OETn�I�͇�~�ČX�(�pT�M�2�9G'���r3�+�Ģ=�LTY�V��6�K@H}4@bp���W���﻽ֱF��['*�A�R�֯�1����Xa�Ҏ$�O��D�l\M���(�⳺�aU�5;ż�1�,?�k��ס��>����Fj�"��Pt���ף�����ۗ�O�gO����H����81r�Ղ,���I�g�6��Hy�Ͽd�P-Ӄ"	U�asHƌ;��oERC#J�턹ڊ[�B$�(�Ej��c?t�6��3��Ҁ->(�z��TJ�ҙ+h��|�b![6���R�ڃ`o�A�%F0��r =q�m��%�f�w^ڋ������;��}�(����X�q�#��9>)C|��� �a����2��t7ۮ��{O6C( Ŵҍ�E���|���,��d��o^��Pb!�~���E��̌6���4�����i�C'�R�$_.2㺾�fe��䭙3�ߎ�[����ķ�׃�2�a�Pc��l�y�~[|u��mr�l� o#�*>�fJ���ǡ&���+��H��7sӐy�SU?���� ��_�Z��\ͥ]J��]r��lW�'���3CW��a���Θg���~��L~��fR���G�Ž��2v������e-�R| �{���x�r=��,��x��}LHTRk�hw��׌t�r�v�b1����A�U�7@��A�C��]��R����e��ץ���X��e@m����=������fiTq������9���6j�8����8L�"#���6:`U�3:���Qdx�?*����JL�|�K%BPY3B3��oN����	����u"f����5]��`pާ����[�����-�X<��kg��n�w%@���Mr�
�P����o��M
ŘF�A�'q�.�b�O�ţW��ͬ�̹U2�ŧ�?�RN�(�f"���	H u�J�0���2נ�X��&MVw� yE�Kh��x���d6���W�Rh�y�[@k��$H&�AP�RY�e�"S���e�.�� sB��y��n�Kh��f���6L�K.��RrM����hvjn-uM��.�����P��Jw�j�Ce���i�WS��Qq����}v��ɭQw%TK��RU������{⊪r�}M6����<���a�dm�?X���6����}�G�����Mr�RSr��_����Գ�0k�%�����W�����1��p� �7E��MC�Y"N=�*�$�"�P�A��S���]�c��TJb^��K��$p�w ��w�6Մ�"��5�V���rgxި"��2GwH�n@!���g��W�)d�=E��ГlDy��C�N4�J��!Y$��Q�iߧf=uj�z�e�ػ(`G	W�����PޜQs�k��z�� 
˗Ǵ#~Q^�q_{����3�QӅ���Kh��&�藥�q6�$aL���=���=z�-�&+Ö.jTk��zY�(�LjH��KXc)9�P�e��>�+u��v�'�,����%��0	�5s静�U��o��_q�庾�s���|��XeR��(?^�Pi��]I�a�1IB�;)������xy[vc]�1K�y~x�jI_~$�� �f��/�{<��/�9�Wf1'�K�j�y�1��肋d[��t�B�{/1�#����YZ	:X�3����44��#��	C��w���H��_�L5�j�}�Q�$uC �&'�.=g<Z�i��PY����m�M���iOb�3GެMx�[��/�iRFj��z"��� h�p�r��)�$���G��S`���*�&��KB��jHuu���~$o2��R5�.�B��k��ur��FLh[�W�1��/<�|�g����^4�����T��QK�_A�����\@������?wW�Ǽ�;I�����n��5�O��� +^�%��&�ٝs=�4�P�GC�o�~��t�:����.�ڰe�_�Di"�	��㭇T�H�Z���� ����֦b���L����چ��[qoG��א�a�������H|�,i�y�%05�����P� Z�}�������������=��5�zE�R����.j��W�	r���Sv+�,,ؾ�K�0�)J�6�Y1�g��s�U�N\\L</�7 7'�p�/�do�z"�J�{�F�bX�M��m!��B�,��+�*2��!R۴y�ʑ��!�	(��\2��Z��7�7y��[��t����.��u��zu���e����Y�5���t���}P�z����E!���q�^KIg�x��ۆ����R��qΛ�͗�&_藯������">�
4>��`լ6�֑Uʫ�k?ls,�B ��a5!�����B`=��j ��E�OҼl���bZlϧ\�Y�u:ͱG&Z�Q�_�fVe@���/������0	(�pX�\�7M�b$��>WȍY���x���������7��U'w�P������ԜS6�����I�G��� :�������ǯj6��d�X��s���;�"�ؿ�4��r��E��1�� 	*�;�T:?��xHC�z�#8��˂&�/����٠���|�#ٞ�91�^5Q�EI�Ʃ��O���X0�v��.*���\ov���^�$>?0+����q�z�\���kb���F�K	6��ȠBQ��Y���i�1����"��Y!���ZT��_ڲ��;��ݠ�i��X�ᘪ��ә�����{U�s�싗�_@�	�>O������5����Q�.�0���{�Jpo!2�3����]bddඓA��$hhn���
�M�*5�-� ��{͈[����.�<���{���vQ��jX�K�6!��\{�q����K���z �y�1Qd���XkN<ܔ��o�-.��c��o5�o�v����-���d�qȇ��?�^jV�}0n�pof�d�SV$�v�5�֘�K���Jk�?�2����r/�����C
{0���EeH��_zG�Mz�lR�"�Cp�B�'���u3w53�����������@�]�ӟ�ěg�FS�p��ͼ���ہ�^���P>�|�){f��7%Et��}����чz�V��6�zA���)�3Kah=?��EB!
B6��QXw�f &M,��{ ��1�c��ٓNMT�h�k��YN�%�Q�P0�\���.��MQ����I�J����UvG�]bh��L�R����]��_k �������D��`�j�m�-󒽯R>oq�
l���������	�o��V��9���=HHĺ
�F��Y:���?��8P	Xʰb~�Y�wK�����9v��F����߮���+��l����'z����O�\~�O�Ĭԙj\���� ��ӄ۝���%��	���I����D �3�듧����ʱ�@���EV�2>i�OQ}���򾹖�&k�R?H�k�+՟��T$a��p!�l�l�s��7
KK=/�a�x	��c�<�Ouk�UOl��YNn'K�'�Px- ���@����[�w����������Hy�:T�)ӵ^|���A��A��׍_s~fbŚ��k�S��N٭G[Ķ�w̎�9��w�����@u^<�k���a#%�ི�<��`2�6早A��.U�1�o��7>g��C�W�'�(3�P��YN�`S�����ט�u]�}���rkQ:�[�������w�����|�W�Z)^�y;}x�1f�u?����:��}��+>�RO����x����r������n���E�"�7)��l�\�E�#P�yI����Qohc�}������HKv��%˾T2;$�������S�������������Ì����;�/���۲Y��ڳ�1$݄�O� ���R����O�~���8��εT��+�p��~���w�0uR���������Qyk�.��F�M[&�=w��bJD��8^�Cה<��.�����W� ��b��cu�n߀�>�k���a���f�s!h@n �8

/%O?�@��E�h��g�4{
N�{�pm��(62��FR��P�x��C�'�$�.U�,[4�{k&No�O�dĥI����M����9QvִJ�c��`�ts�Z��`�K�.���_f��X,yYJ��K��u�bė��E���׿�*��.6���L	8� �CO����oT�\b��v��5�89Ŵ@c�b�	2d��F��)�T�G�h遒�N��>��PL�La{b��V�.:�`JXw�SESfO.㗸�pNW#�	�o��Ω]�ϥ��,V!лHܓ���̏W`=����U�н� ��P�0>������I�Cd]��������+M��������'i�-�\WX�#���O��j/!�3K!���n���ϺJ���6���F��|Ef'%��$7Cq?�{��F�6� A���iez�8(}NJ�'��gvIw�G�]�L�&%�.2�?mo�I���/� ���z!�x��_5<w�4�]��b�e\TD�,�ȪjNTG	"�mQSE�O�T�7�`;��ـR��7j������j���A[�|��&�y9ǆ�[h#8��
�u�r"W�+�ԃĽ2�2U���>ȳ����}=�jü0)h���61�&,�8e����O0$'��8!*3�'3�[�Uv��
�]s���b�EriyHu#=��^'!�ԝy��8��Gg����UD���m����Q�D2��*��Z��;�zx�⨮��=�h�(��Ś���1���$V*}��û{����}���R~ݼ(����yph����\�>����zKM�YE��<P�^�Z�6�I-7G�SH��7)
�Ա���zA�0g�?���q@@k7�_�(OR�?<��#�2|N$���6��o�K�=-���>��3)e�(�����"��a�`�!�������z��E���jD�(v]׬�z���q-啷z͈�ħ���3D�/�5��A�yZ\c���E;�M�8��K�8mH��`b(��z�K��ZkVY�OC���!�mum�+�M�/�e��dԞ,aH�ȷ�O�֚e�ˠ_=��������B�|��ݷLp����'E�(���eG ,"CSt��?�Ʌ4�1��T�&}�6879C��.���.��n���g���(Ȑ�ȁ�X���&i,���	Z���E2��	{�Hx�ۿ�[<߽}�̑ɳ�S�ȱ�7X�v��oƴ��n����q��B[�P9���%BWxP�x@2�!*x�ž 0�0�����]# %����Uf����\�������{������\�����=p�?�h �ID�����ޮ�5���,�	Ӌ�/�	�N8�xў���lQs��	#ڍL�Xs�0K��%����#Hk	�e6��@�g��++l�HF�"7,�v9�R!���c�s|�@�k&O�Ѫ���c���W뫏<9�7�����=���6��8�&���
RE*�i�zu��.�#VG���kz��ì]B	��?`V.�[�kҌ`TVe��w���|=�������F��)���*��c"�"��혛�L/�7JgjR����W��(@�0<3�󪊐�j��	'<0&ͯ�3T�橘i%�nn�����O[��G�'}$Ԧ�(Qon�QA,����>=��������?G_{�e�p��x�7n���R��3e���m��;o����n�-Op�(zb?*�-��QP���ܟB�@Q3�z�Qڹ����iQbL|��4�!I����m����B���<�dތ��cDp0:��i@��yWx���"��^d�̍`��ߚ�[k�<�1=�N��sx�OOSޝ3��ws�1��A�Ar��*jO$9��'�fTW��	�*����K\9�b�-��}���f���mQW��sܸ1����i��ά��NL�*|�
xL�xe���(�߮���iG^����E�<������m����Z�xɅ������"af�K�i?̙�k��"˫�G�5�{+�!�#I�=KD�e��'z9��R�A�~���#*���=�^9���E/p�pR�A��v���"t�BP~�6��Y>��"w�ǁ�]$�@������OT�T�2dYfx�-�x|Ц9���C�J�7�Զ�~�r
�&�}ǚu�+G�7x?:� 9�#
�1�u!l�^��BB"n�R~���x�����TQ54���RP�� O�O�K`��p]���h?D��rS��&�8�^ρ���>�1\/n�MVɵ�Re�'�׹��p}d���k�\�z�����+L���%��ѮG���E	w����!j�Ѭ{�]i#��<.���n�P�${:d�����9(�"�W���>̎h�?j,��R��A�ˊ2�ڨ�JL��!��C5�1�>�z��o!*j�1�E���t�rÆX,�����o��S����=���c�c�ӠT������y���d8���yֆ���Au�%9��m�f��e�E�U��D�p���˯gb��?�����-�g55õ�UPۢ<���4����}
�)�N�]�C~n�Q`\?eS�gqlkE1�h*��S��')WK�k()&�A��;��'�C�����N�K�C�7�Q�U�ȵ	�5CR��L�7����ً}�1��:�ⓖ��xf���6�Y/��x�?{X�\4wKz�ħ�0��������$�d����/��ϒ�[��>U�iP��)�����!��B���z.��k���,�0	�a���׷�ފ��69�xZE?`6Q�Q��q��t�!����:3u1֏�\
Έ��H�bͣ"h�h	I�4k9��5�ǔΐ���I/{�x�gS]�y���I�J�i����kR��;X��h!;tl��Oo��FI�R11��6 NR�k�7��>�}�M���ℵz�>4?O9�'-��Zz�le�0N�M�m&g����mdʿ��`�B9�׊m-�gQk_�Ǜ��.iSx�өSGMʶ��-�#�Kf9�NN`�����R�[l2�T���>tJ�c$h����aO�X��-�=6�?B��g��R��s0�d2 �d}�� �7�)���a}/o��UΐF��ǨLB5������0���X���f2&�XŴ��;2�
Akr��H��Xn�JHd�����T~�	��{7����K��
FQH��x���ah%�����������_��M��s�߮�*��"]���z�&W����\�;�Cy �x��R����ٌ��oj��	�[F(ƔMK3��a��ʮ��#�>);%���£�OQK��k�vI��(\�C���EB�d)×��/��և폺�ѫY�{S�-#J�emz5uiYjwŖ���n��b:Q�%�G)�܋�'aP��\��H[9TUt��Xk�wc%�/�Q��{�!� �:���2�� XA�������x�E��}����e��͢jc�|gZK���׽���u�l��~���%�C͎z\�T��e;vm����:��Ld�! �=O�?�qaCpw��?n)�Z�e�����k���|���w�m�w�ަ�v$8�
-��<5:����.�bPo�11HB*��%'�/.뜧{q�Nso?��?�R��(c���^���5����
,�������q9*��������"�,Dh�2��L�\���� �bb@ۼ��F��1�pG񮭐�ŵ."�E���"ٷ�s��-�6���v����jq�)Y;�<���Y*�����(�Bh
{�*�e��l+y��\r�ԫ�k�I��E�[��� �?)+�eD}aj����T�N!]�B��M/E=\ƅ��#���.A�M ��ĺ�Z|�1m�R
���P�{��O"�d�;%"��a���q���:�NX\%<����JQ�#z�bِ^�ɴښ9���Qn,3�~?�=���6����W�'�ɈgQFކ�uah$��{������%�~�)��_?�Z>��!<�i������˧���:�sM�Z��*y�=G��hG�����W�ӄr����\e��$"��혌�LT�	@�M�����4j��wX7q���7t���Ȥ�.�S!1c��k~�h�����<( >!�yē��G�)qx't��l�Qಚ��zd5>��c���mXp����a�<*��Ȭz�l��몽��=���6�N����~`�0x�F��	�d��q�Nb	$���W-*3���Ȑj�&������ژ:�o1ӱ}۴���AB2i��B0<.)3="��qdI��=�m.���$E�/�Ԗ&�[�����ROB�ά�T��e�&�
(�
��8��v���I� ���̶�-])�{��!������W�S��]����Rn��E�7L���U��'6'4Bipugz�V��\t�(��,b�d"��IN"�$���&5� ]����~���X|��������Lr���,2�d����+5S��fm�;�D)�(E���G�g�Ͷ�{ml��3J����M��Ya�uY�y����"���?o����#m�*���Ak3G%��t8t�}�jg�����Ϗ�Tߤw�;2;N�#��QG/Z�lS���17��0�!D������D�E1n���E�#���`�y 
�S	F}Ɲ��&s�d>/<v�H�[�zR6�aC�
2�LC
.��(����k���@X�7�a|����j�����,-�l"�I'�����t����T����"~6u��D��DAG��N�}�E_M˼#�@b�O��kL�k�[j��|Ԓ�)X���S�ӧ�"�xd�`�э�Ԙ��[)�W���ј)NL,��ԉ�
k������	^V�
��VI�^Vh��>�J�P5�������%==�'$|f�<��&�a��&����Cy���HX�d��E�r��&�k����!��I�����fyP�A��W,^<²ޗG�a2�f�6Dv��v{�җJU�|��.Z������]����'|ӜԮ�֡�v&��aJ�C���4J��]���w�b~�Ys�7ôa�>s�+B�r�C�!!#B	��K���Ab�8�^��| 邎���^�����a�I`��Ebz��VFs�Q���q�

�~���e끺'� ���{>�/�&Ы!���[i�Z^�9�������7)�+����9L��d��og�M=��i������Sm�O�������cf
1!� �{�p��ކ���}̺�,��$o�0o]3Q�G��[z8Q�&�ױW\Ų��@��Ȇ>�G����Z�c�^��Q�Br��&1�5�4�
V4&Ɯ�y��G,�Q^&�i5�2���_��~�	�Z=��ez��oi��ab����[�X�6�	���WxE(I�m���Q�����*{, h�F�	����`��gb뚘�a�[���Qdь8Xg����)ֆ#+^[�&�Z��b^��h��3��"�JzIg�圴�p��91֪�d!?<��nY�`i�vngUka���ݻĝ	��
����ib���v�k#S�Q"v`>Je?q��jW-�}�|4��`�����n9�X���o��/<�W�,,�W��ݞ�_ϒ���â���D� ������8�Ǘ�U�]χms'���������:�+<&���u�L�EYHf��#%�o��|��e�u5���*81�R��;c�Zf�:�9�JtL�F��^ҧ�G��(��<�j���ť�"��X�_r��{���� `,wҋ����ʹ��JV��!�j�;x��5�L�!�������:���5�C-�ͬ�e��n��<Ϭp��da 3�!�?�yb����o��p�5���)����=m�(�-)���:����wU�5x��II�d���V'eҫ�^?���b,:�E�2�W[~�~ %ѫ=���^���z��yU~zMH�1�O�(<�������/ϟ�>���z�G�Le�Em�.<WT0R*s�<öם�c>⒙y*�Y�tI��[�
�^����~ȉÊ��뻵g����y����ᑚG����;�4~"�Ag�c�l�����y&��v�E���0���Pi�֎��w�YH��7I���x���X�P�1HnB~W�!`�^�R��ݫ���i��K3�u��׈]"����ۤ�Pݦġ2b�a5�����BW��N<p�?3��x��)��)2�Ƴ�Ӧ��k��ш��k�!Y����4έ�=��KG����@�˗�Klfױc��H�2�e8�̂��
в�G�1P� ��p�X"�ޏ!��!y|�)Y#��^ۺأ�G4gb
���x�/�x�F��ſ�3��>�䫲�N6Y�&���ʎ�|E���ݺ0Չ�h���x�Q��ڮ/����9A^�x�j[���}FyW)-9w�������,J��m07ܱ�{�^�.� �p�w�6I��i F|fW�*�>�Z\��O�B�-=�i��@�cmC���o%ӿ2{�-c��C���_v/��{�*�)����H��O�R��������]:M*�޼mS����&�N~���>>�W��)y��5�����{���+����x���k�12(o���Km����i�cc�ZLY��(Q�Z�$t'y<>�=Fؿ��q�삃$�+2�rk3W�dc�	�~��<���]�γSɡK����G2 ���j[��8����'b��Z��aO��&e�̆L<x�9	�̼aDoS*&�*��z|���;���s�n��Ѕ��T!������5�BO������W֛M�0��U��r\�`�Dx8%�va"�Љ�mZ5*hD�rƶߒ�wz�<]�)����c��<�'�K�+F��G� >Q`��R��Wӯ愼�w��n�c9eY+�(k�On��\#Q����č�R崔�kjN?��̥1t��j�Ք�������UV��ǩN�=�j�ǈ���}-Z��IQ��jT��D(2�w�G�{�����>0jبT�~L`�2iQ�x�ݝҝN�I�R����83_�+��s�$�/���d�"�Q/�6Lh�k���&x;Ӈ0ː�ENچz�������]y�=��a��nw.��R�dR��:W�}n�k
Y����~�B��ɼ^��Qs��
�8�)�,�գ�]z�yq8�E�u75�x����I��14lM��M��݇d���%Ń��#%x�R�][���)����׻z���@C������ol�Ñ"`t>|�D����A�l�Y�rK��9��0u�@0Tz����֬��k�S��e`��\\��^��|,mG;�CĤ#�s�,�n�E����d��Q�
�cL�1����YQ̤��l:R�w����eqB��3Y*m�;�K����珄����k�h2�%tׇ����n��m������G����G_y���Y��G��)�f_�6TN]/�?K��[����bj��nZd���|�}�T��΋j�q=Q��t8�b�!��}'�;C�P0��L'��Τ�X�I8S�}X��I l
2�*xTT��Z��S����Fx�P
�u�����/�h8Yf�;g�G�VowƟ�2C�e�,�Zz�����r
��":KW�R�v��92#���J�L�g̗���zT�kd��,����+��	0n
{p� )�Z��WjѪ��&���0�X�(�W��Ȥ�47���S}�u揊T:�B��{2xs����k�Eob�و��Sf�}P1fv�!��N�C��Ug���t���l�kWⳉ�>dN!<�K��I{+�-�ٶ/�����dkp���f(J���c8<x�u�褻͕އ��{�������O�&	�k������潞���-]~�Y0�w�n��NL����s�аZo��G����x���Uǵ���N<��Fԛ�,pВ� c��ߑ�9[1�Z�1^6.��7����Z�o����N�9�Bwr���,w�I�i֋��8�o6�s)fR��5��9x1�K��U���:���hh�Q���w��d�t��Р,)t�W���%m�ȕsx��L���1��{4'�Z�^ -\����
k�h/��;oLE��\v{e�;U�]Û��=���<�s�.��
��K�H6��@2n�W���ȺB�z!��8��$���s��Z�\��T�Jq	F�J�5&�u��*f�CiJ4�ue��2UF	���q}XnM�J��o���F���>j�qS���P��=��'�֩�hO�u�]�(Gđ['�7{����O}�����*�Y�@�w]3�A��C<�2��Q�0��N'
��`���E��볔��z�u�+[ZR����{��k��H���wlh�I��z���MS
��w		aYϏ�\���%�#��ɚe�˦�[����"#7q�\�����n����xK��$��&��1^z�6q�ߤi9��n�ߡ�������]Vz�;���|����"n����_��c�a4q +Ku)��V�R��^_����	xl�� �Ql�P��fa��-����u��DVR����7�%��󙸠[������}�Sg��`�өꑶP��Hz�Xl�OO���Cr>�dG���\c��w���~|�>K�C��O��AD�%�+�z^g�w�!�$���n����p��Ѕ��xf���� N ��d�n��\0��̈��ez���)��L�^h��M)����.�#�r�!>)��}�U=�5Ƕ�Qц����^��R4��L�fٰp�P��B�
� �ްn'^7����5��ZArܩ;��[t'��{��B�t?�~4Y{z��i��?�遼I�8�Z�*]�D��(�v�l��L>��3�|���H*U���F�7N~�7v�q�S��-r]��I$n���]/�u�Ԉ>�8�b�z��ZQ�����u�ſ���،e%1��OT�Y���o2�F��(� `����,���+��fu�k������$r�B��-4+�l�U����m���)X�1>�l���Ñt6��L2t29�p�5ؤ�`��:�C��+"�|WR�r���Y0�Oj��+��^�gׁ��5��G�:����/�5	mg܅��nB���k�	BW�'[;�Z�%���aT)8�%���CtDާ�zSrK�b��cqM}`�9�u-�*MM|&�:�1�"������d���f�5��ض�r�ї+���[kFGZ�1Bx�B�l�1�ƴ}��e�?�+�ݰ^ؕ��1x�Hy�i������O� wK^ߡ�D_�/"4�!��s�r2��ٕ7I=N���d���R,8z��KI;��=4]�B%��9���H�J�~~��?�!56灲�C9cw�*4�!�N�%¬��Ha<@�\�g�_�Z����O���}�q��q��-��T�Z�*�<��ŐE`v{�nݕ���d��GW����oW��*хaǵ�N�;�p�\�f3��s5��!���q�7�cˉ!����>��ck�DhB�K��w�
�FDr|J��j���8D�od�Q6����	�$_D-=-R(X=���w22���=R�=��k��Z_�*O����G���6��L��	 ����ct:��:�iCp���dI��������\�f�3�c�l��>VA|�W�6<�V��PF8M��8�NVwǲq�6��v�g�M�[+VK���U���3��׼�H�{џ��5������l������X�d���2���h
ňutQW�_�X���B{~�'�9�m����QM�0�nl7���*�	͞x�s��=Y���Wx��=��F�+3Z�����3�T̼�u�!��13c�	o�F-]������bv{ge�c������s:�j٩7�M�:���p+��5 xh���X5 �^;���3Zqǫ�#
9{ܢ
Q���
R�<F�da��,��:��b�c����y@�w�z�a�&�6$�B���1 $pm�&_�Z��x��L���T� o��來zXW+�$�R+��Ą�����Ze��v]��rqǬr[��YK�3���"�7�`��Ե�5�u��B�a$M{�M�<��ͷ�5�w�h��:)�4]�D���ee��	�r�q3lsa�+>��d;a�.��:aGx����ڿn�~��F��hL͡=]��ucm�Rn"r �r�]�'N�u͌�=��8�bK2��@�{s5�"���,*[]���`ׅ�r�4`«m�Ko"1C=[�2�.��[r6��{�x<.�K�U�LЖ�J�̍��Rd��z��#3�cq)Z��\1�/�X�7���b�vB8&6�^��>�Fӱ�9Wя|`P������PnaL� *�0o��o�m���c���툟�����(�m<��&L�	þ���w\c��V�����K�y:�<�m5�1���+���A���Xc�i�eС�u�҃���%�ǣ��$�*�`��~�f(�#�C�/�^�D1���S�0�3� �}� m�����@�f�^����A0��SJh4�iY:&�n�9���
/퇤�Y�e���%��tT�2�svy`�.��c�дb$��>_w	��tb'�7��h^#�EzB���|�-�r����1�֘�ޣ�OR�n�D���)��K�"B'�v!ls�ݓ�u4���d�)V�V�ǣB:z��/c	�5+)���g��x��V�@�f�>K�܀m+�֐��[I=T鄁T����ϟ�|��
��\ϻ�މ^�&��Ã=�v1N�uw�*LbB�k�/�E^S'��2@�q��1(07��%=�ݰ�:��>X��.�8�U-�C��s�AJ"�{�X�p�6��� m�|����K-gb��a��m&t�J��)m�W�\��8%���zz��r����nRo��q�"*עT�ˈ馌9z�S�y;8�8<�Y�йr)�{�[n|̽�#�ab�b�8�M��eU�A�M�'\�����ņ���2�w��U�آ�9+��aD�.EP�X	��:;	�~�1�/���)<��k0_'���}�2�Z�������K�����)�������kCK��C��c�U+��ޥ>�׆��7Fj#J���M����f6t���"�T�t�˭�tux/�t���	Ց�_�������λ��&MBySuc�y]kے�:q��m �E��6=^��d������τ�j<�nL�bh��H�
�����<�����}C�G2�)�L�|����đ���9t���.�"I8�C����&���I�ɋ�`�X�=�RJ2�5��3�a�>�;0�e��U>���p�mS�	5�1���XZ.�4�ʈ�pO��1��d+���^s�m�'�&y�ز���H����Ty�Jp1�C�����)��� zܱ��P����t&�3�>��֔XeD|:|ݔ���J�RP��8V&D3�##�z�mX�rUm9�Ϝ��1-EI�1�C����X���%yG.H�� ���{�nWn���e��/����ׇ�A���Q��S�{����;�tr[��+�NYԨX�H��>�M?��o{��	�P���� ���ڠЋA]�4���g0�_[¿E+z颶C7jb�7���*'��� �������٥�������Y�#B�i��'O�|��M�V3�i���*(3!�2k}�)\m�K�lk[�G�!)�M}S��(5Nc��i]lC2�������&��W�^���;����&�	<E>��:��T��A�*����l5b�B�l�:�W7�1��"3A๥�u����l<�O2���І����+7����Ĉ�u���5�-�=-�A:��.!��u�(�cn��.�\1mؤq�F�q���Rfr�6AE��-��t*Y�iМ��l�+l6�v2\��[�q� iNzԗ-�{_�u~���Z*>[]�5a�4i�5n�Q�\~e�hWjh��¿xdh_�/Z����P	��/Ɖ�#���R�w��Ӓ��b�1Ɉ��a�
�p�l��8����9!�9��>�:�c��C1ׯ]���`gʚ��"��;0��x�;$W�tR�y�4�Q$w���t9}�@���ٕ�߰jf�k�g�a��#���^��_>[��F���lx����`��2��g�ۇ�U��*����c=Y�0=�^	9�.=ĈPJU������®�w)�։��怄ln!\�)3�V-r2��\+N�:��P$�;AY�JFg�M��S��x�����18�ı�$�����ɪ d�8 eD�0|gaB��yT�I��e{?��_�����=�"6a��\���+����}|0���t,'�S�~�/Qe�m���]�۪[sבa�~dr���O��<r߽�Ȳ�>�� �`����}��2�mDkh���~I7}�B�Q�ԯ���ͣԤXM�6j�M�i� r1f�p�hL��!C�IŃ�����
�����V{p����
��3ؔGi�><̹��� ����IB��x�I�o��#X����0Jx�7����'�:K?�B;�j��A�g;�)�F��������ϰ�'Iz3����}@�4�����׿�t�{I��񟳫Q�y��,�䂱J����Ԙ�RwT�f�rOob��QX�N%�U{@�`����<`�]I��2�N><nj��|ΤM�cF�'k�5�[;q;fRe��f{|��I ����n����������*���ڳc��q�h5}b馻Q��6G,a��p6�Pu�������ݓ^�Ο����t0XCI�q�=��1+��:M*{�2~���F1_��tU��]��x -�3�B������/�#ǁ�1���_��/�E ��B�z[���P� }��4�M0��M� �k� 3ac#˥E�P*]Ĉ�2��y����+-�fw�9����KՆ��*^�K}"8�!�P�l��
��K��06�7��TA]��|�kÑ ����	��)�[��}��l���76�ZR������ܘl��x-�����#C�6<Ѩ�>oF�֫gn�A)�zCu�r&�����ӛ0�Q�-�_�{�~�4�c���leQ�}M�~���f���������)@�}��]�b�s�Zb����	�� ��'��v]WѲ�� .ˎ��T�2De�t�W��KO�-Y�%�%�j)�䌌Nd��u�吷����~�g� \�ظ6Z��)jï��rȕ>�\Mڙ��Yk�	����D�K_�a�b��s��	�j�'��A��^����`Ōs�Cj��5E�� ��±t��5���Z�vq��������c�Om+
{\�,�Nt���in��\.���Z_�5��ɼ�h����!�}�����MUs@�옢N� E�u?5<�^4)�	a{C���r�fۆ�'=:�`���P��g����&L�gB^L��U:�zW!v����'�C}�?���A��J��	��]jY�T��m���d�܌)������2��E��H��$�'2�a�{���S�n��ύ��>U�R��0�;5�s�������߼}Ì�9� ��3�}Z,��6$Ȉ��|��s�>@4xo�F1&3�0_op�bl���ZUI��p<����3:��Ɗ
���lP�D�D�q��^�uSHi��Wo��;F�A��sx���<��_xGxB��k��v�Ǚ��=�E35�X�ޕ����z�XP�LA�k}�V�O�{J���=̨rJ��gl��*��t�(P���nA�qP��0�CUW��9ƌ���{��R9G}=a�q���unFH���98�����w}�d��4�_=]=�2����<@SB���E/�ڷx�ɵ�[]R���ېv]v����L�q���0&+1���A[\��'��p��iN
O�o����r��zĂ!SNJK$���H���`�W���[�k��)��=D頽���H^�2�-�s�ު,��ֶ,�o��t��{(R���d8�y���Ƶ|@�Ǐ�B"F�k~�W>/a�ά�R�dV��8�(]�e��Ǩ+_������/o���U!�b�\��f,1k�
nJ BR9<ҧ�mil���X瞆�s�>�W���0���_%�Ъ�r�����3��")�m��KI��;�2�"���'G(.A��#��.
C/�քܥ�t<w��������P5M�A�6�zo'��}3^0Z_��1_GDk8�e�GtN��if�t]i��}�'ʩ�����/�}��6r{䥛p���u%{��Ӱ��UY-+NB`۝����UQ+/Y5�Z���Z��2�ݮ*xq�5#�y�^hت���X���2��W�&�Z�y�ox�!��v����5���׮��]K�^�h'lT�6��Bķ�i��T�")����M�H�S��Yaz�_놮KU����B�l}0�bd����B�	�f���V�-��'^b5�qwI!襙X��Ε�g=s�k�,{�S��z�[���rͽ�gU	���\����~��^��{@��Z�=���*Y��+L!�T؃��c��Y�{�����cVW-�f�qnd�Xco�&���'i��jM�.���n��j�ǡ�,��yq�ޮ6r�(H��h�&�ލ�G�_�i�b�����H�ݙ�EԪ]�5��"����%T2�q�M���z������
m��eÃ9ӓZv�8�t����&���usy��঄�����F�I���Sp�f�����V1x�8|P݅�)\Ւ6��w�[��{#Z~�漾�z*%j��.�v�[���񵤭���35ú�ق�R���Jq�7-}3`�t�ځ�\�t��i�QWM�P��a� �K�����s����P���?%��I�/��j)�-;X�cg���� nF�ͥ�^D��U�jI�t��X@���z�k��!@,ρ^�Quף4��^��w�Z��q�,O7߱��2�z�58�zc��`c5�S����6��c���V���y�K�֣�'��!JJ{a�X3��3�+JR�Q���`�RtY��JWxQ��N��+�%�0`�BA!�j����4#aHܰ׺t&|M��Mm6�9���o�{eK8�����H�#k���U��g6���� m����Y�`dT Ѡ�Ɖ��r��N�Hv	+�.�0DC�cm�G����K&���_u(̍��	���VZa���s�����i���F��;������&d�']��z'�jK\S��Rգ�2�J� w�b���u����l����1�E�4�qw��Zy��%]���	6v
%,,LP�@EjY ��10�I�!��=K���GKf�a#7�%Swݧ�HQ-�����mǬ�=Q���I#�n�����"z��qx�2���e'Ԥ�<Q	�tS�i�6[FveEO+�ioϏcn?~t�����d��D�A�B%ЧO_��a�M�K9��aR�)�|*|q>��ؒc��OѶ�ɒX��s9/l+m!od{�n�B�v�������#0�jm�Jhg�㮅��+ªM�"��$1gR����K:V�?��ڍ����\�BW.5-�-^nm��OQ�X�������n.R�=q&?��э��Hh�穵mOڜcF���xNvົ�����ۿ�����R����3����M�fBhP9�XC?'G���`D�Λ���rK5�C��W�H%�Na�=1��x���q��\�}�}��.��)�9<����q�?��S�IT�I����8�����nz2ؒ�?��*�g�ø�뷭�dc
��P�l����i�]��^�tRbǳBi�3W�νvA��3�Gj���+�?f���A�,�|�*�L��+6���o��Ǐqfн��@�rwX��O�o����B�>9��Ww��W<XBy͊%jpM�D��2i��j!fl�i�])�ҎA�B9n#�l~OO?��#a7V��F0��羼��h���)\3��{�q�o�0� ��̒�g5����{<�G���H#_p`}=��	�/aC�[%�1M�l;��)޲��/���{��rhڂ9I�b?/1PwK8$v\ԗlҚ!��&�i��ԏY���(
�KY���{`��봷��a���d����Mîʖ�\��V�l	y���W���:u�n[�ƞ�'�,,,���X�}�)�Uq8Ǉ�,s��
�r(�:�u��i�N�!"�>����k��s���-��C�ҕ�0���,oz�}-�3Q�E��Cū��nA��p�{��XCR��b����F5z������?V�|�󼮢8�#��My�В�T�o*9�qh�%wD%����5'i�S�szd��(YSB����EF�Ɋ`D(�8��}��ڋ�����s�D�<�Z�x�Y�䵊��u8*�஧ւ�aSe
X��OY�N&C/��R~�i�gYKE��i3��ν3��I�~��A��N#+�`�Ia��&P,���M����q�������GF�"̶Z#+���VTQ���G�Y
H���^�y���F�60��x]iB��׻Ĕ߻��5
Cʪ�D�j��!�Y�#�l�~'JVI�7��1�KP[���<#W���������o��ŉ/+hI��XL�t��6b�\�4t����c��׊�cnG�1�ɦh�ֱ��P�3���gY��kI��KiZư��O�Pr=t��w��`/�\b*u���#���ߑ����czh��6弸�I�����ׅ0Zz<��v�m����g�ٞ�����r����%qm>�Z�,>2��0Ɠ��q� ��Ac�:��=�;c<�*TI@�?�m߬�~�M�f��^�v��^�`�8�5ε���9���Y{/��Ү�w5b�sY�z���<*�b���[�ǟ��z�"�zͪh<@�8�=�S�e�ě�N;�"������?��a���a�;�aD_M{e��
�6Q߆�f���4W/K�'8yA�xf�H֝�vwxj)��T|��kˋ�Cdx�x��I�#�h=-����$ �~]���6چ�LT.y��s.>7Pki��D�q��_��jh��Rq��1����ky`�6�{I�ys���N���hq[mztWC#��	�j1�ֶR1���.��3CE���ġAQ��y���S��	�sa�9=Rc�>(qOOo��L�f?~�P �4���~G�-G��t�+� �])"���a�$��K�1�f��.R0�����2��tY-�]kҭn�>����f�ΰ�/�=e�=YC���Vw���Cd���,�eVCG%�b��ʲ�5��xhqb.�V����T�;(I|U��5�����5�H��}����+C�_m�7���k`�;"x�V�|�XF9Gw�)�,->$�,�f�o�G	�����9b�¡��c	�|U��S���^-���˼�K��c(����x8�oq�6	WG�dH��q��=O���z��z||�/�C@�����J�Ǝ�]7$�� i<�z�T�6!��f길����4�Xt��=��z6Y� O­����00��Pinު����^PP�0'�]B��oY�%3̤���E�n�B&����c���k,�^�Z��Y�$����Qk�6�#�,�<��3�2�IB��[���0Zg�p��B���+Ӧ�^���Շ]j�b\����g� T���k�S����A�|2��nJQ�ʸ����n��QJkJ@g�g����O?�P־��E��>3�Y��fJm�^pM-х'@�~N��	�^�>�d����)�	�Ɍk1Y~�	�Mb��Ҽ=-?����l ��d2���ރ���}n�Y׌�-v��r��ƈ���3�*�1&��F�^[�m2��	û£��.����V�?HإS�,�����L�����wޖ����:o�!����}���"�y��di�Ξ��Vb�U��a޻���r��`�@�� ���?G�{h�>1�zd���]�Z ��^��x�n��4}_uT�	;����E���)^�s��ㇻ��%�xT�G)s��Y���E}Oc��s���9�'Kԡ1�?���%�ЁHZخ
IH&$�{�p�N�����M��FB�㇏����0ce��RV;_�
�:NͿ���t����ߑ'�*�5��/(O�&.��p�o�9ޭݗ�����=���ZA�r�:��Ґ��o��rVޜ/�Z�s��EW,�\�	�c�ƒ:�Mh�ɕ�6����f6�{o�#TG���03���X��F�1���(��
�5�f�ZȞ
��v����Ε	���:T1c&�&��`L�AHla�۷s��πt?8ٝ`�&��%`��;ER��/��; \G�4���e��.�\{N䜺� =cy4���=�]z�+�9�i�S��m���N�y��킔Dl�%�Lȷ� �ê��;hY��@Fq���Y�c|�E�����0�c��6�3�Bz������X�S%V:���2��}��{6�#<�{ó�?�|�P"|�Cl<񙕵r-��4⡷�2��}��B��{iq��:�SjtP���5�o��j[_����rN�l��z�ޕ1[�#l�r.��������Ŕ��=���~wwx�q��'����x���#�P��z�2�M�BQpQ�hL'�Ug��<�B��i;Ԭ�zZcA�"c��}kw�[hBbB߽}��»��t��Cie({y��ǣ��Sb���M�	w&��V 'W�	�VVRʧ$�hۮ�ɐu��=6��G�D�19�!�+�Hʥ&=�Ge�Y6����Â���f�u%�<[Cʰq�|���U���v0�ȑ�=+߃�8�E��=Rx�y��{�A8Xo�W����ujwR!�{}���L����O����8�g��X��V?l�q�H�zdP�?���Q�����k�?��ShD�f~>��ꔴkڱ4�b(��~O��	`]l�H sqVc?����a蠫@���{ƨ�}�+��V�E�����/hW���q^����/���8�ZUB^8X�YFv���ܭ��!�dB���P~QW�x�t�ꙺ��y��e���!m�y�Ү���7w�BQ��]qQ�L�{�C�]w����>($:����\�.)/��z�  ��&O1cR�B~O^DܠXx��9{�Ж��*�r�
w�l� {]�����5�7�?!6F
�kٳ1Ó�Y��d�	H�Q�*���9������ڬ$�E���b����ř���¨[����`%v&y�6��J���UnpV{Q�$8���'ݲ	�)��~�k�
q9�)8w��2�N����~K��v��g��a���t�t�L���_g_xR�N� �����v��W9�N�{���{`n(�3nF�O��؝��� fIcڧ��0��,�(��+�`�Zv�#�e����X��?��f�����q�f�3�3ߑ%>������i�f
��?Ǿ��}"�D�lkuY�5��)����dT,bL6�nü��ߩd12����m��Օ�[\���F��:��v5�7$sg�^5��E�VZS))����Ә��-KK�r��+U@=#!�W���z-�c���z9�"�4h�PIὒ��4���B��؋naMD�#�Z��͜���d�����8�k��3�Φ�PH!VHY;�b�m1S�T)7O�h�ߛ����~�����4dy��/$����������Z[���(kiQY����R�����megWDȤcЛ"����4S#��@K��d�v�c:�sf;(d�g���l�'��2��g�y���-���xP��%��ı�������}�hG�Yx�U��^;�Z�h����k�����u%ik�P|���9X���~c���C�Q�a�/�0O"9�8�{�0��c.�9�H�e�d�����d
��1�NBkk�A�Ib;�CVu�*M^�0"�����݂�Z$(ݴ_��Uc�ڿ���L>w�W�'�/6���G��1�*FzgL�2��Ċ^ik�7�'a#!b�Oc-~fCi��O�4:7	��zQ�x��GvwׅІnƉ�T/�'�mVqǞ[xl!�<%^8ٵJ��#��m��@U8Zء�_Xs��.�$��9���P���T-˫y�5D��N9!��8�B��x<R!�� 9��@-�Q��St}_���ɿ��\��E�6eR�J�؜0��F������K�N�nqϵY�����5/|������x�sj�f���u|��5���e�D�w����i4�v����@���b��q��j���Oq_��M��C��4X���Eoj��uQ��U�*�8�����G��c��۞h(�ȉ���:>�:�w�Hɝ��#e�Ae��E�@�f(����c�DϹ?������f�2�j��5�
1/8T����w��S�Y���-��u����-����K��-Vi�=:~��ih��W�������Л���p�&���y%7[;�J����%��a��n���X|3� ��R4�d�����~|QS�Z�����91TׯW����s�1To��l�[f4ݣ��VٛqF�z�z���p�w��>�o]�\p���ȴN������K'�w�a�Z@�0�d���VE�k��(e<s�P��-	���͋�x���V����)�ww:�oJF�:֖	2�"���}�;��_�4������}z!��9	郕ɠ!KIɘ�@�n�K��8V\S�<��ZFp�m�y (P���a}�0�
P���%�޼y���ے���WәT*^E/��-�W�R���v5�
����}��뫅� �W�z����tN�c��Sf;��3�%�����n$�;�C������k�k�{���&��L�c.������pеrBY:��D;�C�V��&D��eD�m��W���_/A�����ʖ�`Z��*��*�6#�eUHKYdD�@C��>Mm���u�+�Iok؝H -�|~Sا~��I̺;\�����`�X�r�����&��zbe�[��I$n���}�~Nqwv�!���On����=�G�����8(�_���5��p�a]c����B:�*i��>�n}]��B>܍%+��\�y�4l�M�n\7��}�š�7��־"��2�5'���>�T\7�h�zt]I�Ͻ�|`����V��k�Z�,|6��'��M�$�Q'<�i'{	�6,����T��S�7���L�?D�Ǹ>�u>I��mЭ��OuŰם��a�Ē�6��Sm5�i�N8R��se�-H6�.�J\��~��F�4�/��U>�A�����Se֗�T/��.Uq|����-��M��Э�����j跮��qI��I^.�`D�ŜU��y(�2�\@Y�+׵��86\��
���w��w%���Q3�;�٬6.T_:��}Є�H��
z<��y�5Y(Ā{m*74+|_C+�!>�X��K&�w��,��?���\9c>�%n�Rf��sS��F�s��~T��u�pSGY������7�a��
D��|��h6�S�%^k�Ja���a����P~ؑ3�T_yF2��n���t�TU"4rR�x�twJ�-:lN��D,.8��Op38��4����*%Y�\����!��P�ߌ:�F�Q�#x������nL�SVS��û�ιޣU�U�����5
�
����[�}��4͆���s�퓟�g�|��_�� :*�(�0ts����_�Ҷ}�{ۻ��{�Ta��i�ڤ6���H=�mx�F&��щ���Qr�}X2W�]���
��#��+�z����2t)e-�::���E9/�f���9*4�gɎ�>��<%}B��A�L��75�,����YF��
guA��iO�A�Y�W�|*']�h�ؚ%`~jmsa������� ��;�+T�����9�g��V>m�|��b��8�aw�ʻ]�ۇ1��D����Z�Y��+���d{�~�^�|�q&����z�`!XFO�2�W�����6�{��-��ޅB?��9ڌ�Ӽ�(��B�������Ͽ�g�S����/�$�L��m"��ʪ�#hs���<������!5����4�U���������}����Qd�Iz�.p���汣ȷ��MZaH?~�{�>J�$���iG�:Q$�1��V˛�"j"�fM�n�l�"�)"��2eL����B��|*)������*���~3�b~�/]��@�62��o�Q��j@�ƃ$� cl2��%������	�i��IE���Eڈg�;��_�Jya��u���H���ޙ�y�5s$ZmQ�ՙT�w�QH��,u�m�UNp�0���txd�ґ$�X��G^,�"��Ncf��<��]��q������޾��)��8�y�#bv��1Fn[���"]$�ύ
Z7^k$���z�j*ma�p��:1Yϯ���/��j���F�I�R���nWF��~�1ĵt��*��=��c���YMԜ�v��5I�4RuC� ��/�	���6�a��7�F��)��b1����.��<[7�ks5GQ=%\h��}>O1O%u���P�����䔢��:-�;p��3���K�\{Q,��]��p�p���sx欻'��xg�VE3��X�6���6ڃ�L�]왧��,�=YJ�ɳ�����e�[��_/=U%�Zl���������x��/�&�d�GS���eҐJ��d|]Yq\�Rp����ʆWC�r����9�U�i�Tl�q�ֈ=�=�E��M��e�Kqݱ�'�+2�R[,dz��X���6��Ќ�$��Օ������y��uvJ����|���u4њ����Bi��<�`�5`�O\64A�w�}�k���hU=� F߮�e|R�MB���N�as`C��Q����HQ�]���]�&�p���ZU�`�1��?�&>�g��n�HCJ��S���zZG]�L`�a̟�(��nYy��T{3XcWxW'�Ipw���e����k�5�n�-4
6/��~,n׌�@[8��n0���Ѽ���
�u����
�ob>�*@	~;F%%�Z�+��9Ao5q���U?�i��H
�!���_%�qv�v6:pa=�W�D��^��0�7��M��F��>[���mkj�t�7���~�N��R/,7QgP]������2(��7�^i�&*=`�dH��Vf֭�]u�T����q-իY��^	��!i{�0�e�eRU�3�V�"f��>���'n�����!� 媝�	�:";YJB^x{)���1Ύ�P2l�1Tf��rC?�g!���^����ㅺit*}P�!9�s�5���}���w�v�T(p�:Ӭ����!�\.9���p��]s�q� ��7�i�g7o��!V��e��@0���t�>�)<��\���K��2m6.�==�VV������������%��8\�;y�(�dRjJ��Y��$�Ǻ���6�t<�dY�rH�կ)L��9(Y�5��͎B���X�=Z&2�B[2/,�\f̛!�%�NM�n��v���:��!��1�tJn*0 U�Θa{�X?�K}=�!7�X�O���Q8l����Ï�~{�~�}O������6�x�6��e�m`�#�?J#)����1����5��Ef0����'&ssm��x�F�='V3�^�	hэh�!/NrQI��Z��=/�f��Ъ��|P���^����F}��,��v��E��Z��}�vЬ�����[骖:lZ�R\�D�b$7����l���a^��Ù\�TP�{O"���Fԡ,<J��v�XpF��}��z��E`U���9[K���q���6'������1Ϣ�e��k���ȋl�#2W����ʹ��ʫ��BS��=zm�u�J#�����h��wKd7�9���v�xG���� ��͊"Q�:Q�XT��i�$���Ö�JY���eJA���1
�M�7�{o�YW!?�_ÈU����H6������oe���bL_��	����	�R1˯�Ε}�!ǂ��<����~�/.�Ph�Ev�"�-m'�x����R�^`�f�Ș����W���b��b=ٵ�3:3Ί�.�
��y�+%�$=�^ߑ=U�/�kp.gr-qW���*���7����}z̬1^�%f�p��-��3�M"�K�8�"�S<=j޹p\7���%��L���2����a{�����6�Wz��ֆ��k��:���i5<�Q�SЋU߫�Ԓ�|�W�i+�3A�E��������`�c�9�l�����>����O�&[,��gH!��̹IĦ�*�=Lqb�F�! ��	K����\�U�y�~��8.+u,Z/k`�I'�1��j����:8�cDyd��.�]qk&X���AM���\���쟖R����H1�����u�*�I4/�k��}��E�h����O[��!M�S	�>��6A�fX\���В�T���A�{S�c���w����MD�2��.�!I���(�L�أ�Ѳq������Xlͨ�.��B]S|����&o[؁Ę�Zt6�+�7����4�P��֌}��8��3gy� |�O���U0���!!C΁)1Q��_����5��ֵ��ŵ���j^�n ���TBh�؇i$1p�$��ưW�=���������d�kR�o���ZֱT&���nu:�UZO��7��."R��a,�#7-+�xHY��B�!�lr�#u��k�#P��ō��na셭[L�;Dh���Io�(�eY%k���a���vgH]�ϊ�Je��r�(
~H�&J;�vn�\9ن�nҫuG�1+j/�9j�`��ʁac�.�q���:d��G�H8_�fĝU��(~�}A��M�ԏ��H��K'>�K��4��[�%B%4Jzy�[U讐���6�
�*#nc\�F|_z-��Gͤ��15�w�����9�=��ѳ��5 �����5U4�4�$�fk�i�):!�$����r����7���:�U�*�1I�դ�X��1V����z�V(p���.H�Ŧ ������� ��a��AI
�(!�L���߃[D����̈́QU�9�ŐsU֬�6�nӖ������OJJE��kp�,�����IWܚ�Ʃ���ېP��@N��7{�[��x�������1�dp��þ
�8afm�0���0�4���:��'�4>5�7�^c�歹�Z#�i�v�ɚ��岦����mM�U�*�p�%Yh���-chЊ"�����P92��f��b��a�a�zkc����G8$��MO�X���{;q�\Uv}kJ��eۄ�k�˿iqӑ4ٞ�^s~�+�*K��06آ��yΌ��q(/R�������r��'3�>�������-����ʼ����b
���O9.�Y���3!o̵��� ���
[g��4��>�((���S�9������=�榲�$6�6��ņ�uͦ����M�
k�}�f����B�����ӳ����ن�&U��XYm��5��x��(7��m����e�{��1z�*.L-z_^�S�=�c,a�>�����-�uG^��G���a��Y����s��5e��_4M�5�/�#0Wu�}�Z�]D�Y�� ��a ����܊p��&�F�w�2!��U��Kx����"��K��Ѐ�r�H%C~n��-�w��.��G/�G���_�iM`k?��xm����I��O�8��!��poT;[������t�1�k-��r��Z��u��H�)��<���Q^@�1�q$dd�ƴZ[C*kFT<Hg����Zр�C���L�t�iڶ	���{@>.Ul�Y�L2lF|R��' �>�}�v�����Ơ���:�	pOI�B�ȫ0�����/�!�y��D_�� �qz��c<1ASQ���f�U_�et�Ч!�c�Ә��ء k�G&����>��q).�/K���,�c���5�QV�ZPG�:����F~b�?(+����6q=(���x��5u�2M'w�rҡ��+��vUC@γC�6YaX��Y�Х�5g*ս���Gi4{��	QYkRS��Z!8O�FF�]
�<ilUq���"��g�O쪬<���p��p?��
�~��pwR��wi0�,��3�C���ݜ{w�Ad�u�4t���w�0�|>}�|���I!�ݒ��}�P�/����C����QZ�\�47<`�?�jx��麉�(�����ZY8��>[)ª�!E2��lN�Wzk��4�ɬa�W�lW3�IN
��v��;��:1Z��=.c1�O�*7�2  ��IDAT�I	gݗ&𧁧R���0z��L�n�~�F&b�~�y��Lq�7�(#<��J|n&�_o�����2г��2c�
�8:�p1������#m���"w�4$�o;n�/#q\��W�6��7r#���7����a��&��s��N*��0�A�G�c�q>��g*he�ɍ=l���H��F��gaC*�bR`<�)�FU����K��u��ڷ�خ�l�:al�q�Y1�'������"�E�_�h������8�k@n��8�	�>fn�bCj���N�Q��"T�t����z��d�x�u�0����f3������%�l���Wp'[�=R�s��W�%�^��v�	7#���;��0>s@5�+����J��9h�]�����'�9�,d��x�7�\ϔ�<ǜv�}%���5Hc[�̚��^:���Yp\�U��;e����p�_+,z!�׺�嫇��L���X�<A����6 ��X�>�{�T��ǲ.�Di������.�ME��±�]vv�U��f�!嵆�����k5#NVc�7�r$���z|��)�����a
��XP��˓�b�E�^K�n1c�{��u� ��}u��3�]���<x�=�%����9�Ð���K�EU�̚��l<W��a�����Gf���aW�&Ɂ��i_�2ޘ����
^c�P!#{������Z���e��ƺ���1.wgRUz�{͙�Ƕ��,JN�of&��e�U�+ܕ��>���`����W����/�Z�<'��Φ..a��cp�:��p�d��N�b!e]skޏ�.������y��5+�&��!�,��4�:]]	y�r�i\�ɶ{>���Kn�=���u �e����x��揼��y-Z4K�ć�Ȋ���XkGE���ll��P&yRu�>��R��MM�&P�@-����%�� n��4�P��N�g5����"CX����)*�>�)л�6ɘY,�fL|���M"߁�x-tL�t���=�	o�M��Ħ���r�� �c�>�+�cx!.4zD7��\H�E�Y�(ocH�wFh4\�Rd�!L��.Խ�!�1��u�z�����ڷ�f�JқQ��\;Үkӎ�\U��v��2�ֶ� b��#�U�9z�	�(������g�����Â;�b3�@�5
\�f��$Ù��N�<6/��_Iȿ�nMB�cЋR%��	}?���2�Ӎ5���n'c7G�g])�7��KZY��4K�j�8�����XP�nUVњ���k��K�+��4���G���T�m]ˋ94+�V��=�$n&�����i�7~����V�Bm��\�m�c%21&E��wڤ�u(�X0>��p����<-�O$��J��p�0�.�>���`$��͒<| ���0�3U����3Uo0�j���-Z�N�\!�z���=x(/��<��>M��Cφ��m�>;�Ƴ��e���	u�}���t�/�ӀP��m�^���;k>y��Exw��`�v	�
�@&x>ǁ�1��^<
�| �T�㏯.D�zS[�0S��!�#������r�z����x�aLN�=喓�.�6�-eω�93��>I]ҫ�I�s��:xzO��|Pl��qx~�ؖ�Nʜ� �����:R��>��ub�>�(�8b�+�A]�1���cn����`�� Zܺ�D��8��p����n�7H�Z���C�2�uBX=�Z?/�j[o5#Gf��ݼ0��}��i���ڝ׉>�kC��.�I���t�e8ZCϵz�2�7Y�w������6�]z��q<����xNh+�P�D���M����sYB����~��w��N�H]�ۄAkQ��T�����$�"x�t��BW���g�� F��At���5�'�+�*x�#1��Mw�Tl�E^��ۉ�8,��f`lHC�3B�k�#0�녛���ND�c�$R���������5�cN�z�u���em<R&؍ɭ*8��HgM�B^�m'究�9D���1a���K�}QYbTN]��5W�o'�J(E�h��CtR����voHO1>-��:���u�"#�v��0ϠȆ�n�m��h��S��r�H��y�t]�'��J>;�p�s�*��-miCc��c=l�Ԩ��AX �]���M�T�6�V�F�=�Z�z��l�/��1}Ͱ�qgH�xC���^�0T~YU�	x�+y�_xy�:]]:��`]t��[Wr���d�dR���݉��?��p��JaF6h� B��s<%�p�x�G��'�YQj�!���Ώ�=��bL&a��5)~�^O�kU��#���Lp��V�N���C�8.FM��X2��w�׮zC�*f�F%]�V�1�!�7Dh�1�<ᥘ���v�hAa� ŵYQs8P��^na\�q`�3(��!�mܹϱ�V�à�n&.W�G�p����+�t�5�dmн�.��ޠ]_!�K꘰@c��\;'����Q�a���{q�8b�gŽ��(�̍{c�*qV�.�F�� X��Q"���+�;�$��f!�g/^%�=)�O�],�`��%J�[Ke�zTe�3�%�ۅ�~,�El���2��~{َ�1�BEX�E�gz��7X�_�<yįc���wn�0g��^�����%C�I����fVk&2�m;%ld�l� ��î���h<�������d5����$Gf{*�bC���",,������Z3��K����N����@G_�.n��|;���I��Jщ����F�je�L-�{E9����̯y����N�sgo�{���8�1����Y��e�����m��������>��>�����f]��gQM��^X�i_7@���j�m�U��Q*_�;�Z���z�!܋�7j�{�������"y����!g ګ�?)b}�U��UF�*/��!ͧ��ck�� ��wf�}�M��A /xʪ;+h�Lp�2܍�NcF
<���{W��۝Gk�7�eu+.��x�A�ג�9�@J7@�A3%�u�X�jX'[��c:E+6XZ�;Q�����i������a��g/�S/���H��:��S$�񸸙Ų�UF�AThg�����!�1,ǝ�k�>�D�.�%V�������$}�&�r���1AEC���^��mO�>�BC�������	RQBi���~�^���󅽚�e:T����)G���p�gV���h�02z�H�ﬤ彲
��ۭ�9�][�z��S���1����b<�+����G)���0�����3��팷�v�XA��Y����H��kF�U������|�����5��7�N��󚞰&�d�z�e�� �ˀ7!#����Z�G�o���yV�����A����+���pv�vM<�J��s�"��n1��@-��CN��t�#�9�!�58��Om0����)^I^x}������m�c��W��k�E9ؗkI�"OLV�=��������q�5���E�+�N�r'�p]�L_&m�M�מ���gx}�F�5�j��޴&���F����r����h=�fa�f2�aj�)D{�(�鶫� �Y�2UK?��^$~���e_�y�3܉eu5i��Xj�ƀ^N�u�>j5R���f�apCo��W�!g�ƀa"�}-w��mԻ�|�ӆB�deא���0���J�Y�����>/��tfy���G���8�ː� �'׻M5����}'�g%�9��Y��dF��65v1~�ޝ5�g9(�F)��{|��⌹�*Χ�$�u�<_v7p�x��y��� .wې�\���.�M�������0%v�V"kt*��s����	�(*p	�.����F3v�-:p+�0'�4��ܘD#�f�w�I��p3���d���J��Z������wԦR1<��lz푘����v�f^�$i���6��]1��#_Dљ�]����׼{W]`�P<��t�y��j-�"|Bx�zZ�/R,�K$b�:�4�ȋ<lx]WT��P2ۧ�9�Y�5u^�]�Xb[#MO�a�3�.S�z�3��� s�h��0 W�T-�#*�z_�W�9��Ė��]�A) �אF�L�ة��+\zivdf<!l��K8$B��s��Q�rc����A�O0����=1d��4�y{[��Q�6��F���O�Aw���k�S�����!t?��9C�Zq����R\�V�⫲Q7&�y�{��ʻx?�k5:��8�&�zTƿ��aF)��.����fCq3|��R}*r�Wş��M�Uӗ=�=>��A��<��	R�p�����U;I�y7��1�FQ�M<�.��E�o��#)L�[h�_Vvf���>t���/b�����x����TŚ��{�i�(��x�t��k/�s<�jц��%�A5�ә�w ��CX�*e&>� ^1W��7������>�cx�g��(]և���]%vL,D"T�cOh�TR�t��5BI&ov*S�%[��V��T6�G��e�ƭ�gΖ�4f�6F�=s����'�Y�/C-���2�偶~��t5z�����Pp�F��d�I�u��������t�U8��4(�nM���C6Y�L�9_��;�UO;������z䇳�I���p�7)�Tl��:�7+�SwQ���膕�]ʽ��S?a_��F���Y$���2]r��_�`տ�RMU�����(o�G����/,j���?iБO�l@^K���Z �;�N}M:����rH1P��xw�]���:�M֞��LIȹ��$���|��Yd9E��b�">�����,~d}�G1;B45]ݜkR��G[Dȕ���x>V�)７���b��=�n I�'͑5�"���`ڸ��Ŧ����M-����Ur�I��pL[��q�;�r�b�4qc�ߌ��1Rg6$��b�����SP ��p��=ZT`���N0�z:�	n�h��y>�R�O�t1�	ͦ��q��i�O���	/,�u.(Mb��C��!|2C�/��:i�f<�pΞ��f�]>)���N)�6r��F�z}h���+@��n6�2�h�=�;l�dwu�N9��e�[MB����f� q݄�R"؆�S��tn��?����ʃ����Q����i�����RHL��ӓ�C��;�	K�	�!۪��"I�w�G1��~�'�CD.�h��B�gPO�X-4R�����G	����	����"���v����e��������w�^)u��/G��x`��@� A^H��\a����L��6�n�D1q*�F�D�X�O?�l��47w�|'�?˦����W�1�O����<���c���D�"}�g�w��߉�0FT�	�J3�}��〷�G8��M�
�:��r�`�	L[33�����o�H�$l*]XP��Uįm������E�f�	��L�u�L���M;�L]�N ~�nM0��DA#b���u�p�G�������R;��AL��b��s�M����=xpk� ?j�#��@�g�0I;�v-1٦��'(M����8>������5���h��;��MP�Ă�����l�E�xB��T8@�1�t�1ȭ��� ������'�{Nx�x�>FӡF�����-BUE�#� )�V�|��`����X�f�8O�p/��E�v��E�?��Q����f�s���#�[6�ys�6�A[��zX誅�^$l������q�@)9����^��t�	��ɪ�h$�j�u�
�.EE�(��9Qm��kD(���$ޟ�fd&��y�}�q4Л- {��#���-Ռ*mP���Ml詡�OX���wj�*�Ǔ�}�7�hgޡ��!�z`�Vd��j�lE)��p���~�K��(�5��d_σOcJ�ٌ����L9?�{^+J{�@�Տ������bh R�!ve�1N��D�>H�V�fS'�a��@������{Vq��$e2]�q~�|@����ц��XDĔ�Af%;Zy��y�͹��S����0����Vv9_���٨�|���S�.vh%〳�h��X��ٜD������kRĢ�����*�1���_Ս���K�qz?٦"6<�y�6A�҃��$��ya ��/�]V�6��y�@̴��}Lc�������S=��ؘ��f�US���& e@�h�w��>]"2A�-ǑTC��;�T�HkN��nȉ���R�C�3�� u�徺�:9@P�� q_,�.��{M̸�&��5PKjw{T8��M��t��m3WǻEڂY�nL!�*�������4��l� Iќy��7T5��ڥB�ۃ!�Jb��!׀e�o��l+�ӎ���v��0
e�����͈�`b�&�s��m�vtϝK�3?�|��s���3	��I��#:��B�a������Ĕ��Jz��ɢt���"���1�M(��!�,�/<��c^��b��ĒyBk�t�dβ���Aw6v;��	������`��:Y�S�ObJӋ]�����&�d�K��ן�����S���ژ���)V+=�D�����?g�F/jk�dtb���"M������a��@*l��b��T�����^���$��"��Q}gI�����N)%���Κ8�I@�Y��p8�w�M�az�Q�խQt�c��p� RدJ���r�$63RM���?ޛ��^��?p��5v�EWn����j�. TgP�	 Nϴr�����{��G����L��v�Y͢�d�N�Y�`���\U�{��-L�nOL�H/�	�l�&R 3]WTD�C5����c!��9�4IHDW`���_d�P���v��+��F��+�p`b�p��o ��N���θ�"�r�NG��Y6w{ӟ.MDӽ�������1���ʖ���tϻ{�,�m>�bL+�7چ��Kz[�to�]���3�<��NW�%�!:����@#o��{t|âzѝ�b�fEυ��#5I��y����K����M�`�#�Ct,M#��#��^��f@2yb��\h�����>������ҭ�Rc��c;*���ӥ� �3�#�JOz�?H$ulHr�rI=/�*89��;�����K6�i&
;����N+���`b.յ&�6���$����c�V[�lni�F��U�3��ȇ�F�����{#R�>�J l�x����ղ��0�����>��0C%L�M���ت,���'A��xx��h�$�Ig2Khl�`��K[�\�`�X��b��;�H����`�)���yp~o�=�Nr���N�<A++)@�M�(N���lܠ�*u�:�K	?�QQ}�6�4i�dg�邩����q�1c�������DE�y襠_H��C�7xR�@�i��w�Nt�y�+<�q�l�OQO�{آO���N~���>��Ϭ�|O;��! d/,5�B������;�Ko�ҟ,,���p3bl0]s� r�úA���1��@,-���p�uK��Q�H��'"+�5�C�~����x! �� �TPp�Db7j�w��e2�ƙDŗ������͝�X��� &h�ϒ�v�f������4̃�3�w�.��Y�d���S��	�q416|ﶽln��dL�� ��rPR�x�ܝ'��
�̨�ci�10��mf�us�R�N��Dj��9	��n�!�rѵ�7�+L7��@�̷� ��3j\�$�#�ﶕf��$Q�g�Y�����A���&��<Y'"�#X�d�1���S#i脰D�Y=p�g�S�$�o��N����g��B�Ung;�@DW�_k�_��6�σ���Q��_�<?Γ����.�Ё�nK���+���-���L=BUEH�[��g�\���LR"!^%��.'����'`�`%K��l��< (DH1E{p���l���Z���C������Cc�m]�{�>�v>~���0b���y��㉁���^��~�r~��f�%���6ez��ٳ�a�OM��%ĒH&�*Q�?�gQ��ھ����q��^��&+�_ڕ�9 ۜ�4�-Ggc�Ϥ�BV����q�_$!���+Uԟt"�!�M�jQ.����%�#���!a�1]��qF5�6�z3��v`�k�:B��"po�6H��D�%��2.�δ�FOv�Z���Ү��a5�OD�)u�dJa�pg����A��ۻ�	~CWD�@�3V`]��i$�Q���mW^Bql�����cq>})��L�-bZ����m����\���30��&�,�H
S�[����Z��Z����a"��8�0��>K���,�9��I��"�6��_k��k`R�\6;k���_�RH����:U�c|PՅL|i�%�$Q	��3JC��E���ee�G���'�a���4 >�c ���]S����߲��������Ԣ;���CK�������G��>��PE�;�\b����}1��5�buJ;�̼��8�T3˞M��Nc淢Q��P[��BR��0�VJ�6U=v��{���;�U�sN
�����q�fR��@�����NU#�/p�ֶ4�I3�T�R3R��܏�90y�1l��"~_�B}�Y�ҍJu�>� ��������2Qz8��t�V<X����v�/�׿�e,�oe���������yM&�^�L�d�M�F�xc�s���ǐ��a�&~����?�aP}�m|�H��o��D���d��iLP�>2?Z��cvP�&z>�s×f�ȱ���j�1Y��)�4��J���8y�y)�'��09U��7@*�z�Ӿ��!��h���U-2��g_�g�᱓�|�ޚ��6�|r�q�vы6��v�,a���J9i�ĔΙ��+E��bzc���@�9(��E��e�̆�I�4��S|�_����,d-��s�4��)���7��6�w�X�o3r�xJ㛞��|ǌ�I�K��{�4p M Ou�8�1�飴����u��>������$�r�s���i^1���:���U���4�_S.�JҸĴ����Y'$x:<�%YDD��RP��C�LE�l��B�>�x����N�d�A�ؚbo�}���x&*P�����Ɠ~�4E�v;��0G�jV�Ad52�r�2	��0c����Ǌ�s����75�@.����}y2�h�@�6x�/�`��B���~����&��d�ai ��d���F��w�Q/]���i>ۀ��hFX��G��!`�ý->ӗLnx���b� ��C�`�8Ur��,��E���Vك�D�r� ���P��{�夻ޑ9��ޓ��BY�jͳD;��6�{C�v� G�D\���`�>!�g;�p`�ub�:�>��;�ۀ����?���,�,	��!�8��Tل Ф +tC���N��DTz6����Y��&S/D��
��#�ț&7&�V��}tqA��c���Kx���b9b<�=�;�s��2�����������+������7��������n
�����kRk�����:�m@s��g��2w�̂Xk,�lR1��X���4�.�C���k�8&������@�i@N�46�ݒIUadv�jT�>	Ŧ���[ R�)�l�=4΃��Wa]��h@�oTi2��|�C_b%���?�������d�fH�HR`
�~ro�$Y����N�{�@��&R��wTkzr�(�ɂ\P���Dk����f�sҡ�ƚ�q�?��lOY3�5��g\�}�ϗt��"%
�0.Ztx�8p2���m$Ŵ�DV�d����|�_��W������/�
:c�g�2֤n��nK�����E��%�Q���8�|0���Xǌwv6�x�00	^0��?g�|:�o���_�w�������˿��f%4[{����H:�kp~V7J�E�T��a�;a��t]�����������Xw7��v.%�Cx�g�G���D�a��˓��f�qi�>�c�'��c��_L���?D6~f��œ�������lS��ꙟ~�����?)�	��Ӏ�����d��!�5Ʈ؁N����{j=����L����%?�\w��RV$�������;Ğ��G ��)�^l� 
�جʕ"̏>!���s�8K�jb)�dS9�d#�'6|8�؎��`�,����G۔`�H��;3�O���v6ٸ� ���_��+�/<0�!t�GlQ�����~Q�Q_\xG��Iz0U��+�@Sv�=�D�运I�4r$�u:��|]Rt�d��Q�-��QWu ���z�=�m��U5Ei��k"�t�  Qw|1p�Y���NH�6�1�A�|�f\b&4��f;@
#y��Y5���y�,>�4� Ԭ�#�'�܉��l���!hOl���".��i6�G�;VU���H���B5h�9X-T5�c�7M�g�NyV+�k�8f_xM�B�ϼΎ-(�NO7�}I���0ie� %z�]6���I�@��8�;p�>����:/��_���;o1��͓�I��Z&�G���荥�F5$9ۙ��Dw5�AI�7�^{���vѢJ���6�&Ʊ���F�t�	��q�E�̏?~��b`K���[T�B�rG~��#V�"D�E��?�Ov@��+Qh8[��~�`"��fL�8�<�mV��T�`z;�h�x���T����ķ/jy@����r�q8ɑkƼn4��,V�yO=�us�ЊI	-(�-q	�UG7�9���.~4k�m�KbάS�v���"y��������es5���ޯ޽Z���'��HP��C:oa�%����u�׌��xSMy HY�F���6��M�H�3�%E�˃:���,Z]��d�9��$-��ӡ�<�F��0��t��j���*@��`����p�\�Rs��E���c�J��$���k0��{5OC�+*���2�L��A�����q��Y�|�b�����H̡Lq�,|-�`����9��a��;T�/���Z��/�#���� Rb�Hb��*%ܚ{��X�+@
%+��-H�;��x� �s�!��G�j)��)�����b$>�'9N�rT��M\V�E3aƈA˝�@Ҹ��:�Im@�n.�Fħ������.F���>�]�r�c���l�
}*]]rR��R :�;cGd/��^69� �Pdb(�C�^Z\`kQ���^bՍ�33;=�.����:M�w��%��gb�o����S�Md�l��ID!'�F��`�:{ c�"��p��l���A���ӳJ>����1�/"�Ѿ�I����xP�)b�)lE3��&��DU�aO[b�Ѣ����X�W�s
5M�󢙖l�8�=�)��4���X��zW,��уC�C�F�G�ݯ�2��
�{���I�ݵ���%H^:N�[��%�m��0Pk�ٞ1�ɲ`���w%](��Ү	�Ķ�?���	H�DS���^_n��i�#xF��5�� :���:ݜt`�H-anWjv��i����礉�h0?'_q	�&��O8�l ���|v�]N6�юBP��,�KR���I�N6��OWV�6Mi�Ae�P�	��=�l��s��T��޴��e��,��dfQE'�]a���qԲ���g�A��fa
$�a��~�P�O0���*���ō�Y�lN�Å���q�]�I��)x�t�>�`$�(n<��؎�8�	�뵣�������%���##���V�L�v�p0�}L|�Wo���G��Ǩ}�>�A�8T�)�8��/Zj����KU9J�x<&�fZD_}^p��njJxP��;5�'񝎕�VGě�:���Y�p}Qi���F�!8]`V7'a�f�[<�mgKE� @��&z�"��8���i�K�/�I/����?��z` i�@�T�VY ������*�hDF�zF\�:�0��p�M����/��FM��"�r3Q�C�= RZ��Z�7��&Ou2#}�.���}�4�E���}��.MZxM�6�f�� �}��U�<N�hd'����󠍃Y'���h@-�Ɔ�$�Q=���B����98��vPi ����P�EwP�m�0eL":����b�����ߋ>�2v����� �2~�|G������i�0`�Ht'8z3�lV�d��v�������>�g1�
36Iu��ީ`'A�{�1��,<�n�v�����m>�T��Jz�x��Ŭ�-�~.-���0-�P| �3Fc��и9��Ɠa��;����5� `�H��w��I7?�=�{β��>����c�K����`dAEj��n��T�����G��g&Jl�o�;oܹ�Ã�����K�5�g���EQ96����P�Z<;%v��p�޽#ϓ�ӓ=�7e֣��������W�k�s�c�{�Pi��l a)0VtO�`��ͭ�"Аѳg���8-��0��yhJ���x|D$����h!Gٍ�U.�;4�6��ܔ��!VgD�`�]jw��頣�����b�<�S��a�07���߶���I�x4w)M� ���X %���16%��A��0!�"Z�RЮ���;�0Ə�+��ݫ��� ��VB��ł��q�b������.�n���,�A
N!.^��9���;r�x�V�ް���{m�	�z�xt�P����2���A�)�Y�񁹀�kp}�`�e�i�g�*��G3yz�A�,=�����_�x���*WQ�M��{�s�K��E7�5�8���G�ͤ�a��t�S]5tܐ�I�I*���O���4��e��,������2���������.ҳ@�ZX<�3��S��:;Ȟu����j/���-?N;��ٛ�O �y�01�Dݎoo�}��3����,&b_�6�T
`�.>�K/����b����CmL�������7���?2zۼX\w��K)��qs0�z���n�����>]��Ϸ�p�9�c�C�Q� `U �:�
q=r�8R���&iy���f��˓�ؾ37[�xs M���Y�P���yۡN X��ac$J\���Y�Kp�D�mi~B��5�~D4s�� x]�m���3��Q��`���V����+洺_�^�A��1���$��ōߧ/�Wk�ȓ�v�&a K���*$��~a#��SA<Jv�k�F��@�w�6�0d1��A'� @s�l%(����_1�R�����،�榢��1xEę��.��4+\�	T1��,�����m�60!�~K@O#d�$�175v��E���Z���W��BM�ک�g��9h+�pe@
qv2���}���X9� J����m����\q)nV�fR�@����ޥ�|��w��codT�`%�h��D����|�86E	�#�BkǗb��.Ʒ������E�â�`Tb�#����s*�`�c��z���d�h1�Ɣ�L���	A8���Ul��^P;�/_�Q@�z��ȃY�\��$����,��!��
�z:����0��G�tF���>X�_�N��WY�m'�YRQcӊ7n�x�� �	�J�{���#]u�'�gT0߄��7�z�]���jw-3�&c�c0E�w ��U���->����1�g�A&�%��R�����#�g q	���oR�F��JF�HL�s�4v�X �6485,-./����	{/2J�	C�筒7���K�F)`�# �Q����y��(���Gm0L3g\�J-|�@st~��K�T_��
+��w���:NХ��c[ո�x�.7T1���<a�Օ�?��@�xP�T7һ}AR�����U�j����epOA�I��SO�x�,]ش�sK�/�K�L��|9ɤ�'��i�r�dM�~�n1�x�Hu�1 �F�|H�"e���n|(�4�(Vuou<6�b��bv�.CW�!a�d�M��MQ��)�M�͞),@�O�s�d�J�D|�L��I,��b *y��x��#˜��� 	fzL�R��}n�p�]�?�% ��bFJ%R�R�@:���
���A/�7ڀn_z�dg��g��Ydb�����h�;U;���ݬfA;�NS
�FY��~���/~�?��+���GZ��実��P�oi��@:���U�\���>�\�wI߉��Y�M(�m�)S��	#�;��Ǔ�$�g���D?��O&�}YI!���T��O����%fך9�!�.F(�B����Y�j�[�l�hN�Ic��J�c�w����)������-���=�:��'w' e�k@Sټl[�?���&h���ӞKm��zCq\p���1<c�}Ľ��~�J�{^:ލ��q�c��p���4�9��R�n1cά�#��P<�
�=��8ݬ,b�L��'�)��,|�s��_kI�4�󄟫���Y�O��U���f�O��u��%���C�p��MA_�m\��7��F-�{0K��-�k�X;�{�b�+i�t@Z�M<y�Ѭ#5"0�>��l�����M�\'飙]���JB����a��j��-�5dV��x~TFꢽ� ;P�T֙��6���K$]�6�T����5[(��"&ZŸ�5�~�����Yu�Q�쏏��{̉Gc�����|�r��8����=[�b�Q�j��w�����؁7�&�vԏ�YpƎ"�� ��<�� ��I�|��z�&���c0�i2#�,����p7/�ğ�`;C_6�`�gF*aѳ��pE���_@�����2�� _x���6	����IM mm�!+l 47r�-iL�X���:E{�9lP�l@��vf�.�6���9� Rv�P_�������N2�e3H�Z�Q<]���|�h��n�\s3�!0v0�l^_#�� ���1�K����m��r�����t��e=tQ�+y�נxiik3	��qE��Ů�t��~[?04�'1`����RQDs��¸z�o�P��)�E�A�;�)����n5��	���[�z��(��Dݥ�8X%Jt{��\5`�,�ߕSN�fp�]����,pu�0�q�*
\�ħ�a 5�ɨN��KtW]�Xۅj!l8��c|��P��Q;�S�2+r��&�btӒ4�=�F���oǞt�$��*�h��Z��fx66&i�h��Λ\B/0Ҿ��u��~���j1l��x�q���c@f[.���OyG��p�G�5?�6���%u��v�����:�(�8��I��̶�l�$e߮�)�9� ����`d`��?�M��?�_O��ȶ��>UDxi4�c4���<~j�����-3z��]L���sН���}n�g@��|����8K[b�۾\���zk����\���'�$�iy���F�;7��8j�SG��fZ����([ؚB�I�D-3���:�?�3�����~ڷ4n��|^scs�~�e�<�')s� �a�>³m��%@��v1������?��5ƣ� �;�6�Шv�<G`y�B��u�O����#�σ4J�����	PM䆈>U/���	�˨�	}�٢zȽ��#m�3�rq�)H>�Jl�Ew�C,��飃hX�OdnD?wSl������6a�Q���{��< �t	 G�>*��8~���׀�gI[ly�V!
���D�v��:>��l=#8�8G��{6�v8��\j�y�nF&J���>Z�M#+���0'��,���a3����e�O�v��O�B�6?;;�\�J��mH�~	DGc#��HGj�X�S��6�Jn��?�����z��
�T9����JC��C�C�]�4Jβ�sm�21��i`���ڄʎ������|�U�-���:wo�]��m�> �ȅhA�Q-�q����댯��Ɓ�/ ��wp� ��rI���#�����;b�}�Fuv�p1�����d�b�,�`��j�������g,L$�3��<������"_���J3�΁��AYx�u����9���^=c4�9��Ճ�W,��um���+`;b������ƿo�GW���st�oQ9G&8e6ډ���fC��Lm�����[e��uw�ͯ�(� hj1 �>���8`�q���<a8r�<�E;�o:���Z_qb:(�`��XyL�ܔ�8 �ʢ�2.�e��cp��!#�]���������[���^�7��V]�@K� f_n���f��e\�&k?5�<��,E�:�Ц(�F���rB����la���mV��\
*�Y{�~��9�=���u���Aԁ�sj�y���_�~��8v�9�}i�\&h>o����t �wW����<zǋ�Z�
]��qu����&Z\����G4�L`��7ճ��Y�C�Թ��E6n�S��29��G�L�g��[�lj��Jٷ~4p�pY���[6��MX�`�I�͒�n*���t��Z�.�M>7_�Y��)�VL�w�o�|o���;���M�r�Pl`��U!{g��/��&[far$o<a���:��n�� Ew�zYL��Zb1^�n�Fе��׎,�>7�M���C�ɀY���mp�*�9�����t'�M�jac)����@j��B�r�a^��{�ͦ���{��R�{eڞ�Zw��ڤ�\�^�EGd8콺�z�`~d�G�!��I�� �7��D��u����aB��قwDS+��0�C���=���H��%&�EK߼����E��:+��ƨw��%��#�z�#V&�R�F��<A���R�9�E|��@�؊۞zTz�u�{�-.}�4�5i���i� ������޿2�����?���>/��-%��[�D�$>|���x�� K�p�9�@4~�^�X�� ��~��=/1R��	P��ԘW���n��,V��ڱ�&W�e�4	�د��e'�Os��7�3�����B�� �Xw�`}��5�ՉP 
��&m>F�62п+�Cx���Y1�4���]ǅ`$*G���td=hG��*���f7^L�i�.���h�~׋ξ8h��Ş�aE)6?�kǎ�	@:�4�~�*+-�j��O�<W:0�ة��f�طE/��yv	Qn����c�ʌ���.vL�<ҭ�&��Pq�U�V�PeȮl��)r�]����:�m�������+��G_t�T�a�����K � �O=�0d��x��f�� @Sd��u�3S�9v</�qNxD�w�}89�Z,�՘���C�c���h1�e�fX����������c��Gq!b��m��<)���p��*�4��# ��x}�����$&Lы+��B8�4�
>?�G���q=gz�Y�a�g��+H�Vi��c�xr��^�Ϳ��u�7�=�>��H�JŁ؋j�M6��`%�;	"}��{��f@��M�=� 1�dKWA@	�3��������Rp�kB�[%��s�	2r�Qⳝ?_z6��7c^����v"Fs(�Ntט}DP���5��WQQ0��4L�֢��=O8 uy���(��2�̀�K(�wd��Ζ
C�<��;��#�����zJz6�����C�3�������{����T�h����TO%.��&�F�z�^%�Z7_xf�D����.�h~��K��o�|3������>��q��zv�0�0�{��`Z"C�i�-���F�>Yܥ����+��Ƀ�f�R��d[SH�%�GfJǼ�<3KH�Z�d��ß�WJ�z��w���q����Dk�;�Y�]����'{�l¸��߻���9=�JT�)�'2�N�+����#��O��,UMw|�,7�{��J�{zjY��0j���Z�=Yb�Z��܃чa��$���a�XI�P7��Lc�G@����ٛ��1�����=�^+��k�R��Ō�J�:�X)�P� �'����H@�Ӹ��'O���8���D�1aF!�Ii���D;�kb֠#��ti;�-I՛�UI*QA) d��B"�Ӑ�Vٍ�{��w��zz��u��@�TYp���|���l�{<��X_3X���V��߫���X�]7i�S��΀�Pnwţ����2��M�A�P�����5��{����j<�]I���f��F:n4��Z��g\1S�G�mAk:1}{P���%�r�'$Lц[��� �@���v�~iY&��0)�@����.�U/!|�>/Ɠ�DQ��3Ҹ����V�O7(1 &Gd�3-	�-1��{�u>ivH�t"���F�R��8�J�ܳ��q��גkt�c����i�>U�+a�K�+v�k��%�u���ˁU�rca�@o �z\�O���4�J��}��]-��:N6����ź���"��9�6Aه�	�� �c(y#�Лv��Ƅ����4k�i�s�]ڵ'�^fU��F�����,��A[1Vj��B�Ǖׁ��X���K����v�����Ez���d-�W>\���sK'��4��D=ᖯ��5�x�Tt�7�u�tI<��NbG���@��4�}�vO�y�Vg����f���w�ڷYڮc;#un���}j�X��t�ˮ�l��[��ݳg�ɍu��
q��@m4k=18.�\���hZ�3��?B?������G�GXD�8�:#�X�w����^�؊�x:!��,6��1�K���Z-�[̴�cvYҸ�����������i�<^�׈ۭ���6 �����QL2�WP��%���]�@�a�
s�'��c�3�=C �#91�⟔��:Ê��1"%?�<�n�,ј4��z�e5��~��R�ž�~e`K@܁p��Zߤ�lu=���
u�Ł�A� � ��'j�:�
�a8І���z,��"ѯcvj�;Ϣ�`�1�l��ll�(��w�^�8j���=��C2Cb��Ʃ�=�~�c���zO@
���ryL�Qױ�Ī�%ɓT�S�d�U�����n�x��e�[Ǿjמ�Q����.�xk��(�0v�Ζ��E$�.�tv}�'�c�׵��&J?�$���Ym�Ā����LE'*�}P5���L�bv�b"����-~
��q{�;� ����{��ؾ�^w������$���;�U�5�46i�,�8�����r����Gwǡw�M}�s<~  �Ծ����N\��?��-m���e�n��i����`fRa!�*`�3�$�* ��w|�R�踿]��ڬ�ݖ��xi�u�z�k�KJ�`�I/��]�"���¯��cA.�k�@P�Ϧ;�a���1n$��AT��z��/�čc��& ������6��?�	l�$�����ՁI�8��dկ��8S ���t�X���k��Q�/��ՏetO�W^�
~�\��R� r��p�;�����M�Sd%
r�?��N⥃@ѻ�ٔ�t�:@�j���)9���$�w*�����w��GZ�)]t�y���!1��ë9f��J	���i��֋G��(���F0��/ǵ�Ղ�t���6��E@
���
u,��D���nG���2I= �zH֚��`G��W�滭�A�����G�X���-���+������&�a9Xb0�=5q���s��ݐ&�ף�D��$J]G�@f���Q �jD�$��Z�����KA-h��ͬ�荙����=7�9�"aS��(��̀ H����w��{Q`����<����y�^_�$��5����<�wJ}��T~�����籗��A���D����@ʛ���H�Dן��~W�S���H�\�y�����z�����Lf�O/�k:�X�pr������\Dq�F�M�� U��� c��GRE8���@���&F�
M��h�7��x#�L�ņ�
L���<�~19!�d��.� ީ�����E�L@��^�d���c�Z�8���z��I�d�#��X8B-��YGRJ�D=,<���X�b���z����fOe�Q�ՍVC¹j`2}� �"q����[�:���GuE\��~�>@����EşW wI�t]^��w��L B*�y��Ӂ��Yy�n@���̋@�\��l_w[�1�sSQ��V�|cA'��E6�қ��j^R�Fi>�|5̺6fY!77&j��A�93N����{�\*MǬw�k�� ��%�k�'W��m�ړ�i��A�=�O
�&*�F�y���q����9�l	/�K����$�y�Ǐ�[J#��%1恋��5�:Mc ��	"��{P�%P��f��8�4�;"�SL?�+w6����#�žb��|�s�U���D�����`:YlQ���gi$�޸�۴��1�B��H�U`�ԯ�l�+���Jg���;L"�-�0$�1�[��X�L����b�M��z��&���[��ӳ�T9��&P��r\���z@���V_�{�"8�@��'�qDǺXc��e��&��H����War�@��� !8�v��=�dI���J��θ덉n̠Ӌλ�&�_g�k��n���!�C���ȕe�Y�����u�n�-y|q;�l��B;�{�U��I�##!@s����m "sd0��@��� ��wg�Kki�d�j��=ð2<'3͉��-ň�4����� g:���6�To����9���� ���w]b�׋�y��J���4b֋�?Iu�?��q.�nG|Y�-&��ᦟ8���T��� ]2#��DE��Å�1�
�$����Ã2Le#�s1�9<^ǲ-J�j�U�x�PxS��?�:%�E�f�\R6W�y"�.�1��!�v�Y�l~�Pl��r1.��Z����Z۱�g�N�h�L��̝�.���'�-W���ا���%u>(q1�V��R���z.�_ �f�O%"[X��h���=0�"a�4#]`؜><���c�3�k̮���q(�ބ�e��9��Iw�)��o���yw���6�y&�N�q؃`d�>���3�,��`M$M�����溢$;җ�+.��a��\���j��P�,VF�e�r��b��]��� D��+����})MN2z�@�L�&�(�3��qw���5Ճ� ��l�L>�-�\LV�fj;>-KbS�H�)�|�$Q(2�Rkc��}n�fD4r E[���_�瘞���Q*��+�e[�<�P=�L�@T+�+��:�D9�ˮY[b<q0�����T�P��4]"j�[mA�(a�]�O���6-���9l�A[v�W�i%K}ܺM�#�Y��e�HS�ϓ� �Ya�6��Z<冲}�]=k�.�Z�y��{�N���zk�	猖����_��Q�����@�AȄ�� ��, �[��f����3#%�R)��d� Z#�@4l��!U�A�QM��"�I��+��O����i�ACT*Z�Y_�#�:IY����I��	��C�ω�,Et��;-��Er�].�' ,>9�~�`oL�)�X��Ƭ���a��<Yu��P��E�n�����X��u_��O`�e�p��P�q6	f���o�!QcM9�b�Lm�Z�#%HJ��O\� ��,1�/��,��������3�-6��o	�`5���/X'MX	QD�^�u���D )�#�}
�al��l���%Ϣ��O�cٓho@�hb=�*�.������\��V��CHR�D�k��� ҶI4w�w�$RM����ig[k���XN�ٮ2'g�)�Ӳ��^����C#ӫ9\c�Ne�Ff�cq�ꢀ�M�&}�j��PƋ[1��vI��N�\�,�ҕY7���tSU��X�hX��)���D�����%�K�>R��AU�TQ/	=E3��7@}�����4^��|�[��b���#���R�=oLUＨW� ~<&��ę���C�D]�xR�tڝ��}Y��e`�����y��hC-d�� 1O�n9�����íD�� F[�I\\&U#�r`.�zSm_��U+.L�"�F�ܬo���ͱp�İ0$S�%L�D)t�5��`�S�X���cR�DMn���!IB�~��lRDS1:����^�����hX�T�p�?�	��}���$u��!)غ�[�Y�i�� :Ƈ��Gg�� 13�V2H�N�$�[��{� �����������:Lk�%6�����b ��W̱�iE��B�� �����b6�����PxH1��yt�x��v13���Qi�@�:/��Q�hZ�n�J-L�I]úF S�����/G�E�A�3��I�5\["�-@��y֗�-�D����$n6���	��eu���Ԣ1xf��z�UkW<X|6[dL�V)��ժo&�-�d�U��-v���F�8s�%�=��F��G��*�%���*�k�:0�ثfۍ�2(.�G�D|X0���[1[k:�k3Ь��o�[�=.����54o�s_
�Az�QY�6W� ��gS�����wi�$oDD�.v0?ސ:�����+|d����a�j�{�� ��8�}r�E�4��^/j�L"��%���/�'�us�k0c[����g���7d�ۊ�c�� �n���߾��u��Պ�f�Ƌ�YpR)lV0���G��X� ]M�����1�礛r�7��MXg�����<��l�����tL�~dӽC�	�`���S�q!jz_V�2[lԄ�(ڇi�7���']�b��^Y��]{��m����e������!����r�������h�5 �HZ|�;���6f�����]�&���T�V~ڝ����Y#=ZyY�]�\�nq�,#�I)L���Z&�EAG����{\J�Ȅ��x)iPz&��1e� 5L��@�Ƞ�46�_����\���dS;E��8�4�e�\Nr��J"0�����t ���URq����:Fvz���Wm}��:�Nn�ld�G�T�,.t�^ց^��e�ը?�S]�	W���2.�+�ƀ+J��i�������x~Cɾ���� �]+7�Y��*&�[]�Ǵ�����y۽���>��llPE(I���E�O� ;���c9��me��u����{#�2�A��\�0�*@�mg������ы��`���Nt6����������|d`���Ed��>���'����M�>W�zrd��ű�b`�6�V��'2u������?XT��W�M,Z79҄ �>�QW��ޞE��>���`���T/�Q�������zz1 7�H�:��g�VYad����ԏ �43��N���ʀ�:AxF���(����4ϦUK��U��{�Ć\ש�Oc$���<��1�od
s�RM5�&ߏ6�����f�@��Ԇ �o��A#��@*���q��|���1� �EK
��-�y ���(��; S(Nc�SmkvK�n�����Q�/�l|'�����ėnW+��im6.��4���`1Z�ƛ���A�c|R��T'�<�dc)l����n��iq��:�@X���P	�z\�՘��@��<����]j� ���x��7��6ߕbv�[`Z��4n����� �������B�v4XE3��U����/
����˛ �ag@V�Ӏ�UW�����u�Ii�4c)����  �:#�v؉*�>`��� sR�;���rf;�<2�H�Oq?�St�g��/�l�yE�u�Ha'�]�ە��@8�A�+����T�6"Ոm��t�� @��B�ӹ/w4f5B?_�1/D`��Ls���ؙ�$���%�cs��ݣ�8%��uc���7K�	y<_�9�b���S���Uey^@{}9�ߵ�ї�Qo,�k��H����:vyK�+�����;�� #���&������.1ŨK�p�Y&���h���ĺ'�𬖐wLT�o�b��V�,�U��T�1/����B��9`:n&
�"}+a7ٙJf��ibjʔh#��o� �	��j�� >&V��쎬M�:B��nf�AT&8;�t@:�xA������6Q]j�w��"+���f��= Zy�ٟ�E6�̘~¸FJ����!���"��<KEI��(lg6��e��s#Oʑ(�/�ž��
�®r�Ko��Q�˥^�^w�c��fyU`�Xn�o9N�n2�Ae"����81bg�q�)�>e�@���0U���j�}A4&$f�TS�a�)Q��2أN�X®�PO�]�5�X��P%��e`(X �b���V�uf�b����|�LX�KƆ��nu5.�8H}�o(er�R��#�Ob��X�:���TR��I��u��@h����m۸7Ɵ��5M�M��a�
��7L2�Y��q�S
j2k̂$��ɫ�O$�la��'�.H�@���N�dq���{����*���Z�%��:�s���� J�w)�k�����9XI�h��?��,����?��(�BdW&�rT�P�r`�A �>�����d�Ǧ6���c�4`	�=qd;U�������� 5�,l<�ۢ_6f�hx�M `�>���|��vF���:�za2��c�X̠�50����2�%�����\㇊�Ip�R�t%co��Ԋ��(�`�+-� ��5^�j�ƇHҐ;v`�1�U =���(R��u�y"��S�,��?���3�ϋ}���������ؽ A\��_���k�\�
��ʭL5�����@ �nN����d�T"�؆��ŀ�v�K ����j��*D@et�R����'?�_�7nb�ڊ:h���"���pl`^�:烲���H���ǉm�6���!p6
{ƽ&-l�F��2+U��vuKd�`�	#��kc*3�n��(W��J�Kmb&şL�N5`��
�K��}3� ��x��vaV��AC1�h}L+b�2�U���?��0t��&��w�@z0 �t���M���S�o*�c��+���e�A$oۃ+�f�`��S�	�M���a �F�N��H1�lb5	P]<�;�;N��TU̫�6���,�ؓw0
gw��>&�'�O��M��&����!���3�ƌ�:#Z�И�k�9�j�r���#����� ��<�A6�p�b���-���Y�5��/� 3)��'��<�b{I�6��b�'툷6Y];J��e�8��D�L� x؍g�O5�otD7!Q:���&��iB恽Z��Bd0�T���X�����p��e��\�o��=�>k�^
�Evn���~�i'�5�+N ɂs"��l`���&N�Ln�C��a����KFk �EA�Z���sR-2IO�+ƾ[��վ����@|��p�D0ƄO}�l��q�giy	}+���4Gq
����)�+x氐�f��7�L��+T��=k��V�k��՚z��e��"{�u�̲��H�U�8��L��b26��,E/Z�V[�J�����ԑ-0NЩ.���Ǵ�c�%3B��'�fl����03�5Vߔ�,,�_ї�ɼ�\8�S�l�g��藍e��ĈV{��1���S.`��F
�oԸ�	���)����ph]��jjR��dr��6r�2~կ�� ج�NMM�Ǩ�k/>ѐ�'郓虡th��Y����IT"�X�诀�/���К�?M��6\+?j�#���t 9U�]����t2���
�з�}b?B��ؖY_�8~�e��q��X���c'�Sx�� ���b�?�+z�a��N�-/�0&�{���et����0�}��L5�T|۾�%N�x���;̓%�����0i�S�Q��5�
(u;Ϩ�I�l��#�+�D�]��᢭!�X��~�X�|���Iеgd@ ]�',�<�m�c�� ��l�W�"��i��Vq0qp.�7�?�6D���z��@���@�%��+�F�"i�>m?�G�_,�����-[H��KLxE ���Z�z��-�[��7%����1O����P�`lIa�Lv���N-ww��,�R����ׯ�ą��W[���ͯUl��"��D�R�z�+�bA�U3Q7R9\q�����}�L�����<|�\����f��HW���x\>�7�{���l���C�� |����J	&,KhG0\�o������ٕ��]]d�DSK' ��#z�?q4�q����8�}�
ڴ��-�}����T�@�����#��@�4�0����{���C{� ���^PD�*����YE� SW[#�0* }�Ol��X�����+���%I ��^kT���c_����o�=h�t�ۀ������g���0w�v:\a��%��k}�������,�j��>�����c���3w�<O���1�P_}&��$�̫���&b�1��I<� P�h�x�C����tA&H`B�sLA����YU��HP`Z��?/"�;����N��5V�� 5�ݭ�z���7K�4����Q�yށ}d��N��S�d���G�Q,:vXd�y�C��Tb��G]�+�j��><׼���]�د�K�E���<��B���]�b�#���l�6A�4" oQ����Z�e����b
��d�kx�4XpL�7�eyk�t�p�P�=�+>�@���vn���f:���fP���ÖQ�<^d��մ#�$���WRl�����)D{����� �N�m� �c�;�7��6y�LFś�~.`���e�wtA�!P�?c~(L�D�;��3]�)�Tk���qn���^E�k��zn������:+Ee�s��|X�f� ���\�@�XT&3iS)NU`�H�J�H5��=�>�F	�撴�V~	��\^�/)Ww�m�^x��Mt��^�(&2V�e�tc��`7�)<(Z������������O���w��w���NK)i Krٙ���Np��뒮�SC��%@Z'oӵN��1j8�L�PJ�ګAl�Bװ�������9���q�Q��b��%�R�^�@�n�T䋦�fſ�N�[��Q�C���8��G������
^�>�);���z�0I�w�IF���<��H�X��bt�S�_}��I�J�f�E�ʡ��|`�|�Y6ը�Ѽi�6��Dc6Q�]|G;��ｱ�"�5���S]���`�z������U��:�Jla����u�8�`,����0#}|(�������Ǐ��Ǐ�ݻ�I�e�����������K��c1�������+�aw�e*�:�N�
p�w��Y��ű �r�x�I�V`�~�8^��o%V��t<�R"��!b�G�Hծ�WaK�Lo��u6�T̳��#�aU��b�<���h�;뱂�X�}m�\`�Ffi�	��~o�
V@Ҥ�e,��YNl
��#WŝzyAO:2}ZaF�!��8Oc��^����~D�������W�P�^PFL�V���7G�h1��Y,y|x(���˗/Ogf�^^gf�ylt�,����O�/�RtM;b�"��z쇴���`�
��<1�Q�h�k�.�'w���'��(�[
�1vއ+��w�5�:�(�Bġ=��i�k`¡��1�L`���Ġ����N���FuҧWs���.s��գC�FO1���� #���r�:˱Ks@B?3`�&U��͋n��1��ԶK5]���:��Z�,/2���)����3�bX�$�����	�T,B������G����):��L��ȞŃ���Y{80�i ܟ���i.O����O˗ϟίϞ�ޔ��]<?
�X�,��'Ì҆{2��^����Ϲ�����X�1 jJz�I�8�DxԸ��˦��L�.Պ?���_��^�Yw�[nۦ����5np��s`N�g��g#��pa2���>#op�+(�4�LWq����S��@9���p=[?�^Dc ,R��u��6�%����Z�l�Â3M4�F�H������� ���F�`�e�
�-�$��N�>ߟ����~}W���{��ޝ����G֓�K0���~��P$I�0�|y�R��d))�W��כ�󺲏+|/�o���{�V"�����h��8���,�mɥb|5)�/��?�{<�<=}.��3f������fD�w���R2�-=�	�{������<aխ��I�`��f�Sm���(����	ȑޡ'Gc�kѵ��#�lb�ˑ��eA8G@Y'��*7R޴��tV@�/��������]��xJu^�O����h�0J�Ԇ��U��2�F$��O��X8�`7�R��#�UG�<��N����yޗ����u�O�EtQћDq��Uo kzS��s�������Z�?��p~��|�����/?���3�~�V/�Q��Њ1fi5�VVa̼���o��Q��������K��o��,�k�Ȫ���Y"�F�b���&����(b�r�O,��i�I�X��)��3�O�M٤��,�Va�[�E��h�.��/v���-I�n�@�������̐S��g��S���߼�X�z���&5nЛF�Sm���ꗻ4��=,��h8N[z��[c�@Pk�Zg��q1k`c��u���j��f�H���Kðͼ��N{�K�Ekf�:>H%����s��Z�:#o��={}o�ڀ�Pbx~=0����Qz����N�Tv��|��
 �ޑ�+$�j��<�\h~��j|��k:ˈ�[���ec�]J�\^��{���o�� S�e��w�Ow�1	��)J���:����|����.���S��"�ܰ���N�� ;�u�.Fg�p)����v	�TL��v+�l�٣{q�j�|�x�iK
Њ9]-�V]q��L�A1��6 ʾ�׏�t����5�P8���|�M��A��Z#�@kw�k�n��ʶ��l��`-)[h�}!�$����|�Usvc��Z����#% ���}9�+%&J/��>6~�9B^bi��ؑ�r���Xl��~h�������l�I�<c�]a�:Rp�x��� �u�V���Δ̡ļ��@���L�x� �������,w
������Z�����~k[/�݋ķI1���
�:3Z����HV�������|�IC���	�����N����w��T���Z'�t�:#��$���'	\��K��Teӎ��8]Ms��?w!^,L���ј�TY����g�d&����H�g})��~��'��f�ة~Y^[n�Pz{��u"�Ӈ�0��ꀯ�.΋sR$t����=' ���Z#�"|�E[ د�# �x��k�6��{)��k�0#k��1�G���V�&����x��u׀���F=�n#�됨��V��B��g)=
6�!c�9�(��Fm��ȬPu�v�c��CH �uw��DJ������3�|�� �މh��	,[��&n������oqߦ|���\u]��}�7�P�B�E�I*�k8����l���RR��_�<��3r��2�B+\���GߍV�[����-�A^V[Sd�B��1C@�Y;-e��J��6Ľz�X�EQ�J���K�i�[UȥF>ېv��ԙ=��iz�ݘ�z뮻3�]
�s�7��N���C\:����3x�;��;O�H2�g�H��O��MS� �T"��#L�ޢ|�����Xh�K�� �*Q �>��|>2���� �"6�<g���~sV;�@�g�#��E�%ߡ�*e�X�ԼH_W;��?c�|��n�&{�v��o}�pG{5�1�zQQ3���R%��^� �[VD�0稟�o�wN,rw���{��#g�{�L�4��K6��<��bT�������1�����R�����,�53��A�v#[s���u�5�ì 9'Pt��3��4�]�C �E:�G��V������w�'��/w^���o����/T���˟�߷c����;���}c�^����©�34�3Q~�,T����<��T=��0�ċ/�a�ɞ7 ^�-��O�{<�KKl�?c��i���7��q���� 4~@�o�m�2�f`�� �[��-0uf}2P�	�n�'>���K�����������Z6�c�<������T��U~�v�V|��?�{�����֗�At�3K"<1�;}'%'���,�+y�4��j��1����#�n��T���M�����	���Yd�K��a��3R���4�޳��n��16͠��1��x���{D����l�l�վ��=ՠ)\���=�}[䄅�$\��.��k�������H8�N4~{N (^ Q}�wO˹t{���1��XLZ۲�.V6J�& �=Տ箚�ӡ�q�o�b�@��z�a+m�	w�;�xg���d��d��V��#����H�#'0���F����H{��K�������v�\���u�� ��A�#�@��WL���'j�d��\_���(��u"�@U�J<у��O���\����~z{f�?o�v�|3)�w鴿r���� �3���﻿�Ʊo��62hs	�_�=�*��墊�jn�<~�K"�k7��5{���F�=,���^�ȼ�`�A�Z{8����&_O��A��"D�:��l�����u�K��u�z����/��y�����>�Tx"��S���h!M٫j��� �ob;^�[K��������M��q� ��j??w��wT�Ћԕ��3�H��||�z^�W]�o�	\���ֹ[�M��=HJ�z�Ku�ާ=���}�����+�{%`(������:������F�>L[ɠ�״#C�YO���t���9&RHF G7��z�	Yn�i������EZֺ{�K�z�x���^\d2��(o�#�I�������*����3"�g`����,Ë����Q�)c���x�q��^b��:���G�O�;C���D��'���e�u�{ĝ펯�}�����땍��� ��D��L]�i�_���@sq�]�Z�n{|������|o5z3@}��U���������o�p5��7A!�d}j�\�7��n�6CJ�g��x��bq�5p0�k�߻�rvy���;g�%��5F���"����rS�D��o�!�k"�"e ����o~ΘU�]"1��=�\��1�AB�T]�/��$�u�XVe�}���ۄb\��u{��}�gQ*_��rc҇W �,]��ۖ8���+5 B3��'��JT���ZK�����B/ׁ����
��ˠX��=�o��}��^�V��@Ò]��Y�1d���ϫ�
�� ��g�H�I�C����8� h ����='��ߚ_��s��,�Jo��u�TzpM?��A�ʛ��<<������Zf�ߦ	up�]� �����AͿ䚦9�_G'�駺ү޸!�^˝�ҳG*����.�eN�����'q,�.�{f	�g�<�Rz��ۗ�E`�s�͞�F��R�6v�T/q�o]��"_���B�\���ϼ'��uz�:g���w����c���۸P�EY�l|��`4n���6	��������iF}�gp���fX_���2j�q=]�hAڈ�N�f�a]�K�w/·
����}����W�0�m����Ok��{����W��c�ϗ:+�JI߁h\���ێ �����~����p�����D�M����z\�m� �r�+k=P��&q� ��@�ǟ�Hl׳�_f�9�m����X���IW,7��zU��t�[�_��O�T�	���O�p�j_�\Z�V�Ǥ��=}���ce �<� r/�0�sV �1�S� �{���2������ė�P�$�&Ӫ�~�o�|Q�(k@o������r=��r\'�����`�kF�ϱ��
[�' ��ͨ��/���Q�f�Ժ���V��W*6�q߃���������!T:Nw�mF�z�� ��ҭI���\,}燿�֛���ј	�uF׺��c����=z�A�ZUl���>��|�&ܲ#	�zl�s�3�?sz����F�^���沺�Yʛڑ�W��i���h��a�D[�~�I�NI���[�= ��u�{��=���5@��O�֒/��>���4Ɇk��R�Y}��ڼ.���Ձ��reQ26�֮�~��MKR��K,4g0�`�\�n���F�a��M)�㵀���b�z��&�%]��ѹ�(��nD#���D�c��o�绦'��]���r��Q�~���r�,�>D���y�b���a��s���mW4�c`Y�S��8\3D̉m"я�����w��,�{��@Q����`�-7� ��g�w�:]�k���(~T�D����G �U����ts���{�z���A��-&A~��Kf�u%~�Qu�;�() �����z[㠻1���}r��15�s���y_b�#]�7�7*��X��~"���1����)~�i+끴������%&�븆�&[
`�тF����q}����͆�����:G�%���~�ZL�1�(��l��ؾ�WcQ�(4�Z%�t��CJn���>����%����F��1@Z�j$�c�[4c�r�m�}$��Rz=��ރ�t�E�@o����&V̷�ib)�Z�DCtY��c_���6� \W5��y4n�.l�wP�c����7���55K�#�R-6���V�k�s4����6 E��@j�����ط�K��Z�2�`�uBB��^��y�v?���R��b/�m�h'�]e�%��w�5V~~�
H��z�^�.��{�]�ޗ�u&�������}��6��ۺ�������Wm!��|����s*������o,#M�'��M��p� �W�8�J)����N"�%�-��u�թg�=H^S�X�ݿ\&X�@�/���ҳ_k��A���n;�����.U+�9j��%]�
���$���ܷ�* ��k��7�r�0�y>��\�<��ّ����"��8�4y�ёX�2��k�t�[����І[��t���փ���.�hz���n-ݲ���2�����]��Z}0�os�	@M��u��Kt���/��k��O7��6����"�����2���;h+Q�5�e�`�n)�c�΋okp���V�[@t��8!	�/r��~�U�Ri|Ǜ'�K����)�a�]��7n���@�I��zᘗ ׭j�-"r���@���ko�t�6y_x�׀ӵN�N׮���^[^�[z�j�ƃ���\��}3Ϧ�����'2�[ڧgz(/j�v���z����A�&���x}Em��    IEND�B`�PK
     mdZ��� �� /   images/7b19d218-2217-455d-9a43-b73a208c2c5c.png�PNG

   IHDR   d  �   9s8�  0�iCCPICC Profile  x��||eE���6�ѫt�q�"�����ٰD�ݐd�b	!��l#[`a�.  m�"M�(E�HS�. � MP����ܙ;�w�������w��L;s���;�%ɾc�,�3��$s�-�<��Ǟ{UWz%���K6Jt���-]]	~���{,i��G�i����g����a~���a����_:`���'�}�s��Dc���!z��G��xrzS����
:�jKf����d�:�Ë&ɪ]�i�=<�2���м����3�Θ�$�A"ɬ9���>�Ɯ;����I2��E�ó�dm����}F�5k���6)�L\R��~��.Ӻ���nU�2֜�ff����[��78<4�M�$%Ӵ)KӁsY���L�M�M=Mف����n�ٻG�e�'+�iIW��d��-��N�˒f�J���֎�5��׭�Y�`2���P2�l�4�]�3�M�^�����gI�Ԯ�� T'~{\ˁs1�Y�ѶE{oR,���g�����u����C�f/��@����jM$=	�Bos��;}l���-!����b�$I�`�!������d��c��$k��$��@�y�S��������������)�9�%ɵ�m�ɓɫ��6l� vmاaY���6<��ڨ5Fe���:d�e��]����G_<��1��sژ'�n6v��+��s�wĸV�x�y+�v�MV^��C�LX�;�<Va�+�:c�?�ֹ�]���~�z����rͳ�Zk��������:����i�m����w����~a�/\�aۆ�耍����M��ț�n6c�7p�c��_L�x[�_j����O8cˁ���국��f�/o�����iv��k�}�/��u�|~�8X�Q{���Nݮ�ӷ��C;���_;�岉��>:�;�<y�]���~���t����ԍ�Zw[�}i����O���5{��k�7���ߞ�w��o���)3���f>��}���y��_����^�xs�p���]v�w�:����>��#78���s���vܣ'�w⸓.8����O;��	g����g�t�%�u���Oν���]���W^~�{������|r�S�����r�W�ܺ�����o��󮻮����N|��<<���?^���lz��g|n�秼8��^���]_�ፉo���x�����^�тO��_�?����ڕ\�|���pݨG6��3p�{�ye�A��w�J3W����*7W�^���[��5�Ys�Z�}�:����z^��>�p��&l��&{l�x�S7���W_nL���MZ���լ��ns���������=���7�x�XY���כ�-l�v[5�~�vޱ{����������^8麶;w~l�K������n�!;w�2w�q]��vo�+�+O�j�.����=��/���7_�֊���޺�}��͘3�p���3����{�~WϹ}�C���O�W]�ɢ���/����Z���c>c�%߹��������#�Q����ѳ�Y|�����q?<��.��U'^{�/N����N�|�����?9��3�8�Գ~�c�>�C�=��_��?�`���h�O�^<��/�x�֗�}E�\��U�|�Օkֽv������冎w����C7/�ղ[�����κ��;����~s�o���߽|�w�{���������~�؃?t��w���G��g���������'>�������̎��n������^���F�<�o+�����������vx}�o.}��^����<��'�����>��Ã����n���c��_���a��Fm:�Q���Yc�{����ݱ҂��]����U�d��V;~���8u��ֺb�׹g���{q���0z��7�z�6�}��7;a�K�������Ҹ�Mh�r���n��6�|�'7����[�ro�x�{��-���JfU��v|u���A�زӔ�}�e��C[O���kv���Gwy���]+_���ީ�N���{^�6f���'�����W~����ӷ��{l�&�dm3�����x��C��{�~�Ϲ{�S�^_����٢�Ż/�}�A�����:��e���{�*�m~8;���ݏ����>�S�=���w��p�9�铞;��S^:��察���>��3�;���>�чgp��~x�G���@�%}���.��%���ν��+��򰫎��q??��3����+���w\�����M�����o�ආ�+w����~��o�;w�]�]�w��Y�ιo���>0�����!��c9�ѓ�x�c�?������'yj��s����������em|~�ƾ����x�ٗ��ݯ������?.{���/~�7�x�ތ��ݿ��ƿV|�����m>��x�'�$:�%�5Lj8���Q{��{�}��1?��7��m��+����U6Z����V�r��V?s���<�K׾v��ֽ�����+�_�x�&6]��M�?S�ŭw����O8g��zh뗷�x����m�X��+��˲�ٙ�"q��Uݣ5�ؿm���cvXw�	;�u�̘����I���z�?M~�}��7��t�޹tʏ����\��	���L?b���͞��⛛|K~{J߬��?}�+n����3�����7�>�o�9��m��������?|���.^��%���_?(9x�e㿣���C�]r�I�_r��G>~�kG7�ޱ�/�k9��=~0p�ܓ�|�)�N���CO;�G�~�ǜy�Y��踳O<�sO?����~r��_x�E����G.��e?���+����ّ??���9�ڳ���/.���n��������7��WO��̭�����o���?�͊;G�n�]��W�g�{W�o�}�����������w<rˣ7���]���O\���<���O�磟9�/�?{�s�����x�{/��i/���K_���;���?����o���Vo���޷�}��w��w�n|������~壷>��'� rX8��< �8!I&�+�jŊ��N��]e��X��I�J�s�I�����I2�KI"�a��g�ly0�j9.͹�g�G��1����Ã���צ�L?h�C'�Y<���Z�ޕv�8IF`��'�utT=`M�?���iI2p�{�14��V��@���u�5x� ��������������v`�dc����ߍW��U!pS�0�0{��_�+p|zT/^'����gԅx����xm��7z{�~o�~��ܿ�~��W�zF?�W�3&w�ok��9�v2�@���z�3��i/VJ������hq�>�[�P�Bp�OH%8�����/���� \�������p�e
Ҝ.p�j���|��n]	��Š�o��?If�����W[2%iǘ���|�|�En����&��[S�p,D�2�:�L8�=Ȁ�Au��z�c8���!O��e���7�} �s�;�5-�:��g��?�?�2�\�M#V���+i��A��"N��tm�Aw���$%30����@f$#:W������S�7i�D�� ����?�!� s?�4�@;��J�8�-��SX����e��|�I|�?o:��1� $�)sd���2���K���gA�qs������l��g��A�s�"��m��j�R��������;����2<k�9���9C��/�?���?<kpQu`v���м����������ۧ���:ch�������޶I�ƞ�E����Uf���N��$sՁFL=�����������8�����e��JO���m}��;�zzۺ�'��vv�M�n۳h� ��:z��;�v�u�uU�'O�n���tOn��k����=��mJo�q���E�ա�:	K�ӿ�kx~S�u���Ý���7���|]}�{v�aܝ��zv�6N����Ll�i�k�~��J�(�[OW[kowKGޭcZ'�6;���Z'u�j�5�eƤUkk�k��j��Z��e��2ejwgKG�^m��z���ٗ�i�q϶�����ImS�:�����abwKo��)}]S{z�'v�y���6�TİgGGD��=ugz�Si^Rm�v�����܊ί��D�ڊ�\48�z�Т�A"���k�fk��?oF5?��Ξ*�e5�Xm��a�����)�J�L����=���Y���H�A�;ZZw��!?:��)=nW~3��sw7d�������.�8�����3��z �jc3���s���]F0u������Ӷ۴6K�qjWo{'���	c���S�4�T�2eZ�Ķ�>ld����I=U�E<����og:��JOKgW�S
��n��d���I������������#��i��fZ����A?�c��V�2���'[�F�
+a�ҽ�U�jt�W���^U�ƅIU�����~�������8���R-2�YiҊ�����~�f��k�q����O�����2��~�	f��ʚf�[�O0�
Q1Qz��8(���8:���'%�JM��=����&2�9�Ei)h�V)�T���c�e�k<�R��<2Z�Hוl�����AGͳ*�]��(4�M%�2����*�)�s]iMs�Y4�q����u�r+5�`�Iiy5n�E�م�Y-�)�@g�٪�%�#�%�_������Ό��Ԡ<F�J�J��X�05e��T�B�)����U%�%�1rנ�*Nf$3T/�i%C8ľS�v�Y��̬#�J�F�-6bY�܎>K�MX�6�1�HJ�H�U��&�2l�p�4[��M-5�$*���NA�� �Ժ#��e�F���ƪ�fRn����I�2G.�R�H��
<P�C�G%�Lf��5!�$��j�x�י��5��56��@���0�)l�8�z�k��~��R�Sk+p
��Q�:��Ƥ�ր�{� ��)�T�[��^G0��$��e�TY�#f��p0ZV��dXOp�T�9��@H7�R)�F+s�u���I)@�����r�
$�tMH:�z��mKx��ž�K@�p�D�G�%���ʩ�%]C��T�
ǲ�Gs�Q6+SN�����~*���L���p�8w�9iwRA#�5f��	%�AX���K�uRKK�uk3if=�Fa���K��*\U��y��#2���"�'����&�q4�xMl�i���'~D�T���@+G�$ͬ'������ ���B�%�ZU8|,ܣ%ͬ'�/����;�m��>�"���N���a�dA�t����,U�YUX�ι�:�^��#��0�	`��FA�֕�0�j�:~(+L	��CU�q	Q��u�Dq,����p���?CGQ�h������?�>�����=PH�?C�_�?�*L���ʩE��;�:��*J���+58��Iޖ��	�LC�d/n6�FC��� \��_1�?�$U��N)"�(�4����@���#&��I]�)U�6�2�)p
P{سդ�������z��� ��
�C����{*qR�JM1�T�� �42�U�hB�TJ*t��b5,���h;0�\��Z�F���*p�Z�!�:�t�jx		,��a�`�FT`)��| �#$9bFhf���Q�ë�R��%ͬ'$ia9Eq˒$�TFp\W��a�_G�,Q��$�#�Ru怈�HS5�@)���76�R�Zҹ 2�,�R:J����4��pE���$"��(���p�_G���r��>��P����j�PX��zB�n�w��0#�8y���(�؎$�'�0��C
cB�"�R�iA3R�z�0	�o� $CZ�f̠�p�v�u�!p}�5�#݃[� �Z(|���	x�a�����G��j ,*J�d1����%!�B,a9�8�]E钬!Be��'&���2� h�LI�gD`E��Q����.8 9�([����
�Ԡ�O"e*O%� ��d:EG��e:PFX�i�s�a
���X!�F$�.}0�P�9e,��c}G�U!(kd�FƁ�C&������ܭ�#�i��)�%�j���QĎ��8 ��A�=9X�/ WS���wD<Eg9X�?	��=�ȭ�;

� ,���{���P �K��x�@*�@� Dq��<+֋l�>Y�R�g�C���	r�W �b���A`��SN���D૘+��()���@�vd)*�������� ��)���BN<YuT�Рd�Ry��Dq�jd8��)2��(J9��*3*�0#I�p�BW�,�(���)�T�j2�3G�tQ ��W��(�G,U��bV!����?C �A"�/�-wE�k�b��d�qF p�d�>0� 5����%�*V(��F�RR�wK�;�O��g� "wnX4�T��R��1+���[0��+#sQ��+p���W�@(�"ׁsd��Y�G&+��x�(@ #C^N³!X��
�W��3"��yXE�3tP��U��)����������TE���U%�R)�g�	�����
�е��=�T ,�ܣL��(��q��5 aԹGC�F���pl�{,:
�r�F�s:P�I�-�J������Pmi8a8��Sa���f%=�bIU��gR���TH�>����mZ�6��"���'��DO^�[���"�g�[����� ��(q�Q�3
v�%��(��:��eU�b`���� 	E>��C��YVG.z"�d 䒪3���u�3����w�(���Ѯ~(]-����YVK.zr��T�#+�����jmy�񫥴�CH)ὔs͚`z%+-'�@��`(�%���%�	;��e��ؓ���M�@�=m��=Y�(4�� �1�p�䝡�����KL$J�����մ(u^2@��)�T���2r`K���fN�3.d;��\�I:~$=��@�{�~��*�5z��t�S�V��9�jڧ.q�q���s��"�	U6��eSY���}�eS��)�f�)0�iKzFϔR�I �`��J�+S���@ rZ6�D�ŠU~8��L#��� -���/!o�ی��-[Pi�ϴq��2�Ig��D\���j�yY��y ���%=#A���i��Ǩ"CePڧ,�q�������T3��%
�SOU�5�& ����kAu*�Жt���U���dÆd��	dwH�H��Z=�Z�QIy*�Q0�&+���%^3���q�yBR��w*qpNz�KӘ��`S���K2��Pt��A�����OQ�_S�q�z�(iNV�M�$&H	��1
WlDO	� ��L�Qqr�Ty
��H���cJ��D�7��(�J�¸K�0�0�
=Ed�?'���4��\������`t�L%(9�qZ˭��P�3���� �!����U�'�g��g��=�}�f�P���L�H�EO[�f�����J�r���0�(sy�@���Y�t<�aj�9EV�

M��)���r=YfiNF�G�A�c��KI���I����U�HV��q�Tw�u�J'WyOn4��(K�cOzPĀ%H��H�)a��\�,���B֨W��j��J
o���Y���+�g�łzl��i�S�`���p�����e��}Ҝ��g�'��	�h
���.
�V�;r�p�6��fȊ���,3��	�
���~��C����2+�QT��/zR%�S>'Ҹ~H�����V ��* ����J	�J^�o�O���(��;�×t�R��ۢ'E�T@[2*S�(�I�"�0���#f�̸���P>MZ=DOU�3n�����:=Z�甔��2?�Isfy��V���<�8z�{R�R����K�?�ׄ��ZP}Or 1:F��q�TR��cq����A*0��W�e`��SGeR5��%�z䚹�^=�.iĞP�Y�F��SN�9�O�}~ڛ }̃7K]D�H}��J���(!��P�	 ń�"]D"l�dIt��Đg�(Rq�Q\d�V�ʒ�BfX[
���1����)\�t�����vȅQ.H�o�,�Ӕ��� ���'J�����)[�
MȨX.�#(�ڼgF�L�9�x��=�|�t=��BBz�������&�bR���a��F��q��PyM
�i��!�	I��F����pʤ���<O=	�iQr�q�����N(���)�)���Y&�
27�dqѮB7?���%C���
۳����ڭ�O�[��Mb�rÕMVm�n�y��Ӽ��c�y�u�yfF�~�mD�Ȫ��]:���EP� ���!������&z�Dw�4E�j�������.�=�o���Cs��1���s�.l�6��3�r�VYrIR�\�����$��uH����!��-�G:^�g\DR���ݓWJ:^M7��+i�Ƚ礥��@�x���8�Z�*����ע��b6�K��缔���$2c�tňx��G{�UѩOZ�	��2�-����Ll�HCT�=�����jEh1:��N�|T��2�EhE`t��������9�@��9^ZB��rFO�s[�/�uG��J@�@��Μ��;��?1��N=���%u��RbǫSzt�Zm�]x+��At����n��A� �����,�W�7;���D�I��'qX��E��}+��n
�:W#�V�zU~��x��|H�HԎ�~rAѵM/�@��٬���Đo�n�1�I�9?��x^�$�Z�6�df�r��B�疛�k�I�
z��0������9�L�d<�D��Gb�\�	"o58='��|7�e���,#_$] �����ߦ�3"�d�9��7$��V�$�~�5Г%��*52�Y�u�6�p����,_B� ���U�nЄn��x�Q䭈�~��":Jߍ*z9�SIתa�<�$��|~!��f�i�Pf<)����s��]�kuY�$N%t�����Bb�0y�I-�9�)�r^�?^�V���Ҧ*��X.3�^��`��ZA�����r�_�s��z�Z��yu~������a�s]�ru��_A�xA7a�v�㕩7H�D~�#'�)4]��ym�g��iH�Ck��Y�n2o��o��S(RɜW��H|84�TOB�r��(Z�V#�
$g~�ty]z^�_�r��MV� 	�)��&�F�DM�9'�nN�y�5�\!�N�<
��<	��K* 3HV&��|Λ�f�ji	��6���r�Z%z�@ʠ%�J���7����I
���`o�\+�_�� �K����V1(�w��/�$�c��"ZAx�J2+F��+ϋ�٠.ጵ��S9�k=/9k�j�)�u� (�t�d^��N&2?B�+���
}��a��;F:Mu���v�c�tN�:��PQ&���E� �˱��@������q/�\x���>P+saϓ�z�D��܏�è�U3��PH��IN�]�[\�g��=L��K�)q��0�g�,�"��|	�X�j��_I����\�X�\+�i�z�5{O 2�^�"��­	�2V��~��� �e�_:�˯��7�y�,d�ݵ��D��e�C���r�*@�6tC����C9�*0DAfE�������'����ޠ�{2]|��I�HH��
�L���{��/�� p Y�ܤ�j�N!�d�y��t��n2��0L���u [ɘ�![|΂yO����������0Z"���D��x��0�W��đ����0p�և[�ڛ4'o�<bfl���OhE��yC�@��Z�'��1�GC�8
��{.FW��-0�7�HN�7��Uy_�#��Ⱦ�C:������EuӬ yȬ8��a8D�'��&�V�}��d�0}7�9��1�#	���p~ǰ�=o�a�՟0���1CF��/���{�2{�~܈ahZ�Ρ�2�Z��1��7&�T|���6�WO��er�Y<���_ʲ0��>BrJB��"��xx���ӄ���[`(��a
S!i���+)��H�׳�a���%G���$6ă�D�)Y�D��8A�q#��p�ޭ�L�ԑ���[`��F�{؁��WD�i$�QyI�g�y��g>nR&�]7�����Na96+��n=o�0X:��v�]<� 恷�0Xm�r��y3�yC��T�%|�IY�1t�� �t�6�,b��=�a��>��F�\[�#$��I��ﱧ�BR�UP���h���-0��2��T��c1��[r�S�1kU1�i��R��I���1}އ$��U�5���ɽS �¹�"�z#����,���eIoC"b����Z:pR���E#$���J��] x�*"��y=�T������[`,'�E�	gA7e3�[`,�ER#汧�F�'D �O�;�֟E�0��4��U����ED�� w�n\i)�-0]m�NL�B��)��F��X��_*��AF#�_xCY�&z��-0�>�f�e����GɈa����̼��TH��AF��2���T�j_ޗȈa$2'�}���|��g2b$����&�t����0HWT*�$���1��a\��x�g�"#������0U���x��H�UэPYNbX��2b�n�R�Rg���0�"������K
�y�)�O�%9J����YDC�\�NC7�9D#	q�@j���F��
�xT��XЇ�a��yX$\E8!����1"w�- m�:�ce1��Oɛ@Zx�9��FRu1LL���I�fàՆq�����~܈a�¸D���G����d�0hաbZ�:ݤ�k��R�nP�2�𵷋�a0��A Ï(�㐊FR���`��i�3�[`��S���5ؼJ�x����JB��`��U�0��/sOʀ�1�J��-0ZC�H���С�i=o�a��m`���%�>��������-�'��W�u(�[`�����w�i�k
*bŘ�ABk��MK_�P�(�Wo�
*�}*=��511}ZW�����*b�L�+�����n��T�0���+}���	0��uZ1�E�U�;���>`�y�(�{�!z݁��>�Q�(�[�ިXx����1���?�ʐK��k�y�`AA� |�Qt���Y�0��3�a�*t=bEwȳ� |ȧ:��Q�F�9}(�=F�1�k}~���xo�ȭx�F�3�!X��Ǫ�a�e!��A�@�P�V� �����҆ڕ��ޗ�A�p��V|mEG�+}D媠}p+��a���ح�礦˙��FY�@א��R��ۦ���D�=�?71��k�{���)�C�atV$m��R+��:b
�,�&�&���ǩ:bڭwx��T���WG�黩�s�9i����a�d�^B^�C�<>��h�SAPT��"���k�x���`��l��?�À�{��X�Ky݉F#��O�#���5D�"|2K�T 9=�p��`
�Y<��O�Hn�`
��%@g��@執�a0��nE+���Iz^��FCS���B�J��a�
5��M~M��sވa0E𓚤Zu�Y:bLa}�Hw��,��5DC_�ࡄ�¹�}~�#�q�گ�(N����y7T3<���lz�c"���)'?�:���8d"�A�

Co�2C�R¸�Ak�{����5�bW�G��5T$	�E]��-�뺉�Z�Ã��89o�a���!�׀��͛�a�5���-OZ���Z=ޡ'����%��1�� a�n����/��a{5�C��X@Z_G4��W���W0o"���~oàU�:�!�/H�k�&bËg�=4T������pև(�:i"�!��^ʇ�� �L�0`Pa�z� ^7à5�>�X�¸:�L�0��Z�;��ri��Ɛ����4�<7À�P�pB*?,�[`����-��GHz��kL&b��3���6X<��g&b�{Á��C��x�D�PP!'�q5�k�&b0dv�CӰc��#�1�e� ��]<\��+11��Z!���b#o�a� ���z�J2��[`C�)�Y��z��o�0�M�c f�&�k��+ۈa,}Q^�fC}�����1P�!��.Z��f=o�a�V�<�����]�����{Ɲ3�!7����E1��a�p��`0�c�����Bɹ��l�0"!B
̛��/����0����o����(��2�����xa	��q��_o�0��*�W�����<o�a,U�Āj^�ع�b#���)��R�y%���җn�7@��Oڈa0��
2@*��5R1��uK��wA��<o�a�G%����K�d��-b�3��ᰃ�4�x�-0����n:⃔<&���%�;pt�͇qrPao�XCߐ�I�t֕�r��Xz�x���[��Iϲ��w�Z,]��֥��Rw�$�_�Q���d   	pHYs  %  %IR$�   �eXIfII*     (           >       F   i�    N       %     %      �    R  �    ~  ��    x       ASCII   Screenshot�lK  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:exif="http://ns.adobe.com/exif/1.0/">
         <exif:PixelYDimension>1662</exif:PixelYDimension>
         <exif:PixelXDimension>338</exif:PixelXDimension>
         <exif:UserComment>Screenshot</exif:UserComment>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
���%  ��IDATx�t�wsd�y�y�gH��+��Ֆݤ�5ÝU�P����kc���~�Մ���H턺�M�a����*
ޤϼ���yϹ@��l�@e޼����S����+
���P*�B�Z���~�F��W�e�7�y���A(����{��9����g���O��W�X̟���o��~���>�ߧ�^i?��5�S��B�\	�lƙ�%d�o6�g��nh�l?�)�Z��1��;�O)�K�VSSS�d4��תzϟ]�z�>�Կ�ݞ��h�3�U�Vt���is ��MOO�iS�F�f7⚴� n��� ��y9�p](��}����}�<!�ߧ�S@��$���{���g�~e#�$�
�7 �0.��H�,�
�������~�`3==z�������~��+������R�:�F��n���b���C�!���/���������011!��e�r���I�I �/0�����R4�q�H��S$C|��I?	� �� �kN?�n��a����䟉C lŸ�V��C��Y6��X1`7�(�L�&''�1�͚N{������VWW�~�ޥ���5��+�r�t:��>�����밷�J��������)�E���O�[B�	Ћo|�u�D- 7�H	xIL����_TB/5�6��u�^�V71��tO�r
�)���d�9���~��E���咉Y�nǈuR�?<<�s�./���NDv&��B���?����WXYY̝МX��T� ���o�����mX_ꍉ�{�)�N��,�Ά��#-�an�ۡ�j@P��diE3
���=�W��"�������u:m�=a��j��ʟ����gÈ���#�FNC ���j-�f���Pww����01Y�Ŝ�qb����P0j�2 p�߱��0$�H��)[/ϫ�R�+:�����0�����f�ik���?�1\�r5�������&�`���q\� ����ógk�Љ0k�<cn��c������B��Yϔd��k�F=��Q2��UJ\����QR�6@� F�L���]1��!���Y#����O��wR"grr*,//��㣰�jSԉ�  	�����ܬ��3��a~~^����ֵsssZ�ٳg��Wv��p X��:��⚙[�v�����OLN������%{o�^��3�������i��8(9Q q�X�~�
�� �`�K�+aqqQTztd�l�=�1 i~vND���?ί��77eI�9�`@r���0ʘ���כ�,�k�	 �~m�� ��� З�����W�k�%��`����S[�Rx��w� <Ar?� Y���W��UX{�,|�����\������Ξ]5.�gm}�Ν[[���Ja��>��}+R�U��>:�$�j�8��Xgݮ�+�bq�5�Z-��5�ɥ7�h����,�P�h�����t���-!�ڨj!+&
�X����]����e�ՍZV@=�i��6����ٙ���m��SS�09?a�Z�1D0(����`��0$��f�Z-k�z��Q�+Q��o�fC?++g� �}6��jќ�p�bx�b]߁8X���C�g2�1B���e��ph�8bтtK
s���"�ܬ�D�C�"8�u�)�)�@�:��Dٌ�鴻:_g�ͩɦ )��{X,20�t�ʕЙ��A/_�4��� P�RG�j�ڂ��07LO7��W._�s�!#[ό���߻'N��_�ҷ/��e��@��@�Hy��D�Q�3��%��M�A��lƲdO�$����K����@뜰�1QeE���A�:��b��:�����G����¢�uh��m��)�3rH�N�6P���h��"�c<y�D�2�ƀ�	0�˻�����A�о��vwvEm��R�[�ˍ�F��[3q�L�mr��7��3�+1b�C�Ǧ�^oJ1vQCq�H�����a�D"��GY�9��M����2{S�s�("�gH1 *������ϟ��7V\6�5�+u��ã�8*9��a_�Al����C7!]�OfL2�6��$�rg6wj�Ȃ�QPX	���Š��h_��W�dY�6��Xל[]�&����E�>�{e�?�7����^�a�(JL���-]�rL@Ƥ�z�Ϣ%M����ɓ���o�#�C�j�b׈��7r-�n��S&��-,�cqQ���gl�:�b���P�錾E�a���Ǿ�D<a�E 3����~s�U�HD4j�.���E�h��b�0��c^3���c76��Lb>�'���x��^���KN���M����ٰo� �����p�r��2 @be<c��#����� ��!�5��{��ލ��#}�XA�E�,'b�bn�P����f�l�1eg<wg�C`D�d��j��dW�BxDw:]�^|�����ƾ����.�9��"I��8��(��R�i��UbMڗa1��E�L�C�\�����}���h ��(��-8���|�p��w �=!?�b�`l��ŋ���Ʉ����1����_H!��$&�PD�DKt��P����r�x
ݬ�?����qʚVWW%����{��T Q �{���80��̭Ȋ2�ʞy`�#��H��~i���G#ʰI�r�*�O�l���MmЧ�3Ƃ!k��sm���3�g��`߃��������08;3z�q(�cf Ϝ0�xl���jz��ޮ �?!��e q)AkkϤO�Pj�G}��w���� pNj�K�.�	�������YKY!{�H@���5t�!��� J��`�ez`b���`��/A"V���q�GI&2:���.�ƒ�p	�� brS�d3�(�y �OX�iJ�e
�������ϝ%q����lCnV.��I�;4��,LΠq�r�<t���Q,�g���eYNl���=C�ŋ�Ddw�����gr_8�G��Qs� ���/��3�_�M(��!���(�Ơ":����n����s�$���'��)���x�k����p�K����{* �������w���h!����s�9Q$�B$�1�L�υ)�tɼ)K6��ƽ�Y +����y��C�� ,./���1ſ��J���1q�%l�b/x.z����B$pHh�H�8�q���Dt�,�D�"Q�T��{���B�z�߉!"�L/�O,�Z�,�@��.y�?ZZ��*a	�ƴ�<��ttӁ�� �,$�������_w�i ET���&�/L�`�/��(Ul�ݚ��Zqy
U�]8E�nH���[�1�`���H����(Ii��M�㔮w"z�2x�������x��������I�H����0	 �v���H2��Q����\0Q��)�(�s
)�hp���&�� �3uD,��ˤPA��������r��u��{z����}���ׯ�� �r��S��a�`SljwoO��XGW��]4�����l���d_�<���ϠT7�l��L,�o�N����t�3Q��YB�m�����\ r�&�TAӐ�.��س���MU�ݴ���D� e ɻT����!�zt���b����Ƒ�]�b�|]�|A��������u�`(�n�t�6�����(����e |���)�eCʖ�ݿ��_�����bc#� �#�|��~O�êa[1y6�x���ل: vJ�7V���7�x×2qH�B/ ;�r�V�S��S��ו���X�>l�3A���W5�`�X��B��3%���I65�ӦW)�!0M��6ͺB���X��9x��[)�nO���gW��^
?��Q�X�n�;$ipCr(�8�=N�t岛��cPHx��<z�8�5~ ��$�*�ΐ�:�N�.�5O�<Ud�?�+N6cV�K�Ք�ȩJi����N���J�ŀ{,�T�G`��XX���!E������D�8%��5<��(��H�&�*7G_���2��{ ˈ�@�������;�H6����p��j�z����)d1g�Čm��O��e�t~�嗹8@�H�Oz����ښ8�?�P��K%z��@*I���eC����w�
8k�FM���	�_��ڂ�x�5��@ �p=y�+DI�xۈ��K<}��!`#�X+�4��-�6I��l����D�֑�!璲�[1%�A�Ŝ�HČ[�r��]���0k@^4j�׀��W�j �]]=gb�g��L�	��u,��s�w(��u�]������s
@b�o��:><R����T�]�8��hbṉ��m���Ŭ!{w7��XWL?�2R�E3n
� ��k�{ ��UWܕŸ�ҭ�,G��z�tL��5�Y5�Ƌ��I)i��zAN�1+g{�#pW�������$�5`@aq���B'�޾<Վ�)��Ƥ<�ho:e����O��ggf�u�m,��|E\� �]s�3�!d����=یQ�){�7�|�{  � �?�DA,�'�=�h2����%��#���BO��Ϟ]�ߵzU2ߨ�dԵkW÷�~k�~G:T{@�,�7
�q�L"�9y��.��?#�x/,M����v횸B�h��ȓp��'"�D��/(��ܒ�үU��Z,R���]�.Y����Ʊ|<����{f�C�����+�VM��^"�h�MJ�"�-S���p�ٳ��" ��Ec��/Dg�8EؿX1e�J�Ư�5���8��4�UP��@%J}��n�� ��I]��d#V��!Y6�67?k"�%��������Q`R�O�sh끈��1���^�0�-(j��޸�4-	�T���_O��ˀxy��P�Ke�M��cC��ޮ����f��@�x�$u<��Ő z��LT�����pw?RaP��!�Z��e���Y:���sCI�&�R7����@��e�2f2�DWa�% {}�e,��������JWd �D")0(X+�Y>�������X{���ck��� �1f���ʣ�f�cEL��ɋ<��گ�(���c�π�պ�f(ׅ�}U� �ub�����2

� 7Wb8RXY���3a�LU�ب���0<��6��#2;	A(\���Wo�sAf�YT+f^�}��P�ô�P�+׺LkއS ^�d��Yu��<�Z��Y1|eģ5JAx�Ϟ>�5�6L|c� �@ �f"����ѣ�yб������7��R!^�4��1ȅ�L��(%���P��c:�X�B��F��g{�,,��MG�c�� �T�K��"ڠ����?�x'�4 #U�4F�`ld� e�LW=~�<\0����+F"� z.2��p����k�E�#7���|���-"$� 0�B�R�2���
q:�o�\�����Q[�	D�	��p����!��0����N���!)�U�ߊY�dM�8�9d��Ҋg 톄7X��{���
`!RH��H�1^�����>�j�&i�7�k�������pG����3/󩅚Yep�Д����O�<����(#�4d!R=߰'�� a8�d���+�ޚ�2 ��@2/[:*���AĀ� �˗.�[�nI
�{�%��r<��>N�
"�(�sf���+Ix(�!��Mq! xt�6`x�m{g[����-�E�"2`�w�}W���=��5B,袉R�Ħ�l�y�jǳ~��OHRa2�R-��H��s_h���:�����#J�&J�HfOG �PD-Nݵ�W�����H��� ��z���e�bأ%"-��d�nˊ�rѪ�G�7"���R�0���F|��*̟rH!�����.������h�����X�X���� d`�ݸqS���������!F)$��6v,DVc�'���b3":]����Ѩ�b+���2�����^�m�^S΂��D,\���w� >6�w�}'��B5˧�22��
n��z�psRD�j�{�b������@@O�bs��'	P�R�!Q�S��.�X��R�h�����9�T�X�5$�q��}��1J�8�F�Ǩ���G2Ѡd�T�}��X�Q�= &&k��G��҄u1��P���}/s��Hr�o+�b�ā�j��8�F�(��b�E�$��.6��|��P�v�����ޫq ;y�	$𣠡qg�I���>��t�B���T��_�Q����X�������ǥ����ū�	��%3Y=�'>��]�R�����_� �@۹s���s�6o�T�/%eH�"J�ݿ+'%�#JWl��(D����vd��Km�X|`��j�����w�M�`T{<�ᡂ�k֍�c�T��\�{��h����zݣ�OMD^�v[�=�2e"�{�QE�7��:���y��I7��6{O�r�1�bVN��%�ć�t���1*Cda��(Q��1�#P7�q�LS�>n���<u6�|�Y�w�(�[
��X�[�u����,��=�>�=���S�(�k `tÉ�2���B�qN�)7q�rp�g�cA��TP�QĞ?�補�	�����ML�{+�W�R],T�%N�.r������S/�%eBOv�h8g�ɻy�fx�b]I|�(�#9%ĮG�<� DGt������t)?��'J|<��#�<Q�� ����zD ��Y)w��7���)w�F������ˉ-K�#�@�W6z?�!^��Ck/�ߐ�T����q�'�t��d�\ �_mz��@"\�r]�Wq1Ux�;R_�g�^��y�h�0H�-���w0�"���%Ʀ�-���;,��SF�ޑ)}Ҳ'���Q1���|���TI��rB�������� ���f����u�xp
?��Se�؄C��͉YY�hø�\�3�����EW{"��W�D8_om��񒥆����Yqׄփ����´��x���O��B�{�cx�S�X�`�'8m�K� ����v�PJj��E�.R(��/c�lQ�gg�z�@�A�b�����fdy�Q���q\�~����d!&���s ޻ﾧr~��ߛQA�c@�e�M�+D}��+��;���N�3��dBW�#ѓDxa��?_�|�Mx���M,�#T�Djq����� ��(���5Ǵ���Id��Hj��B����f�&馈����T3�D���3��8[����?w�lTjn�C9�CU�{>ً�r z\���#�G*P�-����tbRU�/_�
��V�������&|%�NGQ%�ٟ��#�<8�H0@e�V���.b
uC ��>x>��3�q%JG��olo��X�F�rl��dN�lI�g�I����	Q�*�]�ES\P,��`���J?D��P�
��x�I_�&o�>!Ԡt��LSj|ɿ��hK_�z.Y38B�C�������ڱ��.�
  �?7�w̪��?��v�Y#���ס9�O�?>�jt�fjo�X����r.����� vMm�SƄQAo�O�,����O�)��?�ڌ���W���i����H��/#JB�=W��6M�M*�5���֒:�����r1:K��%�SV�΢����~%R��$�}�o���V/t��p��=����wE�� �IG��B�^>k[���H��= �{]X=���T}��f�C����*�΄��n(�L����C����+.���Q��hP��!d� ���%"�U#�%C>ݦqcoߌ�I���q��s��l4�" ZLo��H���2?djrB�����U5���TT8��{Ks�p��m�	#ْ���M8傽�3�'��=�,PP�[険��w���r���I[��8 ���H�TE���#Q噅��2@�H�*�?���Z��pbꦊG���gR|A"}��;�U`��8�g�;Jm�ʭ�P�X��1�:|#"J��؈x�dA�ʿ僈!�r��b�I!�+F�w��� ��d*> �HE��۷r��T��*�r����\��萡�+Y��)@PӾ����x��X~���S"�gYA�yA��3y�y�@Fg���LZ����,Cn(���GO"烅V�޵Z���hi�;>'>�A�����z��I��T�ԿFH�tM�G9_�rM����J,n�➒L�8��/�J���ã	!����s����W�U���)"���ɘ�������r[[{.���������6+f*|��w��Ç�m������M���s������bu�B冐A�{+oa��B��	㪙��"���L�U!4C�[�-����aoǬ�U3��M�-I�:�AT*kV'�ًu��jF<��������eEIE���Μ��(vI�L4�S����&�$��H!�RqT��7 MNM��:&��k����g�^G����r *b�
���W��p�7�p�bf�����y�и휙��aŵ�弊^�����cؚq�@4ܥ�E=�9���g�h�x��wLy�ߢ����:����+�/U+�L���5�^�������"K�Fu�9 g�6@L�1!��\�!��,�;�߿��p[[[�L�`P��U@qP�-"��bY֏�v�#�$B٘�7nݔ���_��/!����#Y3�ؖ�%��
�Lfnl�D��;ъ����
@z����j.��~Ĺ}��i��&�fz�15-qI] �8��&8��SQ]��J�L�]�jI���Q�s���(J���k
�ye�RX{�L50�p�����)�c,�P,g��	�"T�@��%�+���+����f��wR�B���y�?ܹ#�q���\>S^'j���&"�h�����Ϗ�5E�!r�\C4$�����1��YT���!�b��>���#lˏ�a�0�ҙ,7���nGa���Ԕ��` Һ��H��S��'��|���z��5��N?ִ��˞:���ce�"
(�&s��>+A�Al/�#�<�b��(z�0*�\����٭���?|����2��7��*Y��pL��typڤ�jeh)J^j=:l�b��]ZxN��2q�}��z���o�����H2����x��CҼp����b���O��Չ� ������R�������I��I�r��Tyr�[
x�;xB��k����OA���b�O>�Ĩ��p��u��(P�Fg�D�ɗ\�b�v�P^�G~�N4�czF�G�j�M:	 *�H1_��4�,.�WR��<z���R�q�Ç���Ad�?�`̺�8jѡň����6<1�J�n[�ƍ�Ѿ$ �;����H�I�.@�"â�p=\B<o�,����Dc��'��X��@A �
ѥ���ѽ�B��L&,2���ԧ�������+	Z�/�R���hـw����( �䱟=}�����eq��/������'&g$ǹ'b�Pz�.Z�9NQkQ�E�<|�P��ԟK�.+�8E���A��˯����
AU�(����BS/��NʎHNI��A�P7�%kĶ"�J�?�I��[�J �pq��333!���mI�d
�	kC��� ~`w�'��Y&^�O]o&G6O�u�3:
 �!V0��M��#ߝ�J/x%�[Gp)�g %���eh��l'GB=��KsZ�@�"
y�˵���^�8z�6�ݱ�!���ǚ�s��qP;�x��q(�)I�!�����e};�44g�]�iґ��*�y����@�{�~^k�RWa�'e�K�JD�;t!�6Y����8������	.*��� 9�օ�����VN
�"�}�QQ9l�D�jiy^�QG@Y�\&:�/���96nE<��S��!�Ì9�ݖ���ޖ�C�M��J��I�F6�ĲW/�v_LU��a4�׃��MJdU���M�x����|-��
}�؎�y�DH�V�>SЛ='��(�K�/y�=�_�cE2Q���ߪ���䓏?�"�(�ʎ���A(�`��Ca@�tsFE���Z�{��8�MD�Sy���'^v�(~>l��Y���*�O�Z����ѡO������JŔg�&�9�p��+揠�[��2jF��"#1���g��(."��v2an�De�hp���2���ئS��8ZY�-:�'RX ��։�X�a�%�"r������TgE��ֆBț���z�-�6^��*LO3J2=[Gc`�Ox
�M��M*�*�^P柾�ڋ��fOj�AȅX�eD��ҀR=cb1����s�@���\ژTE��	�I��Yo(y�v"��3��.��|��ɔC������U��J����{&i��ΈMɑ���i^ӊ�B�� �а�+Z�X����~�3�>��h1T�B><�/��R KE)BMlB��o;;:n�H�6}q��E)O�$��E�G2��3c�װ!��Ԅ��G1y�M[�B!�-s_��p����5��n1��*���
8���* ��F�0H�b�c�$�I���F5{9>��$B
c9wӱ��ۦ�ѯ��W&��P�����J�P�=e*�=�{�*�9��)Ku!F\B)l ��-u�h.z��A����7d�C�=V�4���0������vh*��b��V�����0�1��o�'$�pf�4��խ�@t%�	iJ�f��f���V�9�N���3�s�\h��]��a�P%�/�z�/i�نX��(ℱG�Dl���U'E���KW�h��e����X��T�Q��]Y�,���/?R�Bg�Q��w�F�[����,�'�H�8���g�,}��>K��3K._��� �C�c�����0�޻']	@h4�厬��ޚN!�Z�j�8�m3���8����'C6��"��cxɞ����l�5&�94�'(��a"�X�y�J�(�Z-����+2#Sʕ�ǭ�7U
�l�+>��Sq���H���j�F����)q�][�1g�>�π���> �J�k�u��US��35%�����I�;��`�bQ����4J�,:��pp%ZTT!..-(��g`���l�����d�1'Ί�
�e�����K�F���?��Z�v����Ӏ�<�82s� >P�^e�pǮm�X!fBP��IsCP���s�Hi�D���Q�yy�l `�j�WRwE	?���L����xaVR���$b �!��
����}�ԇ2�pGj���X(*.��l֮����Q�s,�Z��p�!,7D��-������i�sR-�<��(W����*�jiK#X	�1��zd3�ǿ�7���B�tE�ñ#kH�L���Ϥ��uT����\�?ڱɾcA 淿�'��aq8	dAu<�I�CC׎$>��oK�cU��{q��ݝ~�)��n8����pfA�Z�����xޚF4�����MD�[	�}�Ǵ��:�M�Q�A�6����y�����O�Q���)F�B��{R��9ߞ)�#S�d��)��u�F%��=�{�u���[�5�F�� ��]�}��L?ͪ5��Gm��
IB~���W�\���3/�S�rET�C�X6}`��*��&� �h�?�P TH����s���� ����Uc�(�k=z$���4�!!N(�E��B�y�U��łە������]q?�E��"�����C����J��1�bx^�p �	j��lo(@|�cB����i�F�(K�y�&��q�QO�<��ȿ�Z�Qi�du�PP,}��+"�iL���Q��%�B���� QXV*Q�y���dA���/�I�e�_}���L5�wx ���j'9F�3�ڝG�P����1��7a0��f)#�'�B��ʅ�*�1�Ǳ��D)S�CU9s�ٻﾣ�A�^��~��˚!���/�["LB�͸��0��^��W��Z��X��U8yi�SzR�h��P&��}܁����#q4Ā��Nk����f¥�F�%t�X�P܇,K�PDq�q<�WV�b4�yp1kR��!��ycM��H\�,+S�
���3g���\�b��TKh����= �7�-���A>Hy�6~^�����1�k�9T�8�����' ����Y��hB�A��@,��Ԑɂ�L�g�F(j$��lM���pN[5�Q�io]ʝ�-�N�M�0"�w�;�@�d��i߈����K�0� 0���58��ѯ�`�p�H�vQ��z,�%x��B@l�Ƒ��Գ@������/�@/BK�jP�m1A�~���0���d⺷�z[���G*~�=�Bg<� �AD����\ȕ�`T���u!���R���o߾>��SQ(���i�4��z���=��+g�63r"#�ܚwo���{���3%�: 8�0��*��_��93K^}ЦF�}zC�e�<+(֏`�E��I�t����1Z�����ű���5�j�ƕ?.����U��(C2vs�q��(ޭ���8oP�LL$	x�i"�Xp�������ˍ)������S����,�&��JP�:?pg��aȜE��4gC�`=3/�C��^@����bD/�i�i�ٺ���� �k�n(�"��\�\�;zr�TFU��e�ʍ�����v1BlG���B��Vy�K��z(
�9���>z�O|��pc��>�ţ�U�a�g\oq/�mE�m���7�:5`�ؓ��0���ſU2�����N�eL��sG�3D�����6ۓ�T��h䳳��LWyթ�/�#��s@jr�j�>qʱ���E�В�`��R�tAȋ@hj���RG\Y)J&+�������r��Q�$o4�$���� R����DJ<�2��ը q�@��"�1�S��r�L�K�W�Q|��?�I��4U:�Ue�w~�14�G�=I�b�C (e�P����a���?|[<$�����|�b�k��>�k���Y���I���j�&��wzw��y�Sِ�7c$�G�z���.�p~5Z^�s������*�]>D�,����z��P_�/l23=+dj\�!jSs��xY�#��)���8�]� �\U��}zvvU�����3����b��s��hA#��3�\DS?�WK���&]+��<�	Y,*�i��e�a  J�AP6{ �a�%��P*[&���TOhfva6���1�O��4�u�^�)����q!�hT�1Wa����g������p�#"l#i@> �~�g��|d�j��J�Q��\���iq�w�NH�a>b�oۂ)����4c qQ�;��ߛ�p �H��y*�0ġSh�D$lL �`? `߸y���Uש1��B)�m�4��n�{~(A�S��J:ڢ��Ou�Yb��4;;��ý(V��e�*���A�D���{�נ0
�yr��x�x�
��3\.�Í�>���5��'_���d����w��T#R� bP�*���b�C��< ƍ7L�����h�`�|�����8�z�d2�  �Q��)���]'[bޖd�]{��y!��'�����嫗��Ֆ,$5��y�����a�`���Ռf7߹C"륒]�s �R$�u��Q�)���������<l����\�hn�����[�n��?�\�M�	P`wOx���SH�P �ԨQ @�ģ���NÛ��x�(a�=�6�����D�:�*.q����J;�~�0J5c(b͕��$o�����A��-?���<�y�ܓ�Ha^ӄ8C�`�!eɊ�Ќ:<9\��h��"�4v6��U�:�<���z��a���23Ow�ÇO���T���ޡQ�9[k/L��4����K2q��³�k����3
�=;~&ca1Nz����$v4��ņ�$�p�L�=�����N���-�V|iׅ�����/�_I�<��X�|f~Q�|��a.[r,ød�~V�`?�rfn!/��v��j4z��Κ"\gx?ʤ����C���R��GD�K�$ON�5X�`�P�"�yxpO���޶tWC������Q�"Q.�$	�r��=y�����~���ݻ�@X=>j��k�B��{��#Ǆ��8IgRqTC��GSS��~�v9z:0�By�<���- {��mQ>�W��!lv��`�"Y1$WT��b݇�5��jΆ��������sa�9gD���:�ɸ"�����t4�4hmjʇ�������``;0�a�P!x��\�=a��C"���1X� �B��o�Bsg{ꔶ���
eK�Gvɒ�� !�b����ƱTr_~�:�g0��7r	��~��X�.�t�e2y��7oi�o�\�Q4_�D!���[�ҵ���9#Y&A�7�v miq��0���X�@��ڔu�Ӳt�&��x�`O�EW�NL@]41��)CGz>��(�ux8��HB>R��ߥI��h���Q�<u妘V��6���"��F��%�VUD��~�d}�8eƳX���W��L�Q��Sؚ�At��������`�*3@[֢�ݞFq��+��u�/�E��ܗ��Ȅ�1c�-Y6:�������Xքc��	=#{!����#\�^JS�T%C����]M�M���[~@M�0�����;���V�%��7�L)�S99<���L���@�XR��;���Bɦ����|�A[��Q�\��9���Dhzgr�01k:^iG�=���x�Ǡ`�P�ѡ�� ��ǀx��w���T�����9d4f5ҸG��͏��{cS�;O(��+�`Y��V�4O����gC(X�.I�����Ayhɱ�bq䇎����x��^��1��o"�ϖ��Y�*>L>�1
�4U�"�;B� 24 ؔ5Vu����!Oȸw��Nh�k������]9O�uA� 0/��0��'up �"�Y٫��� �	{<7��C)dv'+.���Y/���4��c���vm?8�H�t0�����Xlǖ>��y�R���I)�Pd9�DN��3��rL�#V��r�>=�2�yr>�	c���"%5`&�0����#�Hڰ`"����ȡ��2��Y�:�̀퓪_���L��P����߹s���R�a���3��5�\���T37Q	F��K���:̧���='�h������9�_1�#�w{�n�0%E��^>�3���}/]��[��9?A��{��2(KQG�9���(�@�<~�T�C/bb&���[��AU)IW0��Y�@' L?��}�̄D�'�#��}���Ԩ/�ͫA��qp��#}����ȿ�T��|˴k�(N�rc"�1X
v��ɫN���c�'p�_�/Ao����G��a�H7����2��8�J9?��Q�	;i��B���·���_�E�2B�H iZ���6����o���A�5�ׯ��vO�_��FT$g��L�p �I,Ϧ���!L��A�O�
W�>N��pxO�Z/o��P�� �F�ii�qx%'L8Χ5���p p�`X���'�X/�x:t?���{��r~Iz�n���R�䔟~�g�"3�6�^29>�G����a�c!�M��F�?x�
By��?�y�K�ǁ��X�R~���R�y���˯�T��Vg0B6�&5�U"{!M�Nsx9֔F�G���c"1�:�d����8�1�)��S��NU!?� ���S���SMS~:�-�C�Lj��������R/���xz��v�X5�MO�a�������3��Xa������J���n{˰=+�@�z1�����/r ���Q:�s�Oq�r���顯��&$ܔ�}xt�<ap���?�R��N�1d4b4Vj��,�a���)�F �Þ���:\�S 8����<�A<��{ 7|*�w�Y$pX��U������U��f�g�!��P�S��H��̀�sr��U񒦶!�YF q嶩�hö�+T�h���v?I�N�pbc �GKL늵aXP�����s�J�I�����c��C�?d�'O?0q��|M�|Ճ����d����3�ʘz#,.W.X�M2��y�t,Sb;{�a*�X1��A���'��x&�;H�������?RN�߃߈bge|��VE�`��&�������Z^@���?�ՕN�
	:"v�C|?����������c{�
j�
�Ӝ.�:���������T�r��m��i�.!? ��K�t8����å�#M)�������ё�70�	��~��89uR����[��R%%���$��Ѵ�hz�j�B���+O�%����n���$�o{����/��WR��ߎ��7oݒ��NH�JfN#�t�$�r��K�Q�ra`>��GAy�ss
�4��4yl�(G�r-Er���?����41���KG�a�<%%y�5)]�F,󉥘�XJ?��bkT����F��׏?Ϯ��f�9�����4�f�b�!jw3%^SFo&�C���Ek�ǀ1ỹ���31gY �=^ɂ�j:Δ�	 �0v��e�nD���Y&k|`ʟ�S�e+�1��O{ÚJ"Q�{+~�-�
�!�q,�k~*VP�U���`�L�L�C�/_��s��D~�L%�}@AԽ�^~v��O��\&{�'���i�;�7��W���߰�|.�7~�DE#)2��6 �Q?��:ܤ`AB*W�6�Ή�(��yP)�Ks��-�U���@b6��0�W�����	\�\7$�p�G���Tl{f����9�i����7��A׏���b0���P�eË�C��^�����(՜�a~���@����� e�NF�u0�~X�G�?1鐟t(�8���Q��U���μ�˽t�3qg�^l�����TBa�;5�m�"j�%� R	E}��ǲH�S�~=/�q,#E������8r�D���^I�8WDی�0����d�r;���z�98�x�����hu�ǝh@܉x#���<��u$���oR�kv����d������s���^-W�Ir�=�6�V��'O�1%5��_���i�h?Ü���
���*��8�x�l���.d� ��C�
����|	��9Vẃ󈬧�&*R:�Dʁ�f/���f�2(��fǄ�A���?k{B48�ٳ�Ⲇq����T�� 3�DME�o4��/<ΨH�c ~�<���ݽ#C� n���X?z S����t�	���z���d�CRo7l�؅^�We���(��ŘΞ�P
T�"�X+P�~��%�^�B�FGS�0>��o�FPp_bY���U\T.������l�i�='�|"6�<�P��JU+�#'��7p�䴧�u�Y�.ʥ��}C��g�D$�I�҉��$�`�v"�8 X�[�q�z1"������o��N���*B�0�{.N��L��#�V�8��T���({���  Ԟ��1K)��3D޿�,(s��^��)�D���T£�F��5B��� �HB�l�/�����|j��`
�D��~I�ȍlr#�-�#}��cn�]�N��ў����Q���:��@~�Έ�ڦV���n�{Ko��F;��{�I�+1!6�ӄC�횕�0Hj�X�Œ�`��cJr�v)s��m���Ac��	�Z���`�n�%G��'�Fo� 	�8z�*|8��u��Y�L�I�r���Ǵ������n��3�AF:�7/x��j�Rz]/��{��z ��(i�NU�&]�9'~��A�!�?ͅ䓭s�����T��ls����id7"��A���ʆ���~�sE��w�����s�U�8G�ٓ��p�N{6�����#&�MEi�4G�a�l��i��P{�(�<G�cn��M�t �A��1b��p�}�`Nr`Oj���=2���^Ҝȁ��1��)��,�oU�R�;qoD}��:�t�>����_f��6v6�0<�	����7A@
����Q��)������ |��Е�*:w~2�kYG�����)�y#���������� �(�ſ��d�%�)�~�#�Z����\��9�ju�8�����o�ƳY/���|V��G����*�Y�(���X�u�.Sh��;��")U���b�ח�>l��
x�x��Ԓm�
��!#{�Yu��*��!
��~���o����w:���L�V������Yq ��  dAi�8�l#׽�!o�������������[Y���,�Ap�t*�=�HM����:MhM��i̘��ׯ��QV'A�t�EE������Ux)�gi�n���K'�3�����,�L�l�'�����R^3�.�YN|��产X�U���O�P5�)���R��F(AI���U�Ky�$�w��1�h;m�`�zs�%�l�r�TH+�[@#�ѩ8�s=K2>���CP��G����ى[��􅘯\�����T���*f�uF�?zC3���|��ION1y6�5��Mg��<>,���}�
?,ޝ��w@�g�8y��������+�%����YB�B!XU�`�Tپ!�L���y0�jp���� M��B�f >�֞(�%v��cDi�)�`�#ǳ2;�i��~�� W������,̫7��ZP� �}�]�O�o,Do����G�������@X��p��e!L�.GbLD�F�{��ώ��4�%��B�����?�3f)�I�����.�) ? �#�P@��l��Z�"?O�# �CR���~(�&[�[�؎�~�I�w^�R&W��@�Cy��{�)�݋S��t��ťF�#��P�[:�w Q��P?8����k�zQ}#D��1������>����<��eᐂqJJ�<�0Z�7(�7Gj�
&;�o���,�L�6�����-{�3��+h��O��;ԧ���H ���7Z%�V=�0uƹ]��� I	�X|�{�u�D�#`&7�C ��/�&�?�����Q��@�B<z{�w�[f 5�W�&���)l*�&���ܐ&�AD���ܑ��d" ����P|#t�r)�W�@�g�����G~���J��:�M��Ea�����hQ-i�-�IS$�rZI�$"��������*I�Є=i�TO�,���9l�D�f������^&� 0���j�*��<�vz!5H�0f�ъT@��Z���r�b�@�u��=�������C~V	H�fv�ƊTވ'��{~w͞�qD{u��B �*�;^^�d��œ�3,^Gvs~��M:[ӡ���$��y�I����P����t��g����1�I�BFt�)p*1�T��_�3ߗcE=D��4�u�rz�W4�#'���=�>�ݩs�Q��v�1P^|ǐ5F�P�L�Z[��y �k�X�gWW��~����{�jMc��,Oҏ���?���A�):�Ͼw��۪�e�I(Dh9�A.C��8^��0n��Y��W� �o���$��cM��Py^ޑՋ����|�������@J�| �G��{ò�WE?G��C<��Z��q{G1K�6���>Q�/>�����Y��h����Lr,>�6�i4���ӜR���y,(y���FmPoYJv�d!�
%���z���lqO�=�hb�r���{N�D�QJ"��Ǎ���$� b��$�.Fc*��׿�g���YX9\����Y�x8�⃨�an6�.AߨG������-�˷�&Ș�;�4U�|�.XYݘ�1;�(�f$�^O�x~�7ި��b]���it��y�:5 �kg�[�H�ˏԟ�|�mx&��i(M�4�H�š/<=[���j	�OD$��b�,b�q@��)zP �m��;�}-$�Vn�h�i<ՌǡuOM���W�]�x�qM	�
4�Y��>D����pp�uV�X��v�C?Sf������h:�4N�\��s�7S.F%B��=l�ZZ�8S��G
�`a*�)E�(� �gŚa1n�����{���E#�UI>c�a�2R�e�Y��UJᓏ?`��{��с�϶������~���O�̝�S	�ah칭����F�G��a܉"&��J^�]����q ���B�����k~��Ο_� �ơ3���8G%q\�O*T�GG"zLw�����~B� k�Yb׮�ɳ��x���a=0C�s0�0�P�n\�L�<[͈����D]�S�pv(���F�`-�e���譲2DN��P<Wa{��O����.�W��r�"s�ΔjB��C"
��8�:Ey�ǈ��ٺ>���q�{G$s�Y�߃8e�4��mm�l�D3�	9��\	��$�f��w��H�����OM�N�#(��I6���iE��ڲ��H�_KD�B2<g�QG��^>�EG�&b�����8ٳSt����-�i��9Xk,��0����7�n����kEg/���B|�����p5��S���r����%��|�ng7���ۨ�g��#�Ux"�����F�0�6<x�bC+�2�A�#�_���S��|�b�x���k/����9�>���R�����Ţ!؍#�Ҍu�?]�($R�L4�J��S�8/��,�Z������~^�&�jN��+E��Ғ�Gd`k�O�a����:�e�
Q���N�P߽q&2�M:e'�!�"�E�d��}�3�8)��ޒ؄�1�iO�@�� ��}���j#����A��2�ʊ�f!�|�Ӥq�x��cM�1�@�5��#�Z��Xe��TS
Ċ��>m�2�4��D�6��Y�X�z֑�������A:(JD�^7�<�U��Ӫ���Ѐ3�P��(0H7^:'6|�^Ws�~(Eӱ͏��6=�B��M�����H�U��7��ɐ@°O8���T�TG>}jjFHK4��lc)�s�Ė�q+S�c[1i�m?x�� ~޶M3��C �*��I;�bl�i�T:)g��|���W�~�bQ�2%��sR�=/wX:p��|�R9
��KZ��KqR�y�⤲�n+�ݰFjF�N�v�6�?\�GN�
��8�B8��R,��MCJ��^x&�T}�U7����$�E��:����X�qQ:��'��cCL��gojJ�{�lͻ�H���JE Ka	��N%�G���Hn�z�s��a�so(�C�%�0Ԍɋ��+W��ڣ���<} j;W��JWc%!T���2D��=�e�=�WZ�<Z��ҖAfk�y<, e?77��� J�8#S��&�	D!c�fu�΋=z�A���*u0;-c�C��i��9D��V7�LxyW������h�S0�mK&�8�}�&��՗_�.��Ce>�- ��'����ԁ���|a2U���ot�v������u�O,6e��C���_4�2'T�>�"K�/~�����]P��=u��^�����)�dq���b(����jЉ��zL-�^(��P�~S㧒ŋ�"�Ʌ�̡�n�6H ��>H�1�[�75��A�:���b>�ZOX{�7�dN�P�<)�Om�>�O���Q Z�����+��]^�tvy�O*H�Uv��͇U�Ÿ�b�]lǒV�|�Z�"�=!\=(1�_5 b=AXU34�/���a=�%`�dS�Zd�a\_�O%5r|�DRn$m�:�C7�I�(�u�2uQ��!����a$�dT7��¿�6����]>�,��+Ȳ�pJ�jޡ#c��x����9��J������/�C�F6���hm|�N��N�C7Qϕ�8VY��*R��ͦ��������n��/s�\��~�I�Q����L�(Ɓn��:C�2{%�p:�gb�h�� ���0���$RQ�9(�%�賒��t��W�	�DުʢV���Z�X-%M؄v(/aN���ޅ�}�~�O)�sYkg�e�f��S.!:�W�.��c�J���ێ�q�;�I@L��Ұ�8y�w�����<ܣh�q���8h�J�G��X�>�X��R4Q�	1�Q�����YU�^�'��r�RɨQ�OSM�O�8=�4��[6�Q�T/&�C���ZF�Τ���x�h�[�c��Gc?#���8Aw�Rk�Qt�µIjrPD`
0j�EDZ�w[���45�&������)�T�n(
ϢB�̑BP��L�8�GU! ��#���x��D��8�ӓTň�R�o*YIM�.G�j���%��*��=╅��'� w����ǉt!;rt�`����9m������	�l����- ��H-F ���T?�C�����A�B|�O����|�JYl��XO1��ˑk���̜�aՓ���+�c�ѯ��â�1�^wI"Q��Iu�����\�8�K`|iƲ:���\�	�y� f�J.U��'91=��u���bDXp�D�H�$!˧y���sW�Y~�obo�ꙅ4 7ł\L��8��-I���{�s��Թq�6~c`�C�(�"J,J���rH'�$�����E�A4.��Gt�
��N��E쥂�A�2-��o��Q�>�C���q!	��zKN�A:��9!��B>�0W��8��/ǡc����q4 h�h�a�\�1�3��2��p��t+�!bĐ�P�ȹ��|�0/8p�qDH�#)�qa��u��
9窍-�.�����(s����l��(�l
��O�M�.F�|h�n>������#��rwE�dr��r<�:�W
.2��Q!���ܙ�H=����F�uS,`(FG����{�pR��S����W�O���.����b�N�`��"�S��Qju�iN8�!�7�*�ur2�ʣ,ϚU5@�)M�D����Q<.QM9v\�#����ƈ�4�����T����I��eD�-�,��#��rѩ�R�J;�g��q���5�sTp+i��0��A4�X�&%��d��|�R.�+���2}{2����L��Բ LSsQ�_'b��0{����~�\�霋8,�O���n6�Iuы��+68�� ��%3����d�Rı�f\r�k��P��`��2�ݔ��,��6[*��Q�xr~ր��!�8s�@���;��[�2�M�<�jMJB� ��Tm��yb��룘ױ��8�O�m��#I\�T(��[l=e���^w�AjŨ����%Y)�_���yv�aw����K
��=�j�m�q��#,7�M�Y��c?��3�K�}�������Fy�T/>�+�G����7.�b�^�H�>�#��@�,ˣ ���yM��8�S,�	㓂����~D� :��)GҥZ��J"��눙UK��t_HzF�Ǜ��(�jM1�BX֍#"���KĲQ^達y&1�gΞ�Ę�R��tbM�%�=xDw�y��tF4����ˣT|�r�?���8u� d���*r!�.����٣�>�}��,W��u��m`!,�Q{ۆ�M|���?S<�ON-�u&��>:9�M�� (��Ũ`	�Z�H�L�����B@	�tԏ�X������M���;����O����$�5��T /�� 5�0)y7T:u^�뙔��NN�so��;k�J%)m�t��'q<>�<�9��j!�����|����(J1���J�����^�8Ώ�(K��R,���j�zf���r;ܘ��>�Ps�C��ygR��"��S��l(��� �գC�����Ƀ*|
[Q��8�E�,��&>�A�#�M���Mބ����P�lDg�Tj�P������ Y��VH�'�ݏ��(��
�vj1j����x�V�t�9��e�8?w@('%�+�c���uMR%F�A)��{���hO�(�y�N�b����A�@����+�c	Յ�(E5�!o1��)�MX�{PR=,Q؝�}}���Tc��X���n��ϗ�\�(,���(F5m(5_��Wj�C�e)�xRz�ɧA.6 2רe�뺂��z��he�w~�r�6�l�9��z/[�h������z�5U;������81�cB�Hytf�Ձ�&�ԻPt�{b��?b(c��L]	k�X_t�ۃ� ��m��(G$�*��7�H�7�s)G~GE�Xڔ3��\Z Sv�<�0�%��2�3�i+�^2 �Y҉%G�GvO�A�#�p����|��/��!n�k ��x��1�]�M22�]D�*�*x� �NEי�}۱���u���n�H5�
�U<�NH}+��1�g���N�XYiP�h��k�w�5v��S/e�?�9��Ee�x ���{�"��-Q��b�4��I��}�U�z�>דC��))q���" �+Q��򖷁w��E��S���V��%
�$R��.f_dIp|R:�!��&oWp�u�LT����E9襋�e��$O����8C�G��>�3���P*�"}h����#P�bO>'�)�F}�������˄b%h2�u�m:��"(������p��9m�jD�/nF�3{���ҏ	0��?&(\O�=�	�K0^��R� �T2�K�����n�R}?�f��@.�'��Ѧ�Xn�h�ٽo*��[j٣�8���d]�c��`���_�^ih���Zbab���81O:b�F�7�By������Z
Tn��US�&sG��l'����0u+e;���)8��2t�N˞y 1S��{~�ӧ�#��}�A�3�\���W<�[��~�I.��!1z|4�A�0^8^����熼�~^�X�4~xpC�n���wT�4􁡈A�Z�,G#�z̡�_I����'[�~��|��)oj_)��X8R�iD�7�:�뀊� dAQԳr�
�z�K�aWӠ��y
P�U6g�=<ؕ����� ���zc��p�����+�����~�����bt0�3䝏�r�j����^�'��0R�zfz³���!#Syk��$�t��)t��Gٜ�;�sF����d�{�aKMMH�t���MK_�Ϥr#)�}���������k,sd�q
y_�<���ʀ�qEt��u����y-X�j%f2co޸�Gi�쎐\�x���t0���r�/����^=������cýX����a/�m�ұQ'2�n�K2��z�:1/.M^wG�e%8��i
Ay���Ǯ�f)��Vq��^�8ܺuM%<h�<����ڵ+����Ҏƒ�_|n�xV��Ұ�'�UjJuN�4A�F�/6츣�_�8q�^��8�
�L��|�6�4��@��nK\yaI���hP��7ߺ®�Sv�4@e2tl�^���qˌD��yΒ!����b���@�nw0̳z�A�����~�䄇8b��P��|����H��!0�Ϻv��:�@4K:}�BJ�uvyA���T�G��̲�Eͩ�OL�'bx�"�M	+F%Eb�b>)+��T�j_s���A��g��=&����XM�3q����5�T5�xͬ*��GD�P���YP�u�qM(3�����`]QnI�֡,�I���	��V�&d�L2�0�2t& rw�fʺ�בy�r$�����:Z��k>?��ci�i���\]Z.����u�d<|�Q�J0���	9ч�ǡc�[^Y�)������.����+D4�-p�
�㈔����g����tzjү�a)��,Mf>��ry�Gq���2�����o@R�FK���L��R)���T:*���w5b���z��d�P@m��**�V��R�)TB5;uP�bC�@V��+��b�%��nt��"랬%�G<>>����r�ʔ�7�no)�7�U���J1�hJ,1�U%��h�W@�m{���38�G��G�T�C8A���cs|�DD�8�c�hC�'�܎I�0fc�6Ⱥ�3�0GG��v�Q<�=~�D�dL�k2�]�>�=(7��k���O�G�M���2�
`�WX���䧩t)Q�����]�NfW �E�(EG4�u\���>�,*��$��qO�����e<Ƒv��{���y���b4`���%D���s�O��#gfbn 7@���l3<Y�*�W.���^<o��M���a��x$����`L�Z�,ǈ�,)�F�S~}�j�g�=/6��m��fJ��u�2�(J96�g�Dm�0u��oV]̓���Kx�����`�a���x!�ŋ�,��x�]Iʜw�_�\�����i=0J�Y��ٙ04��?a�"p��I��b�N�'ad4L/i�Z[�9:*K*��i�����%�!.�q�
5�<��3jx��w¥k�E}>ý�c�Ut�jq������������������ZPn_|��q�81�1�� 0�
B��?�Q]c�m&��O���P��V{�����V�g��8ɱ4��h ���[�:�B��Q�z�Xv��f�S;�S�j,J"��Qu
B�z�|t,�#A:���t
�j*}��D���1�i�S����|�x�j5/�ݑ2��2{��A>��G)�4oc�ǣ�Y>j��J|�����y�f���G��GtO�Ϲw�^̗��I��c{i����S>�1�(}�7�3W���Y���J�1T�(2����bE�C=1����RU����v��¼Dia�nj�Z)L3�!���O��>c�Ӕ������s)=����구�b<��S�'�Xy�0#9��w4*{B,�$DP1y�CH���h �ӏ)%������A?F��Ĭe�؎���ɔP��;wD9L^#�����#�e�@�T�|�����PX3:�>z"ЈC��9���]�tJ���=�6����=oa�h�hDF#l�z�*H`����aX__��u���Q[C�@}Cp����@lMS�X]���@�,c!A1�
��Gf����0�NS����8��	��p�i�tcA22k.���T�d�"�i�ǋNGL��2���$�X>��ЉD��z�؂�%\��J>3�o)�#mp�b�������P-H�C������F.eR�3j*�/����6UO��iN��-[F�+�h�M'�fnO��::�@e�lMIɳ�5q�`��J)/�!�=��g⥁��ZҌ
�k����[���!�U�2\X()��Bqd��7
�5�ik'&z�ށJB�����
�t��aL){����?�@�N_ll f�߸~SG��5Q�e����ǰ��əH�Q\a!5�#kҌ
,/��:��~VV�˟p1}(�bgo_3��~�=��85c@���� <x�T�|7���K""�*׎h��
��gT�!�@�SHHe9��#$Q1]K��W�cӾ
�Ǟ�&!�{2˜=p/޸��=ӂ���P\�Z�2��zw!�i��4߰-6�b��G�-�!������Wr��2��6f(Y�1�^o�TU��K>1th��?��WΞ�u4C�������_�"�x�Nxnb	�
%δ��3��{�,N_����.1�nd��B���˕�t��(�3�������~^�>\��U���e?Sо�f�#�� R�z�}�F2?(<���h�s�Ȓ���V���?�1Ί�_:�	��?ƏY�kb²y�ۦP�D�S��A�VT#�J��g���1�Y͠��<��ta��+U��(T�g��D�ߺuC�QN�"s����[��vk�,����!���F�uO�������O�{p�yfי�͡�V�B!�� ��&;wK#��3K��`���[���n���NlF`�DΨTN7�;����n��� ��������ٛ1��u�o���mStey1|{Kb��#��Uök�"BcTR(�b���NoDTBT�c%<|�Xe�-������z���8&����\�[�-�y$�G���WT��|:��s�g�6E��D-ka;�e5���*:L��+4S�[XB�OA��ƚ�����08l>eb$�{p7L�1��f�f�f,��rPatxhT7�5b�����t�ظ�0j˶�A��m�Ėe�Ǆf�4�Ҍ�|SZ��zر�/�s��7|���~8��@=�
l��]��\4~�M2�?���j���V����p���8��%SJ���0pD�yajH�3s!�ZN���|�P�<�ytU�6�; �l)�+���F�V6�V%`Ak�1�d��)��̟�nԢɌ�[,s ^�ˌW�]3a��h�d2�>�_9X��\J��@f[1�T�aO:��טG�A"R��4g���	ᘿv�eGJ6�T���� �ad�tŒZ�}t9��.����G�h~�VoN�E��+�m::pnu/pþ����ͺ"�۷�I���\i��p��7�w�l� �1����>������ճg�2i��˦T����9�g�y�s�^��~!{E�1;;�B((]`�J��5�P)���l��@�*�u!�:�} K�D	���,9> ���܉ ��~�|C$2N����	�٘-v��I-_Gx�"Y.����Z}!Ac�0	�LJFn��8���vH�Pt	���w�?
ׯ��	ڍ�ÿ�7�'��������C݌Đ��x��I[�ez-,Ǝ��ZW��i�nZ���}/�(������p����{�{_��ǟ|bI�n*��Q�zY�
nF�]W#+�oQS�����a*��zͼ/-��Z��+�l���G0���O�ugD+Hh�����)���|�Hj"�!'^EgT#lf#9Ul>���$`�r[\Q����8�I3acNҚJY�~67jB} "�?ܯ�m��$J̔?s�X9��r�rq��P����)r*�����F�!e�8�v��$!��#3��ͪ�1�q}�'�WWkZ`և[�$�AX�j�ـ�q����T*��J[�:W�RfK��(��\7���ZV����[.�9�!枹�&	9���1����N�G���#c!��}Nj	l&�t���ƒmJUfjr����Q<c��ٳy��J�5[����ܹ�)D��VI:E=�E��w>j~�l~H�v�/]��N��<7?���z����6�W Q��X7�Ұ'?�M� rT|#�-E�GǬu�D+��|�4U�@�'�;�ߔ$���Ʀ�X���<���S�-�L���?�(�L h	 ��Q�=�U�Ʀ����|�+��vL����H�d�"1�� :J������ƂrHn@b��q�I� E��a���E)����A7SȂ���LQ?��O��������?�/é��L�A� ���C��6�:���nr�Ty[PV)�T'+�G1�]�"aG^g#��1I���qQ	Uu��&dq)/S:�9����1�<��?�i  cǗ#�X:�5]KP@�%�Fk�~�fS�R]vѰ�Bj~g3���k ]��>��4���lJ�L�Ӭ�d�k4t0�D�, %����.}�Y+
X�nd e��z�g��v�A�,,��YY&�6$4t !�)�*ab|�����'
|���֟���Ǵ[�-p�L}ZXS��/M��)��rY�G�\�g66�0�[�?��a�0o����<t���X5�MKw��	m��ڢ���\'l�V @�ot�bP6Ӕ��e����-�q22�(��8hQO�L�>�e�f� �i�d�ڼiz"E��G6;������j���/�	33S2)����ɿAO808jA����-�G���'��t��Q���%�5cIi!W�ν���V���e�8����p���H��u5�����8��̖�l���T_m1����<v섈WF�,��5����mˀ��;<�/�,1)���Q��ɰ�~0Ts����!�+����H�9����p!�{���ʚJ���zػk�I��v���&}�n>��Ǔ����޼u':0&ǎ����dfh~zN��ܙ���r��|�[�ߖ�$C���Q�E��<�9�w���U�B���S��+W4ǈ	z��Y[̂��>ۈ;����̌�-H��6����k������(�|V+��en5{��h��=~	f�����!
Zc��Ld�#������77µ�W�)C�̲����];T�X��θ��Q���d�\.��¡C�u�@Ob��7\a���}����_=<��N��R�w�ȑH3&�6�vlt$r��zzT�Z�o��*�|���~m\Z��Z��fL�cv8�����<0dڼ_f�(H@R2�522�葟�ϫT��ߩ8��D�>�v/̈��e��� �q5���9�L�Pm?���6�.J��[��{�����,E�������:eu���H�{P��g3��0m���V�z�L�	'����
,<z�R���t;���姦�%SQ����V���\&fZ	L��*|.�u:�Tc��o���+�.$3=������e��0�:3;'à�L�=�HR�k7	�e���F@E1�P%`�ص�j���4��)^�T*&.�8<�T�P�&����:=0�2>�l����u�����%~��φ�Nm��;2Җ��jAע��l�}^T��XtS��^�������-��m�	�x%����ɓ�Tp$� :$��7	��/_()��ہ�����n�a+
F�p�+F*�\~\�+�G�y��z�PC�����ٳK�.�Y����l$u;�N���5މ%F6$��e�E�'�ȇ�g��P��;!�̶Ɏv<���=lW��DYQ�.�V��k����6���'�����RZ��0*�9PZ3+$ev�\�&HΝ;�ȇ���������֡��>�͇���,��R����q1C�)f;|�w����I3��2�E	�x&9>�M�g���g�ӟQ,fz�LQݶ��:d�DyD�B�ح����&c|�!�
	������5P�T�k6�z�]�t>"ͽpV�-���S�&s�%����V���8���=z��!��-����ߗ	,\�!�����>ᯡ7�c�D�C��oߦ<Hbő茛�g���W��{�.�R�,�����0e?#	O�SF�(�:3��z3$*8�Хp��Q�Z���Q	�V�Wl]�,�\�H��x���r0�[Z->;�MH�&_�vټ��M��Wi�E5��7u}�lw�w�4<��ia3�='Y���^�ܾ�(���^Y����*̦L��-��FH�H<��zS�{�� %(yN5�e>k���� �!JBb׮:eW�]~��K�#����Bo�L��BSJ�O-�����|�>Qq��9��[J1i4�8��0�\Q_�k��B�a����̏��*M����(kA.����ĕшk��҆l���T��~� ��{w���H\�E��nO{yI m���踅��ʲ����r�z	���A��aS�d�bP���[��`D`�%�l�#��a��=��8�J� �D!���W�Tm�!ϔp*�����N�M����I�oܸ�>�6w�,ü-dZ5��JV�3�o8�13i��Æ�r��5�*�К�&y���(�3����=3�S��6��z�X����5K�-[�n���]�`����ȕ��n�"c�G�T(���Ǉ�}�JB*�~�&"#�b�fN��D��|��O`���#����E�з��J�ݻ?��^9����ou@H���#��q�琉����b!��ɵ�6�@(�����^j��'��?��S��0�T�	<\TyE3��Eh\90=�z@���Wכ{b˳��ڑ��;I�������z��^��T����I3�EC����RDSo4z	t�@����LrҢ���Q�ՉS��U;$�R�5�.����1�1���k�����J�h��29 ��4 %ZY��px�ZP���&�f�6%�y�0��"��߉�h��w���hkˑ<�5x�O�L��0D�����{�<�8VMohj���R:�E�"M6�n�{�(>[��KP�#U�E=���)G|�.F��9�':EP/�� 	�Z��ʪ�#	�M�?nkG4����b8`\ZU�VXYZK�������?�|iTP!ăA@�@D/|;�i�d&D>��><']�B�&��y�T��?T�#憬��T�m��c����سxؚ��1i@E�eb?˧�й�����U���%���]G$q�=S�H� R�,zr�/f���e��9t�px��u�AV����[�Zh4���..U�ЅW�n��/���=L	t"�eD��Y'~�|V�F����{[@K��kk�2,D���|T���8�l?����V3*DL�����W�
�.^�w��)�3�V�W�'H��~&�sjŧ{��v0^:}ZU_�'aO��YV[a��\jyn�E��q<������Vc�SRR���Ȕ�#��� �N�f�<��3�Aʆ"���qRʀ���9�tj8���~���f6�T`S�V���V�Dp5�Y�3�w����3�U�����yĶg�.��K0Ծ��tUڂU���tj1d�о^��'�
�0��{̊s�CXw�౦�N�?$��	e'<�q�)6�E�C�����!ª���**�֪>�OR��H�Q�H�U��f�q`ǵ��#�[;˷zܳR��On��2f���q�7)1V6i��af���a��frNٟ�j���ܶ]�6��fT�⦺������a(�]��C�\���J$�_>����c^�H���\��䓲&��)���~��G7dHξ�l�6�7��(��GL�@���84r����?�קB/(��o 7'�̒�n�I���:cE"�����(p����)�M!�#�����S7f؍EA�jq����:@7ڷTz�-�CFb�2�.]�T�{�o��w�牪���q��Bɵ0 y�v(�)�:��W�������+g\�A>��b�䷿��ݖ1-��@]����~���T�?�^�GX���9���x�r��&�O��㺃 :V���W��R�ҩ�~�KeV���e)��Z�7-��%�;�����Ő걎r���m9�Ro����5i��o��>	���߈�	�<��t�ٽ�p�x�B�Ǐ���'
Y=	�]g�'o�:�B�tZ:�_]�(�Wa�#�ȑXJx{A��S�#�M��،Z�)�D@�z�L-�29�.J��C��CH՘�R��_�Á�xK��I��n3� �N�0,�"�rc���H0��aC|Ī��fQ�YY��:�~A��Y��/��o8�X�SG%g�FJ?{������>��i	R�����;u�D�o���8�z��p��qs���1�WR��d���m�|�+{������߆3g��e[��}������}��pĜ4K �q�FrK�b���:�������m3q7����z$x�kz^ ܇�������>��/D�#ڝ%��A�/�Zd��w&�����" ��F��e��o۹�%&��tl�Q8�)�:=(��9��]��̆�;�'9��s���
co�:�Ν3�O��w����<�s�m�Z�%j��aͮ��Y�fr�����ۊ��T*99R�B��54��`@���4N^�概|��w�M����2<4��]�D�WOr��1�N�����	}� �'U\�DP8s��m�DA�Z|X�9�0�!1�6j��JN��y�!K��We�>��I�=)?g#��H|�3Fdcs#Һ�ʂ��S�0D�5�y���f�[fw�<�{���_�);p8�<{N�Y�DI:KB��"��gΆsg_�+�ϦB�ʹ��w���Q������HGP�O���5s�͟=��k�v�^1�[�h�����9E�>֝UB�p�3���:���yU��|bfG�"���I�B���F��$̷������DH>�?��ޘ��:[��^ٙ�D�H� 8c�k�%gE��U�L��.ڝ���|�����Ri \�r#�U���ᚙX4�)(��Z�|��8E�;*��}]���e�WT'K�������������X'4Ge�Ν;zY�2�E�7N�yYP�'O�*BLyuuC84:�X 6�⡦�]Y��0Qp�������[�K�К�#0b�24�,�czwՂ�+w$����	������2r^�"r"-N;�F2p�H�fO
�T�Μ&`m_ɂ){��rea�B��Po}"�W����l�ێ�t�^Y��,
�{g��f=�F����D�>�Mc��֒0�XKY�@�c�> �Ϥ0A�gl�/j��z��K_��d�))m���̟h��A/���Qϐ  ���v�u/���u�Zcw����zb�G5i���v2D:U�Wr�f�����f�9�P}��o�u�ٜ酧�sF°݊9:N�6|f���"��`eI~
�/�C[��KG+˥+f�������#������ӧO�$R�k�������Ӄ9z���R �3}�}φ�A�=H��F�5Rx�(���q�4�*�F�%�kd���=��s�#7}Nj�>�������2'j&�\���i �o�^��gs�Yp����`��@k��E�z�(�,BN�BsQ#	t+��h��P}�md�!��ȃQ��+�(Z���|�N�>���'?�������G@���f~�� @������Y^]r	��
,$��cy�*�Df7�nQ�y7�DZ�h�0I�v� ���&�r��8;��J��@m�I��t��*�t"�-�k
����� ���搳�8����`;̎��:#\ϩol��@F ;��AJn�3ā���a�Q���$
����!4	P%�BG�y���dN)�pp���9levN%����^P����z�9;\�6�Iԭ��6�g#}�W#�0m����d{��,8��gy�|���H��<g�OB*�
��nyK A.3碧Ol�50��� {MQ��EnZ�.H*���cԢ$�r`ݐ�,�,R�L2i>;t"���5Cc� p���SK�#,��$�bڶ}TO�I��Y��̡�r��]�-n�tpJd����9$�ΘW�3�p$�e3[��5��T���Q�$�D�v�Ӭ��
��ea��q&׼�MSbY����([�1�l �!�����a�ўH�q]����]/�W�TT����cn0WRHF?��39,������ʼ>�/3�|a^�a$�lԉ�&��vE��R]H��6���Y;�)Ao��l4&`I��5�0����%	>?�%�J(���'�D���:t
�?h�����e-�@�s�}�L������ㅛ��z#lJ]�M��w ?����뫵�ȁ'%�$��&��Nۉ#1O^2��`�E�&4<6��G?n��,�:�}�bJ�3�A�l�.^�`�΢���6^�ȑ
��}{��|L=}���9Wș����XT�	��h[�'yCu������?�zyP������q�p����[�БC�~�~��0k*�on����QA� �Y��x��N��T����3�B:6�ÞD^}b���f`��Aj��8�d;��D�G���zVމr��N?6T������&W�.R�����r�=Y����|t�T
!�۬������^{U�Q6�&�d�,�������%>SQ�ߠ0'Q�L1���):�'|������_�\?v4<�P���_�QE�֭�Q/�-a��j�_���0�{HrA�p��%�Z�y׫�$���&����`(ȋ�^K#��z�#4����|]7���r���g�n������ 	Ǣ~�VA�E���CJ%y-,�&NHP�F�ـ=� q���Ts�}^\N�Ç�\�)	���������$���{W��xͲ��;-Y���O���|C3��r0��C�_�B$�)�8)Ⱏ>���]U�)�xyd%�`N��?1Ŭ��g���jQ���@���V���Y?���׺P�qrO�eJtW^���9�D4E7�Įي�Q��>��f���	�l�:���b��7���];5���1]��Ǐ�g�b~����p��d�'F���A��'ɶYPn�ܵ5L�zX�lz�n�.��SQ�R�b8�ƶ�ο�Ţľ��޳g_�/�r���gN�E��h��'"Y�0y�+$&}Byn]B��;�"%!X�n|�Y�m�ZL�&s��
u�?�[>#�/���!=�����PJIW�+Ƶ�q��qhǹE�,^w��la���nȫ��&�	q�����~;)L1s�K�ᓶ��	4$��G b<�!�����.d��@/�����m����/.�O>�Ğ�����'�Փ'�#q�ŋ�d�&�~���o���;
O������
��:d���1��F��M�)a�9��0وNR�6'��B.�����T���,1.��D�r�;�J�e7'wMD]�EMAu ����K�VTE�6D��?~�s1�:x |���2	8�=�h�J�D@����5պM�.>��~��脝�gv[��P`&I�-��}����I��Ɉܮ�;�N���@*�'}a��t���f�&ë�N�Aѓwb�cef����rرP��NۃnrB�/���~3f�lDXly��ہ��Г�.bˇ���h�5��:��-����퍜���$�v�صW�D{4��՟.�!f�DowS����M�I6���|qU��g���)��{�7����B�8;0&���K+c����7n
x�}�v�X�]�F��ᣇ�F�D���ů_����RtP�������xX�Ϲt���M3�9�2�7j� B+y{O��@��pk!��AH��t$N�|$m�H -lN]�S[O~��0���*Ӄ�n�`�by��Ji�S�9նO�������.Ӱ^_�d\AT�!Mf�½������UA���EH���ۏu�0{ ��X߾;ܾ�4<zz=����m���V�[{��Ec��N����̈́�v'�7C@��޺uCu�m���-"kFނ�y�-�g<z�<�	W�t3ܴ@Rɍ�A�i/[�Q�O3Z�T&�\cieEEW�6`%"*�Td��Vun�ر-)SC$�3��}֒�O+�����ZOm�E�6'��v4�?&"�ݮ�l��`�Ʒ�rn��U�����7{@	B[�N9� ���D7�چBjj\���r�EB7<��ei��l&��� �{�n(o�;各5ԋύw�1\C��-8�t��q�g���m8���[H$��:����#Nz+Va��Di��"�A�aN�� �
�X�X���^�À)%��*P-�o���W���D�N����Y���IHIt��y��Z����e���^��nW�U�E�Iؘ[wnhc���҃]��?�LC�26R�����H8�-�o�6#�o��������e�h�j�}D�<k	g��@�|���p����gD=S�$zT;U����aˡh@u��n����2�tչ5]�������ʪ֢l���z`��錞�e;�U*�_�7$���Q�%�U���O:� RF�&z�_��6N���S����;$fѩ�1�J<N-��2�!B�������h�-yjy��n�[���ݒ�xl�S�[j-�38����67��>[��(�����ʴ�� �G�{�5Ad]	t ���tG���(¥�����"�̍���l3�������E�t�B�w;����oޕȔ�-x��)$y���>\"�g��$sT`;�v���ł2mg1X�Os:Y�z��B����3@��rc�䤢7jW�Q/~�ĉ02^	�͟z>~��2퉨���1�T�Ep�|l6�Az�ϜSDR��5'Wr�0�I(%�UQ�+<{��Q�J#>?��7{} �M��U�/y�9�N��#�����y�$�N\�����E��7���T�A�_l�N�ܱ}��O��Vv�O��pR<$sF�M�5�]���D�����򻗢��3S/]��k^}2���-X��בk0�IY��_M�`͈�,N�����)��_�5փEP�\��lޞ�.=��jY��P�댳�7 �憳���u(�3N���g��k�:�L�5Q��|�7��-�����Jd���8�83����7i��Q��m	��-,�ں� %u	�>�����J�΄��y?�28�HI��l���������{SϞZT��=>s��L7q3`;%��e"��Um�`!�D�Ad�-��%Ε��8_6I�k�OR��As81a�(?�XP��萸L��Ll5������X	����3Y*,F ^Ƒ�N'�ðpDL,�
���GN����s��_��_�_|>��c-t���o�!��'�.|uS>����D�:yJ'�������>��ɓ�Qi�q�S����O��%	�s瞙���5%J��THĸ�]V��p{���uM����3J�hdtT������j�F� ��K��J�ԤM�\t�
>�~F5�x�Yk��L�{Ԇ\�ć^:`��5$����8���x�:+^YehdT7�b�)=~��#�$-�@_)���Yu	��'h���Q!Ů�>a��4���}J�u���)����*��cz�� 8B��N��������Z�3D��r���P�@�i3c�l
�y��.��Lͳq�œb�!}D�?f��A�x�N�O�(�B�fc�%)bÎ��3g�ʌ��=]n��kJ��^�C�Q���ڬ��8N=�n��Y�c��FQ�b��Ͻ����Tg�gc]��d Ԏl�C'�����'�:����*W@�����C�4A&>�k� j�����+S��,��E�DTZ�ߌ�-�Y#0TZ1'�ɚ�CDȩ~����]_0�F��D� "K>��`�6Z�Ul��Ƌ�2���$@C��� 慲�6%�#���T��X���E�D�;���4},l�sx�,����'N����2�8u�%%o7�|�?�ף$�Yן��|	961�����9aq�ج/��2L��N�)k�X�&�`�|Ms}S���t��lg\*��Dm�I`�-����Bĝ�D��+?�U�k%V�ki��ڕ+������� �HG ���f��TȽ09���ı�c#�]���5,�a0�� �M]�p@�_|&���N�n�-�}�:l'��8�dȝ�s�cx���z�w�9�8fֆ1�,x]n'����ᙙ�;���������
�ю�O��q�u�5C�@��~S�_�'�C�f��qțG�\|u*��[���S^� 8��r����㊝1uȻ���z��6��"�!݄&<���ܚ(��/m\����|1��s�	�g���m�'�S�?aЅ� @�[�n�M�m���/���G}
X"���7�юlv{�����kq���h�I]�7����\c����9L�^Lű���,*�"�a��	?���,y�Nr���Bu�ç�Cr�����oVj@��4�u}}Z�SD�*1�ZQWtG�,[LL��@B���3[���k�6��u�-Zlv3���uK��NI����3p��˯�?�h�|S�@�e˝����g����4��y��M	/M@q�~�P@A	@O=�j�@�lKcJ��}B��K��Mi��\���x��|)�;ک���ީKYdd�#�fÇ�A��� e�T*%?��St��m�L��z��wyO��2W�зnH'��%��p�`�٘s���-���?r$%Ȑ_KG��	y�R�i�qh�V�ʥ�Fm��f&`�چ��ɘ�e��+��ڍ���I�S7箓e7�-(�:�%w����C�?#��Ug�8�C(����m� ��k>��YS��	E����s�$ө��`=|(,;&?�F�ɨƆyO��T�=|6�������-�޺Ɋ6�'i��|���)���Vϝk��`aZ�3�H>�� ���/
Z}ue#\�v]�3zd��?��	3���`�CN�0���e��΁ba�>�E��a�drǤP���2W���P��y��rK��`sS܆5�h����&}��?7e��CՉ�Tf��vi�"$s1bcXra����^��M�9bji[p[����@A�����zѱ����S���5��hF�e��2;�V�3��"��k�Y!�U�o��Z`�m�F,�X�L�d����� �ܳk�mD�,)����������p��U]�};��/g�d=`v���_���G}�l�՗_Ӝ�̓�a6m7�L!�ڴ%�]W�#�h�)�#��Io�HK�xx����x�M���
W�7z	ԁ�t=�fۍ��;��%x�BथK��J ���,-
�:L�x|$X3����9��D�PNk1F-�=���C(�q��s@,�s֘%�_|��}�4�N{��e%�(�1X�ƭP��cZ
[{���:�3��ݻs�e��\ ��#�X�Җ��42<(��i�Y� *�� <��K�y��f�0'�ĹBׯ���UR���O�=뮶�ͪD�2�Q%y�7�L�.ܒU�-8��u"��(��/�xYQ֘c�1�xQ���z��g"r��M=X+U?#�̘*)���^���s�|��m!8xD�S�f��-�4����e�@� ,'l�\�A��ԥ8�O�>���8yB�����R�K���U2�U����)��`3Q���҃G���4��NE�� ���y.�LO����f$��:�Q,*:>mS_��6T)ljV����5���Խ��R���EyGև�A�^v�jG{�F^��C�u^�u�M.�y����^u��99z%�N���e�ˉˡ�r�Rl:���ǎ)˽y��~br�|�}����|4 5N" ��$c�3�r�G����ơ���1��O�(�, �g4"t'2Įiaª�]r�8��-�5~դ���F�D���r�>9t3Z[I�Q� ��;�߫ȊM�Hͅd�iu��Aj]u�J�9@vh���2L?#�x9��&v(��fZzpƚA���j#�֦�*��y��/�l��l�7���*��^��D�	GN�|�QrJ%�@
��*�1�����ko�Y���Ĕ�����@УÃ�Y[[��R��"�w�9�A�s>��/����=f=[���~g���t������,IPt�f[�&bt]u����sջ�c��E��=�ܪ�k�=����b/�r���m �Y~����dZ�R��@�:�@+�.C��)A�������yCv�E��,�+>LѲZ���i���>�ĉ�A�(��(�1�� � lH����U<+'9	�D!I�^}��t�F.6����VW��tr� ��	�ǟ� �'GI�$�"��{4NN�P���7��J�E>�/MiY�e�z��E�'�o�ů�b��wĝ�
jP�C��rG�A�o� 7��Ih�W�i���9-r�2�pZlHB�F@��S+(|Pa0 ����-�K�,�`&�((�p�Yʮ�f6]Z��F��S��@ՀM�Ɔ��X��W���0��W�FScE�#r9&����%`KT<1l�z�[֝�iE̗3������a��?�[�F����O�3�	�è[-U��v�ĈN��l���}z� u��M��S*��P�n|���G��"�80���c���:��`9��|7�Ee�1��bNkқ�+LuLD���Uu�k&�A���g��sr�kHP���r`N$�Ѣ �;C+�SKQ��y
���9X)-�Da�uI��E���CCZ�Uшe�d���q`�8�U*9�����^�̙�D0À�!{I� Շe����a�+�U�(W'XY6_���4=��?~���%�R"�SF�-���'��S/�
?��_h�;@��t�}T�y���Qa`��γh}�9A~�!I���`Y��M-4�8�DzC��Į��k��J
L�E.N7<��%���\[r��	�B���8�d9�\ nVr[�h�SQ�I��E 0�Y�	�Cʯ����U۰��z���{Nk76,n,����ŢK�;r��Ȳx�e]�+�DCw�ݕI�{ϭ8z䨐�!��qiN1�Ʉr�l�����F���Q]��܎!KE�KG��P����F��?_��i/6�Ky�P�o�S	<2v�&$�I�L$��q�iYKz5�x���%M��J���\viml,INT�3s֯��3�1h>�F}��Í;42���n�_:�S��������20	�3SX,�e��� +D�t��Ԍ�!h�@���R��l���"f&Q��	��\R#����3��;�S�p��������8JR� ���fcS�EdAbK��LzTc����� @_����fI�̡�u��CR[�_�����g�7׏䆯�eIy9]������:���l�@�D��pJ4mk7fuyM���r:eNQ��W2�o���]�.#��	���;o��g03>T֯�����аc��rG�. ��OY�8����"6/a� �IF�y������Zn'��z�m�UG�"�Q~�ji���ZCo0���7c��u�|ʁ�#��:Uio�
\ݏ�gFΖ�Hß����+*�0��/xyiJ	���P9���'����a%YQUS���9����ݾ{[������-����&mPj�#�@�X�����Y���8z0�濎�!�Mbt�'�b�l�3��l&��_rrP��[�����8�dR�9߽6X���P���ǲT,���Z��M�U/0ʅ�Q�8��,�9\���i%i$�����">)�؟kݒ�fYhs�l��k��v���kW����ɫ�we�tn�T�j7��?�^�\�r%LM?��BmGC7�#���pFs���?����ܣ�����Y��w�M��9ɑ^vscQ'���Oߞی	8Wml*��ϒ����6��t��.FznV�A�	��Jt��nD�H7��RY�
m��� H�QQ��W�iY@h���o�OY��'�U�P|8���Vo������-|��j�O(�7��F����t�-&:�MNUv�@�;5wZ�N2$�<�\���S)Ü0�N����s* Ҝkv:"�-.�rqA&X5���o�����Ci_#�v=�-7�uÄ�~��/�,�N�)>]��z���&*#�jY��N2���I&�ySX���=���6}����6�:���H�R�-�����o�D@v�>�#{չ�	&���`f
��J�_��OH�Dk�]k����ZS�t�Y��왩]a����mA�f����ٸx$��mW�T��+	�.	k�n�{c���bW��������5!M�Uws�PNѥpoMף�&D���^#m�C[2A�`'� �XRdT���Ke3لj�'�.�� 
;_��-[���Ed�rHem���Pb��a	e�\Լ��p���A9}e�9���jL�g�7P�ry�L�h.b+��RI&bh�����ID�ڨo�_�u��JR�lS��dj��������s]�s�D�O���DQ�ވ"�C�M|�*u'�I�� vK&a��:22	��s1b{CR��=r�`�Z��u�U�WVEY������<�M���l�e���t>��F�[ͨ7�����RR�v�lx����R��	�'�ia�0Oj/��f�e�Pʻ.�CAS�2es6#ysG}���X�S����<�W)+�\]_Sv�4��tjO�s����p{��oc��0������."7+9�������U�|��˗ͬ?R��2��Q���iVh�P~�׷/�b�V���*��O8�A]��9G7���v1ϱ��պ������dםT��i�\��o7����R�Ļ�Ҝ8�UYܻw(���V;�qM'?Ģ;zT�4��`��17�K_)_���b����F��䔍?q�4��֭{2%���5��N߻O>%��w���UR�\���NpP�:�(ʹ��@O������.Bw��Ƌ��<KL@��TL�z1m]U� �h��H/w�����'����������^�jg&�	����#�p*j�7��y͎�A�կ���Dm&�ga�~��߅_��*����?������҄�����{�|����֏?�$|j��O~�S�U�V��;�� 5Bz�$��G�2�i�ic�>%ib%`�#хNǵV���r�=ԉz��t�:-��ShK�V���4&%,� �M[���Q9�Z��~1]@M��w����([�I�["9���W���	��9��8�]w@���r���^_^��y������V�Q,#1΀L�TH�$$�I�~ �r�6e|@����w�:t ��2���E�Y���p٩���x{6�����ѷ���=J?'��$���,��r^�T��l���ɾ!�`1=wsm)��iY��v�Y<N��m�J�8U��	=Y�n�����<I���u������ח��f
Q.��6����h&��CI�$m�s^C����l�/�P�P]���~��H�r��~�-U}V�7r�ڈ_�FN��FZp�e����]�'��w1����s�X����ӽ)��x$H�'��R�^�(���l?�Y�}���@I��/��@�(�|As�]�Q�A�IT�K�������`b���hS���$�,:9�+�����=0��>O�7�8�
a�0%v���������[�o)	��^����� a /��,#���@ȌCT,����lQ����݆u��e��OHW������0�}���0-��=`C'j�'
;�o9u�cJ�=޲U�_P<~��E��w��#�@C�$�hB��y����N+N�ü�W���ܒ@q�%��nN�M�ܴnS%a^�\����^~��-��p��Eoq����@�zXn���J���j�8D��Lݹ};�r�L�|.��/u�����N��k9��eՈ���KϤ�?�ֱ��ș"���ٔ�(f�TU ^fZ�Oӽ�'��j;!Ջ�<ܗ�g�{�媲��(���|#����ʈ!`�v옔i���(YAݾ�bv2uBL��d�����s��~EY}Rm[���)��|_��8LK ��ӧU�Y��VK5�FNI�駟)�z�7�1% !8`�U�K'O��X_o�j�J�vBiJ5�n�q9��8�&	�I~�!T(hx��?���{���h2��Dg���Ӌ��s`{�^b�Ad%�v��4�S��>i�/�p��/6�eƃ����l%�����s:QR]�f{�2'Lg�G?�����&$C�����ً~�{��^x38��=#���__���o��I�p�ԋ>�M��w?PO\%�bI���\^�ЦB�3�}�����>rG�bJ�V�I�ZXjU��V{|Z2�(�F`k+s6�wO�XΠ�qfk����Ǹ:LF�H�:5پB���2���ⱓ5��7e� 3����iF�|LV��S9%^A�_~)�M���揟	����K/��'�oiE�Y��3/�������~�.7�ŅRXx��75c�,b+
؋P�����C�O� ��V��mb���Q5�k��f�� ��q�-������j��� �VO�;�8�\�P�	g3��"S�7�d�F-@}�}PJ�?	��<@�&U�''���ݩ�W8���9�;!{!�%������"۴'��HHb���F��XgK���M�"��?R�șB��@>���C���^W��7��W2vx��肋�9uI�N��R�C1f�W�����U?�]���TQ�(mQI%�VH�z��ܽ�7F�+E��TlۦTB��|���N*��:#��!��8+AuR)� u�fHD�|�ں#KT^��vSQ�z?������a�k+
�Q�~���] &������I�K14j?��T{�9Z�8�S�z����g��TvQ�8���C��ƜECpZ؍MU�}a��c���:@x����j#�Hx��5�t\K�[S�lfJ>ty��Dl�p��:�C�����Q�ᠸM��D��H�%>�lZx"�&�qf�,./��bQX�D���aKQW�M�"�h0a�9�8r��G?��K�ơ~~r�(b���G<,/�9u��C{�|���eY�E�]���w��^�^�ߑ�G��3��*�s���H�ڻ庢MBf�@d�r��0OH�½�Ŀi�@T%�|^��ߙ���Jw܇$�V�A�IIxe��Ռi�C���rkF�FE|M����S��"���T�)K�l%^.��eL87���DD �ON��{v�lb*xH���P�%��0��D9⾵g_1_Gy���^Ӏ)��-V��x�;�9*dd�K����	�i<��k�l���M^��'ԫ=	$x8�Ç�`��D��&���e����P�C8��PFI̥�F;[\'��44�P �
l'׉+z��q�J&|�W�
.��U���p�&@0# ��T���]�0uAc�Е9���q2�y�w�r��q�n���ί�?���Iņ�Mߛ���\�)�4~κ
ȭ�]��\{0��IJE>��u֊�23w��U\H��(	�u�f�lv���=������]z�Y���.��H�����m��"fJ���xs�+��E�J8�I���>�Д��M6F'�2��^@LiC�M���2���PS۶��%Z#���ӏ�W%�lI,���S������zVA��eߢ�6s�-�e`�c�W���P-�:�F6��Q��g�ܵ3LK�oA����~/g�hdx<J}�s$$�_E��;�I=zr��x�}�cfyG�g�@�ݎD5��ԅ���r�T\3x�E���#}�&n��Lےec^<�g��0EÖ�'vO=K��"
��f��?َ�
W��yo��D�@�+�3E��a&jn6L�����B��t����͛a����e�<���lؿwG����~�{Im�>bNxL�٘P*����q��U+�έ+*͜�8�Y&�2�޵�f��������J:�%��9����Xߌ$�^����E�t&�%�Ő���c�ָ����>�.��G��4���])�a��\�7��)-� u�J@���YR���A�\0�kLÚ�%4'�U~�]��0-�M{dr��1U߁t���G����������N���q��s;�y�-����i��%�C�v������ �����1�o���rL7��,��AΔ���aL�軫aA5�-r�C��e�
�m4]e'�<p	�k��O>$�^�g�N5�?a�������,��k��'"�D-{�C���v^$,�����	XkY�X1#
}���*���H�4���S�*b�OK諸�?.{����8�(��g^o�)z����]er�N�8e���Ls��{0Q}�C��Z}QJ�U{gpÜtz>RE�v{ �|T�fʗ?c�9����+^��	�o�~]��%�)16���bÖZ��@��:#�	�1�a��� ��Iv�5�@y�Ŕ��%����[p 1asߠ�[�����J�q�U������F	4 n�ޔd)?���.�ѵ�~��0I�v=��?����y�o'���6��
�Tp�7L��;�{�*��C��т&� LG^�m+H�x�gL��\37����b�k�ԉćy��)�]'Ά�~V�6�����m��nB��3 ��P/ǱJ�R�y3-8pgڌ�@��N[�����$B�T	V���f�`m
DVA��b'���ڭq��N좹0rUy�#GN�5�s�ݵӿW_�g�妏�qFS�#��*[g���*�W�f���7l7 �nL�=#��c��l�����b���x��,���|�,���Oj9���զ]�o���Аw4~�}q�d�����Ǖtj�%ѐ��!WD�
{���
:"�O�!]�4��i��3�hAf�9q�`�a }>���|u:i1�b��H�)nd�5��Rš�0ag�`��,��ȏ�hutG2�h��'3.���}.���}^;j��k�9�cAQ����>V�aU�Y[tiUU%��a"ء�3�XJAUI1�-�ګ*w;"=�|4�v�f��N=��$Yu�ےy*�ʒU'�I!_,�ה�B�z]?�%��1�q�uM�GI��ʶp�a�@�0�q����}-������E�p�]o�,�VPBa�XL4��j2�э8'�&�k038qrߖs�0�ֽ�A���vn$u�~��,��J�`��E�q"�,0��wM�p�?$�$��k^*J�[��z�%*E�7�+�5�z8G8\,9_5�y���I,��n�W���Ph�pɖJ��O+b򩨼&v��ح�� E�_؂#A�Q�ϱ���ۅ~I�kYԖ��6����F����s� 3	X��V���Ƶ���Ʊc�*(�r�}Q�=U�ڣ�eͤMckzJ����5���󨹞|﷼y��U�Ai�q�FP�"s56/�ї�Jݳ!~&��[X��qt^W]<gj�~�����!�ނ��I$�Į�3;�W��^ɚ�'T<%Md���9	ɩ��OL�wT9ئ�`���6Re�����t#�伉�&�m����:]r�2"��#�qUDnc�Iar��;�Xl�G�
Ж�A��c=HH��xN~ :��lꅾ���rxj�	������i��pG~��Y����l��X���a`F4��re�D��d�� � s(�(]t%7���M'�p���_=��P*���Q��A�쨏K���]S���Y���B7'��ԅ7��x�M�}�v�T3$���z�	�ygmq����I*щ�a����HK����lܸ�GG@�.H�z���kɊ�<%SRb�4�#���t\�QH�\1,Uk�Y���N[���ZW!�qe拾Iy0�����0��zQS��$?|�3��z8� ��\6P�zh[�>�J��Bbf�T�qf�$�{q�mjw�|�چ��,�c�-�u&���4�ޮf�],��H|��$|kB�D��Ej�z�h�~��f���
��v�W.	яo�#DP1v����VÌyE�>���ؐ��>��D!��3��f8Ô��-U�&�_� ('��5�:\�.��X� �5n7�
���F�9���8p�*��\6D"��G��y}���eͱ3R���2��Q��X7�7�������m|W��3���O���إ����E}2+������mA��a�:N�p����Ӊ�y}��!��Q+%�,{Ϟ�"=��/k�`}mY;�T�e�;��Jߠ� �>&����k}��7�����IQ�j3�c�rg��� ��@��dm.�U�Π�C$��F�-.�(-��u.WTU�pؘ7�3a�cAx_����!�O?���r��v��`G�݌�j7���gX��K���L���̖CT�KPFUޮ��-.��,(��f���\V�fc}E�DQ��SU=�m!Acqv��f��=Q]��C��.?����AC��p��Q�;MM=Q����K�$WA��
1*6�R����y���&	��;��>mV���5����&`b��`��i1Vͯ��5�����k!�2N\�`8�p�;�CV�	>�^Kf�6Dq�G� ;�}�~��{$BU"H����\*��  @L��5)�#G�)z���)���â%u׮|���w��n�i{j���L�K���	@b��-������ͅ�=���8|W���LՄ���>�(�U>��Z뉩���7��@�KP��8?փ��W����y������u��'	����ߢn���u�@��^��ֆh~!�C1d�f+YtL�݈��{w͎�*�����^
��a(%L���G���}��_U��"�LN7��K'�*}f����kN04J$����Kd\�Si��3�=�a9�:}�j�d�!���>x(�%��v�w�K+�!qJ1}v�=ñS���QW�F�e�>׎�X��J���	-��e7��;����E�%Y������Sw��Llo:�V�C��J��5.�)j�0?|_�@E�L��H'KGprl�����+4m$N�
����zU����>o�RиY
�h�v�Nq��!_[���y�Q��M��YELc�*>��Q��f

:p���2�� 6�@$m~o}Ӊl:���MY����� i��o�m���9fn�ڦ��������75��)L"+j[�5R����:}l5N\��ƾ�Q�n6����[�M�X۰��:�& u�O/E,���4�9��@�0�FՕ���O���/���ߔ��VTt�G��e�(��1]U	�Ͼ"�=��b|bW�l}�r� �
}f�Ɯ6)�3~����V�s���N }��Y�5"a��^-�W��p����e�Z��l�t#��S]ZD!,�/h�}G�����_�W�#�Z9D����	�G��8uV,�]�n�ە狉0p°$P��c;�'����.�ױ|���=�v}�k�Veo�dDX�vΓ��$���{���ҥ�4{��%�%�c��Աѷ��
׮^�ii�/���X���cH^SK9��_��ZUdH.E~ѵ��42,�<�������@K��H(�P���C,_�P-�a(��Ą6�*��6O�(��#P�H�V�#"WR�J
��etI���o�q�0W����5ۉ#�Ţ���y�~�b҂#aa� �PrdN���i^
n�|Q�8�����3ܹsWa-��ӥ��D��F��[(��8��ͺ"����M�i��!�L����JvM���UZ��0��>�\QD�>s^����n���xO���gR��ϋXC	"��:�ŶY�d�H��B����T�,�&�x��|!�td"�vU�vM���BمX�2,�=n��6U���^�[�_T��B� ��b����kX3W��y�E)�:E��Y��X �ʊ��9I��SU�+
BR5�Rc❧���Ui��PZ�E��<G�oE(�@B�I��@�
���9����~ex�>:�Q`@�:��vSxF�/�LhL�"�m$cw��Fe���^7J�#a:�d��t����ĭp���ܸf�,�h8�	�@hǦ	��|�H.
��T��-��nz���x1��H	&�cu-����	ϳ&���8L#����N��SO��d������=r�Bg�PH�N�0���WW���:�kɬA���e��g'��\�DA���1�k/4��s9��I��ŭeϿ�n:�I�'O*&=��зRЍ��vT��i�����H�NH����݊�<��ڑ��I�c�XK�+�[Jђ�Ƕ���x9G��A�3xy�j�n��)���?8v���˱@y�ĉ�01���m�: $�� #0�(R�>}��%'6��:^e޽kG��=ba9yLqW��`��#�v���a�f�M����X6��;U"�|��+��B�B��\����3
����R�^��%mÌ�N����w����|���'�w"�g�_�ue�~��^�������-ju�V��خ�(n�_^����Ț���ɉp��I�(k�������^9|����o���G�a���=���?�X�num%�o�'GDg�~뼝�R��/��r�{**�=󲸹|�5<nܸ.^��h�rN7C�Dw��q�ɪ��-�K��������z�~���4�WA�����	�ץ��t�ժ_N�ƀb��E�}��uy����M$>z����#�ѳk/&Q��yHj@��;͎N�өGfg;�MG��r=�7<2n޺!24����>���~�;oi���
���$�#)�0���	Kbɑ<�/�`Bln2���\W�_��v �ȥ|��k:DT `����@t��@��=�V�y�@S����PӴ֢�^�g�A��EK%	��umH"
��Ԯ!Nkt� �%�gfZ�<_��r�┱!| ��wd����@́V�}��������d-(�=����}���~�M����R~������aZt�nؕ�������s����߻�|�M�������ۚ���Er�?�(�@�D�ލaP�������pY����]���\AA]IG#V��4�fӧ��4�5�̳R���e�G��vR�^�.Ay���q�Û�e+��f��A��>%?�(���)��Μ^�N;u,2~G��^����cGUf (X�fYs�#���}�yط�	��|Y�l��Uk~>C2�dƥK��V�o�y��-5���D�:u-���1C��a8���v�IQ���H�P����&Q	���	h�Tf_�{=~�Ă��g��f�Du��r+<���Q��'�lIб#�^ީ�;��Z�}ϔ`��z�RȲ�?`:�@�_׃q��q������j]�?3��ˢ+nU�K�.
E��3B_��@����l�gs��#	%��V��R3�Dg�UVA߄S/yX*����!~�{�W���_�*�M�ץ�������+{�<�b%6�9a����TM*�p��FF���A��a���-���cGZt�����Bᆶ��;͎3��\���E�ĩ'4���eqv��쑠q�=f_�]
����>*?�g�$M���O�,s����̂�5@�L�D8���oh<m���U��1j���`7��@�� ��B%����d�ͣ9�ɓH�:WV�ڃ�h@4�d\�Ň~(�`�=$��Bi]7K�e����գ�#+7?��3�Ȱ��~١�I	��+Hd�\!,!��*@`,!b����p�5�K��zGH@�!���b�B1\w����d���hqi�B����ڈ���A����7�Uc�!OX�n�}yI��g���A�p�oݺ����B�5!�L��~n&�	^*�2��L
s�m�T}�l]`��0O"f �r���;��b$�N���2I�KB��,n�c���Jt-����\G3bg1?t�ঢ���`?��Ca��]�����?�vP�'���[?���T��~���1�d��OW�/~���#h��+8�����P�O{D�����
Oũh�A��{@{���r��>�B�Åz���9N{tdL_���%w���y��s��O��t��m9�5��%��/�H�F~�RO���]Z��G�P�Dtm�գx��/�d�+���&�)�.;4\�Qݙ�sϦ5=D�y�bx�J3�O��ap��GO�����M�Mq����O�D8���̎؅m��s�Th:�5-_ea$�O6�Z]
��!M�I�6��ۉ"��)��c,	��U�Ǭ��>��|�S���4��<"/�m�k�B^�K$��e�f|#�;���k&Ae��)�4#E,7�AD�)��D�m���]+�3s�,Sm��� �����g�Qs���'>G� BM9]��-� l�#� ��֮�Cɵ�W!DG�%)!�~�X���v&�(�Sl;���,	Q��5�k���A�p�fS��Zw���QQu����#6�|F�60$mD#�b��@ 8Q�V�Q�ٚ�+p�1W����AY*L#K%�ܧ��r~�G݈�Y��#ݸC�:.Y�s�Nԏ�nPK�Hԇ��R���x����]�ѣ{��ݹs\}|�J
�`��*��8a%~dfv.<�'8x����p�tI-؊J-M1Ul��!ۆJa�n�&���}���325�ܾ}K4���gG��Q�l�h>�N���p8����H�Ӱ�G앳�q�l�O/��']�X8[I�P=�֗�B��mVQ�2�u Q��0�*��o�
�]y�1�Qm�⌸�Ԥ��xS���Y�#�hayi^W]��;«�^���N?����N/���֞����n	'��1�|�;����4?���f��5	�6��Ս�(g�C�ڟ>y��A��?��L$]K���͈!���i<y�޹�o~�����'��i.�q�L�_�n�*-Uz	퉈�>h��t�V���(�CwޒLƩr�<��LDa� �"��� gzfJ>��M�W����q��e����?p0?�9�D�]"ŶL�!$cӰt�>�h�>�����pТ)"�n��3�T?�geD��n۶�p��~����|�j7Ys��eS
IY�?Y6��{ vڸQO����е#����d��mgϝs���p#��)��I�{瞝�k��K�u8��h��á��p�q���eQ�Ty�uex@#:?�CQ*��a5����p�Wg	���O�)�EU�=R�A�jI��KN��Үs*gf��t�}�m�x;�F�A�'�|cr�v��$<�LG�A[����ǎH+?���������(VR�������mρ����͆v�@�����0��f��~
?FYg���Ӛ s��Q��f�&�(�l�]�&�����)DE�0��	�t�|����C2�����CR����8a5��;NO?��Y���$��<����������&�T-�GƠ������*���L&�2/xPW�Av+n�{B��|E{��V��q"�u�P��5-T���z(R:՛Np��h>�M���}>�t��y�|lܼ��%Q����͛�����;&�������ɨ�t��U�0`��3���*���G?P���ǟ
�J$�ĕ�Q���mc����^G!��bU:AM&���t��v�S��LQ�E���/4����G�`)�)��Ȇr
>x<����X\>߶�zY���Ν�Lb��0d-�ܝ;w��8(�^=�%�����ǁ��yX[��K ��U�~����pއV09�$��n�7�9��>>7���k�n����ۑ��ԩS�F�շ��������z�r�){�=2�T�Y�%��ej��h�0rV���L�q �	>�wfR9P�u#�'%~]�1�-,����,y��'N(<DP�����e&-�%88`6z����%L���in�yx���e���g¹s��-X�I��Ѿ�s�Ϻ~�9�q3���80h�}媅ާ�o� +��NVN�
_4鰙���~G&�\�}�%���ޅh��={��0N�o����ݻ�����h��r����M�8� ��U#�rA>��$i�V�V��2�Lt�lF!o�����S��O�&���+)Ab��g/ �j'�t��n*!I"x���~��_����f����1:y�X@���՛ͷϣH����fԪ��k�n�kd�ν��Y�$7��� _|�m�AM�޿W�I�Dd����ѱ�鍚�Ub�5�l�e�1�u�D$��]A�C*嬦SSs��T��C��#)����o�L��ݓj�5[=Z��%��&��%�[�=�Wg��DF&�Q2�!�t鶦|G����qs��
��m��֛*�(�ܾu3ܲh��#)�0)u{i^� �&�&tE�:L\���N:|��Ө�\R���!�Pb�5l�IaN�� �lzf6|bQ���)�gQ��0\����&(�r:<x��մȵZ����y��GT*a���}�4�����_r]ٕ��	�$@�,��R�L/�4���^3�]�dk���V���r,��b����3û9�}�}	����23��{��{�>�,�!~��������{��]sE�E���df�Ʋ<�n���Jg����C�'�����4ڼ���|FzW� ��� R~k{W����
��0�c��掤�i	,�3!,������e�2:tK�YA=������4g��T
�<����81]�?R���i�3��!� �f�\�v��5]\�z��:��%Q�!p�/��_�|�؊ך�R�Y�tk�� 	��t'��J58dr'A��K��=����,���Dw�E�e'&�U�҈긑����YU�v�j� d�-J��B�)�0�LJ�P�9*\sC�avv;�����KN�"�����I�?�F�=���z;��R�'�	.
$Ԝ�����{]u�j�S����0DgX�Y��:]����ú2˻���|�k*�c�9I"�)W$�����ի��4������- 98�׿e�%܃���=I<zA4����>,W؄<�])�bJ��a��-<�b�Ç��5T�9:N�1�N'� �����-�X�����Y�Y�=�@�+��sR4�3�nwnC'h&#�)�ć�Ӎ�[��}��@�։V|öi���CO�>�v��Sjdww���S3�d��n�[#����"SQ�gICÖ�Z\Wi:h�|Z�H�_8RC���jz[�\ ý�8T��T<m�d
�LK�d��"�7�uv�-�&�u������8ڑxf��ƿAr�J���u��cIg9z�4�T*,�dyɁ55���, �����+�{��%Ye��[��~֝F(�y9*�M�KPWl�����	7��v�"B����/�������L@3-�P��sQ^(���Z���ͩ��ɳ-u��$G�]��Q^LpS�D�㇗D2g�t|c�����2�șs(fіz��A'�GH`q[Z�����	��+�gԂ��7�N��WFJ�Ý�	�����'��Fu�t́ ��1!� 3�J�SF��pp?M����- ��<?��k�u¹	��(A]eOk�#9��X�Q��MP�Ѥ�{1R ����c2P;�X�A�wFN�c��s:�nʓ�{ӾF�L��*U:���������1Kd��͛±���[[���7k��
�k'[�!��Ym�+�+�;�,U��?��2-�ڤ�|^
ϓ��jMҏxgfJ�����iNCj
�@��ϗu�ZШ�@���'E��*M�u���L5>����i.Py���43�;R]>Q�Ѵ m����.N���;>s�d+�ֿwv��0�dhH��!��D���ډ��$+��4�����N�6��{�1�̬�Q�H���ɉpsZ�ۍ�k�ye��E�d�	�W�>�:���U��vt�!:0��8e�M@��sa�iRWi��ө������P��]x��Y-�� (.���X�(UC!�jgcSI<��4���8�E��g�ϴ�<<w�0���aWղ��9i��xp��l1 �<�=����E/Q?�����G%=ά!9,m����LR�u�Q;q�C�S�`������B����eWmxE%��Om�u���E�z^���B>|�@�F��A,�Q�N/ڱ;�����:���K�.k-p��ZE��˶)�� �b�},uU�1f�hr'c1� ���gH���g>R��E��}���AƭVUQ��[�qL��s3ke'���N�d�c��3D�M�i�`nZToΚ����Z�=;9Ͳy4�>}Zt�;5=�%�*ʩ���>3wA�׎(��z�RKl:�U\b�Lp��$4��[����X�T\_��G� ���?p�$��h׵�h���T.g�XG��G�88��}y#�4�sbw�i��%�Ƀ��^���ÚT���N�R����ݒ1a�¤�T	4�a¼�f��C:f�"���iF�Q2&2���;|���֨�z��{�a�����]un�i� ���.�*C�<�RPwxK�T����-:Rme%P��j �	�	�Z�̣E}GE=�=o"�zАj��[4�d�'O�V}^�����CAZ<��d��H��^F���]�ˡZ
��zx5n���y9���q??r0�J��ŷN�n�T���鍜%yqxo�w"\�xᬮ�e*�9,l ���	=�|�;wa4�an4�P2_���ɗ�E/Ϳ2o���eUKlAP��Q�J�n�B�XCt$��ak|���]��� ����'������bS�y�a�cq <���0Hy�8�?~��2���mJ�A��g4���t>]�~M fH(�޿{Ӥ`�>|��@ې�s�8VM߁�GzJW���2i��6����鿿25����W�\�u<�o�S'�K-��Z\�S-c0����8��(�˻�ڛ{x�&^�=r�ד��+;Tɸ�R�$������q�Ą%y}$_���:Ԑ�`"��$Fq3�$4�&�y����B���	9B��u�9x��4��VP(��IpP��)�h���i"�@l��G���~�$����:�O�~�E!�?�㧺��?�Y�|劣�5���Z7�w�r�Z�B��?���C�<�8=�Ϝ.�g�-��q.`�U��(�q���ݰ���3�tFy���+!0�-o��A�����u�A B�4�R�MJ�G���QC1L�������f����R�#�i*J��{�<��)u������zn���7�H������X�a@h�I�o2�m�j�{�����
��T����A�ӤTN����^���%-��'r��>�T�2���@���Ғs���a�x�G>o�B�q�I}h��� �M��8�Q�o6�9�6�3�qU��Dۈ��F��k�򸊊��H�:�?w�t��-ϵL�j�ʜ&D���:C�� [�+��^7�x%�Z�g�%�+J*?y*�^ߔz!���:����1��E$���_�2��+�D�'Meb���!o����Q_H_~��l	��"}�F�S�ɜWW�*K�{��Fy%��b`%?KA��.�*�y*�tO���n����pҚ��6���rL�� ��U��<EN³ @��~�j뵸����𖧑"(�4ۨϧ�>�P:�l�Y;��$�����gSǌ���M㫇����� վn���ɟB�}�&�ל͂���xn~Ʉ஦�ANP�͘p�B��fWQ�}8��y����~�^we�U�u��!\sa4r�X2ߢ���X�9�|.բs��|l+ϺzvU�C�Ɂ��>�N�����c�EA�G��`x� �[�<Bb8�=w������v����7B�`7�Wr�.\8/�9P��`��\}�)g�����;i{���Ѥd��\:t��E��hͧ�������^��4�� �o~����{�p��t��C%0�׫��m�����m��4�WR�#��O�<
��K��=-8����6�x�&PR�t��w��c��C'�'UC�� ��s��7���RI
 ˥�?𸊖65@��hʅ�UY�ޘ��I0���G��ePAp�����>-Bx�����Ͽn	��ͷNbO]���	��+��!0�Mf��=x�*�F:p�pzi�ɖ����Pc#V1�"=�l��Ի��e�nܸfц
E�/��Z%Yrc9S]	9�:�sT 2�T��P��ʽ}��Q�6�7���P*�b�M�ۂA������P��P�f���`��E!>�ۛ�>�*�E�����7�5�g΀V�k0{J� �SP{Ϟ��hϴ�������{AB�d��4�����=M[p�X�)� ��w�9SO��p��Ӂc���%4�9м�~�y�@̃�+_�Y#�>�s#Wu��kR�J�����Zuqy�*�>�IZ=�,���NTS�F�^G����y� gw����b���#i#�y1t/��m�*�-,B�H�+�,���{�ʝ��B[<
uQ)Y��5�2:�>?g���IArqY�p|
Xإw�~G�d��߉��R>x���.�%d��AC�j����@�X?u2W�`��F���Z���^7`�I���5����Q�����`�+@n��vp(>w��ʕ��0���a�xgNM~N$12����u�Fإ���;J���)W�	?���'K��������(��
�F�(������R�E��(l`�',v �B{3�?�7iZ�͓�i�.�&��`��NJ���b���0�CY
�ջ�&o���5�g�8RxD��7�|��B27�K�Z��A���1;lY � ��W�f���v-hQy�� H��-b�ZKS���I	�N� 1)�Gs��K th��v��Z�53���H9��������G�ff@{���U���YEJ)�v�3��jj&��&�MPȀa"��|�K���{��^�d��Rqm���y�{�ܥ���Ȼ��P-����J/;�S�k	�\v�.*�/�F���^����l)§\�~t�沩 ٜ&��L�F��r s^��y�UE˵�EF��8%��#��tp���}^�p-m�?ƚ�,��3������@/�FPpHK�I&�ϐJ��H)E,6C�p�� @�Ũ*�l���=��A]C��ӷ�&pN��Qvjԧ����$�����M߈�t� �����Z8	��g?��a����a}𣫚,���c��@�#8?�����a��@�Esj.���YQe�c��^g�4�q�PoL9�F��81��?�x	OAgm�r&Q��<)�w�f��*�3�>z�kߒg���E
Q,6��;��G�Y�ݶ�L2���7��	�9��;�\T���Gu������1��_��|~�ڽ���.ؾR8͙�����Ϊwc2��K�k��;�������'I���3>S��;r�ŷ�%G �!�AA �OMz��3A�/�-(�_b�������(k��y���N1�(佉=�mҚ�fZ�AB�B]9�	�Wu���d�8�Jk�][��3�"�2I��i��u�4�|+mm�� �-������<�v�,�8<�Ξ?������ǏS�>g}{[��/"�1�淿��G�s�b��n�K�|B��I>�՘K���Ry�,��vlmt�`��_z�C�Jy�:U��r�����N�(����U�0�JG��ύ������OjyR�*��52@͙.�g�^˛z��W�k� ��1���%Z��Ղ�`H`{@��b���%ҿ�h�TV��R�6��J4���UQ��!������i"�o��Ƽ�gf�ү��o ]O��������:�hK���μ{* !D�À��e�I&R�n������n|^�N�O ���c%:�������/ҷ����?��2�7�<ely��-xF�W���?�v�!�f8 mpH���cAXkb2u��Oݜ ��͠%g0���T$,_�Fx���x$G���16�c��~S�D�^wX?s�H>�Ac_�-��P0�T�gL�L�VK�Dm�5����ҕ+�r������b�94�פ��T��^?����	 T#�:z�D�[p��g����t���>n�������β�&�K�P�����f2Q�\��#'�����������,1dj�sY�<�D���uA�V����X�}}P�d�������*��.���
�+R��5uO��ǰ�w&һxP���I�܁����>;���MSߧ���_J�����=Rv����\��'ω5�v9J��yEp��*�ؼ b`;����z��ͨ�@1x��eע�/t
4��l�|�����m!��	���ٿ���Q'����ש�f.�A�!��-,��;fO��sWϹ����ډ���Q�9e_H,�c5�LE����!��n���؈]|r��NE�O�A��s]e���(�H.�sjC���H,��G���0�ZH�
�Qѥ����W�
=��@n����m0�χ�����єk�t,,�f���C�1!:{)�Ŏ���L%x���-�.ᇙ^@j���`?
N�q�G�ş��Xe�J��#n�����e#�պ����2ȸ2�|�!���%����I�A�?gB |	A����
(iq�{Z<n��7Ŕkl�F��IE1�$3�yl�墿���Q��3�x�R5
Z4UsH[q�S�f��B~���I�U��.n��^,���H�*�c��A׮gB��M�ꌄ��$�8,��Z��x:Vnj0���Ъ:�ȞR�lssc^c��4A�G�7����$͈eG�!v�+W�����w����C�uĂ��R�"#Վpp Z\}��߼y���I�W)ЉD�<���>�j��y��^��w:�>�L ��Qڣ���;�4�|ڎ�k��z%������n^���e�M�7�7�B�)�����n�;>	Ȁ�e������7w�߰*��L*��ֆv��2��.[�#Gh.䜰YTL��t�'�>?� FVE��u�q ���(1��4�x�m�2�b_kR�Dd	�ɚ�¦���L� ���/� ��J���PΫv�-�A��J��^�ҧ�\.��y�ˏvZ�� Xc|6����L�0u������?��f`o�5m6��	[\z[�Q�	`g��T�F�v�܊���H}�6�����4{Й�Z35Mək�����R�(�B�&�NQ'Z�*�����X�F�q���- �&�G����>rH�]{s���)��1ԣ9>ǤݸqK��������������0����eknK�5���zѬ#�^�+��t���?�m�h9(�}KAY��U�Pܙ3'-8�-m`Q񻪝������Q�z��)g�t�\�� �y��9�L`�Á�u�3Ft�T�;w�t/�q\�O?�4���h�u�'�t4��W��4�X��s��Qe���no�mkNȥKu�X`��/]zG�I�>}d��"@�m�_N������~��i����;{F���<�;�p��^��?T��kL�͌ax��J[b���+�����z�X�u0t��Oc[Ї
���k+����=3����C*RW�_~�5Ҁ<r��R�P�rTq{i�سr`)����Q�Ǌ3�r� c��w�E|���qɧw#���	9}�zQ��P��6U0I]P�!9��_}`��A�H�B����5{������ 3���!2�������l�M�'.=z\ �O?��l�ց<��8z�l �I����v3�o�G�8:�ߩ��`��bK�g�o�n�������	lc��抖J#���đ~ДΝ=����C��9��H
b&U���x��� ��h[���x���;�˩��N�m�߿�n�v��s�&�Fx�Y]�q
I��1���'���8�~�+��]���9	d*[Ї��fP�C����?N'N�Jx��n	܁���	,W�}I�kb;Nۊm��n;�6|p�x4. �E�a)��qI��\��'A�1Ѝ�a�X�n�HO�<�I;����N�dd���I�c�f�>�/�".�qzbj�bxYT��c��}�����?�ې��E��~�P�fFNMވ��H,W\_�{Ho|g�x�Q��	_�|����b�I�CZY��J���c'<;~���[`��#�8��<:�M:�D*	F���X�(ஔ�q?(P�ݩ��)6��9��a�4�Lʝ�_�i�v_�H�"�ƌ�?����W�1ޱS����//��@K��4�D�[����խ;߇+</)%�%�c^mÄCS��T��\Ť����wӣ���w�iz���J]�����/�'M���)�0�3�e���Z�)�8�z�!��u��4}�6ֶ�����Z�����E�k�+%���qI1]��m	���M���p:��ʈ�j%��1gC9��I�K�LN�>�,���O�v�'�ǈn;굻�Ŭ@��Q�/�������sH�:~��'���E�� �)	���uy/gO��j#�Y͹�5Z�!O�ۻ��:|{R.dY����Mu��,+��W���>��3�isc�N�s9�^����#J�3�� t�ѮC}��@5�r��sQ�4����A/�dr�zE&?�O��&����T������GS���S�z�ۢ�`-�JD��i�k*洮����� ��3[p!����Ddf1�Җ~�6jdj౽���dF��$�};�R_t�פ������3r���n�{��Z3���5�+"��,�ᘼ\Sj���띳���Y�n�O=~�T�\�v��$X͛�Y��B�Gb���|�4�J����GՐEv+���>wؔ�X���\���)E��ݤ��@m\�I��X�[R7-�cIP��޽�F�A8����5�W��1�{ocہh�&}v�jOX��,�JqH������ǿ����ߧ{�t��{J�|��ע��VQ�8h�/@�����:j�ц�$9:��`�ٌs�U�+�&.-v��嫊qn޸)8�'�jJ�����ϨY�)�X7l�w�}��}"�B���'���R/�ߚ|x�"������f57|EY�=5]z�:�lSp�]�%[�.]���]�6큔7wr�)@h�k�d2o���W2�$������4S21/�������,7��~à`�� �X^�K��.�ZX������<�/S�<����v�}�F���mKMΈ8�.�>FZ��PF�1��d�G;s�IhU��6�����Du6�4~�QMm�o-,18�����\�=��N���*�2ZYiҸ�a�i��{#�F�$�����y�>�P�%x�3�Q�����jw�N0��a-�H՜��5�E8\ֱ�B�o꫻�T�K*s��Y���Y�������1նϙ�h�u:~b��¡t�Ԫ�>�������J�Ƶb��5�[��a����j���qM�c�h��6�۔m%=g[��~�J��gϺi�U�)[��'RN��x����lH��@�>��{
SJD�JG��O����H=����4DQS���e(>o�$�읶(@t��S��d~��(1T&-�!�1�	/�葚c �w��yE��fVS\"��Κ6��\Р���J�ʼ�]ض�����ɳ�=� Mel�������pц�hkTT!{�(��{�*�Ǐ=���,j�͟�u�uv�H�T?�80�j{�#uǿA�$��)s�!E D�6��	? ����M�ĀEb`�Y]P�4P�? ����W"@�X_e,��ٞ���=�_�*�C^nTR�����WX2��i��4����9yc��t7�����7�w�6���U�:P���T_�ISS��N��a�`��rDi���m!G|ښ�.�[ڣ����H��
4�B�����&5�ܦ:}1m5�E�?����ZP�<���B���$!K!�͍ϙi�&����6�����������r5�˭���O׵!&��գ����%E��^���L8"����k����Z�զ��p�h�����YP5yp���MgO���tcc[�;���8l���lP[}�=��#aٔ�U�M�T?q�~۽Gث�ǩ�D6B�8{ޖ&D$�!��w�&�J&x��F��ؑ�}Q�W�~������s��j��K��ao���i�3y#�K鑟Q�@���Y\F3Ȼ�H߅�_�᪌=���+t���%z�RI���)��^u�z��6��ѭM��S�HX��I��T�K;����w��[�ӘS���,;bA�nE��c����S�Xj�;P'�w��b��~p��  zIDAT���YZ���$6�L�#��5;@�}E@;����i؟����Grm�@N��[�aR��=�l�Dڨh](����3+��G�0<�z�Gt��!��7�_	��hx����;ҟ�-o��V�Vb����Rr�k�~��rZ��ZԐ���P�Am~8�ʦ�^4b�~���������#	OC�ۺ'@�4�(p��w84A�w��B��n���.�J�a伺1a���醴/^�N�j������������kgX������5����n�8��)�K9����{��M���ǋ�)��T�9��PW�#G	 ;��4ov:v��V������H}i�l�g�r�uw��z�l���'ц�4a@m� �i?��lC���\`N�������_��A"2[dی1���@�,^׫W�>Bv�5��6����-�_?�MY�^͌�e��(ݾ}Cx�a� �j�P2���v?��یy���,�L��������<Y��)j����SD�w,��w�Պ�YaԳAW|�ŒJt�Vb�B��V����K�
���>������w۞X���P�T,�5�uWEy�H3�;�H;�LOhzz�
\Ռ�{&�/�Zէ���}�;�ҩ��+p��O�T0G` �Ra��qyx�\����j>T�t��
�vwwSu:�Hy�2ϋ	��s'Sg�v��;������~8�Ǐ�ɀ�������hJ����'������V�L/�h��C������ZFq�Ng3h��m?�yT�*otb��d����]�w}t^�6�no#����N�3��f�Gl�$?~�6vQ��ܒS�ɾC����gO���)� H���!��J]���ޯ����t�ѭ�3��{��/v5L[�����{�呶4/˄�?J�ע�S˝m2	M��c��L=&����Rr>M�}�u�X$�������gD[����*�U0Eӣy��t5鳬��}g��NoWE�cսb��Euq��D��(T��z�aߋٲ$�f�gt��+���#]�Ce���V�H
�gd`ɤ���+��6S���$�3A|�)UK8��[��>,��p��$�Мۺ<,�h���9��y�N,���*�Z#8_��D(z��U�{�H�'�hK�jA��o�6g�NǊ蕐(�%A��|�r���<���SwFR/�VM��, ���f�ˠۨ9��O�)�`?(���1����^�d�	s^��U��`�����N�t�WD�v?�Q5l1���m�oj���b��ʪa_�:o_���(�1!��?(�\�<R�U�Pɤ�jF�+��]2f'%-�^tQ�7�/9��:��7f$���E$��}��|p�[���aPIN���'��N����g�$j6mdGEj��\WxZ�H�^z��"lo���́8�;E�ԛ-G:�� p��(S�1��$G�,��C��Ҥ���9a5&��嫴t`�;�*S��[���P`�Hɐtur4�~���NV-`�]
��Y�}���lorjO^�1D�'���in�~g*���rzl���[����<҇X^��I���`(�o1\�{ΏB� �%���nG	M��"v��~NК�k�.ܖ�U�QD�^95�`[�@�r__����aT���܏%#���B��D���E�R�t��ܗ�'��Ȇ�)\!8L��e�����v�\�!�>�'Ͼ�ܿ�e�8�&�6d�w��z��źs!��EM���Q*�3�ӀB��n1�(���^
S���t� �{��Ն�)�*�[.;G�;�hދ�P�ks� *`SX�A��asZ8�n�T�7�l ���#y}�v_P��_{���]?)E��5M���-xug�����^�$��M@Y����N�EN�<�R9xq������?R�gb��q����>��M��Inc�!H�/�x�����&*�==���'����|-C�L���gO�)��G��>NZ�#L������]�ا�$��G��tK&����-���f�;� ���;��U����q?7.�Ո��Iwx����HX�q0��f�'�`�����5#�U��99�t���rn߾��?tp!�%�0J���,z�����F��j��!��#NXt�Xx82��ʞ�?����?�/�����7���)����i,\ۼ ��c���E.�ni)���>"�Lqu�k1UC��N!J�@�����|h��i �b6��`1N9��MԌ�Pc�:����_�rrl���*C ��ş<{�,��dy�`���-���Q���BT'�X�"�jq���1̌?��d�1XL¤d{�RJ���O���?��)9F�ŗ�����1�S�����ܑ�C�3 ��SȢ�a���~��݇ϴ��(��(������U����(<�˵�4�l�ӠIG~��w��1��YP|k��꨻Z����5?���Ӵ_�m�q��O_lo�&A�pvx.��ǎ�P/.��$������$[�8Y�4a��)c��}LEY�GT]�v��BJ�p$�G�țM�@@v|�=�Q$����ZzB�#�0j�G��<�a��8Y����$Ѹ����ple�8�Ɇ1�H�;6!�E� N������9�33:�pj�����ť5m.��
0^v�E�	1gJ��u����k�j��;@���V�	�Q��k��{���*�xl��HN"�&�w�7��N"�@�]H'\A�7���#����cg	�t�q�����o,�6�_�(���"i<4�&.#9��ԛLl�D4=�;�3��՟���y�J�t^D�/�"K��wr*R�(�1�ӷ��]��/��)���>�Gɣ�3���Q�����p�ɽ��xnh����zC�d�R�H�|��r=Ng=1>T��~eČ�8�o��&��>o*�B�ݼ�#G�,��% !���TNԗ���,<#��I� �����8=��,�5�j!�hQ�zo< ga�i��1��%�6�R��詶�i��&og]��D��R��w�b79t�a:=����q��
B��	C�/�Z��^TNv�;�]e*��� ��z���}6`�%�<7��/X-xy�$�) ���)hL�mll��55Uo�K��Ҿ$�歛��5�Sk ������84� JjbϢ�,��/�ԧ���w�o�J3��g�����G='����y�&Բ�!4 ���TQ����T���щ�}�����PRi�A�oq��\��j>e���;uՋE��l�� H���qH("��N�����참:���S�%�/i'��}^H||N�4�M�dcX<%}�y[[�Mnʨ*�=��Q�#x5m�B�����~������4\���CS�;�PJ�ՈQ�n���Pk*	/�&���*Pu��n�Ȇ��6!�xo��<):��fx�$Hh�T`�+��� X�nϯRS��unj
 D�i7��%��ǇW�s#R3vrT��u^�9��/�m���]��TI���&��F�D�U  D�:�J8dgRM�t����Y�԰���������\«z�4+26�2cN����SI=IS1��bM��#�
i_P�����d� ��_qC��E`��X��}��z�<��9=�ܕ��|j�\eN�� W�i��4zA<�c���"͈��+$EzZd�M"�0�G93iY5�<v)����R�Læ�}�8����ӥJ_W�J��5gN�>�/�i�7x&y�d�q��`�]O���m*G�I���b�As��+�H팂���GH�qJ�v�!������(<��:g�-(���K!ޗ�q2��\+Ԝ�4�a��ڜae�� Hw�j��B�m@�>�>��J��b�����n������'����Fm:O&���r=%�B�TcXL��]���)��T��U�Q��%��r��2����u/��q�{6�ެ;@B���W9�^TVJsz�8"'�}�����I�C��OUI;̂�wN���T�	OHT�Zw�DmAL:cow���S�U��0_!����E�vP�����c=TFkdr~U�έ�G�c�F�P���j:E��!�k@!�{�LQ���]���gZ�������	'�B�[���%ي��d+^I�'o����gX.ܼ�F�I1�!��WE��q�Nռ��8<���h�E��MƱ�X�J,$�N�T�Z��c�S&B�h�n���@�Y.=E���v.u��|9V���YkL#��v)�,1�@u`�#'Qȵ�ܓɺMs#2��4���}@1�V`���}�8�V�z��Δ�%eDv��1ڭ��# K�ގ������xQ�0�I��a�V�u��>#��7_#���2i�U�|^�R0�j���WU�����25Hn;.}��v����T�(�MC;�&�������}����{@�1�>�Z�f�I��ѯ��*�W���f�\94ŨTu��˳��d0,�7�h�~C4�;���d;�>��R����><�f�vdv���sHl�0�o)�B^�NVY�Z�(�k�_�)oC�����>q��`sK������X��"Cರ�k��Q��\*�W�,��8�U7���%#ٮR�h빂6�*T�MSR������� ��fU'�a��?2ԍ�~�u� F��Z�Fͥ���ۣ/�����A�Z,1N�=�ז0��N����ٰ;����p�s5��t�A�l-�=�dk@�н�i�A*L�2�n�~Pq��K����lS�k��Q�W*m~��4K~�R�?r�B��&�kǨ�}p�OM}�[G��w0�(��WFu�i�ƾ��Ѥ'��Zi���=��E�}��4�'M'1:�I�( ᆧSt�)��m�h:u)<3�e<��騘q�W]p�f�b\��R~Cz5�1�<�� r�c�U3�qD�KʟQ�^�Gu<��ǤP�?�e��,E
��ԉ�t<(n�AjJM��T�P����)�S/���*��g���S_�i)6M���c䈎�c_*X����)�7���)6^��zK��**OݙF$:>�?s��G1�+����B(D�c�N��d�I��8�<A֊��dx.��r�甔�̓\�m�t?0�AU�H=��.]N��>Ô�]d�BL�9[ �ȃ�JMpTk�ϩ�m�mkj�(��N���$����NK�(��u��.�*bjpiv�/����ڌ�����>��y[���H:�J]AW�A-�:�~��@��o$��T�8	W�C$���P�#�f!�'0�5�����"�t$z�tyq>֢*�n�4���h7KSU�@���T�D�0?
@���^�.{qf�|��C2;���{�	CՓ5�Q���C �#�#�
�	���NK%T�X��-���Y|�Lz?�0/�M��>�(z�3]����It#	��"şp>�Уwy���QS�x��I�:�K)E]�=�R��c���d��;:�^!A`����A��	��8�[��6��:6w��C�Hc���T=2���qF�pc�n!KN 3���Z������*b��rsK")�L�խF<�im�A�M�&�f����U�=r=#�>� �4�'�=�`9s�c�L0=����Ź��yӧ��@�R�E�
-�']�J�:AV��k�!�!�����<��9����MI��X�����? �4�#���j�}w�졨�e.$�2���N��aFjf��Q���IN%�r8�G�(�N��%{�p����H1ͬ�S�^����>\[}#�Z�!��Z
���½PU����L//�ۅ�vd"颹���+�S�D����&��6L��n:s�l�,N�X�!���E��"���ժnH$�v��v㐓��Ͽ%�FM�'SIG��>��ލ% ����d�h
Rڜ'G�z#�ǎϥ=����V8�yyA�"$E)t%�)~�z����7�Ƒ��i�x�{s�B�3ڛϤ��m�`5M���I2qf�.
	�$A��F9*���2��&��Ec�����O{ǹ�rp"@Y����Mg&��?}�4�:�x|Ig����rH�E���hH�aC�#"XN{��]���\r�.
_��7�*�֪]�G�L�� ��h����Iԃ�|L��|4ZV�q��8�ЁP�c���p]8u��	KXhtE�>�4����=�l*�uѬ`uy-�*�rd��!\3�Zj�������i�|��1/Nj��g�8CD�=Q�P�'�rbݴ��Ciފ��Ѩ�M`B��%��~UT�H&���?�~���34�I��3i���AmQG� /� ����=��i\�I)�˽������^:rD3���꣮ͩsVЙB=Rf&8��H/m�\��H�v��D~�$omy�],�[C �,ɫ{���"�qT�g�p||�4��a���ȋ��-	9 d1�@��J�� �3�?����ReI�K-ƖrQ�v{�ݻ�K����k+[���͖����i�ݲsm9�{$��?}.'�U�J�!(�fO�EQn�5�ݣɯЍ��:�Vp�hE����0	�=��9h�=T������� �3�TF ��8]إA GA�	�v	`�0J�V��q<j�����"y�WQ�\�.�z�=��У�>x�x"5��#��ҳ�6�mz��xh��=Se|��H'x0zB p��b�1uz��	���Z�ʠI6f��TN�&}~< ����ۏ��6�@�&&p�e�xzᲾu��> �*�O=��?j��]�WHc'U�v���}eԡ��L�ϰ[g��=�\m6E���h4�̪h\m`GÓ���R�:
B�N�Io�uQ�B�Pm��!ahM�25��=�x�!M��e�[W��+i������ԁ`A���,6�4N �w�kjj>:�� �a�����+� 4�P��յ���*�Q���ĴT2:���bY�.rQ �6�U��ZGQ�[�ʕ"�S���\1z�X�\���y$u�&P�d���Vӻ��=�b�4�N]d=�O<+Ȍ/]���z>��pc�x��f��m�#�+��o��)��rJ>��#y7Hl��2���h�ul�Tp{�'&͸�G�D޾};}��?�S�c��fϊ�E�Y8m�9�Ҩi�9\6���|G�0s�Ν<%g������G�2#�>;�� r�3q�ʺ.�z�sKl1��T��J�#�fx�m�~]	�/�L
8�.^�4r��hG�8�t"��_�d���Y|Eʳs��S�p�t<�9>x�c}Tc�=�䨣�P�^�\ ��_����ء+%��\��- ����_��l��Q�ƀK6��g��~>��G��ބ� ��P��-v%$r64xrQ��5�.���Z��h6��\�v��h���Sw��(��Fݦ�N�؂�B½V\��Ulb7/:�k/Ȍ�1��H���g������`iC23�V���կϰ ^oF��z�����p�e-��Y�gؗ�"�F��������s��,�n�mq ����+4a��sT%�����lîc����OV���>�E���Al8Ϙk<\W@s���Z�8�����f��IfIyA)�V��z0T�[�t���v�_����5_���!Y|F=74�B���*���p�ӄ�V����� !C���,>��;7ų�n�SyN8�e�����9y9@(8�4���|Զ7� ���D��[o�%)F�w^tN�j�î�+l��{����5dMm~��M��6���_})0�����O�Q�S����n| �K��pKT@�y�`��=�#�@s3rMi|\��M!��yGHF(e�;Q���L��5	�O@��
��0�����*�dQ@�sm����4�\�F$�{夡6ܙp>�R�9u5�}$����n�_q�<�Lwp�p��[�|�nw�P���J�<�M�!�
!����_̓�&QT�\��b��V��˗�uά�9����S��A*�� �<z9�fB�Q7l>�￿kq[lne��끷ű���\��i�nnaV짨I�MAxx1���������< �,6 o��8 ��iN�����ذ����9��@��I,8'���ӄ�,�`��L|�!�0��9+g��F$3Ȣ�{s�AW)y�%���a'pל�Ш���CM�s&� 5L����pN������:xF�)e�Lz)2H!�"\E�v������M��V�}�����l�5i��$�a9*�3�(?xV6������J3�õ<��ϼ�S�b�|'6�N0��q���>�Nw��w���m|n"���S�J�OvD��CR��	2����)���ka�ƮRl��hNӂ�0	���3 �BC6�����8\Y�$Z¨�)yeS�W&�A9�,��O1��O(^y����CѕK*[���m$��ƖlB*���=UF�j�B�2��a�p�Y�K��Ǌ4�Z�4MtE�Fk3��I��@�S�=�|=��\�������]��Fog5;��r���-1����;���T�V�|���4&'|��׊�����K��\c� 3�j�FGS^���%࣏>��������˗ӭ�7�� �$F@-���
Y�N�a��$_8�L�E8a��o����%���Q���g8��AC];��Dס��g�l����kb���n�e|��\�W*��������F�Օg(ї�h) �!�:��XF�i�/�a�W�H΄o��/�g�qd{UרENlہp���i���t�6����8}괌�][lN�@��S����O�ܧ�����<���٧Ϝ��l�)_\^Կ��k���u�%ZX2�~*��u2��28 Yp�S؆v�i�u�{�^z`�|��$kJ��]`���,����^l?������A	�_�w�*M��_&Uf�Y�HKӼ���Q/CS�����Wp���B� ~(�\��6�����v�*r�KRLZ���x@�\`N&�[0/��Ġ^������Цw�!�lC�<��`S�ښI�sO���q�,�-�In����l��^��io�-�rI�,���q��p�1�LBm��	CC�?��(�Q���Ι�C�J8+Q�b�(*k�R���x:H���tq���2Q:�A��#H�nv��т?~%�����=y�Q��|ԓ'��EqMM��ĺ��Ǥ��d�m��g�ׄ}��{:��m�Q��s�E�UR���L��]�/�	ʪΌ4��i�(<<(�S��ɷn�*&z�||��>�"�^�ԍH��{!���Ɔ8��>��)�GJm&0� Ţ�Kn�I+�c���e��A�ΐ8��^*�V��}���IH���h��(bG�H��&N~�SP�i��Rx�h&N%S7�}� �{	��yz�I��腖	��M��c���Ę�i�4�qTy����W����M���g��R}���pz�T���f�i���E'}���-[�b�!'�N���Ot�y���g[u��Բ��O�Q*��E
��{꼧���W��eXII0��o�������8��@}CI�!c�LTj�[���~�YL�?��ʩ�H��h��Nز6���2*��{�u�,\FU<Q��������cӽz8�Y����N�8!|M��	q�o��`U�
s�e7}����0$ �Dzp1�"�ܖ
a�Ο?��;?#��+A��J]�$&��ht\dj/�*t{�n$�,��-Er�����+ޒ�ͣ���l®���4��'�H�d�Nbc�Q�׾�N��@�sUH�d�K�*c㼯pd���'-õ��&�:�y�h����}w��*�m��������Iơ�(����p2L��P_�0j���@\�ԑ.!�駟�k׮�������X	C�$qp� $������7n(�ŽxHUjq&�A~8H�K�<0����}�$����H�����`�3�g��DGӜWW�<|���"?y�4�r�< ��T�6�~~��w��5PϷ���p��������ZGs8����7������$���>(^�G�C�J��-��հ'+�8J�|/cL�x�13�M��g�#���ykK�|��D���� Di���ϖ�x�7���&�R&��-��[�)ԀJM�Yr	��
h.)��V���$*�'�h�8m�NhE�g�xF�9�K�bC��d/��M���0i�(��Ln#\my�\ڧ�ȹՄӴ�#��{J��c�6����[�	��?�$�k�����	�-F�S�s}P�ۍq|�1�����k��7�rZ8x:�q��`:mۊA�P[���f��j1�7�dL�6�7�!��0T�3�Ϥ��%c�r��Y�!ۓ���s��y�vٔw.]�b�d4H|�d� *����9����7�o$�T�5��$Į<}�l�q�1ب$�M8q���d������I���\��W�H��$����_}-��
�Z;���`?�"�K�R�+��I�������D�S�CB�Y���W_}��L�9�EP��-\QT�Z�#[�=�X���sF��G7�M�io���M��p|]+�� �ǵ�Niׄ��/J�����3ʯD-87r&M���GJ"t(�G��7�^Hu����,<�|of�cPc�Q��nJ����&�Py���85�e3�Xd
~��_�yv��7|a��첻�[�t%q��=  '${0|�����F��'��!,h^�Mpv8gt�c#�z��[����'��d���ϊ8h/�����i�?�X*��o�}��ܠ�z�+�:y���$�H*����䑷G��:N���I�;�M��A�Q�>��]�!$���}|\]�N�7������K:�>�e�PK��|-@��bF:��&#|���3��Y3"�*v�UF�~`�pH8��l�`K�ௗ�މ�=T3��өre,^�w&`W�\��RWo9c�!,)��PY��}^�#[�S]yQ�#ܜ��$aH%7�^e�	9A����O{ܺs[z��YU������@A���=�e�sɕ�9/G��=�&Q�$}��>���؋�<���-�Z����r�9�˵X����͝���W�"U�O�6ւX<HR�,��J>��<�=�{��.ƾ 6��Q��?��2�B�-�/I���v4o޺^лR��P�*�x=nZ�Ň�4p`.�͛7�J*w��K�Y 6M���7��I��2�p���Q�Eu��SfՌ2^؋y���D�:�qVS����9�$A��3�k���L�cF(r��0����1�H--֜&�ʅ0R��Au�6ɕ�}����T0�������ϻ�+i�1�0��W�*�4C��K{&�e��
<�=B��c�=�^� D�C����>}�Lj��L�dʧ<{����&7b0���Q���h�ʌ�D��=|�H�#�O��{Y>pP�N*���� G��g'wռ;�.3�3�?�Uڞ��<��'�\9tPD0�·Mc8��8&����ܿ\��=a����س����8r�qv�/k�d���sX��U�6X���c�%&��2YT;�I0|/^T�N#�ۙ�H������s��9)Q��bE�*�t�T^��M����%O%mEFU�מ$$���#?��BЉ}��f��a��DANC6�"��!Ӏ���#u�!�-\6#WEmO��?q�-Ҫ����iDKH��)�Kl6�����(���W��2i�ِnEW�t����~�=n&y$)�M��6cU�AI��&��d<�-{���{�h��Ұ-�V��������!��qc!s��թmw����tR���s݌3��us}|0��@D���5�ϙ���k��D�,����#4+�Ÿ9����YR
��N,��k9}�y�pmlEn���#��r��!{��i4�{������	��F{0	��D���E�(��z j$�� v�	��~��N�,C٨EI�l�1�i�+c_��'��a�����.��X�qPo���g$5�`����T��p:����6#M��U˚�'u=N<P���;�R}I������u���A��盌�`s'H�G���&���y�̞Qt�z�4P'��kE�ή�Du���O>�D�AFU|�0����]\��,��Z�u�BF� ��-.�t�q��kZ����w@9OWoؕ>'AH��<[�f���"���C �P��h23�˝-ԼzZ�+��{���1�}9,@��r�K�s7�fP�;����A��Ov@�Ī	W6�R ���ے���=�u`.�<'=��vv>It$~��۷�Ҍd�	�N�����;�	/�F�z[1��A����Kj6�+-����IWQ{����pG9�
֎�Ho�H�����%K���[��U��-�A�f��س��^�!GG.I=sz�Nm�(��N3(̠h���.J�)�d�ƙMf�p��A�nn��N��&R��zSS�������M�Un�����%R�����U�͹����,<���==7���cE-��:���%5Iˤ�<��Y������2�����k������ٴjt�ζ�!v��՚>��|f'�Ae�h��DѠ]�X��̅d;���q�s�ޚ�]�M۶�NfyDk�I�'��c9X�����%zq2����H���c|d� ���u
���AT,*m]*XӼz6TJA�膌h׉W��9O��Ls�Y���7W�Sbt!I7�0l�w�'��}�⹂=R���!9.�'���8IO�7�fA�r�I� h��Ӿ�!�S�Tb��u�+�+�9�l��p��-Nx֑��S�J�ãv�|M��J�J)�h�X�q.��۽�\�0mǹ��s�[�h)���a��TI��]D�<uVL��*Αr�z�L���E�p�}m
=w� ���'e�H���Il��k{HM�����њ��q��`���~c��r�X�x8!It�����+Z ��b�9Y}�'+����!e�<PʝQ��X��*��=F�"��WH��?4�z��	�ؿF�9`�WK�JJ~j����uD%UN^,��a@��5�ɬ7HKƛ�f�Pq�R�頨�n0�B]?�l�%��n�u�'#̀b��q-��ی��N3��q���
�[�)l�5�ǌ+A)]��@Z����jFZ�� x��H�l���ٵp��z:����Y�B8_��E����Ɓ��l����gz�'R첳���"v��E|Y~�X�a�F#��Pp�&�O�zm]�{����H7�w�u1�ǜ�N_���q�`&#Y��C2(
)7�t nc�"s���k���U與8�|q�4��t:F]L� �L���;�v{˯I G���`�ݟ���\��<[Nڐ�����IA�V��|gFp1����h4~b�(��.�y{�zrrXA+T��jg(��H�H�:�d��=�sz(b$O;���Dj��xcS�#�� �R*7�"aWp)9�dQՏa��4����q.���h
�!��7�p� }V��쑰lI�R�x��$��) }"OhE����KA���=�I�0��M�G���8���B;�֋��f�2�]��Jo���/��o�ԋ�\Rb_�-i��FHDA%��N���S�\��t��a�r�����M�ίB�G٘k�|�4�������"Lm�H^^����Zz����5�*��X��u�.�S0):[{�|i^�L�G�niaob��k�6?��Tw8/
�K�ǳb?P����ic[�A��s[�j#�: �j�������H������.ʾá-*��x�Ç'rMِL��8�Uu��U`f�>x���y<3'���������;�4?�@�4`&R���͠����sH�A'x���i�R�B�t2�Y��C�)`����L{�v1�̳�I�4�v��*�y5q.8d��gL�7���ćy��+y��K��h�������Y�.^L����n_��>���ͫ&�)AE�h,>7��s�����͐��V��I\ޏ�˜��{�~��m�PrL( LSR����O� ���@mSD�����.3��N��c��h5�p�=sN��i����`e�]����[�YKE�}VS��ozo�
F*6Ա7}B,���Ey�ė��\����)$�]%V�xs��((�T	��֑�==�&6�Oj�t¼'$mqeQ@�ۦwŨ`�G�9�kN��/��f �X��ex�:��<�Y\|O|��=}&I�K��Q�]�}r�=sr�%�j�]q��Ncc�~��Ps�j��ŷ.:�M �1�d	��<�X�
e�xn����3R[RW�Z�{�&0G��C��t��Yi��3'I��if�p��f���0N���~��t@�"6�l��5����� sJ��s����d~�{�︱�2�S�^Q5N%�+N�(�l�޽򮮅Z:q��e�/ⴡ�H$��	@�������pb� 
h�3 bNx��'�\9�E -�ݲ6��ao8��z��N�s���`�-
EM}*��0@�۷n�4�|��J�q����~��󵪁�S :|�<D�l�}��]�0�nbG���G������3X��G��z��zˣ�I�y㺻�A|������n�=�z��{���O�M�ͷ_�+�^ѽ<y���ܩ�(-��%���8/[w��!	q�
dC�\27���ި�
������>Nb7◮�i���>����O~�S�����=��U�Gt6}��_���rp[�#�7gt<�Bb�?�G)��L����%�(N�5�i�x�â��B��u�E��&:)�4�&ɦ ֙� ��93c����>�  a,� �5��5!��8帹)��yr��ٵq>nݺ)!'euEBG.������[�\�e��^0�9fm��"R���ꪬb;J����q6F�ZH�S����8"O�!��J����B�O�{](7�w:=ى��C�ҽ����0��,0^��̙�EC�L�zEF8��E���wGa�Vp���G�H�G��L|��Lr��zk*ե@����;qx-A*����Δ�$�*6j-=�F"ٵJ�o�����=��C���)ӷ������溛���YI�͢^z�L��a����&w�.�f�u�f�O|���7�ҳ9�L�����'�n{&)�a ��h�}!�.)s����$)�m:�/)�^�9��p1�`N�&�Ta�Q�J��8B��5}��HjlS{]ѐ�L�h��������G|`��%�i[q��9�rsџ�ڕ=2U�]ٍfUx��l4�쫬�rZՒ�:�֞��b_`�y��x�����Q��	5�#I֗.�Kё76�@�o�9 lN7�#]n脲PM���J� ���.���p�����,"��o������?ӂ	Nc38ul�3�J��&�--4^Yb�-�a�@�����ƍ�z^�[�BR�s�"Ђ��¯mx�홝|l���@���'��x%�}�k'�7�F�BP�4z�S7�:6*�kBL��gQ4� .óHѩ���R/T9�D�ݖt���, ?O��r{�7*w�N[l�W�:R+������ը���ن�l�wD-��'�r/9������6��+a���qo�(���K��?ԏ{�ɟL�l�����辰aK������F�ðc�p[�?R����_UczCVY���kt%x���L�K--B��߸�>���鬸�2��(R3?�E#��c���˺6�1�ln��x�|�;<�y�Ҩ7Tʪ�+�*.M"����*�jѻ�*���s��U)��x���1h�����
Olg{���;;y'�e4��}T?��%'w&>��L�h����F$�\��OJ��K�>�U1��y}$	)Y��$����S|B�ѣ�1-����^U����G͜S�k�I1����yGۋ�/�@��%K�Z❸îEƕH��+��]}O�� �RT��{0�>�%�A�Aoee&������� ���g��箭y�C���f#��.TtNC�{�M���N-V���H�hxv<u�k�S��M�0�\4GTm!2l�D��m���.X,�_�&M�� �Q��u��6��u����E ��M��o�oJz�,�p6Ժ��%���ۗ�m�{�:k�*=�=v��/�-7�,�;w�9.�%���!�]��eù#ힹ���c>

g��wO(�N�D�gA]5͢M�����|'�r���-����h;�j8�TJ1!��p�|N|͙����2�\�&1�Hp3}���j2�:h' Fkl�=4Q7i�<_�Bՠ&�]=z�D�������m��PO����ay���$�u�㫯�V2��l���)�<�uX`��N��.�u��6������=�3�zMν�>|"}���ҵ��ub����*ZG͑�%{ґ�*�5�l��pb�;K��fy#�HF�M����8�}��M��3��y�JӒ�,ۻ2T��T��pЇ豦ւyuJ����Z��*�M ^���m�����0>�vqiA���9�O���C��C}.Xvhg��o ;f�w�����Vb��؁b�ٗ������ٰ5��~�$���u�p�p��#l��ZÜz��º!,>�\8!��:4M�����(ƃ�#p�IKωs)�M+k(�^��]�~CN݃���.�*�O�)�v��Q/]�f�͑#A��?tu��S��͡�Q,^N�Q8R��$��r����s�`����;õ���|�i�%<)�(:c�r�P.��h̉���\�oW����\v4�6A�-�>�r�lr�~gr�p{�`���,�O�\�4�_X���@��;����"2W���s.�O���3�泧�I�>t����Q$���m{�RH����J�Ϛ�����N�f6[��}Y�'д�`�_��xdK-msJ���'[�����A6�"�B"�xUcf�`��F�BO����Ltt��w��U���.�iő��7�B�J�������4�-eK9��!s� 7N)���
�0e��x>�\���ǜq�(.)RE���	'?�T�8�,�� -�n"ej2]]�g�;�-�;��`�0��35)X�3Sρ��x��l؜B��E%̓3C]ELwͦ�� w�U���� �If� 4�0Q�<h���ްWl@v��AP�7�� ����~����KaT�Z��7'���(�v��Y��q�b4��E�OY��ثgl�n�(N�g��'�[��A�6	 u�Be�k���a�.��R���*�*(�_�	ł��x�'�������zŖ�
�����}�88��XjJ��^�~�3�M��o���W4"8���b2���7��?�R�T�Q%�������L��5a|`Q2�.��p�*!@���q������I�;ܼn�k��M�S	�[�+rd��@��0�-_�A�ƒQ��,^�w��ݘY��x|����	!4���K�Еv}<,��8�^*��1|���A���|6�U�*�ٸ�{��m������S'��6o��UL��e�i>JH87C����,*A_'X��dj��~WYZ��)b�) �n�H��9�]k˂�{z=Ɩ�D��\�.���`wg]��S+�ή����e�1[k�Y3u�Zi~�I���g�@�0�:�4��{R�f�._9+��> �>�Z�i{nj-�U�
��+�7Ri;=�K��a�X#��"9a�~[�Z��ڽq\I3��x�l/�i��N��آ9:�o\s������uB�{1k��$���ܢ�#�K=a��'��yb�6�A�9,�apW1jl�����NH��cS��&���`Sh��X�cKi��R������뼺�������?��ȝ�=1��f��������93���}�5sR��J�J��}vG_�
�������gϜM�N[ƺJK����[R��ϊ:�nB���ك�w54rcmC�Ña@>g%یlC�9pa���
���ć���gC����(ꉈwu�ג@��B�:��tz���\B~$ے"w����,>��jp��z�o��Z����Pr>�,w�4��QO��Lh��w��5l#�7��8���	f��z�����G���~l�n��r��ܻ�@���˞	ʊ98&5uG%m0]�+�R���ͺ�<���߈Ld&B��{����eG��:���E7j�N_7������L��������|H���U����D���aqG�z��ё�؆���������\����?M_��$���w�}cj���X�#���~�D�.��u�f��m��8�����W���k�Ν[ⅼl��<%G��[n����3� ��onx����n�ϝ�%}�888#[��Z���`
p\v��i�J�k%����r
P0��vѻ��QaޤinaIFV����"��u��F쵽ae8��W�;�-"հ���#�-/_>W �ꀱ�������_�E���_�B����<�ٵ5���E=���׾5�q1�_����N?�u�:���j���`�q���XҨ��>�D5�e����Z��k��ܷ�����&���TQ�Kʮ9@lQ�O!R�Ӆ��N��uv��zUWz���<�"!	C�����1�N��I�����|I�G�������*N��v�;1��n�A� @h�hIw��d����yϽ��o�@���^{��z�:�:6�WD�3GeW���U�s���Ā�fr�b3"��b�^aӣ��$�MR���(���g�&�"j<3<�3g�v۔c����j�6�yR�+<�Υ��	��|��O��Y`��YW�w6���j*�$�;��I��vv��_����=�D^�yM bcv�7�hw-/i�P5�[�_�Jr��B:~�pV������ޅ��&1ʎ�6�K�HN�8 5��ڇ��lKww��6$H�T%pf:v�ί�p�uGjwy{�Z���T��8��$¾qsU2,�ѧj�Z;]�.,�0$|F�i6��� ��g�B�t�2�`��Y�,vs��N���qz�_~�g �q�e-��Ӵ��>��gA�97w�׳��y�������y1��ܓ��#8���C��Ս���M���/�������ͣ�j��
����^V���9�j�)/�ڇ�^L��F���r��O����V�\ͻ�Γ/�#v����'l�����&8�{��T.����/2��q|yv�UMZ��gtJh!f�V��Dh#�pF���8���9i#�Ct|������@P���I	���H��>I�!)��j>����_��<!f����=��8���z8����i�F� �be�J:��yU�Q?ۂ�������B���׾����L��~=}��SЈ�D ֳM�ti:�Q����QƩ( �ȁ���5�Y�i}�Mo����8�e5��d7��X��>R���˧_��O�����47����h�d��G���Sgi�������O��"kk�ɧ.���y��x��x!��=�#Yj�=�=�����N��ޗ�Ȣf�nfv>]�b8cN�h�N�A_I_�U���C�n���g�C�<�^�7��߼b�7?��lW�dU�o��Bz񥗅3���c"E�����~>TR�̙^z5;�<��1\l�4o���y�[x垍>rUe#Л��Z��P&6��EG�ƃ�aB��M�FXv�J��s1��撒5����$.�����4U�L11��ӿ˺wWF�, ����/��s�U:n����N���sMW8�7sI#�j A�%��q��^d6V�n��\�G��=��^^��,�粇DPz+{I���W��@�04����)�HT>�϶e#�Hfs��E	'pT������蠍�i�;iK^��+J#�.�4�������~�b��koO^	C�)aC�;�.���5'�1�O��[�P)��^oC� 3.bY���v&�]�TL�.l?�P��3O>����~�wrq��&!������H��vs�����9#T��xO������0Y"^�[��I ]C�pR#�/_KG����_��r)�����9sS��ЧN��w���G�B��eݺ�f�X��65ǫ-�)�,+T~�(�ې�2��3&e�����Q��4M`v�jP�^��{4��R�^`� �*��&j+�2�!O����s �D��f0Ⱦc��)���I|����[�;]^^4���'r���E�"���-�0���t4�Q9B���~�����.%���sS&��7�j�����O����*=��/������\�ҡEC��?pi]H���z:u�Io~5����yeg�ֽ5�S	��S�!�3�^V��)Z& �Q*~�H��?� Oi1��j@q^HJ�h�Ե,��`]L�Jm��7U�[�NU�S9\���o*�� w��i��t3���x�ߧ鹑�'F�7�C���a� m��ż�d �e��X�[�֕��]��"�
�w�y/=���g��m��mar-a�������'�Ns�3Ug�aM��Q��O#�Q��~;SE�]ؐ�(&��?��ڲMcF�q��G�t��~�ݬh�ٮ��>�(����8M�X�����Tvq��]��(u��ϟ�|](4|�~�����-#�4�z��k����.�3�y\�+xoY�N}��X'.fնF���|��(�4����8�	*���ګ����A��h�z�����X(�-��~��kJ����tV��}�s�^*����L��a�ޒ'�ĺ�
�e�x��T��@=���Ta�qkm�-b��7^��x�,*�5�f�呤M��ThSQQ���:I���X���M�s����度�q��.�_I���w���)��/|!=��s2�����t������i�}��i&K����WY�}�z����d��I#N8�7���\��!�r`�v ֙��~);����';	��{�=~�l)93b�	����]�� it��a&�^�n�Z'��S��mDd{�
�߆D
�&>�����8|��^<ʧ���ZH��}���=PT[��՗6�~���=LEm����Ϟ��AR��H�A�y��SD�z����hޟ=1�}�w��_����a)�T��B������Uf��=G����y��ϪB�d3�ŗ~�N��ռ��]z��3�<v�f`��#�s$>*�m��dUF��>w��f*k�\e���/�o���n��+�p�b�0�
���G?65u����!4@��1���qSJx9t�]G�����D>)Y��L�$5�����#��M���֙��4S�Uռ���ڣG�9:*�|��9�;�~���4(x�1�q���u�y�]vd�$5o���{l�/��2E�މ{�DI�5��_������U�vm*61��#����'*
��� ��Y�} 盳c�{Y�?!)���&��b"���pY[ۛ ��.�/������cGus��^U)�:�^�b�i��ܝ~%K]gbR�-�9O4���h�v>X�*�t�ұ{�W.�s+��o��N昨7Tj��/}%}��ǔ&���}/��ץ"���re�����jD��Le^��d���Dpԣ~��\��WO���� 1��⛢��ů�9}�U���ݪP�\� ��S"ٔ�{�[���7�-)%o��$SSm����ʨw��JZS[qR�UN
�}��4��,b�q�p{�>掜.*��Q�������`xj�Ȗ��f��q'!�d���b�X�dSi�/�߭Z�I��:��x7��ގ�0��~,���_~Y��g.2�.4����n�����CF ����R�b�qG�<�j���>�	q��m�8�+�ӵ�g�r�
��|�.y�F�14�n<VZ7f�$��w�&�T^95z�Pl��b[�����$4CU��z~��r`@e\��u39�/�4>��u�0k�8xSw�$A!�\���I'�\��*leWui��E!������K�G�c�*����n�-�΢2��i�fO��l��)�./l(ǅ�ԔAh9�9�ٹ�#�v�َ�)_�j�;Wx�|_���Y4"kl�~��l���FNO�`������i���k��3x:� Q5�،��-k�%Ŭ�����ݫڸ='D�Q�����W��=�|�sOʆ\�|U����P�o��N��#�K�K�Ig3ϼ������)�| ʅ�=���UU�rJJ"ٽ�~��AJ{��i�:ɿ�����;ޥ�W%���,d���OF���t�׷$�ׯh��k ԰��^5M4FKE��mF=() �n;	�zn�v�a�9О�J�߶aZ�
l�J�1O�o�9M�-H'�Ŝ��y�>�`z�D���N���p���ƠF�O�,My�IWЯRBnH��׽o-h�K��j��f
�Y�o
�j��RE����Moբ�tͥ|�.X�:�.��H�`�w����裏+��^���
g3q�� ��Z���~Q�}��׾�I �!˻fʾ�P9�,�Z}��d���B^��^5r��t]� T�Zȼ���;�v�,��|(�������kO��占��`���Ni(�KW���J�S�d��69��@��l��|���pY$pZ��Ͽ�m�?�3o��BvC6ϲ9�sם�"5��0��ݔ�1�0P#F���<���a�T׳*k; J<?����!��4f
�<C��v�H�g�䝷n'�2�B���A�/�Ҷ�|]YǑ������ZבGj�l~��GU�?����H/H���Y���彲Pl��mt�����/9G�O�gdcs����B��1?���2H�fm�aVm���� Z-������=;=�S�����/�g��S	�M���Oq�(���f�ī�&���4
=Ć�?C��0���X3����+�k<��y'��B�ǔ��Y����:��)`��d N'����T����Ϳ�=^z�e�| Ck�j��:�=ɽAٓ;�MY^X�����g9ZV�s��PCaTϠ�O=������H� �Vl�Z��f���q�Q&g�eCٌ�����i�қ�G�Yx'� ^&�Fj4xo�֨T��=vyI 1q���r�*�ɕ�=L�9 ?G���B�ڸ;�09)�I�&@e��$�2w�qb,*v�jH}p]x߱+����|⊶AhhJ���	<*6���7��y8g��,��,t
�vr2;ׯd�.c*=�������埾�^y�%B1�$;������.\�y~�l�3����<&p7v� ����D2��!����YqH�YP�k����(���rhӇM
Q�|ĈɄ�]�y�\��@��>D�⯽qC:<�.�ay�I]�{qʈ�I^�5��Og���̌b�(-hH�^���v�;48��=��x�sUS�:�F���5�SD��.?��C�mP�T� L�/��^�ɋ�^)�'���2�P�L�q���o�� ,y�9em��EU�u��HB`b�P�˱Aw/+U�E����Դ��#�l+�����'c���[��	Ժ�f��H��!��3�9h��^!]o���L�Y��Ii���x�8w���g�{��� T-������6niW������;꺑oh�n��	i��o}K(j�4j�h4��&�n�!�-`�N�|@�TЙd3x {S�k�s4:ن��7�V�OV�8c��;>!q@H��+�ӱ�1�;��.ZvI�`��=��}+m�E^��ZZ�N�0؄Xd^,��䯺=������`�/Xֹ%�L���e �)���1��Z���$�>6�nB��axE���hW�^J�m�@ǽ�����\p�=u�1�Aj� @���/n�r~6�V
��%C)"�8=��h�+)3��r�-�a�|�g-W��f��p}V*�159m�]N�w��D��XHp�4�QqY�j�4/E�"�G��͢'��Ǣ�^������5Eg���9�G�BO6Ӈ�SC ���B$58�W�ʍfK�U��F�K���x��z8obKe`ZӠP�𞬹f��N��=��x^~f7�sg�B#pF�yB���+����%�Y�|�9F����Dvw��8d�2"_"Y�HS�)7�6l�4B�͋A�#h��G��E���X*��KblqyH�kH�2[6o:�<
E��9eؒ�I9�&��7��nN�~Z�&>�J�����VxW�5�H����8ZvEńK|A�"*È������� �VF8������r�����MK���0�6ڷQ�Ua*�n��ڏ�6��ٙY��XW>��]G�:/�=����J��&x6�����5���=r�Ps�($	�ـ�ѓZ�MԼ��u�8R
��vD�m�`� �������Ԇ�a����c�2��'��3�{mH��`"l�����9;����]�Pޟm�ة�u���M��8x�\�`XP�AO6����~��RgY9!�RD�N�g�*�Wm����j�ɟ)p�$�H�е\A�st�H��'��G?91���7+ra���-��M� J���:�5���&�8+v� </:Ɣ�A����3K�%ӳ&\�J�lZ���q�)~���jT%�j��i:$yI����YJp��ά�DhM�������3s�)�6�c�`q�����Os�@��E�&�G�jZ����<��fvcNhH�ɓ�˰��*�<'�FT�f]�m���$���M�hbC����V�B`|):q�5�"���̾ʞ�z�,�.���bhQY��2�]̟a4��"�߳����V�΋$f�w@^��2���Y��p��~v��H�_`f
em*�����@C�m�[���h��,�V��� �L΁��0�&$�N�K�b`�B��c�t���i2�"�)�(𫨟�H�a#�.y6�
���A�r��T3/�u��U���CRK��ˆqM#X+}N�ا��@:���Re|�~ޑ��G���|����暢n��Ն��R�\s�h���+��(�7?�8�?D�Gr,F?��O����ny�'/�OG��"���	H�䭿�
�m�[��RO��s�}\�=��]^8ҹ6Eƺl��,yF�.F2QO�W�uwRܤ�A��Rxnj�(G2� "yIlX�b =��m����6]���ިf�X��^E"��r�tgR@�M]G�F�fÏ���6،g���I�jW�=T�R6X ��l�/���ᗻ������z��8��k��U��d�����߉�Qa�`��uv���q[���U�r���/О��2�����3�= ?}�דtF��ɓ3>�}���<ڔm��1ݟl )N"��1�� c~���v%8m�!�PBa{�7l��h��#�r�k� 5V�j��n�����]�H��؄�9�$�#O�������u��!� �G��f��t$�S�����G�x��wk-��fH�+��{�%<��M��2���Άp��C���B�zF�P)�!�����o�a�_��O�%�Ϟ���HF��sx����C��w�dh6J�{�r{+��2fd7>9����Ʋ�+ҙ���H�eQ09cҊ����h�����x2_�$�tPU�S�\^<K��hs#=c|v�`z�}�jq�M���^�~F�A�8p/rʐx�������������kZ��Y�zW���R#���C��0��R��k�G��kC�l�ۣ��Ȯ=�F��]T9#�5P��ZbQ�,\�ʎ�:��r�����Rk���q�gZ���-��^5��^����q�:�%�+G����}A-�߀&$��n�[�1����{�/�������H]�N���i{e;�fg{ۇ�,9�_�����$aC�sJ��w��7R:�MZ ;�0��?�6;~�� �^���N�e��֋qRa�wސ���L�p4�#m�׉i;{�����lז5R1�PsG��|�i�jzvZ�\i�6E�eۻTA��mv���2�� �Ɵ4��F�Pc8!���*J&�ŽAHb�����j�80v,���|JN�_�g���-E�s��?�0b4�k�>&�SD2�� �����a��H8mB�4uBj��٨��	����:gb�Դ���v�Mmm���T�L��\Aw�)X��Ń�M+, �o`�\7T_ ���t�
XP�A؛��XR渭!/NXF C����`pJ��k$�</�b���mm2]�l����~���u	{p]���qb�F4#{0ǰ�)Ù�y���N�6�������0fsɓ�l�@/V���U�g�"J4NOI��߶��ㆴᚢf�|���]��!�N���]�|���m��m�!=\�"��]V��m�NnF'�2<�)|W���QU,<)���^��(����]��J�	@��iTjSj���*>9;�T%��C#�4/p���H���g��@ᡞɼ1�*�S�4,������SY�ƖCj���F`{����%�� �3�z8�[cG+L�Mb�/h<�$QAc�[�sy�I�@߭&.cw�7t⢮��1X$5d:�P�/OS��R�X}#b���r��k��6��p?5d��M���m��"?�F6h�77�U5�S�)A�o ��B������M>�p��s]�2�Ե���,d 1X��򉊋�ρ��mJ�)��V���I����э����u�^��7�?t�yf�P��Y(����=�.��,���g�����Ą�
+v-G�R�������2Ww0��}��mh��*zYļ�&�:�w�����Ĝv�4��(��76o{�J�܏MA��ݽm��zR�M	M*�]bRji��a��#�O��tBJ����p���w81YD"nz;4��$��;�_0�5��}%��;Ө얌�
NM�;jE�n�Ԉ��q��iP��h�f~�E��h���X����q�7��q�Q"j6�R2�{��֟���>�J*��(�-���7���fώ�D�2L�/F[�~ii!V��3ڀ8Q�����; =�i����Мu4"g��`�����-�~�
^ר��(\�CΗk���"U���������ѭ;�j����CQ�hZ�ں��(V���=�Th6��Q�F���3�9{����5v����E"�]�q�+�o��|%�g�i�z6�@G�|���$w�m&��?yD���Ysx�
���j=r��qvAً�A�n�M�Pgv���6���d��r*f�#u�(0�$٘ �]��5/����C�瓺z��`�G��īa}v7z7*#��mx����Wll7d��t^��f��� ���5��>{2�l� $5��Q��IMQc�T%.,%6��m�0VVAd�9�J��L���y�}�A�Z�ъ�4:ޡ��60IX��<<��0�D6I;Udf"륂�p�	x��wD��i�Y�PC��l��4(m�ٛB��(8�H�؛� �2����I��֝;%�6������ AW���7מ��d8�sb�i8�W� rL�vNK�;����"p�5����坔���G?�sh ���մriE�+6�g��Ϥ�Fz/M:%@�W���F���}A�#�{ާ^:H��S_ �G�p�����Q}X6Ed�RCVGfXD6���,іt{]�skÈk���4�&�f�$6A6e��}�9�p�2�g����F��m7��eH^�)����*[�n�I	h$:V5�s]�ɚa7x�M߁�
���)���6�Z��mf3=��#:�*ߪU���R6cR'��Qw^�9���c���T�4&>��Ӣ�
|��<��s��T��[�[��>��+�!�H��w��Б�������C���o����&��Jc���
9襉�ImK2��/�inn�G�N�ԅl5:�	�\���Q*�?����*Y8�lR|�g��4�ܚ7y~�IYfc�\�w|��Al��?��z��U��u�$�ϘX��ߍ����n�"��U�$��c�[ؓhn��mڼ�Kl��0D�����mw5��b�^�ͫ�D��ZP
��.m+�ܑ�P��n��k�+����$�*f��1r5��w=5�Q;B��>�j=սMM�"�ü~�w�pqEj�����G�e��b����6��ʠ���U��Ơ�j�����j��8	�&�T� �������0u�'=��ea���ţ̽ex0s; >J�I�|���Ȣ#}e2����-��t�X�FUb.�/�ܪ��Os�g�G����R�+(���Y�mM�1N�N'�� �N��G'�'J����L��j=�ZU��}�i�P��.74&�8�=��� m�?�� ��D�x� ��7��h����NvÆ�t"-���܋Z�f�*�!��Ѡ7*��RY��{5�JuD�Px� �o�QGWKj��Г�����R�]-*�\�Fs���5Yh�J(�Yi�(�Յ'��>f���!�S�jgcC����g�t�����<\m������u��N���i�Ջj-mûrJP�a\Q���YX�z���z�4jf��:6�1$��5��LN��}��N-��}y��h8:U�J�|�v7�7��v����5(�V%$�~Y��`U�6#�F��چ���i+A�CxN��/��|}y�����,ÊGjO��=yH[��)���s�.b׶���P��In��R�D@f��4*�b�yVbK]���{c�U%��F� �)Oɪ���^��F.�p4V��5������O����_4�0�$c���S��(�e9p���w���[r�q����AE�2L�BW)�8�3n��i9�p�{��嘬����J�t�sD�8"hk�Ɉ���o4���)�jH�X|FN3m؁����ưu+ �b̷�@���/Y��У��W�9%;�='������g���`�H�3P����:�h�z�����j�:X���.���~�F�����*1��Aa��7��
D����da�'��n�2Ζ���>'(R�:�>�.�_}����e���u�O	��������";v�}_3��X���"(i*x��U�+�\�6U����nLG��6��V���,��s���k�/OPJJ�k�y��	��w}6	P	M*ܞYu4l˄��M�{=�_�0Q95^���d�Gs8�^W1�{"Q��ؠW���pb���m;����K^�lVO�mT��S� 8d�m�­�����M�te�v|@�I��'��4��V(���(#�B����"~l�-R�]ؾ}�дwl�d��@.��~7�r��R�%��}a�����Q� �5q6ʱ ׽��>�� �;a��m�>��Z}{�H��	��Uގ��M���u�D��~,��\�E��z�>Xxd�t�Z�G��[�M7£���Hd/���B�4To�P��x7٬�3�z�+$n-iTѸ��pz�9�=TQ����p�tp3�36��Y�n�V��ꧥ�O�Ƒ��@���@��nM��#�"2_��py9PI^�1�a�6
�=����T���o���WPYt�d�ʚ�-}��ʍfur��#�: ���޶׾w��D߽f�2�q�r�cݚ���Z�g����*4w�!w:6w��W 8>���`>9{Y�F=���M��Ƣ��rM=��d�����-b奆#�u8Ђu����+}�B����9p+j�dc�9
�/�Qc٩��:���)�)��� Y�@�8h�Z����"�t*�@��	)*�OQe��i���b��c�7ڕAj�m�q���	�����J���ӕ7��j�o�*�� �f�-qh6ʒo}?��Xr�}Fa]E��N��T��H�X[uO�S�96����*���F��1V��-�B�Z�99ʊ\�fmdT1.8ݮ��r��Sk�#T��oH�����=�(�l'�6ia��wD�mSЌ�!�;FZ����|�,���Y-�F�v��hY#�y6�R��1�6�6$��֤!w6��J�GG��M����&���k檛�6�P)|�`د��P��p$�MsqU�7F̎�u{QZ�T�2��6��~��ؔ8)�&�J�YM�����y��ݪy��UF!g�{PZ;ND�"����
���L�傶��"����@i��yK܅�Hfy49��H���ć�	充��Q �؋�m�����j�T&�~�}��0�SR�)�i��I��G��*�}TD��F2��UU7��{���<�._�,����;h�|�i��&1�J
�{�֌����B�/fy����փ��	�(�Bhz���G���Zt��&��s]@%��C�,��>x:u�T~���P6����>>c�h؎�ߔ�mz����P�����oR���N��'� �5kj�xR���L����=N�	{
�J�T.x=5Q�.�l�a}3R���RޮWO���/�\�ɴ^�V -�~������ee�LIZ)�~��'���q�hd�c�A�	غͨ�Z��>w���~U�K����D����u����mSw]��� ,3ސAe���"�M�k���7&<�ؤHQ���'|R�~�sMj�3ڳ����[�'���2D�$�1��������>���'5[�6�OT��}��X�˚{<��'�==w�cC�߷���pWKF��_�Ro,T}C����lc��=�kۛRu�-����]O�F������~i�}C>�;�!��]~Ԗ��΢��z��5�SW��������7�����t���3��<i�aޯ�M���cI"������̦|䆘�{]�oH��d|���-w9�e��rI�r_4�=x�o�%�鄌b����Z�S��G�3@2�>S�_ڲE��^F�ُ=%��R��z<r�k�X�(�X%�Dc/Ζ��ޯg��'��U������O�mu�;�J�¹���I���*^�c�FUb�Q�޽�>�iS>vC"Zϫ�?�DDa�٨Ƌ4��|;���f�Ft�5�kσ�Q�s�2������L�~�������z�#��q��;0ݿ���|��	i�b�۔E�?�}�anĝ���y�RQ�Oe���[������������8e�����>�l�M5��;]��<������	]1X�Bi�    IEND�B`�PK 
     mdZ �b=�' �'                  cirkitFile.jsonPK 
     mdZ                        ( jsons/PK 
     mdZAT?{  ?{               ,( jsons/user_defined.jsonPK 
     mdZ                        �� images/PK 
     mdZ�&�y`  y`  /             ţ images/8c2f1315-cf23-4ba8-a920-becb97f13280.pngPK 
     mdZ�����  �  /             � images/6fc4b800-efc3-4a5d-827d-9566cfd108b3.pngPK 
     mdZ�?���� �� /             � images/ae82c023-d9d4-4942-aa8d-ab2ae3c53d73.pngPK 
     mdZ�S��*  �*  /             �� images/cbf7ad0e-0f08-44f8-98a9-dcbe92af212f.pngPK 
     mdZF�i~�  �  /             �� images/85e66502-362d-4a26-afcd-97fbc4859675.pngPK 
     mdZ�  ��  /             � images/b13518ba-21c5-4f60-a735-1d8041d11d7b.pngPK 
     mdZ�+s`(  `(  /             � images/8a1d81a5-79d4-450c-9f72-108cd2673013.pngPK 
     mdZ��/��  �  /             l4 images/aacc0029-e57d-4614-a443-d9bee65b5175.pngPK 
     mdZ�1��� �� /             9@ images/1d90a712-93d7-4555-ae10-1782f839eba3.pngPK 
     mdZ��S�  S�  /             � images/e5551f5a-2fb7-4493-9527-57db21faeaae.pngPK 
     mdZ���I �I /             �� images/ae036c7f-e258-4627-a75d-99715ec815e7.pngPK 
     mdZ��<�`T  `T  /             �/ images/69c28b0d-a0ad-46f0-a190-03e6ecfe42fd.pngPK 
     mdZ?�>�oH  oH  /             U� images/a038ca8d-f9eb-4e93-ad0b-b831193aa106.pngPK 
     mdZ-s;�.@  .@  /             � images/3e0a96b2-ef1c-4fb2-8b57-d71cbe1f3744.pngPK 
     mdZ�.��� � /             � images/ac27922a-fd15-40ea-8551-3be3f9cd5316.pngPK 
     mdZֆ����  ��  /             �-, images/49e5ee10-9185-4279-8a25-10889e7bb4ef.pngPK 
     mdZ3��C� � /             ��, images/cff7cff8-0125-49f3-ae91-9e6ccc0a4cc7.pngPK 
     mdZ��� �� /             !w8 images/7b19d218-2217-455d-9a43-b73a208c2c5c.pngPK      u  "%:   