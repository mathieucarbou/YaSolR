PK
     #{dZ�5,*Q Q    cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0":["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_3"],"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1":["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_4"],"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2":["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"],"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3":["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_0":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_1":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2":["pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_5"],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_3":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_4":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5":["pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_6"],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_6":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_7":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_8":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_9":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_10":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_11":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_12":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_13":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_14":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_15":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_16":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_17":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_18":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_20":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_21":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_22":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_23":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_25":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_30":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_31":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_33":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_34":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_35":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_36":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_37":[],"pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_0":[],"pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1":["pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_2"],"pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2":["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3"],"pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_0":[],"pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1":["pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_2"],"pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2":["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3"],"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0":["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"],"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1":["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"],"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0":["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0"],"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1":["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1"],"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2":["pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_0"],"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3":["pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_1"],"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0":["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0"],"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1":["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1"],"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2":["pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_0"],"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3":["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_1"],"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0":["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0"],"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1":["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1"],"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"],"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"],"pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_0":["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2"],"pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_1":["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3"],"pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_2":["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1"],"pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_3":["pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_0"],"pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_4":["pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_2"],"pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_5":[],"pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_6":[],"pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_7":[],"pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_8":[],"pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_0":["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2"],"pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_1":["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3"],"pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_2":["pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1"],"pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_3":["pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_0"],"pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_4":["pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_1"],"pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_5":[],"pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_6":[],"pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_7":[],"pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_8":[],"pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_0":["pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_3","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_3"],"pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_1":["pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_4"],"pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_2":["pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_4"],"pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_3":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"],"pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_4":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"],"pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_5":["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2"],"pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_6":["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5"]},"pin_to_color":{"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0":"#005F39","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1":"#9E008E","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2":"#FF6E41","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3":"#00FFC6","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_0":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_1":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2":"#E56FFE","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_3":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_4":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5":"#BDD393","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_6":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_7":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_8":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_9":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_10":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_11":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_12":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_13":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_14":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_15":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_16":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_17":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_18":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19":"#005F39","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_20":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_21":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_22":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_23":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24":"#9E008E","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_25":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_30":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_31":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_33":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_34":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_35":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_36":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_37":"#000000","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_0":"#000000","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1":"#BDC6FF","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2":"#E85EBE","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_0":"#000000","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1":"#BB8800","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2":"#010067","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0":"#0076FF","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1":"#85A900","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0":"#0076FF","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1":"#85A900","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2":"#A75740","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3":"#E85EBE","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0":"#0076FF","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1":"#85A900","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2":"#01FFFE","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3":"#010067","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0":"#0076FF","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1":"#85A900","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2":"#00FFC6","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3":"#FF6E41","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_0":"#01FFFE","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_1":"#010067","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_2":"#BB8800","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_3":"#FFDB66","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_4":"#7E2DD2","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_5":"#000000","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_6":"#000000","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_7":"#000000","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_8":"#000000","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_0":"#A75740","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_1":"#E85EBE","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_2":"#BDC6FF","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_3":"#FFDB66","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_4":"#90FB92","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_5":"#000000","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_6":"#000000","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_7":"#000000","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_8":"#000000","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_0":"#FFDB66","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_1":"#90FB92","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_2":"#7E2DD2","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_3":"#005F39","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_4":"#9E008E","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_5":"#E56FFE","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_6":"#BDD393"},"pin_to_state":{"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0":"neutral","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1":"neutral","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2":"neutral","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_0":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_1":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_3":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_4":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_6":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_7":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_8":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_9":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_10":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_11":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_12":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_13":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_14":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_15":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_16":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_17":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_18":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_20":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_21":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_22":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_23":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_25":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_30":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_31":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_33":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_34":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_35":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_36":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_37":"neutral","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_0":"neutral","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1":"neutral","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2":"neutral","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_0":"neutral","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1":"neutral","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2":"neutral","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0":"neutral","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1":"neutral","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0":"neutral","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1":"neutral","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2":"neutral","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3":"neutral","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0":"neutral","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1":"neutral","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2":"neutral","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3":"neutral","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0":"neutral","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1":"neutral","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2":"neutral","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3":"neutral","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_0":"neutral","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_1":"neutral","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_2":"neutral","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_3":"neutral","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_4":"neutral","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_5":"neutral","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_6":"neutral","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_7":"neutral","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_8":"neutral","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_0":"neutral","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_1":"neutral","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_2":"neutral","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_3":"neutral","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_4":"neutral","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_5":"neutral","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_6":"neutral","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_7":"neutral","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_8":"neutral","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_0":"neutral","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_1":"neutral","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_2":"neutral","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_3":"neutral","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_4":"neutral","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_5":"neutral","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_6":"neutral"},"next_color_idx":38,"wires_placed_in_order":[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_29"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_28"],["pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_28","pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_1"],["pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_0","pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_15"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_29"],["pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_3"],["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_13"],["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_14"],["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_15"],["pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_36"],["pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5"],["pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_0"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_1"],["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_2","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_1"],["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_0","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_0"],["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_1","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_2"],["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_2","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_1"],["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_1","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_2"],["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_0","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_0"],["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_2","pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_1"],["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_1","pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_2"],["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_0","pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_0"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_4"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_4"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_4"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_5"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_5"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_5"],["pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_12"],["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_8"],["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_9"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_0"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_1"],["pin-type-component_a8221eb9-381c-43f6-a63c-1fa17c525231_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"],["pin-type-component_a8221eb9-381c-43f6-a63c-1fa17c525231_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"],["pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_23"],["pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_25"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_0"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_1"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_11"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_10"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_0"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_0"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_1"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_1"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1"],["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"],["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_0"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_3"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_3"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_0"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26"],["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_2"],["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27"],["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_1"],["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"],["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6"],["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_10","pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_0"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_9","pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_1"],["pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_0","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2"],["pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_1","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1"],["pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_0","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2"],["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"],["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"],["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"],["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2"],["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_0"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_1"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"],["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6"],["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4"],["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_5","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3"],["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_5"],["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4"],["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4"],["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2"],["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2"],["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_6","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1"],["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_6","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_7","pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_1"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_8","pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_0"],["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28"],["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29"],["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32"],["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_2"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_1"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_1"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_0"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_0"],["pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_0","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_5"],["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_7","pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_1"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_5","pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_0"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_7","pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_1"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"],["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"],["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"],["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"],["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"],["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"],["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"],["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"],["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_0"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_1"],["pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_31"],["pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_30"],["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_4"],["pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_6"],["pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_7","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4"],["pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_9","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4"],["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_5"],["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_8"],["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4"],["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2"],["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2","pin-type-component_ae34f7fd-5bf6-41c5-be78-9d886ea0cf65_0"],["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3","pin-type-component_ae34f7fd-5bf6-41c5-be78-9d886ea0cf65_1"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_ae34f7fd-5bf6-41c5-be78-9d886ea0cf65_2"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_ae34f7fd-5bf6-41c5-be78-9d886ea0cf65_3"],["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32","pin-type-component_ae34f7fd-5bf6-41c5-be78-9d886ea0cf65_4"],["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28","pin-type-component_d357a112-8ce7-4ca7-922d-bae950c817be_1"],["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29","pin-type-component_e754101b-2bd4-45f8-8367-dd2d1465a844_1"],["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1","pin-type-component_d357a112-8ce7-4ca7-922d-bae950c817be_3"],["pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1","pin-type-component_e754101b-2bd4-45f8-8367-dd2d1465a844_2"],["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2","pin-type-component_e754101b-2bd4-45f8-8367-dd2d1465a844_2"],["pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1","pin-type-component_e754101b-2bd4-45f8-8367-dd2d1465a844_3"],["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2","pin-type-component_d357a112-8ce7-4ca7-922d-bae950c817be_2"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_e754101b-2bd4-45f8-8367-dd2d1465a844_0"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_d357a112-8ce7-4ca7-922d-bae950c817be_0"],["pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_2"],["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_2"],["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_1"],["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_1"],["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_0"],["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_0"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_3"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_3"],["pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_2","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1"],["pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_2","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1"],["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2","pin-type-component_ef73fc61-5332-4389-863a-156932dd9fb0_3"],["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3","pin-type-component_ef73fc61-5332-4389-863a-156932dd9fb0_2"],["pin-type-component_ef73fc61-5332-4389-863a-156932dd9fb0_0","pin-type-component_8774d229-a262-497a-8b8f-89515ac3c08c_2"],["pin-type-component_8774d229-a262-497a-8b8f-89515ac3c08c_3","pin-type-component_ef73fc61-5332-4389-863a-156932dd9fb0_1"],["pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_4","pin-type-component_8774d229-a262-497a-8b8f-89515ac3c08c_4"],["pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_3","pin-type-component_8774d229-a262-497a-8b8f-89515ac3c08c_5"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_8774d229-a262-497a-8b8f-89515ac3c08c_1"],["pin-type-component_8774d229-a262-497a-8b8f-89515ac3c08c_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29"],["pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_3","pin-type-component_15115ffa-76d4-4ac1-807f-112999c7cc8f_5"],["pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_4","pin-type-component_15115ffa-76d4-4ac1-807f-112999c7cc8f_4"],["pin-type-component_15115ffa-76d4-4ac1-807f-112999c7cc8f_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_15115ffa-76d4-4ac1-807f-112999c7cc8f_1"],["pin-type-component_ef73fc61-5332-4389-863a-156932dd9fb0_1","pin-type-component_15115ffa-76d4-4ac1-807f-112999c7cc8f_3"],["pin-type-component_ef73fc61-5332-4389-863a-156932dd9fb0_0","pin-type-component_15115ffa-76d4-4ac1-807f-112999c7cc8f_2"],["pin-type-component_15115ffa-76d4-4ac1-807f-112999c7cc8f_2","pin-type-component_8774d229-a262-497a-8b8f-89515ac3c08c_2"],["pin-type-component_15115ffa-76d4-4ac1-807f-112999c7cc8f_3","pin-type-component_8774d229-a262-497a-8b8f-89515ac3c08c_3"],["pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_0","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_3"],["pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_0","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_3"],["pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_1","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_4"],["pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_2","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_4"],["pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_6","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5"],["pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_5","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_3"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_4"]],"wires_removed_and_placed_in_order":[[[],[]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_29"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_28"]]],[[],[["pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_28","pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_1"]]],[[],[["pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_0","pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_15"]]],[[["pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_29","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_29"]]],[[],[]],[[["pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_15","pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_0"]],[]],[[["pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_28","pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_1"],["pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_28","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[["pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]]],[[["pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_29","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_3"]]],[[],[["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_13"]]],[[],[["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_14"]]],[[],[["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_15"]]],[[],[["pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_36"]]],[[],[["pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5"]]],[[],[["pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_0"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_1"]]],[[],[["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_2","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_1"]]],[[],[["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_0","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_0"]]],[[],[["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_1","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_2"]]],[[],[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_2","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_1"]]],[[],[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_1","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_2"]]],[[],[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_0","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_0"]]],[[],[["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_2","pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_1"]]],[[],[["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_1","pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_2"]]],[[],[["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_0","pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_0"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_4"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_4"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_4"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_5"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_5"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_5"]]],[[],[["pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_12"]]],[[],[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_8"]]],[[],[["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_9"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_0"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_1"]]],[[],[["pin-type-component_a8221eb9-381c-43f6-a63c-1fa17c525231_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]]],[[],[["pin-type-component_a8221eb9-381c-43f6-a63c-1fa17c525231_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]]],[[["pin-type-component_a8221eb9-381c-43f6-a63c-1fa17c525231_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]],[]],[[["pin-type-component_a8221eb9-381c-43f6-a63c-1fa17c525231_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]],[]],[[],[["pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_23"]]],[[],[["pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_25"]]],[[["pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_36"]],[]],[[["pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[["pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2"]],[]],[[["pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5"]],[]],[[["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_13"]],[]],[[["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_14"]],[]],[[["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_15"]],[]],[[["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_0","pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_0"]],[]],[[["pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_1","pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_2"]],[]],[[["pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_2","pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_1"]],[]],[[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_0","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_0"]],[]],[[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_2","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_1"]],[]],[[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_1","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_2"]],[]],[[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_8"]],[]],[[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_4","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_5","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_9"]],[]],[[["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_4","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_5","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_0","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_0"]],[]],[[["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_1","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_2"]],[]],[[["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_2","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_1"]],[]],[[["pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_12"]],[]],[[["pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_4","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[["pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_5","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[["pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_23"]],[]],[[["pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_25"]],[]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_0"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_1"]]],[[],[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_11"]]],[[],[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_10"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_0"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_0"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_1"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_1"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1"]]],[[],[["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]]],[[],[["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_0"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_3"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_3"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_0"]]],[[],[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26"]]],[[],[["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_2"]]],[[],[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27"]]],[[],[["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_1"]]],[[],[["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"]]],[[],[["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6"]]],[[],[["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"]]],[[],[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_10","pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_0"]]],[[],[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_9","pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_1"]]],[[],[["pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_0","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2"]]],[[],[["pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_1","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1"]]],[[],[["pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_0","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2"]]],[[["pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1","pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_1"]],[]],[[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1"]],[]],[[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6","pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0"],["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"],["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]],[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"],["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]]],[[["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"],["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]],[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]]],[[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_0"],["pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2","pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_0"]],[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2"]]],[[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_1"]],[]],[[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_0"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_0"]],[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0"]]],[[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_1"]],[]],[[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0"]],[]],[[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6"]],[]],[[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]],[]],[[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]],[]],[[],[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"]]],[[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"]],[]],[[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"]],[]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0"]]],[[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3"]],[]],[[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2"]],[]],[[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0"]],[]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_0"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_1"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"]]],[[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]],[]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"]]],[[],[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6"]]],[[],[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4"]]],[[],[["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_5","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3"]]],[[],[["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_5"]]],[[],[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4"]]],[[],[["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4"]]],[[],[["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2"]]],[[],[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2"]]],[[],[["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_6","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1"]]],[[],[["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_6","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1"]]],[[],[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_7","pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_1"]]],[[],[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_8","pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_0"]]],[[],[["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28"]]],[[],[["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29"]]],[[],[["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32"]]],[[],[["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_2"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_1"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_1"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_0"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_0"]]],[[],[["pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_0","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_5"]]],[[],[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_7","pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_1"]]],[[],[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_5","pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_0"]]],[[],[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_7","pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_1"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"]]],[[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_0","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"]],[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"]]],[[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_1","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"]],[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"]]],[[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]],[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"],["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]]],[[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]],[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"],["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]]],[[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]],[]],[[],[["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]]],[[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]],[]],[[],[["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]]],[[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"]],[]],[[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"]],[]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"]]],[[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27"]],[]],[[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26"]],[]],[[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"]],[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"]]],[[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_5","pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_0"]],[]],[[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"]],[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"]]],[[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_7","pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_1"]],[]],[[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27"]],[]],[[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26"]],[]],[[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"]],[]],[[["pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_0","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_5"]],[]],[[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"]],[]],[[["pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_1","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_7"]],[]],[[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_10"]],[]],[[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_11"]],[]],[[["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5"]],[]],[[["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6"]],[]],[[["pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_1","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_7"]],[]],[[["pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_0","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_8"]],[]],[[["pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_1","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_9"]],[]],[[["pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_0","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_10"]],[]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_0"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_1"]]],[[],[["pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_31"]]],[[],[["pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_30"]]],[[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4"]],[]],[[],[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_4"]]],[[],[["pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_6"]]],[[],[["pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_7","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4"]]],[[["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4"]],[]],[[],[["pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_9","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4"]]],[[],[["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_5"]]],[[],[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_8"]]],[[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_0"]],[]],[[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_1"]],[]],[[["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_31","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_2"]],[]],[[["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_30","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_3"]],[]],[[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_4"]],[]],[[["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_5"]],[]],[[["pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_6"]],[]],[[["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_7"]],[]],[[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_8"]],[]],[[["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4","pin-type-component_fa65e0ca-1b7b-4bd0-8e4c-f8cae4988351_9"]],[]],[[],[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4"]]],[[],[["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2"]]],[[],[["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2","pin-type-component_ae34f7fd-5bf6-41c5-be78-9d886ea0cf65_0"]]],[[],[["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3","pin-type-component_ae34f7fd-5bf6-41c5-be78-9d886ea0cf65_1"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_ae34f7fd-5bf6-41c5-be78-9d886ea0cf65_2"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_ae34f7fd-5bf6-41c5-be78-9d886ea0cf65_3"]]],[[],[["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32","pin-type-component_ae34f7fd-5bf6-41c5-be78-9d886ea0cf65_4"]]],[[["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_5"]],[]],[[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_5"]],[]],[[],[["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28","pin-type-component_d357a112-8ce7-4ca7-922d-bae950c817be_1"]]],[[],[["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29","pin-type-component_e754101b-2bd4-45f8-8367-dd2d1465a844_1"]]],[[],[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1","pin-type-component_d357a112-8ce7-4ca7-922d-bae950c817be_3"]]],[[],[["pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1","pin-type-component_e754101b-2bd4-45f8-8367-dd2d1465a844_2"]]],[[],[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2","pin-type-component_e754101b-2bd4-45f8-8367-dd2d1465a844_2"]]],[[["pin-type-component_e754101b-2bd4-45f8-8367-dd2d1465a844_2","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1"]],[]],[[],[["pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1","pin-type-component_e754101b-2bd4-45f8-8367-dd2d1465a844_3"]]],[[],[["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2","pin-type-component_d357a112-8ce7-4ca7-922d-bae950c817be_2"]]],[[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_0"]],[]],[[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_1"]],[]],[[["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32"]],[]],[[["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28"]],[]],[[["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4"]],[]],[[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_6"]],[]],[[["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32"]],[]],[[["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29"]],[]],[[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4"]],[]],[[["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_6","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1"]],[]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_e754101b-2bd4-45f8-8367-dd2d1465a844_0"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_d357a112-8ce7-4ca7-922d-bae950c817be_0"]]],[[["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2","pin-type-component_ae34f7fd-5bf6-41c5-be78-9d886ea0cf65_0"]],[]],[[["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3","pin-type-component_ae34f7fd-5bf6-41c5-be78-9d886ea0cf65_1"]],[]],[[["pin-type-component_ae34f7fd-5bf6-41c5-be78-9d886ea0cf65_2","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[["pin-type-component_ae34f7fd-5bf6-41c5-be78-9d886ea0cf65_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_ae34f7fd-5bf6-41c5-be78-9d886ea0cf65_4","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32"]],[]],[[],[["pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_2"]]],[[],[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_2"]]],[[],[["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_1"]]],[[],[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_1"]]],[[],[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_0"]]],[[],[["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_0"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_3"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_3"]]],[[["pin-type-component_d357a112-8ce7-4ca7-922d-bae950c817be_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_d357a112-8ce7-4ca7-922d-bae950c817be_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28"]],[]],[[["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2","pin-type-component_d357a112-8ce7-4ca7-922d-bae950c817be_2"]],[]],[[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1","pin-type-component_d357a112-8ce7-4ca7-922d-bae950c817be_3"]],[]],[[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_e754101b-2bd4-45f8-8367-dd2d1465a844_0"]],[]],[[["pin-type-component_e754101b-2bd4-45f8-8367-dd2d1465a844_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29"]],[]],[[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2","pin-type-component_e754101b-2bd4-45f8-8367-dd2d1465a844_2"]],[]],[[["pin-type-component_e754101b-2bd4-45f8-8367-dd2d1465a844_3","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1"]],[]],[[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_2"]],[]],[[["pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_2","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1"]],[]],[[],[["pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_2","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1"]]],[[],[["pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_2","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1"]]],[[],[["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2","pin-type-component_ef73fc61-5332-4389-863a-156932dd9fb0_3"]]],[[],[["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3","pin-type-component_ef73fc61-5332-4389-863a-156932dd9fb0_2"]]],[[],[["pin-type-component_ef73fc61-5332-4389-863a-156932dd9fb0_0","pin-type-component_8774d229-a262-497a-8b8f-89515ac3c08c_2"]]],[[],[["pin-type-component_8774d229-a262-497a-8b8f-89515ac3c08c_3","pin-type-component_ef73fc61-5332-4389-863a-156932dd9fb0_1"]]],[[["pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[],[["pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_4","pin-type-component_8774d229-a262-497a-8b8f-89515ac3c08c_4"]]],[[],[["pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_3","pin-type-component_8774d229-a262-497a-8b8f-89515ac3c08c_5"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_8774d229-a262-497a-8b8f-89515ac3c08c_1"]]],[[],[["pin-type-component_8774d229-a262-497a-8b8f-89515ac3c08c_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29"]]],[[],[["pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_3","pin-type-component_15115ffa-76d4-4ac1-807f-112999c7cc8f_5"]]],[[],[["pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_4","pin-type-component_15115ffa-76d4-4ac1-807f-112999c7cc8f_4"]]],[[],[["pin-type-component_15115ffa-76d4-4ac1-807f-112999c7cc8f_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_15115ffa-76d4-4ac1-807f-112999c7cc8f_1"]]],[[],[["pin-type-component_ef73fc61-5332-4389-863a-156932dd9fb0_1","pin-type-component_15115ffa-76d4-4ac1-807f-112999c7cc8f_3"]]],[[],[["pin-type-component_ef73fc61-5332-4389-863a-156932dd9fb0_0","pin-type-component_15115ffa-76d4-4ac1-807f-112999c7cc8f_2"]]],[[["pin-type-component_15115ffa-76d4-4ac1-807f-112999c7cc8f_2","pin-type-component_ef73fc61-5332-4389-863a-156932dd9fb0_0"],["pin-type-component_8774d229-a262-497a-8b8f-89515ac3c08c_2","pin-type-component_ef73fc61-5332-4389-863a-156932dd9fb0_0"]],[["pin-type-component_15115ffa-76d4-4ac1-807f-112999c7cc8f_2","pin-type-component_8774d229-a262-497a-8b8f-89515ac3c08c_2"]]],[[["pin-type-component_15115ffa-76d4-4ac1-807f-112999c7cc8f_3","pin-type-component_ef73fc61-5332-4389-863a-156932dd9fb0_1"],["pin-type-component_8774d229-a262-497a-8b8f-89515ac3c08c_3","pin-type-component_ef73fc61-5332-4389-863a-156932dd9fb0_1"]],[["pin-type-component_15115ffa-76d4-4ac1-807f-112999c7cc8f_3","pin-type-component_8774d229-a262-497a-8b8f-89515ac3c08c_3"]]],[[["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3","pin-type-component_ef73fc61-5332-4389-863a-156932dd9fb0_2"]],[]],[[["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2","pin-type-component_ef73fc61-5332-4389-863a-156932dd9fb0_3"]],[]],[[["pin-type-component_8774d229-a262-497a-8b8f-89515ac3c08c_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29"]],[]],[[["pin-type-component_8774d229-a262-497a-8b8f-89515ac3c08c_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_15115ffa-76d4-4ac1-807f-112999c7cc8f_2","pin-type-component_8774d229-a262-497a-8b8f-89515ac3c08c_2"]],[]],[[["pin-type-component_15115ffa-76d4-4ac1-807f-112999c7cc8f_3","pin-type-component_8774d229-a262-497a-8b8f-89515ac3c08c_3"]],[]],[[["pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_4","pin-type-component_8774d229-a262-497a-8b8f-89515ac3c08c_4"]],[]],[[["pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_3","pin-type-component_8774d229-a262-497a-8b8f-89515ac3c08c_5"]],[]],[[["pin-type-component_15115ffa-76d4-4ac1-807f-112999c7cc8f_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28"]],[]],[[["pin-type-component_15115ffa-76d4-4ac1-807f-112999c7cc8f_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_15115ffa-76d4-4ac1-807f-112999c7cc8f_4","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_4"]],[]],[[["pin-type-component_15115ffa-76d4-4ac1-807f-112999c7cc8f_5","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_3"]],[]],[[],[["pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_0","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_3"]]],[[],[["pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_0","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_3"]]],[[],[["pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_1","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_4"]]],[[],[["pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_2","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_4"]]],[[],[["pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_6","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5"]]],[[],[["pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_5","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_3"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_4"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0":"0000000000000000","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1":"0000000000000001","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2":"0000000000000011","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3":"0000000000000010","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_0":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_1":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2":"0000000000000016","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_3":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_4":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5":"0000000000000015","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_6":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_7":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_8":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_9":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_10":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_11":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_12":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_13":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_14":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_15":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_16":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_17":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_18":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19":"0000000000000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_20":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_21":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_22":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_23":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24":"0000000000000001","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_25":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_30":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_31":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_33":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_34":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_35":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_36":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_37":"_","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_0":"_","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1":"0000000000000006","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2":"0000000000000012","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_0":"_","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1":"0000000000000007","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2":"0000000000000013","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0":"0000000000000004","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1":"0000000000000005","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0":"0000000000000004","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1":"0000000000000005","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2":"0000000000000002","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3":"0000000000000012","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0":"0000000000000004","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1":"0000000000000005","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2":"0000000000000003","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3":"0000000000000013","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0":"0000000000000004","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1":"0000000000000005","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2":"0000000000000010","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3":"0000000000000011","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_0":"0000000000000003","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_1":"0000000000000013","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_2":"0000000000000007","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_3":"0000000000000008","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_4":"0000000000000014","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_5":"_","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_6":"_","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_7":"_","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_8":"_","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_0":"0000000000000002","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_1":"0000000000000012","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_2":"0000000000000006","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_3":"0000000000000008","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_4":"0000000000000009","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_5":"_","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_6":"_","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_7":"_","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_8":"_","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_0":"0000000000000008","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_1":"0000000000000009","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_2":"0000000000000014","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_3":"0000000000000000","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_4":"0000000000000001","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_5":"0000000000000016","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_6":"0000000000000015"},"component_id_to_pins":{"d53bc8d1-adbf-42c3-9bdc-27d4d2b68588":["0","1","2","3"],"f7d25e04-bb51-41df-ba72-c452c270d3fb":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31","32","33","34","35","36","37"],"32608709-bcb5-4c22-82f1-0b5ac1739be0":[],"915b317b-63a4-4c37-8362-9a35870cbe7c":[],"9e0cc72b-cce0-4555-8c60-9928baea3faa":[],"41689d80-6f1a-478b-ad5a-826ce578b4af":[],"ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8":["0","1","2"],"00e3d6c2-f801-4d91-ad4d-237bada773bb":["0","1","2"],"1c19cc90-e27a-4c31-a566-dce6d12cc7bd":["0","1"],"8b4859a0-119b-4d24-8c3e-f008f1af2f35":[],"eb1dbc1c-94ee-4954-b264-2ba5f2bb6c04":[],"060f78c2-f7c5-4b91-a54e-26722a6a6eb1":["0","1","2","3"],"c483e859-dbe3-40ab-ad85-fdb0e9726a1e":["0","1","2","3"],"786922c4-3cc4-4e2e-a1af-6f582a726cc5":[],"c6b89f01-cd33-4f53-a410-bd8ce0a19726":[],"028c5ed6-a9ce-4916-bd5a-20a0af91ff53":[],"d8ee4efe-302f-41eb-a87d-4235620299ce":[],"8c415f8f-024b-42a7-9906-fa5d9103b190":[],"f0886e27-8ec0-43da-a659-1cbab4912d9c":[],"9b271475-bebe-41b8-aded-20e21ef4734b":["0","1","2","3"],"60b47335-97ed-4e17-861d-700ea31fb823":[],"90939bc7-e151-4981-b49e-514d89d01342":["0","1","2","3","4","5","6","7","8"],"38451353-a24a-49a0-9b0c-182de089686c":["0","1","2","3","4","5","6","7","8"],"6a48dac8-9f96-4aac-a57d-699995a9514a":[],"4ba86a89-927e-476a-9b47-f0cc93744701":[],"3f2e1968-f0b0-44f3-809d-425515dc44c8":[],"248c3be1-2437-4b67-8bd8-26d79162e2f2":[],"5c70012d-03f5-42a2-a7be-1acfd998eb4c":["0","1","2","3","4","5","6"]},"uid_to_net":{"_":[],"0000000000000001":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_4"],"0000000000000000":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_3"],"0000000000000004":["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"],"0000000000000005":["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"],"0000000000000010":["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"],"0000000000000011":["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"],"0000000000000012":["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_1"],"0000000000000013":["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_1"],"0000000000000002":["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_0"],"0000000000000003":["pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2"],"0000000000000006":["pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_2","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1"],"0000000000000007":["pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_2","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1"],"0000000000000008":["pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_3","pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_0","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_3"],"0000000000000009":["pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_1","pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_4"],"0000000000000014":["pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_2","pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_4"],"0000000000000015":["pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_6","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5"],"0000000000000016":["pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_5","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2"]},"uid_to_text_label":{"0000000000000001":"Net 1","0000000000000000":"Net 0","0000000000000004":"Net 4","0000000000000005":"Net 5","0000000000000010":"Net 10","0000000000000011":"Net 11","0000000000000012":"Net 12","0000000000000013":"Net 13","0000000000000002":"Net 2","0000000000000003":"Net 3","0000000000000006":"Net 6","0000000000000007":"Net 7","0000000000000008":"Net 8","0000000000000009":"Net 9","0000000000000014":"Net 14","0000000000000015":"Net 15","0000000000000016":"Net 16"},"all_breadboard_info_list":[],"breadboard_info_list":[],"componentsData":[{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"GND","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[3499.592122094968,381.2251000087314],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"32608709-bcb5-4c22-82f1-0b5ac1739be0","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"VCC +5V","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[3366.1168313046355,378.8059167969202],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"915b317b-63a4-4c37-8362-9a35870cbe7c","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[816.5526985000006,-399.1880574999998],"typeId":"b975acdd-73e3-4b18-a5a5-9b66f369afa0","componentVersion":2,"instanceId":"f7d25e04-bb51-41df-ba72-c452c270d3fb","orientation":"up","circleData":[[947.5,-625],[948.1030000000001,-597.7392055],[948.1231135000003,-571.7030244999999],[947.5,-543.2146149999999],[948.7261135000003,-517.1784339999997],[947.5,-491.1221394999996],[948.7261135000003,-463.25684499999954],[948.7261135000003,-437.22066399999966],[948.7261135000003,-409.95986949999957],[948.1030000000001,-384.5506884999996],[949.3291135000004,-356.6853939999997],[949.3291135000004,-329.4230994999997],[949.3291135000004,-301.56169149999965],[949.9306135000002,-275.52701049999956],[949.3291135000004,-249.5109429999997],[950.5552270000003,-220.39941999999974],[949.9306135000002,-194.36323900000002],[949.9306135000002,-166.47783100000015],[951.7813405000002,-138.01103649999993],[678.5382805000002,-136.80653649999988],[677.312167,-164.67033100000003],[678.5382805000002,-190.70651199999998],[677.9352805000001,-218.5703064999999],[677.9352805000001,-245.8326009999999],[679.1613940000002,-272.4717834999995],[678.5382805000002,-299.1310779999997],[679.1613940000002,-328.24259949999976],[677.9352805000001,-355.4832804999997],[677.9352805000001,-380.91646149999957],[677.3322805000003,-406.9526424999996],[677.3322805000003,-434.8179369999996],[677.312167,-461.45323149999956],[678.5583940000001,-488.71402599999954],[677.3322805000003,-514.7300934999996],[675.4824745000001,-543.8420259999998],[677.3322805000003,-569.294911],[677.9349745000002,-595.913026],[677.3322805000003,-623.7738865000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"LOAD 1 AC Circuit\n(behind a breaker)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[2521.1223679499117,1492.667604045154],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"9e0cc72b-cce0-4555-8c60-9928baea3faa","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"LOAD 2 AC Circuit\n(behind a breaker)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[2767.5835720784066,1691.9991453659359],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"41689d80-6f1a-478b-ad5a-826ce578b4af","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[3123.2036904999995,1157.474882],"typeId":"5ac8a9e5-bb24-45ef-9b03-1161364522fb","componentVersion":1,"instanceId":"1c19cc90-e27a-4c31-a566-dce6d12cc7bd","orientation":"up","circleData":[[2987.5,1145],[3259.5265,1145]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Main line\n(phase) - L\n(Enedis in France)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[3292.519774875356,1084.5794073453549],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"8b4859a0-119b-4d24-8c3e-f008f1af2f35","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Main neutral - N\n(Enedis in France)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[2953.4352836968415,1091.5820712351226],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"eb1dbc1c-94ee-4954-b264-2ba5f2bb6c04","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[2528.8436755,1583.142836],"typeId":"a64016c8-4d9c-491e-ba46-f626b2aeb38c","componentVersion":1,"instanceId":"060f78c2-f7c5-4b91-a54e-26722a6a6eb1","orientation":"up","circleData":[[2507.5,1430],[2544.3571255,1429.1428745],[2545.6428145,1755.2857490000001],[2509.6428145,1753.1428744999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[2768.8436755000002,1778.142836],"typeId":"a64016c8-4d9c-491e-ba46-f626b2aeb38c","componentVersion":1,"instanceId":"c483e859-dbe3-40ab-ad85-fdb0e9726a1e","orientation":"up","circleData":[[2747.5,1625],[2784.3571255000006,1624.1428745],[2785.6428145,1950.2857490000008],[2749.6428145,1948.1428745000005]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"N","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[3393.359241444308,610.2637795986323],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"786922c4-3cc4-4e2e-a1af-6f582a726cc5","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"L","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[3497.068721174747,610.9967802938991],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"c6b89f01-cd33-4f53-a410-bd8ce0a19726","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"LOAD 1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[617.3731045635486,2550.7608732631475],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"028c5ed6-a9ce-4916-bd5a-20a0af91ff53","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"LOAD 2","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[1334.8501274033324,2570.197610023702],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"d8ee4efe-302f-41eb-a87d-4235620299ce","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Dimmer\nOutput 2","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[1690.0171129740847,1041.5458167416323],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"8c415f8f-024b-42a7-9906-fa5d9103b190","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Dimmer\nOutput 1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[1682.0326352223556,444.3766791468882],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"f0886e27-8ec0-43da-a659-1cbab4912d9c","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[3006.71431,2014.5000244999999],"typeId":"5ce5e9a0-0484-4e7a-b171-46d0c4edfd48","componentVersion":2,"instanceId":"9b271475-bebe-41b8-aded-20e21ef4734b","orientation":"up","circleData":[[2987.5,1850],[3029.499982,1850.8571344999998],[2986.6428895,2182.999983499998],[3030.7857474999996,2183.8571599999987]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"YaSolR AC Circuit\n(behind a breaker)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[3012.4637827603738,1911.511553397949],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"60b47335-97ed-4e17-861d-700ea31fb823","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[3442.3552975000002,484.8953134999997],"typeId":"c2a09f2b-df40-42a6-8e0c-c519ba38e9d5","componentVersion":1,"instanceId":"d53bc8d1-adbf-42c3-9bdc-27d4d2b68588","orientation":"up","circleData":[[3437.5,350],[3453.0759055000003,351.3743885],[3453.9921460000005,604.2539555000001],[3440.706811,605.6282870000002]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[736.6917940000035,2642.799167000001],"typeId":"fa95e5d1-b92a-410f-a873-a71d0089e7ad","componentVersion":1,"instanceId":"ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8","orientation":"left","circleData":[[2942.5,-880],[752.5000000000027,2375.000000000001],[782.5000000000027,2375.000000000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1426.6917939999958,2657.799166999998],"typeId":"fa95e5d1-b92a-410f-a873-a71d0089e7ad","componentVersion":1,"instanceId":"00e3d6c2-f801-4d91-ad4d-237bada773bb","orientation":"left","circleData":[[3632.5,-865],[1442.4999999999945,2389.999999999997],[1472.4999999999936,2389.999999999997]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1694.5013439999998,1208.1596720000002],"typeId":"698fdeba-91ca-4b68-9d55-5545583fbf52","componentVersion":2,"instanceId":"90939bc7-e151-4981-b49e-514d89d01342","orientation":"up","circleData":[[1577.5,1040],[1805.7023815000002,1033.274981],[1578.8449794999997,1375.802756000001],[1434.4812009999996,1227.8522630000002],[1432.9845669999995,1196.4688385000002],[1434.4809999999998,1256.7830000000004],[1433.5839999999998,1137.5255000000002],[1434.4809999999998,1167.1160000000002],[1434.0325000000003,1284.5795000000007]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1679.5013439999998,608.1596720000005],"typeId":"698fdeba-91ca-4b68-9d55-5545583fbf52","componentVersion":2,"instanceId":"38451353-a24a-49a0-9b0c-182de089686c","orientation":"up","circleData":[[1562.5,440],[1790.7023814999998,433.274981],[1563.8449795,775.8027559999998],[1419.481201,627.8522630000002],[1417.984567,596.4688385000002],[1419.4810000000002,656.7829999999999],[1418.5839999999998,537.5255000000002],[1419.4810000000002,567.1160000000002],[1419.0324999999998,684.5795000000003]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"N","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[1867.1748476958887,1041.869364359734],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"6a48dac8-9f96-4aac-a57d-699995a9514a","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"LOAD2","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[1484.8216804677136,1376.6664141576466],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"4ba86a89-927e-476a-9b47-f0cc93744701","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"N","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[1864.3224710709637,433.0731522084204],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"3f2e1968-f0b0-44f3-809d-425515dc44c8","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"LOAD1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[1461.8928514608904,775.1707301452052],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"248c3be1-2437-4b67-8bd8-26d79162e2f2","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[387.90041499999995,907.6559224999999],"typeId":"7b6ceb33-1206-44c4-8e9b-79797c6b533a","componentVersion":3,"instanceId":"5c70012d-03f5-42a2-a7be-1acfd998eb4c","orientation":"down","circleData":[[467.5,905],[468.397,874.961],[469.29699999999997,934.5905],[287.71773699999994,924.726773],[287.80879899999996,912.6146855],[287.80879899999996,900.9579725],[287.3604535,889.3013195]],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"-894.00000","left":"273.36045","width":"3373.13955","height":"3857.07477","x":"273.36045","y":"-894.00000"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1\",\"endPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24\",\"rawStartPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1\",\"rawEndPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"3453.0759055000_351.3743885000\\\",\\\"3453.0759055000_260.0000000000\\\",\\\"640.0000000000_260.0000000000\\\",\\\"640.0000000000_-272.4717835000\\\",\\\"679.1613940000_-272.4717835000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_4\",\"endPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1\",\"rawStartPinId\":\"pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_4\",\"rawEndPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"287.8087990000_912.6146855000\\\",\\\"130.0000000000_912.6146855000\\\",\\\"130.0000000000_260.0000000000\\\",\\\"3452.5000000000_260.0000000000\\\",\\\"3452.5000000000_351.3743885000\\\",\\\"3453.0759055000_351.3743885000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0\",\"endPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19\",\"rawStartPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0\",\"rawEndPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"3437.5000000000_350.0000000000\\\",\\\"3437.5000000000_282.5000000000\\\",\\\"617.5000000000_282.5000000000\\\",\\\"617.5000000000_-136.8065365000\\\",\\\"678.5382805000_-136.8065365000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_3\",\"endPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0\",\"rawStartPinId\":\"pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_3\",\"rawEndPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"287.7177370000_924.7267730000\\\",\\\"100.0000000000_924.7267730000\\\",\\\"100.0000000000_282.5000000000\\\",\\\"3437.5000000000_282.5000000000\\\",\\\"3437.5000000000_350.0000000000\\\"]}\"}","{\"color\":\"#0076FF\",\"startPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0\",\"endPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0\",\"rawStartPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0\",\"rawEndPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2987.5000000000_1145.0000000000\\\",\\\"2747.5000000000_1145.0000000000\\\",\\\"2747.5000000000_1625.0000000000\\\"]}\"}","{\"color\":\"#0076FF\",\"startPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0\",\"endPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0\",\"rawStartPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0\",\"rawEndPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2507.5000000000_1430.0000000000\\\",\\\"2507.5000000000_1145.0000000000\\\",\\\"2987.5000000000_1145.0000000000\\\"]}\"}","{\"color\":\"#0076FF\",\"startPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0\",\"endPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0\",\"rawStartPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0\",\"rawEndPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2987.5000000000_1145.0000000000\\\",\\\"2987.5000000000_1850.0000000000\\\"]}\"}","{\"color\":\"#85A900\",\"startPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1\",\"endPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1\",\"rawStartPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1\",\"rawEndPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2544.3571255000_1429.1428745000\\\",\\\"2544.3571255000_1310.0000000000\\\",\\\"3317.5000000000_1310.0000000000\\\",\\\"3317.5000000000_1145.0000000000\\\",\\\"3259.5265000000_1145.0000000000\\\"]}\"}","{\"color\":\"#85A900\",\"startPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1\",\"endPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1\",\"rawStartPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1\",\"rawEndPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"3259.5265000000_1145.0000000000\\\",\\\"3317.5000000000_1145.0000000000\\\",\\\"3317.5000000000_1310.0000000000\\\",\\\"2784.3571255000_1310.0000000000\\\",\\\"2784.3571255000_1624.1428745000\\\"]}\"}","{\"color\":\"#85A900\",\"startPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1\",\"endPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1\",\"rawStartPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1\",\"rawEndPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"3259.5265000000_1145.0000000000\\\",\\\"3317.5000000000_1145.0000000000\\\",\\\"3317.5000000000_1310.0000000000\\\",\\\"3032.5000000000_1310.0000000000\\\",\\\"3032.5000000000_1850.8571345000\\\",\\\"3029.4999820000_1850.8571345000\\\"]}\"}","{\"color\":\"#00FFC6\",\"startPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2\",\"endPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3\",\"rawStartPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2\",\"rawEndPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2986.6428895000_2182.9999835000\\\",\\\"2986.6428895000_2262.5000000000\\\",\\\"3437.5000000000_2262.5000000000\\\",\\\"3437.5000000000_605.6282870000\\\",\\\"3440.7068110000_605.6282870000\\\"]}\"}","{\"color\":\"#FF6E41\",\"startPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3\",\"endPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2\",\"rawStartPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3\",\"rawEndPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"3030.7857475000_2183.8571600000\\\",\\\"3032.5000000000_2183.8571600000\\\",\\\"3032.5000000000_2277.5000000000\\\",\\\"3453.9921460000_2277.5000000000\\\",\\\"3453.9921460000_604.2539555000\\\"]}\"}","{\"color\":\"#E85EBE\",\"startPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3\",\"endPinId\":\"pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2\",\"rawStartPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3\",\"rawEndPinId\":\"pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2509.6428145000_1753.1428745000\\\",\\\"2509.6428145000_1895.0000000000\\\",\\\"782.5000000000_1895.0000000000\\\",\\\"782.5000000000_2375.0000000000\\\"]}\"}","{\"color\":\"#E85EBE\",\"startPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3\",\"endPinId\":\"pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_1\",\"rawStartPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3\",\"rawEndPinId\":\"pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2509.6428145000_1753.1428745000\\\",\\\"2509.6428145000_1895.0000000000\\\",\\\"2177.5000000000_1895.0000000000\\\",\\\"2177.5000000000_365.0000000000\\\",\\\"1790.7023815000_365.0000000000\\\",\\\"1790.7023815000_433.2749810000\\\"]}\"}","{\"color\":\"#010067\",\"startPinId\":\"pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2\",\"endPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3\",\"rawStartPinId\":\"pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2\",\"rawEndPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1472.5000000000_2390.0000000000\\\",\\\"1472.5000000000_2165.0000000000\\\",\\\"2749.6428145000_2165.0000000000\\\",\\\"2749.6428145000_1948.1428745000\\\"]}\"}","{\"color\":\"#010067\",\"startPinId\":\"pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_1\",\"endPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3\",\"rawStartPinId\":\"pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_1\",\"rawEndPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1805.7023815000_1033.2749810000\\\",\\\"1805.7023815000_957.5000000000\\\",\\\"2042.5000000000_957.5000000000\\\",\\\"2042.5000000000_2165.0000000000\\\",\\\"2749.6428145000_2165.0000000000\\\",\\\"2749.6428145000_1948.1428745000\\\"]}\"}","{\"color\":\"#A75740\",\"startPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2\",\"endPinId\":\"pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_0\",\"rawStartPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2\",\"rawEndPinId\":\"pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2545.6428145000_1755.2857490000\\\",\\\"2545.6428145000_1865.0000000000\\\",\\\"2207.5000000000_1865.0000000000\\\",\\\"2207.5000000000_335.0000000000\\\",\\\"1562.5000000000_335.0000000000\\\",\\\"1562.5000000000_440.0000000000\\\"]}\"}","{\"color\":\"#01FFFE\",\"startPinId\":\"pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_0\",\"endPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2\",\"rawStartPinId\":\"pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_0\",\"rawEndPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1577.5000000000_1040.0000000000\\\",\\\"1577.5000000000_927.5000000000\\\",\\\"2072.5000000000_927.5000000000\\\",\\\"2072.5000000000_2127.5000000000\\\",\\\"2785.6428145000_2127.5000000000\\\",\\\"2785.6428145000_1950.2857490000\\\"]}\"}","{\"color\":\"#BDC6FF\",\"startPinId\":\"pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_2\",\"endPinId\":\"pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1\",\"rawStartPinId\":\"pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_2\",\"rawEndPinId\":\"pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1563.8449795000_775.8027560000\\\",\\\"1563.8449795000_860.0000000000\\\",\\\"752.5000000000_860.0000000000\\\",\\\"752.5000000000_2375.0000000000\\\"]}\"}","{\"color\":\"#BB8800\",\"startPinId\":\"pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1\",\"endPinId\":\"pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_2\",\"rawStartPinId\":\"pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1\",\"rawEndPinId\":\"pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1442.5000000000_2390.0000000000\\\",\\\"1442.5000000000_1467.5000000000\\\",\\\"1578.8449795000_1467.5000000000\\\",\\\"1578.8449795000_1375.8027560000\\\"]}\"}","{\"color\":\"#FFDB66\",\"startPinId\":\"pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_3\",\"endPinId\":\"pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_0\",\"rawStartPinId\":\"pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_3\",\"rawEndPinId\":\"pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1419.4812010000_627.8522630000\\\",\\\"550.0000000000_627.8522630000\\\",\\\"550.0000000000_905.0000000000\\\",\\\"467.5000000000_905.0000000000\\\"]}\"}","{\"color\":\"#FFDB66\",\"startPinId\":\"pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_0\",\"endPinId\":\"pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_3\",\"rawStartPinId\":\"pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_0\",\"rawEndPinId\":\"pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"467.5000000000_905.0000000000\\\",\\\"550.0000000000_905.0000000000\\\",\\\"550.0000000000_1227.8522630000\\\",\\\"1434.4812010000_1227.8522630000\\\"]}\"}","{\"color\":\"#90FB92\",\"startPinId\":\"pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_4\",\"endPinId\":\"pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_1\",\"rawStartPinId\":\"pin-type-component_38451353-a24a-49a0-9b0c-182de089686c_4\",\"rawEndPinId\":\"pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1417.9845670000_596.4688385000\\\",\\\"520.0000000000_596.4688385000\\\",\\\"520.0000000000_874.9610000000\\\",\\\"468.3970000000_874.9610000000\\\"]}\"}","{\"color\":\"#7E2DD2\",\"startPinId\":\"pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_2\",\"endPinId\":\"pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_4\",\"rawStartPinId\":\"pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_2\",\"rawEndPinId\":\"pin-type-component_90939bc7-e151-4981-b49e-514d89d01342_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"469.2970000000_934.5905000000\\\",\\\"520.0000000000_934.5905000000\\\",\\\"520.0000000000_1196.4688385000\\\",\\\"1432.9845670000_1196.4688385000\\\"]}\"}","{\"color\":\"#BDD393\",\"startPinId\":\"pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_6\",\"endPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5\",\"rawStartPinId\":\"pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_6\",\"rawEndPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"287.3604535000_889.3013195000\\\",\\\"190.0000000000_889.3013195000\\\",\\\"190.0000000000_-737.5000000000\\\",\\\"1030.0000000000_-737.5000000000\\\",\\\"1030.0000000000_-491.1221395000\\\",\\\"947.5000000000_-491.1221395000\\\"]}\"}","{\"color\":\"#E56FFE\",\"startPinId\":\"pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_5\",\"endPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2\",\"rawStartPinId\":\"pin-type-component_5c70012d-03f5-42a2-a7be-1acfd998eb4c_5\",\"rawEndPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"287.8087990000_900.9579725000\\\",\\\"160.0000000000_900.9579725000\\\",\\\"160.0000000000_-767.5000000000\\\",\\\"1060.0000000000_-767.5000000000\\\",\\\"1060.0000000000_-571.7030245000\\\",\\\"948.1231135000_-571.7030245000\\\"]}\"}"],"projectDescription":""}PK
     #{dZ               jsons/PK
     #{dZR�1FPt  Pt     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"ESP32 Devkit V4","category":["User Defined"],"id":"b975acdd-73e3-4b18-a5a5-9b66f369afa0","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"ae82c023-d9d4-4942-aa8d-ab2ae3c53d73.png","iconPic":"cbf7ad0e-0f08-44f8-98a9-dcbe92af212f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"48.00864","numDisplayRows":"48.00864","pins":[{"uniquePinIdString":"0","positionMil":"3273.41401,3905.84495","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"3277.43401,3724.10632","isAnchorPin":false,"label":"23"},{"uniquePinIdString":"2","positionMil":"3277.56810,3550.53178","isAnchorPin":false,"label":"22"},{"uniquePinIdString":"3","positionMil":"3273.41401,3360.60905","isAnchorPin":false,"label":"TX"},{"uniquePinIdString":"4","positionMil":"3281.58810,3187.03451","isAnchorPin":false,"label":"RX"},{"uniquePinIdString":"5","positionMil":"3273.41401,3013.32588","isAnchorPin":false,"label":"21"},{"uniquePinIdString":"6","positionMil":"3281.58810,2827.55725","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"7","positionMil":"3281.58810,2653.98271","isAnchorPin":false,"label":"19"},{"uniquePinIdString":"8","positionMil":"3281.58810,2472.24408","isAnchorPin":false,"label":"18"},{"uniquePinIdString":"9","positionMil":"3277.43401,2302.84954","isAnchorPin":false,"label":"5"},{"uniquePinIdString":"10","positionMil":"3285.60810,2117.08091","isAnchorPin":false,"label":"17"},{"uniquePinIdString":"11","positionMil":"3285.60810,1935.33228","isAnchorPin":false,"label":"16"},{"uniquePinIdString":"12","positionMil":"3285.60810,1749.58956","isAnchorPin":false,"label":"4"},{"uniquePinIdString":"13","positionMil":"3289.61810,1576.02502","isAnchorPin":false,"label":"0"},{"uniquePinIdString":"14","positionMil":"3285.60810,1402.58457","isAnchorPin":false,"label":"2"},{"uniquePinIdString":"15","positionMil":"3293.78219,1208.50775","isAnchorPin":false,"label":"15"},{"uniquePinIdString":"16","positionMil":"3289.61810,1034.93321","isAnchorPin":false,"label":"D1"},{"uniquePinIdString":"17","positionMil":"3289.61810,849.03049","isAnchorPin":false,"label":"D0"},{"uniquePinIdString":"18","positionMil":"3301.95628,659.25186","isAnchorPin":false,"label":"CLK"},{"uniquePinIdString":"19","positionMil":"1480.33588,651.22186","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"20","positionMil":"1472.16179,836.98049","isAnchorPin":false,"label":"CMD"},{"uniquePinIdString":"21","positionMil":"1480.33588,1010.55503","isAnchorPin":false,"label":"D3"},{"uniquePinIdString":"22","positionMil":"1476.31588,1196.31366","isAnchorPin":false,"label":"D2"},{"uniquePinIdString":"23","positionMil":"1476.31588,1378.06229","isAnchorPin":false,"label":"13"},{"uniquePinIdString":"24","positionMil":"1484.48997,1555.65684","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"25","positionMil":"1480.33588,1733.38547","isAnchorPin":false,"label":"12"},{"uniquePinIdString":"26","positionMil":"1484.48997,1927.46228","isAnchorPin":false,"label":"14"},{"uniquePinIdString":"27","positionMil":"1476.31588,2109.06682","isAnchorPin":false,"label":"27"},{"uniquePinIdString":"28","positionMil":"1476.31588,2278.62136","isAnchorPin":false,"label":"26"},{"uniquePinIdString":"29","positionMil":"1472.29588,2452.19590","isAnchorPin":false,"label":"25"},{"uniquePinIdString":"30","positionMil":"1472.29588,2637.96453","isAnchorPin":false,"label":"33"},{"uniquePinIdString":"31","positionMil":"1472.16179,2815.53316","isAnchorPin":false,"label":"32"},{"uniquePinIdString":"32","positionMil":"1480.46997,2997.27179","isAnchorPin":false,"label":"35"},{"uniquePinIdString":"33","positionMil":"1472.29588,3170.71224","isAnchorPin":false,"label":"34"},{"uniquePinIdString":"34","positionMil":"1459.96384,3364.79179","isAnchorPin":false,"label":"VIN"},{"uniquePinIdString":"35","positionMil":"1472.29588,3534.47769","isAnchorPin":false,"label":"VP"},{"uniquePinIdString":"36","positionMil":"1476.31384,3711.93179","isAnchorPin":false,"label":"EN"},{"uniquePinIdString":"37","positionMil":"1472.29588,3897.67086","isAnchorPin":false,"label":"3V3"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Alternative Current (AC) - Large","category":["User Defined"],"id":"5ac8a9e5-bb24-45ef-9b03-1161364522fb","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"8a1d81a5-79d4-450c-9f72-108cd2673013.png","iconPic":"aacc0029-e57d-4614-a443-d9bee65b5175.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"23.63677","numDisplayRows":"22.90067","pins":[{"uniquePinIdString":"0","positionMil":"277.14723,1228.19938","isAnchorPin":true,"label":"Neutral"},{"uniquePinIdString":"1","positionMil":"2090.65723,1228.19938","isAnchorPin":false,"label":"Line"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Breaker 20A","category":["User Defined"],"id":"a64016c8-4d9c-491e-ba46-f626b2aeb38c","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1d90a712-93d7-4555-ae10-1782f839eba3.png","iconPic":"e5551f5a-2fb7-4493-9527-57db21faeaae.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.69291","numDisplayRows":"28.74016","pins":[{"uniquePinIdString":"0","positionMil":"192.35433,2457.96024","isAnchorPin":true,"label":"N"},{"uniquePinIdString":"1","positionMil":"438.06850,2463.67441","isAnchorPin":false,"label":"L"},{"uniquePinIdString":"2","positionMil":"446.63976,289.38858","isAnchorPin":false,"label":"L"},{"uniquePinIdString":"3","positionMil":"206.63976,303.67441","isAnchorPin":false,"label":"N"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Breaker 20A","category":["User Defined"],"id":"a64016c8-4d9c-491e-ba46-f626b2aeb38c","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1d90a712-93d7-4555-ae10-1782f839eba3.png","iconPic":"e5551f5a-2fb7-4493-9527-57db21faeaae.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.69291","numDisplayRows":"28.74016","pins":[{"uniquePinIdString":"0","positionMil":"192.35433,2457.96024","isAnchorPin":true,"label":"N"},{"uniquePinIdString":"1","positionMil":"438.06850,2463.67441","isAnchorPin":false,"label":"L"},{"uniquePinIdString":"2","positionMil":"446.63976,289.38858","isAnchorPin":false,"label":"L"},{"uniquePinIdString":"3","positionMil":"206.63976,303.67441","isAnchorPin":false,"label":"N"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Breaker 2A","category":["User Defined"],"id":"5ce5e9a0-0484-4e7a-b171-46d0c4edfd48","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"a038ca8d-f9eb-4e93-ad0b-b831193aa106.png","iconPic":"3e0a96b2-ef1c-4fb2-8b57-d71cbe1f3744.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"28.33333","pins":[{"uniquePinIdString":"0","positionMil":"205.23810,2513.33333","isAnchorPin":true,"label":"N"},{"uniquePinIdString":"1","positionMil":"485.23798,2507.61910","isAnchorPin":false,"label":"L"},{"uniquePinIdString":"2","positionMil":"199.52403,293.33344","isAnchorPin":false,"label":"N"},{"uniquePinIdString":"3","positionMil":"493.80975,287.61893","isAnchorPin":false,"label":"L"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"HDR-15-5 5V 2.4A","category":["User Defined"],"id":"c2a09f2b-df40-42a6-8e0c-c519ba38e9d5","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"cff7cff8-0125-49f3-ae91-9e6ccc0a4cc7.png","iconPic":"7b19d218-2217-455d-9a43-b73a208c2c5c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.54331","numDisplayRows":"21.25984","pins":[{"uniquePinIdString":"0","positionMil":"144.79685,1962.29409","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"248.63622,1953.13150","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"2","positionMil":"254.74449,267.26772","isAnchorPin":false,"label":"L"},{"uniquePinIdString":"3","positionMil":"166.17559,258.10551","isAnchorPin":false,"label":"N"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Water Heater","category":["User Defined"],"id":"fa95e5d1-b92a-410f-a873-a71d0089e7ad","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"85e66502-362d-4a26-afcd-97fbc4859675.png","iconPic":"b13518ba-21c5-4f60-a735-1d8041d11d7b.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"39.37008","numDisplayRows":"39.37008","pins":[{"uniquePinIdString":"0","positionMil":"25453.83178,-12736.88404","isAnchorPin":true,"label":""},{"uniquePinIdString":"1","positionMil":"3753.83178,1863.11596","isAnchorPin":false,"label":"V+"},{"uniquePinIdString":"2","positionMil":"3753.83178,1663.11596","isAnchorPin":false,"label":"V-"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Water Heater","category":["User Defined"],"id":"fa95e5d1-b92a-410f-a873-a71d0089e7ad","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"85e66502-362d-4a26-afcd-97fbc4859675.png","iconPic":"b13518ba-21c5-4f60-a735-1d8041d11d7b.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"39.37008","numDisplayRows":"39.37008","pins":[{"uniquePinIdString":"0","positionMil":"25453.83178,-12736.88404","isAnchorPin":true,"label":""},{"uniquePinIdString":"1","positionMil":"3753.83178,1863.11596","isAnchorPin":false,"label":"V+"},{"uniquePinIdString":"2","positionMil":"3753.83178,1663.11596","isAnchorPin":false,"label":"V-"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Loncont LSA-H3P50YB","category":["User Defined"],"id":"698fdeba-91ca-4b68-9d55-5545583fbf52","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"c750f18a-9432-41e6-a6ed-179e28bc29f6.png","iconPic":"3f9b3f3f-db41-4a6d-b13c-7e86a7741a7b.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"40.94488","numDisplayRows":"29.13386","pins":[{"uniquePinIdString":"0","positionMil":"1267.23504,2577.75748","isAnchorPin":true,"label":"L"},{"uniquePinIdString":"1","positionMil":"2788.58425,2622.59094","isAnchorPin":false,"label":"N"},{"uniquePinIdString":"2","positionMil":"1276.20157,339.07244","isAnchorPin":false,"label":"LOAD"},{"uniquePinIdString":"3","positionMil":"313.77638,1325.40906","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"4","positionMil":"303.79882,1534.63189","isAnchorPin":false,"label":"VCC 0-10V"},{"uniquePinIdString":"5","positionMil":"313.77504,1132.53748","isAnchorPin":false,"label":"VCC 0-5V"},{"uniquePinIdString":"6","positionMil":"307.79504,1927.58748","isAnchorPin":false,"label":"PWM"},{"uniquePinIdString":"7","positionMil":"313.77504,1730.31748","isAnchorPin":false,"label":"VCC 4-20mA"},{"uniquePinIdString":"8","positionMil":"310.78504,947.22748","isAnchorPin":false,"label":"VCC +5V"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Loncont LSA-H3P50YB","category":["User Defined"],"id":"698fdeba-91ca-4b68-9d55-5545583fbf52","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"c750f18a-9432-41e6-a6ed-179e28bc29f6.png","iconPic":"3f9b3f3f-db41-4a6d-b13c-7e86a7741a7b.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"40.94488","numDisplayRows":"29.13386","pins":[{"uniquePinIdString":"0","positionMil":"1267.23504,2577.75748","isAnchorPin":true,"label":"L"},{"uniquePinIdString":"1","positionMil":"2788.58425,2622.59094","isAnchorPin":false,"label":"N"},{"uniquePinIdString":"2","positionMil":"1276.20157,339.07244","isAnchorPin":false,"label":"LOAD"},{"uniquePinIdString":"3","positionMil":"313.77638,1325.40906","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"4","positionMil":"303.79882,1534.63189","isAnchorPin":false,"label":"VCC 0-10V"},{"uniquePinIdString":"5","positionMil":"313.77504,1132.53748","isAnchorPin":false,"label":"VCC 0-5V"},{"uniquePinIdString":"6","positionMil":"307.79504,1927.58748","isAnchorPin":false,"label":"PWM"},{"uniquePinIdString":"7","positionMil":"313.77504,1730.31748","isAnchorPin":false,"label":"VCC 4-20mA"},{"uniquePinIdString":"8","positionMil":"310.78504,947.22748","isAnchorPin":false,"label":"VCC +5V"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"DFRobot DFR1073 GP8413 0-5V/10V 15-bit","category":["User Defined"],"id":"7b6ceb33-1206-44c4-8e9b-79797c6b533a","componentVersion":3,"userDefined":true,"subtypeDescription":"","subtypePic":"28139415-969f-45d3-9930-3634e76076d7.png","iconPic":"edf2d60f-7dc2-4972-a04c-2a93629ecddc.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"13.77953","numDisplayRows":"12.59843","pins":[{"uniquePinIdString":"0","positionMil":"158.31260,612.21535","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"152.33260,411.95535","isAnchorPin":false,"label":"VCC0 0-5V/10V"},{"uniquePinIdString":"2","positionMil":"146.33260,809.48535","isAnchorPin":false,"label":"VCC1 0-5V/10V"},{"uniquePinIdString":"3","positionMil":"1356.86102,743.72717","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"4","positionMil":"1356.25394,662.97992","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"5","positionMil":"1356.25394,585.26850","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"6","positionMil":"1359.24291,507.55748","isAnchorPin":false,"label":"SDA"}],"pinType":"wired"},"properties":[]}]}PK
     #{dZ               images/PK
     #{dZ�&�y`  y`  /   images/8c2f1315-cf23-4ba8-a920-becb97f13280.png�PNG

   IHDR  �  �   ��ߊ  NiCCPicc  (�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D�0գ ����d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c�%��V��h���ʢ��G`(�*x�%��(�30����s 8,�� Ě�30������n���~��@�\;b��'v$%�����)-����r�H�@=��i�F`yF'�{��Vc``����w�������w1P��y !e��?C    cHRM  z&  ��  �   ��  u0  �`  :�  p��Q<   bKGD      �C�   	pHYs  %  %IR$�   tIME�WxG  �zTXtRaw profile type icc  8��S[n�0��)z^�8~$R��b;^eWݪ��HQb�0$|�>�� D�h`�dZ@�&F�Ąb�9��m��P=Eec������O8��`��Й�f�
�Q�A:���{�xt�k��7�����������-eP/���\!�����jS�u�mۃ��Qa;��B�["�,FدCl֤�	�����/�&�S�T�c��\���~�y�_���D6:J&�D�z����f5u�R�����Ye:�010�����?1:9�����{��5nH����^υZ�w�R��WU(5G�Ӫu2j�fo�-���)�:&c*+q�y&�"J��G��|/��d�c?&s&]����VG��^q���@����줁/0�   orNTϢw�  [5IDATx���w|e���3[�����!�XQ�	6�g׻��;�ӟ�SO�]�Slxީ��)6Գ��^C��m7����cӳ��؅|ޯ����y����S�y """"""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""�P �t뎇yX��s*�+��������L����>����<�r�ݵ/�ϯj>��ߌ�	�\51�;Z�w�e[�L�>��( ��R�	�NUo��W{��v��	댍
�_�f�|����Io[����7�9	s� W�>����&A����@��H��t@U���"^ n@U���^}z/[�j�[�*)9����n͚?VTV����� �*�, 4 ��{!��yLDDtX2�I�+�|���5]�dݸy����S�NMX�˯����^!"Z�SNDDDው�]8|�+LUU�S�
�n�u=&҉"""�����]bc�L������H'����ZND��fK�<�M��DDD p�ݚf���*(w��CDDD��%�$ϷX��'0���������p��a���ʓ<���#������	E��Qn������iӶ/[�lBaaAV�`�Դ48��vX�6�-fh�	�R�4J)(�L�O""":t��r�];���T�r:��'O�����z��:<7<O�����F�ۍ��*����v����"�_A��jf"��r�|��������Z�����=v�m����X5z4LZx�Ͱ�����QCrTAii)~[�+¹1k���e�E���;���^�&���� ""��:Z،m�tV��r�}^_��✕Nx�^�m�H�Q�6�5�_�6���At�z�^{�7].��#�WDDD������[u�ޤ�r9�q{"�F"""j����"b�-��t:]p{8�Q��JJK��x��.��o�\.x<,�E9�

�i*^=x@w��NDD��VPX �������}U�z<p�\�N'5C++)���r��~S�7}>*++#�F"""j� n��&"M����|��`@'""�f
�����D����>�,�E5AM	��������r��t:���(4��r� Ȉx>�N�3҉$""�������3ƌm��.�x��N%�������/ �y9�9Q���M������NDD�4 PJٍ�������(��@([�6t �z}0z������h 4��^�����(�i�ee����h�����(�iK�-W*D@�1�E=m����R�b� �Љ�����_�� t�"A��#""����+ �ϡ�ʝ��(�VZV��H�*w/D�H'����B�*�˕@LFx}>��NDD��VQY�D�Y�NDD����
��q@���;Q��*]N��!��%t�t""�h%М��J�u�h_u�8>�FDD��9�����_g/w""�h�UU���S�����G:�DDDdD��j5���~?K�DDDQK ��p�tݯCg�;Q4�b��b�W]t�)���(�i�����]��:QT�L���]ס�|
���(�i��LP�0��܉������2�fJ�r'""�j�)(���ua�;Q��bR
!:�܉���� �DD���ʝ��(�iգ�i0�OM�r'""�v͖�u]X�NDD��u*��^]B��܉����V=u��-�p`""��&uݸ�΁e������h~����*w""�����z���*w""��%���u%Ͷ���NDD�4�߯A� �+�C�)���(�i�߯��ϡE9i��5v�#""�~���J`\�.�NqDDD�N��	�)NNDD��l6[�����DDDQ�l65�`@oW�3[j^���&��Q ""#f��dX�~0�d������%سgv�؅��TTT������PJ�n�!11�������dt���D��@��!"�:��i!K�pr�V��"((,Ěu��ӏ?a�����ۊ����^�'��P�Q�4M�f��EJj*�w�#�c���5j��2a�4v":�(���fM�̡2N �ro!���b�ڵ���O���o�v�Z@��hI��� �z������ck�f,��������ӦM������b6��'�#�P\Z
�łX�#��9|Ĭ�BV�C�ϡ�I��x�d�R�=�m|�ɧض5��Q��V����TT�c�o��t����o�����_���{�]-��O7���������Wa�QG��f���x�� ��ZM�mݶ/�y�y��صk'�5�촭ܚ��-�7���Ǘ�č�wfL����/ 6j���m؀_|	�����xp�e�F:i�10�\�˄� ��n|��x�����Ͽ���"�U�&-��]��ۢ_񧫯��͛q�5� 1>�A����PXT�w�{���?�r�
��Gjj:T���d�B�*w�U����r�~�<��S((؏�L�Z���jVb��d�ɤA�4�������!�/�fK!��PX���gݏ��"�|�M蔖ƠNDQ������3�������rV�u!�a���|�8������x����sꝌ0�@n�� 33]�vEnn.�v���D���#&&�*������ �6m�m�6��
?Ȫ�ବ��g�����w/:��3�Q�Q �-[���x6oڈ��/��̀�B����F�}��nǿ��:�^�O�@�edfb�ر�:u
Ǝ���,$$$�j6n�p��(..ƪի��O�����c���5&������ks�"�S:��v8�vu"�:%�%ؿ?����p�Y X�6��҉G}���u��g��Ĥd�:}:���J�1	qq��6�|o�n�!+#Y�p�	���+0g��{�-��0�{=x���w�޸䒋�)~Y�(�(@)��ۋ �D��*wv������չs1�9�s��Q�����s�>��;	qquü����e�&3��G~�>�,r��G]{c
�Ņx���p�B��u ���B��.|l����7��ByY	�s�f2a���x��p��� !>�EA܈ ���p��31���2tx��jؼi#�{�y�UTD:눈�Q  ����]�*w���������];���t9M3��s��3�>��C��K ��f]O���z]�u�qI��g��o�e)�����.��8"�����ޚ��.@m$�q�L��Y�݋�99�3� �8�d���<1P(.*�K/����Bu"�#�D�5����EX�n^|�%���^��c�!�u�,������,7i.��bL�6-d������H��!!DBv3L�ڱK����[�0��<66�˵1l�!{LL $'&��+�D��0*�������?���9�te�:��}8��)R��ys$���~P`��f����+ ;v��']��(�O�<g�uVD��;f��8��S���/5M�����? /o+���m��������z�v���z f�6�V�f��v���G��4x?����|�=p{�����X,�Z��Y�0�L����zo��v��vCD`��`�X`�Xj�o��
��p������v�����������
Ku��6���������vC=��f��6��+_�Q�ן9p����z���`2�`�Xa�Ya�X`�~\���,=F�S�3: ������]�����f�ߚydMi��7"�^@��U�_�V�Z�S+1)_r1R����& 118k�x���QR\��H.5Kh8p� V�\�n�f��}{�b��X�n6oڄ�{������j�"..�ѣ����!''16[�>����rTVV6���dBJr2̍���/,Ě5k�d�lX��w�Fee%|>lV���е[W���#F�@�~����Т������k�d��[�{���鄈��p >>9�9:|��>�{#.6���T^Q�����u��vj����dX-���+*.����d�R�[�;w�Dee%�^o���ƢKv6r��b�0` R��[�6���k׮��ŋ�n�:�ڵ�������|��CVV6C�A߾}���|iN�M� (-+�֭[�v�Z�[�۷oGA~>\UU�z�0�͈�ۑ����]����4p z�쁄��v�ٯ��BIii��RHLH�#&&h^Wy<عs'V�\�իVa˖-�?�W�~�V�������Fnn.�����#==�6/Z���N���w�Ʉ��"��_]�QPX�������M�w8HHH`MBCR�C�r�ϡ+ e��OPU�Q�|���8��qM�Q�0t�|��(�!.>���ӷ/��!C�b�ر�r�]\R�_~]�O?�?��3�mۆ��2��kf�b��%;cǎ��iSq��ǣszzuN���:^y�U��ƛ��PA�Ν�ēO�wϞJ8�v��ǟ|�w�}�V�DaaQ��P0���ԩF�9
^x!N9eb��pj��{�|��gx�w�b�
VO��SV��;w±��/��=��9�Σw�}s^x���"���D<���Z�DFM��8����s���;X�t)
��k���43R��0b�\p��6m*R���-��������罍%K��� ��x;�iiiw�Ѹ���a' 1!�uU�G[�m���_�/���e�q����\}�j��l�Թ3����S�`ҤSЭk�6��*����#f�{����T�Z����o���hpL�UU���_���a���c�8++�)�dAJr2�)S�bƌ��ۧL��>��~̞�>��chZu�Q@iI	����$)�����nGBBB���u]�̙3q���T�� 6�M3�y)���7����DDV�Z%�{��~��i��Vy⩧#�?~]�9/�,g�s������g�Ɇ�����\��{Ӷ��p:�O>���8S��S덑�Ο��T����䤓O���������9�~�����������EV�ZU�Ϊ*y���O�-���XgBb�\vŕ�a㦠i�r{��O?�'�$�Vn'5-]���u�c��V��?�4_�R�����+���RN�<Ebbb[��������s�=_��\ix.y|>���2����kU�$&%˥�_!6mn���{��ǟ��#F��jk��^w�[m12�����?�)

DD�_�jm��x�z�.���9/6ȓ�k��5��t�Y/]-���"�ǞxR��燝��W.�����_8�9���Z<^o�cġ��������W�$&&�Đaß�L����y#�+R���_��ax�euɑ��GE���n�t��oi�t���߸Q�t�%%-�A<�">1I.��R� ~@��_��[��A�dw���V��H~a��q�ݒ�֩Z�~e�&�,�W�j��""%ee���K猬�������-r��dͺu�:���w�(ej���4��O?զ��G�̬�6c%���c�ʏ���$_*�Ny��$�k�6oGi&9a�I�h�v;�}~�|�ͷ2q�d�Z�m<v�C{L��v�Y���E��5�|s޼ꛮ���ify�ŗD�����s5zL�s�m�`���9�] �6l+�=^�\z��횏W]�'��}��|������?Q������UW�)DfBN>e�E]���b�����o����
���ߖ� �9J>��3���%��^�F��W]]�d�%��N�m;vH������n�#��n~�9���d߁�KG���Y�����n�Y���z��q�v���|)���{�%	���S&O����IgU��0�E�V�V.� ��<΁�,���x}�V�Y$t@����""��[�k���u��)S��漼f�π~hzBb��'���) ���X�|E��4�5
I���3\8�o+]�	���j����h�2�>�'PJ�j��j�C�����߭²%���k����~��#L{�R
%�������˯�����뽤�>5�9�K�����|�p&�y��g�tVɳ�o磏>ċ/�����������O<�gf?ge�i�k�O_Kҫ���O=�J�n��=�O<��#(+-#���?�v���k<��l���V���³�<�[n�۷�ե�����Vs�����f��>��Ar���5����Ǜo��nǲ�O?���|vl�Z�/�Ϥ���`�5T�����<���t����ԍe�7z�����c��
�Z.ս�Us1��d^}���طo���v���T����	۟17�p#�6oBM�4���cࠁ9r��� %%�����{����e˰r�J�߿��3X�sN��my����a��q�駵S/V�߇���:�x����n>�c��ХK6z��.�]�*W�����u�VT��:F*�~/��70}�t�\�
�̞�*���vLGl<r��W�^HOOG||<\.v�؉u��a���՝Ϥ�qW������8���o{GB����x�w�rU6�?&�YY��ݻr�� !!n�شi�l1�	@M�2����8��3P\\�G~�����=Ɓ��������HLH�����]��~�z�ܱ>��4źߋyo��̙31n�Q-��χ�^~�f݇Ғ"��:�q�ӧ/F��A�!5-q��p�\(,,D^^.\�u�֡���^fԧa��������O?��G�^�+��+V��9/4� p��!;�z�쉴�t$&&����@����!o�����=�7?�}�]L�>S&�2=�z���Q��i��z�oټ~_��ٌ�}� !>�i�8�ѣG�ꎀTK <d�ˡ�ܭ�yu�kQW�|�_""��J�R�� ��]��E�qy#"�l�
>rt3U=��N��?]#��^�
���Kc~]���b��_�o7��dee7S=	�?`����/-�[�*wM�[u�w���b���㏑'gϖ�+WIqI��=��|��z���R6m�,�ϙ#Æ�Y�e2Yd��iҳw�F���O��N?S�xk�lشY�+*l���T/]&��q���t�?&�U~��v�r�+P��0_Lf��5Z|�Y�t�KU��V�\��m�����2n�1�4S��*M�Lr�Ie����|Qu�㈓I������%kׯ�����RZ^.+V��Y�= �z�}�(��|�m���Z|ο�����_�?q����k�u��r�%��'���?�DN;��z�����������q��R&INN���uHjZ'9��d������������|�t�d�Ν��G˹�/�	I�^�:�).-5L�_MP����{���={e���7ߒ��� �TIrr�����o���g�����҈_'U��_­rOHZ��C��2�[��ʫs����楗_��fx"6\v��uD午HQq��w��m<�����O?�J���bj�""UOu��)�e����8M���v��
����j����Y��n�^�{<�>Էd�r9���͗���ӷ����\)*.iv;^�O���2h�Аy3ᤓ���(�1
���%1)E���FٴeK���˺d��[��$�kwyj�3�?���|��|���d̸�C�ˈQ�e���a狈���;��ԴN��{�!���m�\�����By��g�i�V2��0��)bЛSM4�E�?a�|��gRVQ��^RV&/��buڍ:�)霑)?���;��_~)���Azjj�|���I(��VFe@4x����^y��d`mF����;���I��������W_{Mb�/�J3ɔi�ʪ�k[��""�����s����Dd�G{\���N��E(K^z�U��x������V��s�ꐡ�F�7�~>��|�駒��E�j��v�!�W�{��z]�$����O>U{�nz��Xz����Ss���ǟ��脻��� =z�6؎�������~{��*�\w��B��Kv��2�5qU��[r�麼�����|�8y�ŗZ�
��,\��?ʖ�[�F���뺼��[ҩ�q����Ly��k�9�u>~u������8�����C-�˴��T]�;ŉ�����:nt��	�6�m��{�⥗^FeE�&��0�$<���n� �z����>���f���
��}6nl�����o���a�X��p���>}zXKgfu�=��N8����:e�D�v�ü)(����[�-W �l�⪫��UW���E�2b�p�}��P���>�)�����1c���Z0@� 8��8�����PRR�6��>�ſ�ݷ߁H��i�Ĥ�~���a�Z[tk�z1)�3�8<� :gd��5E���ܹs�s׮��Li�y�L�ݤQ�^����:�L\r�%PZ�c�������QYY����tPi����,p�W����LJr2,Cf����,]�zZ������v+���ݦ�5;��~+����k׮Ň~�E('�|.��RX�ՊI�&!>>�B���p�e�a�)���ՊSN����S�*T���eK{tcǍ��W�16[���I�p�ĉHMKCs=��=�\�}��V.��a�ē���t;^��7o�?���U�|�-�޽��wM3���/�%_sn<�	�g�v���
��֠��t�̟�em�ӑ��7�x:��55�%i�Z,8��sеk�n�桰��]RM��iF�]�H������^�Fb�#��eYE>��C��A߷Xm�����;���_#G��u�]�#�.c�ߋO>����k��� .>]t�SS[�@VV�/�:�v놙3ς�ln�vrs�"-=x��u?���ۜ#5�b����.@���V��O�>�޽[�|t��s�;���k �ٳ'��2�#(..��o�͛7�/�2X�����_	GLL���V��^z	�`�tw��~�	J��ڥ��4Κ9�n�q�>}0d�P��K��Q^V����@4MӚ-��,�+ >�����餶�>o޼K/1XBG߾}q�9g7���-���N��#G���5�VW����_�~?��6�%=-�YY!�9���ѿ�6m'%9ii��RQQVI4�|�ޣ;&L8�MkINJBN׮!�3f���)�@bB:w�l�LEE�z�!�����m��tn2Yp���!77�ݚ�@�=0��i�M���8�&��֩SgL�2fMk�Ͱ �����`�[e����+���n�t́et�������v�M�h�"�ݻ���5�<q"zT�õ�ѹ3N�~�aUdYY~���v	^�G�F�N��Plv;:g�يѣG���>�ݎ��$�������|�0�aÆ!��s`�X���a���0rԨ�Y�ZC!0�_rrJ�|q���1�� 2?��#��`������ĉk�@m/&MÄ	�����7������Ö�����>�+jJ�k׮0����|>����5���DS��b��9}��d��zz�`D�6�Jm�>�-[fp�$��`ʔɭjwn�0q����%���t,Y�eeem*i��V4���`2�[=�i��JHH@�v���b� 6�a����m��3�L8hP��6[B�4����h�a�Á�i�@����.��y�73���}��r�*���>}z�)�F��h���<X��o��xڼ�A�!11��n�SRS`���	H?����%���xU��HE�{ȥ������
@iY6n�h��]�tA�~�Z�w��}���m�6��o�1z����j�����$''#�Kv۷c���tٶ2��j��w�^mi�v�a����ѭ[ז��`;m팚��{��Q�����Ў��� �d�\ߴiS�o^�2�W�ۯ1..��fXD���F��@��r�4MCL��4�i��RXX��;w�߳WO����l����ܾF���cZ;w�j�V���;����iƗ۸��fn��N��:m�v:��m�-�)���X8���(_��~õ%/�e���f�w�.��c��{�n0��ٻg/���߆���vdfd�9��X���ۤ@��TbVJi!�H��J)$��#T�����6�5�G�����W��Ē����؃�̽�d�`2Yj'f���҉��m�F|\<�����q8���9 �)�@�MHH8��c�=D3V������m[�3���Lطw��vA�� JKK���ڪPR\��6m�j�"9%�]�n6��B��v�8m��T�w��)�.���Lf�����t�x��hTPPgee��Lf3����Ih�tɂ�b����$
~���-�;b�i�bs����j|��������l�Z�'���<��~ط��MK�^�O<�8fϞ��-Q�݆�U�ۍ�¶t����G����6��A%f���n ''6�.��N���p:�H	��pQVVVݩ��~
L��z ����d[Uմ)C�u������j6[`1�@��:%��c2���RZ��mP <^o�APD�(5M����P\ܶAZ4�`��5��2�B���9�+ ddd">DUdQQ
�x'-�n�a�f2��#�Q݋�)A��m�Ř�&�ڱ�Б�d2�|�^�V^OscL ����+8]U����J)��C7k��nGm��f�~�m� ������xRTT���o�]�K�1w�*@����]v����9�`>��M碦��E�p�iLGؘ
���>x=��E�"At�vxl�:i��;�q��;���O߾�FGZ�fmTݙn����+QT\]��(Tk���_�W����Y��Pe{�T�����zЎ���@�����G��e�h~������.���?�Ƞ���ʕ+�t���=�����SO>�?���r1l�0�9@NN`2��f����_�QYQ����r��	>8��4�cbjg�"j��M���x���;�<s�O6�f2�K�.�%:�����r��G:��� �>qqq�(����+�}�h���ښ�����_�k�v�ڵ�|���t��@��}0b��u֙8jԨ&�)���i@��������"�t�������QS�z���1��!+���s_������f�s�7� $�znC���#'�+֭]��]Î۱h�t X�~=���P����ʅ���}[�[���郣F�j�ل��m6Tx=h�Ș�������������mSi�Z?8P=�Պ�x�N�U.bc�پ��&�D-��U�!���`����wW�������rE�u֯��n�w().F「�1�2220|����OMI5|F���b���}�m;vT�����l6dtj��̨c3��HO7��N���E����$�/��f[:n@ v��'MBl\��f�-X�e˗G,�
��m��駟AĨ3�`��a�ݫW�w�;�W�����P�t���ׇ���A׃����S�N=/��g�n�6S���;w�t2�ZLucu,��ƌ9
��r��$�iؽk7��{��ko��9֭]���M�7[l�x�)HLH�SSS��c<�Hޖ-(*j�`F�Ôb��͆�$%%��8�D�޽z�f��������o���\�լ1��҉�&��Ն�1�_��.]0i�$(ͨ׫�?��.\tȿ�
���7�xOU]���G�8���1!!}g�Rؽk76���v۶m���[`ti�ѣRSSbNRGҳW/���� ��%%%��}�Y_޶mX�b�nۆ��b������ܩMj&
���a�4�}�L������ְs�v<��c؟�Ⱦ�
�����9/b�0�7�0u�T���ǰm�j6c��Q�XlA�TTT�/�����m��W_c�޽~:j>b���ٶH�{�n�e8߹���k�j��v�n�Tŷ�z�N��3N�g���/�7��x��G�漷QTT��N-"�hh�U�w�*w0h�@�y֙P���_|�^xa\n�!�2~��Wx��W��U������9g�k3�{�1�32��E�W_}��۶��) �������/t�}���aԨ����$
� HMI��1c�&X�����7o�m�/���|�}{�`������x��yx��'q��7�GCE���!Ҵc�:v��b"�Й���z���O���SO>��^zn���u���q���`�>��- e�̙ga��ͮ�o�>}�h�w5l\���|�8� ���ϰl�2�}���aÆ�ܤ�Ƥi8�	HI1�Y�g�~�%K����X��t����7
���!��W`KcƎAff��L&4��XE�9�zˉ&�t�:�s�u�(�_����fw x9�������栢��u��E���K/��=�����/���)^@B\�O�{L�q�=�*<������e����Vᩧ�Fee��{�2aڴi���>�/pth�5
�F�B���a�x��Ǳw��6������W_ᓏ?6\2>!	'Nl�6�H��Ï��5d��i�pJ�S �Ʉ�.��N��C��� ?���|˭؜��n]m�n���G��O�`ѯ��X� 6.��_0hР���ĉ'W_��ض5�� �mk�>) ���C=�իV!xէ��ݻaƌ�T��UM��y�Gl�:�}��'x�٨t�~������u������� F�Q����C�{q$�ڬ0�-���'����9�L��@zj*n����ۯ?�= �P^V���'.��b�2�5�;�ߪ�^���<�}�?p�����K~�6�L8��p޹���, ���p饗��Y澜?7�p#6l�ܪ���k��r�mx��wO0�ɂ/�C�a��iӦ�㏇ѹ��z�ܳ����BQ+{�+z��q�X��Q�UABb2.��rtJK��{�#6[�!x<-Z���΁-��7�_¶�z�����u'2�d�8�+躎_�	�^s-.�݅x~΋X�n=���-�����+1��q��s��#�"����8�N��[n����P�8�t̘1��}]��>�5�_/X �����Ѷj������E���ÿ_��M����
Ǝ�+.�V���$ux�SZ���/��2�.+����ч�M7݌�k�A�0�58�u]���~ß��>��Ð���S&c�ē#�-�L\|b�1�
�}�̛7e�+~]���g���>_�8?3�M)�}��pV:q�m�#��>�zd��t⛯��?���ݻ㨣�°�Cѯ_dee������NTVVb��}X�b%�/[��K�b��mգ�5׏Q0v�8<���գG��� HIN7ހ�k�b�eA�MAD��W_a��u8��p�93�۷/����҉-y[�чa�k�a떼�u5��[�����н{�QZ�șp≸��k0��Y�r9���T��rᕗ_������/�ӦMC�n]g0\���
y[����c�ܹؼqS��<t����IhR������aÆ`�*�ٳ��z����0` ���PU�B~~�?����Zx�_C 1�|�fo6}>�9��!��_|�Ep{<���b��=]j���x�i�zlڸo�a���@bR�6t�\.8�NT�������P�a��`�1������#Z}����1�Y����my0z�g��]x��G��o`���}�hdee!55&MCaQ��ۇ�K�b���عc'�~o�}ё��	����4q�8�ԁ	 �ł���
�v��K/�T�hӠ.��5�W��nǜ9s0|�p�1�3����Ʉ��r�ܹ+W��o�-�֭���y�|�;�#G�0�Y��=z��g�T���G���>� Ji���ǟp".���%%u�<�����}3j�\���
t��	��+VT�*�_l]�QQQ���2��j*��i�-VL;�T�{�=<p`���S�L���p�-�`[�u���;�g�N|�駰X,�X-PJ�������DGVv�����.�I��e��N �$%���^��z�MA�^/�lڈ-�6��wޅ�j��b�����v�ü��93w�uN�1#�W&ҙq��l;v,�5>�a�� O[ri��(,,DrRR�w#z����yUs����eO� j��̳��+�����<�����	��^��=	w������sϴ[0 M�0s�Y�={6F��y>�h�u.��ge%*+*��x�*ԅ-��!C��SO��/�����ړ �����܇��+���{\s><n*+*QYQ��*Wu�i�|��={��G��W\���!��I�N��aC�5 
�����H'?�h��;����Ç���O>�����b�"p��|\�q�2�T���+���;�����[Ӕ©S���W_��.��	�a�W��*���HLJ�e�_��_g�y&,&Z��[�P�+�j:��}�]x��'0t�(MC�`��@5�K�|���<�T�y�E��y��ͭ;އ��.L�s󭷠KvW�$�WTT`ǎ�ޅhn:zs@��4�����)���{������5kQ\T���Z�խ���̒�����1c������ɓjs9XGH <�<3�'O�+���E�����%ψ��GRr
�=�X\tх�4i��ڶ�n<�t�i��� ����4���vj�_�01�N��K]�������X�����¬�z��rI��o�V@lL.��b�;��}|��6o����=?Z�y��5�����_r1.��|dt�Ԧ�]D�=��ů��~=	<�l{��ߪ���f̀���+W���>_+ۨ�ra˖�����ݙux]g@oV�i�='���:\x��X�r%���{���ö��P\T��e0�w0
���I�ջƍ;�L:�F�DjJ2���
s�p��c�ē��w���>ǢE�k�.8t�N�̈��C�^�0��q�2e
�9f<��{���S
�9�2tX�1�u���ܾ0�ZYj����l2��HW�_G��}`j�H_�@�G��1x�Ph����޽{u	�y�6|x�s]ב��[��v���:lx��뺎~���j��b��(���9��_�ѫWO�Z]�S�f@n.f��\x���������`��U(�/���Fs%Jbbc��)Ç����N�	'��ݻäT����d6UUU. "���T8z�V||���Ғ��/8b㐐�ت�6�L�y֙0` ޚ����%��塬��6�( J�`�48bc�������sЩ:�2��w�ݳ;+��_r)^x�y�m6��@M��"(,,Į]��c�l޼�7oF~~>�N'\�@�v��M�`�ِ��Դ4dgg#77����ӻR��`�>�#u,j����Ǝ;�n�:�^�[�n���P^V��
����@\\,233�77���b�����̄�:��~�ʊ
8�Π�[,$&%Ak�ޝ��p��o�j�"!!�p���G���vv����\�W�t���"�{f�III��p�Dee%*&1�-HJJl�픗���r}/��I+_�Q����Rlٲ�ׯ�ڵ�k׮�w��n���!6.q��HLLD�޽1`�@���=�wG|\��;߫�n����=�4�II�߱���xQVVt\�a����M!P�p�@>��m�Ν�p����N@)���!11	����YY����n{}D�_�7<�ԓh�&4&&f����ڳo���P���]��^z1v;z+��]A���x<�z��z���|��|Д����
{LlVk��F��g���������J�l6�b�"�no�6~����/w{m�p����hَ�6u ^�.�^�70��R�X,�Z��Z�������<8X�>(��ߏd-�fa�! ��o�4���p���~���9�4>#�&���b�u����3�Ѳ�m* V�VKBȠ}0��<8�ېF?��z���ЯlCoo��k?�N^�)ԑ�|?��kᡦ��|	��:Q4-�����p�""��$ 4�ërg	���(J�Hӧ2�E9	���e�8""�(&�.͏3�6t""�������Q4-�����:�E�:�5_B�u�����(-�)�D�˝���;���0¿�h�DDD�>�.��V��0�E%DCm�::QTif��z2�E-�$�6tv�#""�Zv/wщ���VJ��DDDQIDD����Љ����ha������(���;#:Q4����3�E)��{�����(j�7�+{�E��&g�s�DDD�K­rg	���(��`�5��E��̶�Q0"��Љ��� ����ֈ���Z�Я�U���;Q��yl��`�XNDD�D��|l���(���Y�NDD�D���NDDtؓ�Oe('""�ja��V�E�0��Y�NDD���ǡ_����[���8�+Q���H�����Ba�;��#�8Rё ���,�E�p��YB'""�b��rg	����c,�j-X�����Vؽ�Չ���V���Y�NDD�X�NDDt`Fu""��ő∈���2s""�(��ʝ����NqDDD�?ζFDDt�p,w""�#B�m��DDD�,��eX�NDD�Z0�E+�GDDt��ќ��(J���;�Љ���Xx%t�r""��֒��։���T�c�3�E%�!"":"�߆.�r'""�V�V�3�E��*�棵��E��c��Z�)�����Yx%t�C'""�R�oF��Z5�ADDD�R-��>s8K�u���()-�����C�D:J!���h]ס (��4�]���������*�]�+@s�	���jE������U�HD�Q�y����>x<(M�b��d6!PFm�밴�����ػ{ws�U���J ��W�1J�DDD�C!�[�* W�߆v�'""�B���Eo""�Ù���G:%DDD�j���tJ�����t@y5�ie�N	�� ���v��H�����ZGӴ����2-%%�q�Ų������#�aK)����φ��F@Ff�q���wy<�" ���j�U�{N�p0:�%@��iͶ�����pD�g?��������9ETM)��R�V��}gm\�a�:����F�~�w��ի��2"V f��b���1&�ɪ�4��4��4�R�T��`B৪��R5WE�T��k�U�f�.�PX�v����RhxW����x9.����R�<\(T�]�R��ԀR����u�V���o5�k���^�=�:Z���Y�~Ԧ���������j��d}J��u�������4��Z��p�	��ʂޠ��^��u��c�o�5��b�x��/=��WD�H�����9��:{�~���������nHBi�{ͪ��R�4����k?���F��w���'��f�!��`geI��5�|M^�~�������4�	��t�cP��V�p��Vw\��n�f�'�z}���`����~i�'|�P������e��e��FK׻�68�W� ۯ9$���dݵ��p����u?t����������K�Y_��]�j�GR/���\�dX �5ikt\��*e�R�p��I�ɋz���ͯ?��ڹ};�~x�W��]��E��O�����FGT},�4��o
 �t]����߯ ݯ+]~�_��D �_W��t%"�~��s��oP՗]��^W�i� ՜ "�7H"XMŊ��>���]���>k��כ����}{��m�9��g���_y�7���4������]�78�J)���x���q�I'��^O���_��5oIݽj��O ��V��b��Ҡ���"5�RR�����R��$5W��;_���U_���BW_]�҅�r��ȁ?���M��r��7�R����d����/U�=}��Li��i
J��MдڿiJA�(/nKE�c}+M� Д��Ai�mk�Mi  ���;�ݨ�j�,��Q{JNIE~�<�쫇q1� ��)[�fʼ^�}>8u14��4��~�AY4(� ~?4ѠC�I5z�_�h�P ���\����k�R
���5��=�j���5�^[k�ª��5�)S��/uWߠ�cG��ɧLz������-���+��s�|6��0٘PRZ��n�/��r�������#F�87--}魷��ߏ�1���d�l����&��-W�ƥd�hT�Qu�T����7��n+�ꭣ�i�h=5�u ́�Oլ\I��������R��ڂQuU��K����[����_�D�N�	�ʹ�p`E���Hmy]�4����P��nOS
�i]��L�u@��lF �X`����*������t�	�v#..J)j|����Kv6X/�y	&�����D|B��v�G�7p9�� Æ��m;v���."�Ꟈ�����?"1�Xi����*���?�㳟�[��E�05�ک���L8�$�������M�Pغu֮] Hk�a꣏?�?���`��������'���Y看��6�sύtr����w��w��[o뒙���a���Lr�=�8"J�""�,\$	tMh��q�ۏ=q¸�YY�>,DD�XB��23�0c�i11��A?.\��Ҳút� l۱w�u֬^��_	������~�o����[o�S�<�$ŀNA���`��1n�ñ�d2]f͚�ض}[���j
@IY|�!|��Wh�p�RSS�>��c^�~��k�N\w�5�N6Q����[t꜉�cƞc�����ݭ�ye��ڎq������#�=.��xi��O�ظ���=�8�#.҇���Y,�SP����٫���7[,֢`�x�.��˯p{�	�>��3<��cpV��q��d6{323������7�Ήtr��Bb@���:�����:u�e�Z����l�2���V��
��U�qｳ�o�n4�(�����G5�I���6nğ��C��MDD�:�>����k猬7��t����N���?6��""���Η���ILL���#G���8"}���ڮ� ��={�]��A���d�'��}��*�G�w��l1A��M&�;;��"���.�sϽ�>DDaa�;��q���d6W[���b��%�r��j�O?��>�,�n����aC_7�Xٳg���H'��(,�d���>Đ��Щs�-��Ш}���8����T�n~߬�p`�^;��11�srr������G�?yB��MDD�>f�s..�������_�UQJRR���oDm���ȁ����f��٭[ϫ����/��F�����EXB��F�����,��>0�}c
%%%X�|y��j�������G|�}�)$%'�w������S&cǎ���D:�DDD�G����?`Ѝ&�E^�����rE])]D��>�N�A�i4��KX5���t���&"":8���[d�tØqGO���F}��a�u���	���`�|�J>r�a0�X�e}r�] ��}���NpDDt�:u��8�̳�&$&m1z=)9U��u������!�͕f����go����s��_o�!�YMD�jlC�f%�$#77woLL���K(���bٲe�Njuj �׋�_��?�F���0��~�j���x��"�t""���G���={?��I����9�|�p:#^Jy��s�vs��Q0hȰ �~c,X�l&"":�j:�6��f��g�"[�n�h@�����#Gs��������w?��r���]wϊt|_|���O�p��Wh�<zbb������v��ϛ����u�ge�?�x�4qR������й�Kq�Eg''��
�5Q�$�=�`Ăys���8�v�=�x(3���"�Ý9�	��CRb"����6
���˖.���D�ÁC*?��x���vW!�8�f�ٓ�����E��p�ݳP�*�R���DD�c/w
Kf�,\q٥����U�f|ڬ]���8�iS V�]������A�`��BrJ��G;��S�L����x��q.E�� �KF�;�j����GOLJ���y���ED
���/(�v󸸄���3<�s& ��>�t�z_|�N�p��:}P|B��P��<��#�$���x�^y��G�k�nn������� j6Q#�#��),�'O�裎����8�-'�K�.���:$����xꩧQ�D��vMӐ����i�Ϙw���`���8��#��DDD�ܜ� "Z�^}�`f�a������^3N���e���>o�IbRʢ�&��k��!����,$":hXB����J���V��f=�R
�v�Ė͛Z:4 %eex��G��/���4���]�u���W_nY�|n��o��B""���>j,N�xʉ�ظ�6kM3�#�=~�J�^�_�|z�8b���M&��[���������\�;�~O������s����GϞ���o����묬L��^ݎB��ޮϣ+ �}�=�x�	8+��txD��Qc�z殿�����>�L�����(z<�������]�u��xxUȰ�#dێ�ZJ�ۺUN8�$�vsh��m��㏱�c  o��v�����(��߸ 0pА�4�,Fϣ����7�k��."RVQ!�\�g1ޮ&��շ_������{���#�eDD�;�Q��ر		IHNN^n�Z���R(--��+�m�~��ƛ�׿^����oUӐ�)��S&M�{�Y3e�M����t�E��3N�̳�����ۨS ��K�UU��R���?�$��䆬jOLJYq�)����,"":�XB���������p�n�ܚ�kPPXئm) ;w��}�fa�0|D�n/�޽�_9͇}�����HgQt{� "澹�_2`FIZz'��ZUB�W��t����ILf�a�\3Y�n�{>�ҫsmW��Z<=��HgQ��UU �3�:�ŦZ��*��}��U�~y��Krr�W�k�����3g��3���0y�4�qNDD����
#G�i�Θ�P���+/UO�K�""�M�����=c�>�d �DDD-u�5��ڿ\ףS�����Qc�ɞ���.�׌Ӿg�>�q�!K��͓�o�-"��v�x���"�-DD�Nq�*��;��O��!�U۾}�n��z�*��>�>����S
��>�0�9g�9S߱s'�v�u��""���[�[3���&�%T)Z��R����󎤥wY:OLJ�8q�Q�9�  �/�t�~D=z���i��pĹC{՟�������V����G�l7����G��= |2�K����HgQ�qrj�-[�`��G#..n���(v:+;U��^���%蜞f8Q��_X��+�-�Qk��i�ҥ�[����7F��5�V�9-*Q�=��l�~{���[��qY]rdђ%!����̺���cBV�wꜱ����;�����@���������7ބ��G�>�ߡ&j��b���n�ED>������jW���P|܉���7��>�t����{ ��S��d�;ĸ]�u��M�>_�`�f�:9j̸����M<t�c?.��z�?f��g8�9Q��vƙ��UW����^���ēN�����t�������J偗R&�ֽ���xc��睏��^�]'"":r�����Y���G��ޣ׶P=�kwY�|E�������ǟ�G\�vs%)�i�Κy�$ p�uk�ϵQ��v~[�,��1�~0�r��~�?�Ou����_~%9]���jWb���{�	w��魷����|�]&"":򔔕AD���N�b��hG�t��]���{ٴe�{�	!{�k&�<􋧞y���7܈y$һKDDtd��変�\i��xC��%3N?CV�['��j1�X6;���k�������W����G��Y����}��l��\@��8d����h��<!1�s����$"�_~����#��DDDG�5k� �Sgddgǚ��OB�������Ymr�	'~4��S�}�y�:�_��M""�#ߥ� ���z�����u�׀���=����:�\ �眈��8q�46�;>#>!��s%�]���DD��nl޶-һGDD�q|�� ���g���[��f�L�>��=���~��7X�zu�w����c���7��~������̬�ו2�8��cbw�vƙ�fv���v""�����G{܈ظ��-
�J�9b���õ֦�:>�/һBDD�1=?w.�="��=z]g2[��	��"i靾0hp����b��a��""��������N8��8-)!1�悹R&;n�޻��Ǥc�;"ªv""�H[�`  ����{7[�뫫ԃt�-��w]|��h�N'�{��H���o��S�L �쎋�L%]w8�^�<uZ����GT:��N:���@$%�"%5�j����i�FU��j?5�Sv�,t��k6l�t�����1�dA�Ι8pprFf������Ė����LIM�ӳOߞv� p��wG:�DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDG���Nþ�C   xeXIfMM *                  J       R(       �i       Z       �      �    �      o�           ����   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��    IEND�B`�PK
     #{dZ�����  �  /   images/6fc4b800-efc3-4a5d-827d-9566cfd108b3.png�PNG

   IHDR   d   d   p�T   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  cIDATx��]	xLW~��d�(%�J"��}�%(�Z���B��_[y~R�R[u�E[[����J����ҿZ��j��B)��'s��;��Ĉ����>���=��s�s��-�37:�PTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��AW÷&��z\I���7�)I*�Ev�Z�:d;iJ�3mtRɲ�������V�$IY6��"a[�d��$}/����~�l���99��t.��$u0Z��d�M��(��5D��a�}0�*�
��?���h��dY~�`ȫq+��L��yY���@���[���������ƍ����0��`�Aк�C��"�|<B&�������r����t�PQ:�;w'N�{˧����a)y���3�t>���ʂ
E@fB\yyP� �f�3b�1�(p�3!�<ÃY=��䫄(�d���?0��&1A3vH�JIi�	�YCd��c,�p?��0���g�Ж���lqtws���%b�G��ɒ�2d'jaxR�v�Zl߈s��S�����_C���2Js;�i���8�f�ɒM>�Q.]�����С�x�g/�5J<����зO̚=�g����f6.:6lX�t]������B��5�D��;ѽ[7���s�p�0g�,�n�=_x��(���E��~/���u{���F�m�6�2�h��!����v����;����dX�i5�7�}�����ٿ�2~޳?��#n������1p�@xV�$��u˖�Ѳe��H�zi��|��u��,�Ν'�����ԩ3�/�5PP��7o���,�_���C�޽ѵK���ǚ5k�t�:>�,^|q 4�XȺ����7!&&�+{�_�~��d��ǎ	SԥkW�o؀������A��n��B�p2�7n����Na��>$3��ARLN�G��&����~�� �����QQ��wq�������Тe+xU�ºu_ lQ������͐�լ�K�.����ԙK�.��9����(�QN4|���X�p&M|�����5�OLLDu��x�"�.Y�9o��&�l7ww7�b�rD�c�)��?��޽E��jO����[���a�0�?B��ۿr6n����o�Y�}��E�E�:uh@lAZZ*�i`5]�ر�u�9Ǻ��<s�4�V���ի۽��1�Q�n�:AƢ����D�?O�F�g:b����a� i4puuÑ�#������W��u� ̜�iL8^<H�Ȏ��ʕ+Bui������®�v�u�zS����u>l�ФΝ�P�U�@.��+��������^M�5c�L�L��S��nW",�Y��e��'""#�|���'B�B�FMТœ8���	�R��ӓC��w��t�b�_G�R׿ƛG߭~=L�6U��?���קў��ݻ[��Z���\�rLd0�q�	��o@Ey.D<kI��
2^U��~�zB�!C^65V�E�6m�W���$!-^�j� ��溃��������͂�٤������m׮j׮����{��l"��e����G�fg�AQ�%{ΫbM�6��F�흚6m"�.\@�ƍD���]P��	��g�ΕG���e?h�V��\��ӊ�����ٳq"m���`1i.�[8c:fd��Y����<P��6���׻�2�sq�{dDG2kd'j	h�͛��)2;U�jW��%�=z|j���)�b~b����!JcӁ�L��+$3�i��ߪ[�Fc�8����2�F����~~���dG��?��%\�9���ɡ���3lw[wGDD���Ç�6�V�Z8AQ?��6U_"���YԢq�0��$��_M�i������W[P��@�nns+�F*Z��@'����!����ǤI��`�<a�CI�>��p������<*T�[�Cɩ�1K�,>�>}�/�h�M�vhD�*��89�-�aq�֭�M0m�t�jQt������5k?C��M�ۻ�Mk5���Z�e����ZSVY'�����L���������'����F����g(4�Ŷ��P�^G�>|<(��p������_�R�VUDK</`9rr��WhI�6��E^��9��~��΁�ʧ(��K�c��K�^���}Ѭis<���b�s���J�efp �e
���,���5��<�5o۶oD��h���%.�sab��F��%a�ȑ4I܍��u�Ȗ-�!00�==̤?�9@���������A��"���K�T����J��2
�������r�̋h���C�Шn+���\�t	�i~`�'t�dA�����Ӄ|�'���GEDCQ��z�5{zP�gA`�@��?�h����\�h*��5���]�r^^^pbb(��1��[ޒbo�ػ^8�s4�叽|�4�@����4}�#0(h�my
?A�#����Mg�<��7��?�il���_ �2Eto�����"����j�37-N^��4g��)�8����&��'�*JBCLQ�JH�C���=d��,���}X5D�2`�����0��g窆(&Q#,���!�.o���e�TF��[���9ʲIQ�[�<l�M�V��|/="D�xOR���vG�_G�3˚��7��aj�gE��s�6��ˋk�Q'I����܊�GBEiB���j���QCG�h4Z�D�$ݢY�-R��By%�V+i�T���I|3����4����ĉؙ}���2r����)���Om�fk\]�zH�|�R�iO�l�Mۗ�I6_dْϜf4G��Fk-匷�ݥe�k�\𛍶���V���_�3���X:�-�b(ڴ#ݾ���KĤ����h$�v!VI~}��+s�^����xg��p�h4"�E@�Ӈ$^N������1���	�����ǁ=j��������o��qbZW�?��i�1��wI�t�G��v��e��^3�x޹���k+�t�w��`-;q<3��rJ�r�##���Κr$55G��޶;�a�±c_�ٿΜ�V�{J9�Ԕd��=�(B���}�\�.1�7����׭w�^v�.\�[��"{x<����̣������{�"o���]�|ҵ�"#��[v��n�ٻoޚ>�Mۢ�̛;[�A���(Ks�#�����@�V�s��I������׸��������gn�fV��8\��@�*e	%F��#�n�����8v� �2�Ǎƙ3�2+yV{<6���ܜ����#d9�¡��ȏ ""�z�ז-_�M���^nzjJ�QNk��i�܇��#��~_�Z(_��?���&��2�G9��ɡ�=�gge|�yx�fY$�Q�/R~�'������ll���<����� ~�N�z�����t
s�PVQ��<^�q�s��mOrrJ@�=�t-���K		粲24x6�;�;�%JHJJ
*�|D��-KKMN!p5�olI�x��ݺ�Ge�F��kǏ�H�"A�ռ!i\�xzz�/_�<�R�u�7�u�����U�F��K0��N�rx����̬L�(B���^b���x:y9��}���E������k��%u����QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB����Blg���    IEND�B`�PK
     #{dZ�?���� �� /   images/ae82c023-d9d4-4942-aa8d-ab2ae3c53d73.png�PNG

   IHDR  �  �   ��ߊ   	pHYs  �  ��+  ��IDATx��w�$�u�2�|����n�����`a���!R�/��D]('��E�#���H(�(�D��5�`�ߝ�ٙٱ;����._���~/�U}�S(n0���hTU���2�&ϿYXXXXXX�7K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�}��/��l�v���O���A��'tB�\
(p�s�?{��N�p��z����@^��MA��1V��'���My�Y�����8��j��<&�㺉u����~ �`�tڥf3h���)�3tpX#���V�w�������y�`��%z߃ �j�T��kwe�A��styN|����݉�v���!֕J��h=������8�t:�}��y�`����{גc3���k���ͦ?P�Q(l9�N|�3�Xv��X�~�-�}�{ΐ�E���E_����ݯ�����L&��t6��[�W&c~�w�V���D,��K`	��0ީ�`;����@D �@��}����4�a��Q��@������d|�}�����u�=� yb��~�s������aǇ�}�}+�����t�{�;����W!~ܿ���qpp_!�x t�έ����ƣ{�q���sC0��N���{���sXB��+�ر�Ɋ�d�<�ө�<�O�*Vb�n��~�6��e"�|����@�J 1�vz6��y��#�o6�r>ޛD�����3���c�$��'ק��g=G�S	V�ѱ�Y�b�W��y��Γ�\�:�o�X#@��z��Žp�b�ɤ�5����Ϲl�Z<��G��\3)sV���$�� ��-�
۶mss����~
���8�V�D�z��w�9"���k��MM�$Js?�h4ۄ����B@����u�sd����.��&	]I_5^S 0��q8W��4�� :6��V��"n7�ɴ�)D��FLa��_I�������&�
)�c�vR�͑�X�h�B��T��5�Mx/�8�v�i��󱞬ݡ�\�	�,�S%�� ��-�
o��&�C�Z~D 6�/^�ط�ti�
%'�����$��J�&���l}��0�S24�V��x�]M��yH�O�7�I�:o���ti�IWaC��s�u�e�Qo��Ѽ��~y��uB���x���������1��e�^�S��w͇���-���
`	ݢ�0::�� (���5&8'6�2)D�Y���T��ik���8��k��X��0R��빬����Jrј�:������.~r����y}��>GHԧ��.Z~�!�B7�ϸ�k��&m��)/Zy�Ga��FkRb��I�X��E�r:�mh�B�L�<kL�:��̕����͠i���\�.���{��~���O��*x��L$XP(|��K��q�8�¢�a	ݢ� �j~�תն&R�g��uM���2��d���$}��qj6WM�Ԣ�sA�
S�U7�� 9=�Ԅ��;����K��浘~�fm�aj��8�$t 1x�d�ڴ�Ztz�i����{�{���W׉�ˉ�A���,,�XB��;d�������֌L�Jp�*��	�U4T~��(�XaM��EJ�I0��P�1��Z:2��%I��.C�j���h̖ߠk�A�̱��륅����J��@1���A XZ�5N;b>����&�V	0�~fO�Ұ��}�y��DZp&��{��V�ږ���=���Ծ���N��!��y�S�U����hPL�_GZ���B��e����5����3l�w���ϸ>.+���{��إ����4�[�⪀%t�>D(>r<�W�Ҏ�:��_I�Lj��|o�=y��y�ڮ�2f�EAgݩe��=�6��z�fZ2*���͠>SCO�����ܷR$��ϜS}牴�����c����T"�s�t�Nxdaq��E_a������6a�@�I"6�I�W:�~6��z�%�L�O�e��㨙�\�I��y�L庆�~]�����AS�1�ｮ�m�0R�z]���M�n&R��cZ5�u&3�׫�0�\�a�O:��>�%t����ÇQ4�5I�$�K��K�{�ٮ���ģ�lS36���)p I2�yH^��kF�����^�WMZ5x �O�y����f,A�8S0��G��Ma���k�)0�����j�W,�[�6n�2�0I�!*�I-7i�N�}����2כ&m3�m���fn7䒚t�s��z�4/i��
o�z�� �^�	S��%8�{s���	�1�L���b���2���=d!8N�}
K�}�R�BwL�Wp��!��րI���f
S�6�Q(�h���'��L�:�J&~��^�JHj�J��y�cA���$f���L�ݯs'�G���b��'�!zY:�L'f%e���*�%t��B>�g2ܤ��4���\B��gi����ܟԐMa!�}��'�H��)D��s暓dk�g�Ԏ�yMS}/S�y��l�mf0[����^�Y^5sL�\� %�@���[���K�}30ʉ5P� "߬���E�� �K��Tq3�p%�{R�OoF����ڬ�)�����f~��vS�W�5�0�#)�$�����:�Y�=�i�=�c�����h4$}O��g3'�g�Vp�Xha�ϰ�nяp�����iJǫ?A�P�ВZ�I\fڕ�J�G�HS�S�2���L��s�(�����d�m����fJ�kZ)�H�~}ՊU�u�)�hs���rYۦ�z��I���k��ΡתB��-�ߝ�>�Z��/�z[�/��u�����E?"lkn+�]ajW�XI�dPC�7��^ڥ�&�v�wl�ӕ�A@͘�L�9v2 .�='���O��z��n�=�\�i�WB6]�
�Z�k5����}��5��Ke�sGd߹�����b���XB��Ctjw'	3������g��+O�i���/IȪu+)���{	���oc�isIj�*�$��^s{w�P4h��(y�\K�{��Wб�?s,�C�Y���oaq5��E�!�i�A)�DD�f�K��MB�yAq�`��&��m�@B#Nj��f�c��^��伽�_�q�(v���An��k�e�0��}/��y0��o6o��<�4�;�9��UK�}�j�
2��9+H2�L2O�%M�I�wR[7�bj�J�@2�,y��ħ�oݧ�'���|���kKV�K�;H�j���n��\�`j���n���4oS�#�|�q�8�|���XX�,�[�%��\��Y���)Tz�y��8?�d�v�;ԏ�����s���\��;7��L[3Mٺ�x�3�����\}S�6�4�`��{U��1�
uZ �߼�$�'�yL���ߟ��p�;G���j�%t��C��<]j��e���� -E����׶�f���nf���d���)ᙑ�Ir6߯t=�޼�=�Ǜ�j��u��B��\�@�K�Q�]����H�O^�)����sӱ=���W��-,���-�
(,Cq�Z2.�W���"Ϥ_���m��U`0	�<i\���}f��Ntv�NT	]I����c J�f�[2�[��t\S�7���Ӽ��J�I��YF�߼��4:�ό�7��4��u�U�0���ёV�-�Ě�kX��Mw,,���-�
�����0�\�$ɋ��ME�饻�+�K�(�@Rm�ok�8?ʝ^\^�"�v�yLr+}���X��?OZL���RM�T!�R��s�V�>L�{&�Cy��a���z�?1[��?�����V��1�C|�" �Ѱ\8�hΔr��dE|�h�H��x�qw廤�^��'),ɼ��NL��r�>����֪i�2��UK�}�\.'O��/<i~�m��)Ԣ�͂+���L�I�:��0��^��Nj15V=�Ft��ڦk��t���do��u�͆ߥ�'�Vi����3mM��$������$)��i1�������RX����=��]��*`	ݢ� ������h��7i��Y����Nw������y�߂�$�D	���$�^�ufZ]�y�f�2h��E�����YtP7��7��4�'�l�>'���O�$o��H�73������X3���NW,�[����=ÚM�҂&��nՄ�c����=y�JQ��D����D���'5i3���k+A�f�l"c��z�W���U_?�^��u-����o
-�y�ޘ�R�sMa-���}�nkaq5��E_ap��e[�E��p���&LS�y���)��dzi�I�Z5P9��+�� ����k�R��f]w��nf�q�\�+խW��^C����j����˥�k�e���?�Yά��$yS�����K7�u��>�,���E_��f{��;�&�&I&	阝 3���M�p�Ji�:D�6���箔{�$N�)��J��N���Z�׹Yo=�G�g�t����7�L�[i��i�H
1fj�f�g�}[�r;��yOL���YX\��n�wH������yI��Ip�q�W-qڝW����Z��r;fh���ڹ��S�@PZ��L��p�.�����J�*0���L����'s���d��%s����o]�8'9�y�3e�����a��Rַ��CXB��K���gS�"m�&��0Ћ�ԗ��i6�˽	lS�79�,P��K�V��[��XL�5�j�}i2�MM����qfN{���v�����Z��I��n=7i�75�.�>�mz{����U�C��;�����q`��Fdpip[ˈ87����X:ik�N�фI�KK�2�w��U@�ք?佇�>㈤��=��|f����d�`���_��U�@Q�rǫ(�L�Kj�j��͸o9�S>��9_���9�g�W(⌂t� #.�T���O�V�x�>���w��kXB��+,//;�\&�n��������`1=���WҲ���^�q�c�ڭ��s���I��&י4�'�K�Sm�;���Z�j�7I�k֏7ה����BLK��;3��,W���8������/�¢`	ݢ��ʝ	$	D����I�O���Ju�M�p/B7}�&��2�'}��b z���[�%�s��W,Ar���a^W2ݭ����KV�3K�&�h�A�_޼~�;�Z	!I	�+0α�e,�XB��+d2!��4�$a�)S�����@���v�}���I����<W�LRF�դ��l�b�W�k�uӥ`oF��z�e�W2N�%y?LkC2��,V
������Z��g9���'XB��+��eX��!{��M-�$nӴ�̱z��u�����"�䚺���� f��&�^Z{b�����f��b$z�zz�]�馀b�t�T��ۮ���t���2�4��w��=^i��K�}h��j�d���1�;� /}�$mF��>[=�q���t���s�}�ꘫ���8VR�0���T*�E潄��9&4�ݴ"`��iu9��M���^Z30����t�V"uK�W,�[���ti��P�r��I�+������i��`��_/�r� ����6��X��\��d�x��J���$�꘽�{լW�H
�1Ɍ��1�T��a��dݖ�-�XB��?J���q��<�L��N!�d�\�z�k��u���I֦��js��CۖV�2�+�!`��6o��t�N�J������aV"� lI!ڣ����en(�N[~��S�H	���"f\Z��qh���V��+������f��g�U��|NJ�������u�J�-ʈ���S$/�Jl[t��k���c�(`�q��?�O��ZG��UK�}�t:%�sdm�I�h�	�t��"�Zq�Y�I! '�O+�u�x����)Z�f���^�����lt�Wa�3���m||}֝8}N�	�s෰TE�W�O�֠~�Z��Պ�-;·����l���0s�3�N�i��抇QP����n��F�V�5�=�J�B�?�P�B�T/��P�V�B!UKU�R}уHi�j�I{����U��)2}����E�-��R�
A���>��������|^ڍםY \Yz�cl�,�e��XX�+,�[�2�l�Je���)��K���V�&Ȕ��n����-�f���^���d"��L�J�}���z č�i�5u����MEm��af6��������Io����8|"-^k£xKT`^.�)�I����*	9�J%*�Ã���@��Dk׌���{�J��o�W_}�^x�-:p|�Za��l�R|]A|ߵ�k�Ր�X1gy�D���Ѓ���D���:z
f�4�B:����D�����E��ܨC�r�l	�⪀%t��B�\��Z����U��cvbӺ���B�j�u�v�6 f�<#͜��nD�EQL�ql��q���
��N5�P��Hg�5\���P�O�6F�D��"y����J����4�� �c�Gb� Y��:�-���ȴ����NJ�\*S._�|�z��c6h�5�������ߣ|�.��0��`�@�c�#\�,x��W�b�_�i5=���ߜ�5#c���_�1��[4<R�K�T�\�[+�.�)h�`�`���,,�XB��+3��Z����^C�p��>�	�r2M�$#ֻ�źs�M����������
�Z��]]�!(ཎ���^�\��n�%�D�a��f���t_L�Yָ;�p�O�:��ځ������ƨ֨�u4��m|�R�JK�
��hv�D˵���g
��]&��3,8��\s�V���C�Y/���T�A�p%�^�
E
�)��X��P�f�zT�=���������mh�E���E_Q�Z�K�*P�)��D$�|����р�(����G��u7�͎��˂�(]l�Ƌ�EWG� W�{"C����FW�N���f�K�����Q�������T�\k+luڸR�޹#�	���@��t���0��!l�����Hí�ᫎ���^�U��ȧa�Vå}���y����i�oҁ�g��=*�D�g�L�͆��QCn|���c��0E����n��~�����4::Fs�x% ����ɨ�熱��F�� ��Ld����sXB��"@.8Q;I�ڥӍC;���N����vF�X����ir�2��'��j�3�'���h*��ł�ܡ�5�f(�j&2QÇ�iEѪY+�&+�%���p*�
�t��f��ٱ�Q�Q�xM"���ic�<p%zm�\GD�:,푲�lϏWD�gXcF�X
AcL� T�����h�"�Ʃf�:�>4F�=�w���iZ^�g��јCLʭ����Wޒ�JerÔ����\��C�R���礩R�Q&�s�Y���_��S���Sgg(�_�c7��"�Ǔ����n$lx�}���D���5[��S.�p���J��,���w�K5��[g����\��������fɩ�h���9�5��?H,��X	�t:8��pj�#�����Vgf&�;wR�q+LX��K��0����ݻy���������|advv6�{Y�ó6�l�����PK�-U�ײL�^~�X�	wa~>�R�L&�+�l�^O�Ŵ�h��a3�O�S-V�s-r!kh.�@֓��s���2?�'��`
�2�����(�y�n@F�j������ips5�- �(�L�C;�K�v��E�eQiV���=Z2h�ȝD����mȐ|R�S��%-4C�����{PEǴ�hӑ����|��U�4���Uن�8```@�aqq^�g�)>�M���L���]/G��\wD{wιB�ѽE*_4���0��/0��dm33s��!Uj.�8���3O�C�X8qe칅<�G�֮�E>BY��N�I��v�����^}�����˭R��e��=�
�T�Qw�0pW�s����ń�.//�f3�T+Ԫ���e�l:I0l�e���7�h�Z�l�a��[�u˖����<�o�㖟�?}���7Α���%t�_�DR_��W?���/gg�o*����`���<�V:l�j��j3�fD�*0I�X\51^s�5t�ܔ35s֩T*��/:͖�A�R?-ϑ������@�F�F��o4kN�Q�/�N19��Q��Q7ަ���du�dP�%�zR��Z����Ȫ��W[V=Ό�שּׂ=Cl�oɵi#�N�t���N{b.���(��IQ�h}�l�5��D�C3�g�EU�"|*]���q~C�%��Z-S:���%r�1�W�5�K��-&v����han�i�.��;����04�������|�D�BN���y��)�gs���S��S�8 [��N��=i�`�aÆ���ݻ~�;{�ԩ����D�O粴��D�LZ~K.\!�-��$� ��B*��w������8i1�|?��gY(��-�n�k�mEv>�[�N���ۻ�9�C����>����{�}�j�W��-.�J�����_�����o7m^�%�Ĳ���޻����˃�Vk��Ç��7ަsS(�C؊���hhp�>��Oҷ��=�8;G���/��Ç�<�����ݷ���=x���?���q�ںu����QYfBt�/
����5/*��o6�`��NLL�g>�iڴa�U�Z��]��뻄��������5��{U�&
.��4�]�4�j�u
�t���q-�q�U�U�?44$D�F�x��Tg��TH0��}]p%���ۣX&f���^K9�A���+�^�㮑�Qt4nl� Yz�=Ք�sI�k�9-:�,QA��!t\�8Co��=�܋b����L�% ��q]�ˋ4�����͛��:S,�s&�Eڽ�M*��Ԭ7dm��ħ������w��G���y�ۿ�=��s|^��[5F��y�q�t�M�Ҫ������7Y�*��~�T)��_�����|�����
���e���������'�x��䲙�L���u'�����h=(R��r���M�������h=!knkdЌ�]s��`��y�c�c�.:x� ���˃��B�A:��r+�uW$0,�Ͳ�U&�Ə?�]>�B�9�0�TE���C}��m�F�'��n�i'��_��K2܌x凌���j{��O(�+��Jј��۩t����Jh���D{Ǖ��C����I�yt�qp žy�\(��Q�$�u�S� ���(y�D��$�>{S�ǝ���^�!���2��B9;���v*��G�����ٟ��-�*�**��Pe��$��[n�����ru�,7D-�q�`�;�w;���,|�ŗ��ޓ�>�K�L~�C�g�^:{�<�v�&V��;n��>��O�\���Q�Q���>�ڵk=�ܳk�;�|��?8s���ƿ�Y�����nqY8y��-_���y�s6��ڝ��M���g��x?TG��ZPah�Z��z�-4:2D����^}}��0Cc<z��<<?���S�\eMr����@;v�$��3�����<�����ӧ�+_�
;v��l�@�K�L�e~���􅳔�2��K�3���C��(�S��n�k�X|��QE.Y����&���
��Dn�µЋ�bf����+���U�� b��I���j��~�+h��#�x�D�~�|�v��|\��k�s6^u^���D@�5@�5�k�fs7R�d<�7@�a��zT/.�C�����8��h�>�9��������o�[L�c��#��)��_�_�JR����!�n~v���[ߤY���B9ֺ�h���q�]�];I>k���~���o�����|?�bá�z�F��|x��b�|rr�F�
�?7z�������뮻Nι8u��1A��Y���V�O��o�C�?��/�ȗ�"YX\XB�����?���W�U6��n���GŔ��ˬ���k6��Ke�"���8�{�t��?qQ��a����!�r�z���l�fm�:�����C3~�=tp�>~̷(�"�j���}�O��H�ť}��ߣ%�Ρ��� !d��� &�������!�]N��.^R>���;Z��sz���i$}L�N\n�UK���H�zܰ�#Iq��s㠳N�}5�������\�5棂4��;7��S�}*�SZʮƝ�P�i��y��H?G�X�HQ����]���@J�j�_*T�A�O,��_`���v��X�r�5��C�}��ͤ�BX6%���2�o��*�*U^kF=�A����{$�vn�FG�i�I�|��w9�2z���k���S�������i��8U��|�g������-�h�����j�Ž�e�ڳg�Щ��7�%t�+K��w~a~�5�T�Y��۶�y<oϞ9Os�%��k��)��-P�	iͺ49���ZXb�g! ��_z�&&����,����>�0]�փ�������O���'�_�":�.��?�ڼa���Fu���{�~�W?K3����=.F�ZgͿ��K�+K��&@d��L��mT��T+��Z�s����(֢eH]-��&�N~{;-�h�jZ�m�N��Nnz`��ŏtJ��K�2���t��9�ɵ��VJ�cAC2��H�v�ֳ6�H�	�4���AT//Z�A} �����?=��E�OE5[���}\wމ��E�zq�G��v�S!��5k&Ă��ذ��7nZO����X8ˊV��Ǟ��Y��>��Gi����_�2����������{���a!a`�Ν4}a�^~�Uq��Y�\3N�6��B�s���*��
y!�j���c�bt���;�����N�<}-YX\!XB��,d�A�p�V49�Z�_M۽g/�izf��߸�Xk�h�+��ã��)�3��r�
�"���Y/���گ�>�OБ#G�'O��.^�(5$�UJK44X��w�Z�2�>q����x��5�5I-C�q��`F���
�g2XM� ��t��>C�Er����/���+���۝h���&}�S��oF�'�# N3p��n
,�@�s�~|V�]4�0�J���"_|�.vH'#�W {?N���	5\^|���#�#�-pR���;Q���b7�fw���[�{^B1���
��D@��w,8����#�<Ĥ��V�^M��������&�Q�C>���5����+L�ȴ��ߪ���wA��8���0/YUG���M��c�{�Mڰi3i���q!���XK����'>��o��;ＳI�`XB��8L�^ݯ�p~����4����H^����j:q�I�e������(�?}�ff�X;_�i��(&����ߣ]�n�����ǿ�=���t���={���̌P�ǆ�}qq1�o�|ʤ������b����<���ùV�R��#�G����j��ٺS�M���� &K�M�H<*�ڹAȏ6{|���9�c:R�NsӐv%��n��Ea�c�y�hpD�k��(�k����t��.Ĺ�@*�}��*�Ǯ�hR^�]��5��ڰG��q���^ؔ���[AJ����5E���@�X�`���T��,���}.����]w�6���� _�"a�#��S�@���D�j�����o�a�b.u�)7��N�?�<MOO�w��g��jV����m�x������歛�ο��𨔞��F����X(��b,�[��a	��r��H*�ɤ��a�\\\�%kRn]����o���h��u�����Kn��)B�ޏh�]7G�p���i!�\.Kֶ�Q�Y�.��\�.��
�*�9-:�,�49���_��s���������Y&��Z���;�hJ��a��p����'��JQ'�V�a���U�5S�L��m�6����tk�:>`j�浙Z}Tƶ�ϸyMf�^�|������y�%�,1��TA�7ڙzq�3���FCo��iA���q��
�BC���r�"h�ș�}�X?N$Dէ�v9�.@xy�j0�Zx����������f�I)�@���Ay�Z�*�T�[^*��=I/�D��̧D �����'��O��x��yI��K���z��H�#E	�k����_����ΑQ��AD�#���n*5��]����������VKLLn�����Ҧ�[�Y��'
�H@?�.^��B2p��:s�^۽�j�
���K�� �k��=�Z�n=���!?����+/��}O�x����KD<L��st�軴qӇhna�G�i��[�!;L�|��(D�q����\�j����!���:��N�Q�? �̀2�L����bQ���A�J�~���6���l �  �&k�n[����x��<"�V�%�ZjǤ�ׄ��K�hPՋk�C���+`օW�@�-�����t,�(`N4�x�������(�)���X��m+���R���6�F�~"H��ި�b�H-M�	9�u�y��Gr$�Eoh��B��p���%*�x�t�}GKL���7R��=��T����c���� �ѱ!j��;t� :�.-�i`x��Yh=r�(��{�n޹�ҙ�r�Mt��ד�ɓ���t6*���tgN�����4<>�F|[\������ }�̅��� �����EZ�Zs�0?؊��5X�L����G�й�)��":Ҏ��\�����/��بhF�3������%-�ԅ�%�����OĜ�;"φX���2�+t�u���Ҳ �6�f���ԕ�l�\��U�k73q�+ZG�6���u*���Y��v����њ������L����;C��v���|���k���\�Kݯ0-m~#Q�q�^wg�-�E�s���y�8XωL�QZ]��RD�5�q�h{�`a�Z�ڨ�'��/./���b/�Tw��qZ3����RL�Y&�\#2&J�������|\U/-�Ňze��@N�U�� �w����7ߤ?��?����!=���i������c4W������|9�<_W�K�`���oұc'����䚍�b6둅��%t�ˁ�Tj�o� �Ӌ��K/��r���:�$����iqa��ܳ��.�H5�lf��&?�Y�	tp4Gy��,E��3���o�IkV���jZZ*��e֐�D�?�O�^GY~����8B��~����\~@�Eg�>eͺ�KS�8��9��_�7�BSr35֨tjK�H㾴�j�&�'��a��@�8�^� z��o�~U?=���f���J�/�'o��5�O] ���ܟ��L�ױM�4�I�����y�%��M.�rw�.�v�~�f�)"S-��`V�B.G9�N;J����4><A�����iav����_b����>Agϝ�7��w�yGb3�x�	Z�jU�KT*-��ci�7�z���P�{n~����O鞻o����(M��S.�%e����O?K_�җh�5�K����ykn��b��nqY(�S�Ԑ|m�.�����w%O;@����ť
k�5~��)�
J���$�/��昨���O�{�?AϿ��<�gYs�,���G%b��AP��͛7�>�j������{��s���j~��x��u(3�E~�CQ��!�9�qw
����Y�!�n��ܮ��ĪdMv�oj�Jت�*�����?S�0k�����rş
"��c�<�w�����v�w���5�N�����։��<�fԒO���Q�zJ��-f)��2"/�`����L����T,��ԉ����O���sHS�s�GUC�*���ɓ"��_����.),��kX���p͠ ,;��!`�����[X��ﾃ����^{�mB����oӳO?%��쀜;2<�6j5��[\XB��,�M/�*g)��d�e�D{�6Y.W��K6�c�J>0JgJ%�zI��a�_D:D�������}�8@��� k���*��U���v�9�����4>4F��������>A7�x��� ���s~��	�n��T^�*k  Dg7�N�SC�?M���XK�cU�N��e�A7S�T��t^ՔM�TI�$^@ק�����?�j�f�_����յ@�2�Y��ټ~��c�V����JۓA�f|�nBפ�)k(�vʦ"w���0kη3����|U*�yg�MASoI&,<�y҅e��۷�Ν;��k��4��[�I���7閛o��o��^x�%:��ij�>��I�{s����[��>��������>*�	���3��7_M�����\�����nq9pʵ����tAc-�^�֋6�.--.	A��Y,���d��$�P�֨H�mDIW�ZbM禛n�����=�Kj9s��L��}o%��^���w���Z*f|)f��I�g#2x�7�����w�:d��%Q��"nq��^}o���ҝ��h3�]�G%t3^��$�9?W(��:��c��Uc7���@�K[�y��9�x]�I��i�4y�>��M�B��k\>f�8=6ſ�g��Gz���ׇp�V�J�����7�=�8�Nж5�d�w�c������4;v^��y�ݴc�.z���rƄ`�9a~G�·�~��G�h-�ޖ��Z��*�\�m�M!P�w��K:ύ�,̣]+���S��F�f	������ ��f��M�F��%��Ղ���|.�J�Z���>{�5�j�$>�@����T�'�|���o��hHo��:?~�6m�D����<T׭�������t��Yj�pL#������n��.ҩS�����t��m��d�噶��1h���'|�(�ˌk�t��L�6I��6S���J�R�<&�������@&:�j�*$$S�ig��6�h�H�dCRy\-b���/���q��՜K	zK��D��ս�׉�@�Ѽ�5�;�j:iu���tM$c�(���I��D�T�tu��(��rs��/�G>�(��y*U�S��W�H��Eɜ���.����򒔃E5B�֟~�iz����W��Ⱥ�=h�R�h��$-.�Q>���4�;�Q�_ST��PXf���i��i�P�����K���r���f��?�
�<!��Zm�$�F��(0�7#?6?�)��j��ޥ�j�F�/�?���?���\��ڨ�m�R�0N���:M��H�^���MN��\���A!{�ߕ�83	y=h�)I���X�M�֓�x@�H��S;6���sӇ׈W+�F�d��e��a�+�w6�&�(H�ى���4JQ� /lG��K�Լ��c���v�w �A�Z��5XOץ�xd.`.�R��@@P��N:���8��M�o�{���
�܍�Gz"\n:N���b��$�:���A&f�{���c�������~�Q���3�o|C*���� �w�&2)�kKT��k؊�ԛ���7C|�Աu�p``�,,�,�[\�t�s�ߜ�����/�F�N��9��J���P�8 Z�~QTU�2�䙤�9L�z���!�:�u&X͛(\���%k~y~@S�lzf��� 06:�дDʧ2i��Y����H3OE�A�ބL6�A�Z� ���I� �B4�.�	���y��ZA�J� �7J��4�q��	!E�����:��<����"�A�v�F�ϝ;'D��@4�V#pD���U�5������/�q�et�=66&���־�~s#�{�ڵm�u����h�؎�D;[��d�ǅ� �m�و
������̸��d�A;�I�ZC��!j�[b�q(*��Nli����ђ������-��Q�M�@Θ5	�z�����J����\+� ���K���:��XM�c#�,�����a�rr�e���@��*��UT͑�A���?jǚ�-�,�[\�V���C1ۦ��*���L ~`��B����9y�#��4hphH���Yj^A[���S��pP$��Q?�=�V6:s�>e>�J��L��ǩ�l	��P�̉�n��D]�🙶%ד����0���)aj�N�x�	Z��	�*�$-O�zzZ�� Q*]���2D�si=55%�A ��8-ca����T����ܸ�07��5a�J��hq� b�T��c��:u�|iÊ��>����Y>k���z�F��ɀC5�'�Z;L�)�]��޸����a���~�xO�/y���D����o5
D�C�y&�3g�IC*�u�t�
�'Ȣ�h}�kb|�D�#���io@R��>��2��|���NU(��r�a��~��W#ԪלFʳ�nqE`	����='�af̗��&��TC�(�_+ʬ-�g��͖�ة��c3�ѡq��Qʨ���gL��:�hA
hԂҚ p����L�\���OKO�ŅY�[UZX���N��w]��ב��x��U|�N�J����,f���)A�I��krE��� a��2�k��3�L����眅v;P��Ql���=^�ԥ�InkA*n��?�a>�h�<>��PFB��&˿�X�d�&v@��T�Q��A�P��0�G��p�0?����l�f e��@�Pī����c���[9;Qe:���j���9Z3���p7�� ��*�6�d�������ȉ@�, ]*�a>M^�y���f<����s5J�4�j-�_��V���:��Ei�[a�gق����|�5��nqE`	���X�E�O�����kV���~ ���^�6hfv�*���F4<��.ʀBkG��t���T�7��s�hQ�ҍ�m�`.���Ξ��'�={߈}�q�r��Nd�ad�w"���|�hC����L�e�`s)�i7Hfp��uJ�І�E���8l�x 5]�O��j׾���\�,������A@J�.�8؇��t��bN���|-�P��=qC��~# ���5��>�|����{�-0���A]Q���fLI�us�̵����0�[o�A�Px�&��'��,���O��@�
����
W����Y�� 7@Y�m[�R>�e��<mݲI�ɞ;{��:�{�=416B��N�!��I��R�AS���w�����+�Hi�L��|�ZB��"��nq��a�dL-�C���m��o�Nk׮���k����1Gg�]��}��x�mr򞔇-H-�r���ڲek[+s��[�J� ��w�#-]��ffifz���g�'��cߣ�'�������[��v�����r�)�r������2�$u]��_a��i����A�0���N����Y&΋g�T-��`����6�����p�q�@dW�Uv�1j��l��x/�&��T0��pm 
�b��64{�?�y\�~xh�H�i��a+�\%�F�@] �R��9
��v����W�y�5n������6�K��,��R�����4u�<]<�B>w�,=��3K����ܢ��M�
,X6�-�� ���K��)�����k�;��X^Z���c��~ ~�jy��n^ς�(ҺM�%�"��"����i��h��j��^۽O���	�����/��-.(��6��26�_G�����k�F���t��������}���kߢ��T(HC�Rm����v�Z�0�!:s�Ů��襗^�`&�亵�jb5eL��)�������f�y����O=B�Z��8L�N<.9�R|5�Z�Jz}I'�D*��ǭ�ps���G�ڦFʃ�����-U��h4;� ��B ��ASq����G�Ž�`<��#]��J��G��k��\��1>ǂ��'�F�s�.Y��A��g�e���5�j��=��0�[Ҁ4UH���=ւ��K#�;Y�J}�I�s�/��, ��,4�<��������O��o�7���˥�T���	*��Wb�ugffN�;o��~��TZ\����Ī���3��*ּ|�A����|?.�y}��t��Qz�чYx�#Gܸc��AӧM7\O��ۿM'��UX��-�[\1XB��,��ړ6�c���|��%���1�X����J��ŧx'k>��[�A�g�����qǪ�IIW{ꩧi�����O~�^�)D���,~���"�D���?7S���I�|^_g�E���6m��[n�I��O���-I�#R�OjJ�I�F{ϰC&f�RӏnV@��r�|����g�-�F��6h��Î�a;7[���A�J����@z�m�#����T�q��u=��q���! ��p.��8>dh���T��k��-�o[��+�;�\��5��L+�����������{k��;�a����${��e�,HF�wO�Q�@��ч?� e�<�w�,m�ϨP�֮R��0�m!��ý��;����sld5}��_��?�Q��_�R~����/�0B�ëijvA������[��i�P$�5�ֻ�{ﾇ��ē�d����[\)XB��,�~#@��T� f�뮻��P��	f�]�yW�!�?�SL>6��>p?��o?J��6
b9@��v"@�
A�m�-c,J.���j������>�0?�ΈFU(f�_���~ݒ��3��bM@Z
�:A�Љj�JJx����daw59�L���n5��XA� ��; ������&@��Zs]�� lc�
x�ڹ��q�@�8�4j|/�z�{ Q�0�C��ZtM��@7��������CP�!@hl���Ƽ��콶��,/�ף�Lw���	ݗ�Jt]C �7��T)U��/��mظ���/�kHf�\Y��G������Q��ځ{X'~{�j<��gŢ�,h�t��i�p�>��l�W�"=� �a�&Z31��E���y�vA~���(��W���;�S����tϿK�W��-.�ۅO;�j����p�a���;y����8��a���i~(�u���7�l��y���K�=K�s��e��wv�&�?$���#D1>2*�#C�Tbr+�1�j����'z�]�b>C�����\������S������P���u@��X�C�<�5�ڌ�6K���u�C��~5�G)_n;X�
�D>�����|��LJ��&'W�M�����NS��#�t�*U� P+#�e���9���j; �0bR�3H�a���"�]5��S���Z���q�q� n�^��0&���@����v+VM�����oetz��v��YS�\7�T��ϑo4ɑ�y5��j���'U�a�r�]��8ZAnUP�J��9���^3A�֮�����ݽ����>�c�:���������]���֭��k@ϝ��o�E��:�o=�m�|=}�#S�筣�L��]K��"F�EK�W��-.���M?d�7*��o�;IN��~�cZ̈́�<u������r�J�ũ!�|~��e��i��7� �ѣG%5m`t�����.^8O�s����5{����ڠ���;?M�cC�/S˯K[SO��衝��{��}�ș����؜lV�k_���,5W�� m5f�5�fv�ݮUڎ9��gMV�i���,�6@	O�X��j� t)��s?�� [	*�ׅlUyC�W�Z�~���ڵƹ��5� �jAP6֤�5>k����jzZϴ��=�֫Do���:������F8�ʆ
���'L�0����R�X�_�T���Ւ�x��)p��6:q�\?���5kh�����7_�u�ޭ�\E��O���G�Ϝ�\6ł�z��2EI�sR�D�� N$�8����2��nq9�0��>�úh4s3Ӕ�f��i~n�����W�v��H�=.��{���{N����;?po��vz�#QU�� �l�N�<A�����4xߪ�	�������THj��{龻��kT]�r{�R���(&�$ȇ響���*�'��-G��VJ�J�J� *(H�y���Ą�𑛕��͠)s:�Lˁ�X�y�puΤY۬O/y���k���OS��":j	��e��v-���ɼ}�,�+��ldd2�.���G�q(��tM��dHd�iO���j�s3�4;=G�rC�06�+�y���O���&��^x�9jv��N���"��5"�$�mh(GC������X0am��p�dYhh6+b�A/��:�l��ŕ�%t��B%Y����A��C�R�jҵ�ma���C٣ֈ	�a ���4�Q6����T�:�Ľ�����7�1ڪ´>5}A4*͡_�J�������5�Il�|��!�f]W��)I8����x�Bk��m��SWR2���6�dj�i7����?��>-���m�u�p�����M��W�h{\�V�L�V���L.۾^5�kKU��לs��߁��ֺ�f�{uAh�\�oj�0�c�9�ɪrz�B�fTX'��a����rÕJY*��9�=���Ϻ�&f�q�֭_O�B���c�i�:�A�/������<���iB*杓 �y&s�\�����}��>x��ZIA\@t��*);\��(ǯ�������8�?�^�y�W��-.!���-��=�p�"�~�ڤ��"?<S�.�6<X@TuY���/��>!�a�ggh`hLH���)����h��v��Z\��k0��S��|���.��C�i���X�g�@�s�Q�V3�������v�Ͱ��	C5Z��}�g���kf[O���������[�ӂ1J�z������4`ѹ�R��6A*�뼺~�P���qJ��5JT;k�:�j�07��R�M6�QAF��,��^�������"���%����ϝ?E?���Ig��>D���,d�0�T*-{��v1���[XZ��������F�~�3�,�4���
�Kљ������m�l�M[�Q~p��<VynAH��{�ї��Uq	�Z=B~˵ڹ��%t��B.����`N|�G��'����LHn0�����f����Nh���rl�T%�3��v��@w�q����K:}�,}�_�Gy�����~���Lsm"D!2����9:��~*//҉��ӻ�f-~��9�̜X�4R� ��҇�'JBJ(&�i'3���\͈�6��A�2�R�v-{��ƫ��U��:U�4��j%�>��5�P��V�3�T+٩6�&6*��Ĭ�T�f��ݠ�ٙN��o��Bh�>����V��R��1�G��:�n�4�G��ƂD���ر�t���t͍7�Λn��3�,���_�N?E�\A��B�K�B��z�6	�3ʝw��g����e�R����G���Sg���i�Y��3�ghͺM�~�VB~�=����<L7n�L��l�,,�,�[\�t*̡�K&E��(Uʋt�0k��52$���k9>�=3EKK%r�R!Ҋ
Ei��t��{,�&�=��o��vj�:��P$��������@���?��?��2���@7��ɚI��D�ݔ�W�Z�ҭ�:Z��+LӹYM.�+����T�ǘ�]�ES�9�i���ꀮI���J�:��6�s�pH��Û�f�5@����(���>j�[�b1�=�*8��L�[����9ӭ���s��"s7|t:�Ha��^qh�Y;A'O�����j� ��A~��%��J :��ZPX�RZ���Y:r�yL�CC#r/~���s?MK��~/�f�;�����ȱA��cg@���\%?D	ڷi͚��v�F���%8ך�-�,�[\�AC*���$ZD�܉���S347��O�:/��+�:kDc��f�R#Ҭ���i�y(0S*W蕗_�W_y���,�2��V�i~|{���r�e�yRK:���˴cǍ����o�C�N/�������471Ӻ(V�J�VikI�&Uͫ�4[	�]�5y�Шn����怦�Z���k�9�'nV�ӆ)J�j���7���樫`���y���ZLBo�Ꙅ-�E`L��G�m�{���G�7��Y]	����Jz��c,M�S��4�K�b�M��K��w�}7}��XGN��<'��V+�4�����bA�_z��bxp@����-,�.�K	Y�I��D[MH�N]��jm�̖�iN�ފ;�W1�Wh|<z�;;eM�W��-.��v3�Ji$��VA
~��S���d�
��Rn����Ayx�3^�i�5p���Jb19(,S��Y=d�
�먴���(>NM�Z5:H�l�D�X+CT�7��5z����=!����FZ9��T3����oZ��a�V2Өm�L�7"A�ۡYc�kQL�МAjp5�@� :́kX�ł�Ħ&t��!L���	փhl)��k�l?t�́�i@� �k�Z4?��k�mWn���j�܎f�k��B��@l(J��(�1�U*���P��D�z���6$����nk��a�o�!��q�tmS��8��L�?q3 =��ãm���:\wq�(������)����±���ޢt� �3�?��~E���؂T��� �2����x��{4�.�p�,,��	�w��?!���>\�]�q��nq�`	��P���VMM��� �W���7�I�S����LL��z���8
�t�J�=i�(�&J��>kU)j�q9Ҍ�Z���m�y�[�_��I��G��g���ޒ�ѕ-��&1â&����a�w��(��+H�Asz<��ig4G�� ;h� q�F��xt@���^���A�C���65_c-*ས�i�=lG����b2 �믿^�}������8�����W\���=!kT�{g��v�2�6Ղ��o���Ր���!��Q�Ns�a�Fj�j�X/����XG�]P��ZF�"(��U� �7��dh�+ҧ>������Q���Q�D����?��,���Z���i�8 Č@�k��fM�N]8����� 0:A_�S�EZZ���6G�`)I;n�V���2��nq9pJ�E�٪3�c��+AO��e���.�������Zk٥%֦KT���\Y�q�)1a"�=�Ht<:�As,2���}�v����O=��>+���	�@���!rR^L~~T��Sm$�&o�<��S�9A�V�7֏B/hJ"u�y;��Z.���F�s���;w
Qj�t����j*W39̿خ)e �� dmӪ٠c�Y��0���\��� ym�o߾vԻ
X�
50��:!L`-����Z������k�=�ڱ>3E��x��uaM�>��u�b>�W�U���^�(���>�~3 /���S:��X��k�;�q�@긞��X���Y?��5I]k֣�>D薗�J�bz��� �Ш�4p���t�a���؀�Nb���/��-.��8�Y-�JMʬ��y1�%W������Z}�&�ի&����� vRQ1�N��ÜJ{L	6���@����.=��T�B�oP��xH#�	������ԝ��=f��܌�ƫvR3�TۡjG4̩����5�\���?҆6��7HS΀<p<�h���p��õ'���A, S�w��@�IA#��0���b)��p��C�W�-�}�Av�
�q��z�5��}hyX-^a �n-=������=ý��m�*�l�sDeg�m�J�7S[��ie�P,<�]-�jTp��e��G�V|p�T�45=E��%vׅ�������v�tj�r�ynn&"�'�y��+�{T�z�"��"� �2�K�����ϝ���Mkaq`	��rf3� ���ԯ7(�e(�� ��يs�s�e�N�Q�K|�yt[.EiWu&M�	OKe-T`�����b���V��fMxl|"����СF�I��}br�F���%���ȡX�t5�}��ԗ7+�)��Q��eL5{��j��󎘒�l�B�7l2��q�|aI�(�DM	I+!�O#�A�Ђ�>:��8�w�Y�� _�	��1 V ����~Y���1��QA@��U�6۰�� D,�mFq}���\?������!ta��������
0؎���p�l�d���;�[�.�v�K��-|ϑfL:�e������xL�˕�\����]���y����@�L6O�f�*s5�f:�G����-���-Q���k�Ã!�:�[X��%�sb�Z� +V*�8�Ҭ5�[\XB��<�|֩=�,��-��Bl��.Q&���ay�H���<?TYE���&�x����Ai��mq�F�6�˃�R�Iz��ML�w���z|O�{����?BǏ��#��VщS�������ж�ү��7z�fW3=��íU�T[�A{��)O U�����V�ѐA8^���Xq��Kƹ�r��� Z�v��{=����\4- yb=�����5 �hx��CH@y]uC@[׊y*d`N������u�ݻ7n5��8B�^��z1�F΃�!X`��b�;�x��c��N��1�M-*L�i�F�ߝY{�y.W�1�������hb5:�-��h�����ߒҷ舶a�&t���o����JK�|�}�Ek��ťYZ31)�t|�^�uӵ��{"�LL��S'�ҋ/�Lo��UYXE/�ln@\@W
��-.i/�_�ү�A��W�Ѻ��Yc]ÚtdF*ϱ�NҾ�(���R�.~uԿ��3� F�w�����n��&��^{�5:y�x��y7�&���)��_��^}����~`��m��T�2�P��3ڦ��Xة߮~t�N5�J{xk5���OM� 1�!�����YM� U<����4�P3�F�ئ��Ad �(�)�kBۧ����؏��G��o���:@P'N�'�	"�g�a>��B����{F�u]g��r���� f 3�,��g{�3۲G~�=�c�zoyyf����i4��%Y�5%���H1@�ȡ�:wu�������/h�������]U��{���m�7��p����1~0>��x�
�yC��a>��1����x=���<�_[���؏���
����WߐB�!���5r��{F������{$��Y�~�u.�t��
@ٛ��r��1����6g��Ћ{6v�O6oZ/7ݼJzz���d�9Y�f��F�����ߨ�^�����x(�Ē@Y 	 =��}��6�\&%����Z�T����5�e���j�$�vJ�0,�8n�>/����8yZ�z-�n�L�,�i�,W  a���k2|��Z�M�-�d�҈m�ss�����%��?��n�enZ�@7��iɤ���w�QL{>kIT�J���O�B���-x ��HaQ��� �q<,b?:c�8�mT���qt��`�ê�2^�Lp\k�� �� �x3�`Ȓ.$�a��F���kIx�7]�q�q�9"k׮��t@�A���((��c�V����3��7 󇲀yc>�s�3y�Ix,q�' c:w|��t�໭꺀�?d~d���ZU�o �ݿH����}��N���Ke��Z�i��`=O�:&��.�����e߃U�-Y��7�~ʵ�����&}�yY����Mal�L�D�c|ܚ����ӑͥ#�n��  z 7"���c�!�bHDK+`-��W7ָ�Q�-��ͷ�*����;����c#j�'�@?Rm6䓟���~�!k��M������铧�i��;���j��Ւ�N������wQ>���䳿��5f���Q�/��H]��G�s�6�P�%���pOs�S�����t,`�2��x �� 4 {�8�:���}�k�=W�6�d��1q�J�o�}��	[x2��q.Y��j�y�`,($��� ~�-�� �
l59��{6v����=�n�]�9p�P���g��kbܸ7�5�T�j�wIE��x(�����'�W�$�u�|�-�$F��3T/�$�M���-j9o��n��Cr��ai5U�ץ�Dc]�I�}�z����m��f�������/��ݻ���9L�]��>7s�Y��ee��AY��_�z:�83�ٴq@��تKT�t߮j���u.�I �܈��h�bc[������%C�A��$��k�����+�m�WR-�n��&���'��ذϟ�`�NLM˥+W�.��
v.��X��1���VT�����m9�ǫ�t��(0p�����%.��F�r��g&�o���d�lȊ �;�����LI�1���>�����u`�B�ą9aL�;�.g΁ӵ���̝D,�����b�Z� [ 9�Ͼ���91�৪�S�����-R��������<�~�<R�r,�^��� !OD�1U8�^5B�Q3R��n�*�rSj���w�]�<Yn�������i�ve�`ӫ��:��x���b	���>����MOMH�<'�|F+�o�}��\o4��Lܼ�&�*X���l�B�}��e�&yg�>I�s��TK	d$ �@nHԊj[[�Hȸ�S��Y��v�:��<kVؑ#�$��I:�77������v;$_���dz�h	I���ߖ�}�s�A�g��w��׍��ʞz�r��I��ްf���o��*!�xaX^~����;��V�r��%�)��BT;�i4e�Gbr��]�~��N�����y��OK�#�@����Ke-�?���8��e&�Y�g	�=�1vk�X�����R�F�rB��{����f]=�_��gC�X�Z ���[��dcQ�y��k��1�����ll]o�����r
g?�*� JW�=K��-˷���Y������I�'N���B�fJ�{a�U���ܼVR��?����MYkU|���\�T�ɤ#�N�F:s����eb� �p\z�ݺ>I��j�/�g������@dA$ �@nHb��'�1�eŦ�z�J�hԞp#6����� �b�ڡ&�$�K� 6�3u����~����,f�?{N��OI<��.���{g����EK��=��#�X�2�K�)�F�$ �V��Ao4��}�a��u���Bv@c{M��!(�rn�k��3��{�{E�P�k
C�f'ر�8A�.�LK�O��gR㘘k�	��f�cl 8��������@���Z��7���M��̇2曼0�nt��r֫3��z?s��T$�� %��fے%��tF�i��rIx��a,}��{�op��L.o���vx2�9n �w��=�>�x�_�IG�oH<��M�2c�j�WGep�r��u=��(����:��YK���,��ȍ�1 ���c�`j�\R�>uB-�W;�֗/_�%�VJ_�"�\�R�+;r���e��2�]��G>"1��''��z\w��^2U�2�a�:(a��{h�
7�����+�!��1W�\�u��>PDM�Y�`�� ��d8Z�tZ�x�aV53�	��o�����-�Ы��gĉi�����N�8���<���L�|q9��9�dXF淎	�t�3>��+̪��2C��n-����{+��p]�\�:���ߐ�)J�k���XƼ&0�rP �#����H�(�kj���9 >���)�#�ױ�M���qDF�4�8x#�� n���+��A����>|D^~�e���;e��-�ç�r�}��?=|R�/��3�N�[��Z�h&�0 ��[�D`,��u =�� ��!i6��rI-�j�a�uɉ'��Zg�Р%�V���&��-��sH��}8�$ m�m������#H��hK�9l	_ ���|O��%����\�s��4��p�6붏��\tk��Ɇt�G��m$5����/����mk
�;���4��\j@f:c�l@��76���c���8��0��3�� �� ��M�y$͑U�$4L@ñ�Nz���D)��A�;��?�JIg�S��;����:בY�%�|\���;�1��/��w[���3Ш����|�N�
[.��RѶ�� �QW�N��qIe�v}xmp�'N����[>(��ה�}��V�0::"��w�����ټ*ӳ�t�m�t��ZWn�*<Q�_W�����w�~c��f2��` z 7$�x�����hN7躹`���Ro�d�-[�"X$K��^�S0k+����l�Y���>�������-[�X��p�
Ӎ�1ʫP��|I��W�l�`�ks��e��$:�d7�Qʺ���9W�|�pƐ��q������;��߅?�F@Cf9����Ը����\�.q =>�Ŏ�  �>$�A	]�T2�99�i�C��@�"�5f�c|�nn��ٞ��q?����c���y���8A�>C
�0n�����\����� ���"�M�{%cW��t�2I���F�*�j]�كb�g	J' ��	�&��߿h�w�_�x�	+���e�0s.�Hw�¨��Cv}$š���
�f۔�}�|�w�����س�@=�� ��i�&��F��lr�`1}�y��2vuʁ_;b�@~jz�]��Ue�c=��o�T�}��5�ڹk���~���G���~���p�������G�J���՗���~X"��D�I��B���xC�q\��<��T� ]&k�"��&�ӥ>11f`�dt%�w��~�qҳ���ZHR�83�r ��f�o�����w\c:��O_˄/(:P&��F�<2�� Б��'�aKV���(=�>��^�U�)[�g�3�pe���a�����~�3-u6��_5��0K^�r��q���^��G��D�m"t<+�u�<t�Ø�0&B9Pn�xg�S09*��+�"w�q��A��K$e�P����c���-rX��|wV6nܬk�Te2,���S�"�/���~����#4Mc���@D@�%���m$.�V-��2Z�V�!S����Ε,�<��r<���F�o*�5���]����1�W�25>�m���'�w��]i7ʖ���d4�.Q��m�v2��*�u���0g��ē��mvs��-.�����@�Ns؁�<0�n���}^�2����ܯX��g}�K�,u�ϡ,@8_�3,K(2$g���|�;�	�������yr��2G<cB� �+�0��{�"��-��Y�w��>���<�)>_���̥jqg(p�Ƈ�B�7&X���f�SI�wc
���V�,�B��C ;jȹ�g�L�"�W��3g���}�h�z7�Z�%�d�˭I;�I����կ|�~�a������ܹӔ34���܁��9yg�!���%K�t����V�����,@����i)(�������P�a��//�rC+��H(j���*hI�27S�M|�I)V\��H4nq�t������h����*@��7�f�M�,)	5��mboZs&~�ܯ�뺙7䞻�Ƀ>(��#�j�d��K|�t��5����puG:q\��b&&�@�% ӵ6~`J6=k��C�=d��e�밾��n��Ų�=��q���,Py�+�1~(� ���)j���*+�L0M���"U->��
�u�s;s挍��*�}*��:!.���.�����L�u�]az5�h�K�h�`����2*0_�W*���b,������e�ݯ��J�e��e�ۗ��+6�?��tqN���)�֌��{�]w�}N�]��c��SO�Z�;ԕ4Z����5̤Ҧ�@у��ʌ�O�șs#�R�$��Y�v���{{��Ϋ2��	��Z�Պ'�{ "�r#�N$�usѪ��?��u�n
Ec��D�`��?��mVzċM�JE�z�M�l^"��T�������Ę���*	U�(�R�������Z�N���ruΔ�_��_V�	ɾ��ɏ~���n��w��KtC{W�x�ǵ����~��>�W��T B�^ԫ�F 2����pX��i� ��=X�lU�>��&�>���L�3B=��t�x1�6�{f6==�Y��B	��NkCQ@> ���Oy�^�����r�0������ �Cс�Ƀp�j�`��ݿq�FU欋M����׌+aH��6�����ܶm�ʣ��P%�c]��eK��E��w	��;����K��F*�����F�}�ګF"��'��Q�R-��,����^`�.�ٌ~�j�GR,U��j��"��  z 7"�ݡ&-��Y+�A�1)K��ܒ����H��;V/���u�ι�bu �(w��"H�R�R�X�cPn��;�Ⱥ�vE�򕿑��iqUk�j%i���=weW�N����3#,@��nn���x.��:3:oX����܆� �{ƹ 
(%d�㸴�	���c�lU��������X A�ɘ5���|�L���39�1_$�qc=�1m۶m��p��rW��}�L��~�^+T֔����{G ����� ��q߬�'3�{p��x�3��y�)��U��2)�e�T���&"���Ay��J�A> ���:gxQ�!�r���Gh�!.�3,Ux���ǭ��,����7�(�I�Y�^�_���ju&h�ȂH �܈�ڭf���jy��F�2�K�<zOXU��M,>��>��,؄��0�F�q�S)�f��U�Y�< �;sХ��~�������P�|�%�P(ֹ���[:NS7��3��]�b��@��0�nm��
�T*�bf�O)X����0hwR�B*��5O���nu�����0���2�O��̰|͟�NN|�� �iUc^p��2߲e��+z׮]�����{g���sz"0&ѰU+����w�m�u���<P ����~B�s�:�����c^���FA�zUb�9AC6�%��~!!K2��q�6z�SO='��3
�.\���!��s�e��%օ���9b��Gd�����m�L��G��q͚Ԑ�����Gm�Y�������&��=�� ��!���nj ?P�:��%B��w���b���־��^]7�e2�? �.M`n�ľx1-�P2b�VK������\�l�s+Ќ\�h;J߆���:�%2?g��,%�H�X��1sl�$���i��}  ���K�E`��L�c���K�3���V��q���� ��x��O����
�6�,7�1Xg���F&�: ׄR��qx�Y��2`~��֠�)W���a%�����G��p
��>�ϵ��]?ֲ��}o�z6��(q��H�B�	)�N�2�x�hX�W�,���rU^R�w�{�'����L�x�]y��1'��9.�X$���g�	oB��G�s�êςXG/�����O׫o�@dA$ �@nHP���,�����z>w�PXM��X2e �%�B�5��Ջ7-�)�Hw Y�`�{�jV&�{!  ��,�a��*��ry�6f9v������<d1t�p����� a�.,QX|���6��Z	��W/��E�Y��'\i{ �D5 ,E���i��|��� 4�B�>���f�6@nn?�K�pM2����5��I�2�kǬ{��������`��&s ��qP"�tH%����p���?k�}�y<��4��yT�:�x²��N�d��K�;�����XN�"�mR�.��;l�!b�/�����ׯ]k��{�3x��)8{�`5�΃ԒJ��VwK���)!ɤ8�d���e�G$�Ey�[m�ld����H �܈�"�1H
����zvnF�
3V�R�V�����4tS��֗ؤ#)�����aZ��j˭��*"ⵦ���{�ڐ�&�zuī��X./��\�����n�Q$l���ߪ���d;b@l|�!�&7oYH lY�	�Z���m�9D:n^d�3+��bdCR�2V!�� Fp��#��	`$�A�5�� $8����j����!P$�����3���@@b�=���������w�m�I�,X1���i�צ�zN{�~�ܫ?�MJXZ�lC��x����j��N 4*#ȋ(��V�<X�A��i��E�I)*�cL��o�v�d�z��v���RG�s^�ŋ�����$�k<��xĞ��*��ƿ�v�Ʉd��JyF-���������g �ʤ�[S�G�}&W%�$�le�ʁ -.�� ��1	�"q�v�V,�dnZ�c��Q$����vX6��d�'����%�8�j�q9y���1�4�Ɠ�!���U�+�!�-�M)�;Ћ���;�+�\Z��5����A������%9�?��p�����4C� ��
Y�,^u/��;��V{	�8X�Q��=F��W����p�Z�^�ޞ�Y^ ) +Y�HL���^č#Q׻�e�Í��t���2nt  �M.�cǎ��ڡ0�4�"�ΘX���u��q|��� OX�P*��^���v{�ӝ�7eF���<��{�^|Φ.��*�M]�Nh8��L��,tT�<��<·��-x�6G#i"L�b����Qɥ�妍i]ǜY�]�܁����bU���굫������ҿh��úB�K�҉����%ƕНW+�ՖjqZ��d��[eǎ{<NF���R-�e�Ҩ<���r��1��G�:<A���C`��  z 7"!݌�a���z|¬�M7�$�<��mr�W,���dSS3rn���>uF���2%s����RP��j�X����W6/^�
�}������eI��M��qyG�Z�=o﵍��Z����$#M��@�(�˚]h�k�
�����k�3����ns��G�@��[�۫2� �5�c��zV��[�2��T�<�Z�#�ֲ���
���`�^� ����l�0�`�kAA�g�6�L07��+wc�>)OI��BC �^��gB��\��}!��N76���e�+�@ؕϽ�w����,S������{g\�b*j
f���Pq<!Ըߴ�f�7���d�Z���.����7�/��/JR���菌ܨ:;'+W,�����g5m�n�V�z,�3��߬�˖�~�c9q��>�)*��3� �=�� ��!A�˄��@���ˮ�Joo�%S�O�˲��-k�;�+5Ś'N9װ�b�Ē��%��_�n�&۷o�\&kn��G�S0��ʫ�)�M�☉�N˟����Jڣ��W*�	c���V���7��k��,;����E����'A���҄D���Mm4�
L�����ݘ��R/��4����IX��c�&�k&�Y�;�T��y�|2�AQ`,�}���N>Ƿ�k����|k�P�w���'���I�k��֕�̮kTh\��\�T�8f�������@`�q���@��җ�Ƶ�M��kEdr�(�m1b����[�����L��M���o}KJ�9UP����|�F�8�O�G��0Z��c���t&-K��e�ΝR,�dbrZʵZ{62 z "�r#J(�����,��v�27;\�o����X��6�7��)�޷��^�z�%_�ˋ���-�O~�礻��Z��ٳGf�&m�5zX� �l%��X+�⬺�_�<*�ZQ~ᗞ����G�<;.Ǐ�������%W��5�罝a5���l�J��\�,iMCX~:Y[X jZ�T���^Z�y�%�b��N'�cM� �{B���l���M�5�&��X?P�Z̔�y8��{8�|�O^�k��h����MNvZ���w�˼B���Ƶ��`en�������+�HR��f�sn�����{V�0?l���$��V'~�ƺ�>|L~��v�	�CV�^��CN/^�
D�*W$��Qp�����Mټ�V�|e\�{�'�yP����	�_P@䆤���!w�H@ʁͮ��L.��M����\�s��m�h.�^�D�Z�f���MĥZ���!=�K&�&��r8l���WezzYnF:>ɒ�˥V-�~��1��M���,O�,����Z��� �������?x�~t/��Y�����.c�N�1s���鍀n$%��I%p�}Ҥ�u�e���s��K_����޹o�ܜ'�J���W����:P��{6��*����خmϊ��E���v�:�_���ӧ�c=$����jed����쳯�L�"S��23W�R7�)�NUkW>/gΞ�����lݺU��r����}J��_������+�}�23]�u�6HF-ytxCr��+�B$jc�m0�H�U =�� ��!i�Z�L2%]9P\v  )����$��F�]�r�!g�]47(2��ݎ�� ���O���d͆u�s�n��޻,�{f��|����Ȩ���8nKϫ�*���5�W_���t�d��=��/ɢ>��b�y����{:�4�QZ��en�Z�v���K�4�q���`�r'�o{pL�c�9�[[���9-{ �fX�αI�J��9@,ݳ��!���5�������&8mO��+5�h��)������? �v�����\�|�T
�s���X��zP<b �����+Wʊ՛���J(ڒ.�sϽ�Q��2�%��G���ey�'��������o����XR#捱9'�5�iB�,}<S�Tښ���KT����lC���9K "�rC�I$[a	u6������C�Y����SO_6�r��1g����|ONƧ�e�P��n��
�g�]��֮���~H��g�IY�d�ter�� �dF��� ���!�j�`ԯ�z�q�(���f�w_����G���x63ȩ �-)��a�G�
�k�Ę�m��c�cӺ���� <�ms��x��d��ǚ���_^fY�
���B�bֵ̚����+���!�]����$7R�
k��Y�9
�'����NǇ
I&Ҧ0!1͟�N$�	/Fԍa��J�z�ócme��ԂK�Z1&Cx��;j�~��IX�HzO�?n4��JQ����UI$ch~.SS��<m����>!�\�)8����Zy�\�~�ȑ �=�� ��1э�ZS+��8�]}q�6I��!��slt��g�Gy�!��mF�l��;v�{w�h��)��%Ṑ����W���d;0w!��d<e.�Ҝc ���R�e��C�Z�.�5�;��	�>8��	��l��E`' ���=xz[�0�qg$��	^t�C`Aܘ��O�[�$�����Gv�����ieS��F��)pq=��2~N.v��~�<=��>��D{Ν�Dyd,�0=Ҙw���mU�V��k����|���ԅ�G�o��O��rd�r��QS���VW�d�R;����y�*Cc
�a9y�\�4*��K�d�a@�d�xQ��� ��H(T�'=�� ��	UJ���hQ`GF�a�n���{O���Z��*R*��
y�q=vb�'7ܓ錁4ܝZl��l�"K<��^x�UZu�����KV�w=z��m+�~-쑣GN�~jnY4�Al?�t�qK��qG3��O�J!(S 0HDù /�yY�F+�Ie��v&��"z�����!L�q�>�����O% �\��	�d��x�� �	[~���}�u�x=�m֯��~πt�[k�j��Oy�������Ð�?��c��2��|��tA�n������jX�h'�u�'��<���P�M���۶�鑳z?I��r��)yg�^�:!�xҔ�|~�LM^�����m�����Ľ�y�w�B�Z��ͮ\�
���@D@�E7�h<͖Jsw3, Q�Sӟ�ZБZ[ʥ�̖x�U�_��]R�%X�T)X�n�ܼy��<qBΫ%�������:26\4y�wd����~,�����lp��墠�0�c��-s��=����TU)w��B : $�x�4�Ԧ��F��&���% �]স�\Ҵr;�\=뗠B�9 �-u��<	� P�=��L~�R���úy�۟R�1�>o�d�#�,�3��U(����?��*2�eg};�
��;D�����i�ܑ	B���$RU��],��B8"�\��
�U����:�:�\��2Ni�Y6o�f	�}�������^�{�q�g_��G�������k��hCu�*�G��o�;�%n�B��H $�rݢuJ����~�6WfN&���𑣶9�&�V�J`Uk�1E+*�͕�ZrXͳs�d�Gy�J�V�[c���/�,o��g�06�F�f�K�Б#�b�,]l�h���?+��)�oK2��Ř��<dt�訆�%4׀�*b��F���'�	�c�l������U'���vfB{����Bi���O:�1�mM���t���	!���]�֝�	dh����E���0����b��+WL����(�S2��J
y�I{�W�Y� Q�ÄJ�?	x�y����p���n����'.I.�+�>�aXak���[�f]�=�~���9I�X!}=������K/�D2�ݒ��<f欳x�3�2j�Wt�Uٳg��^�T�H��XF;�.�<g��r��q��׾.}�P.K�v�|���H �,���u���pR7����/����x�X�s�.8���X�P��R�ძM4�6W`Ŋ���d��ҕ�Ys�tcQ��7����1˵���c�'��/|�jWe�p�Y��sR��Z��F��^�x�m�(p��K�s�ò��FL�uQs�v��&�A����B���G}�w�7����L����aZ���[��]ی�CY0�#����fn��毯qM�G���G5k ��lK�,�����{����LuT,����qY����X��{>컃��^_=;���^�(gϝ�e+V��U���'`�͖���J���� �V7���蕗_�W^yU���%�]85l<+V��z�j�	��r�ʌ�d�^�V�cQE�-Zb-W���g���Ĕ�X�R�,[V�����$�@H@�e`��vq�B=��.������Y��y+;��v�w$�%����ų���w��I�~,�C�)�ŋ獄���'O9�pl��ܺE���o�q���?&�HM��q�|���ܤې��ۧu�W�PK\ˬ: �mZ��g�p��%Z������2'�]�ן�g�&&$��!��v��)~	W(?Ph�J< q�[�҂gR�f$~�dͲ�Zu4��B�F8T:���F��\J ��ֆ�w�7���|'�<�6|���1q��S@�xԭg3��X��G�|H��e����e��we���>��'de�%=?b��P/��������>�=�n��W,l�Օ7v���]����T�!9y���:="=}�z��3W�nqb���Y�S��j��rOO.h�ȂI �\�lܸ��z��c��������n�`����-j��ikl���a\X芮�!�: ���h2j@4=S0p/��u`f��e�֔�\�%5�u���X{z�2;}�6�}胲f��<xD���3R��N\�uز~렁e�5~���G�LFR� A�����g�ӍN��ߘ���R/&~1I׶v�^"]��d4ƞI��o��X7掵#�2���j��L�w�e29�9�Z�ʬp��M7�dǃK>�3���@~���.�9�#�cx؁���0g��h[������N��ݮǾGO�x�>U���fd׮]v��K����a}.ڲt�?�i%�h7��"�͸v���Ti@��fOy$����z#d������i������_�'R��ߡ���WM	d�$ �@n@��=�|�Ѭ���%us$1��ql�
B���m۲Neјsz[yW�%�՛`ө��L�yW6��W cc�d� rY�U����o��@�?}H����N>��}�Ld,���R���0�m���.Ѹ��B����b>P �	����uZ�.A*g��3�����{u�dkc�PaM�� ��8����� <b��.�50w @��q/`:�yȴ��m��==v�^������J�1O$b|��#�w�^���;��Iu p]/��{�O���DB4�Pc�'���1(l�:6v��m_����c�0G�t �֬ ��<Y?z/Y0ߝ�9v������<W�U[��~���)�Vi�8$����)wͺ��LI2�-]��۬�Z˱��Ui�e,�3�sJ�rj��Ԋ�gA����q�-�Ta�E3����I �\�\�x"}�ԩX7�x�k.�=P�F8g��1�!o5:�*:b��
�H	K����d�d,n�¨!��s4b�C��A�Z�VU6�ʢZ.��{�n�RmV&�/v��},��M �b��ə���p? R�(���5�g�8 �p�{<��3�� ��d�10/��a��� �p��@ɸ4:�a���( %������xw�y���dp�Dǡc���+W��� �x���߶y�g߾}66�w����5"�����o�`=ùf,�}a�p>k�Q�����1�kb9>��%���Z���DG{�Z������A8�n��  ��\E.�\�w���� �2W*���fC��<.5뉎�'�~���#�
YXTp�==U�$>pėJe�/!����A��*��p���u5�,���u˹s#Y�l2 ߸nn%l���Y$!�xf����ǣ�)�!ȩ�B\��'�B��Z�n���M-��s� Ĵ5�X�l�\<F��q�DI�8{�%���L�޲,w@��rw��P(fqZ�R��۾V���h�1==i�4��`���?��Y�u�P8`�www)8��2&ē��:�$�J]���]��Ӯ`�/͕���F�cd'�u��x���R��1�(��)�;�j(� ���~��	ٹs����o��в�r4��7l���O�ִ>�X 8���u�"��-��v-r��.�����IqH"`�\(ǎ픎�U�yb|(P`�t�s�}����/(�G�@���r1�sg.I>�չ;�ZW�60��Rv��0ȁ!U���ͪwt��k#4���x�c��dUq��+�l�Ue�����+juW����{hV�(%���
lY�S˧@�#rt�{�{�yX�k���WoRc$�� ��nQk)��S�66��Y$	��8˹m�rc+W%�-3��+�r�p���}m$���d��v�U��m�.!���:}���X�j �eKMQ�4rN⺹'uXm�Zs^����A��7q|�r����X�e�~/q+�e�E��`8�1&6u��I�q R,cc��J�� x R|���pGC�����a����D;\���P$p_PDz�! 
@����`��q����N�~�r�x�2�y<K�`�3s�sa|���pX� �T&ic�f�a�f�X�g|�!�$ r]�t�ul���hl�Q�e�O�?���[z~�8273� �3k:Wqyx2����̸Ta��u��yG�
�mbbJuw<�S^|�Y���仩�+��k�T�;�8}s��*F��H�q�Q��@Y 	 =���t��T*^lVebr\&��S9����ݭ�
�	#p!{�lqN�j� F:11��j)I�%��SI뺆%pk'�	�� �;���C�3��X>�����X�~��2��[�X|��cACB��xv�u)	A
�y�f�T?Ʃa�> �� �$)!��7�h9.����_�Z���c����)��q�bZ���]�ܗ����:�*�5yq�73�-�R�^��*Ir����9�ea|����"��(\���~�F��5���t��nq 7 �c]`��PlȜ�o��z�B��9��"�+��,�0��ón>���P��ʰ.�r�T�J��)]��P��{ǽ��[�n��yɀ��s-�=	fh�'s�Λ7�bkQ)��̙�239!w�u�>t�'��������5+l��#W����d�MuV���v�2���` z �-�����mg��
O{=��d���V�ˀ�kZ6��EX<�l��Nh��n���MNy�t%��m7��Z^���%Y���u@�8�\�g����ޑd�%�xK���k��XU�z͖%�E<�`Cf��.h�6� �c�ԅ���� ]�:~MkPX� w�FM{�kx �l<����������j Tzp,�hc=!�Ƨb���⺸R���h]c\�O��#��`�����(:d����~X� %�ω����!,��l���X�渞��<����e��s��iP��7��|��W���G?�
A��9��X[���@��np�.���6d��p�8u��n�LZ>��O[ܾ=���s�R�L���7��;v��@�*~��8�NϠ��M˳Ͻ"g�/Z餮m���SY0	 =��[n�>^�9v����a��3��:Y�n���eK�e���S���g��+����j�a/]�B7Ҷ�� +VW<��V�N)x�<R2������ZZ��%�:�t%�����l"�kzp�C�-aCG� 9|���]����@��L�93�]ɕHWW�8�!T\Mu�C�j�ݨ�`��9횜 @���!�d0XǬ��ۜ$4<�sc���bﱔ®m,�㹬��u���tHa/��`�2� �����?�n��;���+��{���V��j�s�Oz��:�?�j�zM&�+���8 o����Z�V6n�"{�~F:��6|朼��ٱ�~ٺ�V�Pa�_,��W��~Y��6���|��Ƈ�כ����Z�Ǣ�����}V�_8-s3�2пL���Fi�jGdp(/���j��O_���x섍p8 z &�r�244T�8}**�LRڡ^ku�b�2Y�a�.R@_n�f(}�����:�K���i�h��Oʡ�G�^P�x�$����ǭ�ŗ~bV;Z]|�ֆ�����D�Y�f�1ε�3f�ێ��˵���b�ՎՈ� ` k��ᮆ[`�"; 	1s����醕뱆���wT�F\�V,^g��N�;�h�����5�x�����`��Ď׆�=��ٹ�j�$7~֡��]�7��*��&�a����� T��ٌ��z�]�x	o��\���R,V�dɈ[�V��sK��9J������|G�茗�IA�\YH��?�яX~ �5��^}>��>����zT*e9t쐼������Y�EC���6�O_zQz�{��|H��)�pnR���d	�PT��;�ܮ��1}�.��x�rd�$ �@�[t�O��L��N���Euc\���-2�x����K|����ɶl�jq���.Z=1b�5/�	<6td�ߴq��ڽS����RR�����e�u,9�FaŧR	�+8]�<*����?�a�4Jr�¨��o�G��Y��<��%�K�q���N�{@Ʋ4v#�)�\�~O$B�)�q���=+�Խ�[�ڮ���KNc�0�KzW '�A����1G(��م)��5������7�����0>���V8���&t�s\�'������
����r��mx�3&&=�:�p�[�P����DZW�v(T��s��}�vi5u�H�rFu�0.������� ����<����>=�۔Zܡ�E=?,������lU-�?���`�#�y�Ǥ��C�A9e[�K�Y��^����.�u�Mr��H4$��p z �-cc#='N��FP@���U˥+�gnb�V��$��� {d3���=]��cǏ���JR7dl�=�}��������>�8���;f�3>���|Dz{�2S��g�yF>����cPRD~ts��[>�m�� AluҘ'{w3k�y�� #h�Ӗ�wW#w8��G�4�g?u(  k^��2�*$~^t��A	�O�=	���f|Bk��8~c^8���h��}��G�6�-��S��������f�k��hv�	��P@�̀�

�
�p	�;��xM�\2�%��w����Z('�����W����/-�r�����q�l���<����:tH>��#���~V~�3��?�O�I�x�e٢
'J��w�t���jO��Ы����W%�EW7]�\Jڍ��(��33���I �\����%k�Zʲ���4���O�W�j�ܾ�N�8э-�����e���/yQ )�D�[����^��g�e�-�e��=r��!��c�4rnXĔ�wW����G�|_�{�{G�+p�תu��%�p]�ב������SB$�ML��K<�k�Z*K"3k2�θ�����������wgR�sfF=A�nhr��}M���@`'�,���H�B�X�m��n�M�T6�A<��%(B"����=�A���ϰ���n�Ƽh�۽�g��#�c1���JG������WJH�=~�\(��t�,�G$��J�&ɌKP̴Br�w��F_�4Zu	�5�P����7���lܗ_zA{�ay�]����4��hJ�7�$�����㦀.�M�6��1����K,��[�z &�r݂��l��n�q#�@�o��icJF.]��j��1L˰n;�2� 0�}iw����O~�Iټ�9|�e]��֛�yP��2	��@lC+%f����@k6iY�X�ŎA͉x��V�Y	�ȋ��k~+� `b�V�T�u,V6�|�+��s�<��MR ̂'�+���"f�~H�J+��Qix�9c�8�B'C1"H�����L���6X�ZP����?a͟���#��A�c��s�r`����~W{��/(�Oy�{k�,yS
J:�T���V��ho�C�dL(b�<���w\�;v쐷�z����/#�=�ݼW�P�$�ٙ�]�w�ޣ�="��=��7��:���27[oU*� �ȂI �\���]չ�R5	YF���+2vuB��u������ʩ����o�&���g`4v媵1-Ѭ���s��=���e݆�FGZ�+X�t�k��d6f���.u��u���Pp�[Ʊ�wܵufX��y������N� x�jua3�;x�J�ܨ��� P�G��\��َ��@��V4���.i�t����v{u�a��"&�q�0���	�ժƔj��lLMMwJ��f�	�<��B�z�֟�tf�3��@��Ѝ�D>�,=���,�q}79f�3���<U���N�׋�"F�~n��bE�}I��4����9@���I�n��x'D�I�e�=w˧~�gT�k�3���U�;��.#gϪBАt&+c�S�W%���˺H��*�O�G��+�8��	)L�HN����\C�L �,���u˚��S�l�z�ȑ���e�d���	9y�e��|��ec3{��'����r�d@V�7a#������/�(����EX� ������	@/�Z�hw�w���L1E�ɒv��$�1���86�pM�@IU (��N:�3��qM6���H ���x�T����,�d-��u��uZ��|���
X;����Er�f�20���M�6��@B�>K� ^8kˤ�ŋ�ll��u���Ӂs0 7k�Y��$rSy�9���b�_���i���#T��~e��#d4��{���\.R���$Pâa
B?�r�*��!D>##-�������w�� =)�:�	!��<~X��-�l��~샦��&%K�|�	���M��j�b� �Y0	 =����`���oT��m�HWk]A�nh%��M\ڰT��k�(��$��[W��Z�i1T ʇ :p�c������Ԅ,ZX�,�Z�e�d�9y晧;�@�^����N��*����u˴��女'^�_��\� p s������@?k�{�36 ���Sp]d8��(�x�{h|�A�j�s��Y� ga�c� U$e���h�.bf��ݍ��lx:�l�b��1�Q��ZC��w��Ļ�k����/�y@9@i���3���߽���zsZ�,9�1%����+rMN ��5��w`ߴ�7� 2��?�V���)$l�6vRj͒�'����S�WFj���I�K֟ ���*��~~�ay���ezr�>ǳ���{���q�r��������f��1���U����K9=|D�d�X������/ �rR�MM��"�0tg��X<)g�8�w8�,`X� K�g�Z�T�u�+�Z�ZE���a�Fs�Y�H��80�A��ܳ�C
�5ːA��^p�|o�����t�i�� B��7��ޞ'jq<���MA�-� o 1��Lq�I�Z�����j����4�P�`f9�C( ɫW/v�d &;�AQ��ǚ����ze�>�0��˖�i����X3zC��H�:ָC�H���*�����=�����5![�����z��A���w�L����^�Kj�˝?�/Q����7B�Y������y��	Y4�\r�^>s���l��j^y��Չq`x|z�����D�)4ᱜ�\���g�b�9U��?�g'"�ʬ>tJn۶Y�j��ߒ���;T)������ޓ_|Ir]ݺ�N�C �,���u�ٳ9�ޢ���K�D��ȥ+
 �$�rɎ([?�pL2�Y�)��J���*���믿.1��j}>���f5V+e;r"��:�m���B���F��f\�zL؀���%sybo�"�R�yв3+��\��L� i0��@���ذ|���c�8�IW����zZ�H�B9�z?p�33O���u*� �ġP�=0��p��v�ڇ�vw>�k�u�8������ȅ��PV ���AY�8*ޢ zP�c<\nv�-�`sܫ?��9�ԧۛ?t�3߀.w��X�^��>�f<_C:���BjE�M�[?r^��M}ޒ���jbvvN���LN���ԬT�g
s�~�=2g�e=�;��v��c'Ny5����>iá�
li�)�gd��>U�e��9z䄌^�Q�?0:zY-��=���Ҵ�Ѡ}j '�r�2>>��|�R²���q[\�V�Ѡbs���9 �\,�1�DJ]A ����?3+�����82�!�i��hHbu�^�3]ΰh��Ǐ����{v�!���W����o��C�27]� "��2N0Ľ��(�`IP;v�X���&^�QXڈ�C�ׄ�N:�U`��C�v��h��x���%llH~��W�s���J� ����}�(^X���qk�q���d�o��a��P��	ڬ]g;��[���h�Ӻ��h�Ǳ�˵�m]g�����8���m�!:H���7�r��ҕ햁�k`��+��Ɏ�hd=P�9Em�׿�5=~���|V�^��Z3����N�g9��K�ҔH<'�G&�̅Q	GZ��X�;A�}J"Ś>�����{ &�r݂ͩ\��Dcm���k-�[�����Xn�m���M?�0�W�$+O�N�z�aQ
rI��XK�[w���]ͱ����ҕ�KW�d߻�����B�,_��6�������+��YT�C,!O�	o��찣!�,���JΊ���`	CG�9��َ�aL�j�Ξ$1"q����A�!�;���;��(�C��f�,��Y�%�tw��5\Ӑ�)��񃃋�7��/��@�,U?˚����X5�蘝N�4��1�� ��i�3s�ʀ�h�!�d����sn�!��)s�ԴܵB�%nc�t�c��0z���<8��q���ǑL�䓟�Y��(H42�з��s�^��Q��T�m����e�e��,s<;|N����ӕ�+�t.u�����j�l��U��0�8��	��Rm5�<[�L_�D�Qi���r��@Y 	 =��T*�T˹�2�����BqI�Q*��ȓ�z�;�G/ti��s�[HDa��C�T����P"f%YjT��0����䴬_��xCr
��!K���/�H����J�����6�Utq�$V���������i�iX�pSC�@�z�0kq}��a�Ê��
��t�\� =X���C1������8�)y�q����6w7 �F� ���K������1y��G\|�H�ù�"�ݏk��s��O���a��v��o,Qc�8Z�.3�	��k���5�:y���%��(��9���AE�ʂ��V��!��N[�A���XStSK$��GV*|���W%��ސ������4ȍUP�xn�&��ң�ԣ?(o��WFF/˹3�e��e�d�bWb����O ��[A�O����)v�.W@�e�A=��� ��n�+dә�3�ې�%���[���0���A�R�V��!�]A�"�qs�[Fb$(	�Y�l�UK�Æ�k��%�)�~��������j�}d(�v�H` "�.k���u�<��F< ��qmX��֭7����5���NgtN��-
f9$
��jj����˗�0P�XP$�~��s��0Zl.v(���!Ο���zK>�я�� "ң��`�u�8d�� �˚arĳ8�m��p�N%�d5]*M$�a3�����ą��p!�qI���ԍy^�h'ގ�J̑�X�D:�&��>�m�x�1�9"����w���qryV-�[o���}zF������fe�@�*F�V�V/�t̂ıf�\�T��d3��Ǥ�ϾuDS�xJ�d�4]
\�,���u˪U�CCo�[۳t(��֒�J���`fk4�
�a#4�4A�Ym8K=���Ujã:���:g�����j����`���йb��X��gE��ڵKe��9sQ�ˎR��%M���p͆�ݑ� ����> a�l�v Q�	b(Cb^�a3����X�, �7�E�Y��mYq��v��A���	nP�m�fc�w�%��~��z~��Ap> ��8�F`I�3�[�BW7�#�,^�~�Z���O��԰�^c\*��%�,��pϜ7߷�'^���Um�{���)}�F���|Ýf�8󅇌P�5�NX�j�B��ǽ�U��~��P�,��[/�}��M�+���┈����Դ=U��jW�^��r�(�TZ>.}�CU�4W�T"ֹ.�@L@�F���\�Y7�J]-K�x�Y��N�PS��Z�V1f�E��9��`F7�dJ&\?��iG��wX^��ŦH7�e[7�yV�ɢ&1�Q"eԜ�p¨_C���9��n�F�ա^P� � DXd �T2�VڔY��B'���3g->����%-YԌǣV�����$�5pA�9;��X�M���d��|0Ƃ۟V0��p})�  �7�� � 7�ZБ�0f��p,�	/��Q���b�T�འ��·K�|�(�üp,� ��b�,a� �qM�ƽ��V�tz�3�Ŋ����z�K �Y]�����&պ�7(�/
J����z�����;%$@�jAff�d��.Y�t��]E*��SɈ�]5d�OM�u�2��Ų����A� T2 �@L@�e���̙3�7��x5\��rU�8aV9�t�	E�1-��率 ��ug]�3sŶ���$�T�c=ڹ"-3�ŵg�OZ��-
H|�ǒ��2��B�$��� Z�֙܅���HԕL�oқ21�L�0�ﱏ�e;{.j2��"�B��v&ޱ-*y�8��3� p�{�����hU�=&��7��:�o��1&N��QX�TzX����!�����(c����p�
���sp_�t����4�?G3���\���ʁp,n��=g>��17kL�J"�0�"��vr0z���亐����KT�k��E]���Ւ��-��/R�7/��.U W�m[7�E��l.-�RM��s@�y�e9�����n�z�jU*��` z �-�/g���tetS�d�R���[VPK%����mgmSW96p�� ���v#[�Y� �Jq�ڎ�zn#1N��z��)��x�3Ê�cl�}O��W~"1�?km˺w]RCF�	q����V7�d�g�QK`�`l�=��I�g��f�!9������~ǹ�r�^&=�pd�
/{�\ ���G�}f��� �X4���)�Y\�Dx=RŒ˝�e�/ۭ���4��qm�� i�㇄289t��x@Z�$B��u��bIjz߈W3D@>u��P�@����x|4�x
�~�f����b֫w��.�ԩaU.�w�݊�ő��Ziʺk;�s~6�1e+����*�1�&1������>�W�~�M)*r���w���e��2W�����+����G�=w�+?����/�O�xʊ�kC�H+ �@L@亥X,ER�T�O-�3�����Us��]�F/Yj�EK̚8�J�zu\���!���`�%y����*��D)�,n$v<<���+_1淙�q�t�*3֣��j4Z�N��t-��v��ؼ����� ׂbB>�|w���� p��e�Cخ���z�� l���I (A��`��2���{ B ��+����x n�nn��`=ΰ���lr·�K���'I�θ.�N��f��i��H�q{(P �*���k���/( ��c0�c1���rd�����7���μ+>܉�SP!p��)k���?xV
�eY�t�)��0i��-��&�W��;��j��'�Mo�_��_�W^���Z��ͽ�,��{�ҫ5d�8#7o�lI����<�l�֭����s��/�O��[1� �=�� ��n�����C!���+����e���f�z��7޼I��Y���g�����W_W�*Z��R�V�~�ӿ(?��Oe��jo�e
d�=���s�}G�5+�5���P���;V6�f�r�V��rAP�;6;�5f�')�y��ě�t��ʾ}���u��H�;o`�>W�b�l�t��i+/���! �!��X��'u,�������J���� jK�	 ����1�:��б�8K��v��gxc( �q=~���^8s4?/	k��r8Ix���S{�1�=�����{B9����k�ho:,�E�҅�����{��{���JM\�%����j�3`�[���c'U����qU̦�
O�<�29�$���y��`Ǯ��k��3�0y��q�o��Mij4aɗ������uڳo�l��Vy����#�dj|Bn�i�}��JQ�]	]��Ѓ;��3iߝ�@Y 	 =��d2Wi5�eP��*���ˊ��t3]-�LZAzE�ɉ��k�����c��o�����+[�_�.�jv��9y��~Av���3XT 0��hd5���XԬpl�O��GeŢ^9q|X~�w�oa/?5�<��s=c��$����LciΧeɱ�4-r ��`�� �8�bp/�غ�]��� �c�N[ ���*
��c�Q',s����p���>�_����c�s1uf�3V�1�;3��:������gd�cf>��4�9`ݙ��>�s� Y�2��<P�`i����K�<��t�������"U��\�=Kg�^T ��ҥ�e�h`�dHׯ�p�fl̰Kĵ�z��җ�$�/]U��s����'+���ŪX�����T�|/��$��o1V\��0nH5�Y�����[oEB�pL	d�$ �@�[6o^_z����sgOo���;���H���8��
�u�6��c�N�Z��N?%W���˳f���[2W(ɺ�N�=#���f�<�v��L���|�R����e���e߁��{��y�c�d)W��r�6��wm6��0�u��cΈk �\9�W�̚m��K�kرN)q	j̜F�z�r��-�^"[��o���s�#�@�Чk�����Z:\X� if��}�����z�{t�t�3[>�ՅC���Ħ,C��叐 �
P! �����A�2���Rgm|�����kal�&h���7�+w5��R��F�$��d^��?��P�^���?��*UѺ��vmr��Y9��Ay��7�g~$]����_��#W��g��w�yۈ�Ο9��MFVߴ�y �1����a�V>%��yX�'�,K��tue�:ל�I �\�tw�j,Z6u��C2>6�I�\�i�袑���~��t3����N6�\WFƧƍ;�Jv�@Ak
�`�X+�����P�cA�S;�r��x@֬^&c�#2v��Z��L^l�5� ���5-8)���5Ҙ��0f�ڷ��ڴ��=Ƒ�p |Yo�D9r��5�Ef=�ǵ��ǲ3�Ł�l��q��Y�նz�T�o���k��O��oMJ7<=M�Z��`,̃.��G��$��K���X�[�n�����
gy�sp?h$���]�䈂'c�䋷�i�\�l@X�Fk��[��H�?��6<���T)��� ���GZ�N�/xA���$4<�����/�?����o�������쏟U@�#�Z�ƭ�j&����{q���v/��Y�|H"H����rrj��g�=�츮3�]7�{;7�F	�"	0��)*��$K�xl�=~���qX�Z~kٖ���g��ئdi$R��D��)f� H� rn4�������>�oZ�������Ս{�N�:U<ߎߞ^L�xr��tO޳���;;2� Wv�Ҥ��>t����z���j�&�	��x4F��,��E���KƄ8Fˡf�9ڵ�-*�X�����&;�a���>'n�-��ժ� @�7��p��kf��5��,��[��+���غ��5�]�n]#�V�&S��F-w�8���!�Na8O���A|�st^R>�x`�i)�
����Ph�M٪��~��l��]!�d��k�1�th闞��1w!�a�Ԅ5\��y��/O= VX���h�^��F�5��Њ�_�@�A%�G�?��XV�4b��Xh��Y;�UuZ�B)�V��ޭX�����]TA�!�'�ꪫ��믧����I�Γ	jT����(��q,�)���mx�1(��ȱ��E]���ӳ�2�<��<�螼wA��l�59�cp��d��Ό
�$3tz�-[��������ر�6m�(�Y�^�T:ƖS��������MW���f#��z�$e�z����k�5����~_@�t$dcF����kif:'@�ۇ�S���T sӭ�-C�lD]�ڍL�M��n���vkC	���5��s��,�Q Q*U�i�jǾUI��y0��q����j�.-�R �)�q Xmo���>t�B��X���#[�����$:@�#_�.���0 =� ��ڹ��|��&XGx*�4��ֺ��£
�oB!�v�d<j���RIV���?WXټ�A+,�[�>�rQr>���K��'��z�z����r�f���L�N=Fo��:m����|/Y�J@�2��H"dn���0�y!�ȱ�۟|�I��s�'�Y<@��=K�5�D����ѩ[㱔�d4�$�1z��+��zg���ٙ�+�QWo��GOS���NjT7�'p���޷hF�.Z�����e����[ǥSm�I��t�ƍ�qf��:i͸a��X�����pw���u���n@�� U7�r�kM7,=��q�:{��v\�
��$�l���d�MO��E�x-'S�VU�c�ծ��ʃ���[�qf�B�� SF�T%[Qw�\&yK�T�?P� �x��
�%8� x���Pv�P�����<�E��"���j�� u�����ܺ���y�dZ�<B�}��s~���������K����QZ�fmy�%���G��W_I�V�.�H8�VRR�$�LM��i+�O W��b�Y�X<,��
����8LKV���l���42)=@�伋�,D�W����i��	?,�]���ͽC������a�F��蠴�P���o�Ca˔�'$IQ:;��]��x�����}�Du��mtv�t<����"KHL�3��fز{c����IQ�Wo���4mc����a�]��Uk���[mF4�q�P���PD�:Pjr���od5yc�gJ�b�^jg��+]��&V_m+[V�ܝ��K0w�mc���(]�ޏ��+Q��� ��)��! �€{("��Aܿ��	�-_. �,~��q.J�&�)�-,p(�k�����u���1.>�:+e�&���/Q���
`�A�>���k�40�^z�+E�D�b���a�S��٩i�^N��9@�|�)Z�|%�[��~��Z��"~{Bt���T<N��<e:;�����/�h���E>44H�:�9[����I���w$�p��O�B��'D<@�d!Ҋ%c9�g7+(�1qXbl�����[4;��x+ܬ�#g�M�P0�MN C<H�J�^|���������geC~��?���'h,����^�Ϲ��	 j��{�9�@��o�[tf�-6�V�l��Z�l�g䓤�&Z�������f�e]
2�"�����pS���䬹�5Z���n��/Y+D�R����r�2�i
 ��ĈkN	��-��ӆT��j�k.����a9�k7�,X #\���t��i|[�S/�z ��z@vІh�@�>��Hr�o�I[�n��"Ԯ33Yڽ��v��6�z($I�JA������4��C ��de�Z�����h��7���ҽ�vҎg_�Q~�P�����9~��i�+qGIMHHj^x�9*�<~��������4Y�SB�]�G�N��s��;����:z��؂������/�Y>��o�!Q
E�V�+]�䂈�,Hlˮ7햍R,��R�"�α9��%j�pHX�J����߅]c�Ȥ� (�z�7yX|C�Oѣ?z��A?=��W��I1O����*��
������G᱊�IF�j4:=C�X\2�� o3j�Hn"�4��k�c���Y��vѫ%��[c��Lp��ͯ��w�����q�Wk[����������V�ޏ֨+@]-_X�8O���ư���Ni1�[��^����HT������0��(q(k�J�It��@V:�͆w7o	�s�����~�~�Z�L=]��g�J�)��u���r����o��:����K#?>x��<,�h8&�yA�P�?$���ό����b _��O�Y~M�b3t�,{������K�K46q̪�k[�'D<@�dAbY���Ƃȏ�RF��8o�	ʱ���2o�
GRizjV6LI c���;ʖ|!�5��Ѱ��Z�:k7��8���]�k�� �t���M���S�?��M�>��*z��f�s7hB�S��e>a���!
p����!�!9��^��d���y`^Μ|.�»]�M��[��;�Õ�`�86��-g<\.r���:�^��G�:��c����_`㹼�����V��NXI�c@����O�<)nz-8#6����4�@��Q�B���k��-�/�s����+Vс��Ҟ�T]�A�'r�x�0gi��V�-��L�'�1'Ϣ�xhX��wn�R�N�3�دP�g��A��D_ B�/[*5ff�v`<���螼gA��/~����mi~b�-9��-�I���?�{<������H���2��EbQ
��4�5L]�`��b�,/Kf:\�J�����;�ŋz(7�ы7n�[Kb�ھs@�����{j�����Yz�������3��Z���luek��]ƥ%m�d8���s��Z��r��J�GRO���i�*	���1r *�l������ x���U���QW>��x� ���: NT9���2^���G�xd�����B ��B�%sZ[��z�6u�7`��z�������?��?��ق�,`n_���4xzHH~�s�;�7��L)%y�-}�l<�=BRԒ��܍ [�>��F�+�_����a�!2
	�l��l�=ݓ"�{� ፶:6lX��|�_~ИmT�yJ�['B�).d��`������~�wM,� Xy�Գ3S�J�*._�j'��st����@oZG�?����uwt
��.8��nQ�Sw�[��nP��A}�����D�7|t�oU��k,{�K^�кru��ziݺ��v��w CmO�� ����u���#�.e���z 0��q�ޝ��+^s"�M��pM�Nk�,?~T\��RJ��_\�Q����?<d��q���^
!�-���%p��hzf����@���H( rC!%Bu��	�f]�#]Y�q<�B�W
[�Q��a�kٖ��ū	���-�ϳ�=�0��'�&�ܦ9��Z`l�؜5+���U���ё�p$H�l��XWc�^;sIu�����~�H�*yc�J2[(d�˰�k�@.����ѹejnZ�SAq~�����2?��nV����3-�k�����:�f�k�7Ɋ�����w�����z}����4��@��
����RB��9�1�0��%p��X�;�k\������T��`�P���V���)u��tp �Ѩ͔;��j�Ůk����IƩ�@�q5!�P:-a�<#h{MR�L�/ �O�z�zMMN��1>Gk���8��y�@TC����-�鲓��)����L�=�+x��!+4�1�'�E<@�dA��x�j�Z$ �}��qq7e�E�v<�z��Q��VZj��~q�bS�K����F&2>K8�Ô�E�Ȥ�x� #�/��4�a�9Ǫ~��67Xji����;�>�>Lw�N�s��ݞw�:�Q�cw����Z��DE����2h)��(�d*nf6X� `XŚ������+ ~����������67;��/LD/|?Hr�g8n`�b��>�n��]�L�|�>�9���3�N5D�3a��$��;<�+����b��]�e\�e��Յ�j�,���{B�sߴy��v��)�͉҂k�w�(&�`@�Ϧ�<"I1*9"͆�tH2�C+@�|'�r���'D<@�dAm��l��cy��j6�9rzf3hԪmr�c���GM�n��ʹS2ѕ�L,S>�$&�%{@$|�v�V��*��d�(⿆�~��u�k�����M�+�1��&��=��ֺ��T�r��|ݱw�@�w�\��tl��ݵ��r3 $DK�4�� 8���b$ʽ��K2�V9�&���ذ�U����׬�]o�!�1g 5@<8��;���Lr7o��{�����6TF�:������Np���j�Iwp��Os*�
4���._-�P&�4������(q��N���[��[t�]wR'�KȘ/�����~�|����ZB���V-K�a*����ӆu�������4x�9q���G�(y
M+$�=� ��'��y<�%3؆����Rl��$���I��fK�� `	p$��	�RkH-6��B!GQ��P�c�2�V@S0М:y\6ydc��6��YA2��n��r�[M\�(c�O��p���D(J��kFy\q��mk�MI�d/'v�����9 ;����PK�ݓ\Ig܊��(��x
�����@�1w<'X� k��{d��up,q�1B�Tq=|�s����vxX�������2ڡM.����=39!c�^�R���������؈d�/Z�D�0$�A)@U���k�TE#]s��ŵ���@�z�n�kMK/���>Ip�|f��2��4�D��x>���r��������M�λ��GJ�!��3�Ӗ���K���L�T[88J�|�Wx�(��h���O<� ��'�x<ҪV�v��vG����/���EdږZ���e�	�g���|����3�L�PD����C(�u� �F�"���x��Q{�J�u� {�n  Rt���O���*��3���4��<u�]���0&�Jk�!p-�g�P+\-}=���v����w��ݮx��^7'{�E6�&�q�H�q4Y���`4+])d�Zԭ��mM���,�Q����X��K.�ca��z�߰�q�s��0�C�,s���,���܋6�Ar*5�O��m����)��ߚ����N:68$���/�g],�N:�t�ڴ�`�s�E~��>���mt��J~ ]�)���w�F�_�~�v���9�����������	:|�(����{O<� ��'�V �A�l�[�n�-b�_|�&���h��,�7��E;w�2&�.}�����������䯞�n���s����˷����/��\*�������ϔ�N	�⨠���۵�מ�vS�*�*��Xn��/�tl�j"j��ֵ�������J@�>��J�5�n���#.ۚS8 2g�uN�����-��9α�J��`	67�"���r��v e<C��1Z��↫���_�9IJs����o �_�b�(�j��rP�?)�w��W&:��4)�x"��mO
�i5�BC|��з��99��;ߕ���B�V��lV�PF�g�c���/�?)�	%<P���h�Y��A�S���#�r6U)�/:��a>�t��7�Z�����Z��/��1�ē �{� ��X����I�36c�C��� �%l� ᨻ�G6jl��b��K��n��B����u{�>-IQ?���骫�!X�����(�RQJܔM�:59J~_�V-_��\M�|�ʼQ���$9���Ic��uus+�i���M��jV�Nͺ�Y�r��AQ�h'v���^4�O���G)W�w�<����qw�^�^���(�ntSm�a��9����S�U�]?�KZy�amk�9La�C������5���$9���c�Q�ߩ����e֫�l��0xV�X":<Dp��r���������L����	������kBu�5�=�q� ��tQ��Y�m��&�������r�*
�T�w5��Wl����'r�A�/B�xr�tO$ͦe�b	�R.�E�%�/��2'�da����u9ot}}��>�����}T��2�Z�)� !��-��n�Q�E�ʧw��7�Dbh��I��)I�
��}�#��tvс�G蝽"��R�}AL�9"c���N�s���+k{U��1�]�U��i�� :�WEb~�qxMzS����$3w��\�v?ʥs���;���h��=�#��(pko۶M�e��4�������n�:)/�� /��R�;�'�������hֳ��2.,}m�J��xW�$b-�J���A��R�t�8���(^�`4A��;��f
&���x�9K�K�R�-� �C�a���-^�'J2ܡd��<x^}}'Ba�����ݬ��V���'� #$3!$��;o���o�m�*�Y�\� ݓ	��͛��t�-,�^��a���e&u��A��z�7]l��v~��IL�e����'>NI���zX	8xX����yz�՝�jE�o���:-lt�X������^�����c�l���6���o͹���l2F�u��O 6rX�Ƞךw|p�Cm�v�6ĝ� �n��s%X:77hk�u�˵�V�gp���G=�?��U 0k�U�'�ns(L \�  5~c������3��� ��3�)�T2���o$���E��Z����7@��\�Ƅ ����޴
\����AA�u�9���D�>���l�\)IIٙS�ZX샧OJ5F.g*��PRP��1��q�]�?@,JS㔈�BE�jI����(egr�l�z�?�!����磍ǨQmy�'D<@�dA ݒ>�h���l�+V����O(��.��X:j�cRZ���# 6_�j�h�ǿ7l�DO>�K:p`o�1��C�S���K�J����C��`�U�jՔ�a�6Y�a�r'�0l���]˭������p��dV+@��.+#��.?S0~7:wBZ���e�����q���6?��NxS׽*&�k�RWo����# ��Lq 4X�8 �yxV�w�3r3�c �\?�0W�<{X� JɌwZ�$�Y�#V����0��W����q8�y��F.��9���v�
�s�r笯v��:�_���-]B;_��՚��E������ɽ}���{�����۴%�~����-�z+~��)����Y�H�{��4��;�7B������=Y�0����_HH��dGB�>���E���$e9��>�~���Q�3��Ɇ��w���oڐ����@��<4|F�F� 0*f��lg��+���c��=*;��sx�� A�V(
�JR㶘�-��o~���&�[t��	)���/����C���'�q'ٹ���V��Ν,�Ob���;��Ϸ��U�����{`��!+��c�8��aA+'��7���N@�A�T(_�4�P��o\����@��q�FQ��:'\�Rg���5����j�q2�a���T��wJ -���z՛���AJ���z��<�W_}5����>�)�õ�$u���e�tl�v�x��n��?No��K��T"I3��R*�Q��sKRY1<:&1�tG'=q��oHP�<W�7��*U���'D<@��=����ַ:*�b nXXgEPGG�e������,��3/��-��"�Z.[�Ǐ���s�Y�[o��n��6����/~���j�9���������H���xR�����iJc�a�H0AccTak��V6q+�.wX�)_k�w�`���m���l�ŝ/������Wi��Ẹ�d*����8=���R�T���lɼ���Q,HG�3=�s�7L�O����δ����c��?'�u���f��U�	rj�l�|��`��'$ʊr���k�;���l������Z�6�s�kY�]�6���z���=59�&��b��z��s�d�c��3]�2晑�4�ϵ=��*N�ĖB;h����,���N�]k
c�(<�k������f��낎����f�S��ﯽ�F��?�S��x�f�F'&���G���?I��_��������3;��8_��K��\�c[�"���y,��^_�B<gԫ�2Ѓ'��s�W���ݓ"�{��f���>l�ب<"�;�������UKG�C���ܹS\����e��� C9�2�"Xr`��x-8Ņ=�/�b���N	(tvfd\d8���BI����]��t���B��*Ę�3�l6+��HrxnP,�޻W,vMDS�h�;�)��͚�zu���Ǹ��̍!���N��n:��R����Ķ��6�:�r���C�\��C����s�=�V� �>�G�߰v5�ڈ��Zh���%#��W����R
����;��d�>�t[k�����D9Ͳ��&@�\������������ ��$v�g����o�SgF�+�?@�~�v��Ř��]o�G}�.ٺ�&�'�P� D�b��<�Wӓ��||�G��7e� �A�`Gg�(��H�\A}��_�R���gG1GϏ��޽�'��G� ݓ�e�P(b�"
�l�a��U��&��ϻ�{��ɢ�����J`�g�D��[o�I������*>s�֭]#���7wQ0`��9����Ա�ϖ���7CG���I�U������~w_���&a�EpF��ƤZꎗ�o����BW�v��g�S W��5�Z�q'����1�S��h�ݝ��m�����
� ��ƪ����	�)�@p�����T2���	<mc���&��<m���h8�F��.z�'�h���'�	<W�����p��s�q�6+n���r�oL��1�����￁�%�Ʀf@u$�?����K�xTB'?{���l�*�� ����?i��-�;A��鬸��	�dg��g�;T�6)M���+�c�N$)��*6���������V@���o�"G�xr�tO"v0i��M�X��P���J�{��x;q���o�#��H(��
8�׾}t-o����K�=�B!�o���ǎP"�R���F�$�g�B���Q�Zb��$[�l�U˒��r�� ��N*Ζe,M��֮kJn�=Å7�����2 �`�%S�x�����-[]�u���u�縭}�g�پ�{\�[]��c�Z��r�Zu�+�� ��p�� \�P ��|6���9�=~�x�BV;�m޲E��:��0���u�:B��kz��0����dh}9�7�X�x�|-$�5�)1����_�?���%�/KW����1���:�U���������\�x�&90F��s]q�V��?�"�o�%t��7S�X��_w=����_�Eb)�6ge1��Uc˽L�`���j�:��⧞z�^}�5!�i�[t��W���:���k����'��G� ݓ
[���w�ɜ6]��?����;l� ?l�)���^@�7d���L��2iz��')�����7H�,7l��4\��o��=�3�<C�b�.�h@���<�L�K,8 �Of� ��)�&c��z( ���Ԓ(��0���/�;vP�A��c�,��>�-_�����_"7�N�v��K���%�?i'ƹ��t7������n�����:��������L�|���<q�>t��9��Kd=�}��π��w�b�gi��J���?�u �"ܢ�t�K���H��+h�[u*B��ׅo9O�O����>Mo��� z�����ޖ��Ԭ����-_�\2�7�_/�ƽ����ᓧ�c��7$����~O޻P8�xl��41:I/����h�R.�p��#�u�կ~E�7mB\�s�{r��tO$V˶��(~�٨; ���� [ݰ��Qc���62�Tҭ�R�$3$�Nl��S�[��gw�n���-i����$:9nrX����Xt������tl���^�~bÎ7�,ӄD����X?���~��d���z��;����?}�c�R�}��]�Jc��vw:D�q��ݖ�|�w��A4���L�`�Tu'�Iy��.��Ѷܱ M�����o<?� �(A^+ܫz/����7b舍cU���c,e����rWo�"�GV<�,t��5����{(!���h�H2#+l�~�M��;S�LW�d���Ft�� �yZ�d@�_�z]w�5������Oҥ�7�~��;���w�}�������M��>6[�u$��R
oD_w������1`M���Aj���.�'/�~94,/�ݓ�.�{�a#�e�A����l��jW5�����l�(�1IP���C������*�+Eʠ�4��ykՊ$$������F�#�
%����Z�b	e�����j�R�z�!��\�o2i ��/nx���PwV�%6�v�3�䭿����|P,�0�Vڧ?�i|(%���ص�<L[[�*�i\!�.��� ?��:�Lg��۞�ߖ-k)����f��ۖ�Rq��XWԃ�r&̀�{��d�#+����4��F��C�#I�({`�[�IF��P��>��Z����YMr#�d8|v��W���~IT��嶲��FQ�T�v���>G�2�� ���K���ҫ��q�ѐ�5�9���
}��	��S�I.ބ��x���3�Ҙ����(��,�Z�D	���-j��
��{��U���B��O�ɯZ�<ݓ �{� �D����S�K]�C�����.�o� |&�)�ۖl�l� Dl���5c�a�Hl.�2�=�|����S?�A`\ʫ*ee�Uo N����F�v�/u�Ţ)��,�KΔ����4q;�,��n:��nw��OUw:������t���w���Z��&��z�@�TM��Ys�ו}͝,��r�%����7ԝ\��! }�v��$�����2G���� ���t 2��Ф��]�ַP�R����#�9p�c^X��}`�}��E1)ԫ���ڤ:~W~Vh��7lZ��V��0�Cq��{�r퇎��bb��w�d�c,$���1��g>C�R��}�Yz�?��G�����VX���5^*5$�29���\lr-�����V�.z$y��y�=Y�؍�r@�Pwz<a���@��mAqC�ŝ��	J���w����Ӽ�"��zP�j[s�������~�tU2�W6�v'1�,�f�Wʕ�;�1�6�: �2�^�������Lk�Q6��lY��\����6;��jw���q�c\w���V��x���t�%w��1n>?����owM�����8E�Bwz�O��ɘ(_�k�~�u�ёC�h|dT���*W��x��wg:C'k��%��(?��-����`�Ń ���1� ��l��I����v�x*I$�2��I�3~o�H&'@��}����
��PpM_�F��޷����R�T�c��l��{�K�Yr(�x�����w�BRoD��� K��>���d�C��ɞ'�\ � ݓIö�z�f�B1�q��ٲ7+�έ6Ũ6:P`��'�)c��'��xv�7C�F��z�ħ�}A�Y
���P�a,v���0�6aY~c֚��nKh��EC�ܥ�$������h|^u�c���/w��ɚ�,l��|��Pv4���v����ݠ���d4=G�Y��k�_���7֫ƭ+_�g�����q�����1��{N���`��$�L��n��fn$"�Dr#�ݠ�������Q���`A@�Z,��^!�`��À[.�bRo:�n�1@:�a�xwR��ķ��XI���L7�Q��4=5f%�ԑI�.oՒ��kl�wuw�8p��=����Xq w{�\�$�|u�L��
A^r=0O<9���'���R���!7����}���)IkG:��T.P8�8�f�Z`Ǣ�.�Kq��5���y,��r״�%�cQܨ�G{�E��SY)MC\ܝX& 8��sk�۱m$X1h[Ow[S�����?pNL���ow-9D�j�B�s}~�2=F]��v'չ3��u�:�^s�<4y�+�%Y�<'D*�vނ����{�@�|�*��G�]��hkV -�"x��u����g����g�wDC+��&�i�U�P��Mm{��+x��)��w�F##�hyR� 
�W�_^�-e�C6:�N')_�:V|YB2�J�R�.fK;�'i!��h�����u$S��%,��oR~�D�8����C��[�x(��ݓ�.�{� A��0���,blܚHnll������]�VG�26�D2&�1�_o�+�����mh8I�Z���[�%�4�
yJ�z��^�����g�_Jq��Ξ��s#l�UP��v{��eMP""�X�}��:o�w���[જ &�2���݀�]zq'��q�ou��O�S�WEi~���bא�(.�D-m�<~k�=�c��Ki�w�u ��xR��-־�ϋ���r��qܕ�\C���Nvp�#����qڔ�����]8q�(���AS������0�ې��jh����u�˚
�R�I�����u�n��,Z�]U,jX�#M���Lͻ�ՠ5�.���Yi�����$��g�彃�������@�n���.�(�Yow+�&����^���+T��( *�:�������=Y���j7�u�L:�l�Lŏ0�9�݈m�h6d >�ovufL�3\؍:�QK8���M�>��\V � q\��?�E�z9{��|�gRs�ƅ��m�T66h�)%F��FX@�m>��l��p��~��,��:��M��]�� ���&�q'ɹ����Njj�+ kL��%N��j����YTA�,y��U+~c�5�A�m�Jp���P� ʰ�q���Ic.Hz����n 6��0&���y��a�לX�x���@֬]+�¿Q�ny��I��¬��	~��љ�'��L�m��I���+p��I�v�����h9b 1��L��/��/i�����=gF'�<HO>����}VK�v>��ϋE��O����~��Lx棿q7�Z�����������E/����=Y�X��]��_�he�R��5҄1Ul����X&�]�H��X(�� �e����0[Y-z�G?7l|��N�_q������	���G����a�x��ys���U��*V""U�[��ni��¬,ԃ���Y�M-^\O�˾_�&�n��0�e� =��|>K�f»]����It���	wj}k�\����
�x�3j��ŭ� ���M�W@�0�SY ɋ�R�M��od��,kX���f+XG�ˡ�ֿ���e�u�ȫ�q�\��� �7=�k�:&���X��r�\?��^���[��饗^��)�R��J�$ʀ��Q�����5�;{��1�S��]^���>��O���I:�o?+�Q���nv(*��C�v������^���d�o�d3��g�3}�o��Yy��J�<� ��'��ZMq�wuu�ҥ�9�28����O�GP��n�ի/�x�׿�u'��  %ݑa+g5jѥ�]N�_�Ԁ/_eڥ*�Z��f?[k1�R�$�P(G��x��m�$�����
kS�61�)�Rb���Z��AèH���%��rܼ�87�B����qwaS�\c��:7n/J�Ŗ�o�)���*�ZNC��q� W�� 8(Q�O�igػ�mt>�q�wƅ��5X� rĎq<,n ,�vHhp�*J�_ K^�-o�lz�
��"�e�[s\��`Wap��;��6�cĥ�Ư���ސ� x�Bb�X��h�ʕ��?o�?����?J�����{ĭ~�ݿA��즙�I�ꪫ(NPWw'���� M��Pb�.�zzx�B|��p==���;	��O<9���'��
�K�6nX] ���96cp[')��'>A���/�bG�2� �����K���M��J����J&���k�	�U�R&\���͛����=;��?��MP�aʻ*�9�32���[��ycGs<l,�p4�ve��F0�o��	L�Un;Ip�RQkZ��N-mu㪥�q�|��o�r�-�%>�g��R��)��
���s}`���0����n;JK�햇=k8 �R������R�Rn�:S$�� c�Q���$1�2��ʆ&Ժ	nP�Qg��B \-��IRc<�9��:�g�2nh���i�@�l��2<�D��[ͺ�c�R� ߑi�g�[�Z�d3� ޢl�H��v]y�մd��z������wR*�A=]�T���d���k��B�n����o�L�TLhi���)��^)V��(5ZU�VJ�5�>�9Q� )��}�֒�O,u��!�p�̰59=�Wh���'�U<@�d!b7m�lJ$���VTOO�l��6]�H(L��چ���su�!�Ѭ
{\�Ae�[o�U��O}�S�@��UT�M��瞕����V����F�����3����	 ��9�hN�~�`�R�ʀp���E?u%�y_�bԢ>� GK<�  ��IDAT=��qmP�F�l�RS<�S,�$9�$uHJ�ڞ�l���0����ĸ���>H���A(Xw��İG�8���2�^sb�e�Ȏ �-�jK�ꍒā}� ^�@3�Z] �r2��ՠ!��{�"�oD�&e}k�x�r�+�_:�Sp��W���M�X�~�~�l�Y����}vv��;@�|V�E���Z��A'�?����}�u̕�%�� G�p��Z��`L����9��B���CM��*+_>>���n���xԄ �x}��s7��9���UkR��
�w�������_A��=��WT�������1~���M��]���gE5b4���NӞ���K6Q�.)��sA�"(dA�l͓"�{��;�t*��W�6�U������a�
�L�/ܬ�ûڐ���7����=���{����젩�1� �R	��ݜ� ��kW��y��!���W,���P�"� ���Q���u&�,(�����~��1'�q�[�p�la�"˹R-�\� A\^Cڒ�=���9�����UMZ���9��4$`!9�_�SW���v�d��$R�K��"�����
�6*$��b�5kR'-�5����5����+�A�B��Ut�����}o��e�&$�BX�B&�ܬ�R���xOغ.UK��ĲG�"��%Ȓ*���*�k��2��uv�H"%�~�gg��093+��Cg%N[�H��;	�OZ�"�.��3�~nEz�'?�G�x�*��*�Mf�?��(d����~@�it�����*�����$�y�(e2ݴn�E4xj��ŢT:!����x��M�w�<�����,H�ʵ$93I�O�hP_�Lw����;�r�jZ�~��l�Y�o@n�P�_̠T��G��c�8~`�2�TK�|��8��� [�*�Xr=����٪l:|�!4�i��\
�vOO7%���Ǹ�m۶� n��7�`�~�t$%�Yb��S��u��p��w� E�a��L�����9�<�v���9�da����`$((M��ϭ�El]�~[��xHx��I.(���c+�I:�Yl��9�Eċ ��xxÀ/I�x؀5�J�k3虘|C,eH�Aߕj�O ��L+?�eu$�՜�@�Ȁ]��M��o��Cҡ�(o��IB	q�}N" bߨV0��d:#އw�?��c�o��ü�P��X�9���4���
+OexP���C�Z�y-]��:{R4:|�zR��G?B#�G��@�F����τ}��{������%:x���_�c���Z5
x�y�c'�K�?�` d� O<9���'�?dtәEm�nl�(K�bcE���kN�2꒑�5���5�V��J�ҩ����V��>����Ӳ��ࡇH��'��?��;^k��}��w__�x���tR.?� �-V�C?|���#t��a�o�<��G�1iǪ�+���!�p��b�E���$e��0�X���>�E �@[��)9+�ȴӴA�R��� ��O�Ib�;�qM*�y���* ��%#;(�{0�\�&�P�xL�G��4,��gD�
�p��B�놵О���.b�l�SJV���(Y�����A�
��Ʉ�7��nHKS�������2?o�+��C�}hfrBX٠�4$ҐrDQ�n~�Y(�ihx�����I�<*"P��OIr�����b���Ӱ"V�	@A���������+E-�&�|N8ar,��+��Y^s��;��5�5�]Օ7�fV@����d���J�^y�5�F���(�	^�'D<@�dA�MK��X�;)�h%2A�9���.δ ywO�d����nk�?σ��g� ��������/e�D����:,4dH��;z�.�h-��2�\�H�S�vE��?��?����H�WwO�l� �:�Кe��{���2�#Ng6�ڵ� �|�AS:x�3�W�-Na2�5_.V[Ў2p%ө�u����Ը0��c�Í/���MX$���b����(�k��
�d��{�x|��_��&י�^�ZE�%��
K�������a��x�I��1`a>� ,�BY,f 2~GCAq�7��E�8�Qϖ�l���Y��QP�*�nQQ��(.�PX��|�,?�'�������2"���`m��(�����@q�� ��{��G�y��"�k-MT�)���$�X�8q��a��I�P�n��6ck?ϊ[,��w���*��xm���-���*+;}�������ӿ?�4=����QX��-z���nk��� ݓ���l�M��!�`*%�E������JĿ�= �}_�:tċa9��ba�ݷ�m�����/�"���K��.���S�pj�k���G�!��0`L��ҙ���A���*��)s��7���q��7�.c�F�k�lP��<��	�v��-_7ܶRBf��/�����8,��5�P�p�K/�v�Ԁ�s�L���6>��U���dѷ,�&G�Y[��2T��J�ɢ�
p#d�j�%���+<��o���@K̀��X�-#�)����ߠX�p��u�6*��Kh4[Rڅ<dv�
 ^�BMc�W���M���d,.��OGKѺ��\Wa0���OA���s��̦=BH«�����ˠY!�@P��vc�)�;q�f��@�@[�5�!���7��Ò�8�~���9ާ�T7�����/��l�w���S�*�"rEI�C�_��1���6�4�	���[�#�߷D�(�����N���5���X�N�'��� ݓ���o$��b����]W6XÎ��͠=}fHb���S�nW���1��}��ߧ���tzp�z�A��<����s8�1&��d:DA9}F�P�[E]�Xuh��RWWMLOI��d@�V�����+�7k�u-��ף�.��Rⱶ��Cn�fk�&u�dW��X�H ֶ֬�5�9 #����:j�9&�f ���^Ӛ̥��t'�qh!Fl<�U�$Ð h�֭]N�|^,aű�I����|>Z����,[�߇�8�-�φ.�89(u�蒷z�
Q ��J�V���c�T�NH���U�i�����0e	I��H\��N;NO�x�,^��o��V�x �0 V�п��?!����w�y���A6����ij6Oo��G��Y�D�4��]�D!��5r�x|&��xX'������饗�W^��nZ�%�w���}+!VLg���o}��������0� �CJ� ��4�5�x�%�8��%K$qtl�N1�OL���c��OӒ�U�۳�ϯ���T$:�u\�����,D�[��T����HxJ"��V����X�϶K�P�������$�	a�N� Ha�D���AGeQ�"�D���6ܯ�XR��~
 �a6�wl�dhLSņ4��`���-0Ŏ����g���{�b���7�-7_�N΂�^è�f�lߡ#��C?�d�+V��̧idd����L-wgG7��w�~�Q*�%{�7�e�o���6�QlS��y>��������]�{��R�=������N:p��d��d�����~��l�'��X*�w�B|��]����|�v�m45��l!Oݝ��]2�A��/�Bg��h��e����1w�	�����~��z�@=[�o`�t���%�ɢEKx]2��_���x�q�)�|�et�%[�][�V��s�O�)U�MZy���'����.
�T��T���������z����+[��R&/���
�m�7%��4��M����/
D�P�(ItH������h2B1�������]R7/��HlTyν�cS�{�a)ml�ZR��X�5�m��XN#g�����y1tOοx���BD�Q�d�ޗMd ��q��NX���%�$�	Ԭ��E^��H�\K6�m:���J��o�V��E�M��X�am#�J&EQHD#�M`�=�a?���띛���6��T�7)��I����Ufe�%G��MMy��2P�tvI����>i����D���ʒ�'s�{D,���E��:;��l���'����mI�~5�@H����.�Ơ]�y�x8�mX/�6|v�v�B���<��������u[.Ƴ�t���s�Je[��*U��k�;��o�*Y3����� �����7⽛6m�~�p+'i��ި\ ��
�5��:���{�_V�QQ�&tf������GB���7wʽ���(4�z�-��L����h���W(W��~��Q��l�PQ �	�@#	��5���D(B>o5�	}�x��
ڰa�x�6�o����_��dJ��9 �F˰�S���ߑJK������JE���n�5Y/S����s�����K�"������oyIq�\ � ݓI��-�am!m�i ���A��On�m��4o���2ꏑM&2����}�h4�@��Z�Ir�naQ!3:������t���il�,=���t��i�z�վn��4з����ĂW�Y)�e�>���a�6UbЍ
[�h�a��7v�v{�-<+|]�	�|ߥ�腗_�Lk�S''s�n�f޸g���Sgi`�R,��Hi\���(g�8#Ih�P�V��d�5$���H�ҩ+=���9� ���._��g3�h��u�b�~��/I���-��7����X� �����ٻTz���b��`���Q�Ҡ��%t�M7Pg�b�_�L�)-X�"4:q�v��K�}�q�����Q �`�KQ�a�B�4�;xB�������M���| 3(|S�;�y����J�x�:�h�"Z�j����"�Q̗��^��IRgG�^����t�C�9��t������+.���I���� r(s(M�W ���V�0���n�X�G������v�C��͐�P�C~~���NG�p���Q� �`���+|r<@0�t�� �唒��x Ȫô螜� ݓ�4�j��ʆ�������ĔNUHUZs-D�Q
,\��*IWp���X`��r ^r�܋�[�s�Q`�(R�(�Y�Z��W,C���$^?:>&1r�b�$YIY�.�������3b�(1Ďa�J�)>�932� �mۯ���)��9�������GJ3�2:<�c��d�pI�:���Y&�O��L�Ū���c6K��6b�]�X�P��q.Z���G��Y���]D��S��|�I��|+m�t�(E�b-����AɮwP���^B7�q��<f\ұXT���&fi�P�m۶�o���Q��� @!�V(AC�9I:�x�t�o~J���a,⎾Juw��	]{���{?-�hQ� ��*���xv�b3��˷���={�h��RZ��W��ý���hl|�b���*+=C��;�g��7���x��{���zy��\��M�>Bq�;��=|-tM#?�fg����/ì���f��=_�R�#e�<%���v��(�UC�d[u�vG"$\�i�6n~[і��2�vx5��Oηx���BDʩ�������}׶P�":ݒ��vS�BMwS\�`��;��b�lZb��
A���?3�"nZ���
՛����* ���q�W�m @�4q<�8&�,�����5[b�5��&e�@���|f8���#l���;�u�}�EZ�b-��{@�}��	ڲe�Wud�,[q��l.O-u�i�ԉ��,���R�-R��c�gF��Xe��A9[�Ӂ��r��C���&�&h���⎶�0�s�(Y�M����^�����*e*7��R��h���.�s����jVxjG��3�K�P��{�շ��]��$-_���}��5J<��?8<E���k499.�y���4t�5^���6m��m?:v\�+3S��� ��L6G����LO?���C�����*%>n�	ڻ�8�H<+��Kv�B��.	q��!��"pP�9�=j:�����W�����m��D��M�-p�Zo�I"%�:�@AM��0����	�
S�\�$Z�N�Q<ȊYW��;+�@� �f�&<QB��D0�NZ���'��o� ݓ��g��Δ�n����:,r����o$}و�Z��Q��>Ir��!96r�p�"!���b�(7�����,�T`++� Q>'�B�a�Ih��oI$�ʀ �+��P{��]��v;�jސQC���&}�[ߧo~��R�� p SY�&[�/�~���F{o��CE���I�<�����[c+k���aV ����M* ؎��dgs|�M�d-��=��E\8P��w�ƍ45��&"�&�RZ��赝oK���̔t��fe=���M˓�������$�	 9��`��c��� ��/��=��<߂d�/XD����?"��X	�Ύ�_�՗Yiu�(cKf:��@���V��s�Q��.J�%��X_(���3�TG���ɱ$��P@�c�N�:.JO�&�汖�7������G�֏�r9 Xk���^�΂�/B�8�;�4�U�9)}û��H8 ��+H���ˬd��=6x�0��~	Ws��G<N|���n_����,tOοx���{ް����?�B~ِK� �r��q@m��n	%(���GW.Բ��j&;k��1��K�M_�٬ś;���9J ��IM�Q��C|����m��_Z~�$�:��Ki���g�Rt\�A�W�Y���o�C���a�ǣf�n��ub��)[�9Ðǿ�d0� ��)a���m]�P�5*�*_.2�aE�������<F��TKb�I[XP�JO񀔕��	}��DCq�r�3X�ed$�	���M�V�������oG/om�j� �¶�Jf�P�>����cJ�Y!㼯�O�p;zB����4+E�V�����h4Ӵx� e�]tj�c�j�-�[�/�[C��"�e.��&�{���X���(n~��-�0x�a�<�O/�m:Xxe���>?Ŗs�-� ���P��� [ՠ�Y���GP�`2;A�**�]Р���F�m�T"Tx����9r��7�J[M�� ���y���=Y�����e#V]��*b��>@ +4�.�.Pd��	9��d%��A �q!$95�í�,p��[�$���rڜ����04� |K���E�u��v81	�8;���e%V���f�bC	Iwt�Uh�ƀ
614A�	_�[ZH����q�g��cB��x;��Z�����f�:"E,6Kñ��'�4 �������=B��kBꂸ|�^��fx�P�7>>%J�]/P,hQ�3-JN�R�{I�|C��w�-�nV��T�{$ �d�4幦I��;���k�/:�<��% ^����Л�� 7tzX��e�Iq/�k��xԴ�55�
fB43��ǎSO_/�-�b���6k@yj͂�e��P��Kaq�L����c4f7e]/꣭[�ʸR����w���X��R��� 㽒,}V�p�a�+S[�P
5����˚uk�ڛn��E�t��!�?�]��|M���O���		�ds���4�3�~�n���҇�=�߷�y�FώЩ�hz���v�Z��xr��tO$��ecsGb�:�2��c�Yp?k����l����'ܲ���!i'z�-��%�]N�>���曒T�:k0|�s۾�(�����=�w	� P�[ ��+��:�u6)
\�����S!��c����â`���B 1��N�ak�?�!������͖(@����&w:�I:�q�Mt�e��q�uJ��70���7hY�Zg4֦�d9��-	[�=E�*��p=�i�=�3$�	9N,-n�D,$D=�Y�Ig��T"��ǖe�ǃ�˿T4�x�^��lљkQ�/ ���$e=�`����#^C�1�����Icl5�T�g�So��$���u��2�t����g�}V����NnE��J�k	Ӟӊ9�rA����'����k�<C�$������ eY���[d>��iZ��'L{������Ŭxy������_#��fJ�P
���#s����ipp�~�� �ށ��tO.�x��ɂ6w��$���]+\�(W�����A���+�ӏB,�Z�.1(k��&���mt�w��eK�o���t��
D��[��=��|k�~i��@Y��ua}C�ݏ����(;���  ��/��V�	�ڭWI�b��_�fǣNU���E�fM���F]2���k���,��w8�Bְ��LM��@B�I���gB�Z�6�R�\(�6����.|�!���4�A��>�O�� H�H��ff�R�NFTD6`��S�dZ���a~���ʸu^d�Ǔ&�)`�$���5זi�L9"r�����fg(�Vw��)K�qAUx����e���Nw�4���@��M9W��F�(�I��4��H�zbt���;�g�jt�{����R3��`�RM��6�ox�pj͡���g��N�:a\󁠄�χ�<������zϿ�,�~���gO=M��w��\4�h�Ӣ��V�uW]I��<�,���~��.ɵ�A�kECԝ��y;}��oS��Eq�<����螼ga��|�A��?���������f�Iw�����/���/����/�Y��K�A��;b����D�:{���+�o�r�^�p�r9q�6���Y@|���j�[׀��Wu]>W�O�L�o�#�*=�� W��!Ӎ�n+��$�_��S�־�`��ҟ�ghf�	��� $�"�|�9�8`]k������0�|�
AI�d3�s /@�j���(,>IPl:�{�X樕����kbj�]5���us�c�l�2Y;X�Rg�{�g `�����J�ibr��#L��E2Z�J�Vt����.��l��&-�5Se
 �/I�ȑ�2���ER^���u����yxo��!� ��+n�싵	QFFƄ(k����!���r�B�H7�r;���������]�����A!�e��L��ヴa�
�9OA����K��י��Bގy���=yς����߸Q٪�w@@nw���o���_��-^F۷o�{ｗ���-V$ -������k��C?|�>񛟢���ߦ�L���ڵK@ɸӧ����Xx� ƄW�l�#�x�b��Jk�tZ H�\�#���k'���i��.h��ڊ�[�*���N�U!и�f�kl߰�ڮy <�	ֳV �&��7� zb=�
.��S+pZ��x0S�0�ឧf�t���3z}�
A�259.k�~|��C�����N���4}�Z 8*,ħ�-[�o:ΓX�H!׵��F�(�P�O��));V�ʕ+����xA�M0��N���������������G��s�o�xh����ҾE����>����˶m�C��Ν;�}E�/�k�v4�)I�˖,�5@�}2��	4��Aa-��7��}��ݓ �{��C���V6����a#�k4���X��+<ѭ��J��կ��Ĵ��ٳg;5(�/���/�w�A}=������.�x*���: 5��t�M��#����5�3����eLP4P�t��	z��]���j���Q�&�X��}�ڏ9�:�7�]�:F��8��5Oc����
�5�e�X�o��gpC�yX��N���R�  �g�tq/��(��k�R %��Đ�L;�UxFXWxF$��
@k��c� ����7:��k�-gg=��M���J�wY)sD�A4�����hy*�#G���W��k�,���IRc�6��?;�ա��3�s�h }�}�Q:��2A+hюgw���9+����q�g�ht�,m~�v��L�00��ė/a�P{i�eЛ=��Y�\� ݓ�,�п��6�� $|a��\� �K���.
��ђqOԉ?���Էh� 	2����[�}��t�B�����{�ivUg��|9�W��CuUwW�V��d���A����g�xl<`{�ƾw��0�x�����aB"��$�Z�
չ�+���|���O}�g����;�Q=]��s���h�+��]R��b���z�Fk��9`.(m��>H���c�y��	�6e�mن��2��@n���S�!h�3�!e �	a�5��&����aޘ�%��|1es�������vC�z}�d@�+�<^F���r�K�`����35R)�p.Ȁ1n�lg��NiK�d�T&˝���w�H�z� ��N�����:j�1xہUc�h;�_��╷����������Ӳ����d�k�����g���υ][��	���ɤ)|�0?�P�ݪ�^⽈�����߰a=o4g����%;=#���}2?�(�V��@��sIF�+�����{����::�et�vt|��%���eZ��Wn���5����3��X���p��>08�1@=��0�8!3
E������{�Z�܅�c�N���?�0=���}����#��!�sutu!�l��!P�Ϲ�\[k̜8d]m�R_����+X��c���y]� $�P'd�c�=ݖ~��vX��Ƅ}s��3�l
s�������;�0��E�Qd�8&T�}��m�b�0n��;��^�{�DR�mi�k�W1���G�.y���3���zB�&�o�?�0x���"�Z]P�=����aj#�
R�xsoz +b#�� -rq��
�q֭�x	��X<�xa���0jTa�]gg�g$��"�N�<!}}x�y����l\�ޤ+IP�`���ɟ<dJ��g�׶��?^*G.�M(��Я��j���r��.�Q�?v�8'
;���?~�t���	�5��%��|�+�xq�����f9t�|��?����}�a`�{��ˮ��
p�micNql��G����l�>,��ηRdz�l	=6�J�� ����mw3 ���-	?H	 ��}�х�3�,���?5�0�+�������jߵ��\pM�M�I�0�Ӝ~���'Z��$�">��Qv���y'��</�4��<���`XT� �׍V�����ǽ� �ix�s3���z��'�FMؼQ� �f������<@��F8d��T4^���M�ٲ6��x.\p�4x�h�{��E#X3|]�rz~*�5@ ,�x��G$�c�=�o(�e��#$��ڱ��@����*��!yp��p|te[\\����r��)��Жa����y�W�����u���(4�;{q������9������߬�fʦ� ���n����	�۽m����5�e�/6�/~���i�"�:� v��Q��-�$�~���o|��:��|�ӟ�������$���E6b/uI�%�9bs�!cJ���h�g87�k�殓�6��>6�%W��W��nگ�{���}ZAk���\`� x��7>g۬�
t��9-�����6��|{���V��FL,٭��a
�==}�t�1�u ��Jh�Ӝ�=�MO`�@8! [����(pA��À�����Z)	�k��8��{��[R�]/�;ɖa�����rǵY���À�����} y\�];�4���ݻ�u�S[]�	�)&|W�Y9��)�4r��0����(�HXz�����^#N���	���%5lv��'��_���iӠ���g"u�3��K/ȗ��^S�TV��t�>����������/�+蚃�t^7A F�T��L2�Qo0ɲ3l����w�#��{��06G�\�HＫ!��n��>�����g�zZFGG	L�b���`hГts������f�]Xs�z� 8z�(�� �0l���uR7��X̓�\;��ܻl%��<���[eJIs����es���|0b0OC��������kU�Tf� ���Bu��R��x� x#`�׍@�j���V�M\p���1��C׸y����>iZ��L޼R,N���iң�E��$	".�r)��F 캶�ز@�C��z���1��߃glט|�� �S,���<��јǎrm����Ǜ���p�x���#�BE�Q�6��ܴ��Zu^KM��ر��x2��3�����|��ߦ�8h�/�|0���e���5�	7L���At-�w� �|E&&��3'�� joh���b�g�Q6���:�!ǆ�p��܂LOM�ۇ�9�VG] C�2�������tx���<�-ke��:��>�|ȓzD8iɁ������쿭 o��\����zs��{k9�@ �3��}����i>�q�YG?xi1FZH}����P2��m^����6�����QA��C�Z� =v���n߹CN�8A�#"%D�50�E��y�X�0�.f*\�W� p<�"����n>�2�b?s�1$�5�r�:cȔ�mܰ�9���E�a�mw�����E%=���>�y��R�4_Q�(����_:z\�(�wttR)�H0�9@�#�m߹�]����S|���?����k�I5�R2���]"_]f^wllB^|������P4���
.;;ȿ�����*�G�IR��W�ZB�r�����!O%Mr���l��Jb#��m� ����7�R��9ZP�h�� �?U��Z_ޚ;�<$�
�֋��1�\�<o��wO���sm��[ ��Pxw��5<��WFH$��)��a}�����Ĕ��&vfχ(�A>���W6��مE�o�r˭o�?��)��Xo4���T?�VhZ�=@!�@0��놐<E]rYz֔qEY��M��Ƴa�+�l5�6E`(�����~�tQ�\({5�5Gn�|
{ �!; ybc~xs�v>��ǮSt'F�F�(���S�z�_��:�BI�l��p(�ү��y���Ɓ��ö�͆�u�Ú� OKr�zD �:���拍5�R8^�8r�)��q�&u�-�Hm]��F�gpp�:��S,��9 �5�iyJ���8������& �	�r�[s��m��
q����t6��V������� ��+�c��Y{Ŝ�b�	b�1s0�qХ�������n]�^�nT��L�z�p�NQN�>%�
�{��ǎH�jJ���6�5�|��JL4���������1xp/m�����8��]��;v�/��<�4��Wܦ#0�\��+Ȁo���)����@���oH�-7�D9Ԣ3�є��
� o���[B�~2�LQ��V����wn��sj���@�{WO/#�B����?����k!'�0�� s�dY�W��h6�.�/��ޘ�U���\��+��tK���18$9	vj8@j�J �8�$�D"*���-oy��f ���m�6��qL+ b���:}V���P��g]e�=v��َs%�]뫱�_�	�j�3�����|��[V�5k|���h%��i��"���w|�z���6�fЄ��=@�8���� �h�
�7>���)�֯���Wy����������iI�Z^u�����%N��i>h�kk82��{?�W�,Z�_�!Sv@x�~Ȫ��%���/��U	�׆띛ZKn����U�3Vp��iOp�G�����]��Vi��mV��!��n�,���@��n�^`×x*��D6_��06�����������Woe��J6S/<�S@2�%Xh�j��:7W��ꮧ4^Y4��K�� ��Lp1yjS�ddP�(�߿� m;o�5l�8� /�5���Ы�Q��;K�_-�����o�{�1l��z��k�߷[`�u��}���w�!�f+�{s[tx��l� =�%Z!`��M�=�<�{�� ��������]�D����3�r���y�69��1����<y�J�x�0L=��7�:�����չ�_Y)��j��Xl�2��
%�ݻw�z��5pıQ�������f�ƨyHנ��,|]K���:s�1� h�V1q(�z��x�L5�*���0\+jk<����m,�l�z�g�ډ���>��cMC7gݭ�£D9@�u��3�Q���Cx����dK���C� =��2���ʫͲ�uu� �`�W�0��?�yp��L�>�.����f���JM�א��̓Qo����/���][��6
a�gA܂j븜�g�G/��Uw޶<�R�_����u�w��t��G�&5�!�b�l` a��7ld�uY�ԕ쒜�x�Z �������D���IG@��Ȉ��,�T)@2V��t2�&�AKT0�	kzOY�\�~�6��½Fh��V �ad��?7`�g� ��#S*�=��#* �:��q��,�Q `1p[��k�0ܚ-y��d���xbX��qVv�\c�wt�K��KO_�	��S�C�����t�i�h�٨6M[O�#6�8��	B�W��]IR+���l,�`]o��0V,M����L̇�z�Qg��I=�ɕڍ`i�U/�j7mK��@ F1}�����l[[���0E�R5,h�G���^8F+��z���j��-�֠�����A͋(X�=�����A턬Gj<CޓP�A
��Q�hHtpTx�t:�y�K�=P���vD)���X�K��dh`�l��KR耇y���L�X�ujAO0�Q��[�'����Л����ܚ�<K� :oysH�bݠ�?48`*�\�i���U.Ŀ����b^网�̡gB����������1xL�]�|�n����V�9�ZC��
<;���A��B~^�=�k��>�lA��xȏ����1|@�ǚF �4�ɄQ�S)�ь�b!���b#��GISڰڳy�o�ES3B[Q��H4.����yE�˦[�-v��Q#���	�k��~�.=2�{��{��
���?��8���;����jq�~�VUaf��~mKU*��0�5� ���[�q^.�	z^�G~s^#z�����j�����D�Zq˿ԃt빥`t�f" 5��@����͕�C�RH����\՟w\�:!�eOB>1ak]ܛ�z�}�zyO� W�mfc\�]���-�s�Q���ԉ?<b����`}�j�\��5���B�q526����̜�-,Ɇ�Q�9kz�"�jl�a{�:�R���%Ϋ����Z�+:�tR����D�R ǳ�g�?}�T+�܌aA�dIH5x*%}�t�Q��.���ݿS�_�K6oޤ������3���_8)S#g$V#�Ts��Z ����s>��cM#��y0h���y���(��p������;�M���F7�����4D���_�u�����W��U��׿n�����������O�g�y�D,[�mۋ�C�Q�����o ;@�^l����f�0����䲰�;^7�R,����^QO�aIq���a�p�;���g�W�Wx���[���|ù�=["�Ӥ�!۽5�/-��@YԫC(�
�~�.1ԨL�ƚ"%1�i���*9z�;��V��^DUCI�4�W����+����E��C�K�(���֩
�0h��k������A1H����z��(W�sn�,]S���Y��H�d�8����C�F���TP
��L%ش��0�pm�@C6�둷���nC��_����i���~���}���H��?�+�5^w0�rR��r��>��cM#��	5v�d�!͛o�Y2�mfSv�}b�7x��y��g�ȑcܘ.M+���	���������n���У37��׾�� 
]��G� �06�����9�R��gIT���Qǎ�;�+�-�aZ|�q�z�y��y�A 7Xj��xy�&r�n����elm7�l^k�^|�-Ys\�<~��ф�i���[
�0�u£{\�0�Wn�1�v7���Z�����G�{��mrס�ð3�g`�z������@�.;��`�u��o �ϭyv;_��x��������$H+!d�;�u��/c����)׈p���V`�9lr�7n O�P*�ё���LMLJEA������L�kt4� ��q�M�9!E��2�gG����&���zi��ezfN��l�]ۮ���v�A�+�w�-�r]�z�yY��v���?~�t�i�B �����፾������6n�$�d�\��������>�zw�c�8C�P�;~����~@���:��c�tS�d&��������?N-�M�9",<5=aj˗W��i�x�9|o��-��mA�P��ح�������|��J#�vyk��Jt6��J�kU#�{�[�|���i�h�?q�ٮ����}�،7MϠA�Y0"��C��:�A27�[���˖-ò���r��Y�:C�`���P�s`�m�'J��.���nkV����`���6u�˙�V�"hz�AY��)5y��@�Q�L����RA��#b���z{Q;T���U#k��B��k�uިFNJ�����h�����^��ލ�g���Y��I{w��~�����2��FB�-��9�?�q���XӨ�kRU��-�bY��ݢ������m�2�A��B����t�b77�?������%�zs���	����Q������W
� �'�x�" a�{ʪ��j�PR��6��4*a��~����K�����5�L.N�<L�"73=I0@�S,���^���P�*��Pu�-J]vÐ��ϴ`;AeOػM=�)hx?�����������7j�W�7]�Ԧ4\�3��n:��n� ����3/�m-����e��	i]�#��W;>!A=č7� �>KP���֭[e�SgϞ�rY��|�5��F��l�A���|,Siz�n74��ѿ<$��ݿ����x���nx�(���=����W���СC$G6�$��'@�=��hRv��*��.9v�%�d��yۡ����)i��������28�U��y�#�n��m�d|bYzz@�t��a�:�MΜEd���,�{�?���*�i�YZZ�k�����u���76X4��|��%W�����[o�E�/O>��ttu�{���?���4ù�f���~&��47_��` �v��0(OPT�Æ�o�>���[��36�q��͍�B�8�?��?�0���)�3^#��@�͛Ӌl^V6vY}:�e�l[�e�f���*��Ps�d���r&��i�_��1,n5��HC��Q�4�d����!!�c[[�s�[�~��q���kj�D���/���{�����c4�Ф�(�x��s'��19����G	�b�6*�9�o��=���a�<��u����?ał�G��Q��s�ѐ������f��O����L�1l��F�͸>����vٹc�������7dvz\����ר��K>�G�B�!CD����v�^��u���������XR	Rc�V��m�*z��?�qŇ��X��<�фzT��é7O�	��m�)��P���
�䱟=idV�Q�Q/�����Z��M��}�ѻϴ���\N�]B�W-W��3#o����K��l���m[=��Wu˓l.�O��T���H� ����I��`��h��J�Z����D�4���nU?�^3�I�a�2��y�4�m��j�5����i���+U� ���e.h�a@H�Gd�9q���V�ݜ�R,Q�ϰ�������F����ر#Kܣ��vr(��.I,l���&_�	���ȱ7A'��8��ޖdffNv��ӝ'�[O$LDP���E�[(`��T�&Ԧ�N
p���Wըsy�cM�+G����|����Ї>${wl�'��̙3��kT�C�~��i�O�T�����s�d��k����z��e�����%ԈH![FEA3oT#��+E��+0|@�ǚ�eq7ݖ�`�:u�`�\66��۷��8�4v��Լf#�l���U�|�m���N���۽[������mn� l��cQSS�? >�����\<�v�qwYAɖC�Z�2�Ǧ�6�PC�w�kY�_2��՚'�r9�[��V��)Y�-k�ܽ�W�L`w��cY��\.��lNٜ��*��W��nj�];��!��
�Ș ���f��A6�]ط��^+��_|���ad��7���.z� �h��h/�ʔ[EC�9֤TA�yUBј�f���z�Z�/j���| !l���ٹs'C� ��8}}��F��&����g==���ɋ��X�Q�(��u��۽{��+E��C������NF�%]���y�'���C���^�,�[����r%/�Z�O��d2-�@��,^�}�?�����?�4���(���2�6-����	��D591-�z���w�U��G� �4\�`C^sÍ�u�������%~��������^��o=��fmw2x���m�/-,�[��}i$G@�.-3o�a�8o z{{� ]��Mb%쎕JJ�\"�"��d�bg�l�6��k ���uh��fϚlg�u˔� b �{8��F�5�V|�|�=����eu�	�SBTA�ꖙ����/5(��M��K6�g̞��XHz�*���0�^g�<�&5���뱣w:J����G~bjR��h�����hY�4�P��t0`*�X�X^Z��~*e5j���:�+2>>���߿��b0̬qo{A�- ��O>��fg�=C	�ǵ�^-�Ϟ��+�}Aԃ�	��J��{�����>" f��c��@U����YC���%��Y�����ַ�%i��%��:������y�z�U�4˲}ې�בpD�U�)Sc�r��qpN(�V*���:���?c���5تn��Ŧ51����/���'HX#�;veD����􅍶��\,���9i�2`�:�B>'���7��e����bk�0���'+~G� �f ���>� �s/^"�b��RO0�{4���<���q�QR��g/��Q.;�z�Lڀ=��^����[�4 c$�`�Cݭ�̴6di���a=�ְ�%��0~���0���|<kݝ�[Oo�������_z�`��ॻ5�
�T�����W�i"��Aq�Z]�X$J�iE��p���>����4,t����[���5��&��6���^��H�E�d��FX҈9A��;�6���3��Q��x�0��F,�|Au^�1��hg��;?}�a�Q�:	HBAǕ�I	�ejrF��ѹ�lz���}{�Q�Mm2�Ve�sU�����^�ׁ��
>��W|���5�f3�膉�8�^��Jy�$��t��;︋-9��x� �?���N3�y���|�m���m�߆G�[\��y����҂�)B�O��S�oW�KGw+�P�T��f�)�T�b!1���n����nV�4A��tIC䉋���aj�Zo7�Z[m���j����5Ք8%O�����g[��Ȑ��mLm|Е���$��rͭe�w*��]mTV��� ��b��D��-,����NO����Q�,+s� c�ܨ�,B���S�-`t�BbY�UH0�p�q5��~A�!� wWW���N0�uvu2T��	��!.�HH{g�YI�c}�Wx?a H�h�-C�������{CC�^t����/�Vs���D�=��ޣ?9��s���_j�1�E����>��Fd���n��ߏ����3r�u��dzvJ.����Ã���6s������>����������?���?�4�ߐh8ބwo{~~Q^z�l�&/�|Z������������x@^>u�~iR4�����g�������u�6��|�	��*r�7�FO�Q4���Z $�1S���=wA���0o�>�cs��q��V,�x0�OY>��z�+�᭛s �1�o��G)H}x=d��(�A:���0*�M�S6��a�ݩ#�J�yP���V_j[ƅ�wȕg5LzSgA;R� .s��1�7�=_w�ǫ�0����QO�p� 8��W�O����.�W��*��Y�g:�y�{ט��C4em:��Z�D]x�������4�:4�����=������-2�e:��KGx�\�ɜ>W�r�Ү�x��z��½2�@
c�뮣�����3�=�J��h���:�����j��Ǳ�:����"��a-��ߦ��3��]ݡ�ۙӣ�˖dpk�l�H ?r�y�_�#�5��=��lX�E�iR&g&�S�=�����k���u�o h�	�g:ɬ>y��I�p~T7�i�h��^^ʚf0��I�݅�~�(�?+�>L��h˨Wm�� ��vd�l������Q��ق|���'�m
�������Axmذ�ǄW_(�G����e1=^�^<�B�@�,p��ԃ�!�����6<�&<s��m)
�n�æD-�^(s�M�öyy��r�g��I�O���:��,���o�w$cd@��%ṃ���m���0=�Æ�1 �Ss[�6ٳ\�?�� <�'�=t�ۉ!̭d��Z*r�;�h�[Tp���}�i+�ݻ��gfv���ɗOH�����Ay�-�@����Q�6���I{DȡɟlKJ�z� �Af^=�EgDe�۵g?�?�{ ���s��2�Sn��mN��> +���`�ےQ���k/�L'7��ժ56�!���Iy�N����%i?}RbI��'�ʲ�}@6nآ����25��J��T����?����k�H�V�V ���7e�4�Q���Ar��	��B��+�B$/�8
 ��0�I�8�*ä�2O	d<|ozӛ�����f:��z�h�^��Rf�D؁9���@��V�6dfnV7�(ôd�Cs�bZ��s��xn��>@ǲ�추̦�n�u�6�nAyi���0��$2�P��W���@�|B����.<o�q�6o;�!2`Z�<� �iy���Ca��r��]��&��{i�	b>�J!���}�5L���65A�$���7��55��248�X;��6�z_��h������EN�>+�7�~��\�(%]�;�Cv��%����(�204�u���&�g�ѨŔ>�Q��s4� �8��A�\+��>�N(�C��FF�"%�۰�k5#��`ra}¼w5�*��
��-�|���{�4�D����%Y��Q�!ېD<%�|I��e��I��$[\���E?��+>|@�ǚ�n�
�&6��zO����+����I�� �rC��;'ы�%���	`Bn�eL
d�j�9g�<!�[��� ��52��������p�zR/��^w���h�ɼy�j��MI���<?�<�9e���a#XLE<�ƿ	�֗����K>�#+�
8+�
�5�h�c�{-P]�a�۴M_���껣�1="^�@������_�9ã��gaLDlq=�e�h��LM;^�@��Ԯ~��g�%[�aqK�(K��D�U_��u���� �d<f�T�}�(�r��E��a�᜷�y� ,���=�Q ���^�����E�٣�>*�Ϝ��}����,�4�A��1^������+�ë��Few���xݬtp��&2�;Gξ���Q��쐅��������Uc�rÅ��W�@_BN�HG�����d��������FS��P5D�[^
:�]�{�PY���:����r��>��cMC����n�u	Q �1X��FMA�D�V6dL7C.�K�)�~66Qq�w�b�|'ʶ�j^z��zd�����?�b�摡��O>�6(A��.�yF�ۄ�Q�D)PP���*����֬q��EbQz���V+,�2�j���^��@x^����~|�q�.�° �?�k�4Iu��\P��`�	����i|�R�!S:�V&+�ea!G\*�z�!o*.x�u;�]���C!��0��L��Fʼ�o��]��������4U�@���q�=�5�u�����z��>+��U�0�əI�bB��@�%r���|�vf���l������O��=������g%,h!k�:�!���F�L�&�4X���0�kBA7҄�EU���K�Pgi�4 �8�魞HDP
,�~��W|���5�$��(�{c�ݪ bRwI[
&�D��;p9��ۄ�����֧c#N�gX+�<���n��|��� ��|�Ŭ~G=l΀0�u�B�Jd.���YP�;�y�P.	��-��$�������²�/x�M��o���qYZ���6|�g�H�P5 �H~T�Â�6y�eUM��n�ۂA/� �+�(��L1�\�2�v@�4O�6���������"��p�נ��s2�D)W�v��������^��B.pc����S	ӏ|zfJ�%AC$m�(���S�zQ�%
~A���k�=N���s�@ܛ]�To�&ۆ����	��}�w�C�^dU���r���n���H�jD�pȤ��r���F6u����OkL����FZ>O��{,��%�? �`\�����`�F$��xlouMU��q���2�{iy^��9��I�hV)C[,Ȧ#?��K`AD�����t�i�&٬Tk�tZAP7E���� �V�C����5� P��3mo�.9`B�,!�b#	L�j��
9��Mk��$��<����:���)}%k�Y�lg,�W�y@�T�~zbV=�	�t!��+����S+��Iӫ��'6�3р�фQ������饋�^'74������$.<>(�a�ߵ}�z�������C��Q����'��rY9~�C�����wk�U�wh��tu��>��	���m͍^ ��$�����#R~��@$�9�φ�r��K����o�󇟣�Q��쬦�_��M+نa��-1�)� �l`�.pI$�TP�WKq�gz�ۥ��]N�,�^�	@��_f��uF�.�6�	����c!�Za#���w5���F�@ӕ��y��Z���ť�٠�I�>GjW�hj��}�� x�nG�!�H��"�XX��y�����~>��~T2m=��-������_J������qŇ��X�P�ht��*��KC/�\n��^ �T�I������M�d7x�ꉖ�C��j�F�g�H.��s���3,�4�j<��1��!�;'� d+ �[��V���?$�sFV�:�A��G��Q6����S�AH!蠔�j�4�w�K>����Y�Ruu��W��y��#���}���#��=��#���*k��^s����~�<���tD8�M�T�f	]�tB�6\�ŵ��`�
C�6z�l �v� )x���[���R���`yi^����y4�5+Ive��@�������b��z��0��.��gH����w�y��A�!�
��:�0�q�A�Ȣ'�ta��Bc����0�<Po4��m̰Z��|�3�D'��13��k�W|�k)��:xn�+y�5�y¬$�[\�Z�b��\����#1MF$���w��,[�o�s��?vF�.N�����3R.d��y�$��D�����>��c��̰-r���.,��ع���zol��J��[6@Q��w^��=��ϡ�	r�d��X2�\r�\MC�B^�%���ͼf�9MO'��F�V���}��������0��8B� ���{<�&S�m�vu󭢆H'�:(/�:*�3�d9G�	F)F'-��w��C�do�����/��x��S#类e��낡���`=�͛[�y�����@iҚ�<�aU���q,|Ɗ�@�J}�*�q~�����|�����ٵ}�!���`4F� QJ�Θ�ó���	�4�X�.]�����aF<0�H% �9S��j�Ģ�2�՟�U�z�(�]�������V�{�d�����&nK]Dq6o�*]ݝ��Ϟbi���_�2RDG=��T���ַ�Cn��ZIgT��h��5��K�O����,�g�G��B2������>��cͣQ�9��J�y�ݻ�V0�C�W�͐�������[\���,7�d2BV2 
�* 0�ᑣGe)��M����!��g�s] �
1�t�ؿ�Q�b��A�Y�z�;�)5>�?M���f�B0�Z.��+ez��.sK3�O}������o�>��?a���'C�Z.g$m��cO(����G	��؟�ѣ��G��s�����^�7\Cђ4�,�f2 r�x��`G"�'-����W�8E<@%�i�z!W���'��t���d,�5�-�{MI�9F�F/�5��xX�[����������駟���%��w>�~��~�9FRz�yxǕkֳa0�i��F��`�8zI�7�����0;�_;;���3�7��u��,4���Yo��W��xD^!����w��(��+�K�z���c�|�4���+���QCi
%Ӳ��5r�w��]~�]�?�C9t� ס�/�tO��Pj�Er�{�*{��A
Q�n�N�@�	y��o���я�B�CV��p���^\��?T�XӠ�c 	��[���@�*C�[	�h&�����ʃ>(ǎ'�ՋɤۙK~�-7˯��oɳ�������JF��dS�|�#�ǎ˗��պPn�o�	F�ǹ�X@ ^9:�m��y,����^�����u�����������l	�P�sW��A�B]4��G�`�7��w����FдE�X��C�=9wa�����C�<L��-�~�_Tb�*jL������e`[їŅ9z���?��gE]C�%�
(
���Bj(u�8�=�tMC��&U0���L� t&�Ȕ_a������յ޾}��3?*���mD����
%8����;��v���Q���*�K:ʨ�5;;O��B�mɗ����T4(|F0Z��[�8��nۜ�����:^)!����r^% z uO?av��'�z`-�I�馛Y��>�|X~�C��~H��>'gϞ�p��,7��ZA�
啛7m�L�S�&*��Q����!��?��W��?��_g��_��+?|@�ǚF5�C
���$�l��P$�7^����h�w�L�|���x�[�y@y�Q�NwЛA.��F�1�Q��ߗ���ߙc������}���,�y.�f.n�}7��
�
" �q�׫��w�Ni�J��N'B��W�E���<-[\��dQ�htbC�򣅼l�Mzxh��ղ��B^&����]"��ʳ@.����
�ǔ����qΨ��p���:���wnf��@��I��0�57G^3�gXw��k�f!~�R+��S	�>�29�Tb�� �jE^��e��C񦇼έ�`ڤ\�J0&���^��M�F�ɗ`]�!jD�at�PF�Ȉ�q({[��!�e���O,"���� t�<F�4�g��ӯ�5����0��Cl4-ܛ��d¹��_o:F�'5� J|~$H"������c/!�mo}yP���'�OY��Q~H�:;efzN6o�#���,/��5�*� ��B���|�����/ȷ��	��D*>����������)M�|f�	V Q�۷����g���, 
!����]
zq9{��,N�yݲ <_���S��3��������-s�=}���s�*1��5����4��Q�de=��GH5�6�m�,�596&��u���?:��m���Ș6Wq �3H~ �b~YN�|\A��^v�:��j(H_o�[�m�V�8w�0�K�z�;Y=r�i�	�k[�]A-��蔅�Y�o��N���u� �.��tU
9�Pȳ�dm������߬�/�=պ���py�1�}BD'nr;��i�K�|l* QF�n[V7�`���#2`��j���r�t/t�
ޔ��B?W�A����.u��ra���z��5�x�F&�D)���՛�w�Z"H��}'H��v/ n��(��ϝ����>����c�ʁ����	\$S0���C�%dzrN�}���]�7��&炁��P�988�H����M/p�\���?�4b�Z�Tk�Me�"B���W�9ܼ�(�˞���1K�@�Z�Y�fj{�C����C|�a��[���{L��կ�.�N �nIV��!����D' ؤgg�)���8+[6�JL7߶d̐��3����*b`e�T	� ���%��^8wV��M�a+X����q�dȘv5�u�G�p�.�fX� �z�������>5b(��h*�6����iv�jWC�7~�ר���=�k.�)t���z^�P�jJ��J��%�:���̚�q$�f*���� �(��$Q���Y��:�ޫT��wo� On�X��^wc�-l:�������g� �e�с.�P�P6�G'9����B:7�Z��9�a�(�=jK�IN��D��J�F�h��	p�HTpՇ��K>���p��"�2#�����g+K�j ��E��qGf���dWJ��}]�v�87Gc���G��v��H�d�\.�f�O��Ǖ>��c�����-`X`��GfeH6�1���h��|��?���M�3�����4Jb��������27;#�(7c9P�4�MX7Y�|	X��	�<��&=ƺ�+2>rNA�(��+��T�Nk�� >���)�---�-l]�Y+d~nZ7�H�ʇV�Y��rY����M�7̋m_�ˬ�ZQ��z�󞷜Vp�$iBA�9��[� ���8�jJ�:�u+X�1�Tg=r�;�e�g�n�Oۗ ��zq��R�|��v=z\�]w�E�8��Bd�х`v�z` X��%�Mc���h)���B��� ����[x_ׯ_�[7"P�T�Z���{��7�eF����G=;����A����o?�MF�z����M�:�)P*$�HBд��<�U�OU.���� KK�r�vIb;�����]bJ��^x�9�ȲGI��4�32b����W~���5�����W������U�Kg�R��٧���m;to7�)ȑV�B��zT �)+'�̵�u��jb|\��mRW�|졇xl��$K�T�F�|Eo����e]q����ղ,.�JD

���b$wU��u�գ��4�F�@���AxBkMGj�<?#�BD�ɼi�45�Ã-m�m����/��{I=u�I������xT&�'$��T�dhd���<KW$ƂY�1��֟dh�z�)��J�P���J��l"��,�������[<`;���y�)�}��} 9���Gt)��Q�0]q�,wH���������:��%���u�_/��v��;{Vv��Ő6�~%#�J�Q&�0�b5�"��`H��^q5�md{Z�BFx������/�'�5O��P�F{�*CC�d���|F��eٱm����;���#������aUc��1����H70�Q���j�ƑZ�,���^d�������k�i7t�l ��f'�т�]*V�ĉ�����������o&X �N�:ɐ9@*iw��fy�;}D������(�f���w���<����L����:IQ���Gp�Ў;�˭��9t��g%*K[<(����R��3��lF�6���1�!,�]��ݸca�N
Z]�e(����
�mD��-� ��ԄMsA���\��#���5�rhd�u!�aj�a �c	�*@���]ު��6������V��l � �W]u��>��[n!9�閜�gV10�k0 ����<��K4f>���< x�]��9J���p	h��+r��5�H�����fm7�;�SuE� �4x�ֽc>�|��kt�q��G�:;���V���D��ܫq��%9h�5Fkt.[��G>�����yV�0hy4�����y���^FN2�i#��S�fi9+�{evnZ:{���BC���2���j�]8��<��Is8���D|�8\���?�4t#ut3��=�ϟ��'H^V3ܶ��P.�ȨkF�^#  Lq���=�y����wȗ��W��KGHx�aU�<[lбxd��u�b��0jv��k��k$�A� 뜓:�D$H���"�d��Q E��[�����ʖ.�O�m��J9� 4���T ήh�0,��S5����o�z�祷����uB��Z��!x!�P>L>����w�n}���_8K���x.���+܉�1y��ë�5�����3���2���ؤ��؈�����k%e���M���=�1���>�nc~������M��\<���ʼέ��O��LMN�����s���x�M�Y���hg�?^�"�>7;e��z]/^"Y�\�$/���P�һ8/�$��)�k`y<�V6�~�NP�@�z �.��}��RC�&�TM�yW�gd����;dxx����mˤeQ��~���)D����?�q����X��� 6D��'�ƌ�Y���d��A�]�9�`�%��͸=�EA�H,,�N�����O���y�ͷȯ��W���wI��>��4�<�����hl8��0u�M�v[3�n��*K�����J�Vd[�t��
�(�p4�8%��$ �As��Q�Ԣ�=��Ky���%J�
)�	��=�Րn��8���cc�= �Q��k�;>�P5�Z.�����Ly	�@���_'t�����ko���R܇^��7 Q���I:��W��s(dڮ���Ju�2��)+ ��-�)�;�|�z�{9?#�[f���Q�&P�3�~[6��=w��q6_��P9����fe4�b:��"D�D2�vRC�#LO�\J��['o�ݲm�V���ޞ<yJ��'?)+�շ�wP�5� n�*z����x��0��H4�D���K�R���_�*�\��Yu�k�n���{;�drbZ�uͶl�ȶ�'O��tm�	9u������G�R �T��Ҭ�ү����t�i4��F�Z�c�d]�z6'O�bh���+w$�-$ �z��Y�s���|�BO'�J�8��;����;��vپ}��7c�G~�f<a�t뵚+⊎8׫ss��9R�
e!(�U�:G��y/��W0Y^����V�H!`G-8�u`�c��}���G�ǅ�]c^��p���Z�9�ߵs��O������t�����:�D������K]����+�N�� =�Hؑٙ)J�"b��ɩq2��m#4��
`�]�X�U5�r �
�H�W��5������ ���7�5�;;۽f/5�,�Q���lgu�!:Mz�8�q��;(9="4�KY��-�d��-�Hld���|V����&@ ƎH��s�ۆuM�4��ظn����M���?�jԔC3�z%t���b��#A�e����t�{��AӠ�^?��Q Vm��Ke}����� ڵg�Ԛy���O�a0-#�r�ܸ���mvhd$R�ME��\���?�4B�jM7�jQ=�T2E{U7��G	f��F'�%X��ErU"#���fB҆U�T/�4�h��˩��R�B�
B��U��[���NZaT8	���J` *�r�z�ѰD�;uСR��?����;}�W*��`^<2��I��?��8������0q<s�����i6��U�>x�흒i���A����\��5��nV7W�&u�a�[� өU��s��#��e�fF?.�^4�YP��*p<�t��Y�Ww�P�)"�qY�h<�na����|�l�
p���Q���ѰC5=���H��Ԅ	������6X��tgR-��f�(��J7��!Du������"�kK� Η�<�GF��c t1`��p��֢����RL����?��qIt��E[�-r5�QVW#�[�:�8�*ӳr��9�iF$�4R���t��C�P����pߛN��s�����t�i4��&��lU���zW�*��e��"��ըkV���b�$+%�IÓwL�<�&��պd�&Ϲ4;iJ�j&�l�=�wǭ5���%fa�&Z���ї�pP��f�f8����ˎ�W.������z���^-��.y�Ǐ�7���v�!1-/����D�0��lRwtO�����<?)[�l�TG� ��O�����}B	�,Ǫ�<�����j����Fo�i�#�n�N��W�u�ᔔ�
: o;v�ӧO3V�v������y��S�`���J�H���;w���ٴ~#K�PB�֞1yjq��r����:�x"4Eɥ�za	���,� �0k���/-/�+;��*�DX�o�Dc,�߁�W�TɾG� ���bY.���Y�V�(O0	�{]�UH��229�޻@=�?�������b6+=@���7��0)�l�w�x6ݲ@�F��t,B�LF*��|!�ƕz�ͤ�䭒�AFo��ˬ��ձ[bm!ܧ@U
~�W|���5�H�� ������ag�A0���7O0��E! t[���qB�:�ꜣ��<�*�Q��-����5�Mh��^¼�xD;��X'm�w9��G�n]ꥢ�WФ��1���M"���iCz'����S&�9���J� �K�g�g���X��Nm�~Zj��C�������6��Wox�>���Fl�¦�5�Hm ���"F6@�ꫯV��J����Ȩ���2�~�5��Kޱc�s���qZ����E󛠓��������\���# ��^;�[T��� �
!���Ȥ��wW��:#$乙c+��5  ������$P����T,�.{�\,X�����%�6՘Hv���#r�M���g/�� hC� ������O�<"cS�rn䒫�J�S��+D�cP��G�w����%�< !$&#��Y���UP��ep2b�I��6��tvwɥK#�z��{�����t�i`����GA)
����1����Y�i�U��$CA*C�5�ްYb�E*4H�T*��r�h��+����)S5�&w�r 5��p�zu������|��>�M�z�[*�td:hl��Fn w��A
�X(A[(醭��ut�����':��^+�gQ=V4�V� �\%�I��w���F����u��-Dqۻ6]�q�Z�k�
`� � Y�|�@�%��J�����MCU��s�=�p4@9x��QB�k�5���#
�(jS����F��2��<뮤+�*�x:�L{(�Zq+�cewm�[�m���=oaaY�zz�q�	y<�~|>m�z�l	 �~��ep`�t�AӖLH~eI�;f�b�ոskҋ�[����	U�g{̰�+f>�s�x���z͓�]V�Xt��«p.�lh��'����>�������ҷn���-��|���^H:�p"����Wx���+0�&A�Qb��Qjs7HV�i���6妘͛���s���C �B�S=A���`
��гf�<A�rɭq��f��#<� ���e<`=�Ԇ�p]�_��CE�2��j�l�(��^�{{��H�4�[7�Ύ=W�ٙEI�z<�F	�����D����/2"�����'Xg��Qo�ZB:������E�Y��|�-[1*��N2���a����?��"1F�oPs��
���%b���K�ZZ�9�����VkޜZ��و�a�7��z��V����[>�����_��Ӱ����aG#ʒ4��!�������/:,���;�-�Fq�<>���q�&���Q�'{h�t}@l�46.��;�Ƀϫ!�Q���r��g�۷b�P�Z�����hB�`tp�s����EYX��X�j�Me��Ek��gG::2�4���U�/[�Ǖ>��c�CA�ـ���/�F�G���Je�QsHÎY��遡|���ێ2�is���!8S�DkM7R�]�+=FD�Qz�����	�E��u7���y6FYkldLNC���T�]\�ÄI�2� �ĨS�j�PΥK�$ԡw:j���JN��G\�6��+պ���V�a���K�^��-�4���bv��5�aU\]ץ�z�f������3JxV��j[�^w�u\G���Y�LO��5� B�����G��O���WS��g8YV��Y�>~�!�^�4\ϼ�}������g)#��� �J<%�|��	>�> ���}^1B�US+��I�S�|tL.\���4=s\���3S�$�E�<���{�9
�U��r-�Ȫ��֬�`zJx0�@z���`�W\wE���H�1}fhH���5�@`T�X��J��tv����˒J��R/�ՖK�\���?�<���+XBp���P&r�|݄Y���yt,q
��   `����� �h�V�ȯ:�XG�8A/��� �p�R�*��8۔* cSooK�U��ܼ$�	ܺE6o��/?@R�$>�<tȈ���Y�~�,Qݤ�If� PO=�.C[w�%�XJ�9������J!��f���$��6�B�"��s#���	Y[0g��Y���e���OJ��@m?�nD ֶ[B� S�C�B��>s��돂�`�M���0��M�$���;^��J�ڹZ�����o��L�\�~׉�x_��繆ۇ�Q%�2��w���|{@����g)�+j'"!J�ί���_��du�hX4k�� l�����/�ᾰ"A=tk(�l蘴�s<s�^�-����D,N]x��M%��yY��!�w��۷s���)y��ef��5[�|N�DH��+����t�y4�=�:HF�F9P"i�LQ�l���¢,-�P��b֫C��P<��':o��sG��? �!?�+�B ���!�f�5�ho���*�Y��_ݽ%�^%�bڻ�S�dp�f�g�����\������zva=Ζ�����m$�ojfR�ф�u��i�y�=���Ϊ�0��I��}���BW40����]���a��''�[���58&&�x���?�
�Ü����m u�M7��j "�mɂ o��<�Մ�qX����%�����Y��bH��T[�hq=������|k�`�w\�_��<�&`^����q�u�(�C�8  |wj�]�pA����F�%�鑕|I�(��pj�u]	ئ�[�l�����v�f�H�M��y&K����yí7˥���}N&���{�<s9ٱ}��z�r��z�	��x�����y�����{5�����IN�������?����kIݠ��Ն#���G�8 ����:sV�=��.���b<�-[��3:�@X���mf���$a�E��;�����F1��)��V�����[��f0,>�S��L�f�cW2u��.�NJD7���.zWTwS����Y?�3��` ����p����z�g�^�&<z^��\���n]����;Fu��X�MC�C4� C��j�~P���37nd�^�a`~֣��Ȇ����>����a5W|ǒ��:�`�8�P	i�+o����l�%<o{����Y�Co�����o# 6��,�0��S�#�x����%6��f�eQ5�`�A�R3lw��g�=H&�2~q�M]�MS�\�l<k��-�ɺ�xl���mI�Ӡ�~����P,�e��l�ݿ_>��2��o�n���O����܌tw$�#���x��/<���ڳS��}Cy�?�Ͽ��?���/'?y�Q*�e�#��Y�����t�i���$N�!C���k�b��SA"��2l���c��?~�sR��f�.1ݐ������ o��w�'��������=��Gn~�M�я~T�yɐ�Љ�a����-/(��Ԡ���_��~���_���u��Sϱ�ȴ�9�%?���g@ъ�P�ʱ�'d����ꖗ�gX�^�~R��!*�^�z��<�>|�ൾ�W�� ��wu���#/����$S���:{�< ��L+ЊG�<� �AOT���ȁq�g���)� ߃�~��E�Fc'�r�x����,�Ö�^���Ld3�=&G^w�:�RF�*v�z}�-�cbq�n,�� W�]� ������>�@�i�Z��9�~� ���ٕ�qd�޽29�,�?��z�!2��w$J�8֜C�:�
�xf����ױ����}�g�;���9x�9�������]�?�W�J�z�1�ʗ�����dqvE.���o}���}���p̾XSx��e�Ҽ;qZ�$}�>���������\	��2��#;vl�M�6�溏^�m�NeR)��;\������l�2�(���� 7���	}��W��x:!��v������p�;��`����{v;�5�s}��!�45#���_�׾�f�� T��g��JY�($293-��{/�Ȇ�cy¿�ύ7�ք��+��j�����6*_��W���z\k�]@�=s����S'���۶�~z}�:�r��r�������42���ϛ^�\� �u�B8^����� @p��[P�� /��X�]�x*u0�,Cݖ����՜z�#陜�+E},�φ��ZY���0��"��ɴ��A�@(���,t@F˲jCRi��(�C��-x�:$m]�no��SPc45�t}]aK]7*ck�5A����/�2���|G�G��GDׅ�6mɌ\�7�q�������d߁�dyi�kybD16m�,��^:��Rsr�jP��+<|@�ǚF6;ӯtJ� T��=�j��<2rQ�h^�y����v�ǎ��������<�M�$����}C���������~�dey�� Vaݐ��&<�/h{����^�Zv�ؚ��� ��c?���2=�@��w!W��[�z3A����譣dm@�iH�B�^�@��W���xV�ׯ��	FL���;v� Α_��m	Ҷq���]h*� P�EQ�ؿ�*���5�GGFd9�c{�-%����!qD P2��Q���<�� �����c=~8?B��dg=t�c/UM��j��b_�%��l9���:��U��.5[RՊ!�<�=���A	����z�ջ�Y-�zz��+�l���a!:�v�!�Zض}�[[��D P��H	�6�UAi#:�Y	ڢ)}�|�����������w������Q��յ�:9�ʹCuW��Z���P( �����{���3�べ	�@		ԭ�J�V�:�s�]U]9�:9�����>j�O�޿�1��:a�o{�+�5�|D=�uk�Ȇ+��W^~Q6o�Lo����������I9?xQ/6,�����*���{�t�
	c:��8��НqYcll*����ֶF�%<ԡ��ښ+��;9u�,��0�?��wl��� � 8`a�T���<+�vl7�@���(��D0XGE1���)�+��XT�
Ţ�9�&��O�@��n<�ܦ����n��4�"r���u����c}��_�mjX��ߜ��sTEsY,�b�� <@�9|������e�f�v� vzb\��� ^�p�t�w�;=j(\��_�0��X7x�F#�41���V_�7�|�s��v����3���3R�5�zC�#�����X�����K�p6 �:���)�Ҩ�^�:7���^�����I��ҘA$!p(��ܵ����脇�p_ax �a�#S*W�p��<�/�a,�r�&�����;,�_��]��{��ӀPC ����~��r��)���7Q;?��_HZ׷�i���OMZ=�k�J����U��S2��ܞn�T��IZ�+XwW�RuB�Θ�� �3.k�xV@xִ�ds���WvYŰ�#�����P�s�H����D��O*Un��-07mڤ�[c�6}�g��9۝'M�M��B�<r0�8!Z�h�bJ�nz�9zt �PR3I	�&;9>.c���.�u=��D+���3�5_L�=z��u�]�?��e6=� ��ad�?0�q����O?��y��2GS�NyT ����)������֮�H(�{�V�`5CܺF�`@.��$����MӖ��Ӽ�Nf#E��m�Ҳ3����hY�e76����\*�qi)ץu�e˓f�|�e�{�����|Xa{�;�j��H�"u����?b�׈H��7��U�H��z����p�xdbZA_�s��*!�&z���s�^�n�A::�L���K�Xa>�TO>��454Ȓ�Er�]w�����]���c|zTrE��A��PX��X��	:�e���
�A���8�2Θ�� �3.k���z�5�mz�ؼ�����IY��JpdAB�{�a)�eE��ÓKdR���-���祹�U�X�F~���dth�a�t�sySӮ7B��F��T�w<C�5���R�ݻwʖW_fi�q���ej|��%���b�*>OozӁ=������ܟ�w��ߙ�g�v������}�>Q�_
���ޱ�Y7�!���A��}�*�p��jx�(��u	q���a �`�|�����G�Ҫ�Cyd�M�38�~�f��Vێ^�%f�������ڶ��2y���=rۥb2����VJ��m�-�8�|��l[�j#���{���,K� .T4��(G�b�ӓ�j�i�����yr\�` B�9b�e�u��N�A?��]�.��r�g�ZH�X����i����Y��Z�� �u�Z�B*�<���� ����ݿ_"��4(V������z����gǩS'��e��^O4w ��>@w�e�?�G�L�M�����Jfe�����F�]8�*l�ȡ#L���'Z��.XgΞ�{�����<������7��/eK�
�F�kxRؐ�� ���ߵ�9�l6-˗,�?y��2��K�ϝ��۫/�(gO����s�9iQ����M��c��G,�JQ��V��<�����l߾���/�	\ ���+�6��+V��z\ ��dԻ}&���k���*�ͤ�좆^�F��4�@_�r%{��9}V�F��񇂨U��yp|D�y���6�@E#��9���^�SS�8P�}�-/�.=��ؠn<k&��#H[�x�����X� �K��MD��p�hXS����|&��a}�X����W�pC���-��7���E6�]'>oP��I>�ཎF�l����O�;Z���I���j���I��c.v����} 7����(#%=���6Bt���?r�dΛc��s���f������h��U��챣�w�^R�P����-wg��p ��5
���r��1�K�`��B�Bp�禨����;;�
>=�a幹�ر�D7�ǧ^�z{��p��Ҩ��}�2��g�'����N�#��=�<�Ub#%i�=��d/���1x�`7C'��Y=^���tn�����9�E�2���1�PW�l���i��uk֒$0D7r�P��ȇ�'�u�-��~�sy�/P�{�{d�;;d�+d��w�k4��Z\0�E���'��/+-�2����x} ��������z'ዝ��ġ
�����9x��C@C 9a�_G�(�ŭ>�`����TX����޷����P�~ ��ʥ_�G
�x����4^7�0w���5�A6�Y���Mgj�*�6�z��uk���|��x����M\���z�<zi)dg��9ǝw�)�]{���]������ؿO�ۺ��A�^>��o��sʥSr��1��#?�!# 3�i��;䆍��pE%RA���Q��(�[y�Y4�[��頑V�<7���~�3��?�}t*%q�3fy8���W���]���O�F%iROnB7��,�l�egk{��+yٶe���G?f/�x�ɐ�h��f��y�-Ң@t��7�Lk�sϲƺ���!X�����,b����Y&&�� pS4�`|X���;�HcS������;��ϔ�216IFu1S�B����\���dSY6F�E[,|2�?,[^MƧF��{n!�
a�B�Dm��x�Mb�:�TÔz���6پg����9q��/��<
>.	��;�o�Q\9�����D��U�^ü�9�C�D.�+��i�Vfw6S�]���9|�%�b�j��-����\�������P��:��@Oy]�2��2�׋v�Xs�o�7�� ��^�!��I҈bo�J�t�ӋDm?�=�� [����e�o�M�rQ �W�(�굫e��>��G?�4K1�џ�Q�λoD���1��������hD�#~�h�=�I���THJ,쑞��j�P!��b6%����٭�y��h�c�à�>�L�s�<+o��l��6W^���ݹ��p�)5\��O�u�m�D��{���/C1�?e�_������_G?�����Z{s����Y�;�C�
3�P��/�RMΜ>/�M���fj�SS�C�8uJ^��f��Y�[)��⛂ʾ~���F��_|i3ۀ��o�Ma��z�Vn����:Z�(���5 H0=�b4`���2=:"K�6*!w[��&�wO6��6<4��[�0��_��[_��]�5=="3�	��,�/驊�u~-�M��q |8c������%�ַ�Ź�MN��Y�X���X�IZ�i�C��A��!�kEJ���m&9�PLǹ�Q�	��04��;�8�MrkV#i���r��	��.��Q��F�q����}���(���9jz�%5�J�f��"4�6Kߝ���N5��Va�_w�q�<��R�y�L(���C`�K�b J��P���V�G^Zں�����j��)�J-�p�^���ѭ�n�ͩ�Q���;��<N��?VN˩矕9�]l�z��Y����l��!	�B�o�]Ϙ,��M�]��QkLFǓ29���'@	��ߤ�r��ϩCwƬНqYC�I�M�ԫ`�k�"GƸ��J99v�a +���@��F�
�1���f���c/n�,�v풡���,؜yX������^{���Y��r�8� ��w�̙��w�1�IN��]��^}EΝ:i�=�����ٓrap@�� S�iK65��Ç���U�#G�Gй��+��ڀ�-�\ ��.�0��|�JI�OJC�I�3�~�ٚ�
���|��:|V�z�t��@X��~��)b�y�!j�A�CFQ$c��	!ax�X+��1�پ�y0�qoи��1�Z~eOku1�c�rSs��R�C��"�A�AG	!S	b����N!��=�g���	ߠ�O�]���Ք�ԁ� a�������`�OLIGW�t��U��D:��x�ص�<���.j�g�Iz����:;�$�:()K������|6cڴ�T�ei(�r�����p@�ا��d� ��$s���u�񬍎����D�hK��G����@�|��U2��/V���b�g��p ��5j5O����*LZ��E�;�^eB���+�Ƹ���d!'�S�H���������jx����zex��=��#���oYܐ��,y���?8d�Lj.n��Ĕ~��@,�\Ȳ}�ӧ�5�0(+8�����'��\(IG���c��'?�II��d�O������YE���42|������V����y��Q��\�TM_v�r�$4p���m�Q�ӗ?k���b�3G�m��]D�^z�N>����ф�6IfPB<�c]���=G�+\��+<j����YW�ϫ5��E����cP��T6Z����C�%���
�Q,�:��e0��:�ވL��\B�B�!qz&�:}h@`�_�aD^���Xy}��d&ůbE� ��ћZ;$m�g/��B�J�G����
!-�g�|��(��NA����4Xc��YJyx~kV����LS��Eio�g�\���\�������Exs�ϕx*-�3����Θ��<Tθ�ᮺ�!�m?0�pB��R�>�J����.���mP@-���z(��K�gx���Vj���6eEy�g�C�fdD���� \!�
���C�m�jHLz\tR�&g���7�BZ�S����K���N�2_���z�Jy�������"z���0�|���k�r�� ����?{��� ��P��J�f���������{�Vm@a,!�mj.z���M+S#/�28?*>�߱6��QP���AH�|���9�s�iߚ��z�~����'h�F�t����UTjYS�&k�%r�v;R��i�B�9tIC2����V��hب�r4Dp/��g�$���8Ӊ$���J$��s�xP*��J�>��у����||bFZZ3$G˺�#�J���ΆpI����m�55�������8��"44 hP����T^�ѸLM�p^���Ѩ ��A�m�R@�a&�����g��p ��5���ڞ�-P/ �d�{:�e@�0�y _�z���T���?ۊf�l/ g�4S�@5�ӼUO��y�W�\Z��-���[�����d߅7mlb8��z�J�E;�z�7�ɫ[����
y�������$����麼r��1����Y�a���eV	Y�bt�1pM�9C^ZǺ-�t��+�z/q�cX||��ҵj�3�Y�:A$��(�-�
�������wWM�x /�z�1��\�m]i��'M�R)U���I"j� ]�8����_Q��#;�����^��Co��!2��bN N"�12R���h�À��h�� ?����EA����*qK����{&{F6����Z�B?����ʾ����ǳc���Ĕ^O��-�cײ�
{x��sc^�D��#��s�Z���8��7_=��nV��Z]�(/Ԋ��8��=@w�e��ˋ�$���f#tk�a^2o6P}��<5������P��eB솽��lR=/�ϼ���@���	F���Yb�x�-�':<���o�����-<� ����W^�w��utʃ~�y�ޅ}ra`T^{�m����������W�#.+���ٙ��c�!��a�*C�0���+�j$�O|G[��^��Y��E�<�~��a+��J%��u����k���=���t}$ǎ�0�Ǭ�1r� ��� %mCÃT�[�r����q{������C� W̩�����^�~�ZA@��.���tnj��t2Ź�x�A~Q�����G���AF���H�s�(��/����? �O�����Fr۞w�Ikk;�56g�����t!����U�>��8x萬_���I�c�������*ql�����Fԥ���n�i1��B�ҽ����O�Ղ�]�P#D��g�tJ��\�7�Τ��F�I$��Q�Egf���
��#��Y�;��%&�R!��݆BȺb��Z;'�2��PU%� CO0�fHPs�;6�A�JZ��b�O/
L�h��r[���Vq\��R�`���O�00h��rE2�AV:~��O��:���yw�N�{�B$ �b)Os~�z��}�^���8�%=���,/�?#˗/�?��g$�����u���.�~�z]V�:��)�MY^}�U6��F;$�@��I&Mj� �	qv�3����������z�Q���e	X�h���3g��c�=&����}�s��ŀי�Mz��#��d�T|�8K ���ǖ�h�SP���t�,�PeCi��|�75r��1�|���� ��5:rX��A�� ۋu
�x؏�b�S8c��VԐ;�^=Z�"J3��CS���op*֮�B�9��> ͭ-�>��z�X�˻=�Hͥҵ6���HsS��� �[���=_�P��̈�lѨ%���(�w�3fy8�������"���<)6\ts����z�PR� ���s��T/�����{x���PSl@�l��G���)�d,Ƽb�����FY�`�l~�wK;�<CQ7 s n��m3���u��h8���_�~v�Q4`c����c�v�b=z�^[����^OKs�tv�K.�d�Y�/�e.6idnD�ɩq�ó�I&f�y��a���nz�<��0y�򞸌���<���C�Xc��7���Y���'��������J��ax̙;�k�χ��4�W*��VȨ�65�������?7=]�̤�d��\�qN8am=<w\_D019%?�����½�dSF����I���l���O��܂��4Z��nnl�y�L�N�-��"�T�����Iޫ�I]��ٳK�y��k����ha�L[����x+W%������yz+�z
��O����Ӹ|���d��>��N����\83$'��1��djbL�݀+��3�1��tg\�p�Vjހ��I8�W�H�¾$�asY!wxX3�=�@�O7�h�B&M	���O�я�sU�r�W^y�l߶� �Ps �{ݾ0lmv �ݤ@���l__	g� �A�aB�ؠ�z�)�) 7�t�}|�}�3���˦�Ix��\��nqy�y��P��:u���ŗ_V�4]�i|�_�x1%I���N���(��5aH>���ay[(Ŀ�Τ,���p�|��wf����j�y���[����G�w}^�F��?s��&&��7[���W^�����N�߸�s��b�2��-��� �L���V�c�؆�6"*z2�����G�;�k fCe%c�A�����TD�����ͳ�6? �!���C���z�)�a�w��>19&6\-Ξ�4pS�A�ZL���v��L�����S#���=����0�	׈u,dff��-����4��C�Ի�zd��+dٲ��s�.�pJ�VTTj�C�sƬНqY��������b���Ke��^n��희Î�ǌ�����uG�0�7����h�2���;r�7�|�<�����A��׿�Z�������X����l/^5�8������6�<�zG�Ǥ
�r0��3 ��ƙ�-U\?�ؔM>:_'H�}�����Fz�6����jJ�u�M������a���XБI����Ҩ@���f���"˗-����Ĥ]�@�5�z��eͪ��m�v�g�D�� p#��G��O�9a�Ǜ��Rqk���Xߓ�����˰)�	����KMX_�[��_�ͣ+1�W	�j�)��øh��k��V���zc8�M:)6xa��<K�P���~�S5_�[BM� Ϋ��W��R���%���}9�RQZ�%�����!)B�U�������!����QJ�b�Xa`Eh�.��
�R�\�ׅ���O<����F�n�:IL�3��=�WZ��ok�KwG'9P̧�WO>��[Q�U+���g��p ��=��ZW�o,� k֮�W��=W��E,Q��������g��_��I	�ƌ�Y B�h`�S���X�Ȇ�U��ޕ#��u��i�b�U��bsF}5<���i���?�@���" ���F��y��[.&�T�G��[2�׹/����bȭ���R�a�o!�[�ȥ$��0������祩��Q�4H����k�1��L��QH46�d`pH���]�Z�z,r��Y�!>��1@�o�.pm �h1\�����A���]	��5����Qo?�B!�u��n�ugn��7�w\�y���A��)��>?�C�4Zۚ���
v @��f�����
~��`����4���6��.[İ�a�=.��LN&H�ǔ���?�3�=$������[Z���MNN�: B<c�VN=�{;>9�{A	��#��n+�M�9��g�� �hX׼���$�p�A�M��"PO!��("����}���}���Je��>@w�e��[�-@�</^A�r�Ku����6�� "�
,k�.^Ȑ��mS��x�Q��FV�gZ����+$�����ɓW|T\cx����EӮ4�75�.0t|�n�SgN�=��fY�h����+����i�([�X.�)�X�A��;��zz����!��!{Օ��1�=����;v`:���Eϱ��p`z#� w������tx�1>��ѣ��p�T��#�n���r2 >�<6;�QXŴ�@����T� }塺��& 34@Q�A�@=p��!}����bۣ���nT���=�A��Ax��l���m�4^j�t�Lb�������o�-�S��X� �
�Hp<_��:r��A� ���c�� ����G��D�P����Ul�g����HVDy�)5����: ��&,z-A=/�	�Wt�1����-YL����C4��o~�r��!�5D��I8r�,\��u�'Ύ��%�d�|?�b.�ӯJHL��v��g�Ru ��>@w�eݜ��pDA݈� �A�6���V�Y!ﾻ���m��N��<Tض����;r �a�DX��/��6ѫı�Ի��I4$�#�^��%S��wSc �/*�u���?OC���M>�˕�V��]�V7 q:��k��F6n�J=�݈�V��׾�m@�rɆcq	��A�F8 �ӗ*F�n*�Uc��G����-�ǰ`���nv%��
�)�HF����q�hz��cE��D$\U��o�,0@0_C��a<�4�K�c7J�`< c
`
�������jx��Mc�
z�p�霑{i�l��B�$3�ƒE�h�����w�ex�i����l�5�5�7Q��4�0$v�e8Px����w�X�]��cg��a���Bc�o-�x�HU ��*�BIz���|�K�z�j��?��<��/䪫��_��_���ݗe|t����II�
��Ц��?|\�z����h�o��t�z�xY�Nٚ3f}8��� t��k�4����D "xq+W�R��j��#��N�ܪ�I�Q=#��'Ƨ��}���M���J'���qCf4���Q���¥ 'x�^��fL��
K�Իs{�?�:��+lk���w���ݗ���.C��.�o�\}��*A���	�Za����ѣǥ��C����$�.R�ή���Ъ�8�k�8B��<�bހ4ś���'��;-�t��(P��hmc�z&�p~R��!BcZ���i �!����T���sF��Ng x��&8g[.�ܹRRO������$�麝<y\�8ɰ���Ar���a  ߝ��Xߤ�a���S�%�f2��c�#�FA$d�\�_��6�~�g�
�yMN��#��,s��{܌d ׍�?"3�z�(��1�c�E�� u�tV��GY?��;���QZY"I��J�͐���E���q�,���R*�׾�5ӗ>2�m�5}��9[����7�J�V��N2�������8��������8��<@w�e���S�l&$J�\�^C�����9󥣳EQC<���,
�#C���ƍ������#^����>�Yٶm+�Λ+��x��h[��O�v�2B�G�!pa`c�j ���pCj(x|a�g�y/Y����� ���d篹j���g��FQ<���r���w�PTV�^+��P4����"�\?���1�<�q y�d�U��8F�-۶���� �� �u��yF�� =��ّ�\����z~УG�4:��\�����$������\7�K���|o:����c�� ���:�5��0��ZR�@��`�p9��B����N�Y��WW�#	B9�����>�f:��W�(�~��"8�ĭO��k�
�R�~l��Vm�K�1�I���;֮Wj���"����!��7�E��'>x��ş��Ϲ3��w���FR���j��L����|Q��w�j<554sݪE	�erb��Q���*����Y�C���j�]�V]�\���M���QC]t�ԥ��>�
�Q�
���<==��R��kЯ�5ҡ^zR�h��������뮕��?�e\����.6g��dF���M2���l:�Z%���M��w���9))p�J5	E��sK���I�"���D�U�0� �t�2i�鐪�n�S/_N��6�bq��e�V)@>/���ꥡugH�=��ib�������z�:O��\�: u�w�!
�cht��bnoP���%�w�d�].��`I����	J�S%���:o�����^(KC�`���\�Meh �cX��Wl~�;*J���'����3B�%*�!ڂyn��WB�|��=z��/W�:k��P�C�����W�:z��]�
�^�\�ϥ�Qq�%�����
�>��$�k�&zm>o��P�I%f�U��$�t��5�Y#7��J�Z��t=������|�������� 2`�]�&dIo�L���gd:]��3%��-����	�����4�\O�{��>�wP7t�.g�uƬ�r�e����&]45��8
KҮ)2��Pegws�h�q��9�3��0K�ʬ����?/7�t����.ϰgË7*byؼa,����O���Nom
J������x�T{뭷$����+����GY'�����E��w�/-�m2>5�s�0���><�	ݘ��n�	��JE�j��˟�#�O˻���t��ԩ��ͦ�l�Y`H7�^sE�y�@�lw���� �I����
G���(�F9T�`���`�S��{��:P�C(dE��ff:������X����� ��$�)2��9��]'��C�(�7o3�a�� �z�р�Ü���#�.��5���*����(��e�2��d��ˆ��T��*#�z�{<�<:�s{~�$�Jyv�Ct����@%QB}:� ���'������[}a�D>�	Eb�[���ko�"}KW�ј�u����ys��!ʒE��&Ϟ��[������+��3�1��tg\��U��]C^����X�d1�~e.��{ɒ������1��7�i¶��� Ȫg<|qP����ˇ>�a�����{�Uo�,�����i��Ƹ䭾�v��T����  ���ǎq�G�Њջ�[Ǐ�Q����ѻ#�d믾J:�c���%�<�$�b��4Q���$��ꁖ*e��3w�;~����/X���\�rH�f��`��
���p,h��E����c� F��N��2r�YS	��EA�EI�F�Tҧ^�b���4�IΤI"��� ��� �5�~`�27� Xd����]���װ���.mv��Я�|,��4�m��
Yۚ�l��M�)W�/~����kl���ԥW�0�ۊd�g�M_s�9�s����;R��"~L;W��-�y#����a����0�mT�00ix�QB���:z}g�Lʊ����&5���[7�ƍW�!�2��ӢF]Z���{���Q����1��tg\����%��P�#?	� Z��5�Pr����N>zw�>����O�{�~��������ٴy���{�����m!�%\�3Gn����h��kW���3�:���/������-}�����d����<���{�r#O�\)We��

��M�����#�׮��n�M�~�m�5� �X�A��V�����>���K%�]�v�"���[dx�";o�����	��3���2?�%��5�����<]��?Dxة.�c�d�ɩ��* �	 ~��En�r8��X'�z���܆z�^��U+�����'k\�(���H2x�L �:�B�`��!���Σ^��ظ	��B��j�?�!���f!��j�j1���v��j���k0�pm���w;�O��%�m8��.I����ހ}n�k�����i�n�+r��7��U���O�a�G���i���5���[280.�-���2w�G���>@w�e��[��C�Uÿ�|QF�'�#I�3M(�T` �p��Q���b�A7K°9�ܹ����0�`����V X�7T�%�fL	�D�!O<�HF>�xIo@=s�S���g�����!Vȳ��f)i��l�P'S�06�������3�.��}˂�>�8�>���6�w�X��㨿���wv(0o ���F��z�'^(f��s�.+̍kR��9O��_�����8�U7�1�$�)m�d�2�1r�,زek�)�DbjX-�Aq��'�i��6b48~l#4 P�=X?��Y�N1W	#z�b�r�dHd�M[Ey�HoV#�_���g�F�ǘ��1aT��7��F��Vo�4Tnk��J5��m�� <�[����o{ܶ�o�6"D�\�r�M��U����zw;t	��������V�����_�������TcpP�zk�^_B&Ʋz�sd���F�O���S'�:O�8��<@w�e�j��Η�UR��6Y�/�"�1�3��t�p�_xu N��St�B�0X�]m��Wc��K뱃l1Z��� j4q�����p�q ������ϙ���e5��1&���a��m�t��e�8�	���~���6[��0J(b��B���ak�毠����O<�24�@<f)��x$Jp�d����:v��jh���e�>�}��-v5�b���d>�w�^��� ׎c@�^;�dP���B�_��Zy\������cتr8�i��#��{+
��;�]��ikm�@"h܂h�k֒<�셳�p�f�ղg�Nٰa�t�wpN~5�@8�:@�@PY�Oۺϕ�a��!�Ӹ���k�@��+60��z�� �F[]<�U�N����#'�q`��M��}N�E����^Lȡ�G-�9�tu.�p�QΫѵf�:)�^ĳ�
G����Y�C���	ּo���7�j�k�`���t��;��

¨͞�������6@l��4��2�ө�E��ՠ������qk�ѲQ�����E�BH�D;��3��y���y(��@�.�E��	�Z�(�e �B��p8HOӉ��/��.�{�"�����W���9'T[�҉#�:��������5֟�����%#$�ɦ9�ֆ�L��%VŴ�9�.4QN���ĲjU]UI��;��0b*=�R�e`h��Ćf2��^���0Akk��m���y��M{\v��q~z�(��䡇����I!����Foz5rzΓt��<4�+ղ�}��������Ǐ=J��m0�Xyz���w�2��C>��!�C��n����˙α������������A�J�Ҵv(^�����/�� +Z{��F�F��IiR㳩є�-�c���,i��|<.�W"����Ę��:cև�P9㲆��/z��*9Z�b}3�=%�xF�eF�D�L����f�s4"��R"�VY?���wv�R�D������ɏ�7��[���4�]l���/�H���&��(�I�G=|ݵpdH)F�V�Ur��sVϮV%���H��r��iy���h��C��QS������!�d:#7�|�D�����>*{v�2�`:%!5�ȵj~���<�q�_�1K�9������ԣ���1z�K�>F���PBC=:��m�\ ˶����i��7�e�M����H�K���T������#����6�-��wv�!Y�l�s�eR�3w�,[�B~�O�C`�\�"D��!��N��y�5�kG���-/�K�#���0�M��C�&Oo���/@���]�Z��c��ư�8�M3��������Ź��VYлPj^��5S��\���ɡ;cև�θ�Q�T+�`��e��e�6]T�{H,]���5z�~��jV��*�i��E��<�e�,zl�d��o����#��&�����>Bڨ�P!�ja�y�{�lo	�	cr��B)�fL����B��wn���un!�W��m��{�;�3�ʙS�����r��Aӵ�S��s:���S�+ɲ=x�W]�^N?Be8�E/�ڙ7��
������Rބ��U���M{Q�qW�*�r��>��an�C��DbF�� �� ՠ�	���V��s��JpwAaMLA��~�'�K��wY�A�������s��R)�0T�a��9�cr\߃����w�p��^��O�'s���<!sj7�{0 U��`��g"Fji��b��b��mF>�cs�����s���G�1N�8I��ھ�-9]�I��ʢ��e�6�
Uz�e�4>jz���7�LHCK��kB� N#
Fk tX�Θ�� �3.k�Þ�z�U4a���0��Xfki��52���Xm(���P.=3��X,W)���5�GGFXN�M�56nl�)�[��޴B�x�l{m�mϚ6��i��u0�&�}M�Y��z��}=�qr*!}����>)�<��__�=_�5�jL��2tq@̟�y��W^u�T�>��5�����r�y�ͭ�iW,o��j�3���0�67ĥ%e�8��C��R���5M�$�z�h �F-ȹ���Y�F����y��/���L�\'`�#�B"�r�6������έnh����+$�k����X4,������{4G�y�o~�_���}�Ш ^q�����@�z�86�WK�:���(=�߶��c�+�|�[� ��,#�J!�M��K�l�����鹙*����Ƅ�0�c� �Wb��>gtv<l�Jp�$������?��_��5��LG��`JB��Y�;㲆n��b)_�����eX~Wp��������p��7c���%�+>��O�}�c�°��V�y��ʮ];M����k�GM^=�Z~V�)����;c}  O���O
�T��K���d\���{�֌��z�P�V��(��6m�$ǎ���(>�A8����t�����E� �h��|���1G��m��>*�ny]V�\.�����[��6F
��*�6z�{Exa_[����Sr��YY�j���_���ܱ]^z�%���e��>��߽{���_�9Y�[��̒�/~�"x�<p��q�m�ax=��Gu�?#��.�/}�o����?�������&�Biki%B�'�MS���>�!�3<������Oפ!����0�>$�x��F�t��Y1i)��q;��W��.�iG77<x �����{"2R���9�>���}�����r�R�ÇL.�(ĳSRC4�b1�צϻ�"-m~�W�)�̵LO�HM={�'@�hmm��3�1��tg\�Ѝ����k�LIR��|.���y"��W���wx\%��%B��x�O���{eמ}d��ܸq���_A��{F~��sRIE�4y�p�['j������m�������x=~�˖��0$��nɌ�Λ���o�믿Nֺݛ�z0����~*3��`w�v���rZ�/�e����b�\��!���p��iiX�TV)��)@���wG���jS�c=:�4˧>�)Y��m���򋛙{�xݵ
��Ɂ��exlTV�XF��/�KXo����P2���<p���|�Jg,\��=�m���z�0�Э����Z�[��j������ � w��9xh��]}���j��0�^<�v::ۨ>7�w���G%A(������zo�jƸ��6H{�G����3U�3iЊ~`\Z�v���燞�Ǌ�gHA���M�{����̥�
�3�Ȼ��䆛6Ȝ�m�S����d߾29�������.*�TN����;㲆n���n�C�<���|�ᐴ�w�KC.`��Kl���a}3��[�IO��(,�ƿ|��<<����o��%�����_�Zrټ���YU 24�AL�����Gk&��2�U ,� ěP��n9��X��" rl���sH���I�,Q_��������^xAF�%����1��̨/(���ˆ�{<�2��=��_ɉS��z�U�~/�N*~2!�Bt�C�B�v�.)J� �?~�19r𐴨{���~*o��]���,[�\�y�Yٳ�]���
�y��4eh�����~�3�(+����}^��47�����S`Nw��u�+����nr֍$�<r��o+��5��aL��_yg2)��ڍ���?�w����{���M�|�R�Qo�o�4رіz��H��/=�v4;�D��Sϓ���1���d8��n�j�����<��J����/B�_�z�H} ���y�5�Γ�߲Q"!F*�Z��OP��W�����d�oȡç�]S��T��i����;�F*Uf���y��x�sϽw @.�$/��ի)^�<���
<��c�Y��ںuW�=���\�Z�����KOwER*d5� �1��H�^� x��������O����3)c��Ӎ%f��F�yao���d*9i��f)��)��������:Ϥ\8wJ���v6��X�� ������L���G��Em�{�
�\&C� ��fG�!�W�K�у�u�#F�U�����9TCc��oIT����E��*��k���a����Y5�^���x�0�ʛ� ^=�~C��h��O ���lJ㬼3�$�M�z�Ly�p����u�"�䔰�y�ݻ��^ܷP��d��^r�,�3�ِ��k�;�>M �q]�sf{����V�n�cwC���y��Y����-�������,t.Q�����Ck?��Q��K$�u�WȠ�e�\A���F�/}4�pKE�Ʌ�;o�{5"S1
���I�9��4@w�e�_�z@�&	�խ��*7�t#7`�����G�SU���/�;'O������}���y�����W%o�7�|S��:-��q��K�7<-���"��V�f����e{f��H
{a�f*��n�d��1,
F}(@�w_�b(��,�Պ��aX����/?��Od��iY0�KƖ,���]�l�P�D*+C�3����r��=�Ikx��-P+s�q��9��@�V�v���C^W/���^�[_G'�� �p�@��G�4��w�gr�h�S��'L8��B^�PG�oQ
 �K
F/�7;��ܱ�TxSo�̀ȿ�;˜6^�Q1��=�@<��W�{n�����@���[�&]���k,-u;��zצD��{��6��w�(h�a\��\��`M���X�xS��.\�F�J��}{��=`Ń>C�<2_���5��'+֮�e�7�=�Kjʆ�	4��@"�Fٰ~�<��k�͋K���Y�;㲆_w�x,��ʮ����޻��ȑ��S��\������&����n�W_�b��k���#k��@�ح
s�tˁ�����������v6�v��&���D����ٟ�M7�O~��'B�_��$� ����QA���}������BA��Rc9�|�V����v�����r��~��4 GELj!�`��$s%5z����HC� ��Ks<F �)xN+�������m�s\Kj��k�$@��U�`A�e^�L��k�Yy=V;�
��C$b� p�{��I��ŏ<��g�QCo�U�Y�gSs�t(�
"죞ҹ!��Ⱦ/87�-0n�f��0�(w��M�2x���������{�T�!�����O�(��.{��*T��\��۞4�v�C��Z�ҹ�zVc�,B���V�U��@�#	�J���,���'eѢ^9y�ϵ�ͭr�m���7_����'�Ҹ�6�$W��Z�~�$�)��C�����>��"��� �m�H�Rg8c���θ���֯Y��xV::��ƛ6�&�I21-�(�.���m�0���.6 9w�<ʯeيE�}Db���P�mX�<1:y}�_�%�>���<�Fy��ڼ��u��b���,�\.�� �|�f2���V�x#���Ш"W�Y!?��I�cA����s�9�f�Ź��Fjڹ9��._�ܘ���gN��b�h��Q�n�O>�aI�����o%��P궢��w�N����s�S��������ab�C� ��ym�� ���I��xh�y����Ĩ��J�b�+�,Uc!F �p�<P��ܠV�~�b"�(+0����9o|�����y?��!�{��A�<zo=�ˤ�����X�r�dR3�7�#�2��h��׀05����u�a@��aɦ����ȧ��0Mc"�Ͱd�
����#�߇dp�T0޲����f�����4���6��q#��<�^������R�{�h����$���l$s�ܠ����ge��9�W��|�e�+/�H�H����I|�ؖϱnjj��Ũ���(�z�b�2~�=��&�?��8��=@w�e�����������^��t��IbfJ�ᘑ����	o�Q�e$��4O��"�0�W���/Js{��\�Z��>2��ы\AmA�؆�v�Bĳ����t��m2��@��C��)�R
�n�[E�,o�<5�Q��l�a xtn ǡ�L&W � 4���ʊU�e�w��[��'�T�K1�����>�~�[��L�wv�Թ������N�W�k�N�X�z&\��W�k5!g��b�z� �a� �⑃l�&(+�W���&�����#۷�u�֑�p��Q�����`H)���5V ص��9�������g� �g���O��C��Ģq�������A�� Z�*#�p׽d:&ށ�ё�_��g�����7��*Sj��TC	�����=PC'�1�����G)m��g�R���q�`�Xf���:�1�a��1\ ,T)������ b�[ ���8.����u������oB�B�X2�%�`�/o
����[n��'ϐG�l��L�X�sjX�K�W��)<g8c�������=on�Mw:��cS�T��4��xز�v[Kx����
fy���%�V��w�-�ջ<z���w�_9w���d��FF�5�v�n�Pݵ:� ������3Tߨ�����u%��0y۠����@�`s����ǈ�$SP�cI�#�<"��1Y0�[���Z���eNW+��ăz=SE</7^'7^�����k�ʲ�YK��ȡ=�$=5� �gLo�*�	�lR)2�M��Z=dl���M�H�g�x� ����X}ק���C��6�e�t������ �-�]�X�f�c����Ő<���\��{��["�����)������	�s�.9p@�ٹ��AG�'�C�<��I�5�XN�05���{�C��T����ǚ�؀PPY�n�/@�D �eS���#��#��J⭺� ��Q.,�|��Ft5�RΔ�!o_(����C34�����}�3ʴ�ٿo����ԼR*�dF�Ά������=�T� ���i��|�@����Θ�� �3.k�s96[l�`\C�-GM�*7��d޼yl��:�r�"n���t�iǈ�l|���7�%����K���?�q)��֛o�K�~+i�[2�5j^h�R���y����Q�<22"�#��9���s�yZv����Jz�K���5�0��G�"%���4<����*�4��d��H�gY�C��OJ�+���ѧ3yʯ��;���+8�ڿ�e��259�P9J�pL�����Any���o~��R1��($��a����R��F�M\����=���1D<�%g��y���kX������Yϸ����C}�!qpVyױ'�n����\-#��U*�t�����Ŵ���w��E�L3}��w��_H�ټ�L- ��^��JI$g��N��`H�iF:������`7���n����G �_Z����^���^S(��x�} �ُ'�\��}D�wӍ�r�
�eSlV362D=����=������z���ǖ7���i�W_-mme\���^��{�� U�kf&g8c�������n������|��J~࢜:}L:$��t����L� �ʎ���[���?s�]� �N�>-�?���ww1	ŭp�4� �&;\�!�����
�+�R��!^�O|��-o��ߒH0 s��]ާ�)O�+s�/�����h���0�}�����!�\�|�3˖�7IWO7��Ȑf0�$���̤�6=�������;��Y�&�(po yW�5/ds�˟�B��ͼ6���m�~�ht���p��{ǎ�A����W��3N��11>���s���w�
+�v�U=�Tvܰ��������>����dǎw� {��)������Y�=,{��}�XQ���%�^9T ��e�P�;:i���1�l�Z�Y���g��|��7�{X�4i��&�`������/�� SO����j_�H�V�$�h��4���|xI� ��n��&��׿��6 �|	Z�Ui�k:���8y\�u�X��`�A<'�׃�Ap	p߻�:؏Ǉ�_ϜN�����Q��y=��d��ݲg�.rR��+5�v�֜1��tg\�ЍХ��ʠ��n�F��O�_���Uoo5�2 �0:�)h@�t`p��Ml�� q	�P �����Y�U��)z���2Z�rSL�p$fB�"�%��u��w�QcC�p�45Fd��U�J���6���X=�B�K/����!�b��m����n�������
����%u>)�T 1^)�;������o2��S��"aK���w�)�c+��{۶m��c�T��z&�� p��=�JXq- nD$�<�6miޏ��կ��8G� ��K���в[��0��x�<�-��50
 �E_t|���ԎG���`��ut\{��g���S�6��u��7�,+W.gy�w�&/��U��|��E�ʡ�G(:d7T�yC��������%�M�s��l"�y�:w�������ܸ��D����Jkg���_��\�f��ՠ7��#8L��y��F��ׯ�F���8� i`Sx��dD�A̵�o��9{Zn��6����YP�U����Z��g���F���d�����g��p ���M޳�k��yA�9���%}��X-5��g���lS���	z����k�0�O|�S�G.udl�x�
�k��G�������R�W��J�!*T#�{���!�=��S��sϨ�:.{׫�TU�uX���;�9oeۙS'�?�����.�7J���<�� L������Бc
,
~!�	�Jd�����H��Eɪg_ �/ ���R��eٚu��k[���%ndsA^����уE�n���@�OܖsE����ҧv����Z�Z�ה�.}(�G��l5�
>0����G��� .v��Č��'>)���y��W�駟2�
p�hL:;�����$�L$/�u�]�HK�0qm��VAGwk�C��lg�mOQmp��QiWP}��-FI�X�����=8���̛�D�+��f���+�9�
L*�S ���q9!W��F��5B
��z�\�B�B�`���T�X�*�"P�tRc�!q"܎��M��ٯVae�jAr���R��c����C|�Ϟ?����T�Xɻ�����:cև�P9�2�Dx��wn�ݏ�#<�b�B��g�k]�t��u�]r��A�;q�@����=s�'t ����`�o��d��(������)����R���8'<�r�L�yaS�l��(�
U�̋��zޭ-MrH����=(��88u��^D��,�h��� ���!�� �J�۠_�=CO�����D�j���Y5��iw�\
輽}'��J�4�)"iK��{�[n����O�d��>�;���p(���k�;�Z!m��h5�l�u�v��Y����(�\�]	�0(�b.��H�5����:�5�'z��P��_�<��+���&��IvE�cG��7���/�~�̙3��3�ú��\,��� �x��u��m-2��[����q�d�5���|��߰�J!'F�h,�,.��2���޹�c�����/�� ���O�q�~�����rT,mF� ���&I����ѮUǽƺ�9���_�����F<Ͽ�I�ီ�\2���:�F"�gq_�듸^���&&��g��p ��>9�������W 
�t�Z!uy��y��7į�,<�Qݼ1���/���瘫���kY.�M|NOK��~k�{�1l 8����b���u��r�i �z����=��fHb�� W�X7��~���կ���՛��6ƃ��� :��D�!&]��r�1��Qҩ ����/��sd��j���@y����/��oB�`����?�R3���=�̽��P/� (D D��6���-a�;u�aDẰN��Gc�iDJp,|��ۃ� O�̔ J��\g��5�&C���G�S�%�$z�.�/�Kj�m��������:��PB�uY�;_�X�JΝ>Ŋ�^������3
.EB����d��"���q�s0���u���޾^����$��[m��]5I}�y��	�:��'��M͊���+�TϫTK�w�z�(�@*���ıc\+�� �	^$��{b�iv��5�:��OI�ܪ��>��\��7*�p�,Н��D�����"F��jaZ���gw��t����5`�zM	6���O�k
B~��r��w���0ˆFG��ȡCd�{����v��U$LX���7CѮ��'vKA7gl�02�/곛c��,_>� �2%�zy�lδNU�Ĭ�xc�='��b�������Zs����?v���ٽ[bQ�e��}�A��'>I��_<��Və)����g˥�a��P`�����na6���g�l��;<o���>�W̍����q+ꁿ�/Z�"k׮eH �(
r�۷o����T�E�+ZZ�EFp�s��rM�F`������Rմ#u���񐆩+���<>�u���+�-��O�8�m��-:�$�l~����>b�)��2��=��IY?;2ԯ���czF�&�$�7�sE�{.��j�r�暫��ֲ_�_�L�p$���b����L����µ㳈�@����5�$�������[��lI�nD��eB���#a�֕��8��<@w�<���m������ۅ>�U�k\�y?EI\�n�eZ�����L�8�U@`B��������{��uUYûr��I�n�eɒe�9`l���`Hü�`0����<�,g[�eY��d+�V�s������k�{K�������u��#��ֽ��{}�k�}�]w�S��k�Z�'g�yw?��%y=�@4�O���ܠE
�2Ӝ%R��n�Q�c�A�L��2:�G}T�%�޷�>�f5���B�.�gf��'���6�0�m'����eL�THI��$�}ۖM�{(4��{�	z)	��n"a��i��o�s��S����2j1�0��Q�x�~�/�6���ODJ��tʮ�;�ְ;XǴ6љ$�!ώdv�T\ V��O|���~B����S�`v�g�2E�<ET
А�/�,��<�><���Voˠ{_!�nvM���y=$��Q���pe����*"5z?�O����^3������ �JU�-nOI�[t��!���T���ԲP�t���Z��-"&� b��ky��GG�u^+�(�gKL�p�����싞/@� �vY�'p�-��8���Eb��5�z��*��]�f6HT�-F�����	�,-�j�����L(6Px�Ua􉞐'{\�l��R�t2��l°����𧪛�l5R����+�"֯�X��je�QO=GO3�HK":������N���Rp�#ǎ����us���)��l�Z�b���q�Lim�l)�S�D�eQ����"A��@�Թ�i�Ȝ!-䬲1c� x� ux�X�@�S��k7uA�>|�A^;��o#_�� �Q�kȚ�a�>r� ~<x�o���epȧ�K�1 �R)�ﰥ�^����w0
�`���O�]М�r�r�n��=�K�`E"a�	sC�F��D'���G��V>�I�	�Ct�+�L{�ۅ�.ϙnm�DG�$�>����j����+7nA:%���ͤ(	�7�ms�p����~p̐��ŏbC�LaP�AZT���˦i�D"!�l�ю�~L6�~�BB(�#�:��8��q.#?{�̑l>�VhpB���1�R�d$>tcv�鈅�ᙣ3��� 
�7���kEh=�`�P���t�6.ʋ��B��i���/\OX,X��0��Eo�+��� ���	|�Rѡ�T����G]���Oʴ�3��e���M����9��T�z�%݌�0B�{ۤ�]�vI���g����m��+�G�c��n�')F�Mp@�޳]���Z��m�����$��8 z�`��| $�y>�n$����  H�O?�s �p ��t�ʕ+	�&�>*_��ef=�}e�+�O��a� R��C"#״Y�XS����F�����M� ������>0���%S��H�9V��'��������KVn��J�٫��(�D|��p�`�$&s�;�F��髧k�LC�(��z���Ri��~�����4�����I[��cj���>A����\އ�A�������>}�NJ��|H?��Wy�Ϭ��$�qA��d�.���8ϣ�q.�s�T�4����b=N��8�%�#��^ج��+7�B� A�V��}�$|� C��"l����[ ���xM�9��_�e]��ZV��[�!����������������Y+�p|k�T�G�)�R/�k�e(�s���Co����M�T(tB���eos����|�?'t���K��T��;�BUR�^֥Zω\=��Cx��=����+���f���g��rH�34T���n�aD@�w��۷G�,Y��8tŃk���rm�-����&�_K�"r�0 X�U(�ۑ�����ҙ��&��!R��b�Zu�`�O&R������i��9*sg_ǢDx��kU�w�p�,]vǞ3ݒ�Ee|dX6oݬ���/�Y�UX��c�>��9Sϳy�f�2:���0fUT ���w}7��[[��3�c�]���WK!����TC�|�Bd�E5*Bj���h�@�ʨ��<*�^oLNV�ٷo�n�N[V�X9����cμdm��h9��(�ۆ���p�d&k�OvEcW0s<�|�E6��4y���EP�3?Fƴ*����AX��XW�^?��m�ن��ͯI:>���
Ѣ)��_M��Bո7 ��v��4�H��P��4�g����'���́�9�7�c]rΡ��Ǥ��2��������k�����&�d��L�P0�Q1��ZBM�^��'Ήc�����ڭMqN�<�9s���0�m�}46�C����%��}�&9t��x������5�MY�;�і)����:TE̚���
�Q�&������-�W|�薭�@԰:��ͦ'h'��N[��r��1MV�]�p��Y�إ���7�@둅��)��V�G<z?�̤��g��iҫy���ǧ�^8�Fޤd�x���XF��^ ����yM��Ӵ��zC <�G�_�X]�9��e���<�d����#r��Iٽ��?tR��\L�8K��TFe��Q��x�c,����j�EmYV��OV9��)�m��DdJK+7�޾n�z�)��F=0ژf���K��<���w��V��@BH�f��dZ�z� C�6�\;dlx�z�5��r��tv�SZ�*(��!�x��1w����ߣk*���,MO��}~xm>�ݩ̐�.�`�$���2ۮ���ק9���wC
�bz{��_������Ќ-Z������ �gI\�<�{~��Zr\è�9�}#���� ���cMlз�v���D	���/�'�=�r���r�r��y׹@�ǫ�E��K/�,�^����~�i5z|�r_r|FDI���	��b�ye\$@����7z�j@��,��%6l�������&�^zY���=uj���\+�r�h�[� ����Koo7ea���
5�� �(�+��@������6<}����ݱfx >Q�xg�e����ZJ�!�5m�lX��鎞<��_-E�G\���^}5�7>��lڲ]<N5r}lؒ�ʨ��<*�^o{D�1.��!q��z.N�{����3d�zY+W����f��R���y`������9(�9��둯���r�k宻�%q��)�ҥK���Y��N9������
y��<������Y@�������$S�?� ^/�p���!	��exBdނ��)G$�DH�Z�EӼ�@�s�e̾���u�8+�-g�6wDМ��(A!Z��%�\¶��z��`�d��;Ը�+��!٢�P@�&�l�����e�Vss���d˒�y������Kz��j,?k�*K�.'@!l�Ndl�r�0�m��a<~�fwo��3�����vz�0 �����lY��a�(�/�(?��${5���U���y@=pT,�C�z�
jN��gr� �@��OA-��ۡk�:��!�U���ɓ���{�G�����z#�F>�C��葃l����)M��;Ŝtu��k[_�|�jȅX��~�E�J1[����@�yu��S�Q�t�!3�,d
c<:�B���4�P�Mǥ��$�f���C���������ך��t�y	���뮕��ny��	��Y���+㼏
�W��!�3�s�����5�6ˌ�3�+��5k�ғnh�/�q�_�N�_DM�|а��\��V�^#+� �;���r�W˲e������Ш���)�;!�
�u¶�i���^k �If%py�����oH=�t�"zsc�e��d`pD[ڍ 
��|^����7��(?���Pl�ʥ�݂5~�U�
 �`�������F�^��[n��\�zТ��2¸ �S��#�����Az�N���6Y�F���&���������p<��烬*�u� $ԝ777Rm�����Ϟ=[�=N@O*ȡ*���,O�s��R��z��g����`U���"�덜�~�н��i�]^�}$DR܎ �Dqzz���-������ȡ7c��3����(�<��AĀ*�j��hH��� ��<I�q?4|L��O�aw�����M�9�f�@�U-5u�j��r������d��޳K��	�;q��(�����g�c����6O�E/Y-�f/U��/u�Z5`��N䤘���X�x����{�!�Ta�W�y@���=���D��X�98�7K���
�  &�(�NƢR_�hHm�ID�g޳g�;v�ʩ��ҳ��G>"۶�&7�t�z�U��|�]6�d=0B�۽¡�eJ���w���j�p�ۧ���M;_��c[���ӹ��V���H�0%U��� cB�t\�پ�52�� ��� ���V����e����u���@G8J�z<�tfy�8-T������{��ʤ4�X�"(G�V�h7�6�VY�������P�MT�g=o۶M�C-�� �Rt�21�EGS�s�x�a2���6��#V��<��R�ϴ�t�D����g �@Dbp0�G���ř� "��F%d�c�!0��5�����*9u��p��n����{#��Dȝ'O��x>��ϧ��1�L���X�`M`0���6��	�R��=q�ǃ0��Cn�ʗ���M:H��)Su{YV�w#���;R'=]Q�U��¥%������֭a�{Z���6i�eK���W)�OH*�(�U�y@��s��%��v>���|6������f���n���V`�p�2I�����?r����L�a��
��ؐ�����!�@յ5$��졳�ʪ{vXyxlش!�2:<"����#�����@��3�Ĥ��C�(��2���r���O�[�[���<��3��y�ׅ������hH�s������f�&@���R ���nK��aI�@��~��d�*��sV�T����t�];��~�����,��	�ܵwL�� 0�ڤ80�O(h�Ο˰=���t��!7[��a����Dk��|��s�N��j8%3,|��!���BT���IN�:y�R^�r z~_�G�Nf�(硐M��
���b��ã���X�h;�̙�Ƞ�O��C�+"aj�]��A4"��ү���T�RF�FA���)�rJ�2��xX�+.�L���\�/�G��AP�(Uᠩ��Bς����	�#�����{<��ǔ�-�ؤ��9�C$�H��FE.���O���>*�^�2���d@��a���2U7g���m�S(\��(C�K��<[Xb�̦?(C���M/"/�O�R�8Aю4������;���qXlx�\w�x�hՊ�(�>�Nm��i���T� |YEک����+ܻ�b����}��Kk�}J��m���������a��<��5��<٩�i�����!�����2/��!\*�ɘ8��15b��5�L.����`B�T"��y��l��F�լ@��a&��Q��!�����îvmSejk3�$�3�j���YMm��G���8�RQ���3Ϙ��
lj5)6�z�`1/��(����1]�<zm��� -m�h���L���Ei ؚ�o��ed�d�.��ƶ�,�����޻h,f��腡�� ��hi����t��?3c>@$E��֭[Ձ��Kj�@`�}�\����5F�j$�5���L��~o�:M"��w�A�\�Q�E��z|FƆiP:Q�Q�q�G奪��=�ɑ�����@7J�1kJΰiN$RM��ߡ�6k���A�2��(��x�]� ϊ��8��R]f;O�dP��(����H���
��d &�����d�9>�;=��N��{���ﯪ�
���ή��K&�!��ss���jڇ�ۏ�;�t�z��<g+�!�˲:�&�Ȁ�!KLz��E���/}�K1��  �!IDAT���׿&0�h�2��a�za`��~��,h��R:����z��"���� �O?��\�a=�� ن�&�{jp�Pps�M����qY�j��}睲q�S�[�Dv:�t�~`G11Q��?X����w��l<7�tSvXt�h��#5��kT�[#F㤲�E��!��󗉋8��%"B�`-}0@�$�"ԙ��N��a�5��lP�Y�x	�h���_���6��ܒv˖M����Y�uu��������sF�/�@H�&	E���'��H>C��W�xtlH%����o�o*�2�� ze��1��Su��������acSD������,<����I0`�b2\��3��pVt�E���������R[WCO�NV]x�\}��r�]wJ_o��¥T΍�r2摗��;�ƹ��Ep ��L�"������K�&��.Zg��I���^��R��fP�s�I.��D	}a������m`��=��rި��@H�Bt�VI�PM(��,h&�#��01R���@$@#�����Ѝ(J� o{��a��k�Ex��`)�D��9|��_0O��yG�5@����F_��������֖&�!q0Αc�5c�-M͍��C����kd���V���u�~
�45�赂4���oji�0����9Ͱ�X녇��-����ݱ��X[��i��ǀ�?�q�:��=t|�0��#1�}����ܧ�ᕗ�R�� �'��qih�ȩ�#�6s����^5����
iiE}���d|Xv��.yɨ���W�����ʨ��4*�^o{L��N��\i�IN��{y����>MF�GY�@���ӭoh����G}��9f��A��Ƿb�r���?)?��e���r����� ����!a��cz��?vX
q�����u�־	0G��۾������~��5���VS�	0�%� ���r7���&�KMD=�(����aF'`$`�_9�à����(A �{}C�����܇n^_��Wy}��'i�wۍB ^6�ap[5�s��n���ƽ����g�k����@�W�FJYg�XR�N�>�����{﹋�������r�dxxHZ�"Yvҩ�ն5+�6m�\ W��0��LLf��뮓�~�+z�P�[�`�x���������Q
,�eb��d��ݖ�7����9'&S7��eD(���z37��р�B[��cɼ�R�H��:�2Lm����~��ҵ�J��p��{�̘�B�/�!SZj�}�f9߾]d��[����S&ғ�ze��Q��x�Ý���b%6@ 
��(j��۔)meB� �����;��9˟����ӳ����?J���3嫷�ƺg�q
/kn[�[���oſm☝K�f�ɔ���G�����z��\42��W {�PԪ�/�=��F��e�����S9�u�M7������7�=KІ�x��Ο�K/l�)�-�O}R6l�� ����xP��Teۻ��O�x�{^����k�M A��$�����j1��`y@*��nw��U�0��)��w,΂��K%3̯S2�(�M[ؑ��mx-^���n5>� �y}2]=S\��ǇM#�зo�*�#� �1?�SG����dhdT�M>p㇥E�,x�����$֯_��eΗ3�O�0u�:��˺u��~ "��s�I_� ����y	�H�`�h�R��$�!�)mS���~70�<;u�a,�A(�9��0���$OHC(,;v�k�y���x�O�_�J��#E���{O�=w�F�g���0�|����W�y@���=�Z&�j�O�823�|0ڡr�L�z�iz��fB^�p��������۾cG���7	ooP�������� �ʶ��cCE���<O�p!�j{�����xF�������>�[7�I���b�� Fv�M�u)>hD�GX�/��NKK��C����HQ���A5b��w\s�<��C4CF��-�KK�U~��_���2k�,���W� �Y�t[�� s�f�s�vT��1R���;{��vZ�{˱4�L!���O~�����3����a	�)ȓN����#�u�$����}����Ƨ�U�z?��z���q���d���g?����5���7������_v٥l|SWW�����R���1ft�w���/�� �m{e;#h��:���u6W ���뮻�x��l�o�y2�@>D����q�w�jL�}Z05c�q��C��W_&3�̤���7��'�]����}R����F�5F��4�ފ�^�uT �2��hj�1��⋶t�>q�����&%7s� B����O08~�$��h#�)�5n¹CnSn��_��@/t>�e>��yݔ�D^�ͦ/�r(��?ȱ�Qr�Ժ��ˇw�4 =V="	ӦM��� Wr����轝�G^���Y{����>ٷ�i�
�k�G�Ǣ���[61 �Gi������Db�^%�b4��A�~yf�$,�+B�&�P*G"�:�H����z�J�$���6�y�T.�h�����4�f��)Z��:�9|���Q��a�ȇ�/�c#d�����?}�������NM���J����n���[���������m�5��:�!j���x�B�.����_��e�X4��{B��ITB��A�^=Ͼ={�]�'N������[ϲ�����7��!.X5��:�C�hu�3��ў�Cg�TZ�EOP
��<����~?6��-��]"�Ɍ^�J�j�20�����x�Q�mT �2�e�͝ohj,��Ƈfx��\���86C��p ��*Pf^���5=��jlݼ�̂
z
����+5��r�9^1mZ��Ur���6�5��A�Mw��/�,��>�Զʜ��e2��]=*�׀��d�^�?�A���b.:�>f��y���>q<�q����_(d�S�A8�����[ ���k�ԱV)�4�D/;�,
l�;0�"3Ɛ(�Uӕ��[A��A�������|r�[����^`h���g��SO�SFI\R���tN�U`N�w]�5�WABG�Μ!�_�^^����t������@�\s������
l[��9	oޜY2>2��p<w@(�5c����u{�5�����e��	骼!J��P��Z�*]{���Z�2�m)��:�0m#ѼV� �3{�L�!���_����R]g�ytM�6��J���p��/T�?�pȕ���ȿV�y@��s���ǎ��j����3wY���D7ׂÄ��_�ݼt�N��V��C��H�=��L=OB�Nʪ�L�����cQ�rC��_X���d�sރV4� w�q`T�����x<����*����z�N�!�P�V�h����(G&3�W�pmM�:���䥻ׄ֡�V�Po��\2c�,�S���n=�g ٩^h�Y�]{n6�H�:o�u��@oe���'n�ߝr6⮟!|�ܰ�a��<E�N������h�R����X7�L$��N������Ω��I�5�C&�Q�:�E<nlNR ��.���͞-;��`�,=}�S0� �%(�=�=��`���f{W�L���/^�0����{˥ihۇ�+�L������������5zKF⯆!��)�a������1}w�$�%,��3M$�����hL��Z]c��y����b��_�T���F�+�m���td۶m�qD�%�O7F�<�2Y�H���G�Mݴm�Q���&�;]K�)a��R�I����`%1:� C[� p�9hĂ�-)�F	b�)ꪱ��	6z�5��m�U��q�x���V���ʰ8���Woq���2�}��68��lx۰p��Ǳ�'��jI�^7���@�u�/�Q7�F�5���gXK�}K}�=�{�r�ˬ�w�=y���ӰA��#�ys�C
�_�P � @�ܒH�:�~Q?�¯��@_��2�l�j�����Q?���ǭ�cBBUKM-j��j�/\-����7�������@���~�I�
���u�XWKAT�1�B<X����,��a��|���e��s6�s�2�0��V~�l�t��W׳��*\�w�.�&4�����u�z_^��UҦ��ht���*���8����G:�q�����6��D��ɿ�V����dr�E+t
F	�O7Wt��3����`������ջ����4>G�4:2,5�uE����w�o:�1c��m��[�n��pHl��d8)��wA�Pr����7�X2h۩��%:�g	E�0|��#�>{�\�����+M�8вn;W��AJ®7�`M����e�Q�<W,��=/{�vn㬗.�(CN���Q,���/@k���z�u�
��C�?�t�s�m�T�[��^�=ֈ��l_�¿����X2+��L��nYtՕRLg�ﺚZr|#i0��V�Cy��)�#^���+����X5���|���I���
�`:Zb@o%�� k#��(�ߡ��2�0s�%�Ǩ�(jpT;$���ѱ��_��+�����1]�[��R�q�G�+�m�X,Wz�Lr�*^6� 찑�i��AY�4<;l�`�c�X	�g�w�I	����tJR�\��>�P���'J�|��0kk�8o7�XI�31�uFq��i�00�Zt<���	r�ɉI�M}�OA��B����7��3]��j�Z��1��B�zA�%:���S���B=��U�u?_=Ť�7F�k��u6MR�QF��Wj�a�7���9W�߶��������ڠN�v8���dK�Z��2�^�z�%��7�ְ��TZ=�0?Og3� q���ed�N�L�s��H�C?��E:k�%��?���/!S�ġ#��8�����B
�z�dR�_�N�z�u4�z��0t�D"/�w�|ɤ�A�nIn�D���fv�>���N0_��^B���a-Dk� 쟷�{�����"t��J���Z��������dE����3n	��R��������>c�VFe��Q��xۣ��:��L&s�"=S�}��5jγ�"�N��l`�{�F6@5�TdC�YQ�E
^Yx���[7�n�Ep�C�#˰��6�8͞�w���K�l��7邩A�(B���\$�p���%�H0R#����
ֱ�|s�����)��<D�����Ƌ�W-��߾ �I����8tN�xKG�|�3���'T�����9�h�«����DG��Uo{�(�@�ո�1�l.k���F��3��e�%��.B%Y���Ψ����X{6_,����j �P<k���>���ԖV���e/z<_c0�P��U���*�)���Ճ�j����T/|
5���R[]/�h\�F�28�w��߭b�����q��dB�eR����H��h�,�炪��4u��]�����a��A���9�"�Z�P)np�_��kR�"( x6W✲E�?���]����z#�����Dl�Qg�!��[|ά�L��5J"L;�u�����{��6I��k��k�O����� �)Y���8O���G[[�dG��O<��Z���F���i�ܠ��U +��Vl��b��S6� H����G�t�k��d2��wU�PK�s#r���&\���^:� �s�����Zt��<KC��M80
nU�5�v��Qz� ���!i���9�f��'��Mv��@X6UG�=�>yc������g�q��)����
����ڵK-\luO�X	�F ����Y��y�7mZ�`�T-@�0B�l��5DB�	?�}c��"4�}����v�+J�0g��'�����i���Q j��S��ĩ��`kkkd������XL:::�����;|�0C�RC# ��ʰ�]G[�E>+�*DW���x�)"
~ |��y}�*�O��涙R
�q=/쥗n�U�Vr.C��2�Ɋ���|q�����}��:�&��K�1-�f��F���������D�(��j���X:E���^�yF߯ںF-j \uŕ��X'�?�(#4����)j|U\�z�"��p�4����z��"a}��"/���?�]�m���`(y\��Jze��Q��8��[�pa�#�<���cn��Q�3����07�z ��v�0�F.�Gт�������7� �-1y�|�R~��+[^�f�JdX�\n�bm�vh�&��$/���aD4˴�3����v�':O��L�˶�[���ȡ��G�u��[&�,�T�@��oY ��w�sց��y����{r"�9��-������p����=d�תQ��?>/�����eyz�?�0=l����׌�n��~����-�?�-]����=��#������_n��6����o ��>�1~�{��.%X����(��~]~������/���!��ԧ�������Y�9��/��"���!�����X��`�*�*��{��n��ɟ��g$�-S䦛>*a[)g������������t�p��j^��%By���^qS���p��r�����~9|�0���>#<�J��5�&5��zlZ�G&��G�:���F����v�P_�����}�V;�;��{�{�$�,A�w��:���p�|��|���b)'�aٰ�Jik�h4+]]�R�V����T#��Oڦwȯ����a���œ��*�oe��Qy�*�\�3�H���eX^��!]�t�!��ysd�u�����x�����D�=���W�X��M2�� ڛ�.du���"�|Z7z�=�2?NF7�ܳٿ�n�M�w�����	v�G���=r��X�����{��r��7ʶ�q�>���=X�CGʝ��-�#�'7>� @j����w��a��}r�t�<��sl�ZRGq^t�$S@@:_�fs��7.tIK�s4ka��AI�e^o�OU9D`x<���<�a�����.���{��1Q㋿ñY?�������΀� �^. ����7�7�Z�zڱ�;�����hl2�B�h�jV��k6g�F``�(��8�Ii׾�.Fl��)ٍF-�	�1m�z�9��b/�6ly�q�ԣ�;26*�%,.+��eE���fٯ���ۤ,�(���3Hm47��154%f��0�\��\q�e|nXCD_6>��=zX����W])���o��Mʔym��� GO��r\�z�S�Ζ�sfJ]}�d�	z���\ �Ϝ�9��ޔ�i(ɬԡW�y@���=t��n޴un|2�vXm*�Oko��s稧x�����*FEΡ�d�Pl��������x,*O<�Q���K,>�R��|����5<��;)fR 2��j���1ӯuZ�<��Tp��RC�Z�F�YW�t	�{�A)HA{�	��
����K 4��_8O�,[���V�cE�u��ռ�k@� �H���NɆ���UoP�e��I��$�$��е)�� �L�wmPE���/��;����G�����������w��g�F�w����������P���{�5��uu|4���V�V����g�[� ���غ�e��/Z��!�.iD`��~6mٹk�d�����
T�C%��������~�I����+�g���xB7���g:	��,���и����G}$F�i������,�c��>���D��2�9r4��w*���R�U�.l6=�KLrN�]w�\p�
������l�b��f�?SD�w�V0/�E�6�eW�����S�����ٔ�����%����I��2*�F�+�m�l'N�t���p��f�t���
��?�Q���wѻ��7B��I��?�����{L3�����q���b�Jy�ŗt�N��9SfϚK��i����Z���.�j��Ҕ%H��f��O��{�>���+e���
�9�Q72_�^�|6�x���r6l�B�8@��z��\{����?����r)S�b?���hu˙��׹�"�r9���?/����<v@�["7��������� �4�)חKv� N��0��� rl*Rc�����px�v<B���h��n��v�^0���(�u�Ñ*�6"�g�`����}��ځ(�ɓ�jmd�����癜���j6a��p�Ե4��������LN��"�4h���^%��� ��;��g�bVoi�|w@Dd���T��7٥��·`�B���M/q����y�K���!��D-^)��f��XTF�b����Ғ�LK0�c��w���0C������؍KeT�y@���=Z[[s�-�z���-M^?ac_8��:qLڦ����L�ou��_��1<ޕ�.��w��Gum��G���vʻ��7��u�� >�����~o�9n��O#Њ�-˯��~/�j��T��w�)?�(A*�V�Z�*zy�O�MK��#�^��jÉ�V�f�4?���H��v�<OH.mr� A�Ćk�y��T)p��Y�r%�g�+&G��y�ү�^X�o��q� 5�F�A���C�H��y�Zem6p��s��ݑ�6@˃����|���g�?̃9rH�	���+�n{�;��r���gh�?����?�I���x<Hv]���=H�<��w��P�J=��x)]�H�Z=�,k�!�LH[�t����HMJ��`��;z 8��hH	�/�c��A~�B�z��kO���g'݂z���Ө�Y�o4|���AQpBP90:��B� �6�[0��iB���ys�3���d"I��O��R���%�3��󝆱��xG�����8���q.��p��~�ח/�^�n�`�c�۾��%O(�����%���OA,˰�nh x�;v�e�W��W\Cp���g$�l~�(��]��jwP��6��ޤ�3K�!��K�)����̙8�	Wɐ%����N�OfҬ��B�8�D,�\lM8"��w��VOMI�Vm��2frU�������b~��組drPԳ �t�������Y4C�s��9�K�ێ����{��ӫΛ�=X�8$T�f`���|��q>����t����w�����o|������\}��4>����(�z뭼����^�W�9�{B9߲eKe떗�6'9-o�|��S��bw�n?A���C�)S0]ѐ�/du�]
�x�rE��^���a}c�z}�ԇ��%�<�ɤY��֓j� z��0���ߝa緋/����ӝ�I�e����]��`��y����)k֮V��t�z�}^�`�����'#�Q�yT �2�e��U��z��x|��46dx4���K����̔�e�e`����k�`d_�N�}��/��Ɠ��w��1
��wv[�|΄I)|��vMu���ظE� ��!_z�|�+���{C��[n�K֯�O}�S�;��q�r��>ʰ�Wn�����H��l�E�6j��
���q���H�x8dT�p���H�^�_�����>���7����b�9�`+���$)�}�o��mذ�-@���I��,C淟�G� x�����=2��=� mם��`�q0�x����	p���?�a�P�4��ڧ��@���׫[_���w�����[G:���hiJ=F<��T'O>�y�Ǥ�O��fr��/�嫗��[%?��L�7K>t�$��뱏+H��s��y�d���� ��g̜ɵ>y��:rX��KMk����73�s��qy����(b�gS�b���ܲe+]�i<�R�P+.^G���ǎq=��8'��H�$R}�[)p��&�,� >z=�ʛ{���+!mZ*�2�� ze�큐�O>�-9�% H�X2����.�|R�@7�h4.C#'eՅk	v㓮�3d�.cI��r���ɷ��=��o���e�{d��r�UW��Ȱl|�19tp?�Q���R���z�^5�̃'�uk�����A��+VPS��w�K��أ,k�>�eRS#/1�Wx�k׮%0UG"jd���g��7�浩
��E��!�c�e�<4�|�۷��4�C���Q~�� g竩�����z���#�s됐��̰9�����_�E��ܹs�@ �,�cl� �ED^x�j<��@�%��]h�)����	�A�?���;�x!�Dn��~��r���a�%�mX�|�t�:&c�잆����d��E4�}ة`������_��+��T}f��|��o��/�R:�������?"����\y����}�ލ��c������N�w���+��52ej��{�]$��]��>��쥗^ʴ
R��#�� ���{��#ᵫBq�O@)��]��v�RC!%S;�$��r�HN�8�sm�r^��^�}T �2�u�NW	^�GA,��Wt��U���a��.M�w;�c��u�F����L�U���w����uy��G$:6.�m�
H,>n���<&L��o�Ac� Bκ���)�b� lb���#�������~��,:�A�ddxX���os��wN����y�/����K����,v�;7���U����{���,%X!ߺc�+��w��f��4��V� p@6��,��X'��W#z?lA� ���]��/�`H�������@x�8�9������Gdyp����.m��n c�l���*Ќe�����.�L�'��a��3�<˹X���"P�����'%�T`��������_��Ng����뮗��u���i�>x�5�����ȣ?"�\��!u�ȇ�/��|����;���7J��w|�A�:uJ�c�<���x?�Fx�=�(����73ʀ\�����ګ��a5D�L��"_�kw��A��`��y��]I��ZԸ��T4��zQ^۾W�	5j"2�H�2*�<�
�W�9�;X���Ka�yII��{	I���Ț�6�Kͨ�54D���� �6qR���M��{%�W��/~�����?�/�:�&��ς�~��[�%l��V3<�O����&�����oHl<�\�S'���,�?�r� �D,�F�G7n��TE�<q�j�,Y�D}B=�	(q�(D� �9"/�d�B�E�x�Ϛ>MZ�UArphPB���.���A�kb�r
��;���߰�y&�*�nx	<`_�^���F���[⚸K��R��{��k�/��r�@�I��1;o��~Д��wX{Դ��G�׵���S��W&��hÿa��cG�\��PȩϿZ���;���d��t&bI��V��.��xB��n�>�+�֬��3g�z\�.}���ky����� �{��d��r��A}W��Ç幧�f�;��u�� 0T�n`����~��7oz��	�F����M��%Ԟ��ǥM��d�		E<r����n�8�^�?�3 ��Sv�ث�_�^���R�q�G�+㜆n���pU)WȲ,�`ש^�B�ٵ{��������߬^�@x� I��M' ��ƍO�c�="�Ǐ2g�m�Ay橍,7C���3)vZ9W� ���=�V@��b# !䋰0���<�Q����A�ē�6�y�U"��9�y�7<6�{D������=���d^�#5$����g%><����H�㓆p��wz�t�˔�����6��!w��+0l��#�`�§M�N�5���z�y���Y<c(��댬_����.]o/$QsF�=]ៈ`�-X���nGxv>��9A�aD���Gc����U����@��5��O��
z��t����c��Le~=�H�G
K���}j@������>�9�Ŀ���Ȼ�q�$&bR�}�kx�D\�CE5���U�*}��ɠ�>��{�K*���}j�>uBЇ�����(�(��
���j �������Ts�!�N�*)|�0ŉ��e�+�_�&�V���QN�R��N��8#��t�ڋ�ʡ����/!�Q�yT �2�i8���nҥH����pʒ�Nw�&y�+�d��X�mk�c�Ǩ�
3���P��+����a|rB~����p\Aʴa�S5�ނE�@B�_7i=��Z�~��Ϝ9-���*���
�����z��˛����ydlx��XlC�k��F�=�y�D+̡��O=K5`-�z#�#�^�hm
o#�^�m��Ǟ��ߔy��5�m�܎8`�)\�n�s!�a�PALs�9O���d����� + 1�7ae�f��� p� ��ڹc�Ug_*���1`4���Юk�<Z�Y�.k�r���)H.o���=����u/^(�N�f	���(������!��׾ʨG@�sh�>z���:��-_�t!'�g� ?���K6��}���{d��9����r��!^���#�/�������S���6J�m�`��=sv���D2ٔU�P���zQȱ�Ȏ'�.5B����cR�����.I�2��%��]��r��K2��ѢTFe��Q��8��(8
U�@��5X��1B���X�R?s����ꭍ���db�3Sl7A}8J�N+���FP�P�'@����^��EP�2�|_��רQ>��Wn�� �I&dHAr��e����Z�������"����Bi#�OŲ@HN��y@`$�W��Q�Zc�\R�\/�PS�^5�ﺰ�ڿG��#T�{�٧M#�Y"��Ҩ��끐��v���nwO������~9����� ���)΃|;����]�Ʀ&��Ǝr����>�bx���o����7��^����:�#�u"hI���	��y���c���Le���)D4��Aܮ"��@h@��ӧ�ʮ]��r)f&����!/>���S	��w�Apt�����d�O�p�)�鏾C��J�?��K�բC��e��I��3�}��!a��h@��H�s������D(�y��F�t�Q��8.oI�./U�R���<6$�J#|�!py�?0�-��OIu]�d����8���qN���no��6�nʦ��9+$nJ�|^S�+�u#�r����!;�͖����	�ֶ�S/�.���M&&��ߡ�K��z��x�4-Zw�W��;�2{�<� �\� ?��_�m����=&������fMѐ�X��mjn6�b
Dcј\���z��;5�Yu�&u��Q���D
����i�n�`{C��u�ֱq
��dє���:s;m`�����Ϲ��������M�X���Ɵ�������
T q��e��x2�,��- kww��T�ӵ�9G��X���q^�Q�'85�hЃTD\����4JvY}��H����b4�2�s�Ёߴ�Eٽk'��{�G�(�Z������3�?CO:�NP2;{w�.�_���;g= ��/�G�����	Av7�����:u��]so�أjat|��@S�H��k�XM�y��#AGX<��#���k#|�q��������	�q5bgϝ-C�c���2����T�qN����
�*����
óF8�^ Ox�B�aq��&P�Vw��
���}A���1l�̱;��e�ӂ����T�\�����Y���=���mV�wu�f�0��0�=^����IP �����MM<�k�3�A� 	Y�ދϫ����pL��ihi�l:���^�ð��$O*�{�^�~�"u�SP�g7>�����~Mz�tXح�h,ǑCG�F)�uURWS��ٺe��1�N�:eB��W+����:u .8 �����a���!�ŁB�]O߀�VA�����Aą����
���!�:�ƁC�:�(�;�n.5�z����`
����pt�hc�_AzP����KC�a��y�}F� `
T��q���(�>�����\S��c�F�z��iG�5��ޏֲV�^tҼ�2<h�F)#�}�x�;��Q�3a�A6����[ �Wr@���C#��n�D�h���g���u�VY~�J�#�S�q�G�+�<䯍��!��0���]^�	�'
IO��T�r:��TK�fyt��wˢ&�`�N�"�mT٠cr��Po�vR7^ 8r�v�4����y�u�v9��.uKe��Ùv=2A2o:G�N+��䩓���1C>x㇌�i�l��\��b�}�ꝁܕ��x\~���ȸ�3��U��T¨�Y�l �݌�n�b{�8[�T�f����		����S�8�����$1��Q�ෛ���������L2MC������ϱS�[��L��&����7]<t-3y�-���j��q@�[�"?�pX�I<�b��-_����~HF�Ǩ��~x�h�:(�ć�M
�v��f
��#��}��w�V���0l�����=h�bB�����GD<��u�>FSH�y��)���cH�(�C�����e:����;���낮�n4*�(I� ��M����*9��8��qNá;g&�*a/E	{�뮏�+ ���P'm뀧Ha7K�!�nt^�F�4��,��S�9�Gۻ�$Py�!bMNNЋB]06^�b��O�DF=��H �
�u�uR���ʇG���u�6��ୣS6yD֬Y�?�y/��靎���7�<��߽s�n�.��}B#�aC�O�V^#��^ѽLs�?úb^�,k�̡T����b���u���ڧ�~�v��`����1���#ɉ8l]7K	��'��U�@μ1DUt��N7+ `��~�(�̜%�(Ӱ.0&�Dr�LΩk����o�1�<u�i��Y=�'�2S����V���_HldL���;�)�hl����%�d�S_����9vڅ�%�"fg�)پ�5��z/(,��\<������a��%+@
u�#xo't��<\�2��H8(Y50����@�٪���Dc#$��pҌӤ��Z&��aoU%�^�}T �2�i�|��n�dj��^��%��ƘZ��� #4� �9�*�ON�x<̑;�� �b�4B-KT�(fV��F��v��y^�7��o����!S�?#�/��BZ�zmPT�wjÐ5�3�xy��z�����%�F����=�
���K�a ��>���%����Az�H #�Ȇ4а�!%�<+<:��]e��mL 쑓�����z������7����*Lcׇc�@C^��a�l�ܘ;�Ɏ�&Y0�蟞R���� ):��v}��.�<��� � ��.p���x|&��R4��o����/�ۿ�npjd�Ͻ�wѓF{Q�s��:%����R��R��F+Hà<np�_��\q�r�5W�e���X��A�|ꩧ�5�t�t���<�?G�[p.�" _^8	��|�d�z}/ۼ"
6Sc�$'�RCI=������U�b�2�>p�W�mWcb�<te����,_vA��2��� ze���M��K)� ��-芻��\��d9K<%��0̉&Qv�2���6��P6T+�^e�c����µ���cV���<�3�� ��R���w^r27n`��t���И<���z�4��ཛ�9A��x�)SZ��7HmuD�͛��k�@A��;vJ_��ׯ��B5�)I�n2I�V4h�����<��C�����5�w�e�\���v�O��\!���#a���Yo�H0�q�|�;ɂ���?,##C$��E��V��P{~��W �n�*�<��Qq:���p.'���Y��ϮI�P��t	�"��n4�ry}+Jzl@:,�j�L�"ߺ���^�������i��{t�y�M<�enJ���(��)���g��CZ�J=�^B 9O���A��xh��|�5�]E���2sTo)��>��)2g�,Y}�
�={&���^�B���?��N5t��	����Z���Z�1s����%�:�]�_�NG�����t�K<���S��JJeT�y@��s��;��1��
��Α��l$N�a̪p5���=N �&�P`+2�ij��7���8eH��H�� 	����S�Г7���>�����l�lPώ�;F6c� 9@%n�q����v;o��z�*��x\�z[�������z�	���Ua���R��x�(���QFV���(=�6P+�Ovr��
t�\����Y�x����[���׍�@��dg��_�9�R���+6�	O�%o����]G���'���X޵�g�i�8��sZ��wpxHR���!=���˴3��5�ՀH��:9��بz��I$��e
Egҹ	i4l��FI��(�z,;�Y�yA��Z���9�Wa��9ϒ�+�G�cr�ĉ��=�p��D`�y��>��>v�sy���Z>��O�qYE�fb2��b�!",�� [(ɂ�sdZ[+K,s9}GC~iW�*61�?q�7w��~������|��W�{z��2*�<�
�W�9IW6�t�����Ml��Y�{Fg��s�)�6��9�َG�}�v���<�65��u��r���\��}��YR�P/�bU0��i�	o���$�
�)�}�\uܬ=�qMim�טͨ�����!e��O/.�𱛜0��zp�_�PAtǹ�PF5�}R��/��^$�-2���ǏQ#F<;�."({`��z"�*{ո;]`x.˻4=�kk���GdӦM�� ��b1��9n��F�^9}��Qf�5�2����`��c,&�>��!���
���Z3�]��ᱳ{X����!֖������a�Ľ��@���t����"C��{T����������=�,ǆ>P��g �`�n���K�y�yH�xg��������}��3��:�IFIJ�3  7�6/u�N�4�k�e��7������tK(�����,����~5��̚�������e���a}W�f���E���q���Rэ�G���D���9*�^�4��#\]Ŝ9�a�E�0��eXx�����W�^)N�S��W˚��h�H�"��ӟ���?�u��,7��nz�(�Bx���Aw�b�{� ��۵�بq.l���Px�ؐ�)�;������gJ��3`���vK��_���(�z��W���/c�}�F}��ԩW��|`�OH��`L�Ũ�=�B���k�j07��@�A�4 y�; �z����T�!���CKK3���s�4:��bq����J
�t5�z��G��24<�P��}��]TO��3�2b��Q0�HQ��a���5�:���,k��i (� �&[�R �K뻁���zy�R��T:cU:LH�J�%g�P6�gmK�ڑ4��c����ߓ�4S)N��T�;������u�XpJ"��-������#��)��l����9�tH��q��T__k�%�r�UWHuM��IFr�	���J��.l��S.��y�Oˑ�G�3�
�W��@��s��ǡ��^*���#�v�*je77����n4a��z,�p�G��;���-<6X���%�d�?����1c�n�Ez��O!ת��*��ɶ7j�\04"7���N0�ˎm>��|���!�"�@/�z��ЎՍ2-�>�o��-�}2w�
)�|�+C��F-K�����a���d<F���t�5h������$���6�3X�g[��-涇B)㡎x�lx�$l�r������u�I3!��[[�ȡ�G��� 2�h��g�NHUu��}�F���/��1���p�H#,_C��[�X�t�M�w��ߚ���:eϞ=�O*�f$��������uAR�n��e��|AFF�e񲥲h�Ry}�>�%�H�$����|�h�w0�p> ?J#C5U�Ԁ_�����AV���(��c�l�#��r&�7�#�]wݥ�Q��^}����ʈL�|�Vq��A�B]}�����i���&]�2m��3�E�9Cv̢ٞ�P�[q�R6��vJeT�y@��s U�'<B�E�[�p^~y��x}/	\��;d��7c���v������m�y��C��=o쓛o�Y��Yq��?�����I����9~�(+{��{�f�]^���6���nɒl�r�lp��n�MK�InnnH!@�IB�(	�H��ĕcw�"[��Q�hz=����w�����?�3����~���9gw~�k��%�;@��T�e��O҈��� C�< �R�QZQ��(���icE�T<�2�dϮ��w갸Q�X�Z>(s,�T2MvC�1��(��]Ft_���"��ֿ|[~������>K���&�W�1m��Q���F3� U)�1�k��^c�1ӌ�Nv��n����}g����0���"�0�˞V�?��  ±�y�ܹ�t����ٲ�*��_���/��;�����fd`pX�� q\���<��ȩc�lIus���EN��!Ȧ�cӡ�@��K�}�(f�;fϒ
f�]��LJ����H${ʵފŋ�����I���k8���p�y��/T�ӄ��[��3��w�&o���X/%u �����o�o��5&�ᄓY��d벥dD)e玽z=B�v���<cA�i�̞�)�y���p���y� ���%�Ѫ.�^�d��	]�P/�	f�W�X�1���!����Hg����P�p�<*���g	LX�1Z��楛�dp`�$1O<��<����ls�tg'b1FQ�F�,�H��tՀ����Op�Xt�Nh�|	�f.�Q�:���#�f#�'�o�
�.u���@fh[K�v̯�XR��j+j''���9���g"� hQ,������/�G���g��@.pQD��;ƺ������a���'>��)��q�=y�)���F��,���;���!�Pmd������w����;��F������}r��o���w��~`��׼�g�(G#�`\�F5J��E-���9�';v�欶�rIL�/�=D?J!x.�͛C��i�|`kCV�\�0�9�a������s�.��sX*$!�S�͍R����䝷�.�#Cr��t�>%+�.������R���'��,N*�$�0�!s�.�#y��af>��I�y��019!Cz��L�&b��λ�،L��Z.U=��]wJT���e�t��MH֡��-,��
��+h �C`��E`�h��'Oq�F�۳:g��3ݜs�xQNh �l,�b�P�c�R�ZE0�<���+�a~��5B"Mmr��q���#�pԤ��9�@c8F��ZJ�����j�d��Μ�%x 
D�5�����/���d�5�vq����-����=�|�r��w�#��k��NN�� K�jS�#x�ǽiTcFP>@������)�h�l�>�<R�h$�8 ��}GHނsQ0��MO��kkk�|�C����wHqrP��~��'6]|�l\���g���G�H��@y[��;fu�r��'�Ͳj���$���`��z�i��Iw�)}^\Υ�Z5�ש��3�R��Mfk�/<���WG �I���������z�<��G�'�ʭ.^�@��I��L�NW��d떫����òb�J�sDc)�& ��R�	(��څ��۵}���9��%�=1���ԂLՠ�y� ���E�9����뢚#���ji���QY�d�Oh�b
:�]]�LS]�yy��(����_}�e�Νr��k�N��V��o�^>�������������
E6�!U���Q-�ϧӣ�M���ӊ� �;����N�^�n�ē)C�}t+��0�d�"�N�Mi`��mDA �FUNd��yT{�p�juT�ə�dc0�����o�Q?_����OH^�)w���r�Iֽtx!��c�ǟ|��e-�-������~�C�y�,Y��Mz�;��x\�/��/���fy�Ձ9"��ڢޏc b��^~Q�>&	u(�u�Q��y�0DB
lW_%o��f)�)U�E�ɏ���ޓ�J'��+.�+��T��:"��qM�<����[n�����t8.ڴI>�7#��x�Q�;Z�|]z�&ߊ%K��_��|��T�;�۽�-��e
�;�T�!��nx������>c��mo��(�앧�~R���HҰM��OL#dF��Β��v�:|�NԜY�����%y_P"@�&�I3ˁ����4�������A�a�,	�_8�~�"5�ŉq��w =�Y(�b��Q�mLCZu��%\'5b蓪FX�7��Ex�4*�  �HfY�r>w9��,����+=���[�[e��9r��I���2�B*�)�֭#���?.���gYƼ��7�\�F��t2�D�1a�b�ۚ��o��Ψ�嗷�O�Sը�l�P>|X�{�oˢ9�����{HFsy�i�ɴ/uZRG�Zٰ�B=�a�;#�(0�E�B����G�f2�!��q�R�@�{8
h��KLuh���Q@����&��zdΜ���
޻������.�T��O?,��ֿȳ�>ˈ{Ӧ��7���O�3��W�{��=﹓]�]IƓ��ϗ舁;=�2t�}��l$��@u�ת��Ǡ��l�H��h6��^�QF�W^y���'���Шދ��eP�wǬv�ù@f���tZ�ڷo��3�k��2ݒ��t��3��}G\u,P�)��G̔����(`�WOc�"*M-�
�	鈵ˢ%�J2��}�ꬡ���B�_2������o{�:	o���1D���u�F��1���-Ȇ̟�rRkK�F���hLv����@���j��;� z`3�����z��XZ�D�����v���@zߩ{���Y�FF9��g�NΖcj\H!$��u�]t���\sYΞ~�iC��������i4s��7����x�a��?���LoZձl6_s�{���5�b꾜'hΟ��)nl�h A}�ca��F&iu|��{�M֮X��\Z�.\L5�R�0��p� h���Fd���0���HԑD2BSS��_0��k�g����`1�$J8ac�H��;jq��})��s�a���b!F̔��e��R�̙��}й��3�ŵ�l��T8����)t��#`\�b>G^}|�\D�C��ǏvɂE�%��܋�	Y�p�:M1�3:��}���:���������gg��ػ{�l�t�<����of����W�ftxX��G���˖������� �Ͼj�G�Ȣ\}�՜?_�z�̞޳h<KH�'���#q���"X��{�Iu�z�<�[��6���H���� ߩ۪˴��C8�0wN��W���H��>y���e��#z`��(�SF�$*�{`��@l�(�Ԛ�ܪ'�g�ʳ�|��2h�C��������m\ ����ܰQ,bc�ٞy�{����4^*˷��H�t���^6(�7=��<�HE�d��5�f��t�֍��y�$/��]�ek���j���)�jtC������/�$�/X+�M��F��w=k�/���/�U"=;2��l�,���G��+�x GM�#u��-���8���
.+)h���=F��3� ;�*�ؔ=:֑) "zň��`V+�lRko��hl2T��,S��&(�<�0t[c���c��P`^����N	u���AW<��\�� �1�1�>uZo��K��n�Ɋ��HGM$�Q�~ %�2��Č����/��N��?E ���^�:�#Qyeۋr��G�v���X/�dT���Y���vKS[+�o�م��F8_���S����C�ɔLf����3�P�����h�x���c,��*m{�En���`�����ohh��:��x�2�ݺ/��ٝmr��O~�l"�����g���@R��x�������+ ��Λ�،�r!�R�R�t]W��t�8���F�'uq��4�� ,��X����m W&����(]Gh�G|�T0���S�r�`TŐ�N�������o���R�������={X���Q,�ѮF�al�5�iO?��̞5W�{õ�~݅윏+p$��F8G^�	��g�S�dǞ}�J߰�"��O��]����ȏ�޳S),�#�>6�MH�����Y�x��UKK�d�\3�gv{��K�T���G�/4�f��u��w��9l̾�Y�4��HA�VG �Qu{kIt���ǥ0����80�U9
�Q?�_�T�nz�IY�'�idȈN�WxL�x�F�)uf&�`�PkBA3�ǎsU@�;{V��eѢ���ϫc�A�8 7�t���9:�w�D�Ȅ"�T�h���2�ɤ����qlom��:|���D����s �t,%���作'�����hw���Ks]�6ކY{��~dǳ
�f� ���A�D=��!���R2=�ْ>�!���J7���䋸�)��-��$�����3�<)�����X`��@lF����!�C��(G�V�hqb�",n����M�A��8�p��2�nbjML���-AI,j�سɇ	���U=_��B�rPu�icX�.�H�N(����r��A�m�V0h��@F�o��;�ˈ-�J�a�7[����G�~vpD����Y���b��͌�!*S��n�����	���)�����PA�����`�42H?�,��J�rd �����T2���Q�f*�\�r���(C�u_d���Ld&К�v1��������x�N≌O}k�=R���!����1Т�,����z�Ca���H��4'�9�4�+���/��o���w�/���D:��N/�ߢ��?����@^���?G>j�(W�,�雜dv�����E��욦8�;��%�#��
(�5)�q��1���f�h�ٔ�3=<�L�0�����J��ƱD������3��>��;."���v<��8�"�-TX��lsk;���2�>}+	,��d�6#S��WJ尥´�� ���X ���ъ�.�0�-=�ioD���f'�.�!�����oh��<F�%/8��@�	Mp�yc��\9�9<8D�EC����B\��Ƽ�^&f�*�J2RΫ��ՅuiS{�2�M* �wt��<���f��6�����'`oٲ�s��
���jt��#c8p4�Ɔ�-�SG5µ:�pF&'rr�W�]p���wP~��g-`0��s$�T��C��c��)�#�����g�=h���,��U���m��W�(wͺ�(��XT]�r�@�F��F�h�{ߝ�+/�,g�X��nb�]8rW��;{�Bɏ��|}P*���{ꩧ�ȱ��ַ�C��[`������]G��x����b(|��ᬠ[-�秊Y��,w�^�&��9р2�>@pH8g_(֚���+�k�i���}�x��O
<w+k��*x�"pL4���>���${��(�Ye��+K2����TM�d:�X��o�(�v�, ��fdCC��
�q�+�P[�LfX�h �I�`���"l(�!�I�vGC-���[q2��J���� ۙ�"����Ξ�ś����t��ڌ�щ�"��S��g"��R7*o���2�C�skG;���5b�(��ϥ�t����avm#���F�C���P��B4�f�J�#�Gz}���,)`� =��������/{õ�ʃ=$�3�^�n<i@���-x���y����=^��-X�Q�$�/��X}���)un
����)�'�7\'M����[���N��z��-$Zٻg�i���qL�ΐ'�S؄�>�N�m&�>3�:�����_�lꨞ7���ٍ��&=����%x�9�� u
Ǥ�.]��ԁ����ۿ�}t���^ukǃ��=l*̚�U�|G�R[ *��GĤ�j���ngt�5���:.��xNI�k<,����v��(�d��<��n�6#IV*n�\�0��t�0�ѴƨiPr��1�����uJ]���M1>|Lf'��I"�t�ˆf��c.ӹX4Ѱd8�#,ܖub�2�h<#;S��jHas�M#�R�8!HU��w��Ȱ�-W�g�Y���m/�Ky�ؿgwM4)al��l�ȃ>�q ��W ��k6g�K��/��'���y�3}��ժ�Y�z4��I{��2��"����a���K+,T+�b@].$�C&B�藠�0��qT�|��Br\J�b���7�ճ� �Q7:����2�S�-#C^]c��]���CC#r�=�2������0Rfo�kt{�0Y��9?�7���c����̀�T��D��e"�i䃳X�j��mæ-�ཋ/�X����L�O�R�9/_f�$ �B�sd�@h�T�!�q$��@�i{/Z�s��4p��I��7D����%��� �;� z`32]��p����d�B��� �KɊ�
ծ.�N��Ya_Y,�Q:@!�Q9��W�Z��cǎ0{��A�@�>�@ي��� Q4l� X{���l��`!��E�Z&��E��j�k�<<2���)z��F�Jc'9꼈��	5]���S'��g?{��ph�CP	B���~���|��G�n�� �����6>c"ư�@*�?��qޘ��3w6�p`PC��Z�[�&�n����v=N��"c_*Uǌ�پ�7���`��`�|V{��Fx̨���U��� I�7v�}��_�'ٽ{�̞3�]���P� '>�讟cm�p0p����@F�8�+��L�9B���˧�kg�f[�S����ŀ�����)X��)���A�)P�gY�l��L��w<a���P��FB�?��ې�&	��*�%�lh��uB���F�#_��FB!=N)`�y� ������"����>v֡���夢�$u���ʦǙ��u贂ʻ��n֣1W<11.+V������ޟ�޽{#F�\�m����<^r�&9}���BHD�8�Ijr��F�ji�*S��.�K�[A#ׁ�>ٸi�W��(v���|�{X��t b����u��O��]	J��3��������[�4� D� Iht�v�yp&p>P2kЈ
h(?��%��hif��sĈ��8��Q��9�s�(�R'L0��:L(`��k06�K���t�4���'?�)�#T����e��E|���ַhT=���{���*]4���D��O|���3OS�i���
��V�<�c�RIa"!F� KL- TAT�h `���=��1a��U����8w��H������F?[ú��F>��,?�q��*���/�k�
���e��&�xt��@��vuD\�~��I7$d��%�~�ξ��q��|�}��<Jj�T�EܭBAZ�=1s�v�, ��ffUÂi�h(�8�"M-���x&B4���Z�X�E7�9b���N�x�F]w��CFTH���> W]��ihHt�s�h��&�}``�@�(z*�77�5noF�јQ�#0�3R��6I���.��-;F�,5*��l�
��z��F��@���wH����ui���{@^x���C��n|��K���u���Lm�� kP�^vŕ��1�#���?�q*�}���y�+��/�h�8���+]]]r�eW0�],�(��	�����E6����@��ɧ���'N�m����/|�w��&L�669��W�D�z�GDv"��ǰg�F�8p��F�?F�j�|��g������|Ե8>�;�<ܲ^ע��1N �3<:h�>�
�I+�cAc$@d4�/t�{b������խ s��J|���]0k��q��Ȝ���ڌq�3��c����|���38IF�7���W^*��. QMZ��&S.�喛�s���<�Գ̮�A+�X���;O z`3�H<�4�5u�pu�z��Y��s��ֆ�ܵ�M_!��yaID#��~��y\���A9t�^�)_|q�\����k�5d��Ms��t�",Dҵ�d�s��E, �V��n,�`" @� R����/VB'���b��n�rG1�E�s��
h�bW�;���L����A�u<�`M���n[�|�H}c�d'r�\�I0@�h8�f�əguVp~ ���p��?�����-[��\iZ#���,�L"q���(�|�*��#Z��l�T:��o�f��]%�e��u���Ѩ:_zݲ�㤾����e�~W��PP��j	u��r�	6:���=8f�Sr��έ��K�ٔ��76�U,�~����	��104�����ѣG����@V�^%��M�����Q���^ɛ}�g�զ�A�J��\N�OJ��(�'>x�� hl|X��8%dA����$_��7�iA��"vʊ�K�h���.�,͍ͬ�GÞ,Y<[>������?�}�K8��E0�[ ��Ț��A�AqԸ=]��Q^�|�������PJ������}���~��jݩ�&lQ�C
��!�h�QbwL���Ozщ�1FW�H��Q j�gVC���8��ś�G�,(X7n���jH]b��8�T�Y�.��9�5�c�l8��!n"b��O%R��ҪQn�������؈%F��4�Utq���?L����o�\�ϛ�����p�c.\(����$��7�����%�6˩���ǲ�+�myWD�W_��b.��d_~�ev�#��3g�����Qx):\h�CC�Ui.��靀�y��|����q�Ӣ�k$����s�������1
o�ZF�dULD�s�1C��{�0��;v�`#�W\�y�\!/���+u�[�x-�3<ds0Rȉ���l�3J�9u�����2'(���Y�t)�W׉�����7^w���'?%�7n`drb���p :;gK&ݠ׭�P'3�)�\��g>��w��/ex��Q< ��j`��@lF���G"��F[��"-͍�b�
��+�P#"qȢ%K�����~��ӟ�������7t���۷k��jX)���aini��{�����Z��멄�hż��ƿEfЉ�� "��e�]&-�h�)����{X�;;��jGY�'���NNL�.�&),����s��~�UH�L,#xW#��$'l�'e��Q��x��$	D�}g%��0�1�q�~�6��8��\V�b�̞5� D�k֬a����i���v�7!��kb�JP�X�d�tΞM�ji됵n�,9�߆�F	��f ҆�=F�|�م��av�Á	�c��#�A�E3�`$X#��2�X�k��o�F�l\��{���Z�����H���stv��~v��C5<8hg��z�8A��~�Y��7^�^.X,s�dlb��hQ�=j6H�6��R�Ѩ�����:�[�v���=æ�y�g�Y:~��/�%h�oVǲN2�zO�;;$��#��>�A�K%}B��\�y��^�V�{�e}�J��a	,��h�6#�帊�ꢹ�!G���s�:�Zo[�,�5�i͸�_>[Tp�S*���G^y���.pFV/��`208L�K��$�	x��Gt���u�XPmDgǘ�Dgk�
g�_q�Ul;��+Ԯ | ,��f�/_*�W���k�ʡ��9�擺��Ă�Uy3%F����bDZ�Xƿ���nے� ��-m��1�~`D�VČ�g��� d\d�q�9�t�M�<�ϔ�^���z3�mJ�Z�o�F�n�J��h�x˛o"�;g�Qvn�#}��uj��^,�!���F�$/�DR�dC�/y8�d547q�+�����0��{
p���6*�cy0�+���8G�F � F7����L���絏����<�C��Oɺ5ȩ�]�6͎�`;6��Ʌ��:ijm��;wȏ������[�T��:*���o�����'x��r�lq!�a�-������R#����u2�s�,�?O�Ι�N�^_=���V�cO<�RR0��y� ���%҉�b1�WT#�ʙ�%���.M(�
)���)�<9|p��\IS"x��}���e��92�8ñ8�,��I*S-K�3jW�FG�����;��)xl���� �u]���9r��p :"�|���x�ʉ�,�94�%��it?,q
��pv�Ԙ��?�t��D'��Ҭ�.�E����:1����J�ᣣ�2��Iƣ
������a�H��8���GĈ�}P�r4���?\GP��z��C�)r?r�#���^��78%���}\+��q�t�[�9�밀O�D�N�瓸@�!�>;S�јߠFAF�ǻNr����(�Ȏ�+�s�O��6u�&}�N�͘��2R=�}��ҷo��R2'N�6Y�f\�\k�D� �=�+�?�{��!����&9����#�dr|�R�84 ��&u��&�������L7���P�(�DF�X��5��H*��?%��Σ�،��º�c�)�ʙ���q��KǏo�:iji��0���L��9g��Ѯ�
zI���7�����[~�ིo�.M؋��5�b�̶#�}��eժU\ı�#�j�1����L�U����h���]{���X�O��0��4 Q1�lk6���Ƚ)�9?en#N�\g�O�aCւ�����|@�Mt� ؔK��O*��s�.���q]+
 l+���[�qb�+W��[�+#w�v 0�u�i{��V�e0U �Җ�V�(ͼ<�gѩn���Q3������!S$e����IȚ��F�k-������q3?ڷs�8vԶ�Y�q���ܑ��M�}�������b���;b�����}}��fs�ф����P���O.��b����:O���̓Oȿ|��2:8$�	Å_��I�������#�Y��T���g�_o��ޯ�+��JH�v>- ��fd�C״� �&��E�� ���]:;:�(��94�/���e��)���?:��)����F���rՖ-� t��m��k���G�%IɄ?g�IQ�J\H�����ݡV!��qp*ȴ��@���ܳ[���J�mG'�b>d9�6vz����=�?�]���V�&�c@��;ߦ��;��F�9���Q0;/�� ]^e��d?�4:D-�b ;�Jc�FZX@V2�xz�rc&��:�""Ih�gsct�%iI#~�]�U ��q�r���c�ۙ��.�B���G�C�[�����x�-p)@×�fY�l�Ť�iiie�:���T��Ą:g���d��z\�a��yWMt��Z��q���Эٲ�uĬC�ϣ Uo��6l� ��=�vJG{�\�~��~��T�{�'�J]Z�����i�l{�9�xQi�5W��3��G�h֬&=�F�:v@Nw�D���!	"��Ϋ�،loqĬ����>i�kT����I�?o��s;e,�;�N�9�߼��|��o��_$����P��x�ER�Jj D~�_+�J�kin��E���`xޱH��cIy�2f?��3��*���T6�G��x�G�UC��.���>�N���lԎ�7#t��Y����������L�S)k���k�7:6̨]��=����T�E�H�'ň���Fi�49R��M�{��Hۤ�I،�^ !��k���3�NK�١~7�Gb����Z��#~$TeD�T�+�XF�:ȣ|���:<^864�Q�G�q�ᘠO��Fr=0�Q�M_p�U��8��x$���ɮ�^�����V*���L�>�{�P�5���7�s��/�����Ô䝫�W��%�|�e���?ȴ��c���L�َg�~B2��|�B}�]
݀6��{�g�����u{M�F�A�{`��@lF�'���LV�h���Wf�u����ua{A�����HF�ޓ�9u�[z{ �bɕ�ƸLd��,^�X.�K�E��wJ�H	��tS35�㺐C�
فx,E��2A�
pD�gN�HǬNu8b$q��H=������qv�[����Q����6	KE#ّ�A֏�~'=���n�vm�L���7p�cp�[Ǡd�:!�
p�1�8�w}j\|����ıcSLx��6#p��s �2���>��O�;؎�7�憎����w���Ԩ2��T#��0�v&�����%�/���@�����T�R%c`��g!_�;م3��vg�nF�@�K�w=Hp�G� ��!`K�p��'�ǃF@8^�zߠ����45��:F�=�H��=��K�#����:���I�+7�)]�A�b� ���W��:ҐNq����I���;���$���)xp�LVdpؕ��Cr���'�b%O:ڱ�Y�r�t���}w�{��~�+�L���"�h�̢v^- ��fdH�c��^4���i���֨k��6čhD��?,'Nuˮ���%�8fa�XcM6s��Qmm-�JӺ���9}RJ���ڕR�F=
gs��P��F.[`g4�ЬG�����N�l��j��>n';9�����q��	)\(~a~�z�D�!'d��9?m��ac�F�F�ly��C����{��� %# �(��(��#_˴f��:Q?�?��ƖX��n�|x�~�h_Ɵ���������k=I�� ��z"�s$�o$j�������y���|}v ;+65�3�v�U�̀��QN��b�����V�lN<�H�E�w�pP�COz)쬿�cwL��>��X�`],��<��:&C��㝷��D(��D���!�T>�-9u|�oX+k/\��϶�6I�d��<����O>��?��9�
Mq��_ =��.�n$�J�)��ɢE�dV{�<������ə�I��O�<-ǺN���S�i���WdY�t�����M�g��L1D@@��H��F#���@n�^���m��#��e����9��0"��:
H'�K�t� X�� T�Lq��5:��4���;D���6�f�9\K�㧕s���tN{�3�w<;�dj�7E[����H��?�����9��Ba�)�ӞN1��LՒ���j�Ŀ�M�-3T	�"�B��T&~���;(=W~MӠ�=���7U�0�X�� õsxw�s�{��|(e45�1"��-�XJ��=ʶ���^u(c<a�q L�#o������[�|�#�D�q�LNN��a���:+!
��!L�vFF���/�ɾ�����M���S]�r�|�u�j�Z���>�	'	 =��j�63�d�.ꈌ��yK'���=���9]���;$㓓Lk#
D� �(�����(X�G4:}ꔼ���f�Ȃ�c����h�6	�U����V�Ԑ�Ge#HD[͍����MG�>S�ȟ�rA�X���:��D�$b�>u�ѻ�)E��F�:\6|�Պ�+�U:�=��khF�"M��o[���*?���@�.�*S5{ېW��ᩦ3oZ����v�Ӂږ<�ٯ�x^�y�{�6������)2,x�=��I,E'w�Z�97ix_ͧFh�#�W�f5�؟�F�8:ɻϜ���3��gL�:>��Y6�g/������'��U`� _A���F�r%9t�0���Q�RH�o0�U+�l~,bJ0_��Õ�l��� ��#~��/!��d��&�ʉ�O%�RSSE�<Z ���R��W�H���ȉ"}	 �!uM�L�W��X4�su�L��k+HN0�v�����[��K����n�F��|�:����ҡ��<e�Bm�f7�P<�������.:���E]�Z)I>���ա�7o��k����˦��]�6]N�r�o~c�6@�ejQ&^ ����(3�N�C����S'O���5���R�w}t���Y�LE�qǭ1�M�اt�Q*`��wl-ނ�݇2�u[�R��?O�7�?t�c��a��Kg�4�a�5�j٨��Ke���pl���D�L��@ �a������`��H�����ζ��GZ;ڥ.��x��tw#y� VJE�#G\���H��O"A'׳PD#�:%�D6 ���p�1�������pF��$�T0�)ܫc�ⶠ��wBz��K]S�\q�r���J�ptx8`��Z ���<߰�S�\�3=g%��4�͆�#��<_��HVFa�}54DO`�����x���w�n�S�N��m/I�dR���"
T�RG��Yn9�}������uȩ�Q�0lk��M���g���|� ����Cۦ祝.��̴nؤ����z���87:fu�t�_{�Vy�;�i��:�Z����G�0�aϝ�"Lۿ����3�^�iۭu�O��M�[s<�������ۧjZ���q���5r��1Ϊ�9e�M�4���ANS� ��.���#b�G��wx k8���8hj�k���P�9�r�؜e1D6Q�pol��{�$9 p~x6@�GұC#���!�rG���$�"�-���̠�M��H�4Sz�9���
�"�t�<Z ���tw!R2��$؀�`�m #�Ʉu�2c/�g!JtB��q��K����{X���ҷ��ݜ#�:~\�_��ɸe��==-l�ld�mcp����9�$�W8� I�5���:$PI��+;�gf�c��\բ[ȃ"3�?���Mrv�
�� ��������9����-�/�@��j�=1#j�pV"����&�ZT���i쐿o���o8�3��ͿW�ا�w���mo�řj���1o6fF�ʮ�\�F��	���7������q�11��a{~6mG,d�~��U���i�33���r ���lDVpM1��h��襨�i���L����l���Ƕ����\�Z����Ï>B
ت�k����J��.��O��r,�]q��M��#�{/�_!eHs �������D,�d�yJ�v, ��fd�h��Q�k�(���w4^b���bf.�\��J�0�Y"�&jߧO��S]�j@�H	Mq�G�2�k#-X,e�Li6r�Q+dDY1]lQ@��S��5�8{D�)I&��W#b�À:xq���$�qw��D��#_̯�4r������7\ô�U�u����~��W� ���Fʵr��1��c�՟�ׂ���{�]���n�~�WA�=WD�ֺ]j��O�z���Q���^]2��l�9��L9�l�
ƒJ�dN���y��r<Cy�<�+��fA�d�s���Y�>�'o�Lc�>K����;��3���CfϞ%�����5��=�W\�U�ʜ{�����t�8.�T�T�H����Y��"X�8���X ���(�yX���Ff�b-��B�E�R�0C��4��,��7j�X��Y|��j��[���X@�X�́,�1��v8�QWQ&$���1@g4s�Lƨ�� �e�R�&{j��g�^�;����S���g�P��v4��+6˭7���qP�{\�E�g�KP�{��6�`���� V�����.z{m,`Ow�����������s'&X�b�Z�<f�m���-��8���M�䑟?��r��W�Ow[]u8E�'�1s��ܔ�ƑAv�GQ`�{�J���>hZD��d�ʆH�ϑz�t�hjó���a�����H>R��q�m6�Z��=��}�k_��~���}�WL��;��/r��B0XR�D�
9��~W�P��o���I�2�܌���0���2���I�?����b��Ϋ���,bF�F̑ޞ�(����D�a�?˺C��F� �I�? ���w�ٍ�TqI S� ���
Ivb��l�s�,]_'!�8W{��TZ����`���G-0C���`q�F�(�"�F��&����q<����˯H�0��������\�����{cS=S�P���'k3�V-cs�����,;��f??ޣ6�^/+�j�Ѧ;�N�ۺ�t>zkv���Lu�ێ}#O�˒:q��h�V6�&U�Ow��Z ����,\(�/��3�j8lz
�ZZ\2�M��|����x��?���x�\��*F��:G�N�v�����q'ҖI�u����]\�={�ș޳���{hތ�#��K��gn�����?)O�,�q��� Im>���W�Z��x��G}�5����.���ff��Q�T��1y�ѧ��--{w�bV(�#�ck��W =���a����MB�MD� ֤.h�M�DQ�����$۪A�C=#G]L#�8շ�
 �@���/�u[�����j��(��?~�s���Mr���JE�r�Lǀis�0��n��c�ݭ�"SɆэ��@x���S�k�%s���j�5]n��8�֣�נaw��y�o����PgF����� �~N�js��D��?�O�eW���HG񖜡x�B#5�T���[S��WSѷ=ƨ�%ՒS)}F���8Ʀ�#>[�<��-���L����^u��޽W�|�tP"�u�*P��LyGj�	>�s�<Q�vdا�MRZ+��%���؆F:��H�Ա��9%���&���Y��"���sD��?��t�=� ��ٸ92&;��l�2t싼��l�J��n+�<'Ƈu_�i˺W���dͪ5�O�t�$%����r�ߜ�; z`32��mt�Mj��>%������)�H8&ǎ���zF���j)��u#*M+����|7�L1��}�$`#&��q����,l��X��1*�ܶ��I}�H�p	 �&��j�X#�aw�F�`%��Lj�/�T�d�!��N��ɩ�6��k���uމɱZ�7�q�h�)\�[�|&��`;$k)k�( e�������9�{��a��[��ULu��Kܧ<�H"Ƴ�~�N�E��$q.�가4�f�ׯ�E��ə���Q�	qR R�u8����r�#� ^8O�D���Ԯ���R�.������@����c�rX�y׮]ܯ�5�j� f�恟>D>!dG��<6�wS����J�B���`�
���&�wKʅ
����}� �����_���|���(A9ޯkX,�X ���4��*(zH��{�\-��.��K3m�y�fC�`��4��R����)T���dG.Z"Wn�*�����7�|��t�M��;rT>���J��DP���Mxp�/X�� T_�H� a2mt�q���,^�t�������Ia�gsҤ�A$>y�|w��]�ݴ��u�-�LT�i�3���F�辆�Aj�>����cA:ijl�Fc� f6�G�X�k�~�]����Uj�����5lR���sR���Lב�5ep�#­SP3��v�OP�h��2��!�t��r�7����Wޗ���E ��N4��:8xA^�����5�c�:�)J麔i�s��w8���~F�`)��>�Fm߾��1��wz�p������k�8O�#� Y��~�3��鹦eٲ�r��q�h�%rɦ�8��I7��R��{�F�Ey�{�+O?����mT�z��z`��@lF��R'+>4�͙�)�W.����ˢE(�(h8���}銥r�7�}�= ��=$�E("�뮿A��%9z⤬Z{�l߹��tц%7�R8�|��4�>��s�=��cm	�낌�-�o����NZ�6B����w�G�?�l�&S�c� Tv��!C� &�rv(h�B��$3��lm���}J��:14��5�`���\>��� �s����ݻ�G%@X.��2���ˍ��Lq�s�?�E]~���3ئ��jHhJ
֤��������ʎ�F�����v֜��v]�t��=���i[j��=����s䐲�H��}ý�h�qμ�����y ?�g�
��$�˂��4Rn��'�1�Z: �o�>���ޜ���ر.�(��oP^|�F�ǎw� � F]|G�Α:1P
#�T_Aڿި�G�Ƞ�_kK�r�f�jY�r���Lʬy��Y��g�����i.\���Me�^Ku]�T*��;� z`3��=�!������d����p�*}�"f�|1¸��tQ��[HOH��3~;L���	��7��eނE��?ʮy,�	t�W+����F,#ŋ�$
49!z�0̚5����C$�hB$��M�Y�B0����,]����!��+��+;�a�O��uf�,PV}B�W�M[bHfnٲE�4���!0�F��f;ǭ z�c��vף��}q"��jyx��~�q�߭|����h��'e���Վ���dHǫ�^8�p��#��3)eֿ=�n{�D���:��m/���H&�Se;;oޭV(�b�ma��?�פ���կ~U������O��x�t����:��dW�·���e���Y,Z,���_�f��؋�xC=QP'W���H5=l�Qn{�;d�%�('�♚��!��I�B3s�Β����F�d�>��U��ĉ�)�j˯X�L2uxvK�v�- ��fd���M����~��h��U��[��3�jo�d�|hdT�.[!��-���)7�p�<��S���П9�+<�����K�N7Ȏ]��n{��y,����KϪ�Ar�L}����9G��MN ��"��h�Fw��DZ(�K.����裿`ǵG��#IDr�)��2�'���g�Q| �I��)����=zT.��i�T:Ip4s�.	KzN tS�'���x�l&aFƹb�ǟ�Gk ���������ݝ2�����`K$�&@����tV8;����9��<����^������7�KˆQ��Ϡv���?��4��Ș:j!̅�Mͽ��b8<.��:�3a�>::&����E�vu
�ώ�4� �����t�Ѧ�Q:v܏#jHS���R��ԣ�7����<fu,"ndm ����+8iL�'�`O,���-0�E��>�=$�ioi5Y	�.��T�Ӏ���V��A`���@lF� P)�.�q��Q?�sd���*��HTi�"�w�za�\8҄���S�^^{�Q���t�Q���/]��3��s�ɀFg�J�E����,�UE�|�h_<r��ޓ���V0��L�c��olf�`iol�X]Cc�`���!�huwf�}�x�jv����ǌ=z��|/��jqgz{��G~.��.�(LT�$�.�|����n�i-}�w�8Vb#�CZ���v�8��^/P���l����V�̰�95���{U���O�b� 5�ˤ?��$-8.4Õ*�.�t�l�ݣC��ܤ�^[���B���u�<��I�җ�ĬK8��:'���� �h�9z,�be�B���a��T��y��
�!��#���O�����4z!:�P��r�ӑ���lt��f��68Q�̀sr���́x��p���~���gz����r�80Ep#8���f��NHG�,��3tx�N)�&x_._)^I��B)���C%T�V��z`��@lF�p�&��3 y��aA]�t�FJ��ؐe�Z)����]��*���M�n5��?������� r��-����QX������9qJ��$]�Փ���j�e4�Mcݏ�T���t8�}V�"�88!�� ¶n�.lvpK�6o�O��ͦ7',-�1d$:a�pL����1:�{� ������AQZ��@�:]4�z^ ѩ�T	�8n��Hd��T��L��̠O��ٚ8J�j��?�p{�n��q���]S�/W-�l�_ތ�!c @p��B�p=���r���G��ڥ�&B��Ma���U��;��3��E`� k�8�l�9.eg̍ӑL�`�l��X\��A�/�9z�	���>{�~��]�0�0`T2�ڸ�օK��u�]'��w�4���^�\n�p�$��_ٶ��T(��K7_��{?�>�Of�n�[�^+.�K�q�N�K&�pزz�y	,��h�6#â�А��4������9�۷o���3���{wm��QFg`QC�q��Er���u��y�oQ���'���|JA��QnXLW2c��� ���P��:@?�pL���"�N�|���T�%��C����( ��a��s����d{ӹ�Q9i��������}�s��ё!���7P/�!S/�z���m:��`�mz;g^��l��q��(@Y�s�֧j���n�pdJ}mz��j�}�����&|����9]���8q9���L���ҋ/+X��]�H�3�az��[ء,*�5������{��H&?�{ȕHL��F��(A�f��AD��9����E��p<b1�'��K�L�d�]�p�1��A}}����;�#;w�$MKc��O�2�����#24xV�]�Q�;�����ʬ�=�^PT�nm�%�C#�2��#Ǐt�+/o�����E��̚5+ ��Ϋ�،,�;������߳�]{��e˖��d߾L�R�CM��Iu��#�������� H��Z�J~��?��|H�;*w�+��}F�O��x]*����ڪ��k�:h��Q�:I (�ʒ�� �E��Ns��)w� �����8������6G�2a�:��(�*|�H�[�T���냅�ۼ�k_����r����0�T�q3D�與sA�.�k�L�Ƽ�����_8G�l�}J�|:�@�2�M'���vְW;��p:�B��P����ϙ˿!��+N	�� U���o?Cd�1�|���k�S�QX���m��S�MXډ�����^�:XdAP+GT�U�J�<&&&�TƓ��M�t���������>�%K�pt.71���sTK&S|�~��{���6Ҩ��u�>�2�s�dꥭ����Ւ+������G���棛6m�Wgz�%��΃�،l͚���u�~y⡮744ևuݵs��PPG����l����f�QA}�K/�7�����K2:Z���v΃#E���]w}�MK'O�d��s�v9r�L���9���hC���љd� z��
Rf�����D$-y���-f��x��H������r�ixx���x"�}`�'�jmX�K��L���	ՀRd�k�W*�\#��a��Jfj��%֫�l8��(\3������Ʒ��uЮ{�Tj-�^�I���;�:�Z�ݝb]�����Q-��	�K��ڲM��I,�โ�ݔ L����#�>� ����FTgHn|�v��@����SR�G�(8��ut���ߐUI���2Ci}�6n�H����>X��T�b~Xr���,B!D�h�;p�����;٣o �e�ʉǍ޻����3��9 ]��2}ԏ�%�\"M-m<7�����+_�����>
�3�f��ٲ��$��γ�،Qƃ>�����;�⪺L�yYS,�K/�����$)`A�o�>y���_>��rJ���������.��'?)�4*Z�b�,_�Bn��z�^x����Iʂ�(���!g15UCˊ�6K��Q��&"L�Q���¡*�h������5kY�Mh䅮�ɬFkn��OS%G-���T����:����� �]2���l.��L�|�S˹�������o��!�A_�Md�2���U�	K\&�*�R��h��t�2�o�Ng��/�Zc^�@n��	���)��F8&jQ�H͉�Ӂf��h�.(S�0}Pq�	2��s�=�Mի���S�j2aF]�j������#�[>�ֶ6"���t��}�[JAcu��A��Li��pM��*	v�eӑ�Ϡ!���<������K1���Nt��~��~� �Q�ס��i�n�7g�<��S�h�"f������!�ՙ�3w�w���2o���;� z`3�[n������?���?�D�P���sh����}򔴷w�R]�A���Ȉ�4�"��76�"�Htp�6ٶ��E�@ #7>�E�f0�\��J*��HYţ�&�C�T��qtbPRuW�g�K9��+ ��)@546QU,���UA�Mc�#R���㧍��_�
�0�aH3*����uQ�sk[�46���
�7v����Ѳ��Z�@3j���㧍*�XƢ�×UJ��,����Kv��;[����&N��H>u�^�Yw�������#��g��D�quB�� �e8MQ����r/���9��`<6�ȯ�GC�ַ���Fz������Ty ϑ���X�>S?��O���g�1��bp#8$���"�N��G��zN�Ž��ȟ|�stB,l�ft�i�����
�MwO��y�O�����#R���Y�m�g��~�������&%���, ��fl��u��.ң?����T��K��a����4�!��ʕH���*
�j�Q�m+W]�����nuu���,��&5�uˬ�"B-�\�˞��)})���)b�����R�3�X�Ou�&�p����(�:�t)R�3��E��[)R�O��K��e�F1�p����k���~�\Ʃ��M� Uv|+xP�w�{ $��O{>�����i�sצ�aI\㹾���;��n����j��m�lg;�JV�Lq	}O�Qv�á��u|4��c�F84�y^I|��i�f3�a�d@F=��c:r��>��8�b΍D���\�~��c�2�u^Y��;�Ig<{&N��=��d>���F�q�6�:NU}��T^�;���v���y�l���x<��E/��wtt���475a���hS>
��Rɑё�lGG{O�.�}饛��~�[_�{?$���d�v^Lޒ.�v��z������?~�]�(h����cq$��
�!��:�������A�~;_`�8YL�1�vn��>��Q�=C�j�H�j��`[�jQ����g�ay���Z[����3�w�́�j���a�T�9�5!-ǧx���[�Ƕ9���Wya���?���<����M��(͋�C����]]]����)p�1c� ǆj�� 4� }����~7�a~
�zn��t��6�ՄT¦l`f�C��z[s�����3�W�� ���ԯ86��ʣn�F4h����U���w/\�hG8� Y��J�JAtB#�I���!��!�*��H��.�{���P��P�sL������̏^�j4�`�>9ǭ��7�V]���\��ש�/��.����B�1�#�w�S �,��;�JU�W��Y��W���¥�>�au��b�\i�F���6����C�|�	�D]}�1�X��x����g��u��*��c�	,��L =��f~��]�?��o|�k����������D�p��l_G.���N$	�C�H#6ԥ���)�;�k]�]lO�h�O@��!1Dzۉ����,	���uĩF$�E4���w4BX����ׅ
U��x�^��1W�
�x*�wl�Ճ��U���rK���w*�P%R�}T*јƈn(��ʕ��g�Rz6����D��.[�d�����*�X�钦 �D�-[A�F#�ʕ�Ys�g�����_��_5#�j�Ws�B��ӿ��.s�B�Ǵa�E�,�*t(��9,���X��{���o~ӟm��g��e��8N@�X`����y7�_5��<�C{�F���ϕJG�F���6V�t;�?6\��*u0hm@�;&ǎ�h(Qc���ӈ��˧�>����7��G��~��U�U�"Nm;�!c|�p��X�0�!�R������J��|�.��L��X`����kf��-͉EB���xn��X%o���Q��}sk��i{F�l||��G]�����'�P�&Qf3�&�ȜLm~ӝ�ȫ�.8�t|q��b0H�C�c]8�x:E�4R������`X`���X`���&'+Ԏ/M3�?������G@�i�CC5��4�f4.�+�j����I�[v������v�R�Nզ��H�X��gz�a��������P*��8$/K ��_b��kk�e�)��L�M�����cP��/�O�dR������CW��bӚ�~]=]���W:�CFqmz�}:#~�1 "��D"��d&!n(�NyL4�r9���5����� ��5��d�T\�V��H�.�!P�9jC�B�hHZ3F��R�Mgεy�r���W7���Qξo#u2�Y�ڪ%�)���`������ݶ�K͗�}�<}��<�t�q�5��{�- ��{����cc׏������;�hLfϝKu/�|A�԰�����z]C��Y�e��E��hH��}�Z�}��	Հؒ���s�U�]�a���	����8�,:�������S0�e�2�^x�#u��O��w�gsX`��f z`��F6�wf˱c�>s������-r��K��N��,��8�����N���X��S�H|���f9+"bA�Ε�q�)��W+�Y�ߦ)�ըk���-�ۨ���'�;`�C�>�dÑp�X��[�������}��7@:$��kb��kd���{�F����6]��K�7B>.�Qw�s����l ��E	�I��n͂m,���4жLu5~w�;yլ���W{u��i�|��m�� �棤y����r��ɑ��^s�X.����,_��^70��kd��kd�憇�\��7�4�Z���������"�����l6[� � ��R��Q�����b`�5������5�1ּiҰ���Ύ�Y	U�U�������ں�;;�_V��K�}��o<�_�m$��{�, ��{����}R��Gbh���8�P�
ʍ����>}z�c��{k*��(x�5:&%����Yـ�U�ZŬ[4�N(�:���z=��7d�u9��\�L?W��Q��/8�Nccc^��1 |^�6��S@�ONN�؎͞={��cE�t����X`����:���	}�U�<��������H(`F����� �|�cBg���g�LU�_#iVm�=��g��~��W�n����`X`�}- ���o`>��Q��X`��_Z �X`��:� �,���u`�X`����@,��,�ׁ�X`�X`� =��,��^ z`�X`��, ��,��{X �X`��:� �,���u`�X`����@,��,�ׁ����W2    �����D 0 t :  � B�����`@� 0 t :  � B�����`@� 0 t :  � B�����`@� 0 t :  � B�����`@� 0 t {uUcrC%%    IEND�B`�PK
     #{dZ�S��*  �*  /   images/cbf7ad0e-0f08-44f8-98a9-dcbe92af212f.png�PNG

   IHDR   d   d   p�T   	pHYs  �  ��+  *�IDATx��}	���WU}�=��9��HIH ƀ0�`X�������6���x^k��lq��`#N	�����4�h4�}�t�}�]��W��}�"^���Y-I4��]U����/��?�/>�y%*d�ɇ
�g�B�|��y&*d�ɼQȃ��$ɀL6#%�d*%	�"#��@��,�,�K�e2q�B��	��+��l6����@/#dzo4)Ch^ׂ+7l�|�y��'�=	��8�v'���42<�$&����D����fYK�I�0�l�D�?/ɚr:��:W���bP �d����{{���I�B**+�lU3އɰ� �)g4�Y3*)C�x�C�Ȋ$�U����J"e�#+J����YVT�٬��T��h�Y>H���\.�'�7
I�∄��EbגB62�,W�H:0����,Yrpk�Y��)F���s�ZX�`���}�
aV��<�J�0�d�(� �$h�3j
U4[�.���I���2t�Q(���s��T*Kߥ�;�P�v=}��BU�-UMe�'��4����lN$�4l��m44�p��9�N�������Y��l�>�$0��e��L�I�B�n��5�`+�)O���y��Y�pͅk�s�*� %���s��y�����$c>ɼQc}0�I�ɬE��,�"I�Y�!Y���D"!�a4�D���QUF�O������ ���^YI�|�y��_蘒����z��s�_Ba��C���Bd�����>#��j�)R�5Lz����ItWȳ�=�Á��!D�i��SD)�ww!�;J�=&i��0T�'D	ˠc����lk�� �b�T�N���'>�����`JnwN3��W��p;F�Kp�m��K�ǻo�����i�-�*�_���:�<gO�v�����sh�<�[Tկ�֭���x	�AF*�FZ�Y4�xǃ����0%|EP��]�&8Z��T�Y�p��N\RS��^�,f2��Ukq �A�>����Euu��c>}��z��
�XX���M���S���n�\X�~��+�\q�1��`���`����Գ�CI���r�C�����M~�������,�V��X���sp���^q�Շ���G�����wg����w��p<��������|�n�m#�*����	����U���>fYPӀg_x�&+�$ʊ�q����ƃ}�h�o`*�B�Yi��T��T:%>���l��S�
�-�/��ccî�҂��,k05>�5��lQ<>O�3������z��
	G��;ή�兗���=#��2��I���cA��I$�Q5A���V���U��"��!�cF�-ј����"�;�����cIS"4	�D�8|�~�������C���:�K��誐H\��V��w�K�N�'�PѰp	�v',d% ���VL����'q�qAͱ�C��VF.��L$��Xa��&���$�F�VÖ�ν�Ѕ�X����1�")���W��`�ؤ��� ��Ǡ���I�Y�A~�[.Eg� |3A�-H'b���$��.C���pm&���
��'�}DXGV@:��.��Y��gggdVE����LN���%��� 	���ͨ���[�?�J��T"�EW���aLO�`���X��2�W�a��V4-^��gN�Y_UQ�q_R���1l�(�� ^ӈ�b�����s_ɭ��5��ј�R����BJ�+�7<-��<��d�K�6�7�o ���#�矠�誐L� ��\mkkW'=����H�+��P2�F 5��X��9���am(���_���~ψ�fQ������.+b�\Ϳ�g00؇� �v~�SS��{�<�c~P�z��
q�������K���	��
���6��*Q^^��������l�e�K�3���[���N�?�F"��7��511t� �x\X+���Ʊ����Lk+]c�o"���'�xI���Ϡ���C2bq��Љ�n���0�������qb�cP�>���H�g4�B�gV�z�`���m.�+`-��,V�S@0���\�����L {��0�P�a���_G~d��_������-&��7����.]��)r�	r�L��E�4`
J+�16�!v\���LJ4[�X�%�H$���A�����ő��Y���9{EXE2��{a��E~������3��3t-'1S��r���U�%BY�L��
I�Ė����z�\RY����ӭ`4���]	�UX'�Caa����C�EE�!h��lb�/d{�gccc�3�+f�Y��f�2�����B:;;0�ϐ����~�xP?���X�6�.F+�P���ߠ��\T(�1����0g�L��AqY).l�)��t@���ⵑ(sVL�|+�-'���S'XJR�J�{�ɺ8���Ҙ�0��s�s��ش����#�a�?�B��PE���G?��}�LN�E����o�;��C�~,^�
}�=�������J�j��+`�!�_s��QgA��U����Aq;s�m��PyNY��Z��z��rhp�a$�-7l!�~7n����ص{o���փAo�U!6�j�"+F�"9q]�=4�V�-�F�@?�.�1�C0��$v�1Is!��`e��2X�X����s�:��}��4?����5
O��,6L�M ���`�ӹCO�U!�e�p��#�ۤ��;�v�����K����^*�¹D���2+C�eW��VCn�	b���`1�g���gr��{0\Y,��0�Mz&��J��T9t�,׃m/�Wށ͑7�G���������C�s�ݤ�b4ȱhP�(+�YA�f$GK�ee(�(�!AȖ��I��ҙ��Fn�Z�&��l�Ă.ʄ������(RN�,DXJ2!����٬�jl6;
���~�K��/v�PS]�@0�*+p��׿"EW��;�[�r	����㥗_���A�/\���L���؞��CXN$r�9A
���b̕�h�o+O�PWs��c�\F�_lA�VT^���>��7$2�`���8{l�\}.��#8�v˖-#�6�EW�Ȋ�gh��_}~�����-������D�&`��')2b2h%���H[��Ա3�c�"�.�)-����/������Ur�w�g��r�X�r���?^>vR:�֍U�k��誐��H�������3��L�7���wv�UP�a}��*�#/����<����r
%�+�s�Ba��ȅZߴ��ʐ/�.�qJE���;�E		���m��N�d�㍷�b����S'�E��[�e��ѐ��3������&�0�lg"�G�΢�4Fb�F���^���%������+��U^^.����+� .b�<dE����I�y1W��X�T�����3�ԗn�ӦE��
aX����*��O�=^m7>8r��k���%����HZBFղ�i^���`�m������ʂ8T�����H9x+��O��\���`�F�18�O�t3���PWW�k>q,��*�z���?�	�]28Lxm���z㞩��>������q@�����P^�΃j�Z4�d2� � �3�|�bQs�sk ��@���f2��H�S��=������]o�Bxfm��1>�G��h�Ǯ�M���zq'c���ci_�YQ�@
��3�|���%pY
E�GEe�R�\>*W� 2���[��K�dr��?� �8(�e���e6sQv�7al*��a�ۦirRH�g�S��ȣ��k��V�,�1��.�)��t�'��?���@Ii"� F�F�S#�k\*P���N$)2^XdB��D��J��a.dH��bk&��VH0�����bQC��3m��!�E��z�-ho;��k�㲍��܋;����;�Խ[�%\��3�3Jmm�ܲ�k[6�d['�+��CeE
��������w۶aÆ��k.�� �(�f��	YIKHr֖��CZ����D9?�Z�X�b%+yx�Oo L�[e:���i����(v�Swf�o�=������y�Oy���)"���)1serУ�d!��~��,4�=�I-_��!JG��
V����33WI�N�>���Ĵ�Zv�lNli�\����)�B?	�c0(f���O��S��}��o{V��ޢ�B�����d���	'n���y�
Jʱj�:T���	fDI9��}��"e�Yܹ�h9�Y%��ҙ\բ�s��֬���d0jۼ��S�e��wq)Y�g*�Ν{0�ۍ)�!.�Ѡ�|�G�f�^�-�9d#�����k��/߃w�݋��D�%K��� k��ġ��tٕpXͨ�����ag�"�V��WA��G�q6�W!�b��&@�&�F1��t��1���_(�1�_�	=�ڰn�������J�����n�z��
a���A��H8�<b�<�Ņ��񡴢c.?ފw��K3�N�Z�Q�
kQ�(Z���ɞ$KR�l\N�V��'` ��V6����E��'֭���W��m�8|�0.^�H4%5-�(���[tU���D]m�z������-JK���L�<**`t܃���	�W���7�Z���E�n,$��[�V��0k�����:�k?�eK������l�&��jCS�%8q�V�\�}b;��|�\��uu��&�~c'YU
�z���a������v�0�]�L�s��Y�AV�N+)$#�δϋ��Jb��f��7����,����sx)
��h!E�g�A�Zڻ&����C�4�GØ�	axz/)/��=^
���o�lv���[�߂��b"�c���y�Ld滍���c#����#��&���ܰ�@?��������q�\���2�Z��|f�O�1&�����s\^�(��u"��&�s�k�RS��U�c&r���)�2�hi`Hcc��qa���;�^��-��7>��n��V;|��z/���g����ن��
��Rϴ��4EY\�`�dGlu;i���'���h�[�� *f�H!��ϩEc�4K<�Q*}����"�"������ٳV�O��=� J˪���&�Z�ZJ�/�*N�-�.Ϟ>yJ}����A���^y�T�]�إems���s�k��$�!用j�(#��l�|-��w�X���G�SbFQQ!��+�p���*���{�"II��_ǒk�5k[$N��-�FY4C}�I5�mWW�]�ށ�
�
��bT��D,��K� ��v�koΕ_��(f���S�YY�b�<��DB����B�6��R���,�z{PXP�(�F��S,(t������ÁCm��ýRC�E��L�044����R��NDbi��_`Ś58t`���ZP]E��b�X��kڪ,Jzĺ����dr]��Ė�"N�g��O'㈑��-f�"ڟ�U�f �SK�,'h*�����Q\�������j�ͪ��?I����ޢ�B$��5����!����'��,1��' ��;08<B0f��bCm������H��K��}V�u؊�Cz��3�3����ӗ��X(z+*v�h�t�pf����y_	�F�s��3��[n��	z��Q��Ƞ+��e_}����HS��Eό���EQVY�<��(W>��]my��/�n���oa��{�0��V���������JI�.��e"�I�D �px��]"�M>\��!�`d,������n����Y���Xo�ׇ�����%�y�m��g)��:߃�j�=y���(*-C��U(��k�1Q��lq#��v��FSm%�6+<�#G��514�DB�j�����p�c��$.�Pa&�&���k�Dج�ϊ��M���-8s�����z�V����WwHK7@o�U!	��C�j]ݥ��ի�|�|��?��] ��ru����}9�������$X�U�2�]���uxg�[I��>.�&��B�]�E���"��;;��\*��8Q�#�J��{_4�VV�c�@��+ω��>�'y�D��Z�z���;���?&��X������c1�N��o�q����!�>Wp��]m����)Z
��)ֲ��^�#ַ�D˺��U���������"��z� ����0��/�����Z{ǹ3���I��O ��k�����Š��ˢA�s;T�ק�Rh0Y��!�Ոĺ-���х��6[P�e�U��>L�"0���wZ�5�/H$�p:�[n�
�k��sQD|WLT�4-Y��L�ߎ"�I�}|��MAN4�$kQ4�O��r&���4�.�ҫ��Oi��P��.��#��څ�pd�^��3�$*�ax�BX��P�'��������[a2�p��Y<���zյ�tU�oe�@������@Y���f�H,Kpv�ͷ�p���^E�4������Cx�w�<�o�������bH�X�Tc:�2� ��T#�M���H�&� ���եy�&�vY�=A�`�y�sW��*��A���VBza� �B1���N���>+������v��P�oބ��a�,�艏GBŹ�!�Ҭ���uR͂j�-�󐆦z��|?����D9g:#���v F�"2�ĬO=�ȴ��Z��
�za9�f�h0;�sG7���㉨h -/�j�Y�;r�(�sb����N65aղE�A7[�q��8t���z<���ff�������+���6���S�[��!4��ĺC~���� d&"lFQ&�
��<��O�D~!3>���I��\�����a$�x��a�{?fg���I�Ϋ����E,_�\� ݟ�MRt������qW.@�+���&��'�A����^�b�1<�GOO��Z����c�`� .�R��0Y���_�F�]T���TޤQZ�B��������1���P�[\R��#G��n[6,V�ݙ��l��;�"*M81�ʦ�Ŵ="*��� �܎�*%\��z�ƆQSjŵ�n�ٶ���G��y%���Գ�/�W=Sb0���"�`s�5�F3���҅�p:���m���L���0F~�<>��%豹�f�Mљ�"�]XB>AFO�y�aŖcu�(���T�W�(���E
��֣d!�Q�^��J�5��b��-�l���4?{��-��_?%��7�X��pth�c�)�M�"p��c�����@�߇rʳS>
��t?��7���&����gd��,V�l��K%�()-���^'gE���� m�^�*��+]������e��eJ,�.���@e$����y���0C��׏k?~#���S�MzE%�������Ս�q�XPP�鄑�f��K�!��2�nb�I��s�.�u ��@
�6�ESi-m�����{���ʐ �rin��M8z���ct�z��
i^^��������>�F�����_R"v��%Y�ق��2�T�#��)DFg�{av�!����C��s�<�r���eee��skCw� 9�$��JK�yJ��s����ˤ133�[n��:!G�PRԀ�U���;X��	z��]�&�˖�O���_|�E��`�lU3IX�_��S�Lx��xQ1ƆzE����a�K��;�q�>�İe1�M�m6}g%��b��ň���o=��e=Y�⥍��酛,����#��ލ��?+�j�����?�=�R~^��AoѹrQ!Rl|c��{?��H&��c������D-)J>C���clM��v&�2 �@L4��j`�;Ol
�~��������|�X�5MX��������z	�����)��B$'&F���<���&g��WRb�FgїJY�!��|�|�g��$s��u8`!��H���
ь]C��]�Qb�ee��s �>��x���O�[��d%f����Lb�#���s�OV[VE))����E��L$���gPV݈�`������؀����<��-, ��[tUW�3����H�ml!��©��(,-�e���Y�;.���b�S��������0=�\O7�t	�8r_!�"	��,�g�߲9�(�iD$���(��
x�Xl�������v9ɏL!U�%(�d6�IE�@wѽغ�� =�ko�����j�K����ZAs��5S'�AeY���2a��9�Q��*�ML�.*���h�<�@P�%h& 2��He�h^��+���&DW���kP^Q���ދ��>�uww��+)�s�>C���d�׈�
	�m��d%G[O�Z�G䣵�����}H8��b�N�1Idp��UB�e�(�Y��q���!���p5J�L������0���4�r8�P��$��-,)�bAV�"�9fHF�_��������]�qn ��PLV��#�Ȑ�*x���q͍�»o����d2�����ɒ���R4-]�������F����t���L��]z��Ѱx	�.AQq9�ɲ��Ӕ��a��{��q�q�팀Ы�������C~'���'����z��
��#�H'�R�D�Z��f���Ǥ�z��:-c��C�ɡ��;�׃��j,ij@w�X�����ɓ��n]�8^��2�mk,<8;����s�g��Cl��w܁��^d���j��ڍ$L��op#���^�()5iR/��$��J
2�:ڲ�k۳"�$���ϋRN�x�GS�	L�n�C>�OlL3C���!��7R ��1FS�)���TTV�v���X��NؒLf+)�����E�����w���Ь����5������}��ܡ(4��,�儢IѺ�=$-*��`ݪe�����A1Y�a�2�M����4pє�ID�4D��EY���xR�_�w����.]��6]*��"���3�� ��Q
m�zZ,!��7�u��0>r�����3=�u
�E�M0���<���b�k_���b|��G÷�wvR$4 ���z��h�G��K/!�RaLGQ� X#�w��-8��&��1T���p����=�Fi�캵�4�!G=�yY���]m]-��b3BD����P�h9��]&�u�V�����#r}C��ۢ�-F5��}���;&Db�"*�ɽ��MX�t�	��B�o܄�1�)4�?�w���n�/��&�m{_��]h;�&�	��ƆKp��	�����wcjj�y����i
����!@��C�O��8|�R��3?8<�]���]grZ��^��!�T�[����Y<A>��_��|�۳KXΕWl�G?�]���V�o��;^����0���Ά�~�J��a?��������:o*S��]�TU� ����12�CP(��a�pۭ8r�0�,������}x���E3����~�,E`�R}�%2G�-:W�H�g	�����b6�U�MK	�:��F轃|	��(Y��#	���_w�Up�c��}�!���$[T���Ξŕ�ՕU0Hx㭷p�L;zz�(���n��F 3q��,|o}��y(�"e����;����h=u^r��[���x��!�غ�����Y�u�})���I"t!:�L(-viU$̘���:D�j��f���p�R�	�<���OR�v

�=��S�3�"!is$`(7
�i�F�,2YZ�*��r㺏~�v�Oљ	z��Q�B�Vái�����$9v7ʫK�.r����]��6�.��Z-.�`尲�n'zη�F���sD?1��{<��r�=�Jlq�	��&e~�W,P��Ef
��k�k����J�t�"/��MJ]n�L�_������)%�9u��S\�XT����G��GB�bwn7 9�˖���b�f9祤�vV�UN۝�s#����D"���U���ʒrr���W~�h���G���	�lR0� z�8��"���V�F.������a7����b�~8x\_(zC��4���2Q�;a£�
&�_���]	z:�	�|(+)��\x���LL���XpMϣ{`L�{=z���Z��?�5�r��U+��
��e��7�wI�=��\T�ޢoE2�]���6��?}�0Z\��u�31���^:z_����=���w���#2�q
m�;���e���x�����s�k��+�����W^���E����������5�c�uå����P��gX��l�`��&�,�X�b��>�4[/r��6,h��?8|~���~#���$a���e��L�11�%˘��$���J#�D�^y7l�^�i���IB�[�9O�	[l@<���ᳳ�t"������Y=êb0������	�ӥ��,������Yu{fz6�N����Ɔ��[tU�wr�f���"o��?5Ks���:�u;R^A!F'<���1��J5�,��BcZ�����i������_���l��;� r[s{h���/�����nj�l��_�}���P�%��$�ɧ^��u��3j�T�ɬ:x K֛M�����یw�~Gl%��誐{�r���o��{�L�r����h){�d3�Q���C�wj: Be��j���פ���X_/� x�xl��\PQ��}꼟/��V�%��Ǿ;�܋/Sx�x5*Ii�����l�5�b�zIDEwomen���oJ��Cc��W�"}rח�(����޽S'����~��_�O>�\w�w�TY�M&N�KiY��V�*?�S<�-�t������{�݊�Kq�UW�?���]v��#����IJ�u+)C���Z��#�dI�?knc3��ͳ���9��]��(�+���/���.�B�|��y&*d�ɇ
�g�B�|��y&�(��5�N�    IEND�B`�PK
     #{dZ�+s`(  `(  /   images/8a1d81a5-79d4-450c-9f72-108cd2673013.png�PNG

   IHDR  !     h@~   	pHYs  �  ��+  (IDATx��	�U��Ow�Iw��C��" ��!�@AP��EDAYUa�W�A	� 
*02��8,�2�b�ٓ������K���;I�[����w���[U�T��޳�gp2Ƙ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!�[:	�9%��f����Bw2f1X��D�KhI=¡�5�~ww�{�<˵X�D�lii� %$B[��tϙ7o�d���/�����̙�ؐ!C�5k�S��H�A��y�X,B&X�0���c;�d��3g���������D^�����
�::���,����={��6��k6?�zD���s�PX�.���"���ں+°�ܹs[�O�^��6	GmY;����_/B��-��Q9rd�4i�6�<x�xhw���5�7?�B���3��Eh�1
a�18���DxS\J3f̨	�СC"��V۶0a�gAR�+,��5j�:��!>�6����u���X�7��6����/%�',B�V'�������,��Gb!���LS�N��!��tꑀ��z�Ҷ#F�)S��DM����-[Z���ؿ˯p?�r�����٩���z�&�"ԼDe��q���F V����]lK]]]	a�	����Ӵi�j��ՋA��7�,d˙�l�rk��`��r�~#���B��V[��E?]���m4x�r�x���g/'ӴX���yd�� _&��$a���Y?�_� �zX(ai��^b�#���r�?�J�D��v�ʛ��l�H�FV'�Cp6`�!�!�ۢ� �G��=�$�Q�v�h��Gr�'8�Y�������d�
�P���քo��7���($KD�_V�,�h� Hx�6�c�������}q�����n����
�>oMX����y�b��,����v���5_���D�L�@�u�~�LSaj.��3������F\E-Y>Qg#q"c��v�ob�
��ۙ����g�A��`��չ��ҖQa�b�,$ݧ�[������[Ա��d��P����q�QS�,	�ňe�ԩ�c�Of��C�I=���\�ųΥ,/EX6ClGh��:�N*��a�I�!F[�<0߻�8������~0�B2�0e`խH�dU�U@kI��s5��������+ �����ܯ��B;A�F��$Ha�q�Z����7�[�*�E��a�Ex�Qf���bPFU�2o]?�Y���		R��L���������������F�I�<����kl߀�O��b�Q�RS�5dȏ����Z��o����l;��?M/v5:�p��<�8\�%�����Bd���*���D��"T=$@ji�H�d��D�Y
�(�P�KA���z�y�>��X=_$^'+���B�57���q�$|��d*�E�Z��Y�L�c�[�g��㓋`���@�ݖ�_LQ-���x~N�E�զO�����ܲ�����d!��꠺�6��7�I[V@X@Q-Ȉ�a�?�<���]\7�*���=Ԫ�g����zs+AM���`�R��m��8��y���8�c)5]%m��x�x�D��@pц !�hʔ)�O��R5���P5@{ڮ@d>���h~��^�Df�q:2��o%�U�)�9�&�ZqTB��	Y�6g��Nթ��X��}^�@1���5,��yd8����V�~�19?:'wb�?�M�Ѱ�T$;�pR�54��gW�����/��1ad�����Y{-X�_c����y�Ơ�h��,5PV�"��N�a�56����_I1�U���dI��M�v5Ǩ6�(�8�1u�T�����DVbt�l���H=^ Lbj\T��M�b0������Xj�?4%{ ��Ն�_��S:�*"�F�^�Q�}����"Ը�ճW�(g`�������T� ݈�!����/�H�eɳcWW�ֈЉwZ2�E�1�C�S����8j��.��ԣN��'b�?j��-����'"N�&�PX���g`�M�1#;����{�Y������Q�����j�G�wc��������c���\q䖟��Ν{Q2����I��)�n�kh����d�Pc��/g��	��1F
4��Fûru1tvv3u��I�U�.W��ܳ��OR��~� X��	C�}��Ř(UDg�����K ��9N�r�*�Mc�4e�{����d�P��J9��uKtHԗ;�#�J���d�K�Ո�]]]۩nMC[T���ɢ���3}�)�E�qؖL�M�W";&��H��az�`,Ig�.|UG�s�r�?����"T��x8ń���T��4�L�>�[�����G,�1c�v�(��@k�"}'��1ޮ���Gf�aÆ}PM���K�ئfe7)��s���(�$D1��ڑ}�&ww(�E� ��M����ch_jUDO\Ɨ���7Ѭ�5k}�-�CX���X&�W][�q �-B��������DgԨQi�����G��Ͼe혫VT!�W�Ƞ��y�k��ה��R���ٳ� -7�n#G�L�[��m�0´d�a*V�Fd�%BjJ������.�Kh�G�{h��8�?�)7�<e�w����灲��5k�f渄 QjIկ7�1q=�x�Q\%@*���ٮ��?N��� @�"<-1џ*�s�|E�a\B���Ɯ��ٹ���Q+\�Ov=��y=�p��r�P�D�ArN�./���Dl�V߫�{v��[���z�BX��2�1:$�w�<�����{9��E'�b�Hۢ�R�9��l:��#F���)��^���1U��ފo]ˣ�oE���}����	V�>}�{�eV�PqL"@&ш��\�؂����$4 -��(SemL��1k���x�Kszi2�[Ru�;�A|_E�WԊ�6p}7q^��'S�PA���/��y�C4~�4�V�?�z��ItBlDv�U�
b���B:w�eT�u��F~/FW��UZ+���;�Ϊ��;�6a�E��rhx��$Q�.U�"w!��q��F`vG�&��ڢ_L����%!��?�Aמ�5�I1p3�dg�,�qQDT�����s���T-jiH��&�B�֪�o�䎋%���q�X�Det��`�h�cY��A<6ͭjr _+�I@$$��r�ȟs�)�/�`V�����7GK|�2���-��R���kܙ�C-r��.,¹�{M�g:�Y�eլ��А��J��*6��,�9+�/Ǔ,�zL�fg(��j�A1,,�9��b_*�Ǒ���*~�05+{���|�c�FL��/�s�;�Ly��:��H�Y���s�>Ǿ/UkT�޷?#�S��F��{ǵY�!���=��|�v����#G��ݛ�󼷫�K��%n�����?/����A��2�02�~�	r����?��Լ�%ֈ)jԃ7�|�}}�����j�#���ٲ ����r�;���:J�q�a�-Bv�3^EF��PT��6���,�M�^�>��=OxN���ke�,Q�ZjnE���{��D��b�7Dh%�ݑJ���|��o��E����B&?�����5�����9�|����Y�D�DX���C�o��by�峤Ooz��U^N�w�D_������v�Z�-���^䏼���V'?	��M���i#�Ѽ_����l�MF{�x��1 ��Ѓ�	!�j��g���ɓ?�hy%��3f��o��ƥ��޼�r�;���?EH#��䡫�fe֕C,�j��"}a?G�h����&��X5�]�$D��ɟR�*H%@[s���v	��~�/"�W����Go����?YF�u�Q��-h��uCUr��(��@��d����oGt�{�7-�~�s���]�'�\S&M��z��q�m<���x}d�ŋg������ROeh|�D��e����ya~Hg]e��v��Cc#f�b��;6�ڎ!C��z�d-z~��4eg]5+((W6N�=ߗ�{�{��>Z�t���X.1.d]����* �Y+r)��#�[��
����:«� �}�������q;S���:�E�엻�����r(�M%@���*r���n^��Y�E��D�hި!��������,�����k�8j����d1z�ךC&:�߭�:%���T����	]���n2�����<:�/QY�K>�k^L�O�V�gb�������L�1bĚS�L	�S��}�V�eq=x�k�L�7�c��-�H���>�ǻ�!��i9�/"Dd!�h��p���������1��d�.���"���Xw�@ϴ��c�m�7�߆4���2���1^,;ڊJ�ތ��GD@��k���F�<���J�.��y�%�7R�սK�����p���f���O��Rz)�n���2aK>Ӓ-̆k֮'|Oq��������Z���X�H,qQ��?�����~�զ�d;�/�ٻ����v^u�_?z��`˘w��� ���"�$�5'm�S;k��q%-"�1#�2�"b���l'H��;����u����G ;�W<Ԫ�
�'��!��k��JS��R�3#�E���>�������Q�]u�E���^�h����x��#�ҮW�x�@;>��"BS�NUѣ�#�_W �W�	��	/��K�Ҿ$K����<wX���z�&}��'�[�`_�+�8��^�ճ%%��Z�ukZ���E2�7�����<-�h��"�eBZ>ŲZ��;�[B�YB����n ��0ߧwl�gE巼�y��f[���8[��,DUi�s��*qS��u��?�:3���}�?Dh�1X���!^�ړ��5\���4�Ǘ*��zѵ��cR����z�<^��X��o��|*�uq�S��9�4ە�Nშ�(��*���&h\�ѭA³e�v�}�"��}�^���R�2o<��f�8khq��Ҿ��#�#��Ļq�7���u_.��>.�A��	�`'�r��ǟ�@Y}�^�0�뚞+�'�k�(Z�k��I����,�7k&	�Ϧ�G+/�2����)�*nZ�/������Ӳ&�s�G�OV�`\hs���|�rboNE�z�n1<%����E�gI�l˓z�	��V|���u���VeJ�����"��E݅�9'���1l�;�r��t�"v�آ@B������é�K�9[Xf��Nc��Bs-5��.e������Ձ1��?��?�B��1©<���d���ٜ��o�Ӳ��T��k�b�k��ݽ�8 ����L_��F�j��Q�]���UK��?fi-%Y;�܋���yd:�ng��9�����3~�;ᷩ�ⅼ���S�׾�Ғ!۰�N���DU%�::v�s�1�i��{�����|� �ePŪz8�݌�!���ZgRjxw����=�Qct���E��ԛ��ep��Ѥ��
��B\�Y����߅�5�������$T���(m	���ʴ��4{�x�D|�����K|�<�q�&Mz?˝S?�"�y����}/�fi�lp*�|�/�|0�zZ�*=`F��������԰jj|¼?�L��V��u	�����l�@�ETk�D؞pvi�5Q�v��pd�n��u���s�u�"�'��,� 58�<��xG��k�	[�G���}��}��T藊i�����r���m�E�o/��$�ЇROSs��%�f��^���r9~��K��+��E~VSW�<����� �͎�.�yF���P�ի�ZDmP}}Y]�p������^���G���E�^X\ѫb�M'�|����^yh��h��א[�A�'�C�$}�"܍9��sH�q۱ ����/��z���y�2�3���x�[�F�+S�#�=�=����ٌgv���Q�T��C�I|n�Y3O��[7�"�.V�<*j�7'��--�~ȾK{{Üs�h��� �ٝ���9�ۍ��S��#<#8^�po�3��25�m��ѣ@���a/��XO�%����2/�*9��f/��l7��e[_=7S����<��z�wD�U&�Eyi�ު̅���q<�M�-�4��h��<'��I��j̠��M��F������2���ėZs��K�U^4x:E�^�T@��U��<��ݺJ�����<�ߓ�����<�����r�����N��s k��Q>���D_��W��H��HYH`��V�R� �q�����d�,oO=3dT�a�T^��4�g8.O_=�*b�Z<�;ؿO�i����n)�k��H�5c��h:�� �b�!����>���G�Rt�Рa�Ϥ��ɓ'��Lb�;�d�p-�����l�թwr�Z��BIϊ2���a���@_���"���?�r�$OU!Yx(��dP�Ft�$�����l;�m*F�ú�����qٳ����<C����z���vWnQ]��=�-bu��3u���<���XYH��w/%E��-��P����?,�U�%���B�׫8+��}+�����,��ʗ���iӦ�N����gf�`K��C)����$�����d��5�N��*����X~�l��*�ݗ�%�{�tG��0e�\T�6�J��~/%.È��e�De�P������ů�]7�`~Ká^"�e�}����"��!;���K��ӈ�|���wS`*��x��<�M!3��*��Y6$��S�X�,�B\�c)�l�����i�e�Hl$@��$f�H��_i����s�^��ա�~�q�e��0u!h�y��"T}u�%�=�1Pa(s�lO=��(B!���U-q�
�Y;�aŠQ��n��8� q��R=Ӳ�3�-E��1��
{��'P1,B��>�7״<��Y_�<�^-I���b�b�݄��iX; *m�.b�t�~i[�\+�!���y�|K��t�%/�W��<Ѥz)V���X�
�%t+Bt�(|��H�m������oM�QS��X"8G�f{X��i�,"�`�����&�QO�e%
c�$&�����/�ŧ(�� @�!���z�r4���n�?+Ue����d9���>"�. �e��H�%��:e9\O�u�DHT7����,��X��#_�j�_/\���!�h߮��f�z42��8pd."-���A��H�?U��Ρ�!��6��Y8���;d��S���}o2ʍ�9��㾥a{��m��Q�=iN��3g~'�(V�Pc�G2ƭd�D/���V�ݚ��G����45�
�9^VP�K	H_�+��X����J3�����]���ނ��ԙ�Lo�noo�V��c�}x���L�!�5d�[X��g�p�/1�n,Nd]�FUl�/�~bt�5T'@�o�"n�5z*n}��n���gmc�i"�K�YR��x���b������YLJ��X��p�5����XnT7��֛k��iӦ��s�D�/���L��w������W�c-@�E���_e���_�u"�c�l��Of��tZ'�˝_�&t�����P�1��	�f7���<��c����dފ	��g�ϕ�HUL����t]2�E�!��b�����{�p�J��mpY�����TRm�c%@yN7�prB�����"Ԙ<"^d�3�e'f�D�FR��1�!�az�&��r5�:j���DP�Wt��L�ajL��4g#DXn��y����˭L%7n�O���gΚ5k��-�$�y����/%ӐX��yy�_�U�/{]?��'(n����4�Qk�&a<6�p;�AnaT�K��2{ɀ�"��<L�:���ZQqL�,�ȓَ����o��[�q�<	N�

?ҹ2Z�k�N�a�5>� >�"S� �J������.E��хi�(�œ49�������ȑ#kn:�`�k	_M���U ���X>����}����t%#v�!����¨�r֌���Ū�QŽ�b�|$@�q���b�ip,B�@E������׿6Gx�N-@Йr����Ss#+����h�*���2�il����
`����Fc/D�V��T�Or�2�QXkS4�G�f��՜A�]k�'>Se	�_�\���]���T�P5�1N��}'D�7�ѣ:�)ڍ�G��p샩9�f�^q���F14f����veߓ�T�P��O���p`yb�~��!�E�5X�!:�㾑�],�x�r6q���
�8��:��IDiO���jϤZ!,B�"2�F�O@�n�SF�|ﵺA�B�<��F�c��RuP�Rf�:�ͥ��6�	(��zd��\m���QP�Lb������OF�.���ڠ�E��\P�����%_��\v����b�A�N!�=S��Hb>�$@���m/��&SI,B�f��4K�U0jԨ���z����H�/������������mν~���gm���F]P�B��'�ǧ��T�P��H�SRO��K&O��NeV՗D3�2���iWD�N�$�d�k)�\�o/p��%@����P���b�W�zP�|jf��믬j"ś��<��V��%[.#���欛bYV�*,O �ű�s����ăC����	`,�!,�?y@?@�c[B�gKU\n��Ϥ��B�gm,B�'2��5��BT�c�����5eEV�Jd�<�D;a�hD�E2����V2�*��J�8�wtt��z�r�}��hm�!(�֛�%B�#�{�ߝ�%wI�}Y�� �P����z�ȼ��<�.k(��š��>U�a�{���O��i�osx����߫���\��� �V�Z���r�w��!���T��:_`��=*����=i]��u�".��J2M�E��1Rߠ�W��O'c��b��%��%@Q�-d�H ���,�U�sS��F�ʶ	�Xc���]0��9:��ƾU�M��""2Z�sJ�t.U��ꧢ�=H�=Iu<�����S������,�P�3xȢ�GM�h�g�<�kc�,��wɳ�F���P�h��fyu�<#������N�&tL�S�]��G�#	��1q��-�v\\����mrO�A��&�"40P����,Ւ�/��d��"�KLd�h]bT�,�y��J�N�rS��b�����#�c��%�Q�\�i�7�5�=�\�3`�,���&�If���m���RvB(�i0���N��:����]�_�"��џ'�$XQ��!b�/��W�흈�D���Smz2���E��?A~��������KDB�oC jC�%
!R��H˘RG��(���߅���uq�GRO��_�#L��f`b2Bn?~�@�<��LXkg,�w�]eWTgG�dt4��$b0�Q�fO�<Y��+��ˈ���{�}������.6Z��X���А���;c,�!8�XvR��4�#YoǺ���B�fp�,H��S�)X8�T^Tݎ�}�E�,�p�!5z5-0PT�/Q'V��
��Yv�a�+!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ�o/�9��l�    IEND�B`�PK
     #{dZ��/��  �  /   images/aacc0029-e57d-4614-a443-d9bee65b5175.png�PNG

   IHDR   d   `   �s�B   	pHYs  �  ��+  2IDATx���VU��~�� ;�Nk�}�N&hEa�i�1�)h6�#9���$��A����:�4JEѨ58c�|(��|-���l���yv�;��/��Cs�3�<�������s�sιoq�
�g��8C$�"!�	q�H�3DB�!��g��8C$�"!�	q�H�3DB�!��g��8C$�"!�	q�H�3DB�!��g8��ӧOR__�'---Ikkk���� ��/**zOysssr6�=!rj�~���Ǐ'���I����>����(D�s��}ًlA6A�nd�(-"=�-!���m�t�A�?e����}�����sU'g�:�TY-ׯ#[�^I�:|�ԩ)�Wb\RRR�455eH��%8��3��PΦ���+�&���Zҧ�s�F�c�3
=���ݏ~�B{���D�7�#D72�(~��c����F-�٫�8����7�n�!�*�7q�'H?��S�w444�KdX��w��A���_%���i7��觑#ANM;�&u�l�n;E�I/�}�{t�����Vz�3�^�x�;B��{�Z��p�
��"�G�y�3'�� G������$�嫹�QҚ�����/���!D��0�_���Ƞx������۷/�\����L�"��)�V�����;��@s���E<�0u+D�"8pA�E>8���b��8�1����ݛ�32r�z��>v예�B�7UO�-�6/�I�	1G�a������z$DU��=����?�⫑��]�s��F�[Y㔉8�#��$�bsFOA�4|���N��ȗ����~�rM��D^	�ի�mm�!"�!��zEEEbÕ�ȳ^�K��������O)��A�G��wԕWB̙8f�����/�#�V�!��	��q�ku��wg��dH]���)�"�9�Vg���䕐�#'�,�ְ��z��"�v�nCC�?R5٥{mu�@DJa�t�k��|�I�$$,��V��9RN��2W��R=6�}�~�F��5	ɉ!_�u�P�U�?�_G�+�%#U=�h}R������'J�{f�'N��zVB�6�����9L�z�g���}�s/�]H��2��lޡ�)�?�tϜ���k�q�C�gI��p�u;��O� �	�Q�%�ڙ�S��Z��{�o�7����,k�����'ON�n��`��FZ녆�R]6�=lB��8�/�7(>`=1s��N��Wx�ˡn?�h�s�ǒ^�5�I7v��H�n��γߡw�$]A� ��NsG�eCx��m���vmvG���_Y		��J��а�Q���~[���v״�k��ѡ� �7A����B�{�#2l�뉣��I�Z.�=��9��=)�q�����~Dccu(���Z���t���J;�B�o�g�ڌ��MB>Nن$��!�|�lS"�����+)��5��{��B���%l���9i~U�^�°����܅V�:��5���}�ey�g�˹�a�;��!�詶P=�w���VB��4���
�)ߢ!���		����љ�=0���gl/�QK[S��}y���
io�dǩ�kx�����9eʔk�-[��H�&}^|D�[����r���2k�TP�i.�1��{5���!���1�#ȿ@�v��l.
m隉�m�_-�C�!�V��i�P-z������?1�-4��W�W��/j!�L� ��`g�2�ql�K˗/�f¸��zY�4K�����N��6�!�H/��0`UMMM�,��ty �'����No�����c��
F��!�m��!aVc�y�+0|-eu�&��g��~�Ո��՝u��!�t������i����n�vtq�&��8|�NET3jkk��0 �)cN����QZ�,��?zmYJ;N���!���߮�m���{U{x�[d�cW�Kݱ��0�%UUU�I�H����㰫3}��D��,�l�1| 1���Bh�vz�+d��HjnKl���v�T�ra��<�	����Ӈ��/㐗4u���D|=/yw(T({Q���L�;80QO�n|0���鉕�>��y�:	a�J�u3ΚH~.����PYY��رc=��/`od8����y�@��#G�藫���0�<���1"ټys�/�[��%�)At��H[��)۷o��
}Uer�m�{!}��I�oЎ?��|�!�;�C4l��,$}/i�Z��a�9��q�-��y����{T���y?�JB-�)Sѣ�yJ�<�]�ΐ>?Q��SC��yR��7�Bи�]��HК���{�P�5b���Z�� }�'�ƞ@�	,6��/�moh��z#��-����VGo���U�]�����R�؞�攲��ǉ���-b����c�l~�m�l��?���/Y��	�|�h�.�q�x�8P����xq���e�Y��ZQ�~����	�4�� �d�i�X����lV�s�(��"ذș��u61����ׇ���}mXP&�^c���Շk/�j*6�#����t�g�p�r���n e%�uhmNC&Q���v�.�-h��hX[��\�\�}��a�DkA���~Dz����IpG�`�
:�ӗ!8�	�x���%7�<a=�vSAo�\I�R�&�ۑt��V�$�`�a��'?�S/��bm��� }�\��Q�ꬆ�:�ۀ�[�7;���kB���R�\d�i�������a;�-H(//�,���N��	i96,�2V/R緦��E�ꪫ���	g!B�M�����?��F7W����?#��g��8C$�"!�	q�H�3DB�!��g��8C$�"!�	q�H�3DB�!��g��8C$�"!�	q�H�3DB�!��g��8C$�"!�	q���n*e��B    IEND�B`�PK
     #{dZ�1��� �� /   images/1d90a712-93d7-4555-ae10-1782f839eba3.png�PNG

   IHDR  T  p   ৆  0�iCCPICC Profile  x��||eE���Vx�*�g\�$�{�R�f�IvC�]�%�lv7��l��U����E�4��)"ME��   �4AiR��=sg��E?����d�y�3��)�s$���_�`Ψj�̝�h�{���{�U�J2:�T�͒/�,\���Ց�'�~��ǒz}���J��~֝1�p I�W,��K���- �~��g?G?K�0��g9z�J�'�7q<�ݭ�S�d`���>Iƭ�?�ha��������sA/=a`ͻ����;c�I�*$�̚�x��ch̹���A��$c�\�?<+I���g�\�FЭ�m�Ϥ�%�����2���L�Ve)cͩlf���:�����y��C�4MR2M��4�1�5�kʴ\����Ӕغxx�ඝ�{Y��"��t%,I��ݒ*��,iƫĿ,1h�HZ�Ix�:��&��;�%�6I�8S�ׄQ�u ���M��{���K�<@u�ǵ�1c�%m[��&���_��^[�/X:<4k��j4m��>o��Dғ�,�6�~{��ǆ/<�����,��qA��m�b��(I�x0I־<�m��d���䶶H<os
?>Y/�*����������\�\�ܖ<�<���|аJ���a׆}�5��pm�C��Z}T6jڨCF]6�ѕ�;���ţ�����1��yb�cg��b�?��qG�{`�F����J��x��V�b���X�UN���ʌU��j�w�ֲ�-��կZc�5�Zs�5���'k��k/[g�:����7�׽�+����p�m�y�6Zg��7�k�1�\���6���͏��~1��m��~�u�J~��[l��V�m}�6�}y�/���EM��w��W{�+I�ͮc����r��[O7]v�v]_����w�񀝎���-�M����I��y��[���>���w���η�n�պ���K{��6a��ݯ�c�^S�q�7���侳�~c��N���L6����۸�����l��O����[,9���.?x�e�|w�CN>l��O=r���>z�1W�k�=z�~'�;�SZO}��#N��ߞ5����\r^������{~��ŏ_z��G^���Z��p�'�=u�/n��/�~�˭�ܾ�����;���{ο��yp���,�����ɦ�����y~ʋ�_������ޘ��No�w�����?���-�D�X���3�0
�]�ɇ�׍�`�a��='���W�4n�q7���Ru��W��r�*Ǯz�j��~��׼`��׾}����z����kn��F;l��&�7=u��o~����K_�дE˖Ӷ����m����^�ts�ǿ�B�f�o+�5�zzc��m�n�f�o���;v����>���']�v�ΏM~i�w�>v�M:d�nS�N=������~�w�i[M�e��{�����7��+�Zѷ��[�o�ϔ��s�<`�wf3��}/���9��}h޳��\���*7^Դx�%��ׁCK�t��g,��;7}��C�=���W9�z�8j���8z�1��=��?8�ǟw��?���kO���מrթ�/������'��s�g�z�~t��G�sȹ�w�����'����-��܋g^���/���h��+߿꣟���r�:�nv�6��׷��q��7��r�慿Zv�Q��x�Y�_t�տ��o����w>����z��w���������?���{���{��?�������?v��?|��?��§�yzڟ۟��/��m�����?���^�����m�+����߫�h~m�ק�1��ҷN��eo���s�~���><��?��֏�[1Ɲ��ɿvo�a�&������/��5�ͱ���t�����J�\���%��������k���kݼ�=�<���������������	�]���'��֗�M�p��-w�j��{o��ˇn{rӏ�^��+���gϱW���ߪA�7��5�[���o��rǖ��|��-�'�z��]��o'?������Z��b�W��N]�u�n�u���Ҵ1ӷ�}�{�y�^˿q�7��?}�����o�O6�6c�`�̡Y�g9tھ�w����>5����ko��-j[����t�qK�9誃o[��w���|�f��#ڎ�����;�裎9��s��q��	w����>鹓�?�S_]��io�����=�3�?�}x��|p��}t��?^q�xQr�'?}��]�Ko����O���+�ꨟ��S�>����~q�����ȍO���/_���z��nk��r�:���7[�6�s�ߵ��{���u���ܿ�s~?�����8��=鏧>���S�8�O��?=����L�ˮ���\�����~a������}������m�^������.~��7.y󊷮���8�����{o�k�k}8���Ώg|BH�#�Q�Zä�s>����G�ї�i�_{Ӹ�ƽ=�ܕ����ʯV~�ʕ���ڙ�����k^�ֵk߶���>����_��FS6^���Mo����/nո˗fN8|�s��q���~y���]�i�扵ݿ�o�,;���/W�[�=�Q���v�n?f�uv�b'�������:鲶_����o����&����;�N���[���ݳE�iӏ���=~��s{����ߒߞ�7k�C�O�犁�g<8��̧g�0�͡O�[mΦs���8�kA����p����r������J^{ل���~���C�v��q������Ǭ{���Z��<a��8���'|ʲS����ӎ��Q�}�1gsֱ?:���9����;��������p���s�~�����K{��.?��<��~v�Ϗ���kN����~�ˮ����n����~y�����<s��r�w������ѿwW��U�Y��U�w������s����`����������cW?~�����'�}j������g��������=��#^�ދǿt������W��ο?������k���[;����}�9����]��߿�?~��_�譏��ɇ+���,/n�$����]�b�No'�Ӯ<��wW�x���a��R���k�L�R�H`�k��$[�̱j�Ks����#u�l�)y`��������%�Z�Љs���־w�N}'���ڤ��������8-I�w/3������u]�N�������x�ۿ?���x�̞l�����񊜡�!�*n�Ff�����+x�O@����D���W���������M��Fo�����/�����o��*_��'���c��㎡�m�W��#g �N��޷S��a�! �~ ���C�B��9x�-��|K�_��	�v7����x��k>�b�|�x٘.;�LaaB���}�A�U�����߭+Aֱ4�m�'�lP���T�jK�$�����o��ȍ�7"����T>ukjA>����AYƀ[ǀ�	��ݴ��P7�N7W/z� ���!�)U���a��&��u~����X�~��,w�����\Ɠ˰i�
�>w%Mu2hQ�IԞ�m2�N�Q���c���\��ȌdD��q���C�&���Az���>$d����fh�Z�'���t|
�RY�,��b��O�!�/��Mg�5��d�!e�l4�W�1���,��6n������>��m>�b��;��bNV䝽�Z�V*��zZ�ۻz�vW[�g-�3���?gh���EC��U{��g.���^T�7s������2��}r����]g-\0<�?��������6���ӿ��ٿ��L5��I��d�:Ј�������v���T'��tu���X�i�2���oR{g_Oo[�$1��ή���m{m�sZGo{c���jc��}�Í�ޖ��m�}�Szz��u�M�6���=�h�:�U'a�s��v�o��Ο3�s���B3V����wϮ6��sw[�.��)S?�-=m}��o�X����jk��n�ȻuL�Ԧ`�X\_�NVm����̘�jmMp�XZ�R[˔��4V�L��l�h߫mR_�Ծ=��4�6����X��>�mj_Ǵ޾V0L�n�m�:��kjOO�Ď6�T�؆�����胈����Lo{*�K���Ϯ6��T�[���ՁP��U[q��gTZ4;H�Ty��l�W��ͨ�'���Se����͝8�����6eR�ܕ�{ں��A2˳>�4HqbGK��B;�G��6����o����l��Z�X٥��7��x��}_�Wml���tN�ڻ������]�z�v�ֆc�6N��m�{_8a��5u
��}��V�L���݇�����1�����'�����L��[�i���pJA�������u5ɾ=ܿ{��rB�{�=m�=�L�sT2�v����Z&4�#�dk�Sa%�Z�״jT-���U5�Së�ո0�����|��OV���g�"X�E�1+MZQUvSߏՌPR`M5��Q�)SVWtU���/c5�,SUY��pK�	&S!*&J��%3�GGX8��S��ظ��~R�D&9��(-m�*��J��t,�,u�gBXj��GF+�⺒�И�?v4�yVe�k�a�c��d#T��Q�Qe5w��"�i�0��2��T^�b���Yn���2)-��M���(;��1���"���L1[5�$�}d��������יѴ���(Q�T�1�����*V(3E��A�d��8F�4V�Ɍ�c��:�d��wj܎>K@����u^� �h���F,˔��g	�	�&B2�II)�
���DZF����f������D�љ�)��ĖZwdҰ����X��L�-�z6)T�Å[�)�Q��pH���� �ɌT�&d��Y-���:S#�z��!�&�f��c��3���VO` �rͱZ�o�Z�yjmN!�0jR�z�՘4�\b��6�*�ak�����$U�,�*+p��aF�jR��	N��\#�q� �V*���he���5�2)�r#`��=PY����	I�]O��X�m	��b�ؗ�}a	Ο�贄PX2�P9U#�ġk�R�
[�X6�hN;�#�feʉ�ڹcq�O>�s��#��I����N>'��N*h��,�B=��$�!�Ԓ|)�Nji��n�c&ͬ'���(�p�b�Y��*�5o�uDF��Wd��֑��d4#����� mWp�ďȝ
Rc��0h������ؘ�QW3�0PZ���P�
���{������V0v�c���P�GW�4��)X6l�,��.�9X��
�!�
�9�[G����9~��;l�(HѺ�f�S-S�e�)!x p�
6.!j�T����(��?����g�(�����"��U���6U�TBR�
�#�g�k�C�GX�)q�>@9�(^{^G�PEi���p��A3�6��[=� �i�������a��hH��K"�:�+���疤
5�)Ed@%@�f�0�Ԃ��@�pĄ�2�+8#�j�FZF`|!Nj{���6�8Z���7VuA��BpO%N�W�)��J���F��* M(��JI��p\���mf��RZ�@�H�X�V+1�_G��Y/!��R2L�,ڈ
,E���u�$G��¬�z8;�pxX�2�����$M#,�(nY�$����q1����% �T��qdX���i�F(%�:��f@V
SK:@& {��ZJG�CiZB?&9��ٚD�68����#��B���Bt *��U-
K�YOh�m�f�U'U�ۑ�`�F�wrHaL�>��@dX*2-�aF
VO�&a���dH�Ҍt�֎��0Π��a�a�{p+`W�ϑX=��4�גpp��wX�EE���!&: u�"$\�%,��(]�5D�����ı S�c� ��)����W2�>��E$geK2��[��4�I��L�ɠD�ӒL��H~�4�L
���<p0L�_�+Dֈdڥ~��5���e{���*e����8t�đ�U4���u�b2M^�B9%��W-�=:��Q��:H�'���j*��b�����H�#+ ��'C2���U}GA����#�t�^
�uI���(B�(��(��g��z�-�'�X*2�|]8aC���
$\챾#�#<�Qsʩ0�Ó|3b��%eq UC�AHڎ�,EŔ�q�9��!�������{8VSVȉ'�����J���LX*/Q�(.8C�����<�BF�E�!GqQ���cF�f$�.Z芑%E��! ]�<���QM��|ᨒ�#� �t��
�����[�*d�xc=�g >H�E���H�tMZ,Ք�1�����Fy�&B�V1��Y��%�֨\J���nIu'�i=��u D�����Uj5:f%�@�`�P=red.��paι���� eU�:p���:��d��/�� `d��i�@x6+�XZA��?F$Y\80��2b��T���9e��UB�����P=^���c\*��8xPޒY!]� �V��Ǒ
��"�{��b��2:S��& �!�:�hH�(�� V�-q�EGAZ�H�sN
7I�V�Ҳ�S4��"'g�z
"�U�Ҭ�g\,"��J���L��|�
I�GV�Z?�MK�F�\�5�r���K|kT�T��|�����@��%�5�pF�.��\��\GU����\�l8;CU$��'\zH�=���EO���\Ru&���qFs�U���%�=����� ST=�j�EONY���*ydEU ��1Z�-�:~��6p�)%��r�YL�d���b��e������9a�Գ��{6v������M���'+�& 08���34�=y��D	Q��a�������K(=E��B\Flir���irƥ�lG֔�{"IǏ�'�Hwa��o�T%�&@oq��q��ʼ8_M��%3�ۃ�b��V�9��&S�l*+�AظO��lJ�3��L=��9mI��R�|"	@LU"CY)���be
0@CN�ƔH��
��²��b�p����"�p�1V�5�e*` -�s��6N�SF5錕=��� ߗRM2/��:`=\`��g$�p<B9-U�Ud�J��%^3�SQ��rߔjT��D�r�J�f�d�v-�Ne�ڒ1]�5�JPq�lؐl54����֔@ˢ'U2*i#OE?
��dX����k�U02.:OH�Q�N%�IoyiS�l��xIFu[x�n�>H\�����)*�k*�"�PO%��J�Iт�)�r5Fኍ�)�`ٜ�)z!*N�*�@aX)=yL鑘(�&QBS�Pw���fS������ğ��fya3��ss"��<y�����%'8Nk�uC@���� Jz�����?���\����l6��T�'�/����^II��i��lѓ�}�]	XC@N���e./����?9˔�G:Lm1���\A�	T>���y�U�'�,�����9HZB`,�r)I��5	5԰�
���5��ꎰ.W��*�ɍ��e)|�I��)0r I=%�������V�5�
�R9^I��=� uTCr��X0C���2Ms��}Cڢ��R�l�}�O�Ӕ���27�M����C��
[�oG����U�YQ�Ӑ��e�5�Q��<5ݏ �q�!���[f%�6��R�EO�$=p��D��IVҳ �
�vT� �ߑP)�[�K�m�	T�b�S�`gy����S�[��(�
hKF�`��=�Td��~����]ʧI����Jz��39��T_�G����2Y��>i�,/=��J�?�GOS�ocO*`[Jv32q����0�Q��I�  F�ψ9=n��JCB�4u,.Уz"C��j��V�a�L�F����B�\3�S�+�g�%��
�8��È��`�);��)^��O{��y�f��H�4^�%D�J;��pY��H�M�,�a ��E*3����jUYRU�kK�\:w��9���.U�����n``�0���m��}���7R 0x�D����C�C_�!e�BX�	˥{% R���(��2Oغ� �]�/��'�YHH�С��p?Tc��VL*���0����H?�!��j#�I�:�r?�8!������TN�tY�4ܕ�'�7-J�1�r{� �	��T==�AX��7�DQAf�f�,.�U�&��݁�4�dh`�SWa{�/�_����{����IlXn��ɪ��ϭ6/r�a��q{�6ς��6�̈��-��Y�y �K�U���dPt1D4�;`����DO�讑�HXmރ��5{�������?wh��>&��x|�������}F^���*K.I��K�t��������4�:dP����H���H�#T ��{�JIǫ�S~%y������ h�/��\+]��ܓ\�Z�R��x)���"���D��c�����U�hϵ*:u�I���"x#^�������i(�ʽ���v{c:��C�-F��Z�I�����YF����7C�ܓP>'(�6�KK��V���rNbk������(�V	hH�ؙ�� xG���'vҩ'3����>�@J�xuJ��]�ͰObe~9�N<W�M�|6hDrR�r#����f�5�(=i��$N �t�HQ�o���M^�j�#�*_��õc/�A��)����O.(���� H3?��t�x���4�<	8�G���+�$\���f�̌_�R���r�p�9�?BA�7�F�T9^�2g�)��'�Hs��HL���8A�� ��ۚ零,גe䋤��61��taF伂�3g�������ʜ��o�z��V�F�7+�n��.3s���K��]�|�J��Ѝ�8�;��q�/RYDG�QE/�u*�Z5L�g��t�Ϗ ���,7͜���'��Z�x����r�.+`�ĩ�n��Q� !�UH&o<��7'�4�U�+��kԊ���@�T��eF�����^+h5�!�;^���{�X�C��C��� 9�ίݑ���@�4��u��Y�9��+H/�&�nq�2�	�ȯu�d1��+9�M�l=7�)xh�T8��M���>a
E*���b����
�IhWn�E��j$S���o�.�K�+��X�R��
 ��"e4���ר���?�"��I8O��+DՉ�Aa��'�:�zI%d����ݞ�ys��[--���^ؓ�Y�\�D/H�DR������b?~0I�ϓ����C�k%���Q��y)�z^���!E�Γ�%�$t�xYD+oR�@f�P{�y�!?�%��t{*'c��%g�[�t ��n e�������O�I�dA�G�xe~A�Z�~0Lt�H�����ێpL���T��*��y��`B~9V�`�y|b���<�E�k/��כ�je.�y�Yo���qs��j��
I3�I���y������g��z}`)=%�y�������R��/a�[-��� )� S���]�k�>�_/�f�	@f��Y�0T�5�T��@�ԯA���,�K�t�5�<���;o��̸�6��Ht��r��Z�]�Ԇn�3^s(�Z�(Ȭhu�s^�_���w� Y���cO��10	�)�[�)�7r~0�% D ������A-��)��L=��0��n\x���@�5�)>µ$bk �6d��Y0�	r�y8R�\�<bFK�ޜ�U�[`F�@:�8�!����pR{�����GÌ���	�H�<o�a�h8X�d�4>��aA��y���*����!�����F6�*�y�0ٗ�cH���Z���a�n�$O�g1�����P�D�j����Ѓ��7���"��{$a����6b��-0���2�;fȨr����cz��@fao@�1M+��9�[�V+�z#��6��b����O���0ئ��	2�L�4�g���0�KY��GHNI��[�0o/�p��yxeP6La�#$���pł#��@	£�z1��}��ȴ��ĆxН�a8%�~�Ȕñ 'h?n�0nһ�i�:Sx�2��@r;�!R#�a8��c */I�a=o�a����Mʤ�k�ƹ����0�),�f���խ�Kg޽�.����<��X�v�#� o&<o�a�~�
��o=)�q#���r  ����E�"<�'2����rވa�kK�Dz?)�=��@Hʻ
J�6-��T�⁴<�J�x,"�p�Ap
>fa�J�q#�4Ͳ�aCʺ=�ټ|#�����D��*#�F{���2�w
 U87Z�_o�0�|����7S�,�mHD5U<�Z�CNJ���a���y^)����SE�04���
�~�>:�y��a�=�,�l�y��H�b�<����d�tg�������^��0��>���a��� ��ԍ+-�����މ	XH�T ��ވa�+B7��@B�r9Ȉa�o� �ӤB�����g�ܬ�,t���(1t@z�����Ւ
��>Ȉa��ZRp�*S���1�D����o��/��LF��5`p�������`��JŞ�м"��T;��rO���@d�0�����
#�u�[`	�*�*�I+�<VFC�-�@��W�,�Sd{��^s�C9o�a0�I�$G�y��?��a(���i�f� ��a$!.H�2�|<>��H�_A�*0�1�:���'Dw��"�A���R��{�,#���)yH+�a>���H�.���9I�L��"b��0.`uX}�Ï1ZC�����=�����:tCLR��T~àU��
�WF��v1�A5`�q%|R�HJ��,��4-�v�y3r
8���W�o�a��PI�,ر�F��e�I�:S)���Ak���2:�"��-0Z�<�D�g��sSà�����������yC�}_cR��>���|MAE��>H(`�i�k*b���_Ae�O�gY�&�"��O��@���1���BE��)x�R��ރS�������x��OY�:ӾN�"�Q���p�W�l<o�aEw/>D@�;�U��8*bEy��K�t1�x#�Q��^ri�~�=o�a,(���8��vz=�F�~�!�T��G��y��Tg����0
��?'��Ǩ�6#��v��/����/߈aa]0�B���X1�,0hHj�*b���^��@�P�R�`��0h܊���a�~�O��\�n��>1��9��t9�y��(k���7S*6{���е��`�' ���#��pm~o`��`0�sH1�Ί���{Aj�uRGC��Ҥޤ1��8UGC����T�����a4}7U`p1'��up1r���K�ky����g:b�|*��^$�uC~� /1Lx�����g:b�qo�#�q)�;�h�>^5�i�b�3���a�^�Oa)�
$�g�7bL!y �GP�i��-bL�|��y� H���1�PޭhE�<I�sވah
xU��Q��c1C�FS�ɏ��w�1�~R�TC�1KG�)����ݐ�r���a�<��C87#��/t�0T����i±y��#��!�j��?��M�wL�0�>���[�U�L�0hUAa(��Wf�^J��0huO�2Q��U��(B𴆊$���+ӷ�x]7�P�wx����t'�-0�zC7��0��y1�f��>��I+<^7�P��;�$�{�D��"��V$���SP�e1�c�Fp�H��&b�
�4�
�M�P���-b�J_7d��|�Dcx�쀀����j=~�à5�����p ��^'M�0��K����㐉*lP�d��&b�߇�TW�����>U�ݕ�a��W.�u���;��F�1 ���&b0J�@NH��xC���� �I��}��Dc�{����k�����DCu�`8�Ӡ}�a�
*�=�F�c|��D���zhv:�q�0����w����R�ve#�!��^+��QXl�-0dX:�V�[�AFxc�1e�!y T�9[��)|�l҄q��ue1��/��l�O����xa#�J�>�b���EK�Ҭ�-0�ʐgY��#?�Kp���06sϸs�4�4��h#���4l��C�|l������\�#97�y��A$�BH�y��t���җ���s�P?e>^f���}/,�y?��S��>Y��
Q����-0��Jc�P��;��[l�0�A�0�^�2��8��X�ҍ��B��7�I1��YAH#U�Fj#���c���.Hӕ�-0�h��?�q���ECu��7v�����ك�MgA|���6b��p���0N*�-bk�2=�N8Һ�Q�[`K���y+?�Y6��.Z���k��պ�3^�N��� WuQ���   	pHYs  %  %IR$�   �eXIfII*     (           >       F   i�    N       %     %      �    T  �    p  ��    x       ASCII   Screenshot(/��  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:exif="http://ns.adobe.com/exif/1.0/">
         <exif:PixelYDimension>1392</exif:PixelYDimension>
         <exif:PixelXDimension>340</exif:PixelXDimension>
         <exif:UserComment>Screenshot</exif:UserComment>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
����  ��IDATx�콉�۸�%�R.��֝������_��V���$�XND ���t��v�R���+6�0�����e-k��IkY�Zֲ�)+��e-kY��Pײ�����
�kY�Z��BeԵ�e-ky���Z�/����W�E*������+?�Wj������Z�^�#�� )��~�:��^T�#��J�_��m�P�B���kP�? �����S�מ���{������)��⽭����
�ky^9Ÿ�2��S����,�������.�[m-g����k��6�y?Q���������S"�)�h�;�/�����b�<&;���%�+U%�Y`��$��\䬲2������W����b�����m�.�z9Su���dEȿ\Yu-�+-�{�H�8E-�粒�K!���ŵ��.�:�{��r������31���Bos0]�YU�[9y�s�t:O�%��F�tc�����
�kyvy*�����<�g^N�W �"ߺ�9&���H�6z�~�iE��<W���oVV@]˓�S���cs%�/���ߜ�ܮ2V4�-3[P�>��\�g���M��nN�ƧQ���GY��
��
�k9Z�#���T欴����F�RZ]�S���k��Z5�Ci5����=��aHc�:���yb�y�o'x[�[x���UAG��&����*`e�߽���/O��S����#8T`Z�E@52Z�tx�~�����oT�qt�Y�K�}�3u�]� :����^=�����O�-�>}_O���x��Ȫaϫ��y�c^c+�����Zf���R����@[�1�$L�t,�E��@�X����2��~�����z){e0�ۇ�0�Ff�1���
38�
���
��Yg��L ����T����]�������9�+X�sw8Wf�� LNc9���РZ�9�]��-+���*?`���&s���1͆5���6=���"3@tz?iا��F���v>f,�r�d��M}S)���O����|���ӹg�I���#q� :A*P��AX�&m�f�]`�`���I�(�����^��ȼ}�?Rl&��n���m�й	��k%hg��4ь���F�'�"O�W�ݨ��+�~Ӳ�Z�� '�E12Zׅ0f��
	���0��DxگT0H�~�^��A�*��L�DPX�\�^�T����T�RJ}���cLZ���m�S���f#�&��lz=Q2F�c����$i _������jI]@������B���K�Q��u��YV@]���`Nk<b�:� I���4�Y2;$ #�y�,P�03�����o4 �R��@�JA�)	"�� ���=L�c�+(UlGPG�Z���>ȬC��.9 e~|�6�N�7�}N� u 8�#�8Y'��m���L����F�&��
@s�^k�>eԵp?˩f;P��=K�O��e"���l�>*�ƫ���HA� f|���}��q<Ui�����&p�
��z z�*!��&�a�ߎʂ�32��ޕҵ������'?��*e�T�N����Q�i�6�z�L����n {A�f�1|M�+���+�buV�}ղ�Z�D�(�Q��@�%,rd�0���Yԇai PԖ�����W},t��e�S4��#�c��Nu��Ã ��+Z����2Tk�&+Ƨ͸��ઈE5��TL'���v��m�y�z�}/`K���2�����q�ir �zXUf�[V�~�@�T|��h�򊨯ZV@������	L�k��a�zI��P�'�0T#���u>��d�5
��k�^�؞��C TX�s�h��v�J��O�}�ɋ>��Z�[ֻ�(�2c{���i؎Vo��(D�SV�V+�����J��*��ꔉq�;��AuQT~)S���w�%C�f:�6���^ky��Z�D�aQ0�����ab{�P	0Х&��� ��Ea0��jPu@Ы�1�99��~�*�J�g#���=Rd�������d@X�>L��^ݜ.JӺ]���ưN�h��Y��_��+�0S�t�D!��=�kݧ���U �R/��xq���b����
�߮���/e�;ܞL7�M��92 �u�Q�z�J��`��3�b�����	�*�=7�������H&�:�x>��9�>s<ʂ��o$P%�?�������~,�@�R��r�U{��܇�ɹz��E���aL�� �J��6$L,��>V������nY�g.�2B��?�^S�QHSv��#�� Jb=1у�U<UW	�����۲n#+�iw����Y+K݋�lT��t���!y��a��9�>�=��x1X��3�Q�80��MM�_���cF�mb�}�w�/b��c�.]�B�K�����jˬ[_=Id���|;�*��C]�u�
�?k�
�'���Y��Q4�(�򧴟���CuT_Tb�����h>
uU@1��W��(�H�%����>�u����p ���BDwڣ�R�^ҝZ}��:���� M`�ƻ� /��6,5�*'�[8j�PO��%K�e1١W�t"_��I`�%���.��#�����'�^A���
��r&S��	#�3Ճ���M����������\�9�ol|�&nT' �]�;+����'��A��8�ٿ�\��''꣆�	����F��M2��s�SWj&Y}�AY?���<	e� �~�Ć�"Ʋ���82H�w�����E��Sz�≡�9�N+��NY�g-O��njY�	"^N#�\���$�!�8�a0���
|2�Q��x*`nD��X�+e#����4�L�Y�2f���HH��[���Do�^ �aol�a���j ��L@8�> �q�4�Bn��ս�M��^���U�oj/u��Q�F1��'�8�'VWկ++���%?o�,�:̪���h��i�������Sa�c�cnY�k@M����(�@�O���vy������\
pe�:֬���f� FuIvy��0��Ԩ>�x����_[�]@F�B�R�-�/��P����>?���8��ꞥ�4!� �^���h�����n'F�}����hp��ak*���	�&�����>ki�
����Nr��_��}�1�k>�AY'{  >?	 r|� �-ؽ�xS	��p�,�	Os�5kz�4tp���r��r��Дx���*�j&S�&�l̐� ���ɋ�����v�s�S;h��D ��9j�*Wq����̵��j��Wb���21j�~��t?�S{���ty}�����U�fe٥ ��7���Ze��O*+�����c@��g��TFX����Y�`Qgq�#SQ7)=n���}����%"����	Q��X�$K�k�~�Y��3�k}�VZ�
�NPQ�;��X�W���دS3A���\�UJn���FV��%0����	�&�X/˾��`A�N�<�� 5�8�UY>����"�.��X5���f��r�bi����eԵ,���t|�j�q_�=����c��M���&X�ᜯ`ZԪn��z,�j��������+�Q�;��v{�W��>s����f�����q;	�b�g&��7��^�F���aC�6&=h E�̘|a!�w4�l����q������+��zӵ�\Yu-GXf�Q0����}���(!wib�(ْ(��%*�N��Pr��2�Ә��A�� �� �u$*�of�RJ�p�NQ� ��#�c��swY��H�/Ġ��TǤ���t��,s��vX�
��؍�t�R�6u�_��x�+׊�߶������@�O)\��yj��'}Cuf	v�Qu������O�Ы%^�7 V}7�X��w�^����t�=��"�3 �3v�5˾f����@8��~���$�_ �3���@�G5��<����(��Pw�i����n����35��y�q�y[xҘUN�VeԵ�,5���A�;��ߖ	z�h@J�Y������"�����>�q��a!��7��!u�f�,��f�Ϋ+�{Bl�<����p�&ɐO�ˆ�N:\� �����4w�����8Հ6�S\��Shg�6)���`[�ۘ#��0�@uk������Vl}��ZN���q��wџ�����0È�-,�A��PŵI���� 9�rT��.��T`�����ד�4�9���k�j�Pz�$������L�9��R���ަϟ?���/�V׵�TCӨ*�r��c�F-�K�Q�keF����H��c������>��
�C�E}[~�y�+��nYu-��`��>~���nM`c�6���{H���>]^\�w����Ǐ�N��ٌC�ܬ]j��V��U@�u��y9�+�z)Y�9I�Vr�v�(�7�v���.�����?�d`=��T�ڲn���;��(1���"�z&��v��d��&�3hCe MA0��$�	����X.̳ %j��VM���P���v���:�U0��&s��-�3�kj>�K��~�>M`����]@��;u�Z�0��KՔ ��VD,�jb��W��J7[] �Y��ڑ�܎(��/�>ML���*���wϠ��\�b��u��	#0�W���1�� �3��J�b��龓�`��A�c��X?�Z$⦝b�W)+����=*0����I�����9{K����s�!92�1?�?��/�����ҧ	��M ���]�%�ذ��{��kg~��f�A��EO�ܫ����sC�?����U����1��L��	`�'P%VJ@�ɬx��32r��ov�`-� ����D��Gne	� ����b1V�6JFO]�4�
�/ZV@]��3W�A-����F��]��K�5�U;�2}}9��O�" %y=����W���N@K�U��?쒪X�F���X�Պ�Pw���~�ji���1�ը�h��t�� ���2K=�������y��Z���b.]b�ww��N@�W4��^#�,�`VՉ~6^د�X��چ{_�R�^V@]˓J���6%�G0�@@��܌�j����?�g6�)���/����h:
K��Sā\�r��`ѺXڹ�<7���k@��� � @��(BE���r0%����;�����3�U���/_җ�M��QX!�Qb�UG�����7�@L��î���
�k��A�8rɦT��h0�G�cԳx22}x������0�n���-m���C Q�ya�ǳy�j���>�l�	��N�{�Q��='������g5P��E���,����������/�y;�#�z�Yu2�ʪ�D��P��q�Z�aq������������Z--;4�I��;Ď&������_>��������l�����?�;�B߫�ig,ѭ��k�����XfZ�����\c��xG+�X�����y$�|�.�M���[���gw��j�LSYWP:m|*�,�9�IV����
�kyva��A���g����=�ǿ���믿N`�^���Q@ S�z�{�������^������	rmS��a�t���_��c��� �[Rn�Nd��u�r�Ng��VV��eԵ<��(��f��Tt�M���@���w3��>L�)����`
 -&��7ʤr0�����0K ���l��5�p8C'�Y���+�(�7� ��{%�]�T�'uK�ٯbkU���Vd-/TV@]˳
'�`8ʒ�sԤΚI��x�����4��-�6b����"��1��_
�	a���ˉ��g��텄���L�3M��������s#O/˲�/+���YE��� n�zM�D�R�Zԭh��O��r�oލR}#g�3.����_KP�:����ID� 5�!�Ԧ�!Am�EuGPV]��)�Ϊ
���/��|}Yu-g��2��12��>��_\hb�1Sƭ��	'�3��^�z��^�%�Tƺ]�dݒ��MKA��TS�^\�bV���SUk��L��Z^�����g�����8y�c� ��E3�5�Mԗ�ʄ�9��o�N��>~�-����l��3��fw1�Q���3*�b�$�ww�@�Z��g�P������^ˋ�P��ҳ�~ga��E,ۙ�K���q�aj3�Yu�l9���MY82��*�Ю�9 ��VI@�ȗ���nnnd�BՍ"�ku������p���FYu-�*+���6 v�5[u���fqMa������0�#*� �c������^Q��H
���޽���?��$-Q̷����w��	<����lX�ox-�QV@]��:��R,�S����r��5>��Kiu��aJ���~�-���c��|d‵�U	��)k�9 �^� �D��ޞA\R�&0�lu�p����b�.6[[Rf՛�nYu-GJ͛\�T&4J^҃f��]ɡ�ܤ8����)�S��2|d���qx�s|}�L�U�.m��Q��=,�ਫo[^vE2s��4�J��Q�Xue;Lu�w/�W�/�$�'O	��������m?�7QV@�K����ϩ�Zg�w}(ńS�����d|!��t}}/ ��d�j��i�Z�I�\��o������ˀ����/]�pػ�D3E�骪��y�괝���P�O���Zib�K�vͱz�QH8j��1�w/+��e�1�OYP�|�P���.���3��$��G]ET+X��s�֗��&F����R�ѭ-���8�C�錴'N�M�d'@���~8p�n���jU�w��ny�� �U����2�OS�b�rnYu-M)�w�1%���e���ձR'ǧ7��@�]�G��W c��c�[���6[ ��v�J#�S
����EO4�w�
�!�
�k��`��H9nM��q��$�֤� �ܞ~����L2��`�	5�d,W=�Ǵ��_V@]��%lHݗcZ%�AX�D^j�z�%Jx_&*_ƛ�MN!��uԩOk��eԵ�J��z6����<=#�3P6Q� �#�ܲ��b�L���V�f�2ʮP��,��r>�͢']i��)+��EKT�	�*��ſZU����x6��j^���?cy���6�-=������b.Tk��)+���*�rѣ/�=^Ԭ����9�^��.2C�|���D)�>Z�oH;��5���t��Z��/+��%��O�������H�U\AU���y�ρ�W�8������ ��.��ujߢ~��<�N���*����Z�(=�R����{��T]�h����e��K���	e�49q>Y��U/#���QJZ�(+��%��^>�f~�) �g��-a?��	Q8R@@�T.���K���4�q�XF�Qu������7�0sn[!���P�R�*Yq�cb���MD~�������)(?���הe�_3��Q�/I�$$�'���1������Z�E������:�~�Ė�*'�;��,�G@5bK���U��^�J�q*�t���5IbiZ�g���bv�@\�;�+�u��5�
�kI� ��a�#X&Cj��=i��<ߗ�p�O�a��S7����}�"W����Ɇ*I
B٨�d)�W�>�U��k:e�#��e�!�g͉���8MH��?������1�QB�T8
�tӬ�%M�g��sr�1 m�tmVKky���ZB����V\�ޟqJ�&��ђǷ���ߥ���M[��:=H��O�E�+����4��Z�٧���;�.5&a���/��ۻ������U�h6F�҈ﯮ�����C.�Q_�����gЇI5FDl��$�Po��~��1a]O�H>=�E���5�r���?j1��X�Y�e	�����1j�~��'�����n� ^�Rٳ���<�D@�gs��T�Z[�S�mYu-�.4Xm	���j4!@�����/����{U$:�tq�d	 �蔱Q~O[�*�M����
Ƽ����)��a����s�׿����P�,�k�=by��M׫��h���ީ߶����g[;*�`@����"������-:�w,��c���
�?p���at�6̒��
1Qb��O�MH�7���6ݨ���#��3zc�wK���oRV@]˳�XĘ��:.��EJ�~�����	DiI����������΃LJ-kc=k�9
G�M���;1�>�Eh�م�'N�������ϟYM�T�� �IE�d�Pb��K�P[�������'ʏ<�����g�����72If�Q�SY��J�o�>�T*��I�puy�����XE�8�l��?��^�b��6��1�Ll������f$�qoT}2��8q��r;�<�* �Tz]T �!��u�
�kyV���TG��,H�DYұ�����ۋ-9}ާ�>�뉹r����?�طD�p��bL��"���p�`����g�����ݝ���(���RK�W���t�ky��S��$j<�^��X�d��2�n=I��w���~zu��yi�/7�׿��>}�ȫr^\\�Rǅ+z�L��
/���ӷ�[aϊ�N�vj��4��M��?������N��zg�0K�/�Y(G��&6Q�m/�ar���*��ɬU��疷4nj@�i�eU��������/�Nn@����@�6}��O1V]���֞�L��o%]k߉���.R���ŢɆ2�B{Nm�ۿ~K����͠J�I�
�)��e���
�9c9ѭ
�)c�����F;�^V@]�3����Q}(Ch*�N���n����N��ߥ/��ӻ�k��__]����һ����w�����ߜ���-�׹�OJ��� �������a�����F�|�)�3j�~��U0���/9'���=���Q�vY�(�!��7�����T;��YC�x�"�N�F��<"�&۲'{>�yx����<�F��0��IEa���Kf����˧O�Ç��g����Y 0>O��_��O.��0�(�e�:җ����������Lc�>�OV���,xMPȮ�ib�Su�>�����e4v*�W�.D���,��Hk,%m9�d�Y�;fy���7H�_PC��,����vé���J��Ի��W�4���}^���8*�'4u4���T���t�k㿙�N���O��*��mTv�Q>c}b��b�~����8[Rǋ��b_i7���~z�������K���[���;V���)��9�|�������Bg!�C�I�x�ډBI)�>1�/7_�����>�Ko���~��]Y;j��(י�c����v;MBW�ӧ_�I�C���ּ�F�V+Ћ=.�cT��O�鬛����q��p�:wdDپ!թ���2����縢̧�� ��K-������8��b��N<��I��R��|
u�C;��,��FBp�>�vNef�"�m!��Xr��˒pH	�Db��9��}7�GvP'������J/&�~��h���t��p�Ʃ.{�_�~��"� �Xv�xUR�j������S��:��g3��)g���9Kg�"���7�˗/���n(F���q:�����uY� �g6h��=�F	��tu}�>~���׿�=���_9���X?���(�?�����S{S��\jm������ ���I<߈�Wo���L��U��s�"4z@ ��@���ѷ��%z2+0����N-�^�L� p������U���j	��-1t��vKK��d#h���n�<Qo7%W�a�;?ed�8��PDI	C�$ȝ�[/.�	'f��/�;%q.A��'༘@�D���{v#���y�Olubg��_%�Y�5�]���6����g�C�"F>d���{I���w�N&֗�OߧɈ���ECmyr�	���[�]�V@�� 3�T����ԾW8�ي��|Y\��Ѯ=o���_�1JO-���޶ ���A'����tt��x���R;3���U����S�?�+�Y�+W,U��O��č8��7p��[u������7~|��A��l_+B��� ♁��1�K��4�qRp#�Q�ԩi@�tK �����Yw�NR�� �� ������_�6�����ω=�w�yֻjl:��(��2����.�劮7*S��>	"mN=�1��;;؟<0��N�Gq#@� �d�}�u/1��d�Ԏ���u�Id��&��Kn[ *M�^�~��ݥTCv/�F��h�:j:���������J�H����R�9����3ڱ�.�.��N:�N����i�^��I�"R$߹���
���Q��.�1�t
��p��\Y��%KY�@�t>�V�W�� ����X��Y��[�q�3�쳯���xQ{^L���I�><���
T	�4����	U ���}����T���|�T�	Ǡa�\{dT76Ą��! 3��ª9kTVJɶ%���x�R����$Hf����n�����.a)ӣk�$�6X+OgN E��3`�X;�>�'�R�5��Nz�<��Hi�OU����r�?, }`
#��_� o\��9��^�@���Iy@�Yf0P�b����yǏG�5y����+�\�s�\6@� V��ض��x�a}��:����H����ދF�q=���kre�28w?�'��4\��+�h��	H�w��Y����{)��wiV�:a�����[���Uyb�@霱)�I}j���&:]�$�����6��q���[GF�Sb@ꅹwj�g��`�k��K����9I��44�#�N�t�,5���#�DVZ�����5�=��c��GH���,���b"	���Ԍ�ţ�_��D���^j�e�Ҏ�]Y��ce^�q,�9�u��L�����BK�C- ��T�}����uD.N�E�E�TD��E�٨���Tuˤ&[}��<���o�W��30H��:+�'��'����5�p�T-ꐔ�{G�+Y\�Xt�2`O�l� ��f���ML V�3n&Pl��ܱ�	��TA�a�TW��j����̾�*9Y��ҡ��@����y�����̛(/���:�y���Cl`P @<�Ɖ�r:�3ƚW�.A�/~^bKK��F�_��T��C��zܑm%��}Yط�ޞa����8�|����/ׁ�Xerյ�a�c�c���E�/����R����a��R¬o��	<�Ȥ��}%��]ۑ\�R�)[;��ψA��V�� �*�^�7|��P__�'2�#1��r?ZÝOH�$b�lBxrc�|DG]���/X3�س���|V�ey1@E�!��l��'obW��h�o���#_�\�1�c�wv��>�T�m�`/2��Z��1��zC������&�����1�	�_��Q�5H`�ͺj�l���� �-"�Nܳ�����]���!���3��<�tA����F)���0#��1��I@R��z�M���1c�N�Af:�P�y����52Կ���;πG���1ql�G�.��%�J�q�nv��+�����/*�cq�)�d�ŵ.k���\���ŷ�*fb�.7<���Ͱ7E�D��k/t��G�d�'��稾�A�Vo�0�þ��ƄΗ'�z�%uGJ��O�*��{�p���۬KR�b�fpʝ�`(�����~�:�6���0Hv'����u{6��B�V���YH�卬��;{���S0~���z�����j��e��I���+��@=!��1�Wڥ0��������m�<໗�Tk
ի�c�0��Y�s��+߇q>�G�k]��":Μ��R����+��=��&�B��Ĕ\�D�-#������ ��u�ڛ���������Z<.2V����1W�x[(Ě���٩�� ��E�3V�pP=���v�T hT��*��k���%�/��\4+-H�P�Z�ɥa��d}z��:�Q:��"�9���u-#EI�3�d��c�?�y��Q���硄�v���K��Xz������P��j)�Qt�\R�(貦~��GQ	�dl�1t�J��Ԓf@cU�W;8��V�L1�DT',��D�Z��l�GJ��Ei�5���%2��銁�ٰT]mS��i�"J$�)̔\���W��&�7�0YCTY�J����@f�#IAَ�@���JT15�EW��*F"84"|d�&�4�(���ˋ>J�)4{��E���m�>�1�)�O�i����;j��RUÁ�I��f�=��>�0j+�����U��r��E�E�P�ndP1K�^siZg�
�480� �Ć�f����[�x���-͜y@��u,uL�f�#�w��B���o'�՜v�zv�MK:�xYc�%N�\a���6��^�:�QYc������'�ր*��%�'^�u.��Z���Z	�(�J?��L�}"����	�f<�O˽i?���`�� �uס\��6w�>@v�O�'*��� -��ȟZj#W8G�� �-�]��::��N���RyQ@��!sg$�|��"l����e�ΒC�l���f`��yE����g��<Х-%���,c?����q��!�tq��3�~��p��ejev\	2�rr7�VuPлFܿ�J����7~��:a����3�O��������[`�Z�3�d�H��v���I�~��x�ݜ�J���
�biu/�$$-������g�ɟ]Q@���K\
	��&����$E>�q�¾~�%lu���D%�8��*���%šw�A9[��QTꞻ��u��nd"��Ȝ�a$�cy��	b�h�V����-��Y��_�2X'���%t��� �4�`�i�$'M�G�[9ׇ1��e�5tXڿ�~�2�����Ъ����ĦP���xn�s� �ܕV�A��;7�`b��0$�Ʉc�*|+��+*=�J��� 5�~��C��&� �a,8OP�t�3�59�4fێt�v�sT�D��h��N��A�#�J�(k=l���97�U�@�,p�j��)���ⓗ�9C����c�	.�D�6(ĝa�ib��������#��>�B�:e�����*�ޔ��\���A;���E$K��6nu�K�qڧ k�qm�!��ӛ���<�euLa+�	�<��tT8��&b9d������D�B�J2v���ı�:d	X�&�>�?����Ʊ�-�OJu?��Z�v���l#kT���C?̼�(6;�/v6;U�^OX���T��{�E�!<}�|�:밦�1�9��3��0l9��Y$֝*(V���ƅ#EX��$�".��.���^���z�5�3�)Fu�ȥŪGJ��?c��,�Pf����������Y-f��ji���NU����.}�h��9��J% ,�I��R�L1&A����ڤ��z��Vf׋�`'��T��7UEu]�y�J�3�?� x��/��k���UW0NX�x�yS8fh�{�����Z&�(�QQY��M����=؃c�qx~{o���֓b��i���Qvvx�52:#�̐����U؈�z��Pq3�.�rn��.T̠��_�l��e�b@�װ��~z��r�9py#7�R�x-����@q
PS��L��@)�
�RԨ΀��d���`�hñ��ز��Ȯ#&f�h\����m[�K����:ɽE7��ڗz�v�c3~x������Ȧ0!`��Zo�7�5`ܭA/2��>��6�ЊU����aJ�]�[ĵI�����P��<tϷ�/��s�E��0�\���%)�����0�U$&i���Q\)�����2Z���" m-�fU��}cG�iZ ]pW,���\c��Ů��@��Nc�ǧ\u�Ȏ�D�ܴ�P& s�yjo.~�v"C�{�I��<�#,�0B���=W�F�n��ߍ�Z�
/��a�Uv*��U��Ǚ'�7Pm2�ve�����u�^|ib;��i��k%n��	�Ŗ&�F���O�F�ؚ�����CP���!b,ٖݡ��!� έ;@7J:�T{	|��:	��@4��aS�?3�A"�x�$l�b6�Z&���	�������R���9ӏ�"yj0��Sx֔a9'h-���!CՓ'i�z5��S�sZ:�ߓ3:��_��=8��h~ן���Tgt�{k�%�}�q�,J��4�/.@n$$ת�V����NA��݃�mۏ�D�HT��<U�r��~F<��y�7J81�g��Śq�MO�U�f�gL��y&����wl�G�����O�y���@:*�w˾r���f0�8����i����e�P�OI�1��N�I@G��ҩ�;y�����Yg�.���a�`T(VQZ�^���A�=OdKRe�L�x�e��n5�+�Y�k�t���Q�-� Z긕�"f=�gc��ߖ���a�S���`z���	O���8��x�����B��r)��5B8�ee��|YC�0�g_�7��%� L�xfG�<G۽�V2���.�ٺ��.S7¯��@�k��Z�4C8|�2\�E�pb�4!&�F�4��F��g��ߤ|5���):H0Ń�O$�ګC�����T������e�I�x���:( sS�$0�
���n�Y7��8�� zUѱM���Bu�z�,Z��~�����6"֢.t�U=���y��B���k����RW��p��"�*��6�>aǥW���+�v���~z�>3���@��>l�j�(2�@Ҥ1c�s�Y����:�����2Q�%�����CZ@�zKX�lq�ȈӼ}t��m�*w�S�j�>��������ƖT��R^\�g����.�G:jC��^40���K�I�IJ3�V���$'���_2}	K����������� ��ʒG���=G��ZGAbq���L߫m�t��3W��Nv��G�]�CտEXZ����G�/�r�8��B0J�>���>��U��L�;^�	҄��]ib�~â?9�[�Wq�S2Ј5ok�%ֳi��0���W��%��z��\���'c���. ���xȚOKU�l֯:~~�`�Kg��d�����<�*����A�s�{Z��+=&�1��ɹoI��xnէuj}�n�@��i���E�p#`BU#���I��(Ɵ��A�mJG���ޞ`_Ǻ����i�u;y
� �P1�y=�2" =��z�sPe����Iq�G$ 3��A ]C)����~�KP[��rw����`���Ae�Y�k�j�x+0�=h?�/_1�q�\��ЎK�ij��U}V���&|��J��_�������ұJ�X,�֚y1H��R��F|(�!�����o�T�H�����(������ˢ�=(��G~�"�[?W�BkŴR�����ٮ1(��Ϭ�H�����2K�|l�X9s_A�-9�PN�0�8x�}�2�>Z��+=�2������ o��-�@��sn]/9��V��&o�a�QZ��֮���c�0�s�i��*�������=[}XdWi3��H'�t,�p䙟�R��?�f[I6����C�_Gn��c]�r���G����.d��D�0�Uq�:X]�%O�J��Y���+���o���wؗg�yd�̗P � h�� ӂ�#��Ig>���EQ�~�$:�]�����M�����_��߶�6Z�8�Da�nd����E�WUf ^�!������CCsZ�w͘�\����+Ku�V�����H��W��u�z*�:�rݮ������b� ��$U�4���8�glمʏ�V�lr�2�o1|x6����pK0Yg,e�!|l�?Tq�������Íu�b�_5��=ZC�V0�0Ք�M�3�LXT9kNd<)L��#
��<�rՌ�ab���8����L��N��"�P��ZG~	�|�R�F�L)>��Z<9�=����(�(������+u���,`�5$�͹�d�P�ZJ�:�������"R�e�+��Ѵ�}@��:��K$A�am]"B�u� B=0�yN=_�-�1v�"��D�k��Ɩ��6�n/�;���E�h�Q^I�K��k�;H���t�]6 X�O���S�S���Xfl�c�H��n���=�����b�g^F&c�YMP� Q��yT���fnP:eU'-�;ة�.g�L�z���$,!-}[l2d��~L
�Ơ�B�x����:f즶w)�bT���n�y���yZ,����Dm�oZ�����E�N₇N��lܠ�j��4d�T�m�}���[�<8��A�z��q>k��js�|%�������� �4yb� ����+^����f��� ���N2�嶽rʆ$94��;�<zL|V,�&]>�����E�J�W���X�3�W}Xo�<�s��ļ�	B�'��
i`�����1	�����W��OGx0��,�nNf����˞���Lr+�F�L,���]dr�	���+�̉Z�P�& uum0D�! m�e����<g8�[~D�<�,�^Ȫ�)�x���2�^]_ْ��Z�����7Kf��:�(f�9�����[�Η}"_b�KZ�g�܌$om�:C��I?�?�߾�N�0r��ʸ���.�#C��ߵ��+��4�T�'ХY�"\
�u2#���]���M777lp��d�%��Xa�����ѻ����[k&x�)��"���"p�K�F�4|2�J��r�9?�������#/��/z������xz�p߽7���,���ޥ�������X��u;�wf�z�#,�:�\��%�k�}�K��	>�� �4�O���5-�Y���Mw��[/�����L&�ƫ���{(C�Y^P##�34�x�ۗ6���$GxxxH7�`���?T	 �}4Ηz�.�5�@t��@�Y�'��I/���R��>�0�g"ѷ ��QX�#\�V�~L)�a�/|�9�qӛ>���{�C�܏�ՖUn�1����hr��=z/��W+�s=��Z�/+I�,��#z.����s�@ ����5�|ʽǱ��g���x��BWP��4���2nDh� ��R�-�b9]P���/_���F�D~�q��~�u�N���D��3�a�P��D���k���m�����ׅ>��=P�ds�A���S�i5J1A�5@m%�;��I�!0ݫS�K�Kꉐ�E0�ܼ���'o�b���=E��Xl��eM��È��Aк�&S����r�ֶ����W�_-��1�tQL}�lح�oR���o5<wG�F�F��`��]g: ��I@J�h$���!��%�*��P�ak�k��a��#W���"�֚%$�tN�٠�_��Gˏ#�~���	 "[�Ҥzq)z��v���COYo���+H�-��W�s����o)��%��z� ������(sO�B�%��m�`��z�w�}�Ep0���}�]�o'̷^^P��a6G�X�H�4_��4�_י
�X'��I��1X��Aj�7i�b�E�����|��AZ�UK}�ӓ�3:ӷa�g�Ο�i�sp�gO����R�#�i��qTGF�HP���>�LsAy����=���m,���۹m��<b~�K
���ā�V۲��
+�\��Z&�׿������RS�)�7Z^	Pk񽠃B��E>�*Gꇅ�zU��N`J/b&P�\��W�6��uᅙ��o��=ٯ�&kR�cSƷЉ�=��%��>��K5·��D����H4M�S�h� ��/z�V�m�S�n�o�\	��KJ)?������)��d��v��]jGXѳ�v��(��\{;$�H��k��cSj}yQo���6|��Z�]g��>�h@㳦O���Ld��AA:2z���RI�'Cd��+;��-$��`�(�rhڃ͞��( ƙ�"�٘���V�z�{n9���^���j�Ƨ=3S]B9H;��X.p|�Ν��k���L�*�M���������9��9�'0�Zǚ0�*V�����G�63J�ȟ�1=;\̏#��˷u���kP$����;z1��;[e$Ѓ� ��pq�ۋ��$�$�H��<x
������gx��cS����+o&ϴI}�@)���1�_�������U���3����J=Ѿ9���F�9��9=
����]��R|z _4nW��U]��ŝ�R���G�[J����J�������O.��;���t����k򵋺`TBH����~N0M�dz���֙kY���0�	��K%�>u��hb���R�7O,���)3<�~��-�tT�N̔b�1!��G����T�篪�p3a=�C=�)���)�OX1�@�Dz�	W���U����}�3W���=�Q�+P1,��gi����і�3�ŒF#��egO.�/v^9<���z�}��M$���A�8?*Ysa�E.Ƹ�4= 
U%� ~��S	�GY�%��t�
@��}��;�Z�?>�� ��c��{Y�M<N���\���d�l�R��`|���y�`�BES\�CN=D�K���>�6�g''���dv��~-�urX��/��ҋ�/�S\�o���&?LqP��2��5|61g�G�6�~�D	����i�~_(`���0Tnw����Dz�%�:4z��>Z�T�(b�m:5�~V0X��S��F���@#Y�S�c����n���Ae��%'��9�?��4��D9bx���!1=6���H?A� R쁅�*�v�.�(����L�p��zۥ,���+i]�.�>�V�Y����!qK݄:�u}��@z�.n�r܈���= 42�ri3V�-��o�C}�R�r��ܿ����@�Y�F˘%� ���,a�~N m��&��_~/�ԏP^]/'�%��#%1�k�i�G۽������T0��@'���S#eأ�LL��  @�����}!��י��Nc��h��Z��,��R��*\����Bg�Ԓ�]}�5���B�n���l����_������������
�?��⓸55�FX�JN��?����Ӛ����F���gc��?I?b��g�_'�d}���Z�c �?����yY8ƪը�$w��l�G��.��J�����6b�QO�3��bے�������,�P��l�d�ʪ7���
L�/�.�}ʑ� Lt�)��X�1C@��t�K���@�'u�h�,�����[^���{L��%�窶�X���J���U3�㾩��1����:���
�E ����c������i4tp�k`��N5Xx����VE>�d�ҳ�r_Ͱ�e�(��-��HQ�*�G�	:� �w�5�fj��6 K^�no�^������1��*6VEA}ͣ:��?F0爥m�T����@����>>�ϒo�O���(/�P]��6cs�MӳX�gL��b27'������M,u�~����=e7�~S�R�dY`��}5��0�k$�5�����8�ˢܿ>��4>a��������Q{�#"?B�cݾ�,��0������+	�H���g����F�֡�W�������j ���J��e��RZO�BL�Б�l���$�/�������ʱ��O=�����
��翻�*;u��$)N	��Q��|�W��ȿ���Q����8��oE}�3�Ғm�g��S^PӞJy�d���g��K�G�a+��K�`U�p�ol�s&���ĵ���~n �~����=��A-3�����3 ���X��;��
9 X�P����V�:-��H�Ρ(��o����DQ��K��a���!����X��/�	���m50T���z'���� ��1�XT[�l�7;�w�z�~d����"3�`\h��|Yv�[�ZX.����V�z6�>Z�X��4��!�x�t4��2n+�,꣼�c4F5�)��#�\�~�R�M������5��f��&/�"�zf2���b"U+�G~\��^�0�����m��+�\�F�O־b���f&�/a���Y�yb�K��ۋ�U�������iN���͗�(�'����ﳨ�3IC�|�(��y�K����0�^Nb�ks�����$yȒ��꠫�R|>]�3d��~�T	�ru���Z+AKP��"�&�dm��z�B����'����'H��-�WQ��{X��O�\�'���z|����]ߚ���:��-4���j��n��8���j<[IFm���=ӳ���җ½�x;�3֣������לZ5��_�$=���&Ss�֐�f�Rr�lE\#3]f�U�ٱ����m��}X�8�������o�_L�/����K8[�}CF��:�
c�X�����{�Dҳ�~E2�K�j���.%/���fp�����qH�"�x.Id��C.XS5�юY@���Sr��yL�b �����#�j�-��$΄s���b	����+O�Fot�q'� �?귣e�.a�������I	�t{�uIU�������fle���^��Eqd���x�U�.�{X�A9�L,��AG8Ez�@�=	��P�M'�Ғ�wdB�;�S�[�t'��h�:[_�	��z�ԅa�[]���;:A�!����	�DD���96��y�d��<�^$�m���+zfo����C�X��8yHHH!�+�rWEX�vƜ��o�l9-ufOYO��%��ӘI,$p����+�"��̞��	:��v�r~GΚx�I��'�}Z��d�K�r�߳e��DPѶ��js���R����KEX���G� ���8� o�����Pbg�,�(��^�γ=�$��O&�φà˭'I�S�ֱX㩀��,�0wg�9��p����&����G&�����^`� ��C��=}Bѱ�,s �%N�l%���$��vL��M�� ���b���X��o�
��f�Q�I���z�L�~��'��:��̬��9L�9ko�#^;�-���� �۔-�o�77:S��� ���?vj�3]`�2O�I������Q�L��� �g���K�ԽUrX�Wj�)�c���Y�j��~.�;�9+0V����U0��F�y�A���|H�I �� ���6e��\:d������W$�^j)�lfnD��̸�˜�.z��{I><v�8 ҉��ن�X$�(g�8f�r X��6��J�P�bͶ:�U��)����G����0N0��w��J�oP/����K�5�?���m�e)ȡ����GYlG�V��XԩD����ʈ�!qE�ZA=�mu����&��L������̥��N=�
T��8}�����ꏭ�����-����I7���	�E�y(�u��!�:��@��ʬV��tK�R����c7:Wڥ��w���l�!tؔl���X���(fS�+�Ӑ���`I�� Ԩ�3���u��}ϊK�sp�~oI��v����`y���_[0)�� e�����������ig�9�xo�� M��2�ј��H�0�D�%�[��5N�xN�`��7��~�dʈ�<�đ��R,X�5�k����&�/����܈�GChZP�S
v}K��s�����˘QDU��Y�b�_;�f�'��=�$'�#�ǃ|&��W`���D9ee�c?��d�;�nܹH^t͡�l$�O��-���3�AA������td3��^��n︇�Qn�aĤ�8'�!�����p��9�,�z\��xZ�=�,|-���V2C
���оᜦ��dV\Uà]���I�AӫD`�?t�Rע�0J+#��AW��G&}�'w�k����ЖJ$��%���DD�\�X*ʹ^��'�:p��A�Z�KL5��QX����c��a�A'7՝��V`0�����+����� Q]���::��* .(�IE�biV���f3�~�j
8R�?Y)����ti�^\�Pe|��Ҷ!���\�^rg5�gm#�]��`�1��N�&�r,�y��0q��7�7U�ܐ]�?w�x\`�-s��9'$w���"��}��Ṅ�A%Zی�0�g'�
��X��j5��W��x�t�$v'��Qnhޱb�%<��4��e��ζ��#�Z|�F���)�Ⱦ��vVyq@��s��ݵA��G`�+��X0hM��V�}�}wq �8N����o�$��P�O�Y�H`�c����Nv�P�H�����N�R�y8���C�|~UW``��v���"0ڶ��]�q��i9��i���1o �� ��u�_�#\b��._w4i�J��4%kK��Qg^�֐]����D����ƨ<d8�>|�$<����cPQ��k��,X��������T�� ��������(�	���RO�j{n0V�H�g�e���Q?Vy}��ߘ��C_�lR��E��5R�R=����(��5xܨ��˦S-bl�ԧ~�E�Q�Ww����nzN���V_\�
�r��\�X'���z�:�( t�~d6�DM~�T�POf��� �%���6��v��d9�;�3�6Q/BI��Ɓ��W����X@M�u�i5�o���L0fE۩D�_Ä%��w4�C�n�v8�:���#Ť���G�:St�B*�X�����DǓ*�+k���]�Y�8@�$�4�J ͥ����Mn��1P�{�����~{��&O//�����J���W1���/�HU��L�י�t��iz
MX% � �xE����]�h`�a��FW��?-U�|N��j+Ǉ݃ �AfXQ ,@��������[ln�"k�C����B�L���to!���9��^�ʝ���p>Z��@ld�ո��*WRq�$Yjl>9ó�dI�;�����;�2Ք��=k�)�]:�9���
���>�����A7'������)�i��UQ��n7[/*�q����J�tp���B3��K26տby����80;7d�p�/�M��}�+wqzg��U>�<�9Fs[I֑��c�uT���q�T@��-1u��U@UTX�2^�U7+m�L3�y�)ݧ6NQ��Daj��躑Œ�b�Ds��k>Y�ze ����)+�.����������A�����a�𼸽;�B�*q �K���8%Lx��f�L���`��|����u��0�N��L���ܿ������zc�����<�2�d|��h�%Q?=��`�J:T�����
��R�o�`ا�EWh�dƦN}��	G@%v:5� o覊8�c�lƍ�	P0"0ݲHݱG�ݞ3���uPX]�C4d�=�}�LMA�L���I�X��t�Ӣ�qyq�{4��+nQ#^��ۗ���01�VWȤ �bt��`ME�{�Ԗ߉��<��ǼT�1��Z*2�/y��=:�}�$���tw�(t�`�Q��'�A�SX�}��uʌ�Z7V�h�%zI�!��QV�c���ȒY����h��vA�Q�O/ ߹�&*��Bфgb���� Ǜ+/�w�A�.f}c����i	�(l>uuP����W�d�zƤ��yk@�Cnl�/�T.0a�����:X\�A������	��.jBPG�W5Viup��`Ԩ}k��̪��k0��2A�=7�'fS����{խ��?��Km�e���Gz¹���I��J�R�T�TIG�%%O���Jm���X,fM^I����%zA�Mm��c�� �@T����-��)���XS���K�˳��z` E65�74��Y�dU����J��{�������ҍ�-��3�]�dKi�Z��=;�d��A���~H���r��$!�t��DQ2�!��7����e�pR6]PJXT8��lLQq���̌����. �>du|�.�%:$(�!�C�Δ�)��l�b��I�,T�ӕ��S2��:֤�υ���DDG� kXu�H��fu�zw	������ Y:�:�'��vP���<������J���Uc_./ޱ�:B�~�F���C���{)���f��(��bn�ܹ�����ý�"K1`��E��p��&�UuP_є�!)��f 8z���$��V����LGN�C�Az5F�z�z*�E̚�4����$�:\�lb@{��0���@�g�����)�\�b`���=��X��;���˽��}BO��-�0�%��2
�7'�r�Lm��v�# �ؒ��̠g_�'�e�ܛH���W�g��:��6�������aM��i�6 TFZ�XƪR?l/dI�i������G�[Ӆ�d��A-҇}�����խ/�"�2�}���A�͕ 6�qlE���oJ[��|Xw�[34���4�:��X��H��cm�?g�F��t��+C��ɕ@[��N����X��W�©/��db����vȀ?w�ۊaj�{�����OV\��uc �� ��Z*��S��,�{�*+>Y��)"��/�	P��X���4���`��#ú�D��YX�J��elā�-����pD=�m���Y8�� ��0T�s��A"�Lٖa��	 ���=K����PV��] [�BD$c��6���W�u�n&�,&&ºMgК����T��Rq�٭��~?��Ĥ�$̍���EϞ�:90Ҥ�e�Y��u���Iw�/�4�Vtj[�{����.\�,`@�#龻F7� �]Q߈E���RU3��(ZRl��F/�+���Ґ��W�jd��MP%p������p��p-US� �9x~�1�m���PAĊ'���(�=�Y)eq]2N ��	v �e��n5�#����$��$�1�J�X��F!�B	 e&����*�������5q�z�ሀ5x�!����t���_DՙVM�`�ES�mi��1��x�:U�cuw��X �>�%�S4|�� ����D�Jϐ�a�`�M��'Zu�c`T1�c󃻜L�{�������c�Z�B2�����'r�V���t=��"��
@���Fm//��O��&z:߀�d��lL��-����l���(PA�������S�}!�w����l��j7+�|L��#��(�SQ�=D~���8*3X��Š8ͶC�dz+Vpg�퓊��C�H_�|�@�΍D��\����X�R�n�G�8ۈ`���T431��]�"D͢�C�N~�u@b��:s&�1�ؾ�ќY�4�H�%F.�:	�'��@`Á��`��h+� �(��hYL|V_��
�~}^$��?�{�� �����oLO~���v
���P�_���wPo��zw�7v���M'0	�"�;TY-�����,�<iJH4�8..��|�V��t>�汸�*�n�R�B�KrۄD@(�j	l�"$k�L��óH�Т��T_n���S�3��d�@U��e0���3e��avfw��w=)��<�`� ��Mt�� 08�P@��`@Sp�`9
��@����l�R�A���P?F�\��+Wu�	�`��%�,�O�D�p䗊rp�A�eL<�2���@F@?�26��d�io��j���$��&؇�N�
|Ⱥ����QR���
 �)��S����;>��B���-b���Y<@F�Xu�zIdZ+I&f�H��Aԟ9�.Q��)�$����t5�'�F��;�O}v L���Fb�cɑ�B��d»��Xj���P�{3VZ��ox�~r�~�Z�/Y�t.a)Jy���`GN���cD��ˠ���͍��SGﴓ��Pr��Da;Ӎ�c}6���
�������r�tM*"ډyJ�*��K��~�
�b�ss�˔D/#�e�|4���>7��(�zU�A���� 
JZG�W���-Y&g�V �j�%\t��H )��ϋ����Jw�YL�^�0�����d:V�����n;����DB@I�;<bF�D�9Eܦ��l# �wʼ�J7�%�J��f�:��)}���[�<g�"׸`��5u�$X՗u��xŀ���% �&BZ� E ��T?IЫ����7-ߑ���������&�����n�����6H'����E��`���0.:����������0�}������A��-����bp��"��� �ҭxݜ�$vw�B�b�����D��M�f�;ҽ�9h��Fk7Ĭ/����K���|�1��1��%	��;*3*oQU]�	M�ӄ���hR��ѽ,M��5�{��a����u���K��ɑ\��y�O1���ܛ��PwXt#k�j݇�j�j&�2=�)�%"��jHOp]q�HV���t���>��˧���{���	,�b�!TŁgMҝD v�~��|�R����4>17��#G�~'@-�nQ`z��c.}̎�����6،��(8�� 4Y��흊nce�Ȇ�k"��i�-�٘/�f�.�%���-�.2t���	�݃���Z����t�U���3��p�uΖ���t�"�o���IPp�2�W�,��ى�4{�#TқT���*e�Z���Bi�=Sa��à>��S	�T�gD��)?��]���4!��9ݐޝ��C�1ۤ+IvR�ܾ�5Z�ɜ��\T�ߨ�J�e����U�'Vg�!��N��:�ߦ[c�t/>ާ��w��΃P�)�~��s-�&v�NH#y-^A?j�W��+Bt�T}������N}@̌�49�V��6O�^��f�l����YwV�H	1?�a·���)��F�,�����K�=l6˻���	���{'S�K�#�suy��$�_����6�I�򜲉���)TW�Th*fhto+t�������d9�zmL����:[������5�`{{�
�yD�{�RD<�H��˜�?�y>�܀�����_&0�¾��6z���M.%�O)�,� 5E��S�^�����A�Bo��쫨���%{@���@3�3��{�\��?}���%���O!	K�4P��Q�%	�.}W��%��X,�Mk}��˫jyl[`��>M�K��f�5�UAe7=|X<	L?�@�[�'!#t^��72` ���f/b.��v�řKR]�-��|f�kO�u��
N�2̂4``T�d��_��E�c����<��O���|﷢���A�>��ED����u!96R���j�3�7�W�8�:%؂�o��W���T��MY��{�%>�[��%`c�(6vgz��s&W*�R�a�"}�n���  ���	�=S�aU:I*�'P�ܥ�|��D�M�/?�i-�(��h�7]�/�tщ��	��n���d�OWWW���;��������1�C%d^ꂅ�h��PV7X����?��h,��U���YWbl5����苓e�Ec�\�^F,��$����]E�0ѝ�!À��� ����U!Y9#�w�;����V�L�8 ꢌ��h�Fź8��!o�e�/���tkC�	�7��Y�h�\]yj�K(W��ݻk�1�A�j
M� B#�樖澟긕��R�idU�͏�幰e��c欹� Rt�w{�s)�T�jA�oʢ����!���"��Y_��՘Wd0֕�ޛO(:�?�ްh���F��s�s�3�x�ߘ��DX:KXh�Ɂ	��e��u!�	Шm�y>��s��OO�}���[��K�8��f�>�$���n�G�T���G��S0�]9  8�S��ջ�,�� �P�_�i�L�ڇN}�s�1!���L�.�hˁ�IV!E��+5P�y�&=1�ۙ��b��Q��]B��"u\�����;��i"Xl7�`D�z����_��F�,1�+uwb�%��~��j jݫ�%��s�ԉ)1{�Xt����v�	f�{�����qT6L�A�WW���*�M��o��*�29���Z�{5(���~��*>ݖ��n�cƨ�,�_��q2(���D��+�Zn���R\�h��Ơ�	��F����&��ǟ|<;ū��������]��E����������'6J!l�:��
��'DQ��lE_NR��/����X�i�E��	�`��$-M��p��$�h�>�و����Fa���|�����1IMt��3�0�{z�U�/���!�g�۝�X��ؽJr�{�o��W�*_�ڸ6Ɗ	���M��D丠�Cm?1��-b�"�Z?g�^mk���ŵw3% ��*hRq���r*��;%B��<��uF�ل��4m� ����!Ys�E�f�-���o������{�_��#�a,֖#^�������W	���2�V�K���MfF�rP$���;�P������Fگg�:7n��]:�75)�I���S.g��j�g�|����% 5�� �ٻ��S�ygɐ(�樽�։�y�ό�>��?�g��b��/���>O��X)D}�\��o�^%��ͧsnU�b�ʔ}�gz�������L�B��K��8R�����8���ACW�86Ց���������\B�j���$(���A�]�`�W���V���؝�a0~��^)���;�uauUӳ.�_e���Y���-����e�a�� X���Rt��?$�E,��NU�wVZ�誸
�D�h�~��:r������@��ff���#�$�~�z4��x��R��g],tT�gm�
_>��_$w�.ʩ�������;.��+�ƅ2�}H��.Y]�Kc�(MƟG���oI�������!~��ݠ�M�P�,e�d+4X��|hl��'�"Y�0ܝ<� 	�������dH����D�������٦D_Nm��7�jh���BWt���2 U���NP1�Ө*�=�>��&b�f*��x��]� �w�w���܃��MmMR
Y��
R���ܪ�w���w�z�'O����B�lT�a�rޢ��HO[),y���x�jp��]k�.�&ˋj�ϰQĿ���n��c�4 �^C=�ɳݛ��tk�Q��V]��U��7�)1PIr3�6�@:Y����d�%��#r�M��P��)S2�l5���'[��N��T"q� �D�AAO�	Fv�N��".�d�� s̫Qr�)d�\nؗ��:T��,�	����3ǜg�O���:J��I��3�3J��U�Z)����(*��NnH�/
ҁ�{�=�K7�_����������'�	�(S�A��e2ݚ[���M�% #���2��U��QjR׃��ˌ�c�E�!�ԽK�&0%'}z�u�8���z�ޒ~w�����,�c  /�C(2�Q��{�n:��Lз�"�h=�_�_Ӌg�4��3��5[��今��q�Q���*:�����e�v�jd��������%������+�2��4PF���;h���^�FD�ܫ���z�^@��ڙ)����˗"�,�3Q�
��1i��U���ģ�-���AL��2��v��S���U�Ttu���ԉ�߅�
�I#���Y�{Sd�N̆���
D iY�\T�\��xœ�����E���������W�c���i�8�m������)��FA��)�D�����&'cz�mQ�sv_Y�a�4���/6�G��t�>~J_���������4�X�d�^!}�IX�
��/%3ը�|P7:���m'�/�J�4��rY���>�l�<�q.������bS������*�臚>�oϙm '㛇�3G�t�f(b��h�ׄ(�+�Gǐ�D>�IЫލ�'&CL�~���8HV"2!	�_��fы"��P��\���>�e�U_Ń��u�<�ۡ����D@���Y�'�&x+�M����B#h�������V���ʢ�vҮ;h�eo,�CV��O�7]:L�S�A�Q�"LU���Z��� �~��=�ʴ�C���-\�ڂ,����?��Dz��ӳ�B z��l��P!�$�1�;���D�/"����{5�D����B;�3�(d�4H;��&p'6�˧_������?uB�i�>TE� l8٤ϓ�A<UHj���;1�>��\D��yc5,6z����������d<4PU{��ިu���G��Io����2Ҹ�Б�F��5\ܛCs{*`"�V�®�x��9ZDf_X�hPYRh�}�XJ�14�����d��4�9���>}���]���4�T|��˨���{[�^�9�ʕq�ǽZtK�)�ؖ&�N<�H$�	����d�[q��������A\fh�^YQ�:� s���ɢ3�U�������N�>�e0�_���d�H0���
چC�b�ih0M<������I��c�@Y"��QRn5i���~���xn;������ƈ$'��0�':��%��/��p����G��\�������3%�J�:����I���*]7��D�'�&��'ѭ2�>��QU��0��������QX�C�L�pQ�F ����"8:}�����ޛ��m$I� 2��M����ε�ξ������RK)�ue&s7�dդ�R���J��@Dx�����U?�~1w�+��14LCe=&s�Ci8'C�.�"4�ԩ���pO>�D������B@x!w��5�	�f���k�z�j�mGo�+�£I1�j�����R~���45)f��czƖ,C�z�׫�vܱ�Em	��Ò�1	 R�(��2��К�:����P=�c�	�����Q^X��'z���X��3%
Q�3�_�}��x�m0k�#ن#���
x��캨�/�37�h7�*�b�$h���%E���CՇ�<��4�6�mU`��{��5����Źk9����=�Z��P�)����b~b�s��y���.�?K���f�5daJ�(ZU�g/���Μ�`�S)}v�'NJ�k.�:��gx�ue->�C-a��$�d�	(��0��z>�.�W>�̴��M���z�6>c�ׂp�8�.x{�x(�;�V�y��lrm��S7�Z�e+�N!��TjQ��ޑ�<wk��E�1���9�5r��p�B��v��z&X�Yt�`�!M=�ߔ����J5���0��h�mn2�8�l,Ww؏sm�W=EL���D�$g�����F�Ң�g?���>}:{�o���@g�p��lH�ObSR"&]������**�0�d��2���\�ʒCAT7Z���G?��n��E����5��K�,� ��M.��� ���,�?=}����콙���Y�T��a�u�8LZ	M�?s~�'��ĄJ1�3�󴧟���!7�����S;&60&�$�����S&�0���i��;�[;g��s/@r`^`��~FU��9�G(�cK���hG����	W�h�])�j˒H��B8�cT�,��>��3�G��Nc��`�|&�������ݍ.plXJ'[+��qmj�y�8��u�J���7o�ۻJ��A�������4�<2�O+%1:q�aG����L/=cO����~xf�)��'�eW �W
�zL1g)r����Z	w�{,�^��&��STIR�)�v�/]X�IF����u`�7jU\m/eQ�:[�k�9��}ǌ:�ʁ���V��xޏ�\�|��v�B�a�&��'Ǵ@�n�(��_٠:z�s���;�z2�E"*�p@�t^T+N���fˊ���:��|T9��o֌�l���ZU3�� ל�d��e�n;N�c��w�3��v++
 �:`G.Z��I�JL�!	6/`�'��kڱ���V�k1��F��t���������o�T��A�".�aR[�^�Xc8L���C�p)������]1��X�WՏ�8dt�����0$H�a�y��y���熛�9४q�&t ���k�GG�<����Ј����`���t�#y��|�G��J3��G@�c�'���T��2aA.;&U���gaޕ���\k>o�Ã��1šb�<:E�HG��ð�M��{���8T�@mf���?蟧��ǯgPe�~.���Hub��}��Co!���P ��P'�i��s)�����ߧ��L"�p����	���&��pI!��h���S^G�Ϊ���y�:��.��/�D�#|��v�+��S`��~����NՒla�^����<����//�"�ґy0�s�VS$�\���_;��&�g^�W0s�ѻP�

�3���_J�ն�.bx�vo<�8�d��||��4�:9���#F+B,��V�����2�<�Pѿ:Q���vo0g��v�y<�э5L����S�˰�VJ<��65j�n�*C�j5��9��Lg~��16����>Z�:8!SI$5�H�r��>K�������6�
�m���R���vj��	����Ԩ����������]��'�S�5�^�L��o1�'˥vcL)����ud��X���tޱQ2h;���v�ׯ^�gO�R��O���w��Ҍ!�ф�ď�;�=��0N�*[��ZX;%��O����R2��2�0䧧vM�=�Y��[�ؼ���}�~��>��|}n�i۪�J���l6��20e$xd� p>ƷǤ�*�(����sf���Qy�vdab����8a�R̈́�W��K���Rqo�g����{�4�[vBPb&tL/=�?e���g����{�em�Jx�ɜ��L�);eޕ��۰?�s�q��U|(�!OR��.T>���@m��&�`���j�T�� z����$��0D0�mc�R�!*�P�myS�t� �ٛ�>�����Ym��{�+���CJq/
�-ֻi$�b�ɸ�s�0N���NT".�>���Te��E��X�.b���=��ކ{<9<(	Z�g��*	;�Dv�͡W�L}N�\��0P+�c����+3��Ӈ��D�6�3�����M�!D��
2��.�U�ڢd�G<X��/�|�y���l���q�J�NI��|n��7z���������l�ۨ��`��.�K�u�E9)�]b��Ҕr�k1E���B�E\��r���Tjŏh;vdsvn8)6O�_�|i�5>�|����&���Q�*T؀�s���D1Ñ�By��ݠ�@�%���&e�yS��JZ0V�	
���j�h���.�o��������2i�������(�e��
wl�{�9��=�����<l�U����J�JY�!.1J�o�'��֦��p��Q}F��/Q)U�M0|���G���C�&��N��u��;����W���c��K�?i����;���'O���O���p24��o�æ��n�va<M�i�j8��S�B%�0pKer��K�ǂt���l��ؒ��-�J
GSBF��۷o�W��X���Ƶ%�!��z�JzL���2-X���H�x0E+aeN����J�a�ȣ3���雦�z�B4Y7�	������w�x�}r̔�C����eڠ�26������_�+���[���t�a�Dx���1q�J��,V|Q��!xIQQ�"O���@1��s���7�p����`����n�Q��,�n��\%N�~S�m_,�w~�V%`���O&<�6p�e'n��Y�Z�,��g��K���a��2k��wP�C����0�N�1J�4�DŢz=O:xf�Xp+#E�x,�5�f��9�F%
��o~�[��0�/��(�~0�����fg��+9ԫt3����j���"��̽���5q�]k��������zE�A���H��u�d2����]�����Ci�qt��������ϟ�b��a\����h��.��B�.]gN���G��K�Qa�L�N�U�I4����"�MY�@l�*�����%/�����_q�^B瘡W�mChw#+�rW�+��k(f��F
���Q��k�k�[�We�2l��S����d�o�b�r:������zmu��B�M��[$\�)�wGά8����[��OG��F[�͖p�+�IȈ����m������;n���>��c�m&!j�?��lp���A�D���&��%h�I�U$glB�U4x/�M@z ����ij?���{Ǯ�Ϸ;�,����G]@����6B��jM����G%,n1[��yG�O�Jÿ�O���)�0bZ��)x���і��SP������*o� ��؟���F�ڄ�1fK{��j�E{K���s�&���CaT������e��I��<6��[�8�mӳRb������:�M��Y�(P:O^�ѧ��C�iK�2�g~�%�/��!�pKwR8n}��h+���*FN��}f��y��?81<���h+�*>H8bnS-JE.��W8l$����qlJ�;�ލ���HZ2!z�J���d�1{�8��l����3�~�F�=~�,��%�~��خ��A5o�+���;��ޟ��f]�~�+������M��� ��������`4�!��QEk��1{6��"=����X;ULLnmY��C5�E����x�q�T
�l�55����]��J-jX�%	�K���#��"�x	�*�0��p㛰@�xC����\y�kM{Svjc=qq�g�`�?u�%��p%�Xت�""�"��wPd�}��w�{=[y�v�ÁGA�T��"�w4D0�+������w��і�y��o*8��=u��f�{.XC�h��'g0O-ܺ��-sN(I�j-L��N!�#<��!�ҷ�s7�}�7��ȿ:�A�Ӿ�3`m��4P	����$�k�޺ ����u3z՘��B	R̘�ߘ��EC~�s$G��g}��|S]P�XK����" �*�c��~�2ե� S��BL:x8�p���l�Q=�b6:���J��_�F�� g1�1V��%��</hK������<<�c�l11<_nH�IS%m�#췶+��>��{`��c!Y�*��Rk�3:x���y�'po؏������~g�fC\p�f_�d��Mr���.S?�h�
*a^���7e>�RN�B���X-��HoA�b1S��� c���ᓧL,}ʴfq?S�5qH�L��.=3�?�=��)���0 �ss����4h'�$��tol~��|����5�lS�獹k��yW���lH،޺�����l�����6y�ư��_��QJQ1���5������wy���ۑ_��eզ���߳��VȢ�hGl�S��{���f��K��F8���-F�p-*q�.�I}��<={�<}������{��/�L_~��e�Qr�J�2��<�`�S��״e���Zi[�`"<�H��x���:�J|Ԡ��Ʉ��LkNb�޿��b�=U�#'z����P�0{FJHذ��P�Ht�ʛ���'+���C��-��D��:����H�\F��lP��69v*�[u��!����X�H�7�_�`a�N�3kt*uM��U%L
g.�Q�!�8�:*��68.I��B��}w��Dr�Z���]�L�M߹u۸�[��Ċ?�Uw�v�9��s�9gs���d�@=�MUu'Q�a�@�MPR)�el���W�I�6)��2ԟ���j�3Y��3ӽN��-����g�����8g5y����Ώ�Lo^�v���T���C<�UKL��L�ڥ���|T��#��7�̆�^���~�5Р �?8!��S�Y8�Ņ�Ǹ�*����N]�P�3d�ǘQꐚc!�Ÿu}TSŚ��x�%f�w]`zx�%t1غ�Y����$����T�f�A�gIe�S���b~�<�~�,�#��%���Z�%�.���a$,ԦAp�whڄ8��C��rƲK@9#U���_�Oφi��'f��VE쓑����l��(CJ��Z�����9J�'�����Hs��,�A/+����w�]��/�79�N$l�M`M<�2$:6�˄n��g9;��\���75=��E#Մ�p��}h���1m���/����e���<�ﹰ3WEgN�mM��*����
��}/����[ń3��L�g4�a�-CV������]z���׶�pHn`�M"m��-�Co�zXm.���zZ��RqQMNI�@U?��"���F]w����<��C^�x��熐�Ȟ?>;N!�溼�N�Z�F���:V�Wn��<�iZ&��yP�藶2��.aOS
�⒝M�:�+}�+�g*�K���q3 oTmRDi��w,m�dXl�U��d�oʖ�)m	���w-��+kõrYW��"Px��f�^k��^og�w%HLob`9�m0j@y��뺦h���Oo���G�4���@�6�yc���
;w`��A��~��)�L�p�{�r�C���bx��6���
����j�GrA�#�'�ُ��U�B��d��sR�,	�����ca�`�.�aZ���7������E?��	a�d���t�e�~�16�Ǥ�K���/���-Po��T��x�v��Tl&�x��<~��޻g���a�ċ�XT�>,,���q//"���l�6�mL+�܍.�b�5�k=߫2�bQ��qSs���dֿ��ͨ7/�LK��q3H̐!�S<wHn��&j�4?$�c�~6,&[�3�
,��Cc:ۘ؏L�zҋ���a��4V#�E[x.k����16VQ'�~��si�I���j%����^��)a��i�{�f?��mO�{��L#z�j�[;c��F\Z�H�|�t�P��}���GJ�-�������3�5����n�����)��#`���dȌ	��M��$�]aAa'�2�b-�)��b��F\Na��ә'��8�x�lJ*���׾�*^G�Ս���d��)�J�FVJ�ŴS����ՄJ��Uo�U�/��=|�0}��ז8�P������p��O$��͆�hV|���I���e�+Fdk���
�_W�;?ӕ����ޣ��3-�Bz�08 ���ݺp�⽉����5��`�|d�������y���cNV7����o��8�}/��F���6)�A��BXH�>�<f�;�"�G��E0��Nߦs��e�hs���茆��,7������K�׳�X��В�ڰ��Δ$��Mq�~ʫZ�
��yQӿ?3q�g��~2��ɽH���յ#~z�=��0�²F�v� �����a�{�u���z�����I���H(�a)v�1��q�U�"m��~�!a�Dӥ����'���P�U�֬���	�ɫd��%�jEj�	�I�aP�8,��Ϻ����1<���khi�W����{@��̴�-L�d`	�F~c�w������}Ć��m�A��&��w��ϖ����K�{kT�ɛ��Glc��rs�0j�l<70�'�4Z� {zv���UA<%��F)�n��s�}�6&V �G�_�(��	��>#"0hf���86]�Y�?��rp�X%�kz�S��mx���Z�9.�a0�`�vPՅu��0�J_�ݧ�'&��Ffd�����}+,Fə��EV���s�a��K� lKZ:T5��|�O��ĠT&gGIQ�q*ȄOR��	|���&��<Ŝcbc�X�������nG7��9�>���?|�����H�{��f#��nY`dPSr�=lÚ�O�d�]k��Z���֚��ܽL��'�kQ~G��*�y8�_|a���B�?�sN,�6�5���.'n����;rG��)-��ŋ��ts�U!/�����^� `s���>H�MԜ�[;��QqS�@�Z����I�}L��v�Ț(�?:,�ș��%�E<���8�H�޼��r|cq}�ǄQ5��X۱�6��	Ɓ\Ri,�g�3#;FTP&����3�8��ͥ�F�H�lܑ����"�  ��H��~���ڌі�aщ���_�6S8#��bI��܇θ�x<���̛����;4F��KQ�UH�Q��6��a���EK�ԹQ�|P��Im^*D����|�	��n�[�]��L��Pw���<Y=��o��I<+�6�y�0�B���~��O�R���5��Z@;V�H�B�A�Ob�k�u�wo�y�0��b4�S�Dq��O�����We��8�^&R�s�DE�~��v�������F�F�9p^oq}a�<�DU�h��ydJE�� ��<Je�����������Ed�܌�������7L|J�}�I�mYW߳�'V�i���o��席m�U�)���,�]�q�M�;5�fS��׊�l������ʒ�^�aF#���[�vq�2��S&5I����Шs�M$b}�����>l��0��Z�,�LF��T�C`�a���٣=<0��`{������
!c^j��:��������&i>�qc��.�p��k�1yAʾv����h�!�Đ�Blǫ ;�5�I�%k������Z��0ʃ�����4*e��3���c=��D��%�D���r�'�eq��_A�PI-��r��R�\I��w+�fB�����db���L�I��r��f�>K|����%�Mj��Ϣ�	W�Ϗ��
��6ucݸ�[�����{�s�u�)�h�6�e2���S�H�HUg���DbIjRf4���c�0��8���� Ff�֫-j*6�s� ��n����ίt-���ZK���������u���!��`��6�f�/���<�� u��㨆�l�X���r���Ζ�+1�vM�SMTL�D=T%�ںcSB�|i���	"�ף�(��}��S�,�j�]Pث��F[sAS"��*{ڷ��ݴK�%��A���P,��p�R�t��;��2Z�h�->�35�n����o"|vA�:�G|��l����۸���fDL\(V�h4��I%�?���x�F���M����4d�;� �m��S�d��c����"G��d+W(Ai�27Ei���)�"kja�K��$(E׳kTeXI����;%�C�G�r�<P׿E��;��f.�Rg&x��
e1V����j}�Ɋ��|���Q1͎��~���_�9��N6�4�";��%���}���cgo�aLi�B��TOHX����S�	 �IjW�%	v��\pD������<7unդ�k-�k�e��'�E[�s���w�u��<`�HV�/������&pO�;N{Nɶ����V�'��^��?cM�I�l7��#�>�1��Nwb��[~��]�*�9���P�j�v�~[�������rx&Q�h�� �G�N���M�f�䖚;��	!���JY2�"�.�Ehp/P��b�ok 	����j��\�!�h��'�Ql�k�DC��jC��ŕ'���f�cP�W��c��p�.o��G��4��S�D�O^w�0��:f2����2�b"�}�I���.���6��:E�nx��}�Ml�����%"d�,�ua���Zz?�]x�,Aab+i{��X%^'z%��Z�v�`���ޟ�Y�!�Si�7[2cM0��p�"�o�ݭ��ǎ:S�r��s<�ݑ��"A"�Q����H�Dэډ8��O�ef&-lߍ�)g��I��1�x��تr�5�^ƕ6����x9p}�S)R�_F���߹z�b�`��\�*��J.���b΄O�1&�2	x����U\ۮ�M9l
�ﳤkߐ��ʏcPü4�T���	�[�ͷm��R����˙Y��3�j�`I��6��H���R�	V�(k�R�OSP���%.X��~�W��$���<�.f@�3�ro��ӥ�z���)3�{�N��f�0ɮ�cul�0[�����Z���^���k�̍��G�Fڢ�Hwcl�J~�\"�l%�F�ro��$�'�ؕt 6jb߽{���hW�{}���\��<U7�l���q�JM�d��L6�(����I�Y�ɦ��=5.\��+�V�^�����#)_��0̓W�f�ڐ���<�}X�nvU_A2�ߎ=�A��/q'/���!:�gK\5<��ʚ]���������	Ob"�1݄�o�gZrfU�P���M)�s�����4��w�)c$�ρy֢d`�vs��k�@!�Fb��pp1���ޫ���46�5�F�H�G'�{����)�{��#�Ɣ���LT<����f6��*�T���i�G#�p}0�ɍM�m7���ףO6��懇��/�W�m������R�Ri�Ί��9���a��I�vԝԻ�N�m#�x|�Rs��ʾ����YE�FV b~u5�Rm�=5�K\?�M7Ơ��)B��rR��
��[9��-U6ܤ׼T0j�ɛu([�6�IY��YO��/*OrO��ş�Bγ�c�O?]WE�,Y����Y���g���ΎBQ�iT��%��l�Zcb�&��p��%3���3r�wKZ��-ZDm�KP�*�QG�Gq���ӊ�js��x?0����;��'�F�unB'!U/k���vY�F��N񙰼S.��!L�Sl�F���l��rT�9A7�
�-�t��A�q+zc����Ax�8L g�^1>z
W�·�3�|ΎM�j��/�}�<�ԼD��M����fԼ�=p{VulU�pdG�<���ءOԣG�͓� RT���SR��Q����%&V�W��7Q+V":��ZS4����w�g�%��Y�Y}�̨;vO�*��$	a !�"������5,�w�qAn*�-���<FҥMX�9I֭� �"V�5O��%L���)��Ż�2�D��B$I;ϩ5Ƃt��O��
]�L .�
ɯn�U$'\y��x�tFYb�9"��uY�7b�v>�TE�G�F��yOET$!�h�^P��:������4���Xsp�rhGU�QI�ﶵ�L�����7à��$��B��0)��R`xKz��Sp���ɓ'f�`T0y\l�r�,�ML�)�dKD�ת�N	&�YK�4B�i
��p);�NI�LE�e^��9f�:~;�Ϫx6�������X�W�/�x�Q����V[n��U��3������rv)��J�E�Y3���d���6�E������~S���|zQ�y�;�S�!�ƶ^K}�{�{�,IF�&����u.�{�k�><)垟�z�~��V^f�>�)�.��ldQ�4�h?�_���_�S=d{�i�Q��sa�lr�`�n�k�X�*�]�R5�W��o�1U��nL�7�nZ���>�.���9%�uO�|bޝ)P�����Fm��H��hb�/��S�#�,�uAmqJM|��+�&�+��4U��Z��j�ro�O����g@!j��U��*�q�y�6�z�*�0����C�r�b�Z�g���I�W���3�v��R$��(��+Z��
��!�]���3�yoAj��k�P�JYxN�D����B=�&{���$�Kɮ���7�f}Jx����{7F��0���^24�m���9gZr�u��CJQi�Z�8U�b~��%c|kF0~��d6��X�sp(���cjf܅TV��0�p&��]w�
�PǸ�y���4������7��"h{q;q}��h'�Z� �?UAw�g?�e��^��s�%�;<������~&�+�{�q�M�������|Wx���^��bx�f
!��Y�08®�8�����l�'fS3�����	�RR͙����t�J*.D|�Ĉq �����5y��AQm�U���ĠSu�8��|q�cx@UC��Pc*�:���E�Ŭ���"w5M%�kz�<��|?��t�y��0�����7�f�����~{ZOa��P�H ��DsQT�L���h�����E��w9^{tvj��Y��������9�Z0�n�J8j�S�U_�]U��iLn��z��
��`�Eqvސ�m�W��U8����w�,�F��s�p.�b��6���GȀg>��Ԡ.���%�,[�t�+z��T<^�,I(�\��RX9�TmT��7�H�7=��G�P]�'��mR~4��q����v̹�L�HFq�$\ʒr���^�j�ɫ��W'�{��*|2����c�s>��6<���ɼ��Q'nڭv������Pog/�;�:.6�^�����6�E���2ڭx����7�_d��X�M6�<�����po��^�ҳ$s���ĈBި�+��7I������-[�%\f��觋p7`2�I��;�i��1NΦ�S���;��ݻ��j��?eg�E�':�0�{���ꈡVʗWw���:�/�$�D��#[�[���+�:��d�SYI�$�^�:hpb0ޗ�KpZ�-�&��m��Q�_|�=��/{Je�E��a����I��qcB��h�I;a�I�)�r�y�QUwl�J�B�y"�J�YA"$hQ��:�k�V[����Jδ�>�ݫ``V����c�B��D�q>֫�|>�n��uC��X�A��h��0Rx��P��>��;=�����7����sz��T^g���FŐ�,�-���>Ή!{�\�kܑ��]�A8�yŽ6�:O*��7ޚ��w�����a�� �FC��`�M��ʤ5�p���ߔ�:K���G~�e*��v��OE.��v,�M�W�aSI��k�`�\ֲJ��������ϊ=<:��>Q�*�B(������q3jb�Xj|R�����~,6�L� j�'�ư-�CY��LБ��2�l��5�5�)��O�]��'ɪ���?��\He�@JQ��o�,jw�-�����PKS�g�����}h6�n0���5�r<�J��vM
s镻�L5�rSj��������$d��2����\{BE)U����)�S%l`���׍�=B�h��驧��8��\���M/�����
N(SB1��:O@�x9Rɣ����vB`�)UQ��GO�~�����ѓ�셅<*�"W��!�����ۄ����n����hPe�����T�9-��$��Yh�I���_���ƵA�
�w�d0k���
[�bf얆Am	0��X�d�;z$��Ґz�0������wCyq���]`�B/���N�E���!Yq��40��y\���K�w�^�}�v�ꫯ"+�dS��T�`[�ɚoV[��2q��#���*��K���+GH�U���ͬo@U޲Ċ�]V��gR(q�r�,��w� �l9E�ט]�$�/7!0I:��5�Kżҗ/_Q��|!�g��Rz�}OvO�)Z�ob���g�R�������O(�sa�%�U�(_3��V/՝��m?*\��u��ٟ��Ų|<W�zc�aPn�@����i5ySR�jCĠ�L���Ճ�(J
�_�Ʈ��E!�H�6Iw��D�4[{����;I��D�̙-̵��q 78�	o�[OoM�c�'�i��H�����m�e��q�������8u�4+|BO)q)] �lǊ0kA<5UU̜�PØ���N0J���8zQK�p�����������8�2�\�J�HsD�x*u>��xa������~�"�4�9QЄ���}b������<���ׯ�����|``�V�<ЋoA}Я�s�Q��WlC��G~���#�ټ|��	 �G��ΰC?�=�V/���RƱ6��	��L�ub�U��~̸S�Q�)+w��o�8�3?n�Am��r#@�$������~� ��nnI�T��R���r�EYL�S�5��kz[�񬚄��G�s��q�|'���<�ub��/�=x���w[Fxjq5�������읜6�i�x޲���hV�&��V��*��r��"��m�W�U���
���m��Z�sq�e�ɬp�"�]G��lbyd��0�/��Z᯷�� �nB�[g�L�Y���Eo�Du��b>v���nb2�5&�#<5�N�?���g��s �-^�B}%�px���<b�l1��xC���}i�jT���W���j�#��1M�o����^>!>�F
�-m��M7�7Ƞr3�V�!�Dɂb!��aOE��\S
�P�ca���S��j�N�K�x�]#k�E�H$廇:S$���o�CE�N�~����$�U�(���z89	�!��q��4���+]ڽC�q6�[{�a�IMwd.lB����DR���'����D�]Y�w��3-�U-�m=G��楕 m>��	GkсpÚ�����&�=8�
�£�.��"\?�`0�� ��tR�~��Vx��
��q7��6�j�v�	��4�{:��(C}���o��b�Te��_�b�}7�F�{��������A���j�R�7��"�\D�K�qmJ �)ǘ$y�Y^OM�?�O���{� �Z�{�2�="a�k־��RC�-ED*�^I @��"�;��%x��"4��I�a�Q��t��4�\_�y��6�.�P��l����:�j0��5�õo'_4=S��E"�ײ�)1,ł���bl���a��R�ZO��*�RZJ�U��j����z_{�ٟ9d�jS9]�gm�/��~V}�FUa�̂�X��^%����h:��w�@�)��J~��w��4ajl�Ö��CR�~�Y����0�H"���{�"�)�w+]pBO-[��rj���/����\���䰎�:L$,]Ձm��
�w�k-7j�DqH��8��(�O>�?��~�Ǎ2�80	q�~\���x&�<׉�f���s��@l^g��y��Ք���e�)6W�4g#���'��O���2�-)�BJ*�!=7�����R�solV���P+�80���̸�vQ�o���7�� ;
p[ჩ�'&��<��ǆ��*�d$�`���ˆ]*�q�?�hi�}^Y�m/'Oԥ˺@ͫ������C�cf�!��{;�SƩJ�YT�
�R-UV�c)W�)B�\|�V�� ������"c���d�t\����^Q�ˍ�������N��L |��̉yx�JG�Am�G���+���;c/���d�Gl�P5��<Ø��g�7��Q����
�����ɍ�<��ۓZ5�-k���S�#���Z{�gۍK���`[y���̝�����Oz���Ԋ$Ƿ )'_`�āY_U�H��ϑu�&V2�U��W�^�&�70,���J�첉{b^:��ݰ�$�,/k�6�T�R�lO�����q���T38?N�'.8���Ԃ/r^�*]��`��6�BC�+<�k����z�Zo��1_��M��t��/
��Zvo��9W.������U�GPFDPr+s^�TOI^�n��#�`���X4��ꌋ����
W�f����������v�Ҟhܩ�n���b�Dz"�{��hj>����Ơ�$�k�;�����E�P��2�6�����4-�bM�NڥZ���)wH��HUkm��G���!�싁��?e�jng���^�6���8�g�g�}��r��0�Xd/^����B�l�7�9��s�}�����J7�����'�V$/<B�qe2v'FV��ȧ��<�����o�y�ni��?e�U� ҄�#biH��=te���ý��7N��3�>��c:���E1[���j��	��V.���yY�ʀ-�����x@�����y_���޽���7�C���G����9׆�T�[�dZ�$�����@���~b![9�"�+!�뷪�Ġ�6դ���Ę��p�NXxL�s0&%����>{o=�1��jo�������&�g(�c��J��l��� ޳�*�,�C&8J�h�ڍ]�*J�+o�b������������������*] ʘ��a6�yEA��qBx��ਧ;��сe�ONnY�6��0�K���	>��$XmSX.�{�̮�j¹U�Vм����:��5�E�J3���M{�N���l:6�N�iCԐ�lڵ�����%E������}Ud���Ko9��*�x;��;|���m�.�ZG
�v˚�)�Q�R�o��쪫�	���%���yH~���Qlw��V��v�^�6o��Ƞ5��R�sS҄���u��eA},~_u�x�ԁ�&WuS���A.����߇�u�ׂ��ίt|2��������@h�k�%��pG*�S�_���z4"�'!d�7�t��N���+[�3�;�����V�|�>v�}���kv�84,3ۤ<e�{�.#��zY.]O�������ac�g�!��u�ȕ���#���EB=�\R�����9|��m f�֨�>���������?�;�路o������[\kj[b��u��݆2��lx�p}�$�jӌ�Q��\q��I����G��4�!1�VK�r�{"��s��m�i�t��ـ�̞����u��ᣵ����vaK�~�Ѕ""����4�yd[޳�O��MK�i��'Y�<�=U����� Vu)$Eמ$J^m�1���v[��&X� ����Yb�aB�\��,$,M��6�m��w����6�(�x��v޲pV��Ȅ�i��m�\\���:�)���'އp-��1�Lh
}N�'5��/�z,�T���z�\�q��*�{���nU�M�c�v�x���A��]��8(K�v����M:mW�I�X�Ǌ�����$0�8L���P_f��Pkp䪜d���FU}�U�AG	�t�����6�tyv>���Hvdr��m�(��;��'_}�~����"{��-=�MԢ��ʰb�LP��ۗw1�U��l���^~����ٴq��ߋ�T�>�9��V�!��߷6����q��0��b���s��j�Բ՜����?��.��dU��]�䞎��&�j$\���Y�!�%�:�G�חe����*1E �d�Ol��d�	�Jf�N�yc�mjW��[۝C���ڿV�ō˜���U&�����JPO�G�o�ש���q�)�t1*\A�gfHu�Bj�F��}�'��L�,<׼�  x⻐����܋�Rnt�#C�	{vzf�Tޏyl�c+tX�Bd�&�R�d��ie�L4x��@�1&�*N,�J}Ҟ#5%�/'����n�T�K>M�^�J?��4�|��<Kx ��R������K����O���o,y�>TE^^Cm�qښg�t\��S#�Vz�*�<[DC����p�ɥ��!y-$�aPž�/�b��h4�c}P5i��m���F���"N��a���S�G>����-����Q7��2�*ڂ
x�yxC`��V�yj��>.I����ItR��zks`Ù�l=g�O(������{��Sp�������E��j��c��@�`��ڧ&�b���^R�����#�#��3�^']�gO�hp��$=�O.�=H�@H���㣋��]L{�����Ù�R��0�_���m�⦡�3{��/���fǚ\L���p�t�N�;�I!i�z{h�q�����a�mw�X�����w���w�������_��g�LFŴ?��LT�A	qc�Һ0lV�,$���Ђ:8���V�G�����6i�
L�0�g�b,^� �����QH����đ�/~�n�D+��W$�CD��d78M���|�Mu3�w)FDx��\�pA�JP�^��If���<��Uk¼dz��4G�5�\^����1l4�Ϣ��{^�z�D{�!�X��w.p=�ܜ��S���^��(�nj�qe~������M=~��8-]���P�)7�6O����������`5ޅ�^42�P�G�&�('�x�����nha���Yzj����̸�yK�W�"~Xވם��a(!�grl&�\��".L�n��L��z�g�0���wz��괰�3|��Q�߽uX �,����'>�C	�b��X�?4i�)U�!]O�emjF��d�W_��5+1}�Q2*1�]pQs�p��\"1��Bs��Е�z�z�,���n$�Wa���U�Β�ǚB�(M)�ISs�fPX0���NJ�M��Jx�/�-""�#i��-��:�\�R�SJ1��jGov���d�T��$t�/�:�cŽuQ�!�z�Fb��C�L�%6c�r�u5s"lD��}��ޠ�o4{!�<��˾�c�(���İ�XgZ�j�LL�a���`�Ō�;��9$���{�浽��l}kb��A�|"z�"ɣwk߶7��]c�o=��9�w������`ċl5GE�g`���M,<���򦀎��B��������������O�
���p97&U�>IJ����Y��[7����AIoN5���Ej�Z�k�"���"�V<�?��.g�0���K�Q`�)D�E_ʁ
Ґ�8
 �-�و��0sr#�4�J�ʣ��2�*a��Y��QE@V
J
�56tE�
-vP�1�Z��$����U��T7R�ĕ�j;KDn���0�a�����Q�ǰ]�Nt�OؼL�pI���]��-*T�.���-<ӛ���!�1M͍M^ͳ\2�5ljJ�v� �}ZaG��=������/_�1}6��w��0�n�~l���YW� |�}� ɂv8� L74�x���{lpWy��-*�#*&��F}VC�fN4��B�`�l0��JR�I�:�,nMa�U:�� �����>;;M��������OfP�{у�SqN~Z�	�Ө�_�k� �r@^�w?84�KJ���<���e�D2���F&�PW
<�2�B@��y�.���69?�v���$&>6!��qr��k���u3��,4SQwv�b/i���g�2������!�#����f�Sy�%I�jr�=uURt�M������U����z��;�pf��~���sAT��=:�τ�p@�G*�X���@����LM[���}��u�R�8�{��>�kR��\J
T5�v���h1��h�.l �wgI�?���ԫׯͻ�c!H̆x����VO'��w���ᙺ �g�k���h����֌�!'`%@wޞ����P�
�l��% r!����W�d��pC��E��w��� c�"�`���H�{��rE��'Ӽ���Ȩ2Mr��_q�Zi~ޡj�:�|uE>4�"���`�i޽wwތ^]L�!oJ���e�#�Y|�G�1�F�(�T���W�ԝu��ʼۊ��-�h��V�+~�q�κ�}�ٍ;��GAp�wlj��e�L� *��~O6��0_���&윛�#zhs�7��Ƙ���n%SGx^j�~��5XR�h���T'dZ#m�EO���7�BJ�~w�
�꺀��>�����
�-�B7��x/zWFJ��&ХI��
R�_��"�9'J����"�п��{˸������G��-�-�d�s㨢��4??��]wYdK~0#;M0�n�9��8���t/M�����Х*�l�4_�A�<RE	x����8w@)0�,��&ũ���I��}\�B3@j`�>�YUbS�A�y��(�*�a���̘z"o���4�f��$̢OXI�Z\��M��koP	�'+S�؍{�]٠v�(Ł��k�(���x��ݍ���k����<�B<��ܨJU�E��BA��KyB��q)|�e���K��T��B#�	���*!�揩�����W��U�����ͦ��Jl�/�7�s�%6������װ��5��uaaTG� N�g]�՘��Q����x���-@ ���� [�VM����V�������� o��}V�D�T��RPCE��J/ɹ��=�:�G�m�(�޹e�n5�ӎ�B��r��TE�'����&wG\e����Ŋ3�'��*����S�0��Wa����J���0 ����Ҽ��Z���q$������i��0p�&~��膠LD";����^  �T^�����c5�;9,�S���	cЧ��<�`/H*҄s4�F�_E�Hkz��<��6���ZkR1�ڄj����{�.h`� �������<�g��t�(R�j(o�q�c�y��Ġ��E"�,oV�������S��
[�)���JT�& &���{[\�m�Dx<�?�ǭiZ�t��cM9�Y{�J�w���31��Uv͂sNV���,��n-Q\K��HBGwS�v�H��9�:wR����΄5p�(`�|�����tMX ꫪ���:��U�at��8���4U3�P=��&�\����N..4U����c#�Ta�v^�
���U��hao$hJ���zA�B����X��i��a J	̓hs�<чDy�?��]ޅn�`��#A*8�E0ƫu�@ڲ,zK�nr%*��a�(�{��+����#�qqn���@J�M+m�6L�3'eƷ�0��{U�Ǫ���*�Q�%���6�
��__eoʁ���{R(�O�4X����`��S���{b"~��ߤ?�H�~��-�ќn6��ݷ	�C�Y�m�=z
2:����a�ob�
��E��%�+�!9�^B.,9����7��-w��kqm�^�
�Q0���0�)�ζWޣ=�{�ZbjGa���
��	h�	`�x�<A_D5�;h�����ϟ���kO5g�sohA��l�ý*�u��$�+x��Rq�:PU:w
�g�{c�H0����8�S�)T`�t�dŹXj�V,�7�ғ0ql:��C2������|�o-�K���8r��8IגZ�����o��h�6�aeЕ%Ji|�{�^�sP�����<�O���&]����h�fP�#9��Ul`�F"ܳ�o����㓉�h�RG��Z.���S��䕟Xa6a���SY_����.�<2������O��ܻ?=z�(=��K��ަ�O�7�s��]�֧���MS�RB�9Z%�DL��$8y
��`��6��S*/��e]�������2�OYk�Ja�mC�=lt�l50�imF����"���@q����l��C׃��
��6$,$����F�꺡����m՜�R`����o�ۻ�q��O�Q���|g��/�������o�3�N{�Gg��y�6L� 3U�T�I�HH@��3��ZK�ܴ��y���N	�u[y�Pn,xň�i�O�r�AŸY�r'9�Lu���z��դgޚ|�]��;�� �Ź9`@�oz_3~Sx���`H��j*7��YhU���Z��2RJ�qP�G4�?7��(�{�_����4��ӎ%a���k�T^�Ҭ�$�\���[]���3��<1i`���k�L�x�grc����u�I��(U�5�<0�id=�c�;O3���a}^N�IYڑF����Đ���j1c�>����ݹs;}��7V�䘠ӆ�0>�}U���v��P�C4���ra�/X��zw�	su�;oYR�ز�j�f!��u��`{�^LhlQzZ�<i[n����S^��j�։�L�B<Vc>{T8�����h��Թ����0��9+����,��c��i���e���R�=�(�L&Rӆ!GV\z����rVG�DS�bbO|�!	ѱV���í%ܐ�B��\8�!5z��;���X�L�9��*�fj���9�h���r��\��,)�p�%8N0Rn�˹{��U�r����_�A��J���r��
S9��y��v�}�:�x '�7�_�`��9�C�[&���@Qj�-[
]�T%�v}����4�Q��(k��\m���*G�l�m�IE¹ÐY�|�C�νN�c��V���a\Lggo�0�B�<!��<DE��D�����O���u���$$ �d��+M5Y��Ջ�'���r��{D��5쮬���p b�M�L:�� ��|;oB{��֣{|v��Y��Ng���ꍫ�Şj"�綢�.��./����#�DU�UL_{%�bٍqO��tow���:����b>�1e���b��}����+�t��}$����i���U�R���ׇ��L�o?��X>����6O��YӲ8y�x���w.�b{	N��a
B��O��	%����5����P/&/�:����$
�4����2:��%?A�5��{%7�?P���6[Ye��]�<cGS<����/~��� �u�XQs ���<��Q���� �	j�J���;�u��^G4�n�WQ�ޖt6��7Z�&��x�'%˕_��4��T�hYn
5�w���=zDZ
�31��4��������DZ�J	���M�*�)o8�i+;�#��sM^�ހ�Q\�^�	��R�21��D*�yҩ�V��IL/0��W)/7g�<=p�[H�ݚ���Z�}�)�CyL��v�?�gD�f��lg���9����Ժ�hL�����KE؏C���%bk��_�Uz��M������y��9������=KK_br(�3
��a1��^[)T"N���(��B�y�z��Ax��B���6����{5x�Ą����%��y��!�ٗ��'�WyA�U7JT�.�ӷo�ح�wݝ��Ի�A_�~�����$TӀ{���FUE�Ks�j�q��$��,t�a��7�G�2��F�6��ԥ�ئpI.2�s��HҸ;�"��,Ř��I��x���:�PKx����qbL�����&&�-����x^P�,jP?o0�-�q~^J��.����B<}W��6Mk���hH�Qɭ���5�!?<ҵ)M)����ս�Zm�1�����sZX�&�Q��0�!�����!�<�z�l'ˆ{r"yhNEvTI��w����o�����8zN(LT�(B�(8T���7��"&�š/RKt�N�|�T��ABO,}�J��FT��ƁV�b�[ے�U��b���yy�;[�R~�Ƃ2ʍ��&��ц��#�쭫�7���-��"e
M�$`Tjچ�a8�\��c��K�f���uS�A�A?��t�*M�Ŀ�{6_}��e�_�|e�dؐr�R����v���;�ǫ8?*�Zc��;��،0^<��	�xIH
ѓ�鄰H�A�B�(���<���y���&&=�a��aˣu|����?^e�k��YVF�yw��mD�ztˋQ`DYߏ��g:���b��m<����͛�0�z3*���2+̌`��;��&B�7]�?�۟<^�� Y�^��SV���~�B7k/ݹ��Ixqp�ݽ�~C��R��8~0H0T��Ȕ'#O$�4��I,pI��Ay�v�(���f�|��${�����0끥�loa��I�]��S	ݎ�P��eN�̭�QGfХZ��Lەq]�����G.���
X|������2�$$���G�����{�L��yX)�P?�0��?�ɩ
o�#���t|�B0i��m.���r��K����N�=I��zw�E�Bi��M�ɧТΚ�(% ��Ja^(��<�=G&0�w�9��CpO�F�"�*��B�a����E����E�6���b�j���cP�E+��v���i���!Й6����f����?��?X菶O�=��P`���g;f�#cE���+�����r�����5�|��D���L��<��(O��CJ-(�<X[��^n�G�����s����T( �e�7\�Olb#1��e�F
�1�/��#S3����_���4b�5�[�W�[���s��K�7�E��1.v��{u�D𘞟׽�0 G?;��hX���{~�s�_�✒ޮ,:�0 �pː��=]��0Fh?��jx������g��Ma��ig�;c�
��rCq��h��`^㊨��X����Ն��=����߽w�q�c�d��#�h��	�DTq��O���Ï���p�&Q�7Ƞ6�����7U'%s��Y���B�-I�T�A���B*	<��s(h*N��Eě�篫���\�	W`Kf��Ӷ�̆�i����9����yb!�w4�����'�[�{V,��*.T��HR"�ڽE3�ޤ�	�ͱx���y!�Px[[	�}�H�߻o��j���dH�Y�%�d�	w���k���^�]M��C@�CG�=3>�`� �6��m�x�������#]�;\��l�2e�`�,��6�bc�!�*J����kCD�g��Սd�|�9ᐧ�5W#s�R�}��G*����-з���&h���g�����D%lF0�Pg{�����1���N���~��}�qﵹ�Pׁ���F��h�P[���cP�(��0���O�WOEy�>�wL:L*,�[����o~k����oӟ��'�B֕t�Pm��6��R�J�KI��'u�D��sZ�-Џ���+�OQi5�ނ���P9�����z���{���_K�?)�0L4�4Q~@�+,��ņ�3��UfhF�8+�<�� B}��{���
DnT��$a�%�Jٚ1-���"������{5l6B��ɻ�.��8V�������1�ϛޫ/�2ʸ���U�J�MBq�;�����x1�K���Q8�ko4q��ub3�����D	i0A�E)/���Ό,6`�0����c�=A F�b+ ������̾(r������庪���0����6v%"�)���w��7�A��y�Ch�68�й�j���׳��!ɻ7o����~={�V�\��۷F�ί�?��"�>a�yڥSORY�(�
-�Ja�l�1Zs�{P�І��t)�%�f�l
)Qe�,�D(n�9]�лA���}�����бVSg�=9$K?yl�
��#)L���qa���(���b�_5������&��P�����o�И�RVc;~f�&~,���Ȩ5��y<���6��o�?�`����D�(�K�Ԉ%��#m���ͤ=Ǟ�t+�Ɇkp:�U��$��Q�tx8�I�L�Y8�d7F��a��n]H�\S��;������޳���Q�7υ���9B;8r�C�&����d88��qG����;���cP���M�M<U�Nޒ�0�/p�	�?��<-��������e�����n�S�f���e����Ј�V],6k%#ˊ�cb�0�H~]Z����j)������>���ԟ���[;Ef����]|e�][GOD��
;�Uv&I,[Ki��s����	0>����z��}�}*-U%�F`�'��Jm	S��z"�C��5ɬ+��%��wGl��2�����d7ěA�0�
9ȶ��S�x-����{��/���hRo��l
j��H<��xNO����&���KIʞ~��z�(���\�x�o�^�J
��}bn#Q��	e�p0���b���.��B�ɸZw�����+ɫ�0�����d�&��E�.�J�x�DIW֓�*װ�]r��7B����gT��:�?��-�׃Uz��A�> ���s��Wc:�t}Qd�o͞��0}԰�����jŅ�W������0��33p8�KXD#�i�X{� �*)��ێ
GH.@��ڭS	��=9�w ;��������[x����;�g�
͞	�*��j��JDu�?=�֫Z.�=��6ݵ#�	͸]Ysܨ�Ԫ'o��B>ٻ�=�Бq�j��#�k-)$����G�)�S����6�Q�7p������5I�	_Bo�c�65@�|D$+���Ӭ�{ؘ���{��m�v�;�w��+�l��� ��T�3]������Z��c{o��aH�x�ȼT�tQAj�p�;r�c J{�͘˖j�K���X��8����^�R����y�G+'�8�1�������}0Hv�rb���{������r$�/�ͪ�i�5UB)�P�_F�"%e�z����H�٘�C�
�9A��ݛt�ޝ�?����o��o�o�q\m6�6)� ��OG�|�훅���5�yo��;�6Æ�Of���	l4Q���T�Q�jҡU	� 4�3U��3��x�s.�DY6pS�:��� ��jVwe��.���(��n�����	�4"���s*CcڧS�����Ќ_���Ͱ�v����"�+n��?]MV�siy�$]S~k����� ģ��Z��O�����6Z����o����GG�4��"?T�U����0���M�p6�V������ĹےӜk�'���
��7ժ��+��9�D#��g���F��H�B���mJm���=�gt2���X=fщ�s��.s\��O�c�0ui߲i����֨�X��t��\C�����2McM�}��/x�"j����C��򸊞Ex�<R�Y8/Jr�6�1���,(.b�?d�Ł�bgK�������lg�}��'�(R�ԒOx�̀K�3�}��g�^C���g�k�����J��ޗԃ�e���Z���t�s.&c���	�⼛1������R8���gr�H,8���^WG%
����4&]��@1vp���?��fr(O�*�ئ��dq�h�������vO�o��(Q���i�����2ݭܢ��q��-�Et�%o�6�N�Mj���M�!B�_BBf�c��z�ZO����@�=���{�J��{	!n��Q�6� +�IHl(�˙¿B}�;jD�aj�]�O�Kc�Z#��Eڏ���ROe����6埀~���`��G`v��ZC��Ғ�ƅ��5����{���%�U02��?H_�����������_�5����_UF��j�k_�Lp�ը�j��Z� ����<#�W�joi2E�+)�����#tEk�٘
#�`\Sb��l�j�Z��ވQc=�$���>:\�[z%K39��	ߊp�����]q���c�_����kO�br?�Ǚ^�f&ּ�rC�����A P�u�������Eb�d)V���gڷl��U��@����%�i-ڶ�	�e�[8��)���_3���Wڕ$E�7f�<'
�絨�뢴�$Hz!�7����:����"��J]��ds5��ދ�Q��r@R��?u,x��>�X~F����h�hV��a��z�lf�U�X�(j�b1 �����H�߿����[}�^�����Gs8��P���b!Hl�(7[�����0ޓ�)A%(Z��b`I�I	�m�OZ�0RV�;�ί��k�s˳�_͛�Ĭ�DOL0X�'LR�һ4F݀..�]�J"�K��3սC�:r]R�>_��
c�q��T�A�;�O�4��e`�|���֖��K3�B��7��0ze���{�ڷ�y�P�}���~g�:���cM�p���fyiђ5�$S�
P�.k���X#*�f�
;/%>�N�ITCye]�C�Z;���ڹa��bc�n�[Um���M<n�Am=#���تވ��Z��X5O�]��a����*��7���	�>ThEc
#�	c�P����e,�9�R�O��o�$ͮ�9u�!��^ع�ih<�D꾰,>��g�:����$fO�����wFچ�P]�ѻ�ݠz�еi�L�*hj(1�������ܛ0o�~��`�Ô	�����r�TL �!s�B�yS�#x���C�y�����ӷ�|�I+_$��&}�w^��MN�a-�"��v�]0
�7�%���<��JAckr`�u�ƍ�H�x�r��~���5 �r��:�R�f�^P�x<:5�pY�3�b�M�Z�zŘ��������4��y���"y\���,$%e:
;�uǸF���~G���H����/�w�}�����K���7W�G� �5V$Kwo����ڕ���)|�Ih�j���*%�r�㛦�f�$Y�=0R����<��!�������IƣG_X������^S�7kH/���}K`�h �&����/mM���x�M��@Q�^^��x/���Ƅ�O��=�k�P	<|`����¨yҙ}'<�#J?b�R�ͻ�F�ÆLr׳��Qɨ��z��� F�'o�۫x��H!\���^�djǤ0��[�w�G
Cz�$���3U߄N�!��d8�ttγ���Vc��Ka����o���r�,�Z~��+��"��NO�V�Ԟ7��nX!>�CO��9�W�!ҟ���e�/X�hd��k��y�cҾ�ohH'����;U�o�ͅ�Ʉ)B!#KO��!5������޵K�#C�+N�=fh�C�L��1��e\)��]��:��5��r|������/F�n0u��]��G�@Uf�=�M��JN� q��L"��1	H4{|�N�f�?a߀[Vf�����6��R���j#;�"��݂��nj�+�����6�6��>�Wz˽ҁ���h3�f�ڀ��@r]��'��M�1MW�����<S�h����R�˶eK,��I��|%12�0U����9i^ = ���W�B(x�0Z����!P^�:��3�m�Д�\F!u�V	�����������*����dr)�۠a���]И���KW��\���I�v!ͽT�V�|�p�z�5�k� ~mƯ�*h�-�N����ռ�� �@WZ:���%�`Po����Z���x��ٰB������%[�����ʼAC�$-�d�e$�*_���MY���M���q�;�cd��-nQ����J�����ʓP�6a��=�7
%!���ަ�0����%cz�m�1��Y~�%�7/���2����d��0���8�&��
�*BD/,�3*��0��~5� �|�浵PA���.=}�Բ�;���>s���_o^���@�W=�̫�mnP2h79YI�U�t|h���*�wb��;s��PIBƙ�.5r3�j�{���w":�~�)�C)��g_W�mޢ��k&��R�cA�+&Jl�jAmUh[������I?���h~������+�T�	0,P����O����|�Ҍ�AJ�7�T�ӷ*��B�TF,Η�_֭�� ǶW1_�}V��h��œ��ֽ;�X�z�
-�g+m��uTS=%h����{ē��5ƴ�q��xjT���6�7Ƞ�kC�@:B�O�E�>�8(�lm���-���c�SX�h�p�N3���p�������`������i5H�\����
��)~b���;��(K�Փf#���ڥ�(�w����a!y��A���}�20��j.}zI�-˅�D�u���c��:�iP�0��T����!���8�� 3���V�'�8�``�%�O�������Y'譾����_\�~hM3��;����j.��{�g��ϱ�^�l��O�ܟ��.�F����(tk�F݅�ԩ.���	B�0�V#�)���isC�ƴV��V1��������Y�sZ��;�>�ZR��G�����(,�Pҧ~(2�^��,,��B������	���P`k����}9Vx1���y}�sM�FH��sϊ�Yc�8�p����͟S�;��T&Z��pXGL�\"$�,>k���_x�<D8�ƵR���n��es+w���"X9u�U(g��F��*����0�y�n�0t���W���w���'��7`VP�����A��7�ҳ�k}��Mzw�nQŤ(�V߱c���a�G2I8�ɉ37�8:�B��rܦ��r����վp�S�tߔ`j����t�j��c�C]x��]�u/)�W �����o��E����4�n�u�N2;�n�Bd?]�ɱL|��@%<��t|�R>~��� ���/���T[�'][��6��K;�(G7!��e(D�&y��0אmɷ���55,� �����sf��ɞ��̦v�Iy�'V��#<������k��:����BX�td��	?�F�FH��@�6P|������j҈�:1���a��䭍=恵�g�p�2�Α]���z��15l�z��)d$@����>�Wy�"�c�Q�pӈ�TE�"�������Ԏ�{� ��}���|��Ij���~+M|Ѐ�Y�E�`f�Ҋ��37��$"�'{��~r"Յ5�Dp�Vޑ���Ld��l(]�ךH���h4�ب�V;����ŝ;.\m�k;[��T�Ǩ��z!�'�j7J����������{&V�h�i|#{Oc9�/�S"����71�-�^rd._�����&>ޜ�;�5G��[\���]ӊE�%4I����1�|l,��}3F��_��lW�dj��<�ج�k�l�sr��w.�F� 1C���ѳ`@�"�S��QIϒW�-0�H8�3�׃�Z�
��S�s�x�I���[kw䚡�׍{d���uO��KY>Ӹ��ק����^W����d�(u�X|m&�[z���ͪ��r���[{\����rj�?�,��d1s}ng%�u�F���:��<��n$/^��h�Zbi��g/uϱ`2��/ɚs���x��ku���e����b�,-�-芘�~R�w1�"����]��W�����80�k�^�x]ȿ,����~�;��׿ɟ�5^�h����J��F�KMի��`�0�d���ܲآ�9!	�.#��0{�ݡy�uS�zQ��j��'L+���u|��������b�:Z,��fA}�Q+!������RA���WQ˃~H�A}\��??ZU�Y�J֚�*�s]���ObP+J���TOf��3���:��Liʑ�����[��k����M8��.�t�J���/<�qa���)<]��&GNi�K�ԉxJ��c�ghiOբ޼ky&�S����\]bl�,�V�Ҁ6#��}>����3$���:���L����-$��8���+�{�w׌g�E��z�u<<Y	5�����qW�NN��O�ʧx,�Ѿ����{�O�W��1�4K/���ㄟ��R�x~����>�[j<�^�^���9W	7���	����bQE��;͖�9�AW��+���'*�TM[C�+��D��j�R)1�fU��Tᕖx��A���^�A��{���٤�%����a��4J�`F��W��f�K�W��y�{b�횊�Y�'�S[Ds�5�J6��0�%6�=_��������'�Pm`��z �RǾW�>��Psd@��sb��)�$�-���RY}G�Vj�<�K��a���ޛ�7�3Y� )ٹT�=������t��k�tZ"qˉ��,*%�2KQ�Lq��XP�{�4 ��:������U]X>��;���(�K��^	��Qt`��ud�q@�߼��j��zl���ԟ\������)4�
��Qk:����e�-�-�]R����Smwܩ�&~ߞ#�.�Nj�r��uЄJAvJ���	a��_Y��{�8��z�8#�}q<��p,�!�~��,GY_���u���+�d���&����t|�\���:vrU�r*h�h[!EM%����E���O�Kd�͚Q��O/P��t!������}�I�9(�SK��]g�1����}�`u�1J�!vΨ�6�t� ��Ȥ�s��
����H�CV���Mg@3ߤF�>_�-��R��1�J���4(߰%���أ����}���U�P�p�d ��ԙɠ���2c���N��;��l"���J�$����@ 5�A]����{�紏���2@�.F�Gr�f�Uj���A�u�+��'ZB�qأ�;RJ���7;��c����̼֨�9y��X��RM����1q��pҥ����M5�66\���P�M�c��1���P_� ��>̑�|K��i�Ώ�9��65>�y��M\G9U�<~m2�[��g�R�ժ�Z��}����hTz�UU�p��ONW�F�Ix�N��S�c$jBvM0��m�AU�!�������18�lr�D��f���i�^:lL|��N;FtVOY��n�҂X�tK_�/KS�J��Rƅ'�4gt��Ih@=3c��ҹ;��r�0qD�Jn{
��(�&���r%n�oo`�`УOri��lg5k��[���Z�pPOA��%�ɭ���_a���� U&IY�d�Ԁze��*���И!�[#���޾�$٪�)3 ��؈�z���m�ASO���PK�NI"��C��N�A�pܴ4�~�cZ�EV����ڱ��j�A����T�crNH�E�WTA���R���`C���ou`&]J�:$v5Y8�0�d���:����Y�Ԭ�^;������ ��
�f�����xW��NT��}ä�԰��2�c�<���P�.4:���^���iXjJ�d-	xX��Q[��C�Z M^��Y�+1�媶�4�#��]*XG������e�r��!LX0��b�t���y��@�GJ@�@����ݠ��y�2i?$P��YU'��`M e�5����LvfU���z�H��͞4�N3q��X��v�����q���֜�~��Q�`�; kig�$ޣp��Z������O�4��$e�	���C��6^��̯���X��o���8+���LTt�P�s�6f6+����78T�C%���[��2Z��`��ȧ�ٖ^m4�ڈ5�+�6�V{s:���yx6)P1yV*DJ6�io��g5~9I�����Z�]��HF;.��!��c�۽�P6�d��Z�R ��e�Y@&��h(�Z�A� ��r%@mfqt;�T��&��o�#b�r��ג�������R�]f�.v|.I�ɕ�wp&�#JKz�+�
�Y2�n+M2s�'4Ęjc	6V�.3���uI��A2��@'�`Nx��yg���'>��%��Bo�R�2Յ��&H�!f��hS �:���P��t�� -	�ύE��],��T�ЇM��ߜ�*�@S�w�+,=kU{�����}��bs唣}�=�����&�r��<Y��C|n��1%�b�ި�x�Vtƙl P��5\_`Ș�WD[���OlB�ܒ��D����r��E ���������i�P���Y�h�Y��A�0[�l@n��͜&���|�KϨ���N�Rq�6�\_�׶0육Ί&\ܟ��>�Վꀚ��
m�P�IV�ɳ�R��"�	�-`]���5R�������v����p�2{�=��g���eC+���:��n	 �F+��p�	f���ن�F��;tUt��3�cϓ� ~ڈ���~��V��.��Pg�0��Hy���^9�������\���A[�~̡a���REx����9�C�9o k�0 o��F!�;T�G_��~ǿY(�����nܔ�(v���Z����fך�jq����)_�R �&�^H��:x��0a��+)����VC4�R��:�&#K�Q������r5/?~�!&*�&�h��*�+2��v���EJ2o��k�=�4k$�lZH�\1��=��Δ(�7�63� d@7���x�����,Ƚ�@�)���k���������OR��u(0�z����o}�7�b2,C�VՁzO����˰�[y�_I��"�@�]1��@y�2]�X�O�����,��ǓUQ0�g��ʞ�G6�,2�m�S���ơ�A�f�ژN��I�Y<�gO!�^OY�d����-��3�ڀ��5���{S���� ��tft�Ȕ걯�f���f�چ��3��}�R i�P����,)�������Z'4�7��c�Qz}*i�Y�^B�M1��A.�WΏ�7[9ڢD-��bFQ��9YJ�>Մ4����D��,���H\�	o���9�y�	!�k�c�����0����rOr��R-G���@�A%�a�M�)���χ���Ս�Aƅ��)��nk#���-i�I��uP����]�G�^٭J����X���[X����V�����5�����M�N(��"��h'^-s�|�(3�I$��$�zV��a,�loϰ�k4_��̲'�Pwk����@@d0�%;Z���/	�%����u��P��(m�����$��Kn���U�|�#M�����99C���4ci��n�e��
��)N��-8�)�u�a�03O�ɖ�2���-]�;+[��6��(��铣r����K���ͦ�yf��ɲП+�
#�w�8\?�;�n���#�\y笉R�`��!b]�JB�"*g�nC�8����Xs�fQ���뵣��a����4�2����Z��>�y	�U�ո��i<cW\լ8!�<҄Q:���	Z��@���P�o4N1D �% =���FJtvV��T``�gŁ�~�EX��;��:П-k�e�	CHh�p�� \Z���]ʊ��}��udt�l��?�r�_<@��u~��:a�x�g�t�Lk̸��!�`�O��D�0�,���m�Im莧����q�n/lY�嬢?b��,H����f���{#�u�-xe��=�2z��x��'��Gݓ��jaS�v������TN��{  �]�8��X�������gF�u��r�Qٛ��^��.��z�s�U2��*f	�}=�
�d*�>)tt��dlWM8��V�D�_& �XN��h��掅^9)���d�"�?]�@.���9����&gjuhﱌ�3�2׭;�L�_�� ��G�U����Q�㳶�Z5�j�
��c�6'��v��A���;`܃\_�̔�>KFs���c�`��`�?��ǐ"y�+m��h�4��3{1궦�La����w���S�������C�2:��`��3~�bڻ�����L�o��0S�@B�3`#�3Ń�Q)�#�����58Z7�6i��b�W�ٮn½b`���|���D�]Ut�X��7mA�fg��-��^[9騼aLE��`Z�Ԯa�5���� �Ŏ˘��hy4���ؽ�h�,=�j�o"�ӭlPi�ѷ��ƥ��-F�q3�K�U�>e�{��pGv��߳�$�X��-+ZF�w@�� �5�l3��*�ұz0G�_���`�6F�s���@��D�k�?'�iMܾ����0��MI�3j,[]wPSuL��<�v���:�W�}G}�Y�4c	�*���%�?G�l�h��M0)���ޘ~cǊ�.�㏔�0Tg�O���nܧ'u�p::b+�0�֗f�	{���Z5���L�9\�g����2�5�H{P�~�H�G����iF�y�\x�6��d�bL��5��Z������ϓm���PG[����⚓v��0㨞�����~��P�+�^k;}�	l~��a� J<��/���w��O��9�� ��>	L��k,`�?��2���tol6�8�4+;�~tO`Jr�-P��Tݧ�Ɲ2T� T3o�jN�yu�������	�� ���%`��NI�R�=�� ��U{����##@nԖ=���tOڭ�Z�Yc�^�����&��J�m��pd�9X߷~϶��@���ή�6��=����e�z�I � �߷e[�_|?HX ��O�)8֕GQ�:D7[.�8'rE��ZO�V�p��/����)'��/G�S��T-zNg{h�D�f�\PA�Q$"�cC3�U*�i��*��-&�0�����ys��\=��/����%e{(�Ja�{�q�e��Dſ����5��8�)d��Z�������	�����f�Ť8oKm��3�%u�����f�c��k ��e^��P�_����hj�	�q��8�;�2%�xJ5&��$p�q�%���Ձ��  :Y�9j!���όjC�:�a8��o�R���ru@��T,�E��4��d����f�Hi�����0#��1_hq���a֙Jd�K,b���=)�iJCzKZU�1�'6E9����6�>��(6�e����d:%f�� �5�R69�.y��O�!"?t*@�L�Z��� �����]��7����H;�� c�:�p8�F�Xѥ��Qo��i�6TMCU}0�jW��6�].�^����<̬��/@Fx�% Xf(x��b|��r�,q9�Ϋ�,Vk^8g��U�v9�.3����k7�K����9o:�O�y�f2�
��չVx��N  ��IDAT�2V4K� ּ�`|k�LhK�Xd5T_�-*@sc�{̷�&��!�G�k�z��Ƿ��Z�u�� ̆)Yy���x	�.������Ϋ�`�/����7߶Z��\���wMk �]�Tj���y�7#Q����K�.גM�抝:��j���Q��v����&<�A��Pc�tI'��=��Ep6*p�ar����Tk $rNU@�^�P�;�bw!��y�}�Sd��W�;����;�P��RY��9��.�z��*e�Y�}�^8?fǿA�)h�5�U ��,��| ��y�+�ރ�V	��R4��O:��=v���Yp�Mo�r��+V�1p����Jn�8:PF��y�y���(���T%X0�{���N�ۮt �7�!jC���}�.Ù�)�TU*\߰�%0ӱ{Uq�ɳEαG�%Ϫ�D�j�����b�X�M�%��T& ìPkYu�Tr������ʥ�]�X�;��<#Aݗ�!eaɫ�=�y����V�Y@jP?>��!sR�o�Q�K��!$ឍ�~����?M����XZV�ߒ5�?����Y)L������u�*��w�ܬt���@�<�c6�e;��痩,��i�@[V��-2�f���(�29��^w}H�u>H ����]�r���]��r[��Ku۪��=j��ڋ\��<�>���Q��7�>V�s$o%=;!-v:>�Y}.[��>���(����^b��U�x�R�*X��]�����a@�f���ʜs�)@u&��RG�u6.��n*V�å����&`��s��qyK�-��ψg��Kշ���\��.�gJ\��,7`Y��V�c��Bo��d�WnZ�u ϶�.�����	�m�)+�����p<��S���bm)S�qTM�	��
�����R�?O�F�i����X
 [�S�SY���$K�%7�J��<�,��K�?9Tj
��y�z1ub�9��<<��l��5Z�l� /�>�VfǪ�-�w#�e���kE�u�fW_�PK����99��h)�������N0g]��ʶrź��W�g8�yNہS����K�J����p�s�6�����+�{՛�0���]٭h�h\����Kn�t�u�����8�@�n��+l2�J=�kڙvɱ�r���l�A̏����2�w��I�չ��)��A��j:�oa��-��*F�W�R��/�I*1�g���R�>9���
*�S���yb��x����E��lц�٧�t�o�a�W�>��N��tA�X��O�m��&��4Ŝ;/ʶ��ԡ��eV�0{qΕ�=�`ۇ���/{Ƃ�j?M�m	�Y,A$?�G,a��3�_)\�~ ��$WK0mcS�_�㛎EV:�)��2�G�UI5��Tqm)D0� �15v$�������0v�\w�y��Pen;I�ۺ��!oSČ�Dӈ����Ԗ�Nl�u#�v�*�2�s�*;Wʂfp�H��㢰�q[��b�5IAhW��U�rS����n�J��+ ������<C�:7��b�G��=p׫����7�K��0'��8��Թ+�J�q����O{Hk�� �=
��}6�g�1ܧԷ=i����*'��/�8돨'���˛�|]P,��X�L+e���$N�[.� �~��t~ܔ�K��z$�9E^���n�1�n�k��L 8�&�`�	�������nԤ(���̗h����Ps�����`�2�v�UG����p��p�,3-����h�hí���|�ra�_�ܭ�w��|��K����{��x�c.�hK��&���,Lf�M<��-���K�u,�?�%�i�����N&�z�c���G3��7�c9�M��sD�F����k�k�y�C�@�(�1��-��V��r����<�!���P�<�J� �+�&���D���� ��ht�C�ϖ�~�<��!y��P�<�J� �+ȶM�~t`�C�[�P�<�J� ԇ<�!��� P�%i!�	VC #w���,��X�k!$�G�u�����[�I����W�q_����}���N{�{�������%�?��#��e��ҾVL�yO�݀jK����q�mX�ss]�.���K�<W	&���Y��{�S�|�+6?��x�y"��"Lw�Q�*n��{��P��5�w�O.��eк '��=d�k��(����0��*]�&��{�H�Kl�~�m��=�g�;�3�C�ƽ{�@yȝ�P�(K���|�CN�Py���e���h�X=�Z� ԇ����z�C~y �C�\I�z���O�5e<c�_Qݿ4ֵ<�sY��޹�'�$���Ӕ���\U���7�d�y����	1��>�!��5�����1-��L�T�\Ͼ&��� c�s�i]�C�K�6��E���Yڣ������s�}
���s���r5�
<�Y�jVc:���� �Xs����?b�yA��8�x2���,e�3~zKۺ+�{��Aq��d�3r��J��o5�8n$4�����x����x^:��wKeؘ�e�>klt�U��cy~J#�$>[���(������8贿uUΎr�qw�\_�`�Ӑg6�%�i�Wf���g���� �Ҟ߮*y�#�P_H�p�ڡ;�|�3������lM�}�2�7�/���ϸH;�xM�%KIl�������&����"��~��Y���=�� j9��9r
���5�=~�=0��~����_y�e��vƋGr����2��ru�����C���*��1ը���6n�	x�V��Mt�������Y�Te
fUϋ�t�|	4��ʧ��H����2��Z��۾-W��ǌ��oޝu��m��)r3����0s�T~@`���"�V��)�����)�3ݣ��#�G��R���=_���c�������6�$�m[�w�����G���ܞ��l�0���g���o�!w$��^�6�����bq���w=�!���aS偕y�C��re��Q])�x�㥜�(ݖ�bAr���_m��-�*����k�o�Kk�˝���cO�ܮ]}���K֒nw��ع_9���̀XF������{����U���w�,�<����8ӏ;�t5o��P���U��<���D'�1���f'��s;y|��k"��#�� ��aN�5��A���б5&�2����a�g;���h�Y��"̲K]7�T����>���w��Y��+*[f�_hD\�������x�k�����Z��;ƊG��<�!��ٽ�P�_E����H�}�v� ԇ<��G��+@}�ER�C��7y�㏗�>�!yȕ��y�Cr%y �C.�������� ԇ<�!��< �!y�C�$7 �K�����w�D��4�r��S�������s ���?��h����oGN�Q�ں6wLè�8II�F��R�n)��q��X�ۅ
ekZߺ ͪ��oE�?WEH�vh}߭�ڼ�O�Sk�+$�e�m2��I���,_�w&��$�������^�&(/��xj���ۿG��ߌ�LrӞv�ɂ!�TƑ���#GH�e[�p/S��jAV�N�;���5{�9K���\,�Nք	� %�}�(a�t"�=�4(�S}>�S��Mj;���9}�������8�b��k,ݿ�.{��O�M�W���˶�R�I/Ny�[��h��7jy\"���+�{����V��������ϝ�>�$��%��|7yHz8�n#�P���L���� �K�d�#e@���<䗓_Pgj���5V=��[ mX)�m?�!�5�T�[[��s�nlA�]A���C����{
�r�T5���mm
�ǿ{�y��C�(�.�fQ���1ru��_J�B�J��p(��EY����<�*��*�e�כ�&l�W��?�!�����w����
���>�!����W�����04>�!�4�>���;ö�xFJ���4s�ĕTe���/N�,�}��v"Iy�|=t0��צ����>���l�]����E�j��`7>k��8�,�s�=�B~�����j:Uh�5��-�dv
r�f����~&^ru@Żc�mj~��(+��tM?p*���{����w-f��~�:���x�k��jD��Yp���L̼����d (���d`�u<�4�ŒI�����D%mlp3��"o7���۽}M�w 7��|~����r�b˾�OT�/$�)!�E�0��&�A�����4�kݘi1?_�1��K�s��~�j��V�Wz:������?��/�{�Q�M��Zi[l���rZ��X��h �Hs�w	7���W;�.]�o;'ދ̆�Z�ĮQ]�HQk��U����rf�� ?��vL�W}�z�?C$[��k��%R �5��5�~������x�4��m9���(w%?��`�,���S���i�E/�mL��P˶>��r�7/��{���ٲ��3=���ju�2�D�ܻ��S~@Šf)�c��=���`*����q�Ƃⳟ1��r����5����A+;�gۭ�傦�ކ�ikN��y��ֽa�,!t��f�\
w�*�4��4�z�jW��샊����ܛ/���d誜���w]},�Ԏ�w,��K�]5g_o�Ս�T�|o}%L��:��K~7�2��O(?�.���SN���-�pwXP�f�n闯����J��޵L3��#{P�}���� U��b�������N�J���<[��E�J�V�����w(�m�2���`z�m�1�����J׎�_����pSIX���PL�pJ�UM���k���g�I�(z�٭T�{�Q�U?�f!jg�w� W4�7���c�i�F�?廫+L��	�䀪c>��A5��r�`J�j5u���8�pz}�7�J ��ٚ��n�֙8hb!6T�y��rY��@�~�hY钪�^6���zΖ�Pը^���y
~5�~��J��O5O}��PM��,��?� KN��?�\�å��IO�y �
.O�傭Hcl���/�9���N�7����v��y����/�^cqU[{� �w�<��`Yxhۅn�^-o���:������j���}+X��Q���}��ٞ�K	;*5�T6��)�x��mM׉�x�<��r�������T�����;�E�t�ö=�l�~d�95�W���X�=t92H���Sw3W��{�z�{�>�	8�8��������1ʺ~{N�N%��=��jSuȹ3FWOE���)Y��r�3�L=�6������r���n�T�5��h�ű��業�gK~�W�_�N�i���퇌��ߴ�ٿoo��w#����9���Z �a�`6-��%�I��OɆ+����*�m�=���S�^�@�R�L�Wm�ڵ*Y�{�Lr%�l���~�{�~������k��݌�V��%/�EPM5�"�]egs�Ƈl,ϥ�}eR8��Й��*מ2�_n�� �<��J���Z5�^�W���WC�U������&��4�KO�0e������ʄ����K(�..�Se_+���mnӠܫ9p������}��s;ǝՂJw�������=r�J�)7{NT��v_r��7:�����+S�!E�bu,��P�ZyT���Sh�T���x��kl�J4���O�ۜN{��S�
�惂�����２61�پ~q�;��/��n��ފ�T��<ԧ
�Lw9���=@��7�P7/cZ�<g�����o���9ЙyS�塤�Đx��?��Ë/���_O���%F�|s3�1Ը��|| ��{�s�~��x���:�t�sm-ljƀE&�r��Ln��HL*�;��V���g�3	j�rm��L}�
^�rA-�o�Y���܇�7ӹ�V�Tc�.5Խ��g������	o��L�����?�*�,)�A�n3)mg���7��.�C�A�\y�ʪ���#s�i�E�Y��~���ʿ�����0F]U�u���{k�bN�sg��N���\�{c���;�*�I~Ǌ� ��K���ݵ�mw�W�`�������5
����c��c6m�&�|����� ���v]���O�s-��~~���?s���J����X�Ȗ��s[�n��ݺ��+��D�-�K]�*����ru@5[M���s���6]2����5�4�4�o�q�3�/xӖT�sO�i��'�T��k޸G���{��|���7h������eH���k%m��U8n�E�uY��^��;ɠĘ�!3�[Q
1��V��)�9��#�b��p�
��A�͟�t�T�'�+�Z����t,#9T��l��;�U�ڛfq~�~�/|����O��7'�y�_���u]�]�Als��]�U��^�V���qB��w���ƥz�����7g#+��.[�MH�rtyZ���m3��A�Yy��f{^����`�����y�k5s�J��o��]��
�)�1"��_'�y%�z*C�$)�a`��s/�#C�A��
�� �b�̒�h�-��oe3R\�׀L��6�� ѻ/?��0�is��������� �~�z̨��z���+��-�Jkg�$����7Q!uA���	_;Hm����&���� ���V2�Sq�\M��-]1oŊ|�J)�%�0N�{J��:iuK�n��{ x�(�8����;��VY�nbC�3/ %�����N��=��6hf�T7؊�`i�0e��81@Fi�
���ܭ�bg��_b��uY�Oˆ�垅�o�9�i�X�7.����*�B����(a�6���0TE��~J20�l j����^�°����-N��="6DU?N$ݤ��Aj���������%W�%�)%Tf2�J�,W*T��6Nflt�b���K�$�^���E�^G,o�NP҄��cT�=� 3[g��nen���k1�L�@DY��U�ΗZ�y癉 '�M�3��lỶ�VE*.��
��؞�}��rm{��c{�	���v5��^��j_k����)����O�걵��__n��/�L,Յ*��f�ʪvX�k�ca��Wys�^�����V�Y�hQY�=�C|6ǹj��{��^�iqd��:&�0����ڽ�r�H�I6�3��^v�*g��n�%E�.!֔���)N��*���5�h[�������iE�~Z����3��h4*S�+��|	�s�}�ِ����&���bZ�5���F{�h��L�4��.1@����u�Ճ%��U���{�d�*�vkW��V��0��pk�yejm���1P|�[y��-iv%���s����$>f]φ�2�z�fbZ ��%ҫTc�rj;z�]ƾ><st��L����p�X�l��$F�&���>���$�U�@6�
NmJ0-�U�qC��C�zU�]N��JPn%?lO)�Ե��>#��rj�^��ޙS�j[ j1>�cX�sg��Ċ�V&��f��7��|mӛ_u�w1Z��j
_�7 x���Vj���{+��1�/S����x�����p򲭮~���"��d�'���ˢ�r�*�EB�4\:�YT����j?�ڟK�Jhu?�����u����62J,��,��N�U��`���=�(+ξ��i�1���Y)��BS�p�2G#�X!�Y1����e�聵�ߜ���B�����#���g�Y�5H_�C_��±��Kb�S�'��ݓS��Zcv�L��?j�QJ:1e{�ʦ����ab��p��ޥ�l�E�)��{W�M3�c	���8���f �90�h"�SN�������P 68R�Ylp�%�J#����y,�VY���XI.�鉧6f[rj��Ti?,�J����-Q�#��rQ^;z�Mp�n���[��vM$���o_S�{ͣ/`��M���]���/���g{W=��Q��x�	d���w��nEċ��p0�v
�儺��.k����)�� ��_"&�`��Μ��E)9�l�Rņw���G�ٙ���g�yߵx���x����uK�mb�=lr�_�x^�TZ;�-��:&��S��[��'��P;�������S1x�z^�@�u�H���i�ur�>�Mq�6&���Ѣ"��E[���nǓ3Q�����?�<�����9����K�k����U� 6���:O�d��-$��8T���X��f����"�:�"�bEFw���R��u���6A�k뛭��D���.Y�3��� h�k�s�k
��;ܥ�ί�1��;=��ťo�wu�,	H��F��mQ�K�N�%����Z(���Ѷ��������m��{��s���1j�����_6�o�/�8�����Yè*-�:N�O7��]|D�ޑ�^5�Y:zR@��~f�8)Y��ɒ���:�����}��i��P1��[��K�\�Nۋ6杣�a"�B�9g��Ǥ��C�������TZ38��Z��jn��>�t�Lא�kT�m�l��-����gX��N>�%�?W2X��W+��v�y�n��j�HbYY��;6U.�$�#��1T��(/�XR�XL�����̀]}�6�{^�ާ~�O����'���L��d�����zw"h|a��/��R�x�=s����ԝ^x7U�@@9�ӉڤWv��1��������V'@mXf��B���|�e7��Ap��"�S;#3����`��`1Cu���n���P;�(sRc}j�gi��"����Ń��M�>i��;Q���n϶�.7��`�!c���q��*�����͹��IT�K���Pն��#B�SP���tZ����S����LM�����mS��q=~h9|;�KI[t�2Ɍ`�2��T���K����1i�d�|������;)|i�]��"��1m�Xa���<��X����'Vie��i5T�I?`|�ygV��K��,=�Nޛ�7݃LG��H�u�ÿ�������{p{Ѹ"��B#!����2�A��PL�Ts�Y�+���Q��n����:�Q=��~]0M��B��D*p�Fji�l�,��K�L�6�����9�S����� �ǯp���E����2j����_�<t�;k鳙.�A�!'Vf�=���6C/��3Ry@M���Ax,���pH����<���?M*և�~��k-�:��՛����|��gf#2���t�U�N��E@�\��(b@�op�&� !4���N�B;I�If�dv��A;+�ȀO
�]W-��9Z?��T�שnILt"����8��͌1=��]b��I�=�x8�o�]�zu �VS[�v����L��0��e�l��	y�M���m}m��J�:N����G��S9���Qzn'�<�c?����^�uT.[�uR�<G" G���t��:���S����'~gN�B}�j��˞x���Y)�)�� G�1�b0����+)��b`cJUV�` ��͠��uʰ@r�H��Ri���)�ԧ;�����ej*����UL�v��,�P/*{9@�ޣ��uߘA�1.f��'<�b
�=U�9+Ux/���e��S��G�O�I�f ����Ϊ��ۉ<%c:�����>f�F��ji*K���O	<x��	{=l���KW�X_����<P��!&'3-tV��S�5�G��/��'�s��Ͽ�fh'e���S��NI_�~�"fJ��p����k�=�_�u1� �O��Dm�VHE��po��V;!s�"����Ƒ�`_H����x�U��1��J�FuL����K��:���/L$Q�����H�8��i������<�i�' e�����њ����:N)�1uff��bM�H�zrVg��'�y�,3� ����H�WE�d���-�:MFS�"�-ZJ>���t�'�1)��1�'d�,�s:�O�ϣ�˘,!ʪ� �����}�ԌтiT��A!�6T�We���Z6�Z������~N���29�<��ʷR�ɂefe�V�C��`E�l�W+�����ږ�� 2_uu�:CF7���`=BA���MM|�=]��[ީs3Cv`5���� ���jh�L ���@�nd5���4���L�Y���;��Od�e%*.ݏ@��@�ߑ��̠*�4��YY���:Qa��q)�G�{�Y�B_Y`�Ӏߏ�%�Jϳ\T�T�S=9�t�Dՙ�i7�3�ɩ�r�����Ď�IK��YU;�J�_�r@T-Ț����Tv�=��n���D@���lIr�M?�1Tv���gö�"����{�.��!m� �5��1)CS���J:���{1϶=ل;�Q]�*�ݙ�cp<{a�P��FV�T�Wd�v�>h�+q�]��*��~���h�$�D�}�
f
餍Q�Ŗ�f��1O�����\_��gQGɼ���=L,���Kzy�:ϑ���z�	+�M ��I�'@=���j����>R�m��I5��t������LD<�j�S^������kQE�%Q}RY_մBB��k�@�&-�y@���X�bb�>��ebv���'}{�����B������N>||�q�晃Nt��_4*a�)�&��?O��c� ��4Oi&_�|M���O.׷o����ʦ���}�u�O?�?p{�S��z��������v�I��ǍS���B�;5wd��H�r�7���Or��)��3�4w��l����_�Ec݅��Ħ�msb>��j�i�tl�Y՗��S��&�Fx��t��F�_���� >jP`K��QmP,P����V�Z������hvP��g옹�`Š��Zj$���e��zF���#��U�Q���:*�G��C���<=?M�{XT�d{a`�ze�%�Fd��%'���~�2Ӭ�@������۽h�����g�������N@��:u����q�?�s��gg8��8�8�������ӧOʢv��V�u�6���|�NNj�V~}R36���2�:V��f�O?�u����`O�����"�3Y�e�w�Ug�B�Ea���LJ|�h\p�����
���]����4A�
�����}��y�ݙ�Wڷ$����	��yO��J���4�rL*� h�N�Q� �Q3Nň�-�:6�P�E�v�����������1�:��0�����g�I��Κd���6GU�z���%yMpF��Ҁ�Y�U�]=$����Hਃ#�MU�eeO>(O�;L�Qfΐ� ��1.ϩ��C^�S�XToA!�qfk�NK8z�p����qޫ��P �X�_�-vou����;�8¶:�T�^@�8�>�
b䤙�)�;�}w�^�?h�Щi�h�X�T�Ԩ���I
�x�S�$}�[�:��cG�ij?b��v�z�`a��q��#���%}��=awO��5�oFSOe�oB�|�TqbudW5�e/m���$u��{�eA��j�0�؏�l�����R�%Em	�WR��i�=O�[8Tx�5��P�$���4���y0rz��Nl�$=Ox��������noe����x}�����_�k�M�Kjw��`T����L���s�r�2�i�P�ډ���<u��(`��FG�z���胛%�����*�&�kϝ򩲋yG�ꜚS��<�<`z3�[8�(�@�~؆��B��B�"ḻxN��0!���+����PE�g�~J�@5|	6e��̩}'�aI*�� �46�^�1o��D�w�"�n|����7V/���������f90�]B6�����R��zB�A�T��Q���=��v�Ws�*���b(�l|j]!�S�% ���.WOѯ�7��p��`�D.\�?���(�P6��w�Ol���6ޤ�(i_�-�Ɲ{c��7܆\��ã��hl�ɖKQ?�L@0_�3��Ii�:��?�d@�?;zu�a3Mӽ�S�Q�xK���Nm4|U#�Z7���5(��C藩2���5}�T�#��ԉP�]P4(F`���
I<�I]�?O��3ٓ�RJ9d�C���P9;���es����y�f��.�Q8�0��2�3��tQ�^r���GMn���F�]�	/X�@� �j�Ҹ�81�f�KB� �:�~-u��Hz]C���X71e3TfR�	��}.�O*1]���A��5���6&;���߮s�;�y|�������۱�!]p�I;~8#��,��(8�]�Y�HT�[����4�G�w%i�[�r�����o
;���R��������I���B+tv*�כ�A�<Yy�nEՂ�'=��\�کN��ݑME9'�b�~�	��&9����B �g���A��F��ҏ�⓲*�!ZHW�+��ڱ���J�N��_S�~�@��ǺIE@-���D�	T����C�܈�'	����
�}p�� �8K��]�E����F��+�s�pF��L-@¦Fc3�>�D�a����!�8ry;�n'e	��4g{���Z`]8^�
&�$��f����NT&V��"K� =��?��ZtrBQ`?n�����v�Ѽ���d�����$�LU�md> '��K�~����y��o� NF8���q,>�4���Nb��\WM��K8�2t���N ���*&(�'" ���;�U���^dBRG�j�`�R��ۙ�	��ݢl��Z�o��x�a��#$��cRME�����>z����n԰K�9�ǍE@<B�x���m}�Rؔ�J��ԡ� Mqe_H5���T��沍Lla�����$e��$��p�����U�;zJ��d�NW�P��h,�'��Bm&�A�ଢ଼w�ٳz���Ǔ�z>1�$1�B�S�1�'g�)���_��Y�������r����}�Z'�N2�9$L�xՊօ��Q�B�+qr-�āU�F�k߄w+�k�������1����T`��~bL9�}����~(;�Y��J-:�Ϋ�X\������������D�������LB�ѵG5x�)Έ���D1ƨ,W�≏�▟�����+#"�)=��P��|���Sb�-�N��L�d������C����u��ȶ��//LȄX��C`J[�&���XB�LJ;�s>�_C���?��"�� �5�K�#�59�eJg5lT1�\�~�X>]����1}4�I-eUK-{v���A��=5��WЈ��;�46���y�zBh>#x��Q�a�b��̋����S�/G,~]��Le�I�z0�� L`��=d8L��0�0p#�r[�"b���Q�'?�ϻ#F��=�J,�ep���Ӱ�4�M !���������r=����D�Ղ�|�@��W'�5p�Af�X��t��m<���<q�P��e� ���1���LE�<�qx��{��a!z���]�]�y�V��~�@�� +CF����A��L><�4(Y-F�&i��M ͓ �hv����X�c{{a�x����{�m�r��RhD|�ٷd��X8:�u�Yl���t��$od���|�x��	\�b��Y��*5ƿ�5���\�"�_fG�֎Wݨ��\_�.k�����vi����RI������BdERg*?�(L	c*!�y��z�S���:f������ ������ޖ\���&L�m���c,�Dk4xr�<Tj*Xu�:7��x��۱y��18sR��T�g��6�~�N�D[;�g�\���u37���E�V׫��Y
�[���u�.��f7�����󈉲x��1E��;�������������lYl�c�T����9����������[���JH�=��2�~}c����;!i�8�h�}��,A�s.M㒢?^_���`�QS�z�az#P����7�@NC!9C�0�Q�����חW��']VO�th^�1�����q,�+{�ɾ��l��-jtz(��;���*+�tR��S�O��������ET�v:��' zzڥ��ӧ�n)�頁�$��Bx^���M+gN��ꎲ�آYمih%����f���<�����V]#����<u�8���-��� aG�L8^���݃�I�H�|�_)��Յ�U����&��uv�FeF`�sZ����F`�wV�L�,;gaﯔ��K+����V^Z��U��9���/�6��&u���;%VH�[J�8aρ���	y(T�?������E������~�������P�ΰQ�tq�����ǀà�|�c��s�ؠ��s��I��v/BZ�����������6)�t?
��������ҤD�A��HW��%�C���F��>���9mac3{�Q�Ti��C+b���*���7aIA��:�o/~���$�Y��q�'P�z����K� *�E;]~8L�D+Lv�=>���Uc4��9�|'K��C�4��̣jS~�T6@��e`�qq���dC�KZh������1i����f��lp7l�7�� ;vf� a��ⵍ�ƛՀ@�e���:��r}�w�L�񹣩4L}	ͺ�Ԟ�:�����f��ó-����c����%5����?�$}�򒎼
p�+�TC�'���k�l���<ǔRj��ɲ�5Z'N<1%��K1�P� "(+!�2���f#��bap2��-���6�*WM��3T�0C�Xh�����HHu'`$O�d�dE�(��3/)���F)��=�K���yH&���;��n)��auU�Ӭ��+���J���1;�(,ZL�a�L�L��Yųc�� �dUX���u����j�)I��J�]��2:��f�UX�g��N�i;������i��iq�����+:ۙy$禓C��4���@k�US��W��f�:AT�6f��ZXC��"� �rEY�f��,��33/�ռ61�2~e0# ��>=}H�U�{�S��qJ��ŋU�$��b1��Tl�b��i?�Z%9�"�]2��$Y�^���%e;/�����%���ԧ[�U�@�����и���ҥ��-b�]�f�2��I���.Y�����M������E��(��l����A��hI*����	�MlH����=�j,�d�#;��ç�y�,��}�'�����N�]�<ˉQf��`���
h¹歯e[:�=t�O[n@�A �8XF�� �O�y�,'|�&�e�\aW�S(o��L�DĲvh����Ѱ~��xU`'v�As���BTlR��<�����?�O�P���d�c׽��X쒎Y�?}d߃���;O�(��0�{��l�D���zه�Ê/�e�H�Lk��o�
t]�.CM�� �/f�!�Xz�ه�	��N��_!;LR��g���"�=edE�4��̈yſ�=i�y-nOgHT$���{QN�����Q�>J��ab�̲�Z� TJ�֌���?Jy*v���nBY8��Ճ?�@� ��3�ce�u�c|�+��m�P�U٢-1���m��8�Xj��J�ID@u�c�}_��R����X�� �c޾+�Wz�kH�Z������U�y�~ر�]��k�Umh���sJ�+�
��K�-�Ė��r�� Zp�?娙��M��_����n'�*�^�+�2]�#K#B�˘�6�\�o�U�@���=|���h'�D%��B9Α���2�Ny8N�fT�Ȝ�������f�AV�dK7��9Vn�	�������C�d�;&d�P��cO�x�%��G�3�*�uV/�8���L�+�-��jZB�\/�=�����: W�h*Ŗ��|���s�ņ��i��*�/QM��(C-�K�h�Y/��'LT������5�deͤ�چK�[3�l�� �����V���?�W�C��!¦d�� �Iw��QrHR9���rHKH*:�Q1.����1S$��n��,	̞�����?d�kZI*]������{"G�d������"-rߋI�������Hn�x]�
��?�:H6�2J��0�,�վBd���W	u�@d
@g;�4�d�Jd/�hd >~��wz)�
3(��=!Ϣ��W��z��1/����oNt�{��l�%�2���CY��f���~T�MNr-³��zk������ߕ���}*Y]J��F;ހȀV=n���<�4�}*��GV��RW̜�ڡ�Q�9:�͙�	Ydƭ4�ZT=yv�l�s�'�쑗��E���^L�Qw����] L#QF���?��o�E�J��Z��3PG���||�\��~�𤌷�c����������ͱ 1˄#O�<1�>,mpBʶ���r@�ؿ�[EԌn��N�jlʑ��_�R��Ybx5ϑ��R��xm򷗯��GYCNy���L6��PC̙�������� ���*	���i��r�^��eJ�3�c�r���<��`��1+-���'����ȹbSs��njNX]ֿo��n�kN j�ٽ4���j��-�����>1E�����<{]{�X���3��)���\��m����-�ޚy'] �Ʀ8���>��{\�AU�#���S1ڸ�R|�#vi2��tO��ƚ`�����c�9�u
s����C<ÁA5w�C.�`K�D��������0g��^�����e�53	k���ƑArL/���?�Ⱙ���^�D�|�SE�9���?=�/_'�:(y��A�s���b5el�������t�US�qPzv�y�-�3 Ld� �Q�dE�LĞiq �R�N�Z ����Ύ9,��y�Z<>W�k��[�jO��Ug�$�޵3�s�"��}/)��ݒ=�=�-P���T楺��+�B�W&�Ef�P�ZV��.	�w5an��P&7�{��L�� �=�"�H��~�ʌ��D_��L ����C���z0�j;�"'cb8����O���%$G`;]L��9CG�3̑�+&�����0Fc����u 5g�}	�U{���Nͳ�Af+�A���h�%NP9G�X���ub�d�κ�VNH�BL�bP�؍,�j
�EXY��Z�ʺvJ���=�)︣,�����ꨡ�d��dEPQ5�%�y!��b�CF����amB�Ll<�-s)k ����f���|����P`�h�Ԃ�'a��|*we[��}�Gv� ��4���s��b�Q�+��^���k��~�,��%@p��2n&Nh����7�W�܏����r0&J ��$��$�~���=�a+��Ϣ6�$�U�Q�&��-m�:t/��v)�&[t2�iOU���L�S~��t�Y=.�����z�m�IP6��T����>/���{��Q���0Ԣj�4�M
�Z^��1�m5��U��$"��yV�Fq�X@�+V|Q-F%��:����-܎g�QRڨ���e�ɂ�1��d��d(ҐO���2�{����k�:k�PK)��%�o�ɏ���A�©Jd��	�Cd$�-8.���5\fn�I���l�i��&	 X�����ʯ�h��u�6x���L�J�׾���cx�ɫOI��4���J���D'Yl���*f8�I�X�)9�R[���5�f��H�-	��d�G��������������q��)�v���0��`Wc�8�M�1�H�t<D��G���:��/E5"�]�%c?�%4jH�����S~����0m��1l�F�2�Bɣ�`|?�v!�ؙ���=za�e\T�|js}���(���
LW�+0m���P��G��:Q��*�7ٷ�O��B�3��f�R�AN�
�f�3�
]�p~}���*����c~�ۄ�k�JyG��Jc�������_�E�mDZ���:dl�-�u%;���yl� G_�&y�1���+eՏ"99twhpIQv���?��H�M" N�RƴOHш|��L��u-R�:��K�rо�^iO)���v�ݎ+�¤${=E�8��|�3Z%w��WU#�!:^�tx-�Uf��h6��A>�Ƽ�t�e��FX�G9�*�|���3����#�2`�����>C�~ݥ#X�fґ���L39eБ-M�4Ц0���ٌ=��go������f��{T��%�v��V'宿�91؟3oU(���y/,i�����"�E�{�ؿP>gD5.���@O9� Dx��)��	j���՟���Ǚ%"-��;"Q����{�]��=gc#����Q����0&�k�I"^F�L�m� �F�ħ�T�����xԭҳ%��q��'��V?������y����W
�z���5�����(U2�Z1�X��Q�+r���q��S�#R1�!���z%/?�������a�9NQ����{��}���]l���Ӑ�����G�v�K<Ӟm:� E��Q{I8D�{>|Jm7J�5(5�]��D⅗����NA��AT��gSw�~�����_�}Sv�M��W��u�<�}��YL���ߧ�*G1��Tt�R<�s���4z�Z���sLr��XT%�������KO��~~�Ry���
o��x�)!�Ų"�6���q�kS���jտ�4��mGJ!R?"������6����Ӿߩ�*r7���l�:!�5{�b۸	�	�kHN�2&X�2��o?����ǟ�bO�[��!l ;p�M�4%8_�#�Tt��t�2v�0��]�aR��������b��h?���i��ˁ�9�4�@v� ���(eӐG�A�S�o�GX���2x��j���>��\I�^�l1O���T���Hѽcl��!M���WD��=��;�����ʤ���$l�#cy�К��X�T��jw��R� ������vL-76��� Y�'eC�d7��Ē1�9u|�M��׿����)�U%������#wB�Aܶ�)0���s�u������fV�'׸��^�g���U��,)��A���d��\=�)�����]"�9���`dLpi=�Rd�:Ɠ�KdB �"�=*�3 䜁9 �����$5Ř�qAGv��be�F�.��J���ݣ���ҿ��21T��堲C1�esH�1a90���=6a���7���X��c���c��ɎH�X4�G^8n�#�Q�1���D�4������¡^�!ݵ��� {*�C.�b(�;�e�ǥ��Tr:b[^�Y�u϶Pn̲�F�uf�x9����A�f�B��}P�TU������f��*�X��[�3!ލ:mu,�� ���1zEwH=u�v�";X� |����1-2Ј�Us�t���� �WU6Y*3�=	�Y��N8.- |��Lxp*s�3X����0�'u�qv������%�"3�����.N홓�p��Ž�8���`*�D������ ����{Y=8�����M";$��my�0��9�ٷ�A��+`��6��c���cN�Q�m	��F#j�6(	Υ��@����PS5��E`�Yr������y����B�bQ��8��.1�#�s�~�َt`�t+߂�3:eGR�}ll哂�y�qy7FݤZ~eC��<0b�'P�z�:��9,[N�!^V�Px�0���Ub�<�skj��<�m_9l�K׿��D���l���:d�P��F��	{���aV�PΊ��ok�c�R�4&&/%�2O������$l����U*оʶ��v�sF$��,? J��\좴8�?�H������P��Ǐ�x�a�4�o�M�:�Ԍ	���JY��o��k)1�q��j���w`��飏O۱�F�O,}ͥk�������f�qi�-��9�So��&Yg����@��{1\K��vE4��ԳNl��d���f~d;%peU�*�z�aH�ҍ�%5�K��}�Gt�ʃw�=�G�%@�������>}���}�N����w=eu[��Z��5y�G�L2���7���� ��K�S@��b�i�}L��$
�ın|����8�V2 a[��"Ȱ��lvϢk��?�i-^�H�ubˋ{|��4��Z��9����_릕�pt�{�?�:��A�m�MKF�}���M������_��O�N�me��#�n��0d.x�I���=�V�X����TM<�����ۛ���Q+�MAEw΀]��.��_ƪ��"U\=�vh�+W
��PTW�FY�R�b�ˁ������1Ҋ������; ڣdω��� ����d�|L�@Z�V�`UsZ����8zEPyċ�M=���w������Ug뜥�y��qH����_���� fڬ�u�������2%�<� (_|B�U8a�P�*�RtɡP�	��M�O��R�Ez��2�.�$YT�=a��*���EU9.�u��Z�S��t��՟å����4�-N�+ 4A�T�Q�9�)����?m#����	�ߔE�8Ȼ
s��N�t5hQ$u%"nl+�$`�	l�7��<��D~̄���73@�����l�U�'GW�\G�DŦ�cY����\5*: ���,5&��E��.*� w��W��j<^:ZTm�?����P��P�0M(v~l��v�l��S{݁����c��o��9[��>�K�/�E��R,��o���e����lqvl���1��
%�@����vn3�q����M�s���FP�R�_�}s`��AcO&78��jf,3gۿ�z�]�$��=��	��e\dt<�qOo)�����I'W:�����,��z���X]$Ri#&�"��k����/ {9L�����*�����:iy-Jr��H�"%7G,�Ge��<T�������ڒ�)!g�_�6Uy����������P�[��	c�� �*���I�\�j`Q�}T�ql����QJ���u��K�c�]�N9�󇷴/{ߑ�x�$�������li�(�����Y�!g��J��(���c�v�%�	n#���]H؆Γn˒4	���P��=x$�`g�.4|�	a)α�U�<����Y�4��;�Z������L�l��~���P�1UfsF5abՀп;���m@$s`�	�j_=�J����,����̡�|5O��˸0�hQݟ�ڒ٦T�'?���I��N ��,=��z]�P�����_e3L�,����y���M����y�xl�L�&:6s�=ۨ釖i3c����j1DRm�v�P/�_��e�d7oDR��*�߂�lP��t�|��$ 0+���1���{�&R� �S��>:�S�VR��j.[B���$�����i�b�G������f,5��LptE$<�̜G1�8�d�!�e����?���v4�ȋ:'F[�Uǝj�ڠ�Э���B��q�50�fe���Z}�qo ��R�,�(;��qc�nF��0��{v�ו5T��&�F�#�b��QRF/������9�!C���R����*޴��"P�iU;ٍ�h)4%	��N<�K�-���
p{��&�8/F��x=�"��
S-ԓ�y�ԯ�U�Ϛ{�ۗ���y�>N���[,��b�n�yE�t�	��8��gב,�j�����q�R>T,+��S�T@�>}|N�������((��������%�$����7ǘ�E�L��2�^�.��}�����s,vpT�Em`I�Bglɖ%��4�C��2y�&�컇Fo&¥^yC�Qٮ0�A���3�)ոU�f�+c[#��;�;�j�\4}���,���ֹ�ktC�<��H`<:SA��Rd ��T㱣��=�rr6#'��呂�RN��J��oU�B 	�;lT�/��lҲ�[��7h�O�jB���/)�ʩ�~ߛ66z���?c��!�4��bs���L!)U��8�(%ff��+WҸ���)�NX���[s�a����{��T�����1%���=n���Z�u�1� |Щu�#&ApN(�,^�c�t[�N~���'�?�`��;� �a�W�`�࠲�N���R���`�Ps	�$���( �@Y!�j�@��8�8CV2�uE}��]k��w�z�ꍗ��s��E���I�g;����k�x@�N20I�Х��F� ����j�]3�ǔ�u�2N�-�*%c�E�(��N0������K��Ǥ��\}7���똳~�E3j����VS�DE@�͡_Y�A�����%�hҝA�3����ޝ��u
pq�A&u7�ѳ��Z�5���f�� ��,��64��1G�CA�EYZ?y�f�2.6�<�!�R�W 5��mt;�\��y�I81^�;
���d�������������o/_$�>'ya�AR��X���3�0���_���!�zZ��6{
T�$��q��sA������s������9SU�ζ�.�0l�v��QY ��R���)	��|���f�ޛ�=�qR�2��2d�D*��9IW>�_e a`��b�8%��0U���j�27u$B�N:@��KamA�8��� t����ΣI��Q�33m��q����Ef�&�,�n71Tsfg�ΐ�TS�� 3���}�WLJ�2��ƚT;8j⑤m�K��z?Y6ʝ��&0T��q_�[+�ـW�]���I��8Σ&_э�ƜC;��l�)��Nѣ�s���՜RF
���C�(�� /_�������~�"u����矶�N���=H���t?b������f��=f�����#y'[���x#UB@>���:�}`j)��z��+,ԅ�}g��A3p!*w��;Z|���'�Q�R���b��� 9[�,d,o5���d�0#UK��{#|�w%M�� ����w��A`�Ksp`rR����ź�&� V�	qF8>d�c~r��Y�����)ۤh F�[B�z�4	s�H�����|�&i#�g��5�.b=����a��+�T;+�~g
}���*�,�V�t��rOp{�w	ˣ=
������Wh-2�Kj���/ʀV�y�;ԏ�^ڝsb(��f�Pb�2¯$�`4�����k7ה�{�ͳ������AC7(	m1+k���KJ�N,�ö϶v���d
�͂�}�/T�&�B<�/��Q}P�1�����)���4�ai�S�p��Y�6�B����NR r��,f��A�7VU�V�%�X�.xyXǦ+G���b�z� �;{v��y�yx�Zʉct{��d3�/'��&F�YV8JF�:��j�33Q��<I�mu;�nj�w��5�8`�hQr(�A��=]o1��4]V[�r�ɻX�M&����7���.���m�x'������P6;j+Ʀ����A��J)Y��k�h�!y^o���H���Q��0'ڗh���!ܯ��f?��,��$ ~�����k�����1T��vu�*��U�-���,�-��
��\Z��J�s���j���F����N���t�\�|��l[՜�#�&[dB�K&��t�ۅ�~�% �A6�T���	�k�w�B�l�NV�F � }��z[�"���V*9u�^ى66kK<��vz�2�֑m�;�n����W��1!@��N��h��1GD�h��H���ʾ4���Xof�\�M<
!hsxxȘ0��)�F�/b�|��xZ��i�i��q0�ds:*Sۅ�d�4A{6��y�d`@�]Vf&$d&�&���S*�bdA��ٽ�E�1�H9���x0ٱiL��\��W�)0=`,�*���e˦���&��J㤭L4)%�ޮLEs��L����CM)����N���~$�yg�Z������"k���B���U�QUS�R����N���Y���^�`e��\�]ڕ����7���Ւ:�����bL&t�R�d�xL�(��9��M�������ó՛�<����҄��r��ng�s������?���Q\R�{����*��h�U�l ˙�leö��cl}�����p؛m0��\�$�݇�w�B_�@��2��_`��EPUe]{�������$�b:hRO�3Ϯ��]!���u�
N�X,�i	al��JE�w�I_�F������qp��ɪ!@�X9e5�V�_-X��~c6f��l-� �u�*yP{(���)�}�Cm�ooY�Ý������1�7��Ī%\_�y-�f��-F4TV�h��K\wb��A@��t9��z���A�u|���~�CπÁl���*����o�W������z;��$�(��&�'�� ���������:��(�`!�<��j�x�M�O|���MP�RRU���	�'�,�a�i����.:����̪ሔs��V���Ȓ��v��M��r��qe�	�~ gL�0	`���NV8�E��s����Q���R�o�����#��q����@\��*L�1������y4��h�1��ץ%����&X�6V�G��0�4�\E�6�Paf*O��`3`BJ�Q7��9{�\#*�1��:x�Cfs��B�^N���JܸL�ZJ�܏������������O�>3���tK���?뻒�8:�M����k5mڠ^tN�ۃ��w n8�}'՝��S*�>�頵�i�C5��BFNu�$ӝ�ERf2PN[�=,��L�ň� P��I�(w��*�J�#{�]�L*`�����n ��������͓�R����We����NMtoPǉy����n����+p�j?@tIo���OO��?�i�/`��C�f�xW��puZ���Rߝ�C��O�>�q��J���!��cB����>�c"����R4�u��H��dc�ը��(7�@$�e�q"�ŉ��
��^4 02�+��j ��E�]��"��WU{Դ~�(����u�.� 2cr	��^㬔�s���^VI�B*���GY��C��� `o*����ͬA� c�8U�.}����ExG�����{�,;�(��� �/1<����1�D��$�0����nW�e�w��F�3Q�;�:�d�+x!Ѩ�3*�|����JVJ�ڊx�Mu���\�Q��w�wN����[�yX���V��'c1��OV�$Tw{]���hx�/}yǎD������J╖�9��Avr`mb�z'8j+���yO�j�f�Q�.bvJ��.q����<��.h��v�m�)�=��%Y ?L�����7�6���9i<�F0T؝6x����\�����eae!���[�U������,A�R�A�����<�I�$��=옝`�)�S���!@��!{�NS�A�#֙[��9�i���Фo�X�\���&�0��<�e����SPM�:��!�%�'XL�̳X���eo�;o�B�w�4j�\!���*?�{�!h�yb�"Il���f�p�Mw����'c�X�@B��:Fٳ���b��	K�x�M�z�s�5LLm���d�c�2�@N��������Z&��Xm����4�������c&��4�A���S;ӷWJ���T'�S�~���~�>�L׉������;�.v�	x>bZ&�`z�p�^C���{4��9�3��%l��tJ>	h�G��-���P!2T�5ɋX�p,:����q�˟����ܻU��Tb&��aVʁ���-�غ��}n�܆u-�o&|N�Pe����_�:L�*
�0u5y2ah%���YR3CHꗝ�0iu��k���Z�������NUttDs\(�����Q���Gw>)��tŠ�P�ua�"7�����n<R��pLX����H���!�v{zy2���ާg���v�1/0�\��1,�����>'Th�+X}��rzi'\���%@�G���ᅳ�w�ٙ��M7Y&��F��!L*�Q���E�x��%��1sb�����o�ٳ/��+��1���w
	�2v�'�bS	�L?��_$��Q�O|{��&"[�\0�gj��mD؆6��@u[$�:��*U_��>�C0~�0+���d ��ql�c�] z��(h�[�����p��Zfz.K*ȗ�E�o)���kc�̓*`u�^TF�a=�m)(�0v{�m5�����X^�i��\r�X��Pl��5z�FR�(͚��a�e�4�D
�X�u&�*[OcQEvw���R���*�Wʫmu8*�p5Yx\ՅU4������j7E��,\f�m�����8�`we����*o��	ɇG�+S�e�ϲ�A��;[8���#�<�l��}WTYgB%���ʮ��ۇ���E��S��Xꓪ��d�$����H$.[��LrŲ�1�Cx'yg6�M��<������Eˑ�M�Ꝟsz����LuUe�K�	\��F�Kr)2�&�顗��ˋ�6T:hA��,v�i���l�W�V�!`Es��բ>�>��U��q��~x)I\~�^�����W���$���������(`�!*0��t_z�F���P��*v<ƚt���ύ�Qj�\j�U�V�E���r
&Et`��A�ׯ�w_D�� �����]���V[k&����׶S��W3�����C����b �, |���&hӻ�JE$��D�.n��á���^�Mۢ�{_}߮�,o]$>��\���XFO�$N���;��T�5P���!K%�w,�}����.E�T�Q7�-��0�	0���(�cˬ��ܫ�� �{�۽����-�Y��(ʊ[^��?��u����z[��d��o�?�����xK?
�1�f�͞���3��t��s��:Y�SË�bK�I̅�omѦ�OLC�g��@��G���*�Z��
�$��ׂ��\�ye�n���8cz]z�Q*���oZi�m��b�VX��hv�B���G!���8�*+kP�*mԊm���>�9;k�Cǘ�r<S�2Qy��Dy�����Ō�n��f���[��|���f�ySd.).� �]�Iy�n��V��:�Vs좛n�h�;�:�U��1�2� �2ෳ�4r������W��s��������_�>�/M"��F8�YQ�}��D.�A��yI.B��L�DO�����/��e�ì�
$oj�kƘ��ݷs��7 k��C�Y�5�k���������{<���}L������1���H=Η{�`����^�溄@�I�ԞS���'趿���_��}ۀ�`�Zl�Svc�"�{������'.p�N�������?{0�w�C�]0���TU�WXkD�oi)��Di������l���p ��A5\��Ď*'_�8����-l��� kd�W3_�Ѿ���]M�t/�� х@�#U����;D��-���תbaԠjE4�_-��ڤ�Z(���I��Q7κi�_s{WV�����!ت�4�ݒZMao�сB����dn_o�5�ec@G�X*���W~�!���¤�b0)�E� �c��-�E��-bBT�;�zO��ئxZ|1�I}ׁmᴅG�N}g܁�1��R#�h�֬�}=D�9ۥ�r���Ȧ3��-��r��>�>Nh�|g϶Tc���7�3=�Ǐww����곩�>m��Ǉ�Kw�i}��/��C���-X�������8��|Dt��.bg5D6��0�a������j �C�5*|�U�hư��@ǯC/?A1�NVו�l�۸��@�	��v@o�>���z�#�h؟;�X��<n�R4¦��\�4zE6�X`wONO�C-�T�.����+[Kn�葀���a. �?.+r;�£M��s�6?�7��?���2y�8�h�PN�����~��;���5��o=����$zvK]4<cV����܍	�����ݣ��7��؊?׏;�T�<�+O�H_���P�m�t�����G�4��y�O�hL'��}���ؤj�g���� �j�������o�0��K+E��()��\J�l�z'buv�&��%;9��P�|w�~�
�gX�kO9bc���&$Tؘ �3`G.��Y����{E�]�r����(�nUjA�EN�����l��xV�Ab�ڱ�؜ D�9��.���hgĩ>aq�,��n�h��"$fWU�i,��i�����v�����LSE�25I�IiP�9�Ѿ��cXy�~P�LW[�����U#��Y0�-o����I��M��9u�Rwq���Aqtz�S���^���~�t� �f�����o�âA��/A,��@ X������[�O�#ߋ^h���!JPY|�u��I�p��v��w=D�P�Sam0S��:��� tV���c�a����y*[�]�Wz�x�k7	��,bݺN{`O(��w{�8�CL�0��đ���'	���F���Ί���� f@��8���b�����E��ܙ6��(��I�;��� <�A��`#��ۍk�����E�P�׹����`/���cJ�YHe�,q��[�� �S�H�C/.�믺�y�ަ!]��'1�'���?����V=H��(@͕E������Kwo��XY���������X��PW�׮;$W��m��k�p�rk��L�<�n��V�J��%On[ӻ+
���9�U>��&�����\fڤ��?�r��co���-�����
\�U 8�;X�_Ƒ��a��x�W� �6�Mp�y=(N3}��@��7᪤ u��n����0��@�:>��g��i�����`�6Z���;U��`L>�Y���f��>���;;՘`��!���$dE\�!�F�
5��y��{{`|%�']��є {�v������~��q«�dz�3$Q#&|����h!�>�R3x9	�^��������-�EÇ�B��~��?��H���DTl��*��֏�z}�}�_��v�=`.�Tw�J�������f���TYK��b �Il�Y� ��D������"S!v�Y-qZjx��cA�������+y6	q�@���<��J���� ��L��o� 7��ǪC�E�;�}������Ǉ�?p]V�4Lr� F����>�%^oX�=�O�b.A��%�����*����	�>��>���TVK �	`H+���ߋ�ḿv�b�(���`���1"E�EcC��WI͌�`�k��>�$�%WS�U;7N��m1�n�����|i��UC�#��"�P�T���'�P!��+�}���\�P�ӛ��4B]�a�|
u/���~wG�Գt��n7vɍ��vV�}�j��9;���H���V���`��;\Õ�>k�E"fc�X����s�Pȳ0���S_xZ�ب�q/�m�I҃+Wl/.�Zݡ�'����I�l�����w���C|ףE�B��RL��[�h�X�B%��j|�u���I�Ll[L��5Q�M�a'՜s������~��AAsMU��<S�;�o'	k�TY-���8����G����`�Y���[��y��d�T�*ޞ����}�86�o
��oO�J�%��և���e��S�1�b��|���e@e�Wb��ȹ[_�p�����зF�hfb�G�]�13������Of�<�y��p������x����H����Gq�"��`����!�ɂɪ�d;� ����6��Jk��x��^�J�ar#h���ޞ����:�ሢ�5X q3�3̓V˅N/�W[���! 5T-���3�f��y�������Y?̪�P	d�K��_��C(��
�y�2F�i|��V�]�� ��Q�v���$7 ZhqO��a�G�Xz�h��VWp���U�dK�V	�����/�PID[��\-a�{�P�������ZK�1���>}/���H> ��{'l����8���齎�QE d�\ݍ
b:�;3�m�GE���lZ������!+�Ws�)�x���� ����Z=_��7)� غ>�ʈC�����>��:��ipUgdX�Eub�i� �l2$�%�?"���I��D7�����F}]��U��AG
�dwrU*/�Ok*���O��"0>;����%��C�Z��8_�;�VooR	�L����YK��e`���u�R�#\G�4�$�֧L(��V4T�����o1�r0K?��M��ڇ�����k_�j�\��j���6xK�+���Rxϓ���k�#i���zݎ��8D�/���D �㮂]�hG<#���vu �>���>km�6'n��օ`�3��.��� <���t�.���̂��ֶ(�
_t����n�Y�����G;D����+�����.R\ꓕ��!
C�Nn��X���;C���.C���J 1H�.�T�!�B�%��/D��#���S֎�!�5ư������G����6ͅ�G*�JuE����yV�3�lL���yتGP�7â2 k���p�_�.8���q�E�DMy�F���������I�hر7E��C !H���#������JFB= ���#tǙ�3) 6����)��+1Q�* ��룉���}.�������\0��3�DVWD#�("��g�@��Ǥl~�R����}�޾k����U~{�X�烖�Er�	�b̩?>����걌�ǌe.Ĩj���]�.rb ������`uCS��l����]���,Us����?Ę�
� ��p�	[�ĺ�����=^d�����H�v)�$��g,���bn8KvTgUE���B���T�%"��V��6-�����`�n4��`���������~ś"�V�B 1��ƢZ��~��լ�(��8�����u;�o�h��zt��;�a�B;��	c���^���]۽}��:�7�ɶ����b����������\|�������S�SϔB	]�h"sQ��V������)��U��af��14��V����zF�djup?��Ǎ��}�A�T��F��c�����o��8��ߏ�q�\+��c��8�Tlw�i���-
̠H���Hݒ����P[/��5��ky�y�k��`�`Ǉp.�F�f��Ik�笈�f� -?�:q�Q�4�	�z�������)� �5	�p�d>������Z
����oؘ"��.�s�['�:h�>�;�Hp�5u0�0�-(�tW�+I��k��V#���`@���%�����OR��Xq�H�y��,��k���m	�Gx�4V�����G��ߡ��|l�EW��a��X�3�l^k/4~^���Խ����}�P�j���"g��9U}��±��7�^�)�����z�v�x@]�|����&�9D7%�ے��.~�Ŋ�K".j��վq�Qe�zy�\1��$�J��QMITNP½�(��}����9Vw ������/�E23��r��}�)��' &xx����˖0O�0%�:]Pt�V�0�j��<�6��U7 �N�Y�vfr�v��=��w��/�׌m�Ϲ/{�1A*�%\W7�3�N}�������� 3�������s*{�m�=�~�M���ރ`��2�!����f���{����
6�:��W��Y�K�lE<jw�*��d�˥f��m�/:��s��`<C_��'4�x0��r=Q13b(FlNZu��l�e�G	��%�Yd|ݥ����T!��o�
� R�a�nea;�������}]�ܚqRu`���MNr�0oK
�A$�q�;���q�vҧW�	�k�o�?O��9����}�@��S��?��+�a��iy��2���mLF�h��:�l��d�̭�]�Tzn,V]�o���.&� �1N�?h�J@���R�O腗7�]����'�-���0Ԧ��mˋ3Fkao�PYT$$OH��g�u	�Q��z��t���<��=��<zp���Ax����",��V~,$1Y���䖡4�܍#8���/:�ɬPɀXÌ5�S�{g��;J�k�P~8ɻ�i�}�7���+�tk�#,�o{l������f�µPa@tW�V�=Z��������>O(ގ;nę0@b�*��J��J!0�����U_l�d�Q�ЇE���F�<.T��l�O$
�-�>�0	�,�S�: �x��|ϙ�K,�p�y⏢� �[	�25���3�w����Ў\��:�A$K`���ӭ��ĪC (vP߮۶.U��T��]��ZCʩ�5�(3�Y�Ҷ1�|���o��փ|X�W�zQ��	b�N���m�3��%���Ok��vY\ų�	�hz.���"�* 
�`L��i����ܛ&�#�Y�*$��!�B<+.��{18���@��+��0�l�@�T�Q��V����E<X��ַ�A����T��%�qh���4�Ԡ� �I�|-��"4�+IC�!'R~��1P9A֏}.�F��<�D�ѼP}��ΰX�����Ņ��x*\:�E��.�7퓾ǘPi,38�� d`���� ՚�Gu`gx�\�0{1^�ġ���5Z|�Ƿ�b��;��}łG�!�E)q���Q��m�^#)2F��A��D)汪���D�����i)����6�p�q�٠�t?�B֬�	���5;��5����J�-���h~�,����aA�8�R��X�� �� �{יZ$��rġ��G'j��8d�$��N�-X	Vt{ �'O��4`.
I9�t��`5�'�08�|)C�@�#���Y�5�8>&f�j��M���{dt�v{=���᫕�� �"G�q�ya�sKn�`����й� [��]H�j�U��>V���O�,{�-�?�Z����2'�"���y�}d**3zAE�-�8"��ٺJ�L+�z߷����j����I�����?��s�S��ęB�ZEk�5�����K�����"	�����$ʹ�AG�`b��vN; ې$�� T��>�u���n��GA��cwn~�#6�@�6�����c�fL�$}J�ݧ1H�%��?#��3�h��Ǧ�.ś2��}�4b+��	��L>b	ΰ�w% "�+~�nY=��xc��Bg�5������}A�F?pm�z$�H�*�V; ��7���X<�`�c�:��̀��8h�|Z]Gݞۂ��z?��>M]cio1����7� ޑ�`h����z���������	������Wz;�%�ϵ7M4AD"՝J��gⲅA31�`
�s!���*��h�I]?�s%��n�����	1&`6��������OAU�� '����>l�4���7��F�;�b6C�$�/��XUa5
��nA.؄U�M��M��{u��}i w�p�*�W�Mf�����x,�NF[�j��/H�J��blr���c�W�r�lA^`H,I��;����g�`@�6�=x8��%�����?hއ�ю��[�A~���ނ�g8�+��<6��1�}��ڽR�zWZ@v|�/Hϋ�����h�����@�{w�z�ɫ�"�b��}nZ4R\40�X�[��� ��Ĺal��t�o@�"���|�(��￙��w*���n�(O.���&d��E۾:0g�K-������o ����ʶj�g��	�W` ��{�VP/�)����k�@'��6��͠��ݵ�2�.ݰ�sF���ĤЗi,I�����^��	�]��D���\�����0CB�5�>t������������w�����P[jQ�~t��U����HX9���5��O�U��ܫj!R�m���_���Y�A�}�#$�_{vz��o�铵h���[�s'b�3s�@�+�r H����F�x��a4_�f&R_� �$��eI]�N����gu���Q �;�[t�ys�Q����m��UX� cj �bn7�l�N`�\i�;�	�?k��	AY�a�'Fu6��$���U�,�{t��7Z�3��C�z�Σ����MG�E�W���!uIwG�%�=���3�&��8����,� � Q;������_�%ʚa�D!%�+�����K�#��y��;R%��Jǘ,i�p�P��c3۩����4���:ܚ�t�&�Y*�Y�D�����_U�).^AI�IƤ ,6�t��4p�m���s2�7�!�z����:�%��^צ�׈�łI�B�j�����A��O���Ҋ,9/Tp�P���۠$0�B�� MN�9�=�P�� �x��E��_ �D��~��]����u`o��4- 6QK��
�o*l�;��@oOuPJ~�AH��\δ%@��T0��^.�W�?�[�k�]p*��8�磇d�I�)[�gv�ʅ{�/i69�8(����53X��%�f����G�ʂ�>"|)=ű�w�+�6�ۅ�_�Eu�Q��]^HU��+T�0p"���&U�y���ǡ�q=��-P9h, S�X9ҹN�X��hQb_v�	�'���8�ؿ�����+B$*���7���@}#���>�uq@ų���%�]ז]2oO�e�b�P�]H��@��
���e��l�bS~�h�V�D_��$�������6�zl[�]�#��#�S�1��ƛ��{��Y�П�T�?�},��$	��D���3Jބ���� H��9!Pe)a�S_c����U�� ?�%9�������L��z̃��"qR�7�� ����ų~��[k�;�7�$L�5�_�>�ˡ΃T���ثN�~��܎�]J�˂8��v�� H��?��}�-o���	P��3�ˑe�
H�+���b`�D���UN#�EC��!H�u7�i��CeH�S(Sv�Ie_{��.��DT8ދ����a�V���5���j�ij^���t�K�P*�Yy�Zf#�P�U+_��^�J������Q~1&��G�+"��q�9Viq0MD����"�)1X�(�_�w��R_M�U�p����G1eh)���EP�(߮�X)�� ����k����"X��w{69�қ���� TI�Z�����LBWh�#��[	�W|[a_I��"�r\-�m\6����s�c�⣘�$3D��ϓ��l�e&Џ��bt��:�J�I`�b� �$Rs�� �]:Ԡ���h'n3Jc�c��T>a-� �j���?���X�.��J���QH��*����)��2/e�.z�zҧ;SĽ�v*Y�,�hHW*�)aH���4�a��#e�Un3�K���H<��l\��7�X��RWou<�5�&=�ʯ�8:Xㅶ��蓣�v�¢�c���د��:�/ ���_.�����^[�.���H�����)��E@]T��8���U�/VP����-�H����{nT�E��#����X��87'V]R�@�\5Q��EӋ���.-BVMu�q��t�"Ĝ�xi�>
|�K����/�^� J�|�J�?�K�\��:b������m�V�^�0X��]��O9���Z��������[  C	c�=�Y���Xd�G���D�:���`�m�i�)���/ޏ>N�=[�Ꮛv�;��%-~ǒ�KS~��A�ϗ#� 5Z�t6�ăl�/�06M^��O�C]ݛ�Q$�|8.�ǭ%��p���~��߿}����x ۶翉�o���?4pt�k�8��M��s�h�]f�E�Eu]��/�5�����)O��k��c/?�������j�҂�T>"��>{a�|�:0�!��|oL�>X������a��7��5�耶�i�#��POtvO��� Ф{+�A�=�(�t���ڣn���m���#�k�\�8��ڮ$�NB+�H+��E���mQ���ΔR�J�;��w����}�N��k\�(��f������%vi��Tw�|g�Xf 5*�@��� ŉ�K�qn�Sn���D�m!�9��	p��Ѥ�零�@CU���i}���)��Z�e	&�
}���Smt��}RP��\�f�G��o�Ӣ:����������-��������K������aˢHi�j�D%��o����h;=�crK���¹��w�bʢ��Zg������k��nVk�^��:�`h�/EWu��^Q���gU%]���I�+~���&'�H/��	��@Ww@���V�O
)�b=F�S��=HЗ��l �-�2B׌^��b�ZeuF�$���`l/���3�+x��i�X��&jEY�bۚ�3:�Nxa�}K���A�2�;��b����y�J���ZZ�!<���g�*ķk�'���.��W�<n�V���x4×���F[l��p ��t�GڱU���}��{�]��o?�������-`��q�����v²���_I�s��+�� ��+#�c�6�~o~o��Z�~��3��R;�u���oyk����~���wN���D;�mK-gLg���|���uu�9��²'n�eS��+�)�uJ-b�y����F�A7�k�?�U@&B�zা�O$��#�Rl�.`:�F�?��R�n��W�� A�*�b,9(���l�[rc|�4����,z����Hb�h,�z�E\+�b2�S�s�X��mYT��ߦ~�0��
�<�Yz3bd�_8 ݩ:P_g?-ݕ	Ǚ��;���n_�������۷��Y�{8Ϳtv|�f�&�z_��{W��~zE}�.
'ł�=��寉
}�p���6��e��R=��ǇdP�7�H��	WJ�8�.����3�%"�KLxl�[��-B��u��d���b 
�()��m��E����0��/p��8A��v��).GL������d�E�����n@�NU �!��U:`[�.��X�q��y�O�~/4v��?�o�r�;�R�[?�,�Qɤ�E�Ƀ�|b�q��s4$��V DǢ9l�����i�mE���������?�*����� W���<�) B�-�����m�<���.m��B��]<F��ȃ�3�nI��W��*09�1����ZW����5&��70$��{�'0�:�2_���mP������wka! ��y�R�Ws��?��#@�i�)�>zsLTepY����c���P)����DF�+w� �H��B�������x�Lԧ/�o�L�M�u[��u����%ܕ�~$��b]}k�o�F�.��q��޽>���ɵ��/i7��xU,^_�UcwԼU�I�_�r�3�MY� ��.䤺E��6����R"~�����31�mzV��\Yg� �,����0��7�,Vg��E%0M�0|�Lv Tχ�1On����B�3�c�S�|��~x�3\m�f�����?�1�eX���Y�ci�ɠ�мP�πu�s����f�b�D��1b���Y�Q�F�rP����(?m߄���-X�o.ry���bb�8� ���TØ��� u�x� W�~���/�P�ԃ��Uw�!��t�b�8���`��]�C��H4m�+@l��t%B}�L�'�[[a����Vl�Q�gF"08�9e���6��/&�����;Y�oMi���G�8*S�ig�:��d����`��%K�Mi>{	bjy=q�ŇA} �Gq����d �1��Ԕߔ�G~5VJ߃�IM���	��;�S��>=br�&m��*�D_�۰ÑG���9W;�OF�9�,�_P���:�=���ʋM�Â�VG���-�E��R�Ɇ|�c�{��yW��~!=�[/�;V���x������#���Џʅ?��wt��J��z�э3����'��/���l�u��u%�=$1����������,j��$XӹV���}�Tk�_䏒�t�q�l�.���d��Œ�����g�_�Om�{��F.(�"Hw�2��C��HS�	-��� W�1 ��ʈ�/����C�Db�Ī� cL�#s�؉�%5�I* �?�u��/�d9�v4�L,Ę(�#��Kw�  �3��w��f���S�*{�	uU7&j̹PE�n�j^9��S1�P�i�gg�ߪ��#�P'���r`�Yj��n��۬%]��d\�ga.T�=#j^p�9=��}u�b�iL-�w�)�MU�-������Q3<w�Zb�B����"�]]~�0�FI��{��$��b'y�~�r��C=���@�,2b`X�1�R�6%��P]�6�<�apls��.iE�j���mn�����Ǿ���<Q��ҐUf���rK ��59C�q,N&'�]�%�]<�)�M6��@��3������0#�����(j��TV>3
Z�p�]�`9�!_�X��NO5D�*��I�,��H�Jeem+/!х����h�
܍(�����N�p%��ׯ�䤻���z���!^��&�@�*�AZE�҇II��Vol�m�μ�G�bu��v��MD=�^���ֱ�l�Lrη%��h�c�F���ӱ��An����z��~��8�f>��d�0&�6UI3���"�]�nKeLj��3m媥��M�'dv�����2bu���M������-�jӈ�ZH,���O����V��C���J�����~ʰt�\���wL5�n6���h�2����ܦ�����?x��"{��q�l[��oM����c9�L�K��R�~��q]�*
E<�.C�fe`R�;g^��>HaͿ?-���=R	mVF���tcƨ0��W����z�޸L:AM^�����8l��m[�:f���2��Է�����?.�5�+Z���#`<1�З��~�4Z��j�L���T�N}(y��3�<�+y tݩ�~Js]J�Sy��+�s*ړ�+>Wd@Ex0X�\�SU�o�����C�U�P4��Y��E]5�"��^ީD�Ds6k^���n��*��������I\B��l:�<c���d:A%X�O%ʧ����������y��5ʤ������:i�k	��a9A�ExQ��M���&ou�TmT2,�� u�NE�A��W�F�.n0�q�q���ږ���}���BE;���Ib(�b8�d�*cTf��A����ju VЯw��{���@b��mG�r�3�2-�N�� Zt_�3����l��8������'�
+l�����ʸ����|�#q�0f�j�ʀ`�>�I���������lt���5��|FK�,1�3�#M����GW?�c�u�(!�b�q��\�O��7�. �|��`m�(-��m2uu��&֒��d�ݦ]��x�[�r���!�d� 5���+H(����!G�o�������=z܁掫��=�J��S;�3.���� �k �D�v�@�M�Ѣ���\?Tɦ�n�P��y�(�hNH��EP�\ޭ�Z%��ս��|nN�y�;��]+3�F�������y<��կN>m�lHe���^�[�w��f�5���2�_�^�O�m~�ɽ?���w� =0��e� ��F�"�=���ޒ���?�"��=.5��3����"3LG6�°�\֪��sI��%	���B�}c���Ķ	H�@b�j�'a㙃&���g�@�į�RU�ʋ��c�Zz�c?\�w)�&�9m���,�QJRxO`D����bEj��1��~7�X���59X�WD�������um�˃ߴ^�獍?�/�(A�\��e�����4Q��b�������:�">Wù�o��Z�$K?���R���T@U1J;�96c���%v��8���<!@X�N�*���
��j��X����d�@"�����, u}��6)�)FÛx{ܒ�Z�?ӿj�j�R���ሹ����b0}�&e�B|�<�9l���m�zY*�J�`+U���I��) c�V�`wp% 
��qa+�,!�b��A!.B�:I(W�w;[⤚�x�����J�5�	���O���f}<�,��� ���_;��H��������0�	B��l�̬��PUԍ����" �Lz����*��F'}�<�H����	F�`�Xj.Hܚ�M�U��LavR������DD�F���KQ��J?aT��_h_��ק�y�ݣ�;�<Q�<�$�G�G�����\�]5ɏ�ކ�Bw�d�D�����J^�Jz��/�N]�$�K��i�.)ew2���O��f]���zQ�Ѵ�%��Z������nk\�7�R=�tw��P���$=�F&�'���E��~���!	��d(K�yn%'Iv�d��5>�DV�y�_��������WzSTqDW�*�d���s��8&:V7^���aq<=3P�uE%�LX�q���ș�f�|?�6��nL�n5C��?�\{�s���cy ��0i�C8!x�_/D�H������d�D�����G�0�`�"��8���	���q���:��.�L�)>Y�J�#�B��9��}9�;.�<aL�׏�GP�N���U�J����\$?�}�-����/%�#�r���F�¯!!�My(�a���Na׌��bދ��>3w�	��/���C��R9LJ���}B�G�rx�f���D�i*.�0��k��W"E�Lڞٓ�j]���� �xz����+���l&J%0��A[�{Ĺ�
�^�o<1TV�er��P~�$U��Y���i��YD��F��x{�}z?�<�����*.̾À�s�H�$wmGo�9�PU@u�Ҋ�QA���$��g���֕TN��l���ܓD\JùP��(@��#�g�3��ecI�W���h���Hٵ&D;�]���1v�D�&�T�d�s[hU=�r�����r\]�6N�:9������SPn���3}%݃D�ӡGzɃ�|�/�yT�e�<N!m!%��EL���jX�Š�6���<,�v?3.���S��	���Wz��䭧��ӺY�
~��{��G��5�:�Z��bu�o�Z&�:�H��������H��~���@r /��eEk�0/H���T7�s�6�b�4W�|%="��l6�O��I&z���ޙ��+�ߴ�N3�Oyo���-�����%HN�x8��a!�3�S>A,��zتm�3��u����8-�b%-q�@ ��x؂-�%�eT�>��B"���_Ԓ^�l�Z�骂U
��=&�����΄����󩟘z|��y��P+LAd��n�c%=�����0���g��W�������mK3�T�7���M�=����B;neh�MNCK�e��__�����b�5����6u�qe��t����`��j���@n3>��[�~\�������w��խ�f�iQ��|������`�*%�4b�^f�Y쫓�-9=U�`'�;�8J����I5U���_�Y��7�����Ens�t��K9�� ��6��w�'m����L+;�&���K�ܣ�W?����P��mX�:��է����q<�90�LF�Z�1)��%���smw����Rb���s�;�BP7����T'70��-��i��c���`Љ_��*��� ��_��MJ��1>�X��ۅKW)�p F��@8�@Z�%��V�7�ޗ'7fW��U�U�/ u����NC%�:k�g���J�Y�%uLYG]��ab��/�]qp��� (%2��O�P~WĻ.�B�����*�����Zۏo�R���w��$�\+&Tb,���W&1��>�]-{m�d+ 2<���5��s��N/�۪�p��JƁe�Ku��*L�	e��g��b�U��j��A�6�@���H�'��;�O�&�+�i^=�7�nRF��ܰY��z���mK�g���9�z*#����+�S��]�]uW�<{�W��\٬^�w�n��P�R��T��<qJ�2�yy��B!�ƦP,�� �y�����kl��׆?_�bF+UK,�q\n0����C�u㳩��zF����t��|s� �o�{�R_ ��Tc@x `�}(�_L?��;�(e���2���d�=ꊣ��;(AW�����84��+��_�/c� �.��$�L��*��D�v�t-q����v$���E�U�j���	��&+�@�a� �;�He��A��?s��E���if4�~} ��f[���$4�C��I�z3>-�2ރT�Zbw�$�2wtp�`����W�~Q5�*���:���J�:��ŴםWp�yv�	:T�d��`�
�'�Q8�D�.	<]0�a�� (�C>)�ŵ~[�g��#nK��g�_	\�p(��ԩ�����/`wx~�4�H:���]O{�Ӳ�<�u)��8a���L"3�ug]��r�`����-���o繸D��Bd�G���K܋���u�i���'�fAz�`�\����_�x_h�$���۲�(m���
_���7��U;��d� Z+}Q��A�~a�߄j>�\�s�=�B
)G�l%��I�e*�(-�Ew�r�l����f�:#o���g-�tNP	��j2�����������
������W�Oa���e�5���AwC�yRv�T�[�ѥ�a[����-�H��&Hu(S�{-'��谵���_�U��5���$����t�^���WJ��rw[��e�.���n�a�<�^N ������B.��ns�9c�Fu�6W��JRFT�Ol>�|(�8;�O(kh�}�Ɓ�?+�P��f���#������Wb��M,��]�"ex��������*ݒ�S�>D�a6�(���4{�H�Y����Ϛn���}ˋ�P�+���ϐ������Y�g,ʩ; IJL��{���X�]�s3����a�*�n����WD���p�M���vT����R@�O�L���c�O�ߚ���L�f��o�xe���� P>�	�k��a޻���B��\/�_���K2���4���թ~���pe՘�� JN�0��_T<^��L��8��y�Y�2'.|���UZ�jZ`�� �E��4@�w^Mo"��h +���c��G���u�0���N�qE����Zc ��e;�N�`
���3���t{��-6�|h2��]��� 0�5�=���h���;�1�U�|/�i��5l"wԣ�H-�!΀��W��jӿ���(���&��IN�j� i�7����W$Ҁ�|��Y����V�X�F������[o���\��p:��j�ù�V��ӘK�����	�����!WP�a��Ӆ��+���*��,�>V������������9C�23�$��󀾲͛�L_ڞ�ů��N}^6�����AZ ���ywc�2��n9�|�E�=n�z���,����י����������Y>Z�f\����[���%@�E���4���l������;TP�RO��h��u���i�� )���k%:,O� ξ�cQ�	U�_�~�po=���X�vq��{�ޓ�v�{��k)�i�~Fԭ<�Kͷ<��~�dZA	�Qe���zl����v�̘�_��� 'X���E7���#��)̌4����:�� H+�f��^��bt�J����h�\7c4���e=���IS��U0�Tzma�Z��.�mAX���XP�°i;��t�O��?�m
�pN݉:�2�%^9��;b �����כ�in���?��v�����o���&��T����� �Ou* Q���� ���4\ԢR50g)���y7�\�<����C�6f�� ��$������RU�)������Bp��b����5����L�L��A���6�ی�_"m�K��V�#�?!0=���k�n;����l��[�/e��əbfxPz!��4b��٘��
l$�Q���]�2��%�j������R�=��I�z~2c�p�{�ٕ���c�e������מ�����Z`�i.�n�Pg��H�\�>0��������ｶ�1�Cv7<��T�������rõ��Qu�B��sA���6U��ߌ�f�3���>p>��?i�|&��)����Yf�vP	����t�*-p� P1WD~1P�DTK)�wRYh)�b��="�J�6!��s��S^v���X�|��Яtw��-��X5w)����T��5�J<>-���<�IZH�a�Z���e�Qw�ǁ�V������i;���<���p�@mH��7��p�쯅�=��JH4�/����I�0oJ�C�P�q�&��x}�!\.�9QԾ���Ay��:n���h���Ö����C�_O�	b�H��n���{��;�L�%�WJ���{6������2��mꓭXc��*sc�� �b��=�@�H�o��O�o�j�W������o� n���t� >��T�d�<L�u�o;��J���PMi�W��Aq�V�A�h��V"w�r�_�Ÿ��+v�����*ӠD�<Ǚx��Y��;ѯ��4���S�n?�����_(�~.,��w|u��y	�UIa��8���)����m�n��<��79�.��씁��r#�(��xWu�N����]]A�M�����E�����ݕ���e�تG^�����(���J�O:�|������@`b�"1�Veo&�=%;}�˲�{�0����0Vjz�kr�듞��^̀�c��_���m;H�?�.K1`X5K�1�i�%��W7A�J�IצI���� �����R#��;�XT��4�[�ti��7���;/LE��D�:`�l���Le�{� Ư?3Ų�k���iA2��Wl��jBe�\�.����o�t��a0k̢{�n��6]ڽ�� ���"���o��լ��-��ڮ��_72ݟ��O�-��i'z�"9 �y\�EUP{�c�n7u�:�xS�gt���ߑ��n?)�Z�_K�ߦ�k��cE�l���H~��O?d ����`e�.g�g��~����J~� k�][�B mj�jL�wTQ���_����ޓ�}��}�r�Q�+�L�*%B�Sfz4,�>�F�V,������ߙ����%���r�1ޫvu��CA�꾒�����"�#:���	�oqTb�9ջ��9���|������7v�~~d��zO�^>�C�X�K��X�b�Yh(MN�`���>R%Xg�w3�83�
�:�����q���uw�?���X�v~���a>I?k�'!�s����9ѓ�]tKηo�D>�����4����|�s�� mn���HZ�m}�؉�Pշ��m�TlV�I�L̸�������P�*B��t1������L�O��3��q>V��9���-11І��O�ه,Yl"��5 � <aT��ڵ��i�<x��w0��2SH�t}Mq��8����{3�=w\kA;�W��,ӾX���B�٨/�zW�q]��/7x�8&usq��m�",�Rf&Bx�z� ��h�c�xP~��
{ɢ1�/_}��!��|��������`�n�`.%�у���Kc�ti����-�����@�l��~�g:~���{?���D��%2 +%`)�w��O��k?SAf����Iw�q����5@5e\zn.�VS0�a��,	<�������0��p�>c](��*�r�<E����`g�$�８�҂�!c��s��B��z�2�R�+ ��%�0 ]��ĸ�Y�ǀ95 ��-��뷈*؁�Ѽ�:�������?_�j�>�Y�P�y�r�
��AK���)=P;��Q_N���I{o�RmKY�����C�l= ���$�_��_� &Z�ep/�Ҍ���{Yk�� �-��8D��ec���I�{ߕ͏��G�J�Tę-T� z2, ��n�C�O
\2�yQ�w~���-�+�	k��� �����B]�S�k���a��Z �-�զ�{m����Ѐ��v��� �<E�
�]ʺ`��K'�u�?�(�&�+E+���(��.��A�ݝ�t<���.�B���d(�5���V�\]�(����xt���^����x整qs�.;,��>�BZ�'1��K�_��NF�)�ﵝ��<��y*�2�.ͻ��3B>+UjØ6�k�5�!>KMR���`o���H�0���)���4��w-�x�A���������P��8r�����ϋ�_E�m�ڭt߿�va�<=�h�G�8��%��V|��#oD� �9S���H�@���(l|�%��?c����<� �����U�zz�}���ճ@��J�fYT�%��]�"e���f�=��3���#P������>MZ$�L��͒�U#ܮ��p�ss�IE!������4�j���3��y3ϵ\�2���S����M��׿6�^�.@��������� �)���<.\�wF�y�=���Rr���'������芒����5�T)x���Ź���ٞ۠j�h
�kU�Ϧ	˪�b>To�-�-1��0@�IWRV3��\�{'	��ٳ���7'g�$����ג�ۏS�.-�`�j�j�<�H�
��89���
�G)�5��,�����~�nUX� � l;J$w�K����27TJ�`pxֵ�5&�+~׻N��k���$r1��7��W��E���5\5#�T��iܷy���.i$�������l_�ԋ"��Km�>�4G�qnHh��R��\�1T��i���)��zT���@�l�py��V����)ȋ��x�a������	����P�"K���G�R� ϭ��y��f��|M:\��${L3T�������zz`í%3T��c+�Q��b��=��]�5M曪����� W���?h})�T ��5�70��,���{Zֻ���z���n<�t�hb}��Ԅ#�ȏ���f�i@��WUݳ��z�8�N�Ut�gJ�������������t�S��l�H����
�XIw9�<b�������0��)�����:���[D\t� Tb�aҼV7*�>KW�J�'�o�c`�&?�{��-���y��#��9����y��=~�N�&���Y�\r�EvxV��2��e�5Vۛv`_I�StL�-�,�*�m��� w�ߖ����p�d����ǩ>V۳�5�5�\��J��`�#��r׺�:d)	(zI�l���n䕞��YmY<��s��ސ�]�g>��y�^�zפy��ή簎�t�Z���{LyOEIy������M>;)�,�Y�)�L��N�� ���T����fv
v�V��b~)Tr� ��O3��n{$=����>ر�ͱ�����ゴG׍�C���9zQ������+�@S���"J�wi�b;;j�����Ca��s'�љ0W�=������lT8ÿ5i�o����E���^��˦{��f ��~D�"/sI�E�y���k
�r�'�]-��P���
�Xx�Uc�~�j]��aWw��9钦i�m�|!=P�o�N��y��荰:(���� � V���Yƛ��S�a_�n+"����6�� �]�pp-��?��,~ �Ɋ�:�[Ym�@#���2����]\[�|��� U����~�����0�>жj�B���P�P+T�y�o+�����]���� �i`���}��1��I������j��k+����}{�X�W@�����I�D	�ŷ��-Ƴـ�>v9eqܹ�x��p�\��y�Ϸ�!z8��]M���|-Q��+:�j�C1���u>a��s���-kj�4�����+-T�� �H#��N��T��U찜�+��Ws<�k���-۬��㢝��R�m�f%ͣ.�]�8�n�\�_lϼ�X��k�ˆ��}^|���oL��{��\V�?�zO�jYI]'�V�����woJy�ؐRE�y�N�i�H�?�)�}$՛�
�}��WXvJw�g~pK�N[	�ҪB��ub�� %"J2uv Ԏh�������clq���x<����ӇmY]�.I$C�5��}h���q�$r��zGߔP�'����0�ۨ����M?ס�`��*��ü5A<�/����Hq`�դ�/2 �����Ƕ��60��E�����j��`�A����#��
�W-d��՘.0��Y�TǼ둈RA,���M�&����C������|��<o�'�iKO0��-bn9Ww�x�5�X�"�}ͫ�6�ڀ	/�(U~ݖ��2�;�m�~Z��C��c��;��oE�{.����ݴ,����R?3�NcpoƷ��M�bH�#�(��1�=��8Oη�S6�H���c1r�M�ύ�76���%vS��QH�i55 �l+�4g�gy�+nM��C�IZM��;�V�;k�T��z�ch��:������Ü�����ߏ��N��Of8ٔ�ʼ���*���m��w+��w�j��
T�-��5ס3��i�{��Pi��Q'Lt7�q�xvz�](��f�k��Z6�cf �Q����<��h��[O�Eo��y=]�_,T��(���_UU�Ƙ��vf������~jpӃ� Ug��e�E�jƟ<��e|����u2�����-t�nc�M^�1	�C�&d�� s�(.>����j��'����u[��+���@�5�"-��7?O�1�{nz��JWPiw���z[g��O���0��n���8�B2�ew��gu5��BIMu�F��V�F�j4Wq��f$XQ�W����W�s��5z��HB��j� �J����Y4*�u��f]��� 6��J��P�����ߏ���:��u�:�M�"�3Ԧԯ��������z��Cw"�s�����+,�y�7����R��Q�:����	�$`�Xf:�� ��\��xJ5�T�9�m*���AHE്2�u��!�Hz�d�ߜ�I~N ����v�5V�I=&+:o2�]�:fOF�z$9��d��N��a�z�j,Be���=�>���#�F�fn�
���1�՘g�U��n�y������gX�l?Խ�BDR�vǳ74jK���&7�W6������_I^+�`��BC/ k~�)"
Xl��Ŏ=r�)?
:H�pF�m����O������g��c��Q_�SB��u���:�?{�T�R�k�1�w��(��S0�=�"���6�Ľ��g�A���-HJ����qW�Rڧ�~�=i���T��u3o���T�^ ��KNT�2E�1�+H���{��i��a��M۶�A��@e��>~W�S=�F��k����{�9G����[!=M0T�(��-)'4��`�kl;SW�2BV�4�I�I�}m���N@��~�]���,=&=֘�3^���� �-��{��#ž�!>ˈ5�2^�|b�]p>]�ǎ�T��I�mA��1��t�B�@��{] *����@�Q�LNR���8h�,��M%�ց)]�z����9"��DXiJtr�sS>-���:���Sa����Wl�)vK����~�5s�["�:����j�~C�Y���i��J��*ƪϿ�T��2#_���~�_^���[E^�C�LWE�y��}�oO�+����2D�B�Ű�?L@u|H�`�t��1���8.�%�	ѿĘc��n�>>ǆz��6�K~ƀ}C�V?M����0�_j��+N�@?�[\]���,,�֨1�'��H�JV�_��Qj���D�gQ��V�y��x���-(L��$�+�宺�i�N6���������O50`7�x����TI#�ɒ��P!����_u�Th�t�[��yC�c�6%��zX�����!~���`���OM�s�"F��r���������0v�������A����LW�-�|\�z�=����fb��W�(>=���BI��ef�i��E�"�ܞ��WB�M]�I�=��Qb`p�^��w��)s�*�9DpNn�Jnp�}�C5��Ŷ���Wm�%�� �X�P��� n�R�</8��Ѱ�T���J�b��b��V�w��Ѩ��4��ɶg�a�*�l�0��S(���u���DG���B�ҫ��b��`�4�>�[�����i�(��ٳ���.�x��W�[�~�O�z����G���usC�j�u�m�t��^*`_u�CZ��ϯ�4�Wȝ
��$w��f�t�G|���{����+S�b����yLu��bزj��q�87葦էu%���߫M���e@��vA�O݁��ձ#Ot�hA�����~<��W�w@���~�<e�%&��F"L��w�c(9����K���� oE?���u�*v\�������V��*D�Q�U�9��.i�<���Jm|m9-mC�Yҁ������&�����G?�CL+6�1[�&Zl�*��a�=@�����m��'~��-��������ȑ�Yf�.�~��؄���e��V�15`:W��m�����]̷���PC��,Ă!n��u-6�C��\`�����8"��o�=�[ۛ���t�`˩?��!�éS���-�RY����7����r��ۡ����q��َ�?��!��+ғj�������+��hx�X ؑH���9�*[_tJ��ōW9���k��`HJ�;�f��p�p-i����o-��v�"U
��#��(φ��h-R��{�b�G�p��Q�t�T�z�ZɌ�ו�ꈚ����es��R�k���%�B��G�]w ��UʃV��GL�q�S� ��m��Z�d���Q�D�du�o^	�D��3�,�����k�\D1�:�)F��4�0|E<ʛ�ԇ��KI�)K=��5"ʅ8�D}���+�F���ϰ�GW���tZ16��_y��:�p�ȷ�t��l	��6\>�A���N�7M�}��߇�I��kB<��Sw�6&�a��Yx��N��b��X�(�I}�ni�7����^�e�o3��. 7<Y�sy�`V{B*����ӡ@�$�y����'9��:��,m]M�o����yĞ�
��2�=��*�~���~��� �880:9,��>���@50��P�:�ql^����~~߭����!�d{)�K�u�p�i?9AH�\yj�/�\�AQLr�U*��1xO<�L�e��BcҾw���t�����bQ��<4�S�y5^� 	�@�q�K��������}-9����t]x ��L:O̽����Xa��_B���E\w�X���;-�V�ė�?�'`:���e��_SڸƳ��d1��9q��`���;�6�L��0�.��+vk����;U�.�p������?ޟ3��ՈM*	HG#^ʽ�ͦ�� 5e�Ӷ��F��$m��CFx��1��l��7�'��҄�����b?p,�U���~��$N��wZ#��_o�-v13pO�D7 ��&�Ӈ��^ӱ��T�~�|?�սb�:�Ѻ+�Ua��g�������q���;*�L�7���Ȱx��# 7*��J�s���w4���Wѩ��$���)�l"g�D�@���S`������Z��0H,�����)�����5��DC���/"E�:J�<'�y���ߨ�2ߑ�q��
`'�EF�2P�4�]��>�f��w��{_K�=�E�m(>ѓJ���$�`0ݶ�=e�/�^^�Ʌq��?P���49g�jW�H��$Ų����c��u�p�%�5J� a����m�y��e�K�͔��]"���-�eZ���h��;�K	O���jw�w+�b��Y?2\i�)ѬX�F�~�L
M�IQe;���;�s�1����4i�`	?�`���[�90*����EwB��+9܃6���"p��W�cC�G�q�Gw��Z���ƻIh�Usb�2�>��fH��N���A N`��AJn�2�:�,W���2<'��6kL���m,Z,׭?�S�HJ�ס�^4t�aXҟcU%b�bV �f���D
]��x�t?Vס��a!�ME�h�'�3���(<Y�Oj��dR��q4DmSy�k�����$d�-�V$Ll��#S�};� ���]��M���T=Y4~�5B��C�z� W����m)��?�����ޯ Z\�0g��K[�7�{�:TL����p��\1������F��84L����Kb�Ҕ�i���ş��X(�v��+����&�?�,*�%��D
x�0��B�mwCzd�H"�4�*[ro�)�Wnd�ۦ���\B�yf�yc��8{�����y߯���'��;ݜ�P�Jk���u�uWF�)����r)?�<C���祧���n ��_�QX�s$V�l���������
�yI�ޏ��L˟��̆����瞘3��a ���V��S{,Ϩn`��t��J����g��$��������:���㩋/�a��i���y�[�Dqq�� uH����s�J��s��i>v��-$52��M_��I��yG���(�l��Vʶn±ߝ����2kL��ȟj�N�[����E�UگV�"Z��="�Ĥ���>��D��<g�٣�gk� 0R�������2�|4���7�_ w��Bw�_�&�~�b󸩸�����D�<㥩�������g��gG�[�B�u��I�=.�Ӫ)��g�	 E�S���j��V՟�6T>2!�q��#~�F�WD��Ţ���W�2w�O����b�-���*a�	�~�_Ďvu� V4���%��1���Eq=��Y�D[L��ۈ��O����G�ia��h��s[1�ȑ�O�T�r���D&��y\�� �#K�ERd�w��*��o��i�g[���=�V�X�_c���qTO@Jm�Ĉ�[���j��c\�Ѹ�J]$�ޞ�%dQ�]��JOT�T��Wrq+�v�^�+�-�+��vpN�OE�U�5y;\
�vt�R0l���Y� �=�廞N���U�@�-��
��X(�c��@�/dE &�D=�0�;�pmb��8'��XZ�^N�1C�`]Y��>i�f0��Ey���^�/l�N`�B�3(��)W*����``i��s =�§I7��;��n� W2���Ρ���gd�f��D?X�b��q��FZ:\@����e��7����� ��f�����P3�,�����|S��&����C����ЯYu��|����ov����ʢ%_,0v�d�����z�H	�*�ZyE��X]uV;Y��3h�y�+�����=�w}
6gZ+� 1˿�N=pI�Z��f�)���'_Q[��g�k��Wי�Wi�1`d9ZIw{�������$0Ԁ86@ecQ��>7�k]h���lqo�o�}����	G=.i;�i�.�yNP��G�ո�ڰ!�mA_ęo�P�~0��T�;��N�j �� T�h��b{����������+���`-
�`Kt�J@� ,��iT���C�A�ҷ��X�N;���)B�!���B2��X �e|�X������X�#���9h���U����1�Ĵ�L�%Pt��@.�ޮ���_+�T�*�9`�}���%B��I\#M �4[�+pVU�D��_'(�[H����>�i�=l���M2�p�I/���*�[HI�J���Cg�gc[`��#jH�j�*��$x�E������2�n�"Um�B��z����&�AU��6Pm�1�{��#�L�l/�F'ߐv=�p�X������<��y��=�y���j��I�2�g��;�jp��*K��W�.zC:;�9��L$?O��]�g>���6$���~wݪÀlR
�ZL��8YȘDY�ߛ�/Lύ656�S~,Q�W��,���
�����Ӈ�n [hf�����Dލ�Lky�O!*�X��a�N�`kbι�^�g~�F�C��Z0R?��F�7z��N��o͓i�����'~�4R�W=�G�*��g�h>V. ��?�A��Nw�o�����j�l/�	c�i��C�&�H��%/ eӕ6}m�ٖ��E%�eC��n��O33b��Ql�k��%���T �`��V�3+e*Vd�t�g�Ok�8��@`�����UѠBWs*�Z�s�����} IqFz� ���^�`��q��~�#�nyT5�&�N<�����C*�;n��c���~��+��)?��EFiW��yp�]
l���>�������{��z��|zy�d<k��ߣ'}�\��8]�;#׭�����>;&�ׯN�a��xc�={�ua*�������k�������K�A�Ӭ��Ӷ�C+t9���κ5�P���50������Ũ���ϖ��r��]�)���\����(��?(��K�x��o���Uf��;O߄�{��%�n�%Y�Y'Z��\��@E��"JK©��ϝk����_�2�1�rW��0ΑIp�Q^����5�-2�ᒃ����}T4����1���Q*��}{�w�x�=�c�b@@{��-�cZ�ֱ}�T@�n�:ކ!f<�"����Ç�1%��U��g�*�][��3��+��%��>�����@��Xc���_���6�k9@�Z��.��6�j9��ЍD��@��������QkcFރ�X۽����
ծ;�����v���.O�
s�Rs*A���`��K���H��L���rm\ ���X̪8�2�uu;t����r�/Qe;�*�,pl�n]L�
y�������4��&�� ��9�93B���!6��{�H��Z���{���/�?L�}�c��`�^��uc*>�#�=� ��\�z�E��b;��҉a�͠�\�� ��[7&����\��_~������?z��
]hZԋ5�H����(/�0�Dg�)�u3�ƍ>݁�9/0�vH�jb��;�����OX=�Mim�n{zW��5 ��^�}���������'՛r,�~m?��u.1��n�m�A^�k�2��36�`��`���_�g�)�$3Nl���v�X�'�~v��b.�k#��4@]͎�V|s����/�c	n��A�|�z�f�kʄK�g������"�
 	ۉ+7EG�ќ;�U��'�Lo�W�
7�|��鑵/�z:}�c�i5KaU�e�o@}���;�]��M�r4�o�7�j�N^5�
���X����#�3��H]��L��E�ձn���v3��Q3y��]N���4}̟`��4�ZXL�f�K�ݙ���"S�������{������U, -T�+.	T������cF��ߺ*���w���H�Z�K+
�mT���|.\50�������E���{"��M�r�����t=7��p��[60mgp� D�jz�na�����.����Ed�;���V0����]�%�M�g�F;v��dy���C�!���� n��y���flth�\.��/1�:��q��u�=�n���~�E�Z�T�^�h���4��]�vTs��g��w��E�gX���o�.��-��9�뿘����ݥ��p7V���x�y�t�}[X: .s� �*���o�q�������[V����J��_�M?"���SwJ�h��9�72�=tuj����s�F����	�����}�:�V9�}�����%��;�7i���_��ڇ�,��b�&�3�S�����>� U���z#6`� ��"��uoŎ,�D�na�b�-��s�:���D{�58`�3���d[D`X��e/
���;3Ĺ�w��F�J�c1b-��ь�k\˰ž˂�z��P�,�������l]y�}!����c��c�2�xN�2�nGV_w��T�Z#�٤��"aծC;��#(��F�o������̨��X\����+�<m��̷w�o�c����B��w����J����Iv�l�>������������ϑ�[f=�|�}N�.��������8-Ĉ��vR�σ��EI�{��=ABp]��u��!-J���zp�S�W���[ r_�|�ۭ��w��r�d����ڮ���Я.�W������x��2pu�
�6��51�b��y���-��(��!i[V+�M�����9/P�s�R)��'����)���O��F``�R��1[��<�;�˗A���@ԯ�����j��ˁ���ȣm�*L@ʝ��W��*��r�fEBT���e1��C]տ]u�bbw�����Xc���a��0|�wi�P��]�Z����³�(,��������c����q�ms����}Gە�[�u���v�૟��897C�A	¹Ɯ���[d8��ȧ.?�`}�Zc`��O�E`��yS{9a�U�e+z�U�\LY��`��W��75o$ �j�t+[����͗Q~5�j��|�Pz0-t"��F�j�'�12��8��
&�N���Kl�LX���ٌw����c!�.l�BL*��J���V�=���:�*����-cv��29x�ccB/  �����B��Բ:Әg�9^�_-a+)�헒kunj�NJ����������s*�YP���		�\���>S�F]ME��qU9UJ��P.}nk��Ab������m$�����<zN�2��ل+�ހ������v5 H�(�����< Nb������ kc�E>.����>�t����o������3��\�8�wv�����^e��Tb7IN��i ���?dZܣ$����؄��RQ��ٙ��fw#vl9����zp+���UCM�q�� 6�(4
3��G⪪á����	xE;���3V�u�.v���-��k�ݕP�(��e�8.]��Eˋ�g��`�D�G��2-�]Q�Em�W�|7u��g��A<����2>��Ѥ$5q���p���ʁZ� �sTuq���rU���^9���2�X,j�<cx��d�σM��zCJ�2���+�޵����p�Z�t����j:��-��}&��>�����n*���~c*��$�p\�]K �R�'D���aR�5����v�͊�v}jc��d�1�N�WpTp�XH��m�� �*��[�MQ8�2�J�6_�Rwѡ��7��;{�}3��#�6Ϥ �;`�h��Z�K:GW�v�O��x��{�R��h[����{a��}3T�G�6�PS�1����8~����gU��ms�XR�.���G�i�H��/�dgt�������g�/j������#�\�W���:�&��Ogۆ�U/�΀��&�K��lj��E��\��>��.<?|$���1X\`ɭ���`v|Yڶ���쭉�/o�u�h�S${>%�������������wkq&�c��.^&4o����p�����"������Ex������/H�8�'�eҤ�20�]^���̠��h��ʄpu���q���]�Z`ld��ܶ��a���{%Gr#Kԁ 3�!�V�l������Ϊ��+3� .�q��,M�ĒmH�YI�8܏�U8@ ,@w��}¦5�S��;$��h�<��񝱞M@�rz< �=�E��� 0=�f�v��W����S�\ƶ򐌠���������I�xr�T��"���k�����D�q�}�Մ8
�5I�{c����N�I�����w�P������#f���%�*�zѹ�wʏ-��T�<ָD� ⻲����Y�N��_Re�Xp��"5�<�̭���i��Q��x�Q/�ԅɳi��hA�
}DV`a��߽O�Zr��>�����L���D�X����0h�v�zT��&�s�{���w��`��wǺN�-�s��ui�|jFB�db��"����O�g���i�վ�	X��YkϢ:x��d^j�{J��1�Jjf�e���X��qZ��j�LL����b��9�Za|[����w���ݫ��ze�H��� u�4�m0��/Lc�9���G�j�Э5��q��)Cb��\����V��f��r=�Ȑ�V�g&~6� ̧�c;�ۑ�����p�V"�k�~�}G���5+Zk��p,�u~1�1�Z��*r�G ����|(#�a[�ږ�Oڊq"[	�������-��>wJ��� �L�ZI:/a�Y���W���f��X�|#i)�}�����?��4�]0�>@�BZC�����$C����BM��^�SU7����=��������j�@�-�giS/�9�Q�㎭��Z{1���A��q�{��_%���G����t*��GeK�Ico��h?@j�B�1~>���΄��$����q�����H�`{��2:ZG9�ɲ׊i�v�j�M�Kp�dܹ6N��l"�ÿ�N���չ�U�%��;L�V����b?l?��d����y����#�X
� 6K��j*���K3i9�((<ͨ��)���W*;jl�K���I��nG�m�@B*�I�I�EN��E�o秣�Q.�3UC�vR���l)U������`,͸`��1��{��Hd�M�f\B��A�aQ���Rsq�	�~�0P��G�<H(�TK��wa�u��7�u�U��"�8��N�����=�E�{�/�AL~��v�,�(h�{��,��J/�3%W���@�r��'�s

�U�j�N���Z�%Q��iR�^���G}�lB�r�Ip;��>���6�7���Bm��d���i����h��T��~o��$2��@��g�^s��8��D�LkX
߃Z��jؘ�r�'�?�6�����Vb4\Y�Sj��[��e�X]}��jKH�ԇՈad�I��S�z��x��&�!<����5��N�U�@(��\����/��<��Q\�.*$���6do}	y�㬦j��1�B���$��"L�V�{1)܏c��N�*23�r��,����7�L��(M�iu>.6�Exa|3�]&���`s�"���G���Xk��и��e��{+
��za�����a��gp��3���K���m]��B��~����P<9�k����  ��cE��"�'�k�Q9����O���(�:�Q,ˤ�0U����M^��sR���/fm|���U�����H؀�$�~�h�*T��".i��&#�͛LkF8
�b���b"��L���Q>�V��.����mc��`bC�(�Z_�܌�IM߷����y�$��;�����\��I-/���Jz���w Sf�1�J׸�1a	n��������۵��#��.��{�E��L�A�ެ2W�QI�l` �U�����X�v�u��v��(2��}��6�e������bNɷ"��W�'��7n^����}<ǆ���&������Յ�S͑ʨ�
�ZI�-*Qi[(ۄs�q{�Rx���70�t���yTG�3���^�+)��y|��I*"�9��V4�����Y�� �A��JUs�O	-������l�B�5V6o��`�]�����LİZY��C�"7Z��B��^���C�����z�(+�\�JK58$�4G��F=Gjh��r���k��f�^�_sONQSԻ�J�vL�'l�,��o:3��i��G��en�$��$��Ϊ��A�e6%ڵkCL�k�سW��a�4�﯅�Fd0sRԂ%V:��v�%l>��[>�(�xBՑxg0Z��m:��=���%��v�3�}�ĩ���KcLw�ڍ��Z�O �	_r�n�$��l���~|��[l(�u�V&��j��)�s�U6(ԃt"�BUb�S�bNP�lP�Z��F+�����f���H� ��Yc��,-�ZoG��J<T�����wҵD�B�P�l.�h8�ÀyB���e��_����&��63�df{k52�9[OmhQ��h�}{~ƈ�]��
$ߐ�y�qS��T鞽�z��/��X�����������=k���Gҩ]�	�E4��ۛ�i�t���o{���Ŋ��X����{��_/5&'��f�d�����7����SK�Z�>��L�Y�K�-�t|����9�^^_�ӧOr�g�U���&|��;��:��M^^NV�ں"�3�'KZ9����k��;0��m|��07����T��!�r
�wmG�N��A�A$�!7\���6�T��uz5B���_��w��VE��D���߫��,4	zG7�f�m�y�MR,��/���`c��,4�"��4!ݍw�c'���^�ظ��^��8O@P��ٵw����*��
��4i8�<yoɮ�Ld�-y�zQ4H�#��
6����ؔD�\m}��3F1+� ��l�p�}�yie�H�bƯ%!����U�g�;A�0F�r��[T�z��K_�@!`��G�S��=����ˊ�� ��C�}�4�)Qyͅ�Ҭ>����_`���oz��ps(:���3yAͦ�8�<��ps�_�^ߡ��/��4���/���t��/Z�D�����ϛϹ2Y��oo�o~����}̴�� ��}���<��_�H�<�!0���������&��$���I�f�������_3��6�mC�Y��m�Mb����i�D�3�M��FToe�l��E���I����s#�Y9�P7��{��D�(vGi�ȉ��*�����JG뺵�0v�V�0��v��C�p�s���Z79D��(z����z��gĚ(��z���1�N -�W�O�s$R<:#2 ��������م�^EC`v`�X������y�<i�I2�i�饞��n�l�1����1�i^����,뿝]00�%R�l]�U�F� �m��I����l�0:�{�i�؜���u�UD5=;�b���2��.�f{E�k;}�kdE�����"[pX�I��LM+�y�@Ż�Eȃ&�O�C���0�@%	)��*{��ρN�^�I��4������\�3�7��g�̐��HCM{M�\���*�;3}��Պv[�]�#��[xK���dT��e�M���UyV��	���WL�f4��V*��Ԗ9�kê
�g�����F�����	�G�O"�d����팢�V,�Rm@03�_�"�e����
���^��'4d��58u�U[�4�Q�����ov>��(i�ʊ�C#镡Dy�3��6!�-D�n��|;/l�aO԰ ���{u��B��5���iϢ(ۃ�ִL�����r���CF���ߣH2��ެ��_TX�X�aBL�/vړ����o��L��q��,uq����)xΩ��cOa�4���8��煢�V�Τ�#����U���k��4�'G��d3#S�)�Đ����,��3�j�ى�������!3;���]M��s�n�b#�.s�E2ӈZ	/
H_w�w��	���N�
�҈�<���߃�ڒ�^�K��U�-�p��q��3Ckn�G�C��v5�T��)
V�!��X&lԉ�i�l�I�3�[��R����0A�}��3�3Z��Cڳ���C@}��M�1�Se�jDQ��0b�p�>v�7�-���T	�"W
r-!���4��O�� 
�(E�<,�p`���Nr���������L��a��ٜf�7�c������TU/�^h)��|;λ�x��6ҭ��?#��_Ɲ��-B�L}�V��j�
ڍXA��g�>쬎>x�oK�KCH�B8T;=�����n���hvE����q��JHƊPS5��~�	x���A��tH�i�\S�8�ܼ��嚵M�I2H�I�a�X ���@�(y�{7�W*�),�Sf�ؔHw����r;�0�)^�����,s5g2���c>ug�[T0J�4��q������F�^G���5o;�'�K]���3,s eH΋,�y<Ӝs4��������6[�N���OO���4����y@��P^!Tx䏵9��[�C�N��=�Ǿ��>8sU`�-�n���r��-z���l��|[0�:/��r�V��3�'��#�� o]L�3��T� �&h'R�Z��$Z�(�M�����J6�w*l}z�߫%��Ή��w���[=ې_I�P	�a�+㶷6��YP��LZА�{8=2A!��c��9+KL����͝R9�z��<��;��<�%�L�b_��Gٯ�(�[7�{$�M�060쩯���A��W�LFg���:�2vzn&?թ�#T�O�gl�&�s�D�(,,��ζ>�7���v��2���2��)�W5ѢP>��)�	���1���r|�JAN+��z��_Lêh�`���mP8�F�`�ҋ0�'�{�����w+��&85��5m��i�!��j�|?���+���	��֒���#���X�Y���5��8���=�k�iA��m���5j�YǓj�X�ǿ)�$�k��q��1g����(���m���j�ͷKm��/��Mj� .�P���R���q�(eu�Ӓ�ȀL���Cj�`�p1����]��TX�,�:S�$S���c�j�C�w�+�r�%oB�2�tQ+љ09y��G�B�5��B��5#��%\�~ؼ�L*?>���@�����
��j�F��=l|V.��g������M0ӭ��Sv�d���5�k[6�N�����i��B�%�����mM��Gj@r��{�e��c3��x�xo8S`�GѲ��S�	�\����X��O����,�=��z�מ��	) ���ڈO�]������"Q_v&](B�����2��o��VP�S��x�DT�o��>C�����o�gx��4㪳2�vc������	7Uo��e���P��0�8�M��	Ǟm5Vw���`5X�iZ�B��P��Q�U�pT�獵��1�w	�z�����=���'����i��I���(��߹Q4���7[x񝙽$1��f7A8BOD-R��u�xO�cF�u��$t�
�C
/��U���ڜ5��zcHoo��[��ǯ�����c7���P��6<�/%�5�R�&�L�ړ`,�<�Y7�j	��hc�0D}�}b���/�ݷ�#���QZ���D��L5��a����K�/6��6G��{}���;&�R���輡�Mi�RƐz��m[/�ւ>��i�8\�ſ�x������[�-%�H؍�{a�<gþS2EB7�M�~�r[�ͥ�� l���4Tx*�C�|dTGa7�T[�&��N��mj:���3V�6�{��&Ҝk{�@ja�(��߭��0Uf�D��C�1Kk06{��3e[6�M��iv"��S��EL�2�mX�:��i<��'���*�S�O���m[�P�0���L�Ż�l��Ce�۸h���9g����X;�;1�B��d�����:'Za*v�`'mY];��r�P�T�����5Uu�WiQ_L��i(6�Z��53�Ն<BS��0ܾ}K���+Ғ>�_t쟔aFFR�L �����k�rU ��g��~|.G2b0���p��SM���W��=�T3��p.�~�1Oz��,�.�t
�-�)�sꂖ����F��gI˰i�<�`n�p��za��s��(A�W�Af6Tk�tđ�$�bW�j���ͷ_������G��6�ʗ��"�(R���g0�r.������I�y����_H5v'�(�Z7Fe��D���X�$�#̇�=g���M�<���k��D�;���?"LƑ(TK=`��8��g�W�з�9w�����o[y�q�o=�J��7�jo���FǋJ�g$�󫲠�b#���h.d���&�gf��S�`��hP��%Z�Jt�t\<|��9����N�1g[ B�G�F��e���P\i��rU3T�s�&�;��˟�l�X���]�5����C.>F7AM�Ȩ3t��j�1�������I�銨ܟ�Q���؎f!��6W`�����A�v�i��F��Y��v�K��f��2I���#��RR+#�8�풽�/N�����o��/����o��j�H���C]�0��Sf��1����V��)<�(e�N��{�5�s�%_Z�gƆ�{��m��87ŞiXD,�M�y������k SS��Tbi�a��f���L�
s��}u[��	L5��BBQ�h�l��L9F�3��Q&�Gr�]	�3=lz�6#�_r�Z�?i9;L4@s&@"�l�HM�a��Ĕ�K5�6����尛 �s���eV���f�H�L]	%�����,�Xl�b�;-%�
�$�����n�C�"~���tfꜼ��/7���?�I�����_n?�T�I�e4���4	f���7	�|��zW�iZ�6���{�sjz���S?�4�Vm�5� k`���i6��H�L�,�DbQb��������*2�DnA4Z�K���T��M^N��Vr��ڢ�H/g7���ę�:���
�� @E���9
�����2�Tһ�>�IY���E��|m�y�*N6ôU.�L��Jl�@��?���ȕPR2Iu Fv��ӏ5 �� ��'a�kɀu��H�S���6�=*s��]#eѢm�2�C��� jz�����y�w:%��
[s��qW����ζ5���fF�*�{�)�d^��p��<�J̯3�f ��S7(l	� �[9�n�r���E�ts*9"D|���12�`�k�">t���ט0�=5KS�����p����s@�� 0�}c�z|܄ɷ)�h�|c�_���A�wۗ�M4��sP$PMr�駛'e�[����n?���>��`��s
|�� UU�Y�?�P/�a�t�&�%�^CUDq�l��z������E��?o4�'fD[�Z8�F���|�0@�VL��Qh�����|��k.�)BJ���x`c�6)��Cc�om�`0ր�6pGf�VjV�Q��:l�S��цei�T��oB/bB�NhL�����;)�PKXpV֦%} �����u?�����F	=v�&��b��W)~�S�������m|Pm��2ȼ!�ZJa趒Z��t����R��p>LIn�F�݈����Yk�Ջߩ��j]@�z@ڂ�B��S8i����<"V�Q�٫�j�.�h�fe�+LM9}����f�WE���eH��އ'�d��tA��Dߛ�|�rB#ە�jv�2y���wg�a����E��gON=��(�X�������h_�����y����'���~.��`{�)0�36��2cp�HZS �^֙�~�cR4����禮�}-�����_1�U���1�?.6'���B�p
mɨq_f�u���-Y� �B���3;����,�:ԥF�J"΢} �x�1�J�s����s�
��/�?�g���o+���Q9�p����8Y�����-�3{uKsBn=l�`�ծ�����H�(���c���̠ab᳾[e*��@�Y\C��d���wW����bw�X�*��ZD�����֓�~�kG�F	����k0�1:E�~I���y��::�XQg��ժyЀԇ����a�p��^��~~���l��R~b�tC����
d�f�-��.��u�I]P�0�d�M���
�iբC���5�U���.�����s9�����*�RҌ��YW`Ǆ�Y-�0�8�u�0��w�
��S����9�3�D��;���  ��IDATr��l3�@m��'��N�q��57<�5ig�+���;�DX$KCz�B��x��F�|�?�|G����s{���TO�P
�{0��80.����B�f�M2/y���]9��"h:kg-!n2�`�-R�cwh!�.u퐺Z������z�o��җ�����Z�۞7��A.�ORV}3,�3�k� R�}�_s2U`<��.s���5й�$3%��`w�3U	���w�!�����ΰr���#-�S=<�΃#��1����=�_��6.a�)R6�Pw�;��0�CG�@���5�VB�l�D'Q66��
�$��9��$Ђc�9���b�F~��F�lyF��1�\��2�����%4>�_���`a!�6p1R>*ԩM�I���t�}��A�	< )�:1�ޛ_9�$Q>։��:;��3�i5�LY<zx�������a���2�-jJ`�N/^e��zx_��r���D)xA䌎ÊI�)��%����KE���ό%��P���Z�z����5��������ҙ���s�8��T�ڭ �8��b�j�9��sǑa��r���� B6D9N�3�U/G��vg"���"Ҳ���vH!H�3'#ז���#$!���-��f��������&:"�ڜ̐,�!B��>��{X�2�;{�9-�!�:��f��;4H�� [��M��B�[��q��}��u}R�|�@h��;,L�A��[��Ѻ,�Y�3`��"�;����ٛaH3M0hr��yFM��@�x�?�h��<��zO/t4�]MOm�њ�*���Z��6�J�	���	�:cN��%����~���;V+�@y]�&��b��c�P�O5��P!�8��c��d@�2�K���;<Ȩp���.�p�B*�}\����]R���I�ʄ���6n���b�8�g�[n�����,L�̔e���T��8��`�/[,f�]}D��YG�߁�b�
�T�i�]{h�PY���U�f����r�Cd$Sda�G��&6����.�67�XW����'8�I �%��l���M^`�c�`��e:�)��I��{Tݵe};�-��L�h�`>p�P��6�oJvG�v�"���) �f�:�b��:�lC�2�@'�C�|�!d?���lA����["0έF����j����\9)[W�B�ИDE�=T'sqĢ��8j)7�<��	�$�;򖺮����g��	g��9	fӋ��a'>��[�{��~D#w��6C��-T��qSZh��K��ؘ>7�m��Y��#�����X%�1��(4�3&�<ۣ�HYf+l�Y�aᕠ%����մ���	�Ff��;3�w�hf�Nkez*!̕�<g~H��T����^md!�|7e|ӝ�Kdh|wF
Ĺثc�\�����s8�f+.�.p��wYZJ��򈐰k�%fX�J�:��6҄p򠅃��_�H5�$��U3V��R��
y*R�Ҥ��_vGlK�"])��]	aGp�1gyfc��ha�a!�;`�=3�8�o!�djQQ������)%R謌�������`��^�BM�l0�`�>w�3���m������5v������d�/3�c��FMv��L�u��Y	!�-��e�T����X�v��ח5������Mp!A6���lŗݚS���~E�~����c��s�k�0�=e�Ul
�=��}��b5.4�c'(���F%��^M�V�3n���#[P�m�ݘ*��Q��2ir�����y��y@M�*�"f^F�22,��-��Õ�6��]26QB�>�g읅�T�j��Hp�#���
�f��vP�dl��gs�`si�:̎<%��� �H�.��� �&f�U��xOܢ�Ƹ��� 칹	c ��ܕ��	��cA�0��%�Kk���oe��jn����� K����L4�����@}������J�W�t'�7Ӄn"��J�wD�s�?���
�+9�:�nDӘ��+�"H(J�E�%P̹��@�jK�1���C�v.���.�`ȡ������[q7W+�"��j����1B]�B��ݰc4á����4�m��D������=xh�,��#K��8���od?����������ן�r#3B^�
LT��y�wN)�F�QS`��)U�w�\�G� �s��N:�����e[��Cu;-*+C���sr�]SeQ��5�e����gG-���O��l�1� bZ|o���0	a�^�z/d#���Z>�u�#{,��3����ujRskH��Sؕ@b(r�1�����.=��Gh8�L$i�j��-�V�3ή���f��%�F+��%v�
�Qr�p���@��(�}m7��B��o�U���y^���U��sHK�eBK_N��t	E�0^�·Q���jˁ���\6)�w���ply���]�y�//�m�(�6g�2!�y�yZ`v/�#�������N)���71����̭(��B"[ե��lf�\גQI�Ǿ1����/d���U5m�����cʕ�qsN�:r4b�ք��afվ}��[`3!�YL��]���Ȓ܀��	�?L������&r����;�p(�9� ��Sr�X��=�K����ƒ�GV������Z{��h�cxф{��ZOt���d�]�Qe���,p��ʠ.�)����G4����P4� �� �Ϙ%`���h���ט�>�>��t�
�ޡ�`��)�F�\�I��d:+��E��(��y( /M(TR�qd�r�	��2� �i%s%SQM(��ExX�/���	fR�f�Z���Һ�Jƃ���}�nP���`����=&cQ�$72#-�w�)���Pl�"c��������B+�H�J[he�(�9	��%�}�a�k�<�UVgJX3���zh�����ѽI]w:�90TC�}�Z�����j��َ4�NSn#�*fG�����R[�~Z&I��@{ �f�M�L)I�Vrg \hQ�i$����Ʊt�X�?�a�zT���ɀ-쨺o5K�i������ŵ2h��������g/���$O9<2<?aG�`�x�rg{��3��;K��(�W�$QL�@�m�h�����Ьj�T!�(��jʜF7h��Qu�}��7;�I�*5�(��m��ܛ�sCyB�T�!���c��Ĉ�Pk�&T(����"�(;�2rrf��q�U�9��6���%[*r�{X�K@�k�̠�d�LkW�����[K"� �C;n�/�է�CȎH=�I�K����허��`�L�18^YP[t��=�[��#p���1��
[���mbX�H  @����H��~�o9#a����jo��~��k%>���[�g�����T�:�%|+BH{��ԺS�Hަ��(��g; �G�
��c<0������t�Uk5�*��	����V��8����`�R��̈́qe'Ȭҙ�&���+�M�&�Dj�@UsD���v�=e���5*/%g�-T9p���Y��D�dڐD�3|�QMH�ՃF����m���Dq����pAN$�4�<����F�D�I_#��bg�v��^׊��QH������1�H�����^�l�B��w�����`�B����D��-�0�(��b�H���-ь�k1���,L��Q��T�hu~EU�����b,2+17YE��h�.SJ'�Ҡ5�-��G�xj����r�O���Xb�ff��*d���YդLɃgI�#r��9�V��
�ԯ?'��.�'쯤jQ�cUw*X:i�X���s��м�'ߣIV��?W
�����!Z�J���)�_�g� 3d^#u���%S���408����95KN81�d�ް�{����0^3� �l���;�NŃ<L�1i�ֻ5_ p\;�^������&����4��j,<4��Gj���T�֑ tc��^����X���i�:�-����kV��,�K��6��1���G�(�j�#t���`o�3u��s�L*G� P�f��'�R����d�~ �D� )]��	�R�u��ѧ'G�DA��<����I4P��݈�����X�Љ�bZ}��IK@Ay@#0�=��N�&� &
�DFt��A�K�ʕ�1�et,G)D8��erՂ�#���ω���PQ�6����q�)�7�ݮ�ӊJ����s"��9�-��cF�xv�?R����6䶎%=�1��z�'�P�;q��FEķNz;��sGy�SÊ�W!'e�'�8l��52���lR�zE�e��������J�č�l�N�ړ�����ik]��L��}��B�*��
�W�2 ��S�'ơ΢9����L��;#�E��f2ҖP���LF�y�|�z|��4RR���m�?ҖiDH� U���\��ѱ�eF�JZ.�8�2��瓘i��9�lF�z���qx]�)�(�Z��!	'X2B��]3}lx_��e���@��3^��a�d	�,ox��L��:	%��q�֭߅T�i �f���B�`�+ݝ�G�9l|ي��1�It���b�Z�T"���g�{sr�5�A*aв����F�}+��u����O�s� ��=��(^�xо�0u[z�(��J	]L�ǜ{��k2U"���İ)Y�����o�*��v�=?�j$���8x#OY!�5�*�ã�O�a]0���q����Y�l0�h�z\�¨�:��c����G}1TV�	蕀.��Uy̎YS#���8�̀�)�F���5��)4��Ǽ��9~%�(gD�ȠeǺrP=r�=����L1��sedh��Lԙ��a�<g�Q�z-;
����'B�`�s�\n"�l�4s2�N[֖]�]�^�-�<��+Ѝ��v�&��e�ˬ$i)�Q!��0�E���@�n�W/Z}�Qb�6h�ދ��5;j84mZ��em�3v�ș~����(�A��� *eV�I�O1z�{s77�{��G�bc�P���s$�1I�A����bV����ۦ�;Ɍ���,79�1��s%pOT��S�ww�66h(��Os��|~?�X����-ո-��hMJ��^gć����;�o�^�XR���r�Ek?-�� -6�;>��`F*"�Z���Xx2����&�+&a@>�}T]۵�sI4Θ_U Y���|������+ex�߃h��zB�j�T�eV�Bd��0�)�ܕ4���z�1�!�>���Ԟ@�����������zV�I��!�1���2	���1�ѵ���@����}���L����nӖ�J�o�
��br6�IU�/��F�����Xh@gL��C_����D�(��K&$�>l*l�L����T�gc�H��5-o�*?�Ę-�[J�+�B�gm��awAJ+��J
�Z7�8#,���n�I�*�Ph�}�#*�0G��N�'�h"�r��O-�z�#�;�T�4#�Zi!M��Fg���=� �U�� �ۼ��=�z��8���r���XLQ��u�|ִ�UCʽ���SS�'�+�`K�i��R
O����;V��.eG���0U��,@d�1�c��`koO��H��
"ܼ�s�'v=-Dz�\�l���:��W()��zŋ�ֆ|[H�G���PjyKZ{<i�r�hG�{���t$�� ج����K���.�"m�_� �Ň<K�e8�O�<Nz�[�{	�n əaD�4�e�{j� {�=$�_��� ҄� I�q�9���"��������iQ�'!f:�a�����-��(,Q�L,xQ�:��I�Ë\t�3C������F
ft�B�);3�`x�M��@bf��F��p<�"����aګ�z��\��6Μ���_��]�
S'�o�iZ�r�.�[��<�	�ט?󙠋%�7�뢮2O��fWJ~G}B= ����AՂ�����M����a�aN�oKą��e)u�o�����;ў������V?j�{m�]r������3�t�I�T9��������UU��Ȁ��6V�(�%QCi`a[ۑ%�Hx]��嬜ڔ�f0����a����c�ґ�YB8,6�D��d��H�ſ������˘�2�Vy���9����*AEɎy.f'-��-��`ʸӬx�Ș�,�B�bF��Ϙ���f�^�"�T�x�V)��*���Z�%��*y"���F
�L��䈙�Hb���C� �2Ė\�&�=��aK�佣���?���'B-����x�`I�=�ϑͤ��;�l���G����w=��������L��3k|�TU����y�|���5{
^�vM(�+2M����f�M���@&��-���;bky=F�%ڕVhЇ^齹~�Cg�`K�X)D�B�CHI�V�6-���Kdui��&Q�#���q��f���Ɨ㨮�l�ߗ�+zX
�@(S���,��ֲ�ƒ:S�t�l�A�;Xh5���C���C���W��ڍ6��Ҩ$du����[ݙ�f�B	+h�l�`�#�V�E�		��PB����-�7��l�iHJg@����~��UFbV��7�Q�I(߱p
q�ݴ�f�
5ģ�~�M�N@?���e-}��E^_�2�{����-x�N��2gb�=��B�zeb�~��G�#� U�ɲ�ߩ^<������Vu+�{�T!D	��?l��Vɽ8�����F��0�5��}��e�~�6��a`�y���[z�3w�*xN͢
�1a׍2�H?F�S3�w׬jU�1?���R�]�} ��1�����h�]��F��L`!��+j'�LHܜ57$��}g�0ټRZ���u/H"6g#й���������%�,kج`;���QK'=�A/Z�ǽ��R���F�%��c�6���H�m��. ��qڪ���Յ%�zΖ�{C��-ҼkO$o�9nYt�E��e��N�s᳧����#s����f��ǜ�Z��"�6y�j�-coh�Ã�g;٢M�J��(��rc��������O�׿����"�������&�����R��lW�x�$Ę�64�Z�Pa��PeK*��2\��ϑS�ꦤ�b�`�U7����P�0c��a�c�|b�e?���g2�Iւ �왁u�I*����~��':�33@��q�v�wF�u�γƼ�l�F�T������V�������t�X&��:���s���{�T�h��ɰ��ryex�&�g�ڄy��f#��B�7��Q�&����˩���V9״��p���CC�8YB��n���ݛ��5՚�����1>��r@{�`��jS�~� we�z��i��D���b�/o麻���A]�^Ob��^QŮ�2�`�I�j��g|��}+� �|���?F�QI= �>+ݹ��J-2��T-�3~h\��ss��!�s�s������ÊR[�Sx�o����j��`O��v_�뇿��I���/�r�����������l_sR}I���%�Dɵ��~�xμ�%1�a[T���q�-tH�:��og�WG�R-�bBV��+?�X��ɾI��:;>Α�_]mw&P���)�z7��|�����xF8�H5#,6������6�Ѭ}��|=o�Q��lE���\��.��C�$���̃#���G;
���wG��M@�w�.�q�����`/#���A�2�E�Y�L�eӄ@���6z���wS��{+L�8ɟ���L��Ͼ:B�� "3�?ф��ތ1�J�kv�S�s��7k	�����0L^�A��9킩���3t���|t��+Ԣ��ti���#0F��׾��%J%ު����ߺ�/�iW�>Qj��}�\�&����{����kŭKz���Ǔ2�fN�]s�ؘ @��yф�Ƶ���P��n�d���g����b�6���R��2�.����y�T)Wv�
MB��2�z���=Yb�j�,��;Q�X��� {�_Y'6�ΝW�r�(��̮�P�%:Uޮ��QVlct$��	��CVk�*�f[U��xC�����PO~�}������^�={�o�a�s�mm[y�˦�m�m��Q�OY����`ӂ���d!��Bbm=� ч$Cu��b��|����Mϻ\^�ǳp�jr:8���6Yvjj\�Ր���XO_�-i� �
�t�i�V$�ҜeV�15�;S����Aޣ*��$�{�Jl�; ��;ã`�Ɍ�F{I�l�: G�<��p(� ��cߏ��oN��%���j�9C�z�gOrJôA�u˙���dSS0�/�5R�t�t�������S�D!�����XN����\$ ��\╊Q��RH�F�eʪBP���q�*H�}].��Ԑu���eQ����b��!Uc����k��jHZ�:{�?�n5���_�8��K}C�q��ض�*�]J��ʣ�i�8�4�d�������Po�Cf��q�����\s�o���x_bf��JsY+�q&Qg2#�Z�r�ԧ��Z�hqp#�C�Ȕ��蘰f6ψ��%(��@躮�XKx�\VdG���Xr *M�>�Ⱦbe%��A��o�ccG-#p����u�����&�1�~��}-�ǳ���rEHc����J�x�S�6� <ae�#�@�k�i��D��:	/���,�+��hq��:�<����}���S��)X��F���aCɬjA\�GDh�7C�^��1���-|,��P���	�f�͋�|���!x��VO�y)BUY�~������%Լ/�µ�=�2�;`~ "��mANa��0����3Ҹ�('5tb��y�)��������x�9x��oĳ�Y�U
�s|o��l���A�`�(�c4����)�w�5���G_6�j�Rh�Ҡ�%i�
Ҙ@�X\ˉ�<����A��N$bWǎ��p~�		NW彃9��Xl33X�D�s��n� 8�Tg���=�5��<gYh�_��S ��x^`?-`��ZdBx��>�Sr���fz^]%���Ү�^��� ψ�Azά�BN�B���
���wW�Y�۽�5�E��.��������\��qԧ�p��|:%�(jP�@U3�v��M����[t/��$���mp�z�lF.suK��H:�	qL��
��C�#��#m��&��s��P#C��87VHQ��+TdV��.�v���s��;�v��r�Z�9�t����v
��W�68Ɩ�"��!H��0�T�����Z�SM˜�ӧ�3�շW8��е�̏���TO�����iN�V���;���$�]�xdC	��)�XȚPo�t�I����[h�lr������~]�=@V5�H@�:W��s �B�r�$���&���m�����ǹ*ĭy������7ԧ�)�D��I��v��0b���~c ר֎���B��1�^j��W��v�3Tr?�3�sy�>��9�(J�A��g��l�zkU�(C�"QWR2�-�o��f����������l��Q�_�}�<j��U�@�L��Jǐ�҈y� ���/���U.t*ر㎦�����sn粙 V�גr�FvWk��aP��h�(wH5mx=KNц�B$��vur��S�+����dT���R��� 
t�uRL!��^����_?]Q+���k�ֻ���`�ޡ�B����w3�x͌%	 �T��G�`��S��Eӌ�5��(�d1㛵G���m\Ɯ[�������4a�'O-0=���'���STw[�=�+�"�T�{/�_o���&ѿ�.����:�eš����6x>���vZjeذ���03=��9�B~Z�4��*9�1P������J1cQ��V'�������j7�b�a�s���1���Dt���	@�ʄ�P9�a�iK�Su5�4��W7E8�TO�X�����_=�Ω;a�1�f���{�Tb"�0���ֽ˥.λg�8��,�U{cd���g�| �2�&؍Q�Log�h���a.lNj��Pe�_.�S �TW�v�N����X 4 �OO������/�g!���f�)訜����.�}����C����<4�L���g m=� j��>��-�p9�<�Ϫn��i���ۃ	�g-�NM��rc�/b�H�}�ta���V��aX��vc*���M��T���oa����MU�c��V��Ve�[�Cf���y,޴X5�1��m|@|K7�h5&UvZ���{�����c�����n���r��.��4Y��u���r��-��bv��s?�=�;�\C��%�Ԃ2;���M�}1eؖ�Y�c�pG��Y�X�[�c�����b{_6p;�mh7H)�zFE].3AiKP�m.Ȅ���-��Bbp��E�3��Ȱ��k�Ac^>�<,nӆ�7���d�S�y�߄�u��	�ZڍC��F�8�<�KSg3����YVRUв@9j�:hra%S� S�T���z{�n``�*��&� ����4�Z�MI���!�!T�@�>�ΰs��RÀ>L*{<�nD���b�jۘBL�K��"9[�Kr5��+\���s��g���`;��3�S��p�Սi�W9�_ѦH�B-�����6v�^��d
���G{ثA<p`c-�b�x�&d�z2FU$��2=ӄ��(q�M�t3�.fȎ$}���vm�3)u�v�Kh��q]�t~��I�'�F�@�_��Qf��vИ���e?g��I�#��!�̴r�C�Bp��Q{?�!��$*�{F��{`s�d�+��l*)���ZF�	����A�1���)�о�+7�TaJ��Y~�:�:�Q�*0pV_�{��3�'V�����i���E7m��������[��rMd���H���'��Ӧ��=C����Lc��PU��О=ԯ�����U��1��tAe�YTD(�@jc�{(C���	���db{H^SK�>��/�򓈲E�X�һ^#��4ML]!D<�U�!L�*�%p�mے���6�&3B ����f�YMf�á�͕e���>�bzڱݡV��fatD�P��Ib���t�j�c�!Ԯ��l��=b��KA&�@���;�[��%
չ3 	!7��x��U@�_�NQ�m�+:C��	�˞_2��o1�1������_����{&���J
d<3u�>0�9ɐ����sHa;��<�fC5��#ưU��ܔ�U�FS�ͻ�)n ^uF�=�~�*�>}�K�xX$��
U���3��m����*�5-s�>"�deo��Y�۵j۴X?犀n�yli�
ݳp��^�%;m��c0�1C��x��$@��B�'��Y��SѮ;�Z�%�<c+�%�-N$�.xw�8�KĂ�)9|��k��0f�zrRH�%zw��Q�^sh4` +K����oI��/��f"Z2�M5bl�s/����� �P,$����B�~a�D=���D�P���npzҹ���s0]~P��瞪�)��έ%#��)�*�av����=��]��s�4m�*�� -�6����xK�m��(8�fh(0���A��Y��R�����rc?�[�������_b�ZnvS]�J��9��������zH�(E_#Ii[6,lb���Ü֓*z���%��|�9z/E|�p�z5;���jɣ�86.��*���qd�
�odS	u��3�\��6�(�G֔\�|��m96����3<Ƀ���<���f�A7V��4�L>9����ʩ�	Ɔ����'�@�1�
(uA��I/3�Ia�hPt}��fS�( �5��B�M�"�|u�9���0-��s�b#�`��y�����8���萴&C}��u�v6˼C@h��v1T~c��P�R2����<�l���.ծ pV�W���ݬP�6+�X�l���ﭴ
�α�{&{.�}^��۸^N�:x'h]hm7���~�I�O�d�#�z�}w2i��v������ʧM��^q�|FR��c�����Z�X}� �c�����n�Z �wc�w�7�����B8x�,[�U�>RE[�4>����Qm��K�*�Ɉ�e�פPQ���8]>���Z�L(1J�s	��\��u����;4�6TMd�*ԩ�.�j��lf,r��}�y����^��m��3(�t��6�A�����Q�s�@Fv�1�y8R]>����T�1��'3_ܔ>X0�
7kɉ��ywεU5��&�m�!"&�dsgYq1ޗh7a�1�J���ʞ8���Vf%�&��������~�.�o�{\(yش��e��l�HPX�#�S�h۵Ǒ!l"%�8d�Y��
L�$��1R���>�^�x�|���b��[������������m�E6F�0/����V�u����YE�B�붴����<;��-j�*r�}�p�����ZK4e���n�7��d�L)��.���+U
��*ӹɸ��Vrs�9��{�H2��cǋ u2d��,���k�� �IA�E��TZ�#f�d97�={
�0Ex�����͛,�f�>���p��b���z9�Vz�脣P��(��Xh�v�x\:����?mT�c~Q�ϲ��p�kZD����4kiZ�@����-�ԏ�V5`�����gOsJ�;(O��/�?�6�{fI9W	��]���v*���]oj�6����8�bd&�6-�����������rcb�ʋ�\j�i�I�$�Enq��^�C��0��	{1����M��*�~�.�?��@����D�@l�D����֝䎂Q*�8����������Ϊ��H1�Sڔ���#�s4V�wBsp0�q�	J�akY�ž􋬵먧�L��#�զ�uj���[
�$��/HJ��⾡C5��ݎ�#�� ��BoD� �Ղä`�����#9��Vx.L+��y����W�jfBH�Qг%M���kz[��q��K
��e��&�px��"1�O8���}�wA��-����!)���)M��q�\Z�s���TsuVM��d��&��9�*ZJ����� ��q�[~�z��TץA�7�۹ǉ�ܤo؄�l:y�:g��Xm���3��W�r����k����rC"g|���ɶ���M,5�d'��,ccܹ�I�J���"��?��ΟP�X-vM\�ʄ0�A�pTqv�W����L�oOr(�#�7��y<�.�.��0	!�%��{E�`�DUaUC�n��l�s�T���iqb�
ķu���+.[�ŗF��D�'Z���w٣��T��i��$��w��3*`BЎ��t��\/-�MЉx��nnib �O�x>��װ+c�����ѣI��K����E�(��:��6d�]ӣJNz�jxM���Ԟ�Z1�
\�V�d �/%���>�V1���E�c{�Q�#��0w�/��LO��q
o>�X8�]"����a�8���%J%�՚��Uz�ƥ���<������R�@93�����TBZ(Ũ`�T{ْ�.�07/ �b�L�`�PF(��&M����L8�I*o=�փ�z_�v���sO��>�A��e��A�=6S�ˮB5�|r�d�V�!4!��4�*����%�o��ڒ|Y�Ghf(����f��6�n��I��6ԝ���0�}�q��r���$�����¦��2�����Eo��	�p��HA�/����g�},-�ix�3i�0�\�g���b��b3�:��%K,$�mj]�V��L�,�s��=z�g��D�t�y���>%b�E�!@̄r�l��s�<|���gڔ��C(�\w�ѯ_�S�s�!*K�>0��{�ƅV�fWьq'Cd���njo�)Nzfن��8�ZT8M�J0v��0��=��N�b���ky"�P����ƶڻ��,�Z\+S�7�:%�K�q�f0��7팡��h�6��q[{h�'Z�x�&~�w���{���L���D{@��� <q����ٍ�?ec���@CGԴ=�m8*jC��c|w���ǿ�P�������O!-�:��o�*$3t���&y��o�������D� �{nv S��l�'T��k��|/L�B��7s�z,E=Z�	�;G�Α�	
4wKI;��##Z<�4[�$f��|�����ג��a��)�P�ܭ=ƞaF����9��zCh�`�(�2@/��C�{���c���T�Z��#j4�J�p�M.�~~@ �f��L�:zF[fq��!F���D�n���z�*`�traЭ2ّ~1c��n[��Ϥ/жx,�%����D�V�U�r}�kj��UX�W�M���.mt�}]�L� ������GtW�ydf泏'"�N%g('S�o��&c,W��[�XS'͑Wf������ݠ�	�"T��*?��Tl��\�ʉ��e i��ˊ:=�ef�2+	�BJ�M�4"�g�0&SCR�)�i�Be�w!'�M��D�T#�'�lR�ہ�Vj_�hI����c��.����o_Ƒ�/­�;��!�9�`�q2�3���v�v<W����x[[穑1�0߁@�ڄ۽����ƚk�K� �Ƒ��8����ct�b:���6���&�Y����#XMP���C�MM-h��ϣ���`v�[7�w8%�@��}��5��Q��2��r#���eQ��&�����|&��Z��S�ߠ�svޜwk5b}��$�J�^�Iy��k�>��eor�+�L�SÉ�� �a�sV�@���]^O/7��dt:mKк�$���A�>�ڧ��Dᑮ�o�R{��B%{�����裸�`51�
�^0�6�Z�x�BB,�Pm���ϰ�'�3	�>����^�2'�v]<��h@��0A��.�0�S<��N�J�-!�2c�є����S�C�M�����%���n~N��vJ:ט<#�Ӻ-��*j��.L�~W,k,����\I)Nw�44�ƃ��F�ן��N6�|B�n�
 ,�R������l!R`����r�)-Ju����_I{�um�R�4��Uh�5��Wc�:X��?ds�7Oc�`��w{�/_>�_��Wc��?���}����3�ώ(���dFe�V6U�K ���zDB$���MՏlh�۟&��5���S9v��>���=�3l"H"d�I�b��&I�Mb+ƚG[~�y��ACh�1y���T��V-旑�5����9$/<�=$�ޙ����G��1�a�Y�|��ފ��m�٫�?�4�v<IA�-|�����o�.Lǁ�ؘ���5��6�����eO�|2i�Yo�1՞��N�h�j/�����P�4���l�,݉�*�]3��5W�!ñ5�`^�fE��1"��h�?LZj����`��MH�����9����.�U�	��N�ׯ_������o��K��M��g�x�~S��E�l�筧֙�
&�8�fÆ�{�f%��V���b#	*-A����*<C��=�&���d�$}����s&p@��k��t�FJ�*RڗZԎ�J BVw�s���A�(�����/rp��zK��f|`F̘E����.zd���mf�`��n;���}��]�T�X�,� ���f����dt��xl��]6�N�R�,��g�6�pr���-��K��0���W�2T��SU���S[4�0�{��o��;��Z�
a�qn����YǷ	����*�=�<�qKhH(`�sG��e��,3Vi%-du�׎�?�xC526�(;�Oʟ�|���bR��uJn����^���j�6ۓ�=��ç�9YϤ�ʯNU/�a]�����y�0�^:�Q��$DJR9��\L�ɞD��vs-��v�S �\D��6q2�Y��;jq{�ޭr�s�Sի���c�!�I՝噕 X��3����A"�pږ�R!m	�
�Ea��4Q��_���Nh����A�X����`\�(�c�V!`�{x���������6�hO!�A�`Vq������xA�~~+FL�0��N�̈b;����$�-��5�^N�6W����e���c<��� =j�A���n��jw�#��K�-���=�[C+rMo�g8�,��Ѕ� P���'���C:z�񴮧3�K}s��P�/J#��t��t6O��ɻ9K^n3u���.��ʷ�{�+a��~��ח �Ѫ��(c�t�,H��c3�����6"!��H4�y�^�����*ŘPJ�blD�gb*X^;g�G,6�*�=y+�?݆��Y4�qڌ�D�Y�(�0#Pm&2�#���
��*����'Q�1���A��;�H��/�/֑ޅ�v]�tDɊH�b'�MA�z���a���9�IC��k��s�?͢9��R �
�$W�ې�(&^ڂ�nhk!hB��
 ���ɵ1�� z��LD�W��g8t=j�`��y��4q��(^y�s�i�*�n�y�t��j@�]k��}��=G�`���_��̄���_���X��y*b���̟����E�Ү�����[����P6M7��Xp��o7)�.V$EQ��6��/��;i��3
�4R��I��q�)"e82I�j������n�mA��F�ql�"TI�b_�����Bh����N���FfDa�ޣ�����E(�?C�)
�p�G�;QV�����=2rz�:S�*��m��Lʖ,���^��HF��ϲ���Ÿ�wH����X�9*�!�@o����I��J�-8j�#�@	�*�m�ns0��	�z]�iT�5�,��B�84.V�"<��Τ#���q�PG̱;�|"N�f�\k4�έ4�V�Q�(�,y�-�'�
��)v�E�%2jiD!�	a�ӱj����w/�t;O��_@�W����Oϫ�/���Ž�ׇ�@��v�W�h�*S�p�C�*In���_n��f��ʤ�y��m�n��8�nz`�5 WS;!�ň}`��y�n@��w�A.����a�nj"P+���s`d��-�����`#���	1,���l�T�?�/� ��w@�@�@b��ñ���lF�t�̾R����G�"��*�͌�_0 � �����t��;#�]��������@�{��V�]��*��F�y�"?��V�M�^�W���,aO��N��:�FGW�_�����2������Lj{~%�˙n����#yMԹ�EO�p��u�ۼD�X�uBG4G���6����8TV/����ۛw�Ժ�C껕�R8ne������]=9N�ʤ��P�n*B�`���'����q1#���;0�#3�q�aD�t�;^'���?�����ױ�@�"�os=nA}��~�N�Az�N9������k���
�����t��`?���i��}�d���]V��u�}�]���9�������oɬ��Y��yB,,~�j9�ܑ|�`Ӷ�Hj7�����Q��0W�92��P�=P&�}�uX�ބP�xw��o��!��0%�uJڱƂ�l�}��������f~�]B�}<-��%���B>� �U�iqZc��k�b�I��Y�ۏ3�k��K5�Í�&����/�F��ɔ�߸���M�ο�X$�x�ܰ��f2]�i�`��E�����9���Cf�Ϧ��G0J0�R�ټ!˳�lm@��y���屧�u�-,��4�L�ĄV�YϲwcL�8c�����%[�0����V�
�g8�u�ю��Hr�:���0:�4O�}=¼����lˍ��<+��>��x�E����>4��̬h��֞�-�G��p��S�-+���E����:���*��{�C�o�P?�B�ۍ,C����s�ַ(ͦ�e�t������c��B(�p���B�CHU�� @?˵"�p����x����=�S�%�z$���#���Ah�8� ���#�q�~to�g��.��+d3�]�s(1]'Q��z0+`)~�m��uS�����@�yA4��3��VF�
��0�r�Y��N���!i��d+�?�׼�%��!��)�T	�l�3=�����F��"P,8��?'�0�����:��7>�[�3�<�x��/E��R��-�b��]틭Z����u��q����ƪ�.V;U�E%���2Ģ��A��G(�Pdkɴ�x����#X�1ڊ��w��[؈`�����d
Ta�3#�[4+�(6�:�՞��]�s*�9�����	1�dic��r�C�6�-��$���9����#��K�k	xyL�����ga�a&$�4�D�j��4�g��V�9^ZEs葎�N5_K0SC�X;r�,:hXc�1���v���[�{��[��������xC�#	`Qbb�`�~�gu�-Q����fZ�V7$�����&#�ǂ��J�f���m�E};2;����������ʊ`q<�C�Z��Xyc��~�~�� �Ŗj�l��CF�LzA����]�W�f��bF����o����6x:��Ӌ�8�:3r^�a���y>2�ܼ�1��Q������q'ظ�̱$ Z������Av����B�$�=��Q!��L�"J�%�R��`�M����Wj7P�)Lo�9�s����D\U�+�F��߁fb6����A�5m���l��<�x*C�NJ���e�/��� �k��Ѱ��i@\Y����OH_�m���u@�G�d��2�g�6g���5!�)t_�{a��s�Җ�k�PwvC;�$[�G�{'���ɇ��JU������ILuf|��G�:����(��\����Ym�Z�����7�k�wPM9yd���lS�P�%߇�F���G��Q<�1���q��F���L!\�Y��_�(���[;�kFM�m�����%jO�j��rOt����_Y�W)��*IχM�Z������2T��A�T��E���Ơ�+fT��أ[��sTOW��P�:���o���B�#�=��Oz��<&�H4�����|�7^	~a�"9j��[�^�A����1���� �C"S�;Uf(�`	�pf��;�I��8w����=0] �����\�=%�4ց���Z{�~5+�]2hdL�U��<"y����9���w�1'�Ě/����x3���y�Ƙ�бO0g�EtNIg�q|�yW�z��c���ؾ�|�.-�f�L0q�b�8�
��b�#��;�(O>��Pk���@������'���f1��o��N?�ꔵ���x����xQ-�G�/D,t͑�.���kB�|O|wDw��4�2�.������T����31;9O0/"k&����`��Ӏ��9�J�x�3zVn���e�?��nd#���ֽ��4�Ŧ,�'��GJ�ǌ)�n�q��]�l�
Si^��53��>�%5�4#D3B�߲		��XX
�{Y���7�<I�345�._���u�;��FH9R��� ú6I�5:�{����`�ǵ|��\�J�tL���P�a!W��m����o'}R[�����Q�rC��k�^�����礣���k�X���7y�l�����c�G?z.�X>������Y��8	h�����9D�����z	S*;�z���c>�V?B-��������N���ȸ)�bT����G��Fs��̿�<'&�4�qެ�'�$h!�=jǲ��($�����%	AS���4�Qs8�֘7�Bљ\�(p�댽�eS��xwjQ���0����֏;{7�0��8G쥺�7A�MIC�����*�ќ�i�����ʈ���tЙTy\�O�9u�2c���;��ʱ��������ϙw��(����|:����!ʯÁ}��}�L�Xr��C��db6Iح��w�ϱ�\�>`��꽔sCH�3������>
�0��xE���.s��4+c��Z7�"��D�b`>_U�"��nxF}��FrO?����j2T��,�+��tODo�]aYYR
�F�t� �*g6�9؎�bb˂3�̰��Q�,"�Vh�Sc��X1o� YA��& `���3��W��h}���0�SSO�Ӗ��/�G��f�����*�\Ė����^�O����M���낼}��Ջ��.ݔ�K����[b�H�-��{iQh%7\��&][�Ϳ0���)f�`1!��0�'�H]%�g�ji����GS 490�c���I�[=�-��r��c,���_r1i�y1+qU�P�+z>3����fF�?֙�ޡ-���"���dz:
�@jo�sTV���*-�V�y�O�}���١յ�nk�6���G����Tf��&��ZJa�e!��a�$���Z��=�?E�	=.QuL�=�$ kݲgq��GfT8�Z`�|)j�/_�9ޒ�iD=��~
�TA?�n��x<�����jQ�L��^#�z�w��0u�2^��h{�{<��-l�����p>�5%?��%��F� ����=���Ẽb�D�w2:����q���m Hvp�րg���b��K:��d��� ɽ����Nt
4F�Ȃ%.��B�|��7͛�/�����Ѽ�G�q���x/��#E�L[���ڦ�Xe`*�����B�
�3�D������&�2$�-h���<��a�e��l$��0�i���
�У�iP�֭:V&������O��/�y�1�v<7l*(>5��i �ZF�<[�~6��p[�H{ǰ�FS�?�,�ڠ�	F��p�ad�j�MUs�Ck�w��J�X�
�����9�D��	�S���#��jc��a�V�!����0f~7�L�{p��3M���}��y�L���gX�����h���q`v�j�z��5ң��(���(�OR3{�d��8l="���	ƼtCC��Q�}xI/6u�s�c=��,Hԗ�4��tL=�Ǚ�a����^�����쨪�&��,�[T�������i�H���㩙R��؋L�6��PE�Q�rS�O7��!"��7���L+�XRE�h@�#����z�TE� 3e��bb�!&�,BY�]�e�B��w��o��L���V����R� ��XO�'fu����'�ȉm�@N���� �Z�q��|������\3��4�l�MB�nn��A~w�e#��L-^}�!28�~\��>!Gs.y\�v��I	�`<TM�����@�G�奔��I/��V�j���G��;���s0�J��e�!����u�`boHn�C���E�%�Zo����W����Y5�(ş´�Ê��K����X����lD�r��\�Y����61�:�PI����^��؟}��YH82N#�;0��j!3�f�l�19@f9M����p����&@(1��Ʋv<�sTap�[��;b|Y߀���P��9�4���Q���x_�25��=�o
�����q}�������ݽ��KMW|N��MUo�g!�يwm�[���؟�8�kZ��2������ {n�边1�S�Fq8fM��
 ǒ����3� �n*��z6ț׬�d�N����ސ�ke��z��6m�;�t@$�p�c��v�V�B��S�;�&�/��̔�U&�7W�������S��m\����� �9sSa�e��,�'TH̛�W#���L�Z~����լhGC�q@���=鞌RM]G��i�87��fj��<�u�E�ѻ�3H`�z�7Ơ���&�4��IQ<��Ԣ�9�]���9���֨����=��3Tܛ��.к,5�O���V� ��a���S;�L�	|&R���7̗~��|�*d)	MV"C�n�E����7m�$ǱAUs�Ȭ�s�WfegDvV�����/-�[]��nJ��x�#M=�,�.��0wӋ�� ��'Q9���z�/��~��1+���X��wl�f$�ʥo�>�	��d���2�EY����4����ֻ����-��"��_3�>J���Q.���$�����|�o]�2�E����Fj?��.�Σͅd��m��U���T�zO��K�%#(d��7T}�V�)3E4������E9�^X1P� ��lYϕ�s
Skn�����Z�
2�iv} �4�L�ԗw���_�f��O>����r2p9 >�A�^;)|Q�{<~-s�{'�q����i�@K�S�1����I�Z�gq׎���}G�L��[k5��Z���@` �qm[�13Cߍ 2�2�r �aiפ~�!)!����[������(��7�4��|��E3��c}����:>�
�Yq2���̀v����5������AN�;��'9	Y��������DJ�#4�P;���&��^��FP�1�V�F��Ms�V)�u��6����A��瞌Ż�]!�~O�w�@����F�$�ĪKJ�r[џ�~o|}x������j��\�:Q�l�=��Ou*�ڟ�wtD�dҺ������PG2X��0�0��
I�f2 �@m-լ��4h�����ێ5 $�*���Oq�Nm�1��Ll�'s9K�$T-��n;�lx�	�uxO��H�_(g�vi�s� � �V�V����0f�A���W�+ege��g<��N"6k[K�8kw�{�%�^�%��C��&��ڔ��	I[~�4)[�?�����2н|2���o5.!R��ֱ�c�_��n�����`q嗽�MQ�}�K?0c���%������� ����^WG=?=�����'�N��*ǵO�(�� L�Z��R:�����300h�#�,B���@E����}.��{�8f�u��7�֖�Ƴ�E �=\fފ�6��O��SF@̘�R���}��ڌq7a��'�[��uQ
h�S����oj��9��6�8���/X#�M���іvD4E���ܟ��"9��[lm��"B-��`��%�g��퉊�R۞�Q�\��=�)��RwUP_��ǧm�9F�G���c�Ɔ�QG���d���L~�֮.�����N�,'�n�DW5���0ѡ�)�V �{�;lS֬ G���<��]�dCN����VF8��-�֨�YN���0)Q�	h����vt�]K�]N�=#�˛�-�)0��)�W�� GL��w����D�ԶV�D�v[�e���L2�h���u`E��t��4�Q�^i����$�k����!-�K�3�'���߷��$	َ����n-��P��E6�O��<�L�8��Pp����#��n��5��J�� `��>�V9r�Z�h"6Նw�l�O�`:�k�����PUt��ņ�w����E���g�x����P��\7�e3��y�@m��| "�(�7��:؟&�
�h;��Ŧ~B�u�cnqO �1��`o<��](����6�m��C�o�ɪX�f�C�w4����KO�.̡γ�K���hp�����d� +|����SK��RP&�`��)O2�3�{J�]f��*�ʐd�C�@���"��`C��;���[��o�\+71�Y�s�)�k;z���V��~f��W��Ɲ`l� Þ�4jX
������PEr�O����\V���r�ɻ2�����EtA�F�;X�wX?�r�<���FZz����ouݲ���;J�
�1��ۍ��T�H���[��w��F`Nt�EQ��"���2�<)�����>.�a[��5בZٻ|l�bʭֺ��z1���XƠ77R#�x�*p�]0���
�xDֹrhj=8�b��O�3P�-�(!W�E�x�6�?�X����@��H�V�,`20���r��=Y����H �3���g�[��*�G����{I�)&C$��E�^K+
`�L{���Jd0�T�h�\p�c %�� ��oQ8��z&��!�~ޥA�7�ҭ��e����!O�����7���x1�*;� G�
���E����٦ܤ3�
 U��T&H8������Z��~��b�PL�/��ɦ��Ŧb ��YC�w�[�D����`��C& �%���C$�V�7<�XFp���-rN� �ȸUf*��{:�����-�^`ΰv��hL*�i�rU6�9�y����O��V޴e�`�,�ˁ�F��������q�նX��ʄ��>)<n�2���(B�q�@�%�h�� �>O� >����̲=�����&�)�&�v�C���*�p��u��K�� }��)�h�z�u��KZS�-A2�}+vkq���F�`yx�])��GyE�\�u歲Y�$����9��8^�W�y�H�ǫm�䶔������WTe=���F��t<؇ھ�7A���"��Q돓 B��N�z���ec�,�7�>J��ĳ�|&�D��4؍�n:���<��qO���Tl���w�b5> n��e�pzrh�i���2�m�u�p�o�0��G��"�P��4��=��QέWZ�������[b&Bmπ% �g�<=�zP�|�M*���M�1��0���ց���S�vMfo����KC�5�[��� �}Ꞃ��]0h��m~~d7+�k'��7Y?�d�Q�N�wf[�  ����RkU�5ν��0�:���Z����(�u�;������'��p�X���t�98��3�4�^/��d'd���p~/�/'��?)�ټ�^�%s�u쉠�/5wh�-Ι��;��	+���F	 N������ ��]��{�I+�3�ۿ���:�&��c�Zi�㘵��hp�����\3,��Z��I�Mv�\�	�$�}:Y�|����aWKٓ�M�-ӳ�v�]b@eG�1��\]���.��y|�DDƘ�g����+�N05<����;|�b�Gl�����f4'2�Xt��C]7����9��M��鎌P�*�?;�����ZI��X�M~���%�M;4.��,�o��ᬕAe���}fQ�Ҧ ��� 8�A�
���;��D3��9]��`����&v97�4����2�ao��$�yӷ��Y-MH|�A�e��^D��"��H�¬9AjL���v:��ky�e%��(�Hƴ�Uu��lyUz{N��n��SΊm��̴3[�db��������tM��z����W�~1mYb��d�ɀ�rPnx����g+����i�*qF��?��������]�z����.͇�w�ٲ��L�-�S��2T` Xِ3�w����e�;L"��� V� -;��)D��E���BG2�d�����&v����)4�X���v�9F�K��1��4��2[X������P:������w�3�΂٨��Z�N�" �EAL��2)B��	���8a`Q��ދ5��S���\UE��`���U�6~r�{j���k�*7`���`ڻ���US�кD���Cū�.����Yx����.`'���w����P�VT�DZ��q��p����_0 b�<�u�؊�1��f�]V�A�Rm}-�x1�͉0�$�/��WK���z2���t��ܒ��g0����m����k� P�g��/�a@��l��
z^g?h�����j�1��*A�v��0�򚼾M�����#�!�(� #�a��%���*7����>]"'�IfS�.��1�Ysf���T�q�w})�s*Ѩ�M�"R���'�30���',𴰠��l�+@��?혌��v(��p7/������] �k��FoM�Y�>t��G��ܯmk2LҌ|����>t�$v[BR���:�=eֱ����Ɉ�o�3�w�l��v. ��b��q�M;��6T�4��;���� F�u���lW�I	�`M���^{	 �׎�O3'(m�����"�i�KXY��d���	Р��]N1�}޷4*��Mr��U�3����CF�����Y�	cN\�/�o�jQ�Q)��<c�Jj�ű8o0���'�=?������?1!��<}�%�N�u���m�����y����_�������7;��; Nq��`� �b�.�|C �j��!e&O�X$3-h���>Y�ȇ[K�53�;v���& K������f���ğ&t�l�V��=� ��X���D]�=��\����B��}���QC��2b2��X	�rZ���O`�:�(p����.�⩏����\�Ʒ�bL9X-���.r̊tʭ��O�!8����h�1� ���fb��M.�3�%��ju���O�q�f�.[.$l�.9{�{ #G��÷E���O{�����r����Z��1���ƌ٦ZQal1�flF�@j$��!���`����X\i�ü���ϗ��@�@m�Yv7�갆�轶�]Kϭ���Q�l0��j���J�I�����*��i� [A�9��^�2��2K�@�&�F]|Y)�&e�g��zD���O�9Uq��{1_3=W\)�1Pb�k�۳BΊ���3�����u��I��#�qY3(�ƨ1�ST��q��K���[(�d���UuC�r^��Qɢ��!x���e�O[xq��c ���ɻ�@��oU��j�w�������o�1��^�������@i-3&Z|�zTCJ��r��E;��H`٠�z�C]���l��9U���2�uǢd�O`�� t��x�	kzN8k�s���S��3r���i���z$c�2k�j�~%nEBqg�^~<��6��S�9�Q�6�"��޵���#㉹�0�� )�� cjGza���K��dF)�T�'L����xّ��s�=<�E���wV�-���YX�yi�ڲ��Nr7�-Zz�w2yz�@Yd,[� \�
��4d�B�������>_���
�����2�=�8�����p3����z�O7@�W �FPƪf�L������̥�H%g�`�� ��S��Ҽf���gґ�������d~.bb��`�cl TKge�2�i ��b�CdV��ic~6�J<#��
���0p#s[��?�\�a�H�/����X��%�����t��������Ƌ�և�¨��-�4�)�AZu_���@��J����ב�B0�(k	���h����t��6)��Kfl��Q6}��mTm�"�j��	��=���K��6�/����CC(�P��Q�gf����l�K���u':4Gd�ǀǡ�+{t���2�{���H���i�Rl�­��,��Ԏ��ކ$��O�z����/gv��P�^-���� �Nޑ�&�C˚��Q�x�� OA������--vG�z$��M9m+�������e[A��|�`ZM����M��^r��!�i�a���ؠ��p�Ȗ�^"W�wZ��ϲ���Q��]�=��bnۼ������u��^�J�(q�#�4��-��?ͺ��.`3_*a3�܅`m�T�B����[i,�c�fL8�k��s8ɸ�RtS=�9�64��۾l���a�Pͽ�W�rn<��]`t阱�h(h���_��_��zr?��k�?|�`����%߹�V��vmHc���̰��˝� 4�����g��L�B�>b?e7�,o@1;d�����`�о����?")�iO�������Y�3gw-tu��s����`��k����v����X��9�0b�k�&��waHZ�xͼ>cw+�z�
����R����Q߻��d[:��׼�A����Gkol�zry0Y���Q�BvF$4����ۈ��'e��0��k���k����=¯��6f8Y�ʤʌޯk�5��k�K�j��"ë]�+� <���Ɗ�=�xX�>�A��<�RG.�y@64	���}�{�0_�R�#ˍ`^�"W�O���9�ڗ]??�^~���|����|��1� �M}����~;�%�h���'�Vp1�D�4O���~'�?}�O7�_����Z�8��u���.����A�蕱�M�D3�ׄ�ff���lG������4uA�-ٔ�Z$Wix�5�c���)�Q�
oa���������a�)�@lqu	`�M���6<8��t����6��WD��з�m)�s��7���C���I�U(�'�m���������r��038�Y%F�z�r�F!OVOu�ȞTj��=1F�#/��	
	�m�Bж���K��J�\v�+Rl���Y����`�8^JD����3u�[n�V���
�{��r����Z��70�駟�_�/���Nf�;m�'	D 3Y����W+��S���u��Q�><��T�4���곏��fd��߈=f��B����qy�LL s�̀b�Ȯd�rL@���#������ut�Y��'��0L�'�������F�=�N�i+6���6�`��]�	�[��#32��H�����C��6�
�TQ�TD�k�L>OE��:R����^"��t��^m�u���!����2m�A�bJυi�	KL�Z�5��I�G��>����~�muln9j�JLeėh>�X���� ʓ�D|�@��M
e	��$��$c�zd�!V���dۏ��E�)�y���H+��r�en1yc���K�D��Տ?�(?������SǑZ:ۍ]�5c�0�A?L��{�,��uLɉ��~������Z_~���z��%�U�f�_<��эYKm8ͫ
�a�3o%�Sd�cM��7i�~���`��ɿ����X�T}����R�L�&k�$pp;�v��J�� ���u�9[�|�	ܟ �_�TRIրxКq%�Ef	��W)?�}�"���[3�]��\�YY�D􀸩8�/g�"�۷wA#����y����&�M�����E��y���00ԉ��t1D9�H� �zk��;����l�9h8@�Y �2�y�)�^��%���{�7�C�D�0������8o����T(6.Z���� (�u�-,����U)�*�� ���}��'>�x,CM�)s1�{7m��/y\z�j��?Z��(7`��9(O�p��ˋ�[�s16����X�#)�w�Tb�;�5�94�A[��4 5P$fQ�>U(��L���lD���{�k��
[!���ڰW��Lu�v�(s�A�%�޻|����=�MLJ[�O�D��Fɜ���Sk �������~)6������K�,g����ǹ�.�����L�l=��}`ma��ǧʻ�Գ�Ve*B�Ko5Q���R��vL@\*��.-X�Y<� <��u<�ˇ�:��}}Ѽ����H���s�{����_�"���nf��L�y����=��*���2�͟�U�L=xR�Çg��
�zaR
�NU��ٝ�,  俑�؉�=�� >�W��{|#ޕ3��~�΂Tۙv>�Qp��bFu�k]~�����Ͽ�kL8���8E�h�_C���f �R�a~�1��G]20��� �Fu=b�'�ۼJ�M@�&����I�`�2·z՜�G�0Σ}� ���o�ư�
�G*eg��&td�9B1`��5�!E2]K����G����
P��[�m'ś�d��-�7��!�}FiuW�߶��|@y#c�o�rM_#�M
32���ǋ'��v�P�j����s�b"��@=�-#���-�c���&�p^��[D��j�mQ�n${�	�n�o����?�Q���?��~�Ӎ��NfHf�͞�wy��.>T�$��6�D"�1���/	P#g�L�F��&�	��r�F��&��_���iY�(@dF�kƅ���[�yY1�d��0��	-���3�T��׿&y��G�m�#�p��[��=?�W�;����(W��Җ�,��1`�x�"}}Hл���V�+(1;�c����D�	��C3�Orc.�mL;.�k���>���K*ƙ� 4�e����͔��Tq_(�c��n������	�IBӊaAi�d+&�%,��}��po �n��D�����r��[={ж��`�0劾G�VZ�Yv��R�k����n7�e�"��ҥ�y��
�7V �
�����At�,��2����(}�+���x�Z�!�[鉝l㻣��nbW�5���L=�=N�����>%���,��s��fb�dZ��[�#���!��u�U��-}��Y.7!�=r��{��x���ۋ�X��0H�|��/dM��~:hC������0	1���9?�>^��ۜ4ʦ��P����.�$.���*��)���-���'V��?����>b��7���Bv�:	��A��> �q�~Ы:M�x���4cj�}�iԘH9b$�1��IW��t�^#d~��;�c��OX��{�T��8U8��l&7z~�2�@ 8U#X���[�3�"�%���� ��X0ѭ���}���-A���E)�:�ź����PaΤ9�NZ�D�M"��VB�{7Vb��n�x龥���1�þ�
ѩ	�|�	x��*���x۠�R�u&�gQ�ıZ&�Nˎ ^��;|GLU4��_b�g�%Z������_)��4� 0�@���R9Z@���Mq���ͱ�~O��No��� �T�aJ���p��l:��v%�]@�@EÃw'HB
��|�%���7��bl$�Lvo�����8 ��-��}ߣX��}�2��"��{�w�P����SNX~7�X?~���P�b�[�"MĘ���lQ�R���z��~z�~�}qM�0��^�V�ɂ���l5�<��s�#8~�SAh���X[�ϛ�d�*��t�������3�5�&"%���>`���M�� ��1��i�h��/������m!A��b�\ N��Ñb[0��N��l�J�[,�Y>���g�WZ�ä0�rv�����l6���`�L�r92�6A�C��V *�䃵ޞpH<����td#�9�_0zS\:)�O)���E�j�a �� F7')W;BݐTje'l�x�s�|)�P��dF_6�J&������i��\*�3X�a��)�������)�j��2�g[��-a�� -��o��W�Ev~V�bm�Cc����ꁥ2qw�ڿ>�]"�@�Ј�7�l���wa��&�������?=C}�H�%)" �'{
��l2�� z��塝\��%X�M�f�+�:�߉���u �Bbi������,��h˲�>r��ol9	#1���`گ1S�W&��,��ɟ�gmU�S�OF�0��E�{�G)3�i�����
nֵh+X��Oqk�5l_�L�rZ�@��/�J��R�p�J(�A���	��$�i�Ba6Y�A���3��L(^f5�:Vd�Ǭ@'��N�V�ma�(������� ��	�KȒ��_srJ�2�s�ٔy)�`���,��)Y=&�J�L�#�D�weވ����GY&��~Y�-rY`��0z�oO���G���<m3�ȝ�+����gy_t<P��߭W��Z4n�T8��S�2�hWQfLw?)h��=X0X$/��!��8γ���N>"W�������6�b��~T�7��H���l>T�~C�����o�Q�#�F+0�@�6��Jw-^Mv�A�z,��-�9`>{�k����P�b��bx�Э4�9h4@�XR���&�L&��ď\��Q��^�����q�5�T��>$4G=W�jZ��Ǝ�XI�ڴ �-�ϖ^ޔ�-�?��z��R�}>"w�.��e��T����֯�ڏ#5���9WI��Ji�rD�%�O-���3-?iL.AywX�=Z����j>��{Y#V�"i�+I��.�'��[�	� g-B��#՚&@�g� �=��/ C���vb��V�'�L#�>�2�`_Ua�m��o��l?n[��?������C�$�:�#�]�,E�i�&
�A�S�m���V0�\���8�>b�U^>J���� �ۓ%H22k�`6D�ꮥ��m $7$�˛AD҄�?vd��<� ��K�_u��
 O�3"���&�D��=����.�dܣ����X�>࿌o�߷dN
����m��h���X)
 m�=��1mh��Z�xt�G����-��8�����<��Y������ ��P�'5��}s��=�e�vT��Řn�;��C_�j��vuM���L���\��e�q�K$p�c�����rR�'���x�݀�2Q���򹹠�l�p�x�̱y�||��?J0ܩKZ\C��5SO��´��ڬi�W
kÄR�&|�L�2+�U əq�>L�"|y\��K���XP�n�Pf�__�z�[���~�Y]����?��#�����CM?+c�ml)mF����%���5�]�Of,�0�e�$׼{-�abD<]��wmg��4_F[^��x�0T����0�NN�%�O2N2������Ϥ#M߯�uŀ� �n�k�L�M�lP��b\lUˣ���YT롷?�,��o��[��n�:!��_>锸<}|����g{�^>^rr������[���K
��
��J4_��$!��S��aB���qX��{�xk�  ��6�, ���C.s%˷=�MԵ\�x$y2���� P}��?�:��������,�z@�i����OI�5����r�3���7�)��Pp�qWҬq�u�qhUfU�~���r�3De�b�.�Cs��LQӹ7f}���7�Kۻ2���P��Dx\*G�A�N�6�3���e��2*	x��d�,K;�p8;�tg䤤�O�(Hs0�b�c�l�ltd[�qD���"���duO99��_��l7�K(�`���]��BH�&��CN��q�p�7�y� ����e�w��C���b�C*��C��,�~Ǆ�*U�6�g�q0i�Д6��[���[����1F� ӿp� /c���O6�(*���N�Q�MD�%���v���P[�F�gs�0	h��1�>؜�h�Q��M�M��F����E�p)	ځ.p��i�����x�
�u�eD�0`LW*���ā��Z"v�8�ov��j0�+�)���ƭ��9�2f�	wd��W�����'�cw��xҎ��C��M����el^���P�seߊd
��Ou��%�(�swv�d"��}����e̴E��q����$*zN���
��^�7�W���L�)���� �J���
���	��I��MMFJ���x*=>[�g�;�)b\�pg��r���X���cxR����iqǠQB$�qj�1r��czy\�}��o4��.4m��O�4W���Z8�A�4�4�,1�l"�{�HYA,������N�����$����$5�DVҧd��^�	�fϋ�W)�)��Z�}�l���@ 0���}�
4{���>����F@���/��n��SB;>�ܐ��%��!`�(Y�ٲN�v�N�35�yS�u(]�U��z�/ٴ�~[��j	��
i��U�31z�4֖�i�\9�e�ZZ�T�@��)Ֆc������\�%#sw�N߅%�vAR��G�6Ř�?�
S�P�V�T���(4�)q�歲]z�Y��fo�f	|��ӊ�w���˖gK���h�uR ���U�=�������w���"`c�?�ی,:�5�&ǐ�fb��a�}����s�-1N���f�����H�{Td��(�+52��z�$�$ܬ�Kю���i놶x|��K����ƌ�v�K$}���`���_�`s��U�_4]���~�T��@�ա�2lj�i�`��P �rN>�6;��M�V���GI�O���VXkyO�O)v*�9'M����a>T>��K�T8��g�a�όr�.�Y_���q~T�$i�x�̿�,�O0���c�T���Yٷ�~O��>��� %X�H��	0�w{H��Ђu�b��I��w�!��V��ZxT[`��1n�&׾Is{��ϩL��&n2	ڒ�e�\��7ڣ���heV4
�sJF��{��SA��2�~��޳��we���KvI���V�~dK���LGd��c�2ލ�7
�"�&�j���RC��"c��� �(?L�ON&���MKd���~��n���[���B��:0f�G�f�X`o�Ȭ3�ԁУ�G+�ͯ�$���3P��Hv`�|����16�	,�.�HZ�Ͷ�r1KY�-n@��-At���6�g��!�y �s�l{��ʑ�U��\Yy	��ٶ�Й�-:Q>y�dbuh;����I��
�i?	ψ�(��j�d��PC�݈��n��� ��lB�@^�y0�g��?a��r�o���˃H�)�8q���'�h�<�
 ���ol���d��&��9,&���=e1����\�w5ի��w����^����XFL}4+��8�q�Ԥ[B������j�B��Z�����k��$�	� D^ő-s��<NsN�AY������׳9��I�� D�U�Q1�l�js\�=����]�ek`�������˂u�>Мa��bk��z{n�,0h"���V�%�[X�=�[d g#ʭnfm�i��|X�٭�ks��+/%5���w�J�r�
�΋U&7J%_�s�����s]=�6�@?��y�%�˒�MQ��j�{ �iS}�%����kӸԝl��1��1���lp¥J�D���f�{j�xn�V.�b��zy����K<i�l�XfI��Q�d�U?9�G4*��Yj���윯!fg�nQz�~4�#�@$H�|��M4�S0��v��=Ǒ^�r������P�2cP��͗lJ�ٌE�(`�iy� ��\���Y�$�# �����beQ ꁄݡ�l���zS�k�i��ڗ�f���T�%%Z���,e��P��ᰬ��4����Y��~��a��K�h+� #÷^^�n�s�ܙ���9���!3B��|r�[�yj��^	��8񁞱>6�n.G�+��${��&p�f��ɩ[�C���/6�B}(��<���-r �Z�Dg^��b�s}���]����c��������lU���<O�\�%�W��'{5bIqH�.lGq{�܏I��̧�jj%�C`F�#�����x�s;�P�ρH���y����&��~'3��e��IF�HfK��]X��|�k�:�@��F�����>��T�X�i�j���/o�^�4��O-Y("!��_(��(T�*���nB�UJ� �IRIf5c�A�%KjOj
iS��{�b4)���a��NʀL�*�:N~7�Z�:�t$'@�f���X�7K�[�S����_��W<���}����nu�keл7q���y��ny!c)g��2�A\g�J&3tO2��!@�^��N�<�>���
ж�o:�[
W7��S�CU�� ̪�G��E�\��O-�'�z�(}v��|BaP9+/��;�Q�;���rԝ��c��lS�Ӷ։XrF�<�Wq��i��RK?_9��A`�UL��gZ�%��֦��)	�aTCr�����_�MG��#by"�w��B��P���Թ�,�͘�^��x@msC�A�	_0��3�7~<f�W���HK0��ݲ�<���2�s6����e�Dy�e����E��eF|Z	`�)�v�6���qJ	����|��ܥ���ȺCY���䚯�nI<�2;��	���i۔`:��ɥy��ew�D�s�cpc���n	x�h�q4f�3A�V�� ����#��CHqp_CK��%�KB��,�Q�N��I� [�GMe۰b�l�M/�n�]4ź���+�aX)�R���( ��b�����8�+�D$`� Q�\�������?#��D�@[����ʻ�)l�P���J���vq�i�B7*L��d����R�F���`�&�G��.�?@��"3���G��|C���f������lY�MJ��?�W������hP�%�؄���]�E�QҲ�1�m�X�^��e=
���v�����U�`�'�t���{�<b��p��}��P>���Y � ,������.,~r��` ��m�/��d�p�S�pgF�1j}~k�3���XU�ٟ �H ��/�T�������+g��ե}!I�A�8ʗۨ�����{����`{������G������t�п���	D������[�וS���V��MjAI��+��HhK�����r[ka�gT��2@=}��a�>��Ta�ǱL>>�x(C2&A����U��<M00��ޜ���x4����:����k���C&I6��9�ybߝ�Bt��&pY}�S���-�f�/��:����ac��U�!�]k -r@n��:D$3#A��Ռ0��Xjys���|�w��ff"��I���@J��} �y�L��ni���|�;c)�B��̽��	-��w׼�$&� ?�H�� ��Q=�k����m�ݏi��K�A��4g�&Q�����M��6����~�а��[�ٵ�l�ܠ�q*vT��	�(&���<d7,z�>Ѧ;��-�=b�͓��r�k9����ö@9��VOJΌ~�9�t�񉤟	��I�{m���z`����P��Lxlu�A�Ln5APsO����� '�(� lY��O|�u�:��Hz�IMh �k �MƄd��Y4`m�fɑ�@�|$�负ԆN�S�T���cv���i	+^E�4�����;��1�	Pl� �u+���"_ \��3ʣ��ϱ�9 �mNf1h��^�nAn����摫ہ��z}=,K�ʲ���r���dr�[�h��g5�2W�0)
?q���Ѕ��)\,3H6�Gs�ۡL�(����2�X�
������b֣ѿU�w����>ԅ�np�7c�Ok=�A��k=�v,�LT%Vs��6гG��~��!�5���#�)��ւI�?y�o5�l�*$���
���#c2H�j���`T	s�X,����I��wm��gΦ��������"Q�ͩ�s�c�`�8G�B�e[b���H�Y��X#��?c��f
����ONn�. 	����L,��*#���c0�#w�d��}�X�&��A�-)~�M��bsIn��05�e�ޱM�J�{������LҒ��<����G�T��{�t�b������Qm({�n�r�y�Ǌ�_�9��@n��i0Pkئ_�����dV� *�?&>{m�0_}4X���1{G���۟��Z�~����J�T�gGX�:-��<��ÿ:l"�cKs�aH!�g
�}��k�jŉQp6��:�.&��h$$[݄�s�/��i�I�"�bR� �^;��]�OZ�	�Q������PX��6�H�av���d
��_2X� ����+���[f��b�N���M�[�4�#_8���ٕ�Q߻�,*eQ��j	%?W���UMS����=��P	��wvn�Hb���N�k�����Li	���\~����'��Ɔ`�N�k`�`^nά@���3���*;������pO�%���m`lr՝0M'֩e�4�Gf�J��9��3��C$ �fj���
�z�}��7�`���<��P8�'���9�*SQ5+Dn}�>T+�.l�x
��]���Nƻm��7�F�@E�p�	�K�1�)�~��������{�7O�|5���cm)2g��OO�kw�בE�|��b]��=�.�P,��7��*&� ���n�J�婯eq+c�?C�ۋ	 b��c}��ܯ��y��y��dIR��I���@����d���Ԃ�5�`d�V��b��k�V��E�z�e��ּ]�x<���=����J���3-�����P6=g�����=+��41)7�17}[��C�JM�
��$��R�:
��"c_*��1�y=~'V;m�H}���L��٪PyEJ��U�K={O���a�;%�n��'9�~ �m�~�.$��J�~�|�7P�P~����2�k�
~���n�!1������Ϙe�Y�����Z� ��{�E��`\�7�/c��5�25�;͇
3�˹�+�3�fq��}�%�����I�D*"sg��3ۓ�Aφk�10�}���<��C!@ Y^��Q����M o�'�.>@���Lt�O.�!J�@;�
YN�# �1�H���^�حu���v�k=��M���n�rpу,#\N�t	93Wj[�W萵��b�b��ݗ�ɤOD09�|檼ը%6�ji�O�=����u�dɗx�M\Ҹ�����P�E4���8���Q�@<y7�/�&�OX,�w@��O�zg�S��2�A�A�``��H��¦�����11S��4'��i��X�[�\öԩ��ͥGG;\noU�
0�`�}���#��{�0t/��g��P*n���F ᭘(�!4�=���b	k�k�dzU���a�L�� O뛊bnD$����rX �=�#M�YL�bgcG�Z-�n�`���`����2��_�& o);�h�q�E �{�HN&=�_t�������_���C�˿�k,E}2k��ɨ5|�.�Cf~Ac��NA��6��p��/ ��X4�����aHL��V$�W0Ƨ ��K���U�E�σ�*چ����5��:ޘ�ҿ\��4��	�+�����>-7�A	�f��2��l����V[���I�a;��D����S�kr?]\�	*��Q)S�#�m��P_lL���t�T�RR� �M�L�%3������g@�r��4ݖ�ʾQ X��2��#�v��y=f��>�&.k! G�tD�ղ�Ȅ׋��z�L�_v�����b�c8�{@E鮟������7y��9��&�W(7�' J{���~G���#�=4�2���[������/�;
�N�Q���J��̬��OY�$7��j˘3��0贳}�`I����f��A,����KY(���t M���R,8�*.��u ȅ��/�N�({��jG��m��Ѹ�}x2S�Cb��C.�oc��Mr?%����#�dkB�eKc=�+L�9� i�JDHȣo'm5��o-c��g�
��+�J��M�8O�a.��?l��<���/��W���:�e�����<�P��lsȱ���Z) �e�C��ld����T1+F��z����ϟl7T0�U���|����1���"�1+�)țm!'�?,R�Ɣi�?HB�%E�ဵ�~h���Ϝ�٪��+��O�P��H�в�x�8e
v������c�������M�hb�-����7�x�
ժI���NT�*-��p_ni�T3�����
��s�Ǒ���Iۛ�|�~�}E\7��\��.��w @B�_�ը�����h�d�+r�h����y��߂jmd�� �ag@�G�����ׂI#����o7��P=|�{�l���==���o�ٷ0Yd��^�����ADRf��	m�;3F�Lyt�n��3�(ܐ�=|�:Q��s�*dy �V�8��M�I�-w��� ��n��k)G�����B
>Lwƈ�15�6�x/4�����c$� +���	p+X�T�%c��Tq|�Џ��a�<������G~���ڒ��M5��8�:�����ˣU��x��R���HM��Z��2���GE���cR%��mO� e��*��d6w�W+3v[7��@(�;�m��\���rGo��>{�j�l	�h��<�����[�6��w�K�ơ��X����r���]r�'��R'�3��>��GM$����Ķbc)� 1�<	f�z��b]V�dZ��Q~�����z��26Н�t�^���0ہ�c�v�5eq�u ɉ��a�(w,��*Y�6|���B/tO�n�L��� D�gV�w8�&�������K@GL������p.��ʞJ:!��a�X��#��
��*�ɏ��rla=����D�?+{����M�oh�H��	H1P,w�2ӟW�;]sX��5تO\R�9��|z�0P����������Bb�����O��T5]��0�J�vݓ��"��;���E��nޮ��5Շ�9:/�{Ӷl��p��9e�"KF�����GBO����;LC�ij�?<ˇ�oe|�Y{=.����G(�-�ـW|�����Y�4	)����G]/����ֆK�X��QO�+	e�ˍ����wD"쑦P��w���7Vz1e����A~����í�?o�l�0�E������F�6f����5��?i�F�\�+������ ��f\�')�"U�e����'��uI�"�͔��T<����/=%����'�O���m��葆�XҀ� ��@����1`6�@��l+w��m�z&��X�A�b	|:F�D��V�)Z�׮�$7�V���6����~���>9�{��5�c$�k[CVx�nf�-&Rz�%��n��Fɉ��<�s�������R�I@��*��l���[.X���8M�FX�D�n��KK?n�-h��7�1*d����I�,z"����ω��|��Ű���t vA�����,1g��/���V�9�t<~Qύ^�|9��..�<?��O�!�r2G~�P4���D���˵�O۳|`߹�X�o�}٩��z؆�����_1f�I��WS}���֢m��_]߻�ڦw���/�A�p���,���#/k-�v���g�G��bp{Y���'�tR<ify+���16���k�tJ1�f�H�<��b���}���HN��E�c�D��ܒh�jg�$����4�]�Ok�����V�]m���P{�S8l�h�� ��MCy�@��=�Uw���c�g%5R��n��K��ܽd�1��m9!ŘC�y���LSge`�r�b�)��,���)_���B�`����^#K�g�G�?�	��&�<��m8�����;�S=6ſ�b�1|����o�0z
+�0絭h>_�}�fT=Ty�Oa�?c|T��u��)=7"tg�����j�G 8|x��'}n��3g��̃��t#ԍ���L��
Y��Fyx%(=���g��<	��.���n�5C�Y���j�I�����7u-��^(���H��~m����>.99v��@��p��b���40�Azn!M� ���ߟEˁ�N����;{O��k���������R����Y*?��ٳ��b�ϟ�bG�38j31�e\.�&�su�������>���-/*��|�x����=�D���<�Q�� pАok��a�}'l�������5�.V�VPi�]��&1��	�
6=�Ć�f-���?pIR�L�vA�L�=��+�>�9���w���X	��7q++�LP���#�^�zA�L�ⱥ� IY����1"ݑA��PQ^��Ї�P����&�5'dz����8̌�%`����L�X��~��$���w�d+]�| �����dT�ǹ,m9h�K�3g�㎥<+��s��f��a�,P��ɽ���8`������L�
d䝎w�Sj�Ռ��A$�`��Ⱦ�nbTY5��_�Y���jm:�ae!:��I���(�_�ݘ��V�����`�V&^�������q��X3e��o��lJ�l�[m!�ף���>�\���
���r��M%&��'��X������3�[�:�������ἢ�Hz��T�`�yyy����n����W�\��{��
sb��|���l�P�-��a�Ԕ���"͠�k�5v������?�����/�������l�Ĥ���Q��%K4π�m�@����W�_�Ch�SP��k�6��)�v�x����qo�>�x?j6j�Bq�7X�{�S8�5�� ����4��^��c�P�mw�|�,�� -�{��FK<�B�hi�xh�2 �X����C�Y���#6���k�)���x���/��5j�Yg�:|rN�\�4%���V"J��>�g��z�i�=�`C�&��^{���F\�� h��:y���w�!��;)p�O����	�H5;hs�*(zT����R���5%��.���e��ʺ��<E��ʢ_����������������������h�!^&�*�H���Eo�&�� �WJ霅��u@��H�J	�-�>��<�u<8l�?�m�	X2vf�a˝p*(��t�V�������o�MCɢ��ϴ��g"4P�ӬOHkE�<���ұ�a1�J
-�b����`�H2�s�\��%�J6�J1��V�����b��ƌ�8�=�&7�#���NN���o>Ɂ/�(r�Gн4��G�}�ԺXl#dn ��}ϹB��,z((V�([��ٛ�B��W}|�a�!\�r�� �ǃ^�Ƚ���n��al�������	���͟���KL�����|�&s%�a7җw97�HL�nYP�=�n�s���@���0-ө���i��\
n
?�<b�<h�O�����X�(�Jf�u�rxW� �S��{*u#-=�H��A�C/���ƊP�����>$L���*�X_5�3�naJl��� �t���q� ��H���i@ ��S������[�F�Y����	3��%��=��+������1�F�����Y�d�
����ev��?�g���"
�Br�*����>kl�Zv�E
��Gism)��>���N|��[-j�TW<>#2���|TA�|� �>����(�ۗ�<�xj!jI �� av�kH�
���"�d�b���J����C�}�9\�/D���E&;�L�2a$#nss+÷zΰ���U�,w��Z��Z)Å$�N���U4
J��K\sPK06Q�n�yOuʲ�!�x��Y}#P傶�|�ɉ2�;��o�g�S_���,XB�jqt`]$T�̻H�����XL��,�,�?��N�z�����E��{��au�]�=T?�\��f���/�?�᏶��y���
7r"�?�ʚjh�N�F���Պ\&�ڊ�sb�LØ�WLP��͖�[��b�se�������)a��`�Tg��A����r���"��:�]g������L���Y�����g�ڋ�����e&;5H�x���P��ˠx��#Y��?�����&�c�7��9��ho�C�2�평�N�jԏS9�v�����y�P��Z*���Vc�b�(a�9K���"$
�t$s-�:��Em���XQ�G�i�-�ǝ[��;�a���#.sB%b�i�i=�&@3�Ҝ�e�~Uf���Gc���J=�j��,���_X�Lu:���ҷ��
��ɀ
��~��H�U��*�Y%�����G�4)�Ȅ�����"a��O �i�e����;?1����.�u@�k��ו�рX�#���+Y��h�j-�(��������Q �/�9ُ0l�V�������B��e�ڹI�mMD���Zk��Vb�NC(�F�Ő)a��5Lv]�#S�Q��v���Vr_���������K[�g�2��ҷ��[]|Ǆ!^z\_��%S��G����E���EM���6�+ە�N�0)N/v�'�1Iu<�2��W�E��)�X����f�>=d���~�� �2�����Y�������fj�ځD�KF��H���.q���H�nL
*����Z���K��N����Fو)���60^�3�/0����{������"j[H�&
��:t�β�Xĵ{^S�F�����ܛ��9���z묿�U`��A`ŋ���^I&@׌K�x��p�� ��	M�c��	���JX-<£)�P�(�)��>%�UL?��{s��J:����'J�@?/�U;����a�Bs�2��f��:��^��+�E��T5��ӧO2�7��7t�j��p�ڟ�\`��h�א-~��u|��������RI�O5�Lw�ٛ��-���EV�w�
���=��Kǻ0Tf�8�����l�4�a��gڞ~�$����Y
����';;�0m��g'���*�kW�q�O��KT��Ύ���T���PsSB6���_��Cks��~SS��}A�%�p!�ـ�������Y���G��c�䯗��#.�\ѻYP�v� E�BPY<��7����+a_�Z�������� r�C�Q/��TTƜ��n�Wg�B�&�`s��P�W�J��<_����zTf���6P���vj]�Ӓl���J?�~���|��,&�4(_T��ȱ�(����L�O'��*ok_��K����-��*�i̇0�����>����m };E�?rR웯�������$�4��t7�"�����Cү��$8/fAw&��*��g�==��a\�����qH)|<,�4�&�%5r+Qwp�,�5�Vtbm�I������,�\I��Ԣ �$�n0�e@+͚����.߇z��0Ϭ����ϻa��u��F#H%ްs����w�F�߭T~����B�X^amK�i�@60q�nZ���2�9�- �m��Nm��*���	�ԊѾ��o�����}�HW�l��'���f�`�ʻw��M�0�y2 ɍ6ިYa�H`�{�	�9ج�����;5��濥.%M�¹��M��I�[
*̟�6����M��=�����o�%Y��K����}_��y�,�|�Ym� ��1(�L�'�nsX �	,1�\�"�u�q�O&�{��e.S�K_�V�[�?�w�rr5�c���Ԙ��~˷�E��R��5>�x8�z��r�g=c��3��|�c�drHK����z/L��2�q�rG4O��pG�Iz�m��W��٘63N��N����ⴉ�� �������� �Nڋ�&�{|�,�Dݿ�:����YiDn#
�b>T]Ǐ-_�����-}�>�X�7ط(�ob�wJ����e�\S��(S�i㲒�)�"o�9N��ǻ��F]��h�F��/R�� &���䠬V�L���3���~�3����ڣ�vg�zS�F�d�,y�=�	����b�t�#�����_����L���$���V�PJY�(08�X�_\
D,��:��ϺI�����?#dL`�I�U����������X� yv^f�������l�U���R��x�?)�Ɂ�d&��ZN�4�;��9�i���vD�g��M҅�f�J8�޴���yO�7ah��{,�j|�!�u����kQ1��1����d��mS��j�a!�3��Te�����s�%Q� �f�L2V���L1��s_9��S��xC�S�|���c�����]L~;H�Wy͠�C��|0K\g%gߩ$��$��}�� 	�˯��mN�,��)��r�"�#*��΅0��o�&��GlY����M��w�d�׎oQ���]�o{�L��kW�X$�w��O�n��E�ۈ5-B@\o ���.?gvg`z�P���^W�^E��$� �	D���tz|Q����C��1J�%�{��)��5ƈ��a��	h��nsX�T������zNB�T���tA� ��������[�7��̉����g���`�}/ ��ߛ�#��s��"�l�.��	hM`�� �_��A�,v�E+���PK��% ����.�&Y��N��|6+�/�1��òM�/3(b��8cP�	���}d��P�9p�G�����e~��-�n��",�A��۰���A9%aX�ܘ�� �~'Zv����<��=�K'Zkg��=P����)��215�`��x�j9��n��>?[T�� H
,=�m�.]X��.�[�6�epBV& ms��_]o��6���;(
2�J�:�)�Y|�n��wZά4'��3uޘ��e�{w�`Zg���\�%}_���<�N�|YJK����<zF� 4r��3��ݝ����A]�=ǺG�W��������w��廉'o0@����'Gyz�,S��'��F(X2D�ݶ�C]�-��)[߼�O����� ���O�=�x�-P�}���� �](3MS��Iӷ�$�fj�+���ٖ�-Lt�.��TW���Tm`�< (�7��%m�aY*�(��M��v��٨f�Ζ©�|Q�_�dtP��-�U{�N;o"S�&R,`HP ��ūz��P���b�(9�d/���k��14o*��Y�K��1R���5=�D%'M�49�'Ӊ��rjKN��$R�7�h� 1��t~ �V�Н�Zm8ϰO��c&(�N��o�)�`�gj/�?kz�|'���؂>TG��c�B̎T4�?�R*q��v�>��P�n�Q�=��Q�&�Z>��4�D��i`���r�R�^h�t4�2�,���d��/�D�]��%����o�S�ޏ�����S� ���������ݳJYr�[2��]��1֔�hǻ8胈$�=��L�@���鍲K���Z.�k�|���ȷ�@Ւ0E�{�,䙖l����k� ;�2w}E��-^?����)
0���WK4�5|��,m�r{�9f�2<m�냶��Wxz�4���U��daV���I���s�[������y� ��v�
���C~��g���_n�_3s��njh�[jG�,�J+9&�E;��0m$��]��d�&y�j2�R;��!g0,6m������.�ůͽ�z)@�wh����m���Z;5<�x�6�-��k�����v���d�N�������~�w�m�^���)��,{�1{a���-H
Z6��պ|L�B���>Y�J�0�g�bܽ]���A��9�"9���L-�~/�lsV��N"C���xBj��#<gT���"~bɀ�
�9�U�8��?P�d(6�!�2 ��su+?����o	l�M*3���m��
\�\ƒ��^�.n�	mf_g%BbdR�(�x2�����e��Q+��ӯ��*��~>�|����]߯ϵD�1a$)��;
��e�H^����R��s
��-:�e��Fd"��I~�Z�ҏ�^�z����x�O�~!A?��5�f��|;�0�����i���ѥ6ak� "L����A���M ��&S60������ngL"XH]�-A:['�J�4�E�ҷ��2����z"3-����-G�o�nN�?bc�މ���6dR���9���ۜ�n7�X�r52�m;hݤ�����2����i�r�9{?�(��$�Q_o�P�en"�<i_��,d����A��K��})�-`_�c<&�?��O�lþ��I.�ob��u������9���6������ �i�Q�����T��)�Οl1�$vg�ήS��l{��x����@уX�	���2�{��э�J.;��n�i]�:3�kU�מ�$�	?T�@��!��{�UE#���B��7j0���:�~==�ܦS3�(<�� =��o�GQ	���i�6�Q�Oi���|G٩Y+�>IMOU(=��w7$in�Ʀ���5�&��yޞ"#=v�[�:Aig��e�-�v�G~�0c�����-��=�_��OrV\<u��8��k \/���3�������Tn�]�۞�X�rV�q��͖��5 �T"�+,�K��k4.'�-����@�o��el=�����WVɆ-���ҒӼ�b�ǆM�1�n����ۜ�x�q ��mo���&�[l0�l�-�W��Ү���Á��v�߃��:E���б얉X���ڴ�r���ۄ:�C�V�Zl	r�,�P����P�q:N��O�jq���dy��y"��`.2K# �9�xH_��E�!�G��:o�{"%[2��LK#�rumn�MJ̶��^t�V%����R]<�C}�d�KO��p!��#�b�u$c�F��ʟ-X�����]>	�}�-@�.R�M_#��
�K���)�v���P�)��K�R
 ��ԨM�i'���Y��k����Ï?�>0f6���N'�eN�V��^��ַ�>7��Lz�lR����b��l/�r3q�
�tp�391�P�X���_�7]�Cgj�!<��6�;\����6o�6���)і	��H���wAMfv=r��xiZl���Ep��a��-m��8�y�ة�Mm��]�ιJl2��`A���sX/���l�u��P��I��")3�#��&}���F��c>?��C�"�p�e��Ω+�� }�}����m|��֜��1b��]c�����t�������Lh&yI�/E�촱���$�2�d��jO�1*ы4�%#�c솀�G�����q�x���
|<.ub#7^cߐs3^�}�"��r  ��mވ�����L�덥�fd�?��lG�`8Oi����C�|@���[�g��1N�����"KP����#ho#�Kg�{C�U�wO�6|�zs�V�P>ͬk��". a�{�����}���q�,^c�U'����(��ۺO����b�W��V�F��@�>h���K0qc/��Զw������hZ�I˗�%+ꦼ"��,Y�T]��Ii��z�O�_��0�5�H��H�/=�7�kYO ڶѿ�W*�:�"�>a֧"⢂�r�� �
Y�����yA�v����ˬ_�ge�C����q����W��߾v`��)v�	���3��>�`�n�������Ϋ����g
�Y�b4�p҉�����e������!����=���k2��~o�&:]�hhO΢u��{21����Z��AZ�P��'3�} 7�����ox'��Z���_���ɖ�5׉�ushm�훼��r�2���ɮ������ ���O[S�r�N������HR���s��۶ |8b�����!0d�����=��r��6B�ox*���BP��3���-���$Euqߜ�H&Y�ET|�S_/?�.�sn�����=?��E�h��]����\�R�ۅIR�:��,$�p�ڲ:=�/�_r���t~���Br֨g7�ⅽ�r��Z���2)4g���1�{�K��ߐ[�60T��܈����M�v��S0��?�AxfWcZ���`�f3�b�]ˣ�tD�5�<��V��%ƚ~2�b�I4���Ckx0��&�v��D{i[�!+�^�v��5�
P� ��걟-�qa5D���5�����P�#�LUɘ_(�ُ�c$�t�b�&��6��,&��R�x�{��J~�|PJpo|����ܶ����q���9<&$\Z�6�+���������W���#�]"�6��2LOv$�?}������=&&��gR �vODHM?��7*�%.�g3�u��3�}��!w��=�/1C���F~m���EJD\$�4�w�Y�;A&㙕�3��������`�W2cq�$ޣ6�O �k�xO�"�xR	�o�h�э<8-����̔�hSh���.zJpԨ������zZ�6�}��V³<a�k<,��]� n�}��de����� %�	>�� �+�	]�W��[]�L{�$+�.;,�+kD�f���5TNj���w��o�`P�E��[�8z~~��u2�Q�c u��(�N����!��¨���Ev��0�K9�}�P�j�`�M��R�~�Q y���L���5����_��gf{��|��n�z��q������RJG$�T�W��@���~?������pU����tL]u�	-��Dyz��{��\-�,_�|P�+	$�1�UϜ�[�_��/qyA;9xG�V���4���W;&q ;l�16=o����4��b��Zb�'Fm+�����e�~�v���s�_�j)8���S&{֍M��j~f)Lf�UXIާ�,ZȻ.�e��Ɵbyj�v�Յ!���<���n���Y~���w*��X��|�z0��Ӊ�\s����?ޮ?|@��(z?�'���|G����'�Zjݯ�E��GF;p�j�x�va��k���et���A��p�q����}���f텕O�{�[^vg@�%�Ĺ�������~�*�>~4�v�^�}N`/^X������pSD�>��|f�?�S����	��{�����M�cf�!3/�/7`�l�g?ŒDw��i�8�n�����r~���ϯQ�٥37]����X.9+�j(/���*ps����A�5"�r��Ty�$)���m���)��Y!(6΍��e��ݴ�k2�d��#�>:�P��=F,Z�k3ޗ�FFz|�U���Y��AZŰԫyX
��ZP���~�����Ab�)���w�����7GY����su0������	���o�e:����ӧF�,�# ��dn�|}}- ���MaX��f�0����"$�.eM����"(K���Lz���N���V�+����q���>�"D.av�8��a����f���O�b�33oS�[�x>M��r�����(�_Uu�2۠%wX�H0��xy9ne�怷�_d��\ ������1�j%�w����v�E-W�7o����ٶ4�>���.;�~P��������/�����)���7 K(]$I)e9����l�����J�$��b��)�4f�W�e�[(���/n���Ė-�^`��ճ�[~uW8i���@]_VY�v<P������M�iyhC��Y˦)�j�
�'ty]%�)�a�Aq�����\kv� >���=Y+]H���zl0G�R�6q��*c0G�>/�gω�.3�'H���|?XZ��! ���䰜4ۍL�kG�X
-�7����?�=���+���f���؞I1<�!�	�Hs�w�-�ݞ=��H�($��*�,�ʘ�͎r�[c &��{\�\�	%lq'@�G�'��M� X�R�빏?� �˟����[����2��V<_���i �d�d�Pg0m�l��O��3���e��߷�*9� .��n���ܑ �D�E!e���p�xĽܟ��^oZ"t<4۔�6sxG�MF|=l�@�?��Ҡ��'�����QW[������A�N0,���Y��ߡd����a�ϙZ� �-�}�?�|Ѕ��E��9�U`�.�|�V7թ]#��|�b����L~��G`�kL���.(�(f2�

'� ӋL��L-d��%}�sj�su���{� ['���ʜ�]@�cf��-�|: ���7M�	�fj��:/�A���b2�wm\��m��Y���]�}��2|����\���"0?��,��.j�z�{���N������^�q��Ly�왏����u`��o���ӧO��.������ARP_˨�o}�g���R���>�x�]OG	����;ף��]$��q��k��P�;ԇ�/����!��L��Mɡ8��N���!R&�?�|�2���ό������ߙ��F렀�"�ھ�K�Oa����zY�A)oY.�Қ�kk�Nq�`I&�?��r��՟ح��O�)�<|��j>+�&���,���U��%&&����%u]��[ ]$J�m5dcXa��o����"�@M�D���@*'V.M
aBJ�<Uw��H�!F�\�x�+E]0��C �͑�.r���<� 0^�j)�2���+�>�eda
t���잫��R���Q6m�	P[�T���Rx]�a���nz�Z��� ���zcC�&@=�n/��8�l�e����(@U����>|�魁���?f�bU�ޓ��&b���O�ی1oS�����.-�����	�b�D[�:m
��m��M��7�`O�.mK�<�J�a �����`'�F�>�=�����d��5�"\
}
�>�&�~ʃދ	DǣRu$�4�/��5?��G(����6MX�m�v4[4�Ҭ+��:.2L�=b�`e���Ƣ.����pLn�WP$����m|�؂��������������B��ax�3E��)W��,�,:�x�L��
���_��oa��\�; �іקk�M ,�����_q<v��/�r����
e�G����i2_����`>�£��㊀_͡X��ͽ�N]>�we�4
��h��ta�e��i8��C���	�X@>���	�m$@^CȲ���� �W������ �F2�Ƭ�f��l3C��l�Y�/�E�B̞��q$�Pn��z��i�N3�)Gcfj� �k�=+��~����ܽg��F�-\� 9A��׻���x���zoڵ-+It��p��Ar<���h8$4:�>��e~.s��yPY`�����d�������(돺��ct����n���q�_]��Lm�SZ](�W$�#�K�L���޷=�O>�CZ<�7�|����#�D7Z^�,�3�B�W �����`�� ��gÌ�kh�m	���q<]�)a����X�F>���p8��o0�m� �1���X�y���G٬<���&�0ܚh��$��������H+fg 1Y�p�Q�=�����l����ͪVpm����	���sr�D���DT a� ������
Pm �XЙ���x�{��@�ʰHC7x�ͩ��-��<���y�vJ����x�s�ٍ?r_���<N�]��-�G�Wtc�l#�,W��q�{
��{,/61��m�A�D���/�� id�ϛ����jVi�N��> �@t�oҔg�����8)��(���1�+���zg�
5MÁ@�I�77$������~��ɌR8`��0I��S�͘`��N�b\���&���kw���$םf�D1�7��3ʜۤT ��PQ�8��N0�e��`W!�/ �*�%5�9�c�bRc���֮V`3�4����-`�G���Q�%3-V�稳�үݒ5�~���ɋ�Z�����p0ө�T��%���!p�a��@���9iÕHK_�k7��X;�槊�H-�槚���o�/�`����X��M����J�6��  �E�-l�
�
Ⱥ�H|R��9�-u�����l����ø��P��k7;�K�o�O�f�$ui[|�~"ڎ��h�vH�ҀQI�nqI��k˜	_	Q�c��$�@�'�aă�K<�1W[Pj�*\mT����"l��ȝ�Ӝ�3����6ǚ<�[{G�k4[�*(��B�7�C��4��"q��%��0� k>�<��h��q=�?����c�at��f�N�IeQ(��Ĳu�'V��-�1�=׍�{T,��_�(B·'+��SU��sAp{X�]fC ��J��`���8n$��a �k�����Rv5�6�C���A����>g0�5���;a�07F�$V�Z}ײ�:��CuT
��T�_Ir���9Q�,g���&�$�c]I=XO5� ���J��O�CŢw�O��OU�zA��,����9�m�gg��.��ґ7�K�|��'qƿɞ�[�.�����t��@O���Zw��o1��,�a_j�2_qs����L� $aj���{r����0���.m��x�k�z)�q\�4 Xy���n�:D���Е���;��Wu1��
z2uR
F�qǳ��#��"��]��c����� �F�I)xF�֜�KiPYg]��/XI:�I`@]2g� ��Z���ޖ����+��z��zLm�o��5qP��+�滑=C^[!!���`骔�w���PXH����:V��;��qV ՟d��X��늡��J �_�"��+�f�8AA�f`�j�%�Wv��d$�Rl�B�v�٣Ǣ��;��"?�@WZ������*�@Kh���������S��y;�.���&����0%*��:��>�~�)�zѵ� �z?�'���z�؃����)�IZV�C��i��ֹ��<G�C�⤌���7>?٠�8zQ�i����)�k�xt�A�Y?�ǌ��?V��"�/zs�������T7MH�ϴ>PӼPE'�@��9Wp�<�b�C��理�y�<��$��}��5�$�ZǓ�P��Hҡ�+*�NV�g=1�DEˮ��)���a�ѩܻ�j6w�FC�ʍ�H�=�����Ħ��i���Y��I�4}���C�G�дv_KX��t���M�H�\)�	؉�)�#ё�,����zI�Y�V阘�F��EC׆тfb�(X�l��/sc��zCaz]֣�>�`t�H/g9W�;!:�%�Z5�Y��X������ꂲ�`i2��_�R<24fU$zoV��p8Ж�����'���֭o6�\�+MT� w����8��ã���XEu�F�E��R;ߠC�w��3Q *P�t�u>�e�x�s11T;0�[�Թ�㑠~X�Ծi:�C�v�=���O9).L�3��������A�K��]�o���&��>&P #����>�t���ضu)+Q/S���1��Q�Xr+�]�2�j̍��Z�b�?n^z�"��h��D���-D���3%R�aqw��FH�]� U>���z���0�K�)�	H�>�?�{�.8?9#���=�����R��5[څ���$�6�܋��!�y��o���!x�j��9��|H�-�,RB��v~d��~�[X�#136w"p|J(�ٸ@$PK
��~c�E�Z�M���x>�2�~>ᚥ��5㋶�E������u��rDK#� �mǙA����X��=��u-^a��bQ����VNa(�/Ʃ���"�݌S-� �b��L�?5'�>�uuC����/����%�lt��9;���?�z�d�	U0=X�+&Ʃ�����?��d���]�] I���/�k�3a�fK��l!!:�;�i�?�ĸ{�>��Bd֏"�/���u�J0Sb����"=Ug�
��z �Js5R�YUOj�9ct*Bvc
����Ƴ�i�۵{�х4@���Pq��h������ZҬ`E����W��U.y+�U�1� &�?�Iن�Ap6V�5Gvv|G$��X�h���U#ł�#�$K(�����U(N<����Y�Y�:����A�$�SjQ`���qo��0b�*�Mޯ�Әd��D��R�O{�?r<����O��}�C�R�	�� `W��u!���s{�w�����ҹ>�D�33��h�f�jb��=��'�+�C�s���%���	b	?"��c�ú}N)��"�E^���G�ᶂ�ԓ���IQ @�� �_D}�n���y�J+��d'{¢��k���hѕ��{��b\٘�d 
k?Q0�<�zPΞ������d�Z��%g0��@�i�Du�B���e�%"V�p`�=����6R1nR6�$&��B~���iu8�����N�cC��s��h��9M��g��{�ܦ�����H���4�£?���}�� �I�x��Q�� ����'%5ା��	�hq��be�����"�~���X���Y֍J�b����rm+��EL�P����Ը��C1)a��Ϻ�'R5A! �&/XI���EX���E�p#2�X`,Ib\bɞ�luOe-����i!:��t�K>#B�s�Ƈ�˳%�R])��b��k����0¯�Ũ��+��p���T��4����U��{�����u1����w���W�䱾���V�SW-�����y!K+�����g�	"0��L��'>�C� �T�@�%�{2	�5��1/�r�Dp��K���� �t�>���h��!\����ښJ=�>B�J&� �U=�de�Ln������,�NZ��%6WA}\s��	��C��U�R�7i�����i����ˇ�Ws)h�^�|��秤�}��s*�fV@���ռfp�����B$q�~2�1gρi>7��i����`�>�	��f/� !�5���d��i�+j��x�BlK,!���~�Im��ζf.�|o�
;"��_%-7}�8;��U.L!([ �T'�����&�����8dMW�b�U����8�R���<mp	h�Y�����!��,i��v����kx9�$��OnM��1(>2�{�����J�u��2��S��p���9WE�:�`��|<c~m�Ε�L�=���uS{��[�����W��睼��yG��΀���������'�F��N�4�eLpוs�§���v����䀊��u]Q����C�u:��.�X��,.>�H�K�Ɏ���k�|d�}�.�(���xY'��?s��s/X���=�&n=vF�Yl���`���!~?w\����@/��F6(0�������%bi�8��}�����p�EgK_`d��w6M�����T6���Ikn�G�')����ף�n	�����i;��&�zr����F���U�-p�S��'��� K�GY�Q�R�^�8y>�^}?w�@\>���� A��o��@�<�����Tj@��ɮ��ȯ~_��1�S�<+��KF�0̈�`���
���ݡ�������i��=.V��#�Ùa�uTCĊ�e`l�Y�X��a��9�Ԧ�2�˓�A5OȒ��	�-_3��n�؊��^QT9��z!e��Y_�[�X%�=bsЗ�(\�F�P�����_^g	�}x>��Xm�]��@)�=I4��y�5�Z ���:��f�j�hh�{g ʕ<��Ͽa	�����-���P�S�2t҅~:sLu����÷�&o|�m�ŹV���6��j*]�B�>c1@��v#��%��!�̇A��~��$��q�P�g�Z�I/7�$�oov.���g�Y�Wi�|������n�W+Q��#L�`���"4Ry�D}�#%��=��t�x�>��2Eǆ*
DBP�8����6r�,QE��g93�&kvĞ}��:�,�����QA�ޑ͘�Ԛ���B��ԧi/H��S�i���ς�mXH�c�/E!)�!���b�:�����B�Z����i)�4я�6�DL��i�\)uJ������
T�{� � ���2I#�XM�����x��� �Uu�2&�aT�5��Nl�4`eQ�'�*�N����"���NI ���ꬉ��ᥞ���ک!~���-gT��
�KY��. �ޑ��G�9~P��p�j&.���k�S@(9䷴ W�����
B�'9F����d����J�*��?l �`��'9��x�͐�,���V�����u}��[��!5߭䈾g�x��g�+6���)�ˆ�)�G�{X�EG��k@��O�j8�>[��z��n�E2em[�<0耑�'�څ��X�'�������4e;�	��XtJ�v���}S���u\W�'�V&b�:��L�=[�,)� �gq��/KU����H�%� ��>�%���B��+e�������tk��}����|D�A߆8s~S�2�;@(+�]�/J���DQW5wm��rw'w5M�[��:�=���U���
�hub|�%X(��`���X���8\X�v��R�t��Z%��N�g-�3��i�A�}?A�<�$�Q �)9"ɧn���h�h�^�0ɸ�F��ū�$��g ���7OO|bٙ���D���Lі�B�Z�ɛ���,��W���ՊřGٔg��R�$n9E��#�.(��˺I,��yn
�z�m�g(eN�k�4|~�c��gu�2�&�;�[�oXP9�R,�}� nB$��Y�oO�Uҕ�Euf�W�nJ��üYte���B�M�:oO�A6'�K��k��=0$<�<�*�0�ƛ������J
�-�9�����ՐB��A
�I��)l��.DPlH5��\��6D;<�R�v�?t����5�<��h���.
�|���������Ȕ?}@��XCh��E2iO
�9SO>�t��8��6E�̡&����Z�]c�9�T��0 8��Q�Ĵ$�9Y��7��vf 
 y>DdG�t�#��3��"kӲ�?��0���R,֤x�k �7��0���3۬�P��h��JHzQV�I ��p�g�2S���1�O�i5�OI-��Pd�j#���.�T;e�RW�x�lM1���:s�bB��6�xjY��sd�b}Lih��� 
�hPa5�b���-u��:	 j m��?'�&���	�pԬ��y��rT�|D�="�)���Xڠq���8��kU��~�������]���\*����N�\╕��$�
�C��c]c�E�j�w��3�߶ ��關u�Ǧ��.����b�d����m��`C���|��Z!I6�/��ވ�lՄ�`T�V�d�*�����O��2��&�4apq�����{h���H�W(>1nS� _Y��	�?H?�\�V��܄������Ϥ����X���tgo[d�y	h�S@��nc���9��R��n˕,SXuP��Ml�'O��3�O����,�V�E+ �x��^�xIϞ=�g�'1��n�}�Jz鰹��:ҧ:Ч��{6�6!�X6������:��s&�zUu.������Z��p��ݤZ0���.�sD
#�7�/媞��eT^�=�3�����ҝ������ș٩����'��}�;݊��p���kB!3�-H�*f�\x��E���H�b�Zwj�{XY֣�t�iQ#uZ�.H5@3\�lx��d���g�{�_���a���b���(0'j��M�����-^[�'���AI-��j�(�j�H���bN�q8�%kް1OLY��bg�ϑ�i����"%�9\DR��p��"'�P�7@�|Vm����W��A)I���V�|������*60U5����W��j0�2y�d���u��2VشJ���cŃ����/#��6���nQ͢�@��\ֺ����C]c|�MŲ�|$�,V6 (�}8�'�8b�)�2�{d_�:��܄8y+q̓�~�@�u��q�<iv�L:�y]�C��.}TLWfI!����=�ٳ!��%[{�ۖ�7�� �.l���E���A�G�&`����.p��Dy,L�#���k�׻�N�j�n�4ۅ��\��Xf�mtk�z��d�>���5�t��B�6�m�%]vK:I��#_O1'�b���
Qܲ<��\�0���B݂��dL����V����I�;���߃�))��1��G2.�^�&�й�p^
�&���
��n�Y�R���]�!�M���_c����5�'֡��"KSY\E;ec���]ۆ��-��F%�XT�ŇE7�J��'� z���3�L�Ѓ����4I�pd0]��ho����%[�$	��3�EȮ��#�M�"c�3S��$c(�i;6{��,�����`Z�I�.=���نl�L�g�*
����TUY�����$R����K���TQ��LQ�"�&n�ʘ9��h���������<�)��������Tf��C<���G��DY�#m���@��\�ҭ�qZ�U���F1�E{Lݬ֨��2�M�<�:k����� �w��3��$�fn�]]�b��V�p�<5Xm�l�5�'�6�	Q�0��:@aP�OYLlb��
ȁ�&@��BXJ��:�2���w
���K}õ�O"������~��=��R׸O�](����V�Qt�ƨ����=`	�N�p1O>���l5� �˝[��I}����	���d�H���`0F}t7:��댈ն�9k2u����j�����4u0��Q��G��ȯ@�F28ro���ˬ�*������]HL,ʓ͢n5�PҚ]�p2�1� ���Y��@3�J� ���#:P�	��/{ɻ���Ztp&$G\;�\T��j���s��,��f�5���/�����
��4)|Mx������O�C5�oB�b��wZ��_&׀��[&[-�ң��X�^� &����,���$b���zFta���u ��Pu@�=e�����|�xAo��:?f0��3t�E�����K�:g���Xl� ��YDg����)L���^�Hs��-�ˌa.:�H��z8��Vl20��j�j�,�qvp%?ޔb�j5�sϭL�Gu�i���6[$S>J)���KaH�}~uT0bf~�����bLB͔tq�� )��6S�z9��(�U�n��ʂF()�@r��ڮ���З $n	�)�vA�����l?2k���;�:��liʳY�����A�綳�c�TH|��1CTv�J��HHt��	E��>�>��ɻ��gN�,�rˎ��(և����iG�2����y���Dq��ҧ���b��?2��\Z�\�OU��:�R�i��j�n�Ӽ�L&�ju3����X��$u�>�`e��!���[S��;6,�c�B�:N���nS-0�t�L��3� ��d�~ϋ�5K\B%0zP�نd�# @�I��E�9S�4곗-�ʙ\�4�Ҩ��Q�( ���`)����A�
���,Ku�&r.��Ȃ��  �vS�X�|����z�5�=��A�E����:��\΋�_#�]໗�@֝����)n��%j�;�(�X�|��`�sM:�kq�'s��p��ź�e�eFԷ�j�1oTg�O���V5�>���	!TT
�2�'C/��˻֥�~|z�0??��1��5��A�������Jiz���[� ��wZ�n��1Ƃ6��"�Z�u<nnvt�ۺ���y{�}��="O��������J��h&$����h�ju"W��J�0����ʶ�OK�16D,��#�R�c[zh�L;ϕ-ϕ���@�����!�+�/���O6*�N�Dh0a��c�Xך)F@@�$c����R���'�rMXUmЛz�" �\��<� �m�b�4	`���{;�j�}��͟g����+D���_����E�������a���AL�E��z�ֺT~v��5Z2�T�#ܹ!;.`N#��L���|��k�|��a�ј�sc傭�P����:3���� R<�,�,��uH���Z9�a� u��Z��o�F^3q4���GE�I@��>����H�E�&D%!�td|¹���3-#b����c����7 <��p`oD����Xd����g����>Gˀ��I>��K����nS^���!?c�;�ͬ嶇hu�̶ �_�������7�y~OϞ?���s��̆:�73�G�Ry�Q�C~����	����v!�7�zӕ��a�Sr��`
��5�'w���P<�-
.���}�-��M�	S���% `K%����Ui�&���@�LU���`�5�{5��~�^�C�P`d�"}��	�Q��F/�=\����,��X-�US������Q�;䡸����e��.��`l~����V{�bඁ�FS�F5�)�7�7��u�R$ON������\��Hn�Ɵ.�;��I���؞�*͋��u��U@�{��Y��r��PE�g@��O�?��g�R7+IrT#,�����[�[��E� ��:���N�*�`�q<~�`��?�E�/���2�p��Ct�Yep"����PY&���k�X�g��@Tc�����3a��ذ�o���4~��0Z]l��_�t�� ͪ�h�$��Y���dB�KX�����	�ʋ�q�OϓE���Y0]o��snl'�_v���;")��d*��o���+:�!ΛP���U���mߨ^ja��������	]�����~Ɂ}5Yݰ+l���~�B/���u�a��J��~p�KL�0�@���� �X�ӹ��@����`�E�65���IJjj_m4�]�ޛi+��ס�`����nׇTy�H��Tc��˳r�_fG<n�'��ғә6A�i2^���s{�G�@�)�������?�����_�Ub9<��x���^g�	�3�G��Z��y���;�9�0��2�oL���t�s`몏�Z�qp�ٹ��7����ryy�	F�Y*D`��W��nF�y�M$�jނ�lu����k0��9\{L�?{F?<!N�3H� ��(2�YD�	�oŀbu+:V��y��D��7����y��F~�G54��'� �7�n.�d�e�g�YU��c��471t��u��`qxw������}�糓���2ag^�6�2��\���f{�Ev2]�9���~�z�)��[��
3ݙsx���Le�Gug�m�wwN
��Vwi#3c�:?�n"��9K<No߾�òq������b-��ۚ�¯�ڝ����7:���f�-� TW��|�׉lVI�~���J���S��0\���8�F)�\�)3����t��gB����rQR�T���?M�E�d����9d\�A���͎��z�90B !�=y�e1�u_7l����
�b{NR�; �@MQP(���N�Ɩ��7�5W���S,|R�� �E���ea2���je ��$��f4$cj,�N�ɢ�\�nv<�XT��{r{�V˞�!`J<)��C��yب�"����~E���&h���Ƭ� B-e� {�ۘW�����W@�W���'�M!:��;��[ `ll��!5���ʖE�17W%�Q�K?I�R��L� ��Qu��@vA\���~?�}Om��醙$y1��� ��N��	Rq�u�eǣ��S�-e]1�;ټV"`�)�r8*L@]�b�<����\��w�x@�<t�6@�pg��h�cs�6��<tQ@�|�߆J�]C��''�SL$��j��9��u���a�X%�̓18�2�ԇO�#^���y�}4��Uˬ$�(
�Ӭ��ܕ���ީ�<��4���ivI�q���,/4u�Zؕ��V~w;_�Q�
�,�o��a�wd�64DH�D�\�Z9��r��ˢ����]��2��6\W��g.���Dt��[%��I��m�♹�������.�D�M]�dc���i`
b�7eK7�D=T��
�Z�V��f�D ��g�J~���Ƭ	���"�*g��np�|8�k�K����e�dâJ��v���1��Qڏԁ��A�nry������zX��F+ٸ��l@&���m�d�E�l�Yja��Jgq��h8�d	괱���?�x*|�(p�G��FbRc�$�-��G���Y)���uS�n�w@9�2�o���+�����+gX��wLt$cJ>����.��6�{a`�vL]rDVw�8#��0�2�e@BVl11�r�R,�h�E�N�˅^T'�2D�"_�T�W�SQ�U��E51{4
����Z_�f���c�X.Ѯm��{�χX<e���� ��9/;�֘���.l�ls.������A(�򨮏���iލ�*�Wѹ�.�5O�VUtc"��0�am�u|nӘP�nr��^LJv<�K/�6jȔkU2�{U�ٌ!�,�F��QZ���T}�ǧ�u������K�٠24R&U����'䀥HR3��7�ڝ߰gJvm;�zA.V�gO��M�~Կpv)�8Ku��X�9�GϏ"6ts���J-L�"qG,P��]��t����78��b�E��l㉊�\fTuv�w����&$�@(^M��ٜؗ\y�n��q��z��?�T��g�"���j�gb7�ɼ��	�bfU4ۖ�O����!n�n���V�c� ��!/�"�
IgfH;I�dpٰBs��ތUBs|8X�z-����)*u�O�~0jw�*����4��3�2���tR�A��ƨ1�Q7�$�;�aсۤŬ[�RY0҆��}͈gƺK����x����،|����i̔uF9��,<C~�
Nlc�/H��r	;z<��vJ1	;~��ǿ���ْ-�9sR��g�|��+P�r�� ���z�4ՠL���4^[�SUْ����h&����aʟ��`Y�
��kYj:=I-�v0,1 YD��8;;���N�=�2��֨�:U��k	�2��9J)%��y� �gS�9�!����g_Y�gHL��&-���}YM�@��R23���}Q������[�y�<��-�:�c�{�>�ޚ=s����[s�Ƴ��?�ט!#�U�^����m��s ��k�@^�����N6r1����v�Ͷ�Ͷ�cSiU#�	�'�z��2:`��6�h�|���x��N�\��2�|���1�A��D���۝֡�92aQ�����lq��Lo�����¦�%\��!i��m����6��#M\gUX�p)��f5}\�|Ý<�Ϳ�M���x���%���sS���ԧ(��P&��Ȳ�$v5�P�@���9�7���-�qf�k�kULܰT'FL�q�hE$z����-	ΤI�(�Y�;�F��s�nsD7�"��A(mRkd��Ki��
������sHR���IJ��c&B���3������k�5l���@�i�R=D�������� EВ������E~a���
�r@��t����4�؜D�f�����؍���/�&.Tᇉ� T��?Q�,vu�C���Z,|�~�i�������hѩ��л�_u�����P���~�4�6Mgø�ȼ�������!%���|!����sb��|T��f*� 0�^|^����9�!��<ϰZ��!�b�_{$�Λ�˹��*�҈jl��=ȮCXs��e�`�)@}ނ��'t�,06������W�M���
���5g)�S��9+r��Ćŀ�<j��yI'�ҩ��cǓ�Ps��)c���?P������ �+�� QˎPgF�6N��N3C�������3m���Ѽz�#�B�n_J�yә5S>�<k�.)�+� s��V=��������� ��߮)�����"��f�$�|��Z:�����u���������6�ʁ;��I0�M�� ]�	�`�>�x1��(E��~������\�*�����LyH`+��f�}�7خ"����ə6�38"N>��������|��Pnonh�F���O�4>6:����5��i
w.��Q#��=O�qS<�ϛ�*�c`��{:��OV�����QYUCA̬�/f�m��odk�B�G1�I����8�v��|�$��L��V%�j������]8�.����hWl�!������G&��˺�����M������dD>L<rV#�W:��I���X���-V$��Q R-C��\/�T�W�4*�����BEgl��C��Ǯ�∇��:Z�Q'��^מ4,�6��̮'�rS������S�=Þ_Jd�"��+,�^�]L��c��vwt��^\�$\��z-Th�܂�{����.]4_w���~����O�qf1|M|pb�,���}�sַ����5�t��mr$�zv����F��
��ki��v�p��M�yއ�9�`��6��dP�����\�����J eG��i7�=DLdg����r;2dv��?���/D����{z��wz��A �'���UdɟS;Ң]���z-��;  ��IDAT�1�7��]m��(R���&���b��c��G�(���7�h�1�`A���͚?� B�U���tr�@H	��,������h�&�P���F8d57 u|�X�/� }��:Q�w
�Яථ���h5�b��)f�P��=��C�s������Y�*j6��k-�ؔN�O���wǍ'f�({�X{0od,��ou�>�]:0�p�� ?�Hד�p�-�.���a�t'�F���9��	,�l���A�H������L<�3��g��U� �^�37[|6	
��� �駟�?��?������_�)��>~�h�4��Q3Hi{�=e0��ή
Y��`���71+�d���.��NV��jl�ŏ?��ϥ���eC`�q��t>0�r"��>Їe�������A��� �
�	�i>����I����ؼ!o�n�!�*�D�i��`#�KKjܣ$Ll6yc�Pa�Y��0,�3U�}Y:�R-Tzj�eo	�����9���=����1��6�2�nen�"��W��K~/��D'N�	�����pU��h�����5��e��cQ��OL��DS��@G$��&�"�]�O�6���4:�QߓD!��ᢨ1qy��*܈�'���4���	���r��mޥX�)'�`@���/�3YM�Yj܃�Ag��9~CL�c+�� ]�׻��Ɯ]���D}P֥�X�g�������������^-m�_�6뻎ǘIv������	�������[a��Z��A]�}	0@߷x|S���M.m>z!���$Pͬ-��Pb H�L�z�{_[�')iy�iS��5��73�>(��e.�a�
xgF�.t��6|$R���l��^���	J�z��ӧW�I:�X�Q��N�X��ײ�>C)�)\�������(��S��U=M{P��<c3������`a�Y�L[���nS�;��͖���lmA�ގR��BYG���KZ$v�LR�'2#�8Ri֔u�[7�wv�0�����naq�jR���0�h���'�T�8�>&�`4Q��_C����|��o�/_���Dw���/�+��?�.�=v��m��ۅ}�c�-tr=ٝdq����w�R��oۅ�oTE�1���˛��7$a	}a$YF�%�gt����A	wr��9
��,�d	��SھR^-�l��d�}��}��%G�*�������;�÷l�_4fN%�1m���u���cp����Ա]G�6���p�#d��5h J\�kIa�H�y�?�ГW�p��:pˢ��,���A�S��ά��A��x|p�{�o�A:����8���4�?�M��F�h%�|��qX�I�3�p>lB]�BJk櫉�����|�.>��G�â�ra��bAG��6Y�s�I�S�I��J%�KG_��� @��F��ǵ���j�~��.�����/��?ӋW?J���ہ7��L��Us���lWm9��ݝ��N�����X���;�>-������CwC!D3N�eL=�-lr��"��1zB`1� �y�CB#�=:��U����w��T����Y��a�Ho�ͦNQ7��l�9��%=$��^��'��+��H�Z��/������_H�-`U�v�^��GJĴ�$"N���ħ��q5�v3��3��?x���!��V}Sf 2��	�=�N�(�s���^���x��2玲��_�d��U�u�{X7i�1f+(� �F܁̐�L����$�^W�)v�a0��n����⪢��H�]l$�ߣ���yk��8����n���{�*T5�f�1(-�a� ��/�����B?��[�L�n�:Q5����ו}T$��S�
��xX�^/����$�������Ŋ��5�#�D�2 �R'���9,m`0)S+ئ��h�2��c<�����"J5�>�6w���Hq��e�}X�����$��P��%���-.g�qq��_�du��_8�/�S%B5<`�2@�e���ܯտ�-j2$PO�:�o�#y�}�>�u5��E�&�ȏ&�آ����,��߬O�w>�j�]��>���=��Àŷ\�l�3�ήY�L�E�׆T��B֣&�7֘
:�f��I>�����t�q,��9�ߜ���˗�Ï?.L�N��n_�ϖ����w��n��#MM��2��\����NRrb��FY;�����),"g�o�`L�:[o\e�4���K��;6��hd7�d���}�	0,��{�w1��>�R���F���)����ԉ��L)�o��b�>~�����g�M ��B_�{��x��Rr����X��`�6VE�{�ۈ	Bq��!���;֍~���/ΤS5Tq�����w�1��ݓl��[����s3V��G�wVE��ӱ����^�u)Ooױ�c�1�� ꋗ?��W��3�?c��Ç��?�Z���;z��ɏ�O)�Y�z+������]*� ��x)̃= �%�f�w���|E)�"ꤍ~�)R�q{��ޒX��-%�	FUa�U{�0��X1"���h#uB+�W�5��6��^���[���'��q���F����ơS.��oi��5>5��9p�6'�=,��,Wҡ�b�(�)0/����t1����_����ckf���B!���ߺ/�Dm��I4�z��D���(L�8�j��Y�*���M��x����0� ��s����,�����P9���� I=�.��ͻ�"��{�û���ﴵ�/�����;1lqC�v���N������~j5~��^X�$"�^��Qny^��ifwS���'������e_$YK�"4�������~����'��r�}aHhu1h�Ƴ,�kC�M��u	k|=>����ȂT�~�Bš�6gr���N��ϟ�
�v�y�;+��VwT��E�j��hUh\�}��9E>�UJ;��� Z7o���LꮔG�h��K���uO%DɬwS����L�\uo�C'9��A�����{:uH��n32&UW9*��z���ؕ�`�>.�ݛ���۷�G�Y�v�;�������lt��`�U �K%R��i�&��0�ْ`��T+����>����Hr���.i�,�D��|Ĺg˹�%�K^q}6X��7�c���:e�
 i*z?�4��Ȝ7\�����IH/�3���b�8�1=��zb��pi��#���|�5���U"3�6�pD��B]��="�X��+�3�P��[��̊���s�P���.���3!&Q���Qk��θ���$
�a��2��J�G{�;���."I�:y z��i5�V�����ҁ�����fgڿ�ce�XYDg4��,�?,�9�b�A���}����k�Hu�qN�
�m�X���p���֮���Ǐz��g ��)�M��/���3�>G���?ο���/��~x�R�wʃ��.u���?Ї�=6�! e7��?Ej��C#�X�q��kw&
�$�tYl�p]�y���H�(�*Dm���|�:Y��6s��%%�g�ZTq=o�-]:��ʙ��@4O�z2\Y[��m8���c�1R K������)�P�_���1�(>�v-%2�h]�^罨�~�(� }���U�it؁^��Z���UN�]�����%��V �YT�X{", z����퍈�B��TR]��e9�[�=�U�5�J����U-��/��Y�|rӺR�;U�y`�1|�W?��~z���a��g�-�[z��+��_�B?/?\�Hr���Qˑ�;ֿ��Oɚ��eX�׫�(�'��zQ���nN(�p`]�K����A���t?R��6���/�	G���Sǚ��~���U����=��&�u�L��u�v;߅�0����U���I��/��`�N/���h��{t���n�������E|�&�ƹ�y��{��7�����
�ƺ�Xh�s/�E�_����O�M�z��=m9Z��ZB7��\���!�e�A�Esf�H�'��G�2ڵ�)��<T���@��\���u�|�:㴀�Ze�O6�I������N��@���y��ai���.u��r(��i7Z�!��g�-����7td_W��m�����u7s@�������&� �rõ��b�A/���!�a]��T���g���=3��Lh�	�4��q�Zv��}%9��0�v�R��Z��'��7��jx@�6�H]��F��1�kӛO"�P��o�H�:��u�ܧ:霸?4�ʈz�`�M�s�l|8ung��8��4ي����Eey��F�⯃U�F#��HW���j9eu�귱�[*�h#i����3?�S��u�D�QU��}GI$n��Uo*�_vYj��Y�iv��JF�=w��٘�(�L*��o/'^a���.�xU�����إ����
��`50{m��z%l�:U6)�N��j�D>�*6�`��T�[��Zt�@�o	��L�y�g�/iiڛ���Ԕ/>L�_Ʒ�a�i e	PͲp7���%n��Sc����<�q]@-&�z�� �o�
��+t�-1�W��@����@��XX̲$z�-�R�I�3�l��<!�I=)��m4�X�K.�����%�)f��%���ɶ����lm�Z����ŪX�}��!>�rC31/�]�� �g/ ��*Vt����V]��E���`_v�Z�^���}���C
;QhRI��4!K_�zo�������o^����&�/��-�����}����ꕰQ6��'��U�^���,��%�����$�AZ�=��!�K��ʄ@�c����e���ӉQ78��y���#"����A�w��g8g,�|ӹ��h]3#s��a�7�kWT��#��0��yH��IZf^�6��n4�Q��ҵ���dH�5�%K�T+-�PgMO'�+�qJʻ�T�mqT����1%+�b4��|��.�-aխ�m�$��?���o�cf�_~�E�0�����3���K=d�Jyd�w1�a�N���]9Xa���o	�.�n����g�x��J�m.9��\T�)	.�p<����^k�����"�Y������������ͭ�g�A�̏�h	T&�aK��K�,i��/�$�"r=��%�+�yJ$���2���!����1w��ԡ��^���S��8a���I�M��X�%�紞t���
p�Sm�+ �n���OQC�13s�������|V�f�'\�>-?�0�i�k~������O?���L'�dP�2s;j�T1@�������M�,��0sk�a:�����~_�ux����$ᓤy4y�;�D�ɢn`�_�Z\I�9����̐���׀R0��l��f�a�h�݆u�U�`��%����͎�E�X�+����N����<�N����n���"�k�o
�l�������K�������"��⸿���/��˦�x�Qc{x
��4ӽT@�͌�%�*�p��ټ��	\�YB��϶l����A*kACN����
lkv�c�LMf�g.��>z�ӥ�V�R=��ڤ1j�1�g�ʹ�{�R_�����uy�N�?� Y�G���_�C�:̯�e��'n#؝[�������
�k����ʜ����Ή6�m}\������H$Bf��Y��r'GՑ�c�xf�9K;�/׭|�#�!�[�^t��Ã��3����v��;w�ADg��E�?d�� Ơ>�Z���4��ncm�R*�f�|F*���	�g�LH�\a��W��N�$�f�E�,�|�*����|��#? ���@����~�о�����3�m�;�&����h���A����l����5s�	���^,��$3K_�����X��ŋ�!�a�G����� ���k��/�htZ =*���d����x%{3nV}�{(�rf����,�'�����Pf��}M���z��G���Z�G�D��Z�7Y�[;�S��݁?-���� ���Tr������ >g_��uܓ��U+O.W3��6�c�5FJH�p֮[�;D��?\�PK��N�U���a߀�Bq� |i҃b�{��ݹ��W0�>��R��u��[t��G�~�eb�Qc��	�g�"O���OT]"��u������(�L��לQ���<O�1����F3Rx���	�E�.�l��p61���l��,Ϊ���Htas��յgn��y[0���~|�ra�7bH�<�&*`q�Bl�)+~Z�]9�M�����x4-`��r,?�K;-����a����A,9�y= T$+��^6�ya�}BI���s�����d�X�ᨎ���EQֻI�թk��Ŝ�E����R��:�������r�J/*�	�,nw����uM$��s$#��b��{��(#���әK��O��~�̕>�W���t���*ْ?��1a�4�qC�}~�Bexb��9Wԡ�Owܙ�<�X�EK�^Q�"��(6W���Hì��󶋲RK��'
J�^7�ךg8��kdng B�9>�����T��EX����%��+}`�[�$;�W�ɺ٪.��C�F�A7@���Tːp;�Z��������0�0����D)�(��R��2l!{;�Ja�8�s}����̢�Yg����E��\r7��X�$B��a�Kx\��8��r?��A�'�>M����{��n ������Tn�\a{v�ɒA����H)8����q�.z{+Ǽ
���J�sF�D|ͱ�ޟ�]���c�3������=q�����2���Ó��q�j|<��4DTm��qmͩl�vY�ۦ[0/pI?g���j�?����P���ލ̊�`�`q5�N�ͭ���C�P����Z���t�I�?OC���g{c�0���w�_���۷�����>g�bc��t�d�5y����S��{jv�W�u���7���\��o��￳�� ��L��4j�>�;�/���4'K�̌Y�Q�$�nj�3�dvX�{��ӼF.e���a��y�d�=a�v/��(�f�r��]��1�:�N��_��� 5�'�4W��T�r�6}F��(����`�U��yR=���${�l�C72�O�??����.��e�'�
�-��M5��(k�K��U[���ナ�K���Tn��1ES�9wf��r�ׯ_�o�={���$`���+r��{	�/�6)��M���N�����?K�(����L߾}Co߼�2)�3J=�(�nn&"[�@3��T)�E���Y�1z���m��=W�[�^Kd ��@s�=t���Hɧ�X�}�`sQƖ3u����Uu��й]b���n ;{�r�+����W�~uP�S Uu�%��I��'˖��?}�׀��س�n�%r���%y10k<�iY�d�-щ���r�[�͵����{��[�p����3��I-��*c>���|�������X����c�z��-������/��ka˓뢊e/i�J���o.Ë߾yK���?���N2N��?W�����`�ZQ�e`��S��bs�u9�)����wz��K9_\θ��l�|9��:�[�>�b�$ђ�(`�[xC�T#�jUDo$�JuF�8��k���G��p�S��L����F)q�1Cc6Ja^�iJ1���\#=����Çq�z�����^���r��j)��!EOs���g�q�����K���h3Y�Љ�_f�r�P;BG��)�2�
S�O��;>E�2��5Q�9�8���_n�s���3sb��W|)�k��b�}�å��`]��IJ4QI��L�p�����޾}G�?��$��,�`�����x��Փ1V�C��ϹPQ����������"���0�����=�%�t�����GN�'b��������n�Z[��϶�h[*�5�2�@�sO+}b�0�f+9PA�~�z?�:�rξ�N�`��<hU+�Y-��2y��O��IU���XDV.Q90�먏Ɯ=F�&��w��Կg�����|{�ABa�#:���B����O֡Q�����B�M��������sV�i 3���a���\i%JX����g����Pa�қE�eQ�l:c���Yٷ��@��,�KUؙ <��G�����TU7#Ts}/Xi�zl��x�)��$L��y�LA�c�=�75�����m�ע�e�0ڽC�hφ*n����񱱠Tv7���X��oLdb|�R<bh[>�]��>a�$�I����l�ɇlBEY��)
�����/�Qr��,f�3ʦ��JV�6~�o碠�Yl��RhC�����QNfN߄�Q曟s��>Ѿr�w1AO����O]Ӟ���t�&�k9��ܥ��
���8�/���-i���k0���j�rf
�vR�7iȺ��=ji�ٮ��T�c6�믿��k6gIz��6��ɽ� ��4x���쁪`40�I����-l�/�?����K�Ø���~��>�ua�N�,��j�%_�#���7��]���h�Qo�YQ>�f��}N����2T��k)+�^X�d�@�Ռ�Q��j1B��L\�,�ڴ	�%&�����Uy�j��~�L�":�In�6-�cH)ARV�lPxY, ��s���Fj@�w��f'��򳡳�w��wd)���}�����L�ͩ:�|��x��O�2��d��ku�_�=�_I?�b�:�SP����s���>���P�x�Jl����q�Ȑ�&�9Z�Hܧ��0A�hm�M��)Q-��.V����ۖ�.5:����q���'Θ%���Z4�h>�
�R�u�G'q�7�ԃ���8�:��S.o"%��/r��^Q�����hY��۱�b��i.�acU�,W|����]� k��ހ#���0vnR����b�o�H�ctPu�V��6�K��'<2N�I��4g`�~�zq�]���9#�qH$@횈�{;ʥ���gx���]f�eP��u�r��N9́8|�1�Z+�~������zȴY ��j��&sC���32H%}.Gѐ�w;S�ӽ\�`~���=�u���Qf�a �f�������f�����FJ�����A�\~�H4ł&&���8��fY�A��E��I�|����8_��]�
�^PH3���ndH�Dv�&Uu�j`����7+V����_�=�V��+~���\�["�����#��:O�U-�q5A��u�llj�pi�r����z�ێ�R�v�pr+P��Ƥ�a�t���8��� ���>��h��x�l�*�{�|��u�Ϯg��.�P?u�n1:r`���ȹ���D��o���;���
@��#?"_��8�]�ɝ�'�	��C��AFM`\��� �=�wM����
*���O��f\3��,�}4�1����r��H/��7��x�#n�'�(�Ժ�y�PK�(`��A]�` c�Ȁ5Ih�$?��@�N������obo1F�?���r�j���[���-V�Hf�"Sw+Y�Vtn˯��|�&��fŒ2p����\�e#�}LC�ס���Q =��� 2�VuG�{ݯ	���/��,*�{Pݱ��u�d�4�v�@�����}��ga��-�`���Q�ZA8m*ד���P����;ϰ���x2���ԯKyt���LCN��3��+�3�c��� qy&��
c��KX�ԅ�9�c1V�(�^���t��#�]4E?�Ə�f��_eD,i\9�٠_;J6�f@��i�)oV�ْ�0��uH�
�J>��w_MSW}u�lX w�g�SRNS�V�
T��a��`ѕ|��V7�Y2��e���Z\����G73�f�O���	�gҙR�T:ݔ,ξ�{.�ۃ�yJ<�5%J^2��̱�#���.�#�fdӭ�i����O?����<�-��=0��)���5���wǺT�5��_�����lLZ���L2�yR����4��󎧏�wq��S�IT�@�IYR��9�2�_`�1���c�P�.J �N�v�Gݤ{�v@'�N��^?��=#����ǺV�e'�ɬi3����1=��Є�8��c@|%�
�W
�qi���ZMdA���`�q� ���&�*����X����Ⲇ��ߩ��=��DYч02��F�l��2�-Z��P��H�y7�Y��� �32�g��bQ��u�7�к��>zUU��ꀍ}��S� � �9����W�/��H�GRBہ,*�J�E�9kRdۘ�*���.�<��~c�Y�\��x_�|A�����^RQ�i%�<o!g�O�K	�����G����>1*��}��(k]r���>ڹnkGM.9�Y���6>��&"��T���uTRjg�S�;�������>>�k�T{�_���P!@�(��.��	����T1qb ��H�`��`�&]�<����}�>U�?�7���~LBWg�G����h4���~f��U�w�R�s�GQ��~����,P:�6c�_A�\���>G{z�'%7�eB���r�J:���7RD�U��VM'��
���u@��u��N�d�P��3�U�~v�7��J�/��l���3f��Iz�㉜]^��N�?�29
�?��ӟ�f�3�����=��SW��b"��}�I�ɔ,Z�~r��	s�u��`Qg���5�uDu��#��K�ʧ��KٖK
��q��,5�zc�1V�bg��@i��1rhC��	E�YcsDJ:QUxi&&V���䉶E��ZqcS�a�~�MR�'a逃�"�:���q��{H�7��؞�@U����P'��M#"���)Ƴ��@�C4�Y�]�$�?��ru�[M=�H�in�}������[�di|�j�⨂������y�߯�Ǐ��PO^؟��_u�X��=X�EsN�����"N�V�����Qt1.̏��f=���G�ߧ<��2/�Y�It���>1d�	9ky~�P�"`(���rR��st=��� ���	�ì�>��iP%Wqh&��9�e��1���� ��@��W�
Ʒ�����"�A���V+��J���0ZIy#K}B�|���jE֫�U`�`��r͂�����Ү��()�@\��6m���Z�+�]����ck������b����.N�Ǉ�o�/l�WO��������εU��=9�|�~�ޕD�p#á�5)��gK� Y���6�e���Ա�H�<���}��>�S=��jē�9���J������:�&���ۄN��a
�����Uݨ��Z�?|�����J��p��F�9nY�� *3�唽��-B����������b�c܂E����Zϻ�`�FF+���|r��ì����c�4?�,8aw5*oJ6�Deqa�mf!)�{2}���l0fjnT����O\��A)޿�:��CM@
p���y*��MJ}P\nW3%�g�������(�P`u�D'�W\��틸���>D��}q���fBz��,��U4�����L&��Wύ-=�bd\4�ڨ�z���ٓ��)��鬟�l;�5��fFn�C%�dȚ�}h��Ǵ����^�Y%J��ל�폢ED�G�ݭp_���ђΐ�+!���e����v�����*k� �kx�H	�5�v&�Ƙ�����7�fٖ߳I��c�Y��-Ue���"ϭE}yt�%i�"�+ï/b�_A�x�8���~��.�Pb�W����(�n��t}��>u��K��|�B�c}����x�/�����k�|wV@�o.�Y�	p��Յ,�B�2���,�0�M�ϲ����A��w��ʠpX��^͢�*ڧ�;��!�T�E���'���Kx��Ef�&nw�( Gv��d~��(��+v�}*[����b�J�=)�P�5��iL����������)�@Zn}`���^d~����Y��D��v���j
�t�S�<�^,?�3�����p5CʛO �݁���P�4D&=���5g��3��}��ƀ`���w���/��ң�vح�-$� ՏQ���~�*�av$1]�Zq ��E t�ł��r������m#Gͭ���,T�OV��b`Y,� �Z`j���~���;�p�I7�'zţ��2k�U ���-�D��-���I�zo�*�I�>�ǫ�כ|㾼�������:ՓOqL~x%�c��U���c
��_�Ṯ��'p8n�A�>��r��%�}��M%�;aϫ��{a��7f��r�e��j�z�p�n�e ]�G�t[O|Ĥt!D`�x����hCAu:�;�`���5���L)g��E�ʐPC��7*��^/c��5@��9E^u^��SO
��0��ȹ~��V��&>f
p͇I�=�Y3E15��A* �½�Ĺ]X�����ˋLu�?x��V�w�`�G�戅^qARg�5pe���Nic�)�ЌY|
�Ւ�=��z�|�a�@�Il-ᓯ�USӃ^��>�*u���@z��������*�"����~x��;��s�aB~�~��PĞ�ͦ�zT묊��NM ) ̟U�%`5nXkZ��b1.�Y ��tw��'� 	�:�r4 v�YB�57���-RI�6������h��[�� ��O�r���N�� �`��R�����>O@����s�bUC�%�u���3 ���D���#��x��?R�@YM�yN%�*���<I�׻w��Cl��Gv�-0�=�[Hx#��~��4��������J`�'$ ���u�o����!Ɇ��?��a�<���|?���eӗ�N��~��s��X���?n���}�0��߫��I�Y�a�
�!X��ܱ_�������	o"JO�@]�LV�Bd� �q��u�7YL��P�ذ��?�����|�H�Y9GE�":b�^nû�k�D~A�c�tw}���=��*L��K��u�T��栏sX'���\�K<,�Cƨ@j�C��Kw-'��u��ߎY�&+���v^���񍒣�G��񱮇?�/۾�X��L0q��MpzI_�F������ǧ�� �:�c,��,4c��1*��g�]f�7<�X��Lf�𧫓e���ȯ�DZ㪻�
��,2�����ߟA�"ƭEyLm1�3#t�t���%g�'b�;T�4;QS���U����m9���bO*1M�|�}ڪ���_�|z��+��G��yXj���*�-'�L)MXa��Fɓ� ���eSDj�;"�-�����]�D��f���-��2��2���ܩґ�蒬�h�.}�X�1��;~ן�>��P׺'w��NnL	��z��ĳ>B�+[�VF�փU95������������ɏw����%2���㰹�;�?,�$(��%�>��zS�(��"��ja�E�+�v4�����P�6+�B͢�����bg�h7c��;d���c�
:�4�<ߦ�9�YP��3�Vu%��9�S��&�ɲX�վ��α%C����#AT�=k���۲��NR��X��,�ME��nj�R�h/ύ��60��/b���Ħ�����̲�H�,�l��n�~;rV�㞞��ԅ�a��.XE��J	�)���@�}x�3�����y���SqY�]��I��: �q�ń�[s�o�q�z�@����m}<�� �ݖ0�N=|3��Rz/]<�$Q�fYTY�k�%2�%���_����wfӗ ��t����C�U<�=��t�A��ňK���#�.@����PEN)���A���2����	�݀(w��=* ���0�y�h�R��Y�T�:U�)�S�V;���Р9ϯ�G4�1�i���|R�����o7-��T�!�����qb�c�����
_H�C~U��x83MBd79�����2��v�5e��)���_��K�)��)��.ǧ?2I�G�p2%q�0�Q�����KWL��)R>Te���],L7�2����h�}B�}�s�R�Y��/�5�����;a#�F�r��W�~�ϑ|��y��+��n�?U؆�]|�?��A�&�\�S֕�~������TA�vY�p�W��)e[+9� �s&j� @D��{L$�/i�����κ��	*��k���'��w6�8W�|�K&��3#�AW�k!q �^���9a
@�L�ik�r�`� B���|��\�w�߸��k�R.�Tӳ����7+��d�Ғߞ����A���Zr;9�h���#K?��y�L�W9�����t�H[隭��'����Ӑt�,`������tE�&��r	g>�ml,ᆜ�����������ʖԽV��r�n���DO���K��e?���i����}RmF�Ҟ�K'�F���CP?�Ey�h-n��1!�?D��?9�������f񎯉�P$��{r���@�[� �#z�e3q�#$^.�H%��qO=mPWy��O�ِq��7�,z#�s���L�� }7��6.�O��);����'V��g��ʫ�� �Q_�M� ��퀚k�b���E.���)�?P!�gQ%H٫$Ο ���=��Ņ� |����3�+��`2�`@����nv7����?泻{�-ٗ� �9�ɘ'e�*�O�!5��ds1#R�T܆�`X�X�\0-eP�!�z�v㌩��'�����T��i�(�i��4]i�H�LdN`{DTs�I`�Q#��<�H1@�O.�X�o�6�:$�i��4} b$&�~����K�G��e+:��̐G˴U'O,���"ѓ�-�%�bc���������BfQ?�@�-]��f�1��zljP��Y��!�^���:��'2T:�x=���|J��� <�n0�̷͵���c���b:���ݭ���ͭ2�4D��P��O)��"e�Q�2����8]>��m����fúZ�[6�-����=Gˈh�9��O=r�"��(��K̟g�	���( �^'m|%]�D���q�H&�~�̾�l�r���Xn���z�R|�������4��>6�}��*i�J�!���ƚ��D-3i�1]�Ly��d�X����:�<.=��ke�`Hk	�\�������z��+߮L��4j0�/���D�Kb��"�0�>��������a:����F��|�v���$�8�s�Q5���
r[K?ǌ����#(���Iۻ���s����gi��Ǌd%��Qe��
�ie:Q����L���D���e��dA�i״�����f�� ��f�k�N�_�~�>�5K�޺m`O�D����w��6�� N6W9P �&�sT�Q	�-�_���9�M�1�(��\�NTF0<{�c ��&RN���Zǟ�P�� ��.��b~O]����O�:fz��s´�t��Nf�� u�g�5(�� ���%�6�* 'T��1�.���{z��%�x�B���۬�*߱(�.դ�Ia��[�QwWf�q�}�O^�C#�u<���	w���+N9�Y��>���'jy��$�4��\��x��}.IOˇF��m@5%�FI2�[��(��"�5F����=U�z�0t�14,�á!}x�Fi������y�?Pa�]������l�����E�(I�z4/�񗎳���I�侜v�f��]Zl�OЫ%#)����r>�P�HXd�
823�������_~@��!XX��#Bҧ�s�:B �t�u�٠�li:6i|C�j �BD^��G�y�\��w���&�ɯo�i�V�j`��$+th�;���5Oi^]����GiCT���}�}�T�(���[�|^<'k\��7��7"OQ�G=��p����Kj��Բ����d��P������b\�x��D�q9�%���<������/}>(�NJ��8ß?�>���]�R���d-�.=h�V�dCP��L��X�>J<�֕Oo߾���rʌ���	��/���T��fʠ	�������s�����+b�a5�j%���SN�~vm8���yx�+j� 0�<?
%��&���\	_ݒ��/ �Y��Ӹ[���.~��������W��@PdD��"�Tζ�4o:��S���oQ����-x~��y�+��XU?�or�6��G:<I
��'�Kˀ�s�J�� jZ@�[��2����y'�vY����6�˄�1�cя��iN�j�l��[;av X�-�F��zo�p�8�c���$'��o߼�)�΋+��hb����={�̷zL6�I�j�h�:K�;�뽥#���� 9��p���}/� �;N�fϤ��0̶�'�f��:�,q�Ci��+�5��l,~2p�� �D!��}-5uX��[�ꮝ,�b��,���K0>�M��&Y�w�A|�%��vc:�4璔��nH@c��^������؋��F�{�=�̇�)��J͛��
��D��tu8+o=e��������ǏO�����r�S-,�`'�]7��y�V�m{�PY��G-Aͯ�����8o�1&0�$N�?���D���S�zޏQ���T�ZB�����z�����>pdmy3�s�[��"|	 ����	,�`[�D����Q�p�XSZ�k�I�=U]�ⷼo��1^���I� 0�<,磦d,�e%�՟5����43t����q�?@������ۖ/�S_��9�o��#�/��`�l���"�3��z,F�.g��Ey�}^<>L��޳͑Y2I�i�[-3ұ�ew���ؽs�<�̌F-��wUE2�x�!���"�� ��L�D^��J���l�L:�q�_�✮:�b�ȓ���$��"8gbg  ��=�'�E� ���<��>w������������ᄵ��#'~QΕ�}3�ɻ��5��
(�2w�=)��A$Gv]�̚.j�@��*I�U��w,!��Z�w��s�-�Uﾞ�L�o����q�u�?��Y#Q½�ſ�&u�m� �t��̂%?�ڀt�6l��QL�Kb�닚V,�w6®i����f�-��\��ȋ^v]�����W�U�������[�k��>�]�����?���]�K�G�\���8�D��s�e ��ǥ��f/���HX%�O�
����-$���&G�A)���e�R��ԇ���D��h$*]\8��+N3$�L��'�7�N��H6�E�]%v�.u��x�;��n�[P�~��B �/�N�e�ҿ��V�ڕuV�O�d/;�[��֠��X����=pܾ�:u�⅍��j��q��q�>��`��Vt�׳�[��zz�Jm?�,V�K;:��%8�;�� �������]����S@-��ۘFX�3ڸ�_��X���q1Jm֯ў����!�\�ջD�z��G�T�<����:�Z�iT�&1��-4���%��ZJ	g�+,.K�yU�?��E���G�E�:���&�7/����5CN"FQ��܉vq�if|o���>/
�p�~dR�q��Vz��DK�?�zgl�� /:Y_�[���������/�t�z\������ҋα�?��	�L��Qv�>�۔���i�������Ƌ$�7��m�i�K��Ns!h)J�c�Q�p�������q
���_ �PL$y����&-��G#i���W��-�F�j{?��J%��%jKh�[OW��g��*�E��1�W=��Y^Ċ�I�/Z_W�S?����z_�zY|��MTc�-��.ʨca�vD��4բ�}������}�~r�a��;�Kj����(h>E�"��l�zS'��<����P�rM8���]�b��M�d�*U�\�D�*qS�ʥ`��a*r�e,z��_�
���� `���j�(y��S�C,�~V���!V�-�B�\�1��'si������z_w΀U��X[O��\my6���>йsF�a�U��w��@exA)�3m�R��g�/��rS���.e���0���V۽��ۦ"o%��ߪSu�J9,��s�������i�ZOt��;ʭ��u�'�R8Eٳ�>��5�T"��}���ߜ(�D�$ǝP���� }8����p�ݟ��[�Oo%�fx�-��9 ��흹M�a� ��yi���7�C���h�1����u���Rur����z&�X�Y"򤠴���"V8���)w���z%�����G�k�)Z����H|�V�}�0D�\{�Y�r��6�Bm4&~ѿ9՚:3&8e��l�`�3x�4S�ip�XK#��������p�~���K�W���_r���&� �:kgƭz]���xB��A4�Ȫ����U�N��p3���	E�rS�$=��~�C��ȸ�q�t�
�����_�o� ʡ�s�h��R4O�ў{�:p��T/�:�LP��V�<�z�Z��uJ��_G��K�c�0ձ�Eu���1Pm�G���M����ZZ�͋����=�?��~~3jE�:W�z_O��8��(3zy�+W���6
���	��h �sp�s	�d���DeM\&J����<$�|g�d(�>�FX��<�Ӊ%�N]o�w�m��f s��:�Ps�)H)�Tq�|���nLT'2f�w��Ond"q!����n��͸��ӳ��V`n
\zlR&��Ts��gi��+���VM@���uۖ�Z�Mp�Z��Ӊ�5|=�{k���jYNwv������"��r�_�+��U�➰Sn���wܙc�9��<ƙ�59� ��Lq8���KE�ѿf���b�4��^D����'����
.O�b�\V,�>�t����@R0h�����i����6ս<�"+���[������J�eMhb�":U�T��"doL��hA����@+<z@u҆�[lwIeT��S��[o���J0���/OM��?�#�"u��(\�tT��t�oM�7���_�E�^++��;mQ�� �s=�;��>'�mb$3cA�m����D�+q�Π4d3�/�0�h��0�>4T�nT��.�I�'�:(@��iP)	H�q����b@F���N�����њPK<���ɽ('�,W(�z�=O��u��nME�E�?v���*P�s��U�����DI��!�h�Aoam(���؊�1����Ƥ{�ܻ/G�@
��Sq�aw��M���)b�r&�	���K�'0����|�5�D��r�JP'v�&�'ɍʾ�|����oI�V&8�Q�S������Mp�Y��8��{0���b�n��(D'���,���C_*˾�J�(`�8�)�q)I��=}\��$�	:QB~�W�a�����u��c}�@��?����-:'��z/�T���N�o��~5<��Ӎ+Cڗ֔��K�޽2� k���LԸq;m�V��6ʗ����i�!}A�-�+���$�L�_"j*�ᷖ�hE�F5�����0iZ��x�z.�����e7�h�smk�G%"%���DMB��X�P�zhxQ=()%P��-.:�yQ.��S�#�	�:��*o�g��U�n�X�t����a|QA$HZ�f3� �"h���X4��Z����9��U���T$Ne�_T�K!�������Չ�&�s�ٽCu�V uпX�D{�U��X�ݤ ��D^JvD�MS	(�8D��w���;7����m0��+��I�o�&��Q;��Q!��DܥZ�䯓���$���"���4$Q�%a�#y�s�8M�K�!�Mg��	dLyB���O��HyF�+���u�<Ȟ1�1�k�~�g��4��g�"��m�]A>��:��^��q�~�7��n7�� �w}eѾ3���vY��;\ >2,��'U�� �_hfuA�k;å=��zC>���S_�Z�V6ǉ�c���
=��&��F*0Ÿ��;h[T��������_�!�"o�P�_���JD�]��BpǺN@'�}��
�ׯ���n��DW��/�X���B#q"�B3�}��?G�ڵ��9��T�e�R�T"�d����u�yQ(����N��Lf�D��M�[P�Go9�Ǯ�,��y��z�t^�ό)=F�Q��x_u��w�sc��E���r̀C�k7�L�~=G��Eْ�m�y ���|��]%e4�w_UHm*ѫ/5O����_�2�9���s\1H���4��|>%Z<e���ʸ�wk'�иN5���<�4"Q���[ؘ�ݺ�o�W�ǝm�rV�}z-�n�U���+[�s>�>����:Z��x���n1B�<��'�8�9�\"���
��&��V1@�����H����U��fl�EU���GV�c�(k�?$ջ���|=X
���B�p��q]$�kt\��r����\��9�
!6�X���<���N�r�|Ba4�++�Ή�'%
J&�iBK��%�
��\/��\
�k�Sq�#��ƁXgpE�n��h��c�]*����z�7�y��#�h�7P;��[�So�Ͼ�_�ѻen?����a�x*��~�ƺ'#t�oԘ���[�{}"�aQޥx����ʠ-׈�6S�X����}�f��>圱���>n��0녥�o�xT�����Bsծ�������|yR������~z}�X���X=h%�����VI,�>�y�t��uy�xޛn�m߱_���5w9¬z��y�q�	56����'h0���)���Aa�C�bs�j�e�l���Z�]H"�&�b\�ߏE����?
#+|ӏV�~9�;�D�(�4u�y �(���>8(���cܮ\IQ_��.�'F��N�U-
�׫A_�jI_�UY:y2�49P�g�ݴ�t����q��(�Z��B�[l���=�3`��dȡ�}��@0�l��C�?���*���g@)�`;�a���y�FN���C1)��I���Kt��H�Ro�0�S�U��+���)=p���{,�g�\]�~�
h��9����2���{�_���c��\h�d�L�\��v��<YsA�����M�Q��:_��x�P��ʝ����{�ש�C�����(x�?=��bR��	��}����z���>�~0E��P�Ϳt�fzbԕ����Qm�$��[]�ĭr_}ł{ZG�<󹨻̉j�$�����H�7�3��� 5�R#,�{V#�i����J�^�6�����W�icE�z�� 1�!q�o�B�^$֖<��I){��V�PD�N��"\�-ѾxP�3��To�i�%zXyVG������x˻�r��w^�wᐼ���'�6�>
���獄���b��T�aS1	qp�O�>[����a�U�:���X^ZF���ڇPQ_�[���j�&挋<g?�&'8�
0nR]���ל��x,�CUˮ��װ��� 1����µ�oiI�7��j��⣣*�q�3�ܵu����`�?��;���2���W�S���|��,�o�8����&��=X���sDs��#���{��\�?�QsǺ�"V(2��PD���q�ol��c�r6��=��:��Y_:�G<P�\�n���cl�*��)v�q�2Tв�)���nK���Ձ�X��~�w�U�vܔs��v�=i�����&&�^�1�_jϳ���:��E~�w1:y]���/nb6�(\M�5�f!9ໜ��e0P��5v\�;_#���\�x�ۦ,>�->ɭ�Q��ɺ��No����8�z��_�x��ED]�F�R:�=\5q��SZ�ܫ'�@4w�W}_%!Uꌾ�?�g�@�cǈ�5@â�]��}��a"vD.���K>R�wYO��~��\����2��=6�M�fJĝs�F+�ôfQg�7��֡�R�$moM�s���{�RFn:��l����ܘڭ�����{�����q;n���I�]�ʥ�d��]W���=�����~Vå-�3ʵ!��yu�>[5��0�	v�[}_�mu��s�x�:�/�C׺V�(J�ߏ1�[��7<@e1���k��F�;j���m��LK"�Ƞ�-Ke�{��f����S��'\�����z���ޙ^X�L5NA\E�z�5�}lJ�6Od��r(��@������+8!�{ml�8c�(H��8����_ O;vd[��,)Lk�;�rO��]�7U�v�g�y��S�=��*ef���5��
�j��,�I�RF�F����.����>���`��uG�|@ã�s7��[j
��=�O(�H9�d�(���LF�lb�Q-\n��ZVޗ�("`�~i�Ȋ~��9qi�N��r��HPcq�n�K	dK�"�����i�lJn�Vg�^�R%�W�N=qL��\����J$-�}��T���+�@�^��6�
��g��~�A�Qш�����n�x�^ߓ#��� ��62N~��CV�K��$\�hW��1��O]��O���Cd���G���?W۝��)��c£�+G�^�����!ۃ3nU��>�pD�k�oĤ�ͬ�:a5щ��:�a�i���'�f�׺O��[T�v+�Sݩ����g�K����g�!/�WV+<�ܟ{V�w�I�^��1��\��>8���q���]�k��9W@\_�䡭�N�n$5��B���.^����Nr �A	e�g*}���F�J��]����$ب�0b�҇�Q�^�;��0u(y}^E���gLWm�E�*�V�7#�#�d���wд$0ׅj�� ����kq�M�POp�	ݜV���1^����-���fQ�$�8��z:;#"����9BӃ��=,��(c�ǡj�޹d�tPW���s��JU��$�6N5j�¥֎���E�MR�M�����WO�����W)-����6w]c��T+�[����|M?'B�Y���ÍYo��`C�5�Y�Tʋ��]L�0P�����wb%0�J�[��s��E��L�}���>����W���@�h[K�i
b+���x����	�g�	��K�;
f��8���t����m�(مl�4����"WO�Qܘ8��a�d�v�B�1��+�!CD�L��} <������τ�x-�>�d���R�����{Ml�W��ӡ�g1=�{w�mS�t?�e�Ux|���V$'87Y.4�m�6�a�����z���"Z`�>��S �R��R�ґ�LTeP'?Arm�^��,�v(!t����*s���=K�0���Đ�MJ�%
`�Z%a�u3V�k�S�{s%\���]=�Ym;���R�59DF��/�B0��T���&�M:�t�^'���^J]����&��R�_�O�
 .�iee��K%�q(�G�=?��)�y8��'�Ƨ��ކ��^�w�X3(���C�Gm$M_�XAUK{p�o\�ܫ�O���!�M�n ^��F떄��2��-[6�Q߱���<����2Imژv����y���7�}�Ǹ�Ҕ\l EY�C�P�"�Ƴ����쯡��ٲ)��Dّ�R�vږ 5Y�G4�"��_l�q��p�DG{'�_d1��}���}�b�P���8m�|4ݿ�~�:�]�0[z8�6��݄�y��Mx��yx�����ٔt�L�黯moc�j)��JvPu%���J����)��)�6Nʪ���9�}hT8�{�Wذm��q�x�҉�v���0dc�\S=f*�8q�c�X���a??��4l�l*��ծ�PO�|\kۗض���W�X�vPrd$N�k�)u�)��� ��P�b�D3p�	��+��c)Is��T�^���$z˻���E��4V�^��/���tvp��{������ɓp������c�Pg�=�J����.RK���r���j{���Kq�%,t�Q�u�k�6&��-`귝P��j���z7�aj#�[�S/�6E��/<Ź]�C����a�o~ʴ��mz[Á���i�ѡ�D�.A]� �Zܹr��$�-�]K��DK��Gp~r\���N�X�@&1,��B���4�r,r�"g��&���L�	N�DS��'>A�����w�����>Ϟ=#МH)5<�=+@5(PV�����	�U#N�.ba�L���u�d�{�3���f*���|J�|��uZ_?Z�xA�EPF��1@�wN��ΥT���')��n"�[?F~��VO�s���Y��LT���
� �tR��O~5L��&%�y�((-�.�l����r17��Jd�L݇*rr�{�y])1lr/�{1��||�rI��0 � �s�&�2�x�X�g[p��H�K���,��tt�^�f0($3��S��WN���-7�r1�� ��~���K���c��`"�f7ٌ�-�����n
��O��w��HZ���{DK�S�0�/��ө"N�.��Ż�Ho���m�.է��:0��P>g۲��P�@��7o�Pyߣ����[�{�9�Y�~d� �/ `��O,�(�a��T1�?�s��	D���\v��ŀ����P�@ݢ��s�|MO��e ^Ȣ�����/��W����}�ƥ˗��T�?�T��fL��|Oť:��8[��<��Mu�i�N�F<�d,���6}>~}�6F���>��:)P(��Ѹ40ũ�Ե�~�c�gj�?}�Xۮc
�%�!�-��f@=��������ի�>o��{�><��|���'�C�N��?����9��* V{��uˮ�P�oh�,�ͪ�;�cݵH�V��Vr�p��KZ��6���H�D�|�F�_�N}�޽s'\�v��O�U9oT�i$�2P�(I��J����6k�quzJ����,mد��s肴ɳ]�f�p#�Y%)���w����w�~���-�z!���<"�h����q�4�T�����})\��c���L� l1�0��\��,�{�.���?���>��dN�$s� �y�����h<g��A���|S�#�d۬���tF}�cُT�9��9L<��o4��0��c��$���0�!�Sz��S�����xx���1V_�u�v���[��J �V���"��N�2��e�z�Ę6���Ʒ�,M��!���q��҆����Z������sz5m�V[�.U���D~mc��9D�3[L-k�_�n�ʯ��J��? 'X��"uppnݾC�I-����(�������l5��@k�Ne%b`N��Z����q���RUjıP6)�@g����q�網��@�ntJ`�J+��^�.]�k��V�$-�>밚.XU�t��O�d<Ne��m��]����:��m5n3�e���Q���T��71sݦ�H��@��t���1;�b����ߟ|��o�mPe��U��p�3�v��Eڅ�0�t}&�%��/&��s���Ws�W���v��k(w��}�Κ;�{����T�!�S� LM���{G�c������%�B�~���\�?'Q���DU��Y���S�sV��V7�69�\{6�O�����6c��S��O�vw�=b`�T�F�o_��]�F5���b�&7�I�g�����m/j��Z����.\�@���ǧ'=)�V�:[�= ���NA�sM!)��+��@f�|�#�t�$)�8��Փ׫�hsÃqˢ�ŧ�`�w���\�����Xv�RW,��� �����sp��e*�gN/�L�fT]��(?]뜳���[�Ul�8'����2I�D<�f>�6�v,(tɬ���er��Yѥ�<�ꜵX~W�wr{7V���c�S��|�������8Ԩ�9�X2�g����U5�)����u��Q�_�8���2X8����-�$pSK�.���U�>U+ n�&���K�x}��4��.���-:S]��$-�1H��} ���$'ꮅ+�ϰ&��� &��z�֣,U[��
�����M������*P� �I����Q�6�G�x�QF����5�g�E��������t�u�G�qSN|��0m�AtX*LR(>�^"-N2�`�����\7����(o�(%��θd����������]	'��Lw������Rr<��{�]~�N|�i� 4�����c�(P�P8pS7d�_\��X����425��F�0
��V�K�Vw�g=S�W��e���~��o:4�	�C<�n ���H�u��5�W�_DGƤo�?�%�!�]�W(������s�>@A�mt夵�$96��f��Rn�cy��E@MC�WiMW�S+�#���a-/���������J�ш]W�MIl��k�=X���җ}��
��c���ݘ��تs�1��r^r��'l�=S���v���e���>�{f��1�4��L�1��%�2i_C�%�n�mJ�� ��^5�|D3�g����,�B_�t�Nű˾���mYAП�U�^
uI�?�Λ�zQ�������ǥ���4z���/��Y�}1�V��G�e�/"w��Oa`)���ʦ�j4�Y�~	�)��a.�/��De+�;�W�mZs� 4�����7y�}P�M`�&}��U�+
w��f�D׻�Y{
AT��cPk��48��mk�J"�H�ʡ�I��"�cZ	�&'ڦ1�U�������l�=���m�����ݣ�S=R��
F㌶���B���1Nu�~��c��O�=on`���2�=�Y�k��f�Z��	�j4�ax�3g��}�l]�O}�߶�(:0�3I}�����"3xP��8
��D5�z�zc��~.@'�
�t����B��ڧ����ԸV��(�Z�_��͋�!xZ����FO��l�
&����n��έ��2����ǵ���`j�iϿ�EU=s�<�T7_D?Y[���j���V�����|��m����(l`*�j�h�7�Z���*ZL=w7v�9�q�A��m�������yUK�㪃6jt�f�/�i����1 5"O,;m�����W/G:�jSoУ�!�*��۴�kL�3OX5�[M��B�6�J"�����뺱�?r���Ʈ�y�7��z��h�s?c5���_�M1o �$�_�_VO���ډQ��K�a��B�t�n*�9n?9�s���h�Z�\i���9�Յ���K��0z�x�o&Jo1�w�#�ڞ�Zmc��U\�*Q�wz��D�I��]��Zf�G�5����v�M߇q��ES%�(�b5�}j"��e���	���5^��U�]��	쁭�M8��OY���ȯ��cpˉ^!��F�����0��-��W�-��e5���>��U7�!�-:V�-�=��?��h��]�R�5*X�Ł�Yȹ�;h[T߬��Gx�l��$�U]_�n��=��G1����U���0`c�� Z�r����\������~Ζ��j�����]�9Z�GsT������]۾�_��y��������&W �G�w7�O��+B<>\��JN
�(ɺl���������vnE�J�̭vvm}N�r��+�0�X�Y��� ���eA��\%-���q��r�����x�Z=���%ɰ��-M�O��#-�X��izڱ]��V@�)��v�b3����N��x�j_O�.�������|ڍ�}e�rA������Lʕ�3��p�a���S��g��z~�r$Ϊ����0K��
#/���JT����yH�xF*��?�ǔJ�����˔�٣�$dኪR�-%y��ݿE������Y��˷L�g���:V������lY����#ъ����ci�T�H��u������s��c;�V�I�	�я%���m�t��pr�����/�����N:�a��Q�sxy�0*�ڢR35���g7��^��Y��U��j.�m�����(�b�{S�O�[���d&�&��'��&^g��\]Y|���S��L�=����s��|��y1bɶֹ�\S�����''�ou�$h��]�.˸����t�k��}=����
���M����뢽����Ϩ��1p^����U�ۖBx�G`�D�\��Q��ɫyAHV�Z'/ˢ�e�פ۩J��V��\g�	���~�H�@���v�Dw!�d�"��G�i�&���Ⱐ}
�>/,g�~j�C4M�=[H�W��E(���?�:g�{���^�>�z#����zlx�ݹd>��t��R��q�7^H�����k��~G�NQ��T�HѤ��9X$!�8���N��� g`��Upu�ȑ��i
W�!�q�a�uێBO�mi�����Db�*�8 їǃ&^���(�����S��P	���ϱ��`%�K�6��Z�f��<�^tbN!Vb�Of��X%�}�I������U�p$L���L�)k]ƴ[��'��g�H�1��&�V�_R]V9aMTC���i�|m������^���;G��ݗ�QV�"	�-v�1��At�9ްt@���PB�	ԙ/1u�r�E� �ܴ�~����D�Ui��4��Z�3�|��_�>3�*6��PH�+""����Bx��
j���x:�<֔�Z�V �;}���h͗s�����c�I􍭉�ZVş�D�Mǃ	�c�Z���K�l�����â��=3�Ef�^bL�g*p�A_���
��O4��F[�ȶ`�EG���Z�?T����ߌ3M�oC+:�@���]��/j�;{g�y�;[%&NK��U-��.\����+&��B�`	�K�O�O�Z��+.G\�|څ�'
\�����(y��U6�g���˩��4�K����y ձ��ɿt��k4�/��o��rp�S�Qi�ϵ�WRT��"��9@b�	�)Q��z. ��Jb[���DD&��YT�05��,�*^uxғ��#�0_��Z��!G�M7 э1q�2�t��I++?��/
��O� ��3�D㡞���^[L��Ts�]�E��=�}�6��O�`&�k�	���PR��{zW��|���NU@�H��UZo�E+uږ�*�	�
e�`�E��nى����a��A��Y�X�ߎh�q�cJx+"`Dl���5�P�խ��_�6Q�5�9�*i�+�e wܢ>
ㄈ��+)/ &RA.C�K�qJ��8i;�S�l�W-��i[�P��n$�]*G�6v/oDS���M"	ՠA���>��r�:>8��`??��kj���h�>pTin��ڊ񸨓����óg�������Ix��u��̍����Ҏ���Y�x�R���'ݥ�ẁ��fl �d���Z�ՃA'�$/Jҟ��h�f$�`�/D�H]:�U��[Qm��};�t8k�:TncR���	6���h��X0�ɨ���k��^���
��������3Q�Ė%����$ �ϵ�_��Z8U�T����8��G�е��OĄ��^�)��:]M�.���&��{]�~����ӣc.��r� }\%�����CA-�P&@j�g��|��J��|���z?�&d��|>s��|�I>�M~�c)�rd�*�b���жS�:w;�~�m�a�m���;�65;�6��^�
��^�w{��C�V�e�[���� Q�:�@�y�ƍp���pxpH�ڋ�T,��<�`��~�,�����X-���E_^�z>dp�	�~TS���/^�Hۦ2��V�{b�N��;���^�\�C�@P\2�te��Bx�C�L*v |3�J:��0����R�O��<��G�.T �)�P:�i~������T.�s���>d����Ho�8�^��gb!����Ȓ��y�o߅��A�d�~!�a�����{z��TA|�._
7oޤ��\��+U\cd�A~�w�އ����丘��f�tg�%���I ��ǏIt<��߽G�{�}�v~�k����t?<����j�����"����KVټ�4�(��g�.>��@`�ğ8�㓻F��jb�� /����y�Ύ��T�@oO2�\̴��A:�ٌʭ�C~��Mx��q� օTV�~f.����$\�r�\�̠��͌]����g��H��(��֣���Gl�Qu��0u��ZtcW�8w3j�'d@y~��?������H���PEx��(d ;<��"8̼
_�p%�# z&l'�P�{� a���������߻w�t�� f��DtTV]�NJEs���ׯ�O��>ND�z��"F)��ɓ'4y �Ws�p=��2h��&W0����E����������<_�u����N�\�0���<N�3����Z��p}�V�T%c2�k��?���Tei|ߘ�u����
}%
G>}�� ���q�׼ 7��֠�"Ť��� n�KUmb&�MK �?�Jt����[�*�z����_���<���ǔ\���|��޿���^�v��c΄���0�C	Z�r�"D~4{������gy�j�D��Y&#	�ݍ�Kw���U�Ko���%m[�n�T��&�P�t�Tu�Wc�=�bO'��f�p^d���?o!����Z\A�Ġg�|/"�q���]ȠN��H�Mqo	Q��os_�xAAXX�nD�0"�}ޓj���K����%�>�\������_~����_a�y�9��1��ϟ�>�/]�d�8\�d�\��zԏk1���DǩɆ�w4�����!���7���Vu�#h��Z���a�j�/�-^�~�>�U�:>|Dt���!1]�v��	��a
��T���+�a xE:$�lhL5��P����;"���m��畊,�XR^C�7˓T���Ҿ�}b�zM���I|� �w4 K�5���؄+.D���\2Zk�`n �_�5�: V�@,�eD�s�=B���F4p��tP��/(�{J�"���5�t�Y��q��V8<<�F�}�;���_~!.���؎k���h�^����S��ܽn߾MtsX����~M�\�����Z��6o�8�{
����,t�cH�Y,L�Cq�B�j�][֧+���
�n@�y�L�X��k��,�p�U��mЕ>{�T�vn޺�}u���G	hsj��Y�z��%-��2�N���*�yAӢ�ҭ��D�rS�/
H�=�%�NCU�ٛ<�<��:����`��@ \����%pwy�O2�%���oџX�MR?5���~h���J���+�y&"��W._! Ұ�N,� 7��!X
������N��
���}�V3�B$S�< ,�^'��_�sA� )��m%r���^��d �J��@1�ײ�?�Zb�'�|��5�MI$�T_��*��i_�;��-Ĥ�sab���G���o�y~����?�b��I�;s���f>�=iM��KX`5d\ã��t�m��Y6śFRK� ��nJ�c}��L#Б6���;�L�1�͘IY�ÛL�/�"_�v%���K����L�٦���W�3W����l0(�g 
��,�迿�!���j�i�2	�xD~�K�����IbjTev���/�[��y�z�?�3���l��;�3�<_$�$����e��r�z��'���!��|������&�������#epM��h�CW�U`�s��e�O������;$�R�C?�-f1`�&�,o߾	<����a"�p�Ѓ�#iE�S�����Qg�<)�dB1>]�+���^t/���T���Gp�X��5���ac#�Y>��sߡ����$.���3�~}�^�z�*����L����>�ܹK y�/���@�����?���+����l/�*g�j�y�7�bq�F������G�@[m8��� C1?�ă��B:�{��S�1�Hs�LCqMd#p>R���~�4�a3-�̏Y���^!K	 X�}JX�H�3't�9�� A�翳)/�)�L'���>�P��IK�ӝz���������fJ]d�~<�&I�-r�#��.��_)n���;cHCWJ������U�J���ɍm�L)3� >>��M�b߽�|ٽi/�.b���� �:�a�?�{Z?�j�z?T��O�H��jN��o�������$#��8�|� "yAXЊ�&<����}7�� �}��ع>�b�G� @ �k�3������I	o>�'$�-����-����	~�ӿu��(�NX`�ڿ���t���)��Wl0x��I#>7�����߶8T_͋�
���	M<"G��U<�A��(h*�m#G���$����c�C�=����sV��Aq0���C23��V��!�d�@�ǔ� [�FB�Z%���$@�Q8ݥ���:8�Բ[p�[T���rN� ��}��r�X��HtCEFѶ���ԉf��{��ۉlG��!��I��. ƍ�y�h;�: (��F�$�G�8!�b ɂm��N�@�}��ӷ�\FX&��,���)o!�������y�n�W�.*�M����AU��)�-�)���A3��O��фO��\�[����A����'��A~���T�����2��B��ɋp��
�V�Ebiv[I���c�͒��� :���3���Yl� Q`�}����B% ��ɓ��ehoܸN\(�8jLU.ĩ�*�x��ex���j�?���U}3��h�M�$�АX����^�I�m����J��G�|Q�ߦ#�E@U�:Ъ�eC��h����@۰������3��G�,����M��fW?1��3�Ry�T�X̡�j�`� �tט��[��Q�>k��0a�@V���������ﬕ$����x�����U���j-�P�I^�4l%��b�EW	�����D���@�D^r�tX.l�P�Jr��u�C2�l5`��$Kgo(���	]*|�<6���I�]"��x0w̺�VR�a��Gs�3����}>И���֘R/^�?�t��q�[�n��_}���2C�}EՁW�E���	1����W�R@�� Tp礯������⨙V�6��icnO>��N�X!�IM2o�0�Ӣ�Ԁ`F��?K47��$�h� ��_d:&���`��A��˗.S�'G���YR���_IZ#ϑ,eMg��X��g�&� ��n��|>?T����ѿ�� SpZS	�$����>�9p�'DnU�J�����?�s-2��I�7�4�b<�Ħ%w�X�Y����_&\@�����`t��I�K	$��������W��#��kWIQO��D��*���]2Q���`IG �S�o������ŋ��x�W	"�c�_��͛�X����f�cDN�֘��q�G��u�ac����W�P�����VI�=��;��J�:iu����*�x"���	T��oM����r�1S]�.^�Hn�� �~E�	�=�CsMt�<�yo���	Cm��|���|).�C���| ��--h�(8eo7�#_��Ԙ2=�"�k틚���#��"�Z=��+�jS8�*�_XLO��V�׫�-�2�t�T�X쑸 �C�pP��0�@QEY8���J8_n�%�bפ4&�h�����?�"��X�[
gј[���gU#b .+=\T�s>&b��?�B�?L�|���!\vZ��(�A��I
���ϘxSϟ=���5�ql�cd����8�J��s�y5�I'\g���?Q,��&�y6�
�,e�<�h:7�^�s��s||��Q��<�S$"�
�ɠ94���� !��ܥ��(-��H-yu�J ��TՕ�[�q��6�lvj}�S�7ש!J�����ޖ�5�˪�D�o�.+z
�f�$+y`NS���ZNE�ٶ��L�%�&���=|D k��C��_���޾��*0weLl�p����x���q. N���q����G�����}���'h�;8�j"�3Y|�O�����&������ha/S��d�p�]_�7WC�/
CRl(�0�/���%Y5�p,��T�>+>K�|[M79ɏ�A4���k�|N��.:TNn��b�B��&�~�+���u	��s�Y��]iѮ+�L����P,�
ܩ���|\G;�b�U�_[���ѷ�Yl���y'����F� ���� 0M<@��=������ �R���[���c	��ʄҡ�����y���(�lP�����ݯ���|K�xGǒ�Dߩ�����Z^XR��U��p��?+E�<e?�K����9{�/���L穡�唢å%;�26�v�� ��;�a�9ՑB]��E,���	d3Mr`��I��e7�߸>����D)�,A�fc�)Z�l�}V@5}�nW���o*bG�7"�,���T�yr�(ⷲ��=�C������8<0�6��f*��c���Մ`�0�#4�:C�/�L OP���<���x
�Q��>��D���W���'O��u6�g&j.������8�VBi%e ��p��z��a�HA����~��3���`�~����	O�F�� R?���n'.�ێ���D�?�J�wl2b.ڐKR��*q�/~�D�����C����m��p�����'"uQb�'O(�|�����WwI�C )`��r,O��E�B�5ʎ
'�6����M2����mʚr��"��L�K̰z�d̡�m�'�wɉ�;�(�+�Ke���F(���e�㨅(E��k0G�}d :��i5h��uP �8j2Pe���h&XB�G �' Ap���u�V�m#\�eZ,i2�mc�r֖�-:O���~��O9kD��Ȅ�{�=�,�#S�f�{%1���?��� D2 ���O��AD􊜋t/,���Ç<5|�~(���_2���u�����k3=f��� ��e����C�7�����a6�,�U��}K�`M�\��������^S�����{ugrǨ�в���{����I�|���[�q0���� *���eՇAW;�,hp�T��J���lU�$s]L��fUG�At��mJ�P��(@:%D-!�� _T%��J
�MY�����\o��HE9[�����\z�t��6&e�!�=}����+|
�y%w.	�����?A3`u.M���2����c^<�.�ER��/u���9U.������pO���/X����B���p�WH7z)\�z���@�a�(�)�}-])�	d��~*���f�8Tm�=w*�6�2�6�-I���E�����B�ĭ]��?b1��j�E���ͺ-ٮ� �z�  W�n�4����2��Jy �z}���;���8�1�SE��O_������f��Di�:��)bKt��O]`ba�G�R�y���P����^��O)�_b���U��Yp#P`���ỷ^� *�&~��S�G�J����U�V=�&?7ݽ��V�~�ꍽU �h�'b$@��ר?�\ɋ+\���`�k���n	u�4h_\��Mk��Zi�<&zR�Nr��٢�����GM9�J�P.-�5��{�pw�(J��$��8	H`�J*J[�B��T��{������8SuM�Q����󂸞��zO����	/]S���ϣ%�U'�\,e����[�|?~B�>��_}F�����Im�d%��$�ل�ƨ'�Z�.�s�HZ4�+�A� FJӖ9U��Y��q?�wd�� w��*
�}Q5@� ��y�P��eo�ri���^����2�A?Z��
�,P	8�����m�Qۀ�Gu�RN�}��3Ƃ���f�\�H9���M	υN�H��b�e�IA����#�k]@Ճm�.�6$)�G��e@u��Dyo�ID�g_Α��D �bi.7VA�ďNqI+��A�R�,궤uċ.�s>
 K�iߩϧD%�����K,=��9X�5'��}Ho,���G�4E����."�!�g$����Tj����V����=Қ�yA�0`��k�χ�)"Z��l�H%(5�U�>�W���~��|�·n�����RA�ЉB�  ���N�-PB��r�Gj�7���?�L��:
��0�a��4�~%�a���g�����-�O��H���q��m�٫o:Ozc��8��@eB$)��J�=h�������9�:�VTF�"��%N�T�d�~�S3����m¸��w� =��V$�hQ���΋���D�)������Z%�'~%OpҤLI��{[��k�r��$��5����t�<N�V��P9ߏ��+F���u��_��$�`�g4F-ł�L�^�R�7mf���:I���@I�ˠ���)�������� ��W.!���T��T�R ��
����o�o���R�a�=z�J���G)�+�����0����T�<^剢b&r �W_��	���\�����%D��%�0���8v�c��~��a����.�Vq�P)S�M^��cB���ف��˜��a?jɣ*ю�AW�"�4AϚ��И#�?��GK��R^ P�:)�s��kpj�R�y��t�����t��[EE{��r���&����6g�������UZt�Q!Jl����K)9��gX������Hp#b֟s�Z�@���� h�38�7���)% y$�J�b$��}����"��<����wT3����?�~��{��T�p��W�M	��>$�0M��u��ăWqx�˭dQτ(�����-A��Y�w��i&�u���$�-8����I$��>�F+A#��M�O�Z�����k1�k�^�~�C�odp�z
����Ph����ܧ�t�4��ᓭ	R��U.)�~��5����<7m�>�K4W$cWKp��La[����q��\�[D���(�a�/lL4Yƅ�c� ���W�������NY�N��4�H�R�uDB谊~�ݷ�Mp��GE��8���Wh\R(I
�mT[�������E�����O�]�ʩ
3�� �9b*c�+&�Y��B�I�s9x \&	&,�$�e��>�-�x�2{����+E�m���b��QM��׵��Z�q�1�ۀ�8�rC+��ds��J�Sw�d�@�5���+2]�>5E+��r���@�VC�Պ.ׂo����$�4�tþ��}^$�?�i(���r��N�^q��ߪ7u��ؗ�V
ߏl�nR��(�뛨�۝�@iNu{�D0�w�㤜��ߵ�m+��=��S���$�(��1�(����a�9��!�<�``G�p� �?}�}���o��e�x�.Y`����0A)�+W_��"d؅L�!G���D�5�aq���m%�~>0U�"�8�U�/��M���Gދ���*��Ze1���zo�9���y���H�ʘEaZڙHV����<�,�2�%�0�� �]l�v�ND~�<[�k�����ʁ��Dܨ�o'5>�c��NW0�w�׵A�}�)��C��ѥ��S����}EYv@d�� �d����>��	D��@��Du���k����D\�"��D�D�ą���W�]���}���0��\����?SF)��p��k\��	)P/��Zo���_��F%1q!g����+;<�q� up� ~$�=��΍�f�+���Vj�INt��&��Y���]�u�$���)��[�b)!ԇ$�PJJ���Y���m�;�X�t�j�0�y��K�� �cb����-��E��C=��[D;s�PMU����
��'d�'�(�ۦR�s��c�x*5"r[���9�/)���D���yX8!j�>�����mJ����	˵��ˇC�t� �� ���L��`�W�5ĈX}2BeМJ�Q��(�B�Ir�gR�D"��op��,��h��)�D������O4/�7��,aKb��&#��4���/葔�P�`l�po>�"�Ph���ϥ�u&���U"��0�a��?��@{�O"��D{�v��c��qց��7Z��~7�^K��8P.ָ��mg����ۢ[��X���>�/�uΒ��j�	1a���=�(��)��Ը�$vqJt^����=% "��;�I_y F�jW0ItB�H�϶%��)������K��Ԉ���(�/T/}
УDذ�Cω}|m6&�p�B@�{I�lW�T��1��ip�s� .^�㔨f���
+�\Z2����/���<�>kSfäJ��?�^�T;�k8�J�2m?{p����t�h?R�}��ʦO�mq�fI�*e�	�HtZ�H�z�(/T��
!�i�d�T��(�˾|������h��%J�+"�Y�V��#�Y�W�q���xX ��787#m��R�=�rʜS��F�������4r�H�j��<�S���H�ʼ�r*���ω�8�,��ZvB�@P��_�J��p,D}��������Jɇ���u�&jb���"�:U��p�Wҥ6��T�8���Je7{��F�S���nc��V��D�X�����ӏ�2��D=���	�������jw�T*<����r�kN��@CK���̽K���uN�!��(��.����:r0Ew���1��~��;�B-����(\�r�is��Q�D�� 4 �v/^���/SkL�o�9j�C��d�w$�E�\G~`	���Z����S��DP�#6nH_���\� ��͋���jRe�z\��'��w{� �Cb5�_�^� �Уb1�7�}��.�(�8������*���BC)�br�_ ���7�~NPX�h�� �1U�X3�R��KT�H2O�gJ
�RДh�A΢�����^9hQo�)}�B�"����]9V�ay�纋!ߩUCG�  ��x.��W�.�+-nTu֛��e�K�(VO�9�E�ZXXq�%��I�Of�o߾�?�Hw�"���3�ׂ8�g�=��z��l%�n��Nh՞͘�}�6��"�	��huH1�7�|R6�ٌ�^������I��suע�������1е@a��}Y�%��%�C�@-�A
6�b��(�d���ϝZT��>w)�����"T���ӵ<_
�C��H�8��Ą�����xu���k��Ƭu�S8*�}�&��rC��ݮ^�Ծ����e�sw�����*�=�_Ǻw���Ƣ�Q]e1h�j�B:�ӹ�8�l��c
յ��\�4;�����RJ��O�"-��'�(�E"���rQ	+������	*� ��8#YPs��$#E�@|��E9�����uQ�P�.�믿���)%:�����ұo(��$���x(t�l��+�Q! �8W�o��`q��	�#��%1��R�q.g61CY\��ҩ{�#��~��2���ۖzÊ�#g&�K�R�Q8T����!���4q�f�ЀlgR�ɬ~BY�iޖ���.��DA��d����	�}rV 1K&q;�轶=j��͍�1+�dW6����I �Pt���T�����%O�P52C.F~��[R.*�r��er%��Z̜��5�������+��1�7���ʤد����Y_ ��ף��%Nެ�����D��ǵv�b��.P�;�K�����tf*v�?wnߥm��Zb��!Yt$�#'jp�y_'o�,�a�9}a�$�V}�ơ�I�P�K�
�M?zRԍ`�a��j�������⾃�S�8#�m��CN�����pbg��md��6E���"R�8�}�t�z���a�@g�Y���Gq�O"U5�&S(���r�
��Ld{���@L_�I�=Uj!7�}�B脩P�V)8E��I>���t|�@E2y�Њ�6���0t�X:?f���R]*���E�_�@�=i�xӨL��%��bj���~x�0�.;N5G���).R�+��RJ'wjo�2h(\G/��(J�\P��ɩ�x6�T?,:K�ń��n3:�ǃ���r�h��I2��1-�3W �C�ir-�r�
�T	��ƞhE	P;�`�F����<�9�ⶲ'�ۆ#(��� g�-%K����PC�R�/)�0�ri���X�p|�o��� ��w�Wtj�U҄�R*9�^p�CM�5 ��@&��W����m¡����$�Y�LJ7A��h�6�V
:쪪�Ez��E;A����� ;��\�ٯ\��̅h{����%Q�vn�<��|Ga���|�>g�~㕊���A�5F~K�:.����?��[��	5�X��B�/Ǔ3�8���ىN�Nլ��8qv��Vs�$K}q��'iP�(�î����?+�XO�LbIe5�Db�<�apb��RU#&6նp�@���Z�(�TC�-��r	-/��T��ઞ+J��7��>��*z�>�&�V�T�Ē�@��0.�0�}�/��~��9=�e$����1ZXW��T0:h��$�����?op�mf>J�|����1E�>"��G��b���ytrL�!=$�&����{�:ʡ�-)�s�y!Db����<�y�$��uA�Q�Ч7)��b{M��3;�ǵ��Y����GU(�hAߵ��]�cR�l%�u%t��B��-�ގWZ]m��g%(AB1��S�N�Vj8Q*5�9��2a���jYH'�A���IXo֌+�C@t����5]�����2���E�p�8��v��'�z���4�{��i�����M����e�H␜�E�)�.nB�X��4x��,�,�r�t$���O������U1�j��@]fM,��T��Xh�i/p1ᬛX��6�gT��7;��Z������@��`\,sjC�h8���x����r���S��FVЇF-���T]��":��R��%��w�| �� D�7�x�s"���5c��^�ܰd���=s��"bUn�<�:~���<�X�$�+`�	����t��{'z8�z���c���K4�-%>X9��q�;,Q�A���D�`�L�MU���h���­�����C�G��Z�:��Ad5C "_<{N%�o����W�`��iE�2�]{2�#Y���t815���gTav�mX-U�(�U|�D�SR���
�)���]'��{0I֐�R9�"��k��H˹A,�K��p��VR�� M��u/b(�a>���8��Œ�Kx@���A��bT؊`���7+lb��kD�B��Dʘ����8.�ol�#�"f`��8}u��\x�犱)\QƕV�$E�"p��_o_�~)'��"!�`�>�T?� �Zo�Ҫ���:]�%7���BQ}pˋ��%�5Wf�I��b�3�b����<|� \�t�\
�A2�N�j,X��I�J_K���:�0f���q���������PT3]W"���B�����U�`�[q�B
NG��S�zTNH�2���9.��׉�M�f�e��h'&����L�в���t�HO'L��,��Ju3������=���@�l�I ,!�I��;�O�X�V.:5 v�0V#+zm����+��4�M�`�/V�R���\P�r��j��m��Dy�j�;{z9���"��^��Z�)D��Z����W_ݶv�ќM�	Ҙ~�'z��
"A�>�N�O��?'��˗�eP���$ę�1�1�y�8	E].w%q|"Z���
�CJy�0:��L������c�ӪA]n�$V�Ӣy�#g�'�g�>r�� 8���-��.����� 7�E�N�G��n��1ȭ�u��fǱ&����v$�u�z�E��.h���4��ou��1`�f`f#���$�x�+���]%K�
r�f�I�Ul7G󶔳F�-E�:ӥ|X�+U����P��tq��,��v���R!��7�1S]z6?-�*�P5j?E֪��b���oI*{�����"�L�V���������|��K�\���?�{Vs���,A���N��@ߗ�m*��n*J-)R��Dy���4R$�4�fd~6�]z,�*0M���x��3j��@y�F(�ĝ���T�>��̉D
Gݑ�с���Dm$u�4JF'���LM,N!T���������+'����3�/:U�$R-̦�8���Fǅ*pgqg-��X����IX*��w���ʴ�:��FE�t�薡�&�r��0VT����ǚ�	�� VUq90�@1�w5�:���"90��d�T$��ܙ�Yw��d����:��>\
�Q�w.�h�	�)8Vp�0h���yQ]@�x,��~F@-����aV���W�薽������1V/�D�X������&(�1���v��
uĽ#�
�x�2�{󆲏/]-%��#W�<�2����	�Fj �(�3��S�6k{`@%"_�)�4�q���DY�2��0����px���Bb���}�D0�E��iEV���7|��i���(쇬Wȫ������_�,Ɖ��DNH�o��I�)�k���J��S�jL��C��Q/���M������-�hl&�c���7�����KT�pt����D�Z�K����eࠐ���ܢ �W�^���*eg�
 ��
�`H�s���⅋���(�Vm���-��]�/�(%<E�*x{`����!(C�/��m��^}5���g��Z�{OG�R\���!� �����r�+x�8�Ku�3� D��i&��E�y�)�j�dj�n�N'J:6�dc��)?P��^�krgy���~�;�4l�ʧ )���/�
���%��n�D|�a\j2�@9my�ՋTH&C��>�`� ���}�PO��5��΄3�a!�� ��a���Dn6�V����Q�C"F}��JW7��L7dj'Jԣ�NhWY��T�cE��N�*N=������TLm)���J_t�x���<!�鈀��:�J�E\ʤkM+Uɉ���v�N?�QjŮ8�U������9�������YS]D7����`u�V�J�����u��sr��N�g�@�|H?p�\���m2��9N2p���D 1�	tMHf�lU3��T���gQ�܋J#�z*���x�D���1e�G�^��t\k:劓 ���iJ�5��vBݡ�'s~^<#R�������B���
��^T]��3���G�c =�EYk�@O���%�IA�e�����w�q�⨊�6R[A��{�;W'zS�ƒ,��+4���($,�T�4/����}W=ӣ�̌B�8�Lf�����t<� 		��f��%ȶ��J��&�T{d�?F�0�9ǋ��u��b}&�ڱű?��ױ������%����}������d�x������Pf0{G`�(��.C�A��G�*㐹4ҽqJ>*A���n��d���	�V�`�����	�(�����C�v��G�U�h��?�z �;�)b%�;W8�Z��Ľ��6������N޿dP�����jU.�.R)y���i��9��T����AG��6i��޸�M�X]O�>-��XQ���``�S<�qn*��7o��\ �,%ݧw�a�¡6���!� "�n\�A�!�p���.��·�����3T� ��:���^3���D�4����jl?��P��f��r�>k�R[O�TSs�}Db�#e�Ղ�~����Q��P�9���B���xL%�) Ȝ�;q�	� +џ������~�'qs ��t.��3+Q�ϰ4gf�y��ɦ%�Ŷ���N�h}�^��ƇI��ꝉ�Y-ۻ�o�+����U}�cZ�
`���H��B_.^�j�G����3��~H�}+�ddbF�N�	�Zp����?¯~%5��?q�F��K���M����!���u�Ë�	j��|ɺ��s�`4q��3�(=��S���l�Q.j2U��R\���K�����$�4�q�;b�cc4_��D��Y#"�T����۲$����΀۾��3x�[ݔl-�X璠�5����"��HD���3�NJ6�̫�s.{J���_�I8TY�N!�8$��ҡ���w�۷H��=�C��Z�a�ވj�}�T/��Պ�}������ ?�uo6���?�B�����3I{F���)�������ЗH��2w7τr�^_)ɬ\�Z���de]���o#���0��ء/l-�L�N[q{��:���1q��8���d@��'���Ts&f���A�
��5 ���g�u󖉄���A������O��
c��/G�N\��+-�a��Vl+$�F@u��s�3�]�U�����U7��۸�U��W?��L��A�]�p �s�������p4�����S#ゼ�d��
,AZcΖ+b@�\h�X��fK��޲>�}nSk4�v����a�ߨ�%�FV]?Z)}̺��O���)ZI��"|��4�u�~��>��Y�锤P�>鄮4W�Äo�V�;Ҍ9V� �_~&�< �{���������q&�I&���o�E��G<nZO
��ݿ?�����N�	YT?�> c���wI'��U�NP�VW*��ͭ	τ� aH�*K���TǊ~�\"a�֒.�`�Y�������O�������_�9?���|.'��{��ܔ�0�8�R�͹�vJ�F%o�>7��h���W�I�­�b�IUCEE�)9M/ߥJ�W���&���
�$A�Hb���^�|It��û��6��%��	�!�@]#$��(/ ��]�O�������g M��l��A	�����ȟJ�F.7��Qϥ
���O�������&
��e�=?��)<��bȠ���gfd�a	��MXu��4�|N�Q}בh�� !p��|���H&qY���^<�9���`�d�J��"�i1���@�ʍ�R~+��{�(c?�� � �h]�Ɔ�G�н�en�`Q~Ic���K�.�kD�	D@��o�q/�{Ρ���0���L����-���T�������0�EK�;ƂT'R���ӫ��pxȺ3)_m��(>O��t� �F�4m]k'�PMV<#�Q��d�k���2Q@���k*^+A�o�"�jp�>��0ׯ^���&q�P1A��~x�`WO,���8|qH ���_�9�RMctB6H�MM�Vsj���F��X����<��K�"�]�����D�%�D �x � �J����DR�!94� y��p3�%�,��{b�gC�}���3�u+���4�?��%D����[C�=�<2Xv��Ŀ,��e<Gt�b8��������T�Oݴ@�t�Ŝ~�m$�N�J���/�d K`t}+H}+}/X���@|�� փzVp&�}�]���L\&8x/��X��Zd���*�����ne R�4=Y�1+l��Ɍ�����ǨN8So[��:w[��`0�X�c�Jx�I"��0*H/D"�$�lP�]c���$�<~�<:`�W���Y�Z
4)
�'h��;J��8�p߿#�b=�ܼ��#����"�v�� �X3E?+B�Z�v�L�9���}ōf���X�E�E��1�?~BD�;�3A,s_�A��D�K�1_�8�`���b��{eq�����  d���A%NP���ݯXG�Ŝ��  �1a�#�z�d�ӟ��~u�V2op$]��b��� n/�� 0��������	�}������P���5�Xd~����:QZ�Q$#^�3������������Z!�k�`���P�,�-W�]�7�9�_��1��Gp�cb��6�"ƕ�a�ſ4��I��]�=�X�(y4K-32��c
l9��� ��0������;w)��8�,����cq�ӟ�#��|�[2��[���'�����V/�z��T��[�]���jrNhјxM��Ǉw�6FUٌ�bT�9<�[px�TS��T�LA\�^���#���Q9�Fyb���2����_�
`y,�s�;��2� O�2�{�����[�'�<P! �>�cp���|����@-���=��5�4��D|sBqSB���3B��q'd 8�q稥�\[��TJ_���)~�1b^M�H�ء.@ZW.���[�I��%�`M�RAdW�Z2�a���E 
]�0�c�!Xq�8�ܴ�T�eM�Eq!�8m�r}1���7Q�)[�S%��~5$���i(Z��N�;�շN���,p��NA�; '	���3�����W����X����b�5��Ot�D�?�J��/JT=����S���(OF�yyw�~3��+hIxbnSd���P\��$Nz��M�'�+B����Շ����'R����J�VR�ㅼ���)|�.KI�9����V�_�!�f�)�a�{a�s�6)tO��#h��譄�B�@M\c�-`�3�QT��O���q���I_q)��Cu�:(�o������\L����ܦT�"_o��*s��NR4P|W=%�n%�����S �;��� %��й�<�mx+@���T�HD?u:or��_��NݕF���I�
�)E�-?bq�bn���V�V(ã>��Dq���h�%�����J��\+�K�td�w�y��L ��v�����/�鳧��Y���!�tG��䜒�Y�7���)/�����2��\��Y�/�MZ-`�l�Z
:DX"1�A��nߺ���Lhz�p` 'r��ۏ)V�D�qa�8������:��^$q[6 :D�����{rB�D��� I\`����lA�^+�ҋ'���'����WA�G�c��I�!Vc�8q?�`��vp�j`ڧlAd�SR��>���J�pe��"�>���'.��m$ �����{����%����
|��i��
ԍ"����L�����}�s����Rӈ��K"�P�w�K*�WjO��mHpI¡6��|Fa�"]g^��aR�<id��{�zh�.�Z-	
��W�FU�F����Ę/��Xh�L�a��~C�j�l�����K�cK퇻��:V�x���c0B!&�T}e�ۧ��*��\Vz��SB��/I�F*�!��M-�:X�R\�����U�i�@��\R�U �
�%�I˓d)�����?�՛Z,9 �S�Mh�87Rl�8U	p�_JZ���	���9rI�%l
xoF|00���F�,q ��Cc����صʪ.TM�H2����97��J�XX:IC��Qj�}�#x�1jo{ٖ����0�S<�Hs��&EQ��X���To�fҹ���dqo�;b��B�����_�xBRc��B��o�rN�w0��n��� �42����o8{���+��E�S���0��6Ki&�A<X-?yL�������r]�8��=�D7GJ�N&8�tM��Du��9a��/�C�D�/�gb�R� �|�	e���"���S�|�B�:��Z����R�&��*Rb&�j�3��j�1 sJh"!�b����alR�b���\�z��"��\ ��g�Rғ��Z;�~�~Sq��{c2�0&!��+>�N�A:kxQL�`�3���?uL�y):�3N��0�|ڒʈ�ԺQI��ʤ�K� �D+� ����C-�)����_��
���oo�0�KjK� I䊇œ��_� �;�O0	`0�ozFz�%��L
�oaWm{���YjH�׬��>Q�R�P�&����H$Vkl�-|��[��`0�$4'%;>/_<'Q�&��X�|�-qa ���٭�L�~T����U�ZJE�?\�2v"� t�~Š2�1�*�����Mp��u�Y}�~���\����"BG3��oݾE�DAOW����.�g��R%����{G�%�UER��ڼ��~��������~߸۶lI���Y��� 8DV�VѤdϝt�EV�8 ,���.%��>!g��uSx�V��~zc)�s�oq6:F��׬���q�g�x60�BV4W];4�b5Wg0[<g��^�a��&��|'���1�����ߣaɴQ#���j$��f�|��C����xt�R6�A7b��{ɹ?r�ݻ���+$���+�����Y0q��#��3=\��e|�n
�1�r��=��+�Cv�X6�U+�tV���j���Cl*3�I� �մ���z�'�����ʘ�3���ZV�T�Ȯ5�IB5�Yu ,z���X���'�;����_9[`�p)F�������%)���}dt�A�f��3_v��RB�h�����w0��U|,��*� ���F(�sI�u�����[wn'%_Qs�aW)�Yd [Ӿr�P5���H��*��h �}�7.hU���M��
gYi^eh>�j�M?����:Pڿ���2�PQ�����8����%�����J(�32^&w���;|�u"7i���ϛ>ϵP���
�?-{I?�6r�*6R>��=��_w>���0K	c;����*�)z�=�QG$���/�ڂV
͒I's�mFE}���E�.Dp�������ü�
�=��n�am������M��{�����GN;[5�2���B����-���S����0X�vS�I�V�\�f:
�β�+H�cQ��i̍�a1W,p�deϡ[%���+g�S/�x�L�J�����O�j�Z������0��Y��M����Lo�G�� ���t�R�^whs�88<��4�1��_�k��@���tx4��i�Õoz��)��O' 0\8��ДwD���ǳ �i �E�QG��!�A��5�?0��k��+&67*����k��;��$qh��x�Y=g�9x+���n����9>4ݔ���>F��M�n����6�e�9�3*�߁�k�8�fF�Cj�*ʘ#�;Λ er,L�?B�#x����\���/]Lׯ\MW����/_KYih��P�t<,w´SD��/�a�
9���v�1�p�,�Β�cm���㐣����P�y������N��%z�nɅa8Ii��쿇�wZ�N:�i�Z�U˙�~�RL�s�*�N����h�E���>���߯UPU�nY��������/丠-Փ�T�LM���$���g2�5�5{A<�?�Q��BWxL��7�l8Y�Z�N���P�E�u�%DM���ʊ�i���8(��G�}f�%��sR�x+��X{F�b�*(F�j��1O�
ܨ�u�模w��{�x������l����̴e�@w���eg�#皒��R���?}��\�>N���:.[��(g��Y ����Xh��R��g���5�2! �1�z���=[*�8ą��"jB�zX4�����@��"��ϟ�&(�	n��F�h�2%�����-à�-u�/Y��R�׬x�H-�a��i�e�x����Oq����yY-m��^\pRY�"{Y-=�7���Z��<�#4r ܚ�=�"����c�Pɯ�(Q�2��g�8��#R������V>�6%��R,�i�����2�I�M�R��RcJ�r^mbi�dO~o�R�ǰI�&���uu��$H�q��������-:�����fpQX��y�Vb?AM���sq��Y��Fl�=%�^J�:2J���'H`a��IJ�'���5�aӮ��čB��<K�ǉT��	��x��	�P��ug|0�� ��F����wn��-�Q�%������������Z(�؀����J�}�␠���>�� TA��#�0}�����-�M����Qw����/�m3�X�;7<��|cwe�t����Z�F٢�2e"ĶiצsS��N��i[��ʎ?vx)��f
���G�l
��x�#�	�3
�{d�c���g+[��-dl/7�~������^�MG�7�U�;����z�X������gJ�Io@'d��ci�^9��n:��6s����cx�NA-K�k����Ɔj`f���h�G�+)�H�U�U���˗U�J/��r��& �]�"�YbU*,�����8�7}5�?쀣�%�5g�c0��B�������f���)oǘ�g�Q��Ń�W�$i*�9	-dF4��0M��+�A%�	�wz�����*U�sJ�S���搚9�f��{��1�`:� L�ǔw�@5�ʸj��fsvJ�r�®���!T�3��۴	!th�:R�ws�-���N.n���b�@�.Wi<�
J��fc�i���C�P�q�ڍt��5	��ֹk�T�4!C�{�z��+E0�a�7o��y�Ze_�3�������<ix�Dll�Iǘ�ĈN@���MY��l�BH$?�IIR1m�@��G�M�^<%�F�Q��2�r�zX �	|���M�eҼ�]����j8�T0lM�m:m��>dW�e>/lA�#��M�Ks(��i:������؁�!) ����Q�9���F8g��C#^f���Z)➇ٞfޥ��Bl$��������5�?��?�ݻ�$��t6�������.�K��D
�?���<~,d8Hxx虊�H�X�����F��`��v�$~5���>p���n�-�����"P��D�D����q�t����)��������2O�q�i�� sRja>�u"������S+��	n�o��N���w��D� ��5g&Ou���q��z�'-�WMK�2H�G�����m��
I���/��/��N���y�2h΢觠#��,�,sy,��ת��˔�n����?+#�.�ijh�T@�zE9pE3U�#��)�\	�q��RA��B��@�B[ݱJ��O9�����MB��(�����Y��vQR�KV�t*�}�$� I�R��3[���<��-�y�A/�C׼�(
_�#���K�(�TC3����)��c���rjp�"�U�
G+�$Yk��B�����~+�������sp�B��!Z���2I-����#[Li68#��M��Z6	��[����Ѧ<p�����[K�H굇��M�7')��h�� �<4�)]b�j1��=+ H�������ο�����g}�m�;��V�c�B�	S�u\�ٵ��j�� ��B��*(4=�Q�)��]k��l�0�7	�s�T�<A���7K6#�	���'O�� ,@��޸Nq>���VS_�.Ꝗ�~�>l#�Eg�$��+3K��!<y�&������F�ϖ\h]�������a8⚈	 ��T������2��0	rp+!�I�����i�m���5�k�����G�
9��+���0YU���+Z�zy(�R���%P��Z�6jETٰg�͝R]���G����ݟTVd�[%Mɲ�"�S�$�3�&�Q=�	��UԢi�FC6D|p�N�2������Ҁ���?�xc/x$!-G�I"q|�(�w��myo�M�}�i.�kK4)�G��dcY@�%��A�-+ьg9cb�zK�{Jۄ��;2G���M���X.��_[�w��S!�r���_���j�9y�
��P%�H�gn1���.em�q��W_K���'τn��۱��]%g��7d<���:,'���}�k�0*@�������(P���ݫQk�k��KP�~N|F�Ӛ�8i�㌛[�ڱ��
�$�`�.�QR��G��ɽ�t����4�\��(_�&Ę�.d+��L�_`�Õ�QC;}Z�(�ZPl�L^����U���o�I���R΅D)������_�@$�f��H^Ѵ��	)|���̞U�f�CŴ�iO����}����[�'�������{�;�fI̪+��xz)�Gpȸ��L�.:�4Fl�����j�R~_I�0�ף���L~�u�
ԯD�.��r���g�8h�X�FQ��/�G�M`r�u���]�v]1�2���z��
�3��p��ɓ�I�'�7��&4�4TmD�g�z ���Q�@Ǭ%�gVMс�`�g/�[�փ�𚉖�o3~��~�2nr	�����lae���1�II!;�c��8��,���&l����]MPʻle�w-�d�"R��*Ʃ��\,���Ke��&|q��Χ����R�	��Q4��pU�=�>���H�i��}��Lˑ�s7�̬� ��P �F�6����p':P۽�Vx�tF�����)J�!�[�Cn$'!++�5����-���m���):��)��O�0+�>� ��`i���~#5���@jp�v?\����%�/��*X��ѝ:�ׯ]���}�>��@�Ii#4H@9q%�?%�I���~������y�UC}o�$nײ)�����s���P)l��9O7%����&�z�<=ML�j����<���M��M��K��!�WE?�X��It�m�;/�{�MRzKSXP
Ǚ�9�~!�{������g�vH�j?f�3�e��;��4�z ЊY!���=���Xn�� ԌGL����i���Nb�`�G�^�_W�����d�c��8�XZ�pc,3��]lr� d4�H�Ki=�s#Qa�8	�����G0Q��r�Cˀ��B�'n��ɿ��m�FKheT�S���K��a�t�n�U�p��M0㑉�zh��@�	�+ -��@�Ar�B%.0�Y ����]�|�wp,����KWd��$C�Fc�b	*:3��k��T��!��:��OJ�g�Y�`���g�O����9����O�}�	�p	#A��m�M!{��^�Y꭫�Y��Ġ�״Cm�z�?\T���bĕZd���$�j�9���@N3SD[�U�0�p��L<2�w��:�ciB;>_J2[(�(8	=x(%~���	\Lrh�0�P$�)0+)�b�>��!%�M�Xh9���p2��;ڦP�0���*P�K��A�炀Ƌ�k��c0bk�pB�g�>�z���1�_>���W:\�&�G�$��fO�:��pn����F�|��WŁ�7"،��� \Q��ʪX�X���7��J�H׮^������:,m^�.\�|XS0���s~�XY,2���"Gf��R�iD��s�����L&X����`Z�n��g��&Z
[�-v���q��h"Ɗkn�K���W�?�1� E9FY�Hj8���N�Ѵ'j�q�nm_�<b�8�V	�!%�W�'U� �2�'�=��P�yӆq����B�)5S��E\߮�Ok���o�J���?E�"#
�
5�K.Zg)Zd�,��f������Ŗ�)����i�\�r4G�hCGK��j��~f��c�k����ګ.�?������ڦ���,8b�tnъ��VJ?�tW�Ik�鹘��s�źcm+Nr�U� ��~	����K���`QLh��{������6�M@׉>kfZ�����SO'3g����q�m>o2��㹆*��7�g�p�mX�{~��0?���F�X.���^/�p�V-�,�ì=�5٨-Z"�Ԍ�0��@E�Lt8 X._ޗ�;��(p��;E(��<��W�D;�B�h���IB� L�;kC£����ߊ'f��@��BJ�=m����0�#b׫a��2hy���(�L��ʰ�x�h����!PǕs��v��H�y�n�5�a���bS!�?*�r��N�oq��lo�x�ŦNO'$]�{�A�Gxu1~�?͚�P�*��eK�s0�A��]��a���7c,0�p,��8884%jaT}:wD0�
��>E�ߔ�����"�/^�:R�Y��>��M��ٔ��Qu��B��?�5z�Q h�KR���V�O��gr��`�A��]'l^A20$	�Gk�3�����Q�*�I�>i�X�x-�#��{�@RB�%�_Y�o����tD'�i1���H)}�~��*�)�X�0y���;��v������l�3Yd���`״I�C!�u�޹9�Tƕ��]��Ls��ll�;����±f�s��TE�s^�B���e����v�.�+:}'�G)������2�Q
�mx�`ަ�K*砖���ٯ�`:w���G�� @�"u�6u$��whP�6�g����Q�3u�
Q8��܏:UדV��1��΋����Tn����f�3��-��y׍i_�y�-3���üs�Jw�x����26��Tɴ���-ޚ�d����	��N�b�0؎w E]n�:�"nJ�K�哛���D�ZQ��ǿ���yIqO�>�m':�p�������>x��<y"�?��,�?K���B��p�]+�&aO��Mj�d�j�4ŵ$���Ę�D60P�C_OM ��el�T
Osč�pĒ~��S�;��%��A	�!��k���P��O�Ov���`��C[��+��s���,js��/�l|��%`�h��!�Wu�~f�$4+�������h�0/����(P�86�A���Y1H�j��w>��L5�|�]�z3�Ï�&� 8Ҳ�D ���U�:C)�y	:'��"���-.��4��s��)��[��:�(P/J)�]��vqI�{���=#�V!ي�y\j0O�MW5�G����bE�K.�+�l(%]'#��K�S�ٲ��"�ӏ?���	
MA���{@�a�7_�nߺ-Z�6�cc(��,����V�<�cmʘ����%<[�er��9�~�CK7�+��\ʹ�U�6�%5�S�㦉ϳ���X�t����P�㜃PaC���_[걯�:�ÿ�MZ)�BXb�'�P�?�8u3���9ax�`��MR
O�0ƸA@jl7B���.5^B^�e6w�VF�0����G�M��Cg��~�1��cZar�h9%LX��M�,�%��Uc�_u���_M9m��"t�x�
�\R3���>�`w�\�i������v}�[� �ϒ�ࡘ`(��ة��/��9w�3̙[��Ջ�|������$4E����D3ŏP�	�E�Ф����0��KMW�dh.�x��f�<� @��j���4dj��"�,f{}4�)5|h��I�
�Yg���H�@t���18�'l���~�-��@�]cN͜���y��h�k�{{��ˌ������}`e�A�[�N��@�H"h��&��P6\\]�G6��ӯ�~����k,1�G�s����g�d�*ԑ��?�QM�����0Eh�i���t.4�_���tW������{�fr�����+H=R�U��5�df!oM\�O��5�'z�Lg�����oH <���QwTh���$��۵2�1�<��0�f.7�d�$�ڠ�C��j����&&��.^��+��l5w�����4B�`!@��A�~�}��=%��ZC`V�19'�K2(�6Dj3��Ա��S������Ov�W��`l����\�����<��˞V��4p�'�PF�g��fs���~,|�HsrB���,�`?���ƼA�n	���#�fjZY��h�$����}]l���X��r\�@�c`�`sݳJ�d��=4��gq�Bb�޸~��~U�%�b�x8����gqd�
���;w��cOxs�)�q4�q���Y75j�n�R�� �P�p_����)�B#��>��?f�8�k�H�gv,j���Y�s��{��Z�b�?���H�����)�^��.rgT5�_�	�����)��!��ф�C��Z�__��u�
SU�NX4��������W[f��W��3�97'd1�G̈�j�^&�8\VM� �|�.΋�/�%�~r��2Ύ����;&�:,	��b���d��a��Ӑ�К괿�N�t\�Թ� �l���p�j޽e赥���J���:� `��` >cq�#)e�^�Ï8�����+���#e����?�J	�C�/ugw!a{3ې1���bӼz�����6�l���\_����æ�9J��i)�P5���u֧U��=Y��UQb!���Ԗ_�q�E͘�^���{�{��5�N=�X�Y��ʸW,�em����]ٿ���L��4�<�
�#�H�{F�=ާgϟWa�D����3��Ki��7��, z��zk��O�>�f�C�`���ʑ�����!������
d�'�VFlb���ciy߸�0�l+uvH���0�U�&3�G_"����.&?��&�d��y�M�Ñ�%ơ=�M��ʐ�|�&��u�m��d�EPt�i���8��8��M�U��l�"r%�n�����k�G��{���טgBJt��GÝ���&kۈi�{/>�b��S�[��!h��_<7V�ך@b0Zm�UHh8G,��6P%J��~�Yg*P����b�`~�:h)r��Z� ��s0�$&'���311F�
+���\VV"8�"�Lv��;!���&����L�	Zu���1P�^<V�e>����uǼ��g"�`�H��W� L�g�����`U��['���(�1z��dNd�'N�U��V��G�ՋWR�g�8_�h6�P�
��
S�.�r��`�/�?�l���=Gk*f~�&��;w��ݬ��H��h������GKR�Y�s��Lܚ�L<sR�Y����{���>|eq��0�/]�)z�,��^}���s�K?�ZB�9�7j��;�B=i$iIbcK��;7��̏�S���ͺ4�}�C~|BԆ7�]�������m�0�2�:_ذ�Sv��j-\���F̜�X��V١��q��{H�:�,�ml��a-@5�Z����H�.��z&���woe����z�M��`6߂B<&X�2�?�`��z��(����N�ח�6 �.�U�HL�&��� �l1,4h~0&!xP���	)Z���UbEp,�uGf��]��]=O�3\�5���s�Q�N׮_K������￯�Ӂh�R޸NV@���]���b7]�T5�K��e^N�z���dY�%"Ӄ_���ߗ�Q���;�L��C�`�~V�	�c�`G�AdA��5��� ~�*�͠%B�ޫf>��nߺ����z$��Hj���n���E�H�r�Zk�3etF���oG2�TCD�6pց�zy�5��Y � ����Bɶ��X.EP���o�ԫ��o�/x�nf_|�U5��9Ɯsɕ)I��z���hu5�|'��9qf�X���|�����7��3��	��>
4QS�y�gY��t Yt�*ԮݸZ��-I�x+!yi̮!ʼ�:�l�����`�-ϾX�1e�|V�zb����.��]q<=��?�0� x��V��RB��@(}Avє�Aփ��I���[�nF�Ow|�T�pB�S�i���}�d����]1eׄ��X���r�؄6Y�A�OZ{rg������Q0c� <�Y�<�o޽�Ҹ��D`���䙤v޹}'ݹ{G�|�_B8b��N,]�$8���˃RC�D��>�x��^��n߹%B�Β=b������+�;����#�0�!� d���>cB�dӲ�[Y6��C����y3��� 4�s!�Z%	�E���?�����.w�M�\�0tq����0�|�gYhR��PY�`�"�k���+���a�5ee����Kt8�כ��Mן~y��? /�Q(Mk4�{aJ+�8g�3OW���q^J?~��W2�Dq��G�il\�3�j��Ν;:�H��%��T��)�*a�0-]-F�XKu=$%>�p=�H�mIy��5�1�=u���)��z�'"�&^Xl �'D3��v0�[m�B�lp���E���xA��oAb�ih���\A ����b>�v"���I.&0ǥ�������|�B�W�Tv�-���%���e��eK%�� ��UP��Y&pX���,�^C��=�Ak�E���:L{�}�
���U�W�A�)8����XL~��`�V�W�"���[|������Ǝ>$�
���"9bh�FY\�X�r���qh!B'ǟ�x�?3C�����dEZJf!lb�q@ bIrG�����j�����@�{����y�g���]��0.�U$⤮�K9������3q�NTn�����G�9��3�����M�ib���r��j�����$�+K�-�c�Dsڤ�d�ɍ�X��^�~��
�גƉ���A�"c�ƅ��(f�M�U�@��Ź�$���������O��k��c� ����~������Cqj7=�����b�"���]3�c�Z
��Q�GHk�o^�y-׃��{sY ��|��	95��PA����������/h�O��8� p��n�N�}����4X⊍s`��"����x�Դ�d����Қ��"�7ٟ�ҟؤ�uW�{d*�>Zj����GI#.�s!D�8GEt:�!� �N��\��t�����!u��l�W�W9���?�@����n�)$'���V{o� zG��h��Ip����eؐ�K[l�+WA���%=��az\M�w��o8L8��zY�E����y%��+����E��[������7��;����?D# D�WZI/��IrAV*h�0���8�ќc�$Rb�Y��J�F=��Z	�ܱ0p���&�I1���D�����|��1 ��p����qcZJy�#u�9ś`��}�o\Ow놂�ܓ�\dy_�������3��&��ZHU�X��'[�/Oj�ʹ}v
�ln,
3�~�^����L�͎7�D�ږ D=�DA�yr-NC
=	�$}�x;��0
�i��,�2��V�'w�e6�3>>�@uAy�ˎs�I�F�i�v��E��kY�'B�����s6(|ɒ%��2u��/�ᚈ �=4�*T��y�N���Y]�Y-&MQV{`�z����5�;9�Q��?��?��><+�gox�����d����V;}%��UH.Ŭ��й8�>�\iv� B�L?y�Q1k+,zPR�I��`6XM�Ɖ	m,ڍ��Ç*�DM�  @�����kt�w��M_~񥰷C��!����5���o�����k1�S�z*a�9��Lk<m8��=��J���p��]R�T¨Bi�(�M�.X��/-�1�1�����(a���lU9���x�!�ֳ�pd�����F��8-��i4Ԭq��O�)l��05��&��(P��S`��&�����5�m���X�衱�C�I&�k{`Z߸v#��_ߋ)�4Th�B��z; �w��L@l/_�pHB&᪚�R���ś7�7�~#���
�m�vBAB_@�W�!�,1���0�!� �!pᜒ8NI�\y����0��|E[�z�YcM���^� }	��u3�^ūo�7 �[����sq��7*�r3ea�R���-&���u�	�����:����ֶ�t�M�h�V��xl�V���E5�1���in�jՊ�)s?)�|`�l���>_"�;��h>�X�������j6���0��j��i���
��{�_.lj�c3vZ&���߽�
���i��N0&W艹f^�;&N՟���W�RGf	;	7U`}!���Ѕ�A�pX��G�2�`2-y]*i��52�eެ��� �}��i��VE��ƥ�_�!y0��K1�/]�SzoG��W��shaVKK?ݱ4�,���LP-ĉ��]q04Sx��6���9�9 ����17ě�1����ژ�L�2��ʰ@��p��X��1*�&��U-uF4�q������Ι8��=Ne�����F	���aR��J�D�q�Z�|Y��O
/
.
�lغ?WM;f6N��<�ب��l��s�!�5����2+r�-C߳
�S���П9>�S*�������=]�_��[-�����~7�x�i:��c@C��ʌ	j�Bh�/�x���~�(�ǟ&�ޏ�1ߓ<�V��,�"�l3
�ݻ{OIF,f�0� �/��)�V�vBcE,b�s@1Ghtv-����D�gi�AԿ���g3�Z�>� S[��>'��.>���G*"���
H0�Z�@t�l��pH�E���}.x)��X6��^�K-�(�Hh$�bT�T5��ZY�a>����ƹ����s����q&����"��'*p�Iǐ���H��(��2�r�=�\*4@�H�|$1��L`���������+��]���0J�fˮ���:�>(#�*y�e,��Z�=��m&�WJ��NC��=ۛt�/���l��wr��b��̴Q�]�|Qr�>C��+��I�X���͛��)j��C3�W�(����X�'���Ȭ��\ 6{�\Ⴐ"�:�)g�2�q�ʃQ�����z�����X��:蚩>rg�\����S�%_�6����0*@`��;��i���B�Ҝ�Z2�_�� �.U�����$MS]߯}������':�����:�m�N,��g0�KgD�}���f}jk���)���:�~��$׎�
P۬�a�]c�z�w�4�by�hm�;���N�~�:i2�8�(�rZ����:QX3�u�Z,�� ���M^�61ΰS�d(�����k�fx@�b�\`�����,�N@kՌ��A�4��'�J�j���p-J Y��*�3i^q�:>mݕ]d�"�F��X�
'���0����hP1��jƇ��?Z����N�"�m\�D����8�~;:�eMi��f�fFm�lme?u
C���$���V���"��M�M�I�W�27�VR�41OAE��m͊]�Vݹ;���`Bx��a�	PMi������w�8M���Ͳf��Q���Zdw�$TsnZjbg6�+.~�V���'2 ��P��2x��CR��"HYK��Aj1)����Q�,D��b�?�|�J�W�+�)����,������;���#�y�@��$�$�Soּ��0"`
/�<(��(��ʲ_f!dep�#��24[�:�,��"�-���`��Q�hԁ�UPc0Lve�nE����n���� � ޵n]�!��CU�pF��W������IT�6�-�M��i�y�"d��_L�侊��u��&iO���t��5��N�Lp^ͨ����?#F��*iNNFT�'� %��ʨgu�]	�J#SU�)<��-�$-���N��A��Z���*V���.n�����t����8$�a��h(�v;�,څ���k�I��$eP�ՑYnbΈY�4)j�Z�~��9��z�	%vg��7��L$Nŀ�<1Yv�V�,7L���LۭM�#�S?'�DP��a�ʘ�Zx����k>���~@}3�>-�G�z՗�f)�S=�����5<l`��(���}�w���IװƱ��2����i;aɟM�y�N��8��g85*-L�RZ�/[o3ü��H��'��b�U�Q�A�i^L0.,�~4\4^3�K���  S�k+S���{m��v��L!�g�&�3j����t�ٖ@�R��h����D�����ꔝ(�y�m}R#Ӆ�va�NS/�����z�wơ��=#�2?qB{G�K�y�ڔ�(��
6�*�X\�!e�`6׀
!h�M��q��^����_ � �f�����6�-wPLfr0�p�Z
�?%Ιql��F�O����o�P�Q�{h�c�&��&`�s͕�T4a�]��z0�O�3�s����w֮a*&�-�L��1���y�:ޅkf5j0b��e���_�­/���{&�4%��E�&P��J�{t��1O���2��=���^:��`��?��V�'�Pه[M��Bj��nM�� $��pSϝ���q�Hr�kKa�ۯ����$�H�K#w���-y�"j�]�&ro�f���V��I�e����'r�	�_��p�I�Y6ez~�m���g��X��ht��.Ϝ5�q,��{v���X�h�ك�R�c,rL,YZ�����>���fz�ƾTI�N��.����K�`�D��f51d�ֈnP���X�K5X�i�_�:���E*�Z����������s�';�;Wj����N�(����S:�1�`c�;�6�G�{�F�f�&j��1�⚑�N5���F6�ډ��/�����&�*:$U�Δ'��-��0�8�~Ӧѷ���L
�:ng�WN>b��`UsW��)|0�8]�f=��.�fOꈖJܼ��͖sQ�,cM[���6���K�������w(��1�=���16�=��1�I0����!�1�7xP#�>K�\)�Bu0���x|B�:�NrX�&ͣx�F��Vj�&��v��5g�����;J6Am/�����ő����,��|g�G�m�6JQ�3���R�>Sش�������k����2{>��~/�+��Z\6�M>�Q���Q���U��|b!���~]鼢�q׶|�f� ���ZC2�� �ti�C ���M�vs����{���J	�dC��,7���*������55�lʫ��\o~L!0b��ߦ�#�2C���w|2�J荇�R�IᜢN�o6;�/}�C���k�ײL��w��co
�	�S[��^�{���L-l]�C�Ѳj�N���Ԏ����0��̜�3͜}~uh���D�}7�I������i�8���־؞ܵ��H����:.Tد)!��"*�%�	22A�!�&��y����%�۸d�ćB\���9(1M�M�Yo���q`�J��䊙���l�sd�ny�f<̊����{���m�m�v	N�.�>Z���;���7�9YQ^R�[ω'�ߍ�����l�8M�Eۅ��}J���\jl:)�v�V��ǣJ*S/g��g��qǚf9�EY�(HHG��2+��w�[K�0��@�l�,XWE;�c���J����l��߈�*�"	�����C��;剛2U�A޳궹W2���&<c�����`��dLV+KT�2ވqf�b�b~��ϛ�4$����J/KR�S������&Ȥ��)���������&?��������;�:F���)/�}�QC��K}�tS��&��ѡa�E�`ݔ��4%3hg�T�.���b�l�pL���~'[�b^cK俓LՍ�RG��]cg��)�Ԅhg��!L;K~V;��+�����$���3b��Z&�>l�QR�N���LB�+�d�!�q��#��P�9%i�$Fؼ�y�ɴQ�� �Ӿ����kZ�b�Bzs�^cw�~������f;M�7���~j�!������2�	Tj5퓍&wIs�nz��4���&n=�_�m�ꎟܻ��"�lh.�f��*��5�7.�Ιb}�ߏ�4,�=v!X�SN�����ф�.�4��'2��Uq���k^v��@�������w�peXAg����~����5V���l^�8�M˒�YV���ۿ����py_��f�'��埕�L��/��l�N�\.�)���f<!�h!\�3���К�,Hǡ��Y�o�.���m������Ã���U������'bC�A�RgN-C�������f��"e�Q(g�����&�\t���TM�5��ؕ`b�1
��1v�6s�K���ʉ0bN��%vy�G�k<��P�4mś�~��{�_:�`f���%��Ǽ���k'P����o�H5���������*��W����l��,��O�c�p�F����К]`��q���ܨ?��l5��IL�a����<-�����Tq@�X��B�1����8 �}p�*��zdｨ����G��/���P�m�]�� G���
�5)�^�8va�W<�RU�T�IL0�^eh�L�T Bc�e�S���'&�0����9��~�-�;��w�(Z�RV^�q03M��qB<�<�:$(z��qC�[銈m���Z�h3�ᴻ�����Yk+n�ӑ@KG=�v�0BÛ�%{��*b:�Q�W�g����ɿ�$i�d� �f��S�����+R�z�TV��Uo��U�L�����62��&!H����I�=X-�	�h�S�C�{�>`�����ϟ�H?��c���ߥ(��؂6��E�">���P<�M!���&����y�(v^���υ8�j-��t95r�'��X �A8�&��{{{��w6��q�5j�����SmF4��o�9(������w����qV�s��aG�)&(آ ,���lLAӶ�pO�0ul�4��`��CLA{r�����xm�7��Eq+b��F6"�S�u�W0�Y̧��m �[�������1e6����٠R�M�y���w�m�Y���C){�
�/��J� ��_]���bv*-����9��&���I
�`#Y��n��H�δ1@?Hs�\.�m��؟�]��+#���~����ÿ�]W�2R��ϟɜ|�����v�:g�g�q��
��2�����m�N���v�"/�)�_XoR:��?��H<O6��C�L���8�V�JOv�L���$�YH��3�UUU2+Ⱦ0�9C�|��ڑ�þ(�,Fi�O�p>-����~<���u��˚���(+u������Fw$_>� aP��/z��N�Tt ��i��;���uA:����q1��j )�"YI$7��*b��B+�t���ى~�ju��2%
��[���<pv��Eud� h$-�>���.�s���+#��B����a5c�	o,�U�	BKE�&�i�=��%<!������|���ψ3#�_�z�x�G>t��?6Z��fV�Ok���R��ѣ*��X|�XV�Łs�5C�ីӅ��B��U��:WQN\�SU�ʤ�v�D)�a`��-"�qS�6�9�	[�������M ?P>Ƌ���B�Z�b�}���ˮ���3ժ>n ���H��W���m�ݳ�����Q�oi	Q��b�Z���&�H�V�iw�+��3A�3��MH��&�iO�4�&({���b���ga2jg֓'Zh&���1&����[�{!}��w�̺��J�͙kd��[�5_T6�v��������`��sF�#��A�ᅛ�0くA�٫�p��D!<�s����(d$4Ch-tj3��ʨG&tD��+�:����#���L_5�GL�"��Iۄ��~ϺP�Z�.#&����X�+�hj4�"�a��(�\�<���y��*�]`[U5O!  `6���]}�����=��ϒM�΁K ���Ȯ��d�n
��y�K/Hd��^�CÄ6�yۦ�b�?߿_��j�ߦ�>�%�`P� ss���'���G���m���[�"xv�VVkhge�Y����Ê�q�γ��c���H"�UC8::�~��<�\�gl>x�r��0��ԱAM��H�l\��cw
NUխl!!,M���)l�vN��8C��Q˜���	��?k��b��hL8yV����d�"8L��/��nE�i�1�;���b�� ����^�v#ݸ~S�l�!0�I�9��ɭ�U�R�-�PZ��`|�♘�X��H.�]jAؘFub����,�������LG�8�Դ��s��u^\�����ݢ/_<�&$�O��͛7���:ai�ϴ"j6B�2Hi践��xR;�#�� �J@k=��܇ڐ���Lnct
�4S*�q�>t��@����s ��g�L�5�f\-�}�c=^V3  ��IDAT!C�`�d�k���я��qГNn/�R�CC����m�"�/��&}�ͷR%�1�q�S,���~+N���f�3S��F6N�V�h����Aύ}�t�����V�֠W���F)�K���?~R��t�
Z��.2�χ���kL8D8�[�y�	�ꔊ���c�S��bh_��頶���{6'�&[*�S�f;���lԌ���pX�EB"��������٠A�#+1���I"��g;?L=hy��,m�%��;�ơ�B�������h�h��-��}��1��}���Â�V��ѯ��_�Q��i��d��h]�W�^��f�WGJ�Xt��9pN<x��am�sߘ �@N�5n�?߯u�	eйἛ�O�T�9tf(�) h�9��j{���d�駟�K�J�hl)Ê �Y)V�Ǵ�%������R�y�	o	6YR%R����s BUo���˪�~��.�����>{�X*�P�6'\��%�d�Ȼh��n]�����@-6l�Z/MQ��.@��K��m��u������V�9�������P'�r��99���GJ�%�& G��pk�Ү�c���:l�b����
ݖ�T�)�٩	Aw %E_��b�-#K,7�K�Sjg��>��k��4����*�~/���`\,�G<��N����_b"�{�X��Aͧ��oR�ߡ�43�;>������W�㵇�P�a���"���o�ݻ��s��fgWk:�C[p/��k�E����%���[�����pk��ls��8gm�.dmb��Cn*̱�Ѧ����w�z)j|��j���l\׮^K{Y��$�&y��;�i�U���kR�ϊQ�&���B��!��ի��!��1>�[��z���?cr�Fl8aUh�+���R�����k�D
���ul�^��@�X�FAI8
J��s��>��bs¦;�_OW����R^x��Ku˴��9�,���m�w(��SJ����YT��}��*�Ys��;}&U��w` v�p�R�!�v�����4Tmnl��pbL��Cٍ�ѺI
�EH��ʄ*���6͜:51�0iQ[���R��!9�i�f������j�%��w����@5Qh0��B�T?۱�kj�8"y0��'�l|V5Shh_~�����dTa���˪��*�N��:x���x)� ��/�H7� Z˓��Od!�=���\�$�e�5j�dG�z���}͉gK}��T�-�x>�0�ꫯ�!�xh�^pܠ/��J�Yj�6o[ll�w)��R��ʬ�tj��v�A�g��A��7�y���^7�Cl���;�Ox'l��X������ăE���b�B`�mb쟿x�~��C��W~����!�;��846a�_���5O� ��~�}��+4v:�R��VdLnq+?����8��%S�N�������l�m<��5�������i��Bi�U�#�3���"t0����SN�����Ζ+ ��gx6c|��w�>�(o!�R��]��R2a��A�(��}(<�3GM�{@��q�
@:�o���UJ����b(���&������{ᜯ��*]�rUڠN&5C��Θ	�ʨ�3�&4Q����ݷ�	f�k4�Pq���X��wK��Һ�C�(�k�_ntZW��R	1A��8���#�c���P(I|HI�D�*�Fh����|�^hN���w�eĄX`b��U�� m�)�sf�{���s�E��|�����nb��n,��2��IE�ӷu#~R�����_����6�բ�PV��Łv�,:�$@_�[l�h'�SD`��~�p����N�R6�����A��4�?�(����f�S+u��7�uZj%N�L�5�^�R���MQC��i�m;���-Mܛ&���d�J��#1�TL���3bk���^%{h����/D�@˔r�A��ϚiM���h�gp՟K����Έ�{� �K2-Z%2j�-�"A(���z]�/��P�GՐ �	\�����B��`Zu��ćb�e3���,�Bh ����#��� �$w�H�ZJ����Ii�ݘH@�����*��ܾ]��KҮ[�o���e}'3�I��C#H8>�%nҩ�.��-���9�#�y��I�}���0��"��+�l�[M4h��,4�	s���Ï?ԍ�7qV"��*~8���^D;��ע� ��`ΠO�Rmm l�؀����V�e��ք���G:��˿n��Ǆ�����n�7���薾�4��̻�ACQ��~~9��hj#�ϴ�S��I�*��L�����'�b�I<��˄Ƥ�{ﮘ�X4R~�$�tZ��ɉN���>g���X/C�b�(&>4��z��.�h��D//5k�7�y0'a��D�v���8���Bx�T����kMj¬�	�w،I2����u� ���w���" �e�z�m��+�?�͍@ &+�!H�R6;-4��۵Z���U �+��e���.�o��V��P�=��Y�5����ܮ�ĝj�3E��82�~!�G�;̿������`� �M�RsJ�YU��	��_<sE�P�u�M�1 h���֍�V��B5]x��8��V�l��Al�a8������N����&7������2�Nʮ�L=��1�O<e�l�n��4G���<��:k:&&����{	�A<߷�~+&<�`��1��0��&F���3h�4��C��d�BkQl��f#$G��f-[�e�!1a������a�B�� ���OC;^%DBŗ��`VZ��ﱄ%{:m2S64�tfI>���3���7p;���Z������X9T��"*v*|f���������|�����q�`)-�z*\�SB����9�����mVX��,��#�	�Z�)k&�
Tu`a�={*��6���~�{髯�V�{���wfC`�0�/4��JC�a#����[���Y�+'�kG���c\�l���[�G�~:���0G�7�.�6��0*ӝ~
�8�Fa;يE�I�&�Į���n����J�NYv�&��CXv��	�)�(��^���\h	�ijb I2px���LC���Th��Ы�u�P��u�`1|��g�A(9�
Ly'���5������l����0!̰�mp�$�:�����nH��s���U�ͣ%�|	�12%f^C��6�0���2�Dê}�_��_�Շ%��jGpH&�vz�[�{V��w��5�l�)�-&O�B� {��XJ���J���s��쩻w�v9��ٕ�����G|0``�/���>�����w��G���o$&�m���M��גz��魪�b����^�sBW��L4��W�ӶG��hU��|$��|N������g����S��.�o������)O(�m����z�b\�:#�A	��Ǭ'w����B���|?h������qw���J�f7�:Z�����3���U�4�Is��6�X����@�pюy(F�2���粏�5��H�x�:�5�g}����M^��&��3�f��.vH������"�]d��6��8�'K���K�I�-��06h�B������@mN�v���w�/�<f���`Fs\b<�
��0]ٿZ�-��I��y�+h��T�'���/�fe*6�;a|'�!7�����Z�}h�b	��cS��aZ1�d�(�
 "8���؝˽p=���k��s����-[�C��1?�̝}�o~g|��@m����uN�m������9�JUIi*���?ٻξm��Z�h�	^Z|�R0/��0o������G������vp\��h��T���"�V�5b����6��gfAC�f+���^�D�3	m�� Li
�am��@�a���)·�L6P�a�}�l�0���B�����G^�Y��H�i�Ԝ�9t����
iE�m���FK�AA��u,l2�ú�R�7�e�xg��6d酥՜b%jJ=�i��o8�[���Q7���|(��_|�e���?��>F	�x������	bLp_D0@�II��ʆo�#
�=�TX/p�}��w�p��U�<e�f3�{]x0?��@�%�W�HKqo	˫�DS�q��f�3���xS��� X�O���Nq��@�	��Cj�lX=�X�G�f�x�C��L�Ri&>��3ĺ��G}�p!3���yhG+�"�A���]�/��DF���M�)�[T0�����X��!%A@D����N�_L�b�"�	YDX�G�
!��/Ne��[f��.\C��oē�E �?��3#���o���.��
:���H�ڪj�*�,�o�:��x��i������߅�ͥ#mE�y�&���#�sF�؜ -޸��ԲП4�GR����	9�"4R&馶�C�`�AJ'"$!��}�^�p�0������R��/.�(t���Mep�?��,��U��y�x��{A��/�@U���r� ݼ�΅+�Ly`���8gO���w�w#�PC���4�Z�3l4���P.j�p,"��]=�w#_��$m�!h���7u
�La��r橷6�b-���c�}7��h�Q��n�N+v�F��v�)��3��V-s��7��떡5rڑ��d�0��Z̦�6����*�{�E����9*D %�!5Ar��m_�ZOJκ��D�9�BegxF�J�P��B�L;Rh�����+���K3M��"f�O���z�/���>���8���2��@��.2a���}�q�{FG�^� ���Jd�����tW�������ٔ�yД�	��eUF7�hV7J=�V��T�
h^um�q��?��� A<���B��zdRI�R��<�Q1�d�,Fx�9a�,0�7���_@�J�_nߺ�>��s^{ڭ����k׮�@E��C�!�y����hd
��(�&�g�R��2*F����Z$柰H�ł��"�&>6a��������'X#
 �1��ي�  �gB1�Ïyr�;��v��?�>��"��"��L�KM'W��f���~��)��V�COk����p���ܞ��뜭q	�V3G�i	�wL�D�%�~>��"2LF1���T��S[��=���.*,<h�8���DB�V0S�a���V�-&U8v�܂Z��&MuZ{��}Q�nf���9�dYv���*�H��-}T�M~��ר�I���P���+����L/}&/B���2�v,|��R�i��oA�4'��Y_L>%��(ϤO�p:6�lۊ12-��N��k؞�������@ӆ�!LY�YW�cX���N5�٥˦�&~�E)p��5�+�I��V`R�!;X3�:@��������L���[�|�Q�e�c�aRqImN(d��!��T�d�o<�2���A7��$&滑_՟��a��^|HLe��|ؑ��Ǥ�1��3Ϝ'-�(��I�L���g��9jՅL�&�f��?w,@�T�KjZ}d����Ex�^�cq�$"��W�h�a�v!��/3��V��-�kV�H-D�Cw�L�Qkh�E)ˡ�j�a�{Sc���+cjYSaC����6��J#�^��J~�Q.Rj%{�>��o�	�Y6�$�����P���/��3���	��s��lz�g)-��E���>�Ӯ���d0�����3��!����D����v~YL}�7��� ~����+�}'B_b�_�w)��eD)�I�4�@j]-v���}�x�� �p��t��U�"����#*\_짍���.
��L�F!X��i�i��ύ��^k�gߑ.ܬ�6#��~{�SIC�79ޚ�NɤE�D�)��_д��XwGL%�������鄠{[8��a���.w� |o�bH������4X#���
�eP���*LI\��ba�Z��)G*AѢo�O����C9�W�U�Ь���e�mf�]�<c:�����t�39����^N#Vy)����D��^A��o5�t�x/�A҇��K�ϒ���I�<�^�Z��B�lLsj�"(�F��f,��3% ��h;zn�1�����M:]%؜L���?��E ��~����<�{l��x5�X��L����/���pĵ�O�ޠ��}�N�/����ŝ���_X�=��y��O���A��.4�F7��N,c�J����`�-*a۵]W�#���o�Ҷ�q4�P9>��aMJ�A�xV�GA`B;`J�
͔�|eτ7�}`�ǂ�)���;qF�x�B�c8.�,�]'�{%��R@�l,B4��W�"ƹ�%W�C�D k�8�A�T*@教���I�+IMT�kɮ������!��u�~�/�q�1�E"�Ԣp,��~#��FR.%��Z�����SM����cO�	���B0|��vZA6#��Cv�m����m�Z8�>c�>�Wh�Z�s��`���P�0�U���S�\x6��_�5�y�Z6Qh���1����RH1�����%��Ν;�/pU���0��V�u5"�^j��z���i��/���3�s���Og�c�N��D��1��&e�*a�������h����¼�⠘����L����ґ�c�
Ќ#|�q>�y >ɔ���^�o�"��W��»:����K/�(T�Ґ��k�Xp~�|�R�\��R%��
�V�6��(>x���~4Ȩ�=�|��Q�j�,Q��%�g�p�j3��)he�G��X\����
:���e�ءO%u:>{_�M5��iR̴b�0'	6�����m��~z^;TTæ��~��\�h4�gCt�$&Yl����S��4�e%�=7�V��x.0�+���\X8�^���Ҩ�X��%uWRl�r_�����@�H��ۺ��m�-�/)A
�MA3��K
i��_~�p5@@3\ߡ/R�w@��G{=�Y�g�N�����<�*t�2>�)�CBF+�q�?�\"͚����(�y�����F���L�UT�������� af��ӄ�a6�gf�)0��1iR���h�/�-$������������ ?ĳ5���W��bq�AB��������Vq �x�=@@�M�`�e�0�+�
-�Wq��F	�m��x�����o:��	� t�6E�$hs+�(K�g1�-�"��ˆ�MЦ 5�M(��M���Ԇ]bL `���ƥ����R���:�^̌b��ԣ�/�@�	T����7�ފ�g��U� /�>L�	����Il�!W{l寵P�:��`�@��x�L+6�=�{:u�p�E5Ә�k����Q��fa/�1�bI�Ɏ�Gc.�z�*]}wU�%��-�Mq�щ���`��wpJ����1ԖO��/Wͧ���Q�X�=��w)�؁��d3�����zM$�+�9Gg��[�M�#g$��\�Q8.M�V/6&>Bb�!񄻻���ZQ@����M��܈(�y�l �%����˖,@���xBI �S��c�k�"��(8����(+I4�i��3��@#$�� -��o���ǒ_oV�J�0�L2�`��KR�!���	IS��ߋ��m�[]�ёnn"`j; nߺ-LK��4{I5^a�s��ȱi�fj`���+"�IƲ�G�(�$����3Z��z�j!6��	샿5�t�bUJ����Ԍ0����]K�_�L=T���,��B�r��p2

�K6��J7Ø�y�1\�vU|�I}�60�=&4%�֨��9�2Y�':��OS�$������
F��s�."���Qn2U��D�	6������i���/9�Z$P?T�7�"��ݛ8�Y�L�������\�}_0֥NV/ng&"�g��W����ԯ%����Q +оV̤'�L9;3�
�U3�M�#��>_����x�j�W��]���U[��x��eYL0�h��z#!ipP�R����jv�K&,4|�4���|���A4pFC�w�h���,�_���RJm�� S��YLjw��|�&MW&L+�27v,��E��P��&(-��A��ٷ��W�^�[7nҍ�p��]e�ߕq=x��8�`M ������*�d0�|67��xB��k6� �A��N�_-�"�%��0�̪c9ouB��r�bs�s~�M�'�P�9�wq�ell�A����k���Y��M�mtٜ�d��R��K�㦅3�=%��T3���,7�v�v.��D��)�NuQ@�B�3.5�i`�^��K��p����G%�5l��炠��/�t�����L���k���$%�n	�a��-^Z�dh5���xЪ��V�;`h:��Z����㫑%h�]�|���� �f�"��|!i���o!�^u��ņs$0�a7��k�8��*a����'7JGl`o�HM,8�0���K*��J�!D��;6Dh�S<,�*�:Y:+ݾ���9�FP���߅}
07Zh�p&�v�/s���|6�HV+f�$��BK�HYȧ
���gZ�!:{mM�&a��)B��#�)�iGn�ױ�5�})���f��������\X6�����\T���P����GpvqQض,��͋�Q
�[�d�̈5^��B�7{�s�E{*�+PRt�$���l4aK� ��څ���)�ͬX�Y�Ҵ���/ O�f�Ɗ z�´�&���'���zd�ȁ�_R�;�B���٣f��#����6jL� <�1�/s��fie��?H�Ms6tYP�1����h��2߼Ѫ��+:��ǦY�Moq.�8�T��A0��~�@=88�L7� '���g��ŘôVrh��	ݰ����G�>�'�Z\���+�� ���%!���/{X�B�*�u�Ю����
!��'����E�_�=A�~���gE����sgW��הAa���aS���ϸ��h��(CcY�l`G�r�u���OzC�s�q�g�4E<D��7u�h&o��Q� @:ݻ��29q�h�+�3�0����@'�΅XE�=~���aV:�������eq�INm��SY���;��<�/p�jUQC�?q�(&��Ѩ�wr��H�������e1Q�	G$�f�X\tR/�����K#5a�?=���U�hR+�[�\;�֊�9�qҨ	}�H��)��,p�LwU���O�1ycsd��+�ߠ�b�D{ȧ`[���2_�OYa"`�G ĩ� �o�j�ڃ }� 7n"��N���aݗ|�CT�,��s���+��|Ŧ�kT%�iO��#q����Q��j�W[������0���bp�(C�枾{����[��Ķ��o~�=�XC��R;�Ƕ�C +��~t��㵋��RD�Z�ѫ�N\���&3���Ke��ef��;�X=V����T�v�q=Z�/,�03���Z�J��	�Tr�x+ON�s �X�� IP`M3rZ��gE٬�K7.�,�>��g���ދ q�3[�Q��9�$�2�"�.�	Bءb�C�~g��<�0g_D�g6S���뉡��/�e�b����?Xj6�Ss� ��=�y����~�$Q��ZT��}���B����[��Q����H�K�\ZRQ���E	���3�qh��:%۬��e�M�W���^h��N������?���~I��ۑ�Nط��I���ݽ#�'�⾸wO��f��l�#nH���&}O%_��>��Y}���f6ؚ!I5Iv�)�p����?v���~_eFݱh�ĩy�q&U:i�����Sn��]�� ��ގأ9��o�	HU�"�Ò��`�_%�j?l^jm�C��m�mj��), �@��{�v%ڥih�4
=;���HNΥ�'���q5I�Ӊ�λ�s��������]%Q(lQL�x�	0�B��p4><�7f�pz�vZ)�|��4uϟb�à!cوy�o�ێ��p�i����{:Ϥ���jM���l�b�x	e��zn}m<��4A��ߦ
K�V������mr#F'��������ŵw��Y>�pA=�L"��h���%qd�w�j�RP6ɢ��bG�'�|n�����9%��6���n�O����{YC�Ȝ$�9��%��fLa�i�ݩ��9�����t�S !����p� FH��&���rK�l
BX��x	��*L�^8Z7M"� �g�<s��	���&5;}���u��P X~�9���6X����)'&��ɹ8���mLܭfo�ȁ�vP 3��� sW�1~t�h̩�c���վ*���e��ډ��8ęA�J�A&8�e���B��-$b:4�`�c�)9���Jؿ��-��fCs��}DhY��j�U\qD�lBs�	b�L{�J��|�`qs����w�HF3��-��W,x������t5j%����m�XHr�W���^?���f1�j=�i��䁲��7S���F���f�PjJ��t�����Եk]��v���L�ܞ�YJa�e�j�����T���3�u�{�M��'߳)�*�����'y2��b�p��쇕�^qG,��lV�e �=�װ,ӛ������<�&�)PY?$��}�V�XK���,�����Hy��dS(�f
�����K�n��i�А[z/����SbR�ʲ��h�E���H�ɛ��� �6ȨO�Ώ}!)o�[�w|����D�(F�T�L�G���&Ƹ�|ԓT��n%H�y�y&A��V|�	n����}��ŸZ*���
������Cԛ��E��ޙBe݄�X�_3�L�i�)�G�N��{���:v��%�������u���f��F�L��m�9�a��������x/�k�3������X��8b�N�[��ĭ���'�wd���|
fIl�unk7��A��6�:����iz�d������e�HKioE����v?�u[�t�:��Z��C���@��M�e� .S��߮i��G��:Y|��͆\�f����x�a��ͥh�;����ǳ�	�%��$ǐ���Q�1γm Mȑj-j�Qh�g��4)j��6;��a�'����Ip��������ۻ~��bM�YkYx���\YRs��yύSK��zD�<�9~�{Nӥ�Ԣv7�3��0ju�-�t��v A����M�����VY`i�U��侦�T0,4b�y4��6o
KZ1z�
�&���ݜMВ�"Z���mN�U�m�+��S:q���/}�3M&��|�r����^g@J�ݞ�2<���	K:S�`{G
�ɋ��;�������ɍ�]�G��ǹ������i�y��i�p����"�]�E�i�A�F���/JX��� ��*�K#R/��{�&cW4f��E|xs��V�[	�Af~��Za@
��36���y��So�SG��o/Lo9�����Ni:"�bN�a�c�6����Yl�>��Ij>��& M����-9k$�
v������km���|S|�9<9��`��b�Dੱ���P U�@�����4u ��s� ���VN\�y㯛�ik��(���K�N/%��?�M9�.�~��ߡ�>�ot�����ޫR��Q��{���hK��� m~f��-��J��YBp6�f@+u>�StP���fq\X2�F�yܛQf`�V��)��
B�Ǿ�A#�&��q8��8�R�=� ��`��x}����H }wM��z����SH�����Vp����G����2Tb���gO�5Î5�tTGˤ����c���8Ͱi��ҧ�t\,CCv���a��柷�i���M�(������O���kMs��D��M*���Qyg�fk�o�e��
�4i�n)!{���GIA����lRI��*-���k�z�:���Dܿ��h��Ў��֤i�blEh�Vdq,5Zz����%�Gl1�-�:��u�ǧ�)忘~D-��A4=\30�r��5�?�ny0������-'p$�m�˔�4��oN�a�L��Z�e�-b�x}{.ئA�]M��p�?m�s��n�����:w���]�<��%#v�n�f�/\����ڢ�\{�<}-$I^�!����i������ڙ����78ַ��Á�Y�,�Kٸ�t�U^H&Dyt�0td�"fE���	7���17Sj��1�z��߾�y�ֵ�c���F��;co����
����ݺ]�ػ�U�g�L�}�5[���C�E�%.Dy_�Q�	+�1�g	��ĸ�>�3�7����$���]�	���Ɖ��t�W]�Wo.��Y3�8�7	��,�=h=�ݓ�Mp�Er�'�#^gZ���(e��̭�<��׀�������m�@m���VG|�b�m�dn=�i��8�Iؤsn���;'Js@5K"���s�����ùM�H��~�3m�LEjp�DY��:ǧ���0q0�/�bB�q��Ʀ�1Gؑ�;�+p�0��"���@#
T���e��uc����&�\3B����u~��^4�z�z��l
k�����ЛY���֎Nk����5޽Yw����R/4ܒ	בe�sL�-���[ zj��!�������Y�W��C��$�f&j�����w�K���8�4L�����z�i�zQ������*'�L��a��hJ�`��n������>,�2X��_�8�V��g�qߧ�V01ݹcE�T�+\`0+c4�0Y�U(ʦ�SA 5U4�0("R���N��)R���wg���r�B�8?֏��?T7s�m1�Ȧ�B���%S�ܹbfX��ڂ{ʽ������r�Cq��4{�8Y�����9�	_ �o��B�O((��*�r���!�=��V�>��Ӷwq��a��S�O�a��{ns��-�c�{�'ZBܬK�*eΛ��M��v4�ʻ��qL���������>�x5[��L�ԝ֜�\�Qk�Mܩ�$z�����2����q.u}:��]c�/�&֏Ql�P2�w:�\3���	�'�L��eZ��f�M�Q��VNoui� I?�^N�:�Y��ƣ���M��?������z��֤�l��c���	̊���?{���ȍmA2��Lɴ�6�u��y�o���'s��9ݭ�7%�MCk;l @&�����e%3���E�8�9n��[:��5�����w����y�I��ԁ��n}G�_�2@�uٌ"N�����b'�^t���cqV� ��_�-d^:
�w=��d��G�b`Oo�T����P��$w���=*r�B�ĩ�)��B��\Xft����w���=cO��,/�*��?��}���)��j*I��8F�)�.ʶ.WޘRZ0��:g�~C�r�T�:J�.c���e���%	��/P�t(bț�yNc�������Nl�&:������Q~Չx�k�mT��z�""�p]S~g�6"�m!��Z�C��Y�c0w;Nl�0@UI�'�E]���޷b�W\.P�^_���zƶ���'��H��D���c��zc��[@�	В��ri
yv�2u��}��$>��3f�qڲH�Nl��W�`�hoi�q^����r��Uw�aٲ('��i�P��B!�H�e���k ��c����S�F��ω[�2�E�jz,�� �٪���*����f�՚��&U�Cq��͔��m8O� 2�Y3b�'�ύ�����r[���|^_�欚�y�:[�s@�\�p5����z�d#���,c,�n���h��;r +/ɑ��/����N�2���&�hJ�b����P��>�Nf�K�x��������Ь:�	�k�3$�>sOj����o�]rnL���X��YO�g#[�@��埵%��j�#�{���E�}Q�^�?��<���%�K�sM
�F�ѾX'����������駟Y6��|�}�5[�Ю�`��A�)��o_���)�$N���_Qc]��V��E��B1J�X�ӝ�o7Gu"}sA񕕿�T�c]B俤F��B{.����g lF,<��`V�0��:? \�Vi�ЉrU�R��.���ӧ��~�!���/�/	P�������<c�-lӭ��E%���Ъ:�E���-������������A����n�lr���^���=Ǩ�!�m/6�k7�CZ�'O>歉��f��M�i!��\��3s�ظf^�:q+�,GS4�ܽ��}�����a��g(�θR���yx�����Y�ٷ�����8��/ip 굔�+C��}��^��}`�V�T(�iذ��5�+֡��q��}L��V@�i�e%�7��a}�	`�Su؆�t� L�=�#|��7�Q���і(�g���3�Ruk�A�����i��� 1٫�fy�0�/���YW=V�f]���4z:�=�ݧT*�@̋�yx��%�'0U��;"�)n���so�ͺ�Q��2WG]K�{��¶ �Z��|�1�WQ�-^�	f'j��x���>4q�����4�`��3hb���ǳ���?���E>a���b{�'O>	O>���Š��H6�H���=��ڻ�׵�e�^�vs�a��JUD���4& �c;�3�1R�B�Á���slۗw�4�y����#&��߬WR.��7g��q*���׫H����_cekq��|X\�uC}�YC�H�Q��m�yK�{[��qB{ů��.,s��Zė���[.C��y��M������a	�C�! �M깴���z�;rL�`��W���:Z�xpbH<@m������̊pe��m�K�o=g���oq�RN�c�I�"�LY�V�����he�-�� o�T��y����-(�o{sК����� ��4ȑ u���������n�����a��Q��H�6�m��\�����u�%S��닂[�po���ǫ|e�ͤ��8��S��Q��.�Ey�h�!������B�^�s��&|A\���֣���zM�CFU׭qڪ[��v�㮄6���lDd�8�#q��P��~﮷��ߤ ���*M4¾�QS8�U��\�p �=~/�AŘ�ԌHN��2�-�m}'H�U��UDW�Y�aT��^�����U��n�GB�U�h(�0����FITB�' ���_�-�
���J�� �m!;%b���f7c,�V��K��>��5ZcXR�pԴN2�b�u8=;��QX��!�;� ����0<|��H̑K�>�q0�0���~nQ*��F�Q���
G�iW��ːN7���Q��I1̕�
�>H��4MwԤ��$�	$�6��O �&��ld[�D��,BCf�粋��ZS���)T6O���huLz�A�N3�C�c�G�Ċ4�6�f���&���xI�:y}��6���|���ܛ�m�X�O~[�s7vO@�8x����D���\K�zD���^v|O��^1w"�e�@m�������>_�ϰ�0��CY�TʡEdaϨ�tky��ryL�8��o�?���NQv�]нy�1�Q2���.V�54���/h.�䶾wt���UN����az��n����-sQPjjŕT*i�KdΛ���'�QJ_	*���+���wEXA�B�4�	�(&k�懗Kf�u�*�*G�+�� �� 5��,V��� ��L �<�h@�Z)I߂l�k�'��<	V� <�	��3�i��X��o�BI6Nj$�Cbf��D]�s�<G�´0ᏗGR(g��<؋��zx7,��� B�9����(�7�%��8��cX P�	ȱ��h���k�]:u;_0���ek��M�y�@j�Űb�9��<>e���gd�BcnL?��V�9,%�P�:� U6gS���q��+����+���!��դL6�!��脋�7�+ԡ��n����%]�9Kg�+�t���u�h/e�)��mla�D5�Hm����u�:d��`A����s�a�R�ֽ�)G{A�B*����d:m�J���m=�:�gOq���BT�U�R*��3�H���^��Jq%`�ŉ�gHw*.���6�ӿy�ִ�N�`Yb+h�eJv��6K'P�H����s��P���i����1�И<�e�9O����4�Me��uCAa`�����S��|�	�e��!�^f��dp8=���qJ�fU�ނ�Σ�H�Č&�h�I�π�����-E"�ԁy� 񘪍q��)n(y,��Ld��e�Q���&�&w :�LC:��2���(�G������KuDi
�I�?ZbxI�d�-O3�~}���C��z��&�&Κ�PKh�3[����s�\I����Ҽm���X��~�~�34���7d_zZ����˱rmW�)��L���̓�S:�)��Iv8�{�=h+sgeLz���4EY�R�NK�{���
-m�a�{��`�7Ib��]�Fe+��2���X���X�v4
���#�����a��E3�Ϻ@���XV֒�Q{'�:�uuy0!G�ZS�-�I�n4@iYg����rq
4��
i�%��P�TV-��,�v5�jN)�Ny�g�:����,,2Є�PݯN��NVe;kL&�����2�s���P����[&s�&`p�P��u��@ܧ�����3������A�Z]��yzr�N������x�����cѧ��e�y���������g�4!�$ q��=���L�m�_�z^�|��U��'��G������=�������� �\�l ����\\s?�be�yK�ٳ�ؾ����ً�<��z�*�I~�M��>]��G�=p�˗/�N��6�}wt|D����yx.�'�&��7E�	���f��P��K`J��U:�9���}���!'K_�b�2z��u9��ǹ��Y-#S���.����d���qU˚m�cd�gꉠz`���w�Ők�e/�{�@�4�A4�х�����3��7���o���dKvf�݃�j�� ��NJ�؛?w������O&��uL$]E��ցl?�/�N!=dR�I"���2k�=H��P2u�3�(���R��z��c� ���a�Y�@�,��
��5a"���\��PY��fz�.3�^�IG1��&��< ��% ��D��e�H?J��E�Fshl����P��,&:��9OP��	��Й�gy�Cܼ���'@-��\���/��?�~���*�{ƅ�����f�{�� �a�{`�G��h�y @?��s���o������D�F�?��#
����Y`d �P�������_��Wx��%-"h �|���!oǝ�_z��ze�nLO3���0|�6���;TV�������_)���X��P���ۯ|_��T6��x��b��\I/2�L&p�":W��t�:/��lx,�z6'���ws�S�����>��ʔ|U�T&�}�k	<�$b�z"�O�MݿX��*��v����k9 �U��T�R� ��	���A�Gz7Z��/�O3��#9�y�� �¹u�r%��4���t��H~���(CjU��k��m�RE� �?��GT+����ϟ=Oό�_hR��K�5�����O?�4|��gP ��d�_�o,&(O�d�S�/D����	��ӏ�Yf�p�"�xW�- �����_�X�J%�ڣ\�����"� �,�ϟ���>����d�����΢u�w�.L4�s���d���느^���?�`l ���q%��>f0����O>���Ԙ%�
��������#���s��ˌ�_#����(ba�h�*��+�����ȁ��WT�'�Ë\�?r�������ᗟ&VN�23,����o�E�7�ɚ�m���������Lv�(LR�2Ii�`{���X��� �֞i�y�̫d$<��}��h3̙(���A��P~/T�ǪaR��X9�O�* 
��窚��[R�V�OoP�B�$	A�B;�ty�?zp/������$f/�X��n�%Wlg�휼zV�ð̬".�h�}	��d*��Q�բ����3�^
zP���{�߫�o5�	
�!��8
=�	�7�������w�}�Y���b0A�nWK�_AO|F�	��}�E�?���n�(i�bq�"=m��`h�e������(�?~'�ƹ�E/�攐c��w����s;��x�����/%�d|���6�G�UddR��m��� �W��e:�5'�QP&������>����<�5�{W�%���[`���;��a����@�s��Ԟ/:X0y<� {�y���9����o�E$���ӧ� K��E��D?<��)1֔�M��6��0����9Rc���^L���KO�����	r9��S���ms�Kv������-=�UpC�P�^D����D�N-90�m�r�xu��oPKs��"�#��r �yB�5����pz�!}*��2$��1��>���1B�	�y��%ۊtO+�`1J����4�N��Z�-E�$����e�������B>�}-��A��#�x�>��?��A�{b1���1MնR}a�p��H�����}���ٟ>'VQw%��^W�vҷ���=���g�>�7��wXO�����69y/]֤r`}�fŢ�!���ܸԊ�����u�>3��E�*n4y2��t���YE��K�68��mS�����("6����n�|���PųB@��b��ږ5�2�g��?����u;�~�w_���`����:T�Gfu�N�i\�[�5�V~5@����x*�I���So� ��\
峛��I=Txw�p��b�����M��~��H܎��CM�!�]Y���o���CF}O58�;^�p�eRr�ץ�gN@��<���*�CĂXy��UXg6���l�V�db�3=1�<hO3;Zf� vx��A	`�N��QI�Ʌ���)�C�`u�	���w�*����U+�Z�5�%>� ������w�~Gb8�k�|ad%_��%��,�`� E��102 *�@��-* �^���G~���,��8��t]�=C�g� I4]��$0S���w'�QX���O���s�;��32�A��g�ŒM��-وcTXh Bx�(�#Ó��#aC̙h֋A�f*�����b��Kx��_��\� ԏ�r=�=<�,�ۇ���~�#�w�� i�;�~�{�)xweܐ0NN�߿w_�\�]ISuRHl�:�����*��NĮP#�H���Ѡ~��LU
��U�l|�L�5Tתz�GO�\>�'��ĭ��yZ虑I+{�d@8��QV�%���jM��4�s��͑��E�wu-
�o�q�ߗmЊ2��z�E����<���v�T�|�y!�|�� >y��C8�$CƢt�l8'd+z0��&d���PGT_vb���`#p�I�Q�)�-�����4��e��&��MDLcf2���F�?���M�L����q�e�����R[�� LD~\W���	������(��1�,�S��rE�Nݤh��]
C���
m��MF���1酿����y���t`q`��^�2�|��j ?  ��	��f����xb��1P��»��w�``��t�A��,	K �/WˠN�`�P@����C_r�,!m���_`w4�k�,$'��8y[����w��s��@Is�(A�+���d��ҁl谁�	c	Z��8��n�8h�T��Q�}�NEwځ&5~)0[���4�y$�]��0KN�f p�EB�͂e/�l�V��JMt������T�%+�s�<ȃ���GF�!�C�����Eƽ< 2��fѕ({ �ҩ1��8@�%�8�ݢt!�ډFF���F��g�"
��������瑷��X
ۯ���>e�/3��(ޣ4m�Ly�'�-z*���o���xQVhnb~	LpL�� �O��za� �6I��}'��;b��lIb���	-�+J�XdT��$��``�A[X��q U��+|����/�_~�e���O��}HV|��y���t��	��$����z�nq�:X�Y\�A�ܚ��$"��O@4���@Gz[�*����ft*,{-lXT�� ?�� �ot;��W�ﾥ��E���5��>~��H�Ņ�ƻb�Ӕ��e�B*#��Y��#�"�"R$�hH���R$*2bnJ�_������H�&���YI����*��t�;@e�l��I�J�e�ѐ�wX�H*���{|�E��=rM]����ZÂB,����PQ�QCŴ���Hs?b��E��0�h��FdP�`YFV��i�9YE� �y`�����H�b���D�ď�As�;2��"��*8�1Fdف6%3>cR�`q��B��D��b��_�����_@�8�z����T�NEQA�IaB�'YDV�ƀ�d�B�W s���3�h���믿�1�ַ�:�`��XT P d(����&-.X<�`ȁ*�qf�����_��ȿ>|@�$��~��G2����O�f�z&����(��e^��3��#̏ ���y�����f��^����q? �~�X@��UYQFq�WR�o12����t8��ի�t�G������S2�)�ճ�oP�@�/��m�"^ ib-FD�x @�����Sx��3$�u �&6�I�}Jcߒ�Ś�;�:Ό���BP�U��G��dzޖ	Z���?�~qa�>A'k��X��~���`(�Ev��~x���Q^�@��}>y��^��.9��r��j"C,�!�P(�8�x"�8��XjDF�2Ơ����iH���w���I��$]C�g�����X��yp塚W���K2r��>��R��6e4P��Z�,9+�dD�1{��R��1[��
v�V⨿��Ւ]�4���,���S�T��>��qDbj���x�c-u�&]�Z��������W�3=��T�����j�PQ'��}>�@�ş�D���}���߅!��؛��1��=�=K�IEE0I�3����%�V_Vb���x޿���q��*T���2�A<�H����;�
@�&��F}9�}���`:���G�O�����9`� v�45-�G��d��ܢӰ����ޕ� �@��:��>�`7�����D}�'�6��y��=O�5U�# ���Ə,jþ�<?������uGK-#�pS�*TQ��Q�O�;�y;p � &dW�рiZ,"�9�U/�{���&t���(it^8�Q�S�w?��a��,/^����B�^7��-w��b�����\9C�ΐ���Q�dV�?�u�D�(�Q����.8����GyUBƩ����~�b�m��:�N�,T��AtN�ٚ�9Ƀ�E��z=|�(��,>������ zV�q�z�!�Wpp�Pj"�#tlQT��7`t� �D�R��a����5D]���O' RH���'�Yd |FL����ڳ�uK��q/ 41�?O�[�3ƍ=��	�������z`P�;�1%速�9�xWf�P��9:d�/�:�(A��C&������$ �AW��CL<��?��?����2� M�H�-�[}��"1��?7���:F�Z�9�{�9#w-���\�`���iႤsĉh���[ڄ��kQ5��T&Kƴ|?��g�}�%��P�+ s�U��ǟ��K��(����^ 5QۓKj`���ʿ��c8��- ����"�i�A1���g�Zl� -X�i��"��|���Acn3Ʋ���ċ�B��>�PQ�	T�w�� �X&��E�x=��ȓ!3�\׳L~���瀨�G��'u,�yp�FD~29Ex�Y�BL(-��`/=Ϋxe��p2f�V���=(��V]�0��Fu��M��YXg�|��3���9
0����5�%�c`� �$X�3j(�����J����力]�T��%�F0����������s��|A�X�� �+�_�,yE,8SX@Y��t�`�؈��\r��a�%$� �<Z?$Ƌ���ً��u�����e������0�ί�rcZ--�V]_ V��7l@�D�
����0� �^�+ꖍ�c�I+�(Ɏ �Ѩ��V�f��+X���<��}�ДUm�&�j}�`�^�J �v���ɓ'�P�3���dĂ4 �q���b�J<1x؍����4�GN.��3�b7�Y�[
�_��ڮFWU�RZ�["ŨٙDX6����6_KQI`�B��֡2��T'*7�azO}NCs��1��������d���(�QV��H��	�Y�p���t��s���-���(Lh���^��h:f &�f�yp̆
1��41>�_g0���D���G����V�3����<�n@d%y�x���,�VL�����H���(jf0;���8���
5��Hb�1i9��1���ù�F�7�3
��a�J���0h���L:gU_H+MZ�<�9����Sz��(��*H$�ȣ�������-1bMF�F��:$B?�0��h��2֦"��GH����mX9���!�F��g��Ң��H)�,�F����Z^����I��?m�'��f��R��fѲD+�U.An������ʈt�>��"?T$5�Q5��_��������ŝ�U���1��0U�Łk`f��5�EKy��c�$����RY����xǅ 0�Ml,WQn���>c��ʋN�-y�t5;Γ�񇜾���,<?G��(]��X�`G}9�y�,�'�B�E2(-��Γ_��%"gp-�h��N�슒��TwU��_���i�F��M4M�K.�,��Ơ�Q9�tN)�ǚ&�J���(�2�X�R �E�	a�d�5� cU'���G�̆��[���	R��$Yuq41*��fX0�o%���e	�\2�I�R�W�O�R@��&��L����������D�X�L��ɔ/��R��m�@��ho�����>�XNn;�,����#D�8T��3و��|Syw5��v�����hL���uBe3�?�̾���פO����b���Om��ς$�1���X>������wNT���A3}Q@���1H��h�J~,����Bq�R��Ƞ�C�4:���r���H�u����(I<ƴ&��WV��+��Cz���,���S�7� �4�7"�Ujm�	��L1��
��r>Er'�˂|U�S�a^��CQ6�T�Re}:�����sb�Hp�J �D�������4�i��u�n<xPG�Rg�VlX�1�e�1�ġNYp�+��d`�!�?��y|ϡ�`�e��<dRJ}!����^�Fp!�(�,(k��u��p��'��E�����J@f
0F�=I��ekoU��b(��i�aZ@5�Fb)J���={�P?
j�䲖 Օ���;)���Ȯ\P������'�_�{�{�����^PV7?�mf�ߗ�/x<���x%ޟ�Vs�O3�ܠ������w�Q,��LN��ƍ�g����n��a:D������M��D� �h�9�4��sƲ��эǅ��Q��U�T/"�飼}f� �I�@�,��{,A�E���`�j}FII�SA۶�����R��>|�E��$7�\�C��fm�.�B�ۢ�1yCWR�&P������}_&��Tjm�0Q1��peO��]���
��xr?�����|99�ǆ7{��T�_���rLR�~���0��,� ,x@��M� ��Mـ�DE�u��E~�x���J�|Y�MEeʒ%�](�^/�m2hB,Д�=ܕ5�Jj?S]�����<�H�1n�n�HZR�^����$?��\��0$�J�(., p�A�ls�]
� w� 5@��@l�U �u�Aq�U���.k�X��j�	c�*n���e��t�`b
�݋�� ,�Q�s���*�"g��d�C�#"�`�Ԩ>���4�~G�]ӡ�T�pRxu�
|h,4J%Η'�*�ԇ���������WY�Mj�r+�.NI%�E4b?�5=�:r`���q�h�>�Ě(�G�qh�V�Z)�r���5���b���B��G����c��x����x�W)<ً^��Ǚ�|��禗��`��D&������A��C7&7�)cC�T�-_�K6�b��$�ą�v���A �թ�(G	�u�D
�_)��I�6��0�T(zRMy7:�����R��,(+X0ݤzN(i#=��ǓS�yo�w�l�$����W�YL���+���V���ʍ�Tp��XP�Ht����xhF�(��,?g%?d���8���Ye��R^���(X0�,Be�;pL�=tbTsđ�:^E�[[~��^$Iu��0��'�|�>��BiWz����@Vd�����W��q��ӅU�"��G��+7��hT$�]
hp�XS꼳<H��@]�8���4���+ʛ��D��u_뉳�����nD�"�z�FT��-���:�p$�TqEg����${QLam>w�3	G%��#bG��34�.dP@��r0O���Nп>�����X�Ŀ�2�AIca�Fq���L�Q����)��UaN�(��i�8ⴟ���QR��{��E���W<��NSu���['n�}���[�-���t��.4s��}R�����/���$��R��Ou#۟�	���RG)f]� �Oϖ|��&4�aL�����*jS�睧$���L�M2�36
������;U����ֽ�m��y�Kц M�(�z@���K*r�1�y��,��X���#�&I��4�_n4۔�F�ʉa�$�Q0�Qc� �ny�ْ��#����E>~���e�I���"G7ɺ�*��a ���gu��5��4Vz%3������Y����\�w�"$F	�����'��	C���	 �+C�(�
�S0¼��E �3�t��o�����G�e5�/�l����SJ=2�p�8L��S��)m#3V�0�՜�3١�㨝(Y�hRl6��HZGuvq,q��܏��E��Q70R�꟒�<�R�>�/�Qi���:�$�je�:T ����~��(}I�s��S�,��-��_~���&�����/�z"�h
��h%G�(�{Z���$Y�x;��l�#Xd�
Mz�>����X4p��.2�"@�y�SF_��P�g������:��hG��vzm�F�w�8�N�d�Ň�5/z�٦��|�~��4�8�|��e�Kɨ��e���S*�J7Pe]K�tZ�b�^'5�Wd��������>���0"?'�,�ؐ�^��X��>;)��"�F�v�ӃA#Wr�P�!c��A]�6
��Ⱥ.�U+o>�D�Jh)tjH��Te��D�v͝J�P��JnL��! �(��)2 	��*�	�ԐW�!ļK A�R�d��������Sm���4����Ň}<GۢE�m��X�*�0��,/$�L:P��EHQ;=�q�}�7X$(���I�B�%j	�"�lL��D�1�F�:�%a}b$d�H�X����pO�%B������N}Y�\�E�¼+�.8}�
�h���K@�:�E{s�|�G�(�`'����s;�"f~�fd��X�E�Q�G�K	���Q����'{?�.���u�H���Cs]�unk�R�Hz盁����bu̞+ N,����k��7�V�ݖ�S�)j���,��RfƧ��F�[g��$�ʋ�`y�8<>zB~��Xv�������73�;σ��ޗ"��7�D�VЋ���ف���Eu]b�`+�m����O9��(�P1�G��B���a��/�D��R�K�K�3�iF��P5IE�P}��"7!t$>�+�jL�Ȏ��T�3Bz9Up�MfwdHf�a��$g.J3�8���-���B�3�2�B�p���(j<��������� d!b9�7E�eвJ����ͬxc"��t|�xB`Խ�ث`(�[�@Y5V��/ʢ���C��.X��8�R.�~F�b�+�.eAձk~���l�҅��i�����>~HI���,�:��X��dҮT6�H��0
Cg>@���w���
��� +����j?Y����Ư,���!_����#�I������V>�������$Q	\�
�j u�`l!�����;(ڐQ�*O���v)ڏ��#���4$΀�|r���Ӏ���`b���q�����-K�3dB
�~����xvt̫$Y2�V�'u�^Ȩ�	C���i���%��~L���>e����ҧ�`B8-9z��o��	It�Q6Oc1鈶$yD�
H�pġ����~���9iL��bQ>C���'��E��oQŅ�,L�P_?sm_��~��%+����Wf����_�=��ӏ���&���i_�Ȫ��Y�F�̚���܄.yiM�(�Ӷ�⣸��Q��i�3�\�V��";S<���A���-�E�����x.�W��ҬO�%� "�l>ಏm?�MIm��8������a��셅�M#��2G� ��DJ�����`���*{��:�������C�K�=�yPT�7�:��j�/%�9}|đB�����щ�8��n5G�=���.*W �Řd��52'��l�nUo,�ڈ����4�
|=�R� ��ºA�X8<
���������S8]�)�	T�>��l&?:@��ê}��q8z�0����p���o�H�'0evA�āqi����jE1�eP�DĨ��5�������o�ὤ�>%u����0 ���)^�w}>�����W_RRҡ恴L�����>����!�o�����ݷ�&}�H���N��#2�I��l�ےR)JT��,���p&G�֍l���D&8>b0��aM	W�
 ���������Gg�_���������\�u,9B��Cc����&#�
���(�������A���&zM��Y 9���Y.���2_�zj���d����>���~����ܿ��>���ꑤM$ϋsk��qm�<A2�s�FzM�A�z ���T�?�����
���R<��$��"�o7���ϛ�iS���0Mm��U��z�@:�)m��Lj7�9/���SA�H6m���J'Z����R�T}���ʥ��O��3��]4��Ģ��MY�v"[�+w0 ��r_�B<����p��i>��SނDҟ��|�lQQD|�|5���ۃGI|��]#�p0K�VK _�T
c[:�R~(�; $~�ظ�a�Y#�c��ybS�)��$��,�5��\L,JG�(�\�O2�~�����O Qh��Ĳ�~��aaQ�� wv���d��/[c2����Y:ʒ$��u��f��c8���>���y �.�]��N��ɀ�\��O�D rUGp���8��%��2$@}�	�b�6�Ÿ ��%���Ph+j��"t�������]�<���>����{�d��?Gs�?�Q	���p]{���&�L� �s�4f��
-���=��p����69e�4<A(0l*���ȳ;�\$��B��;��<I����ѕ*$t�5?V{�`�b�|����
D�"3�J�^���>��..�+��}�
�uF���(D]��9�\���Z�?���AD=Z��q;Ĳ�B���V�̪��AD�Ɖ�1�$&���K����X���DY�(��&�) "b�a�03�jz-����"]q�!m���T�|�)��[�(�R��ǒ�6�Hj�$����XD��dF��g�_�=�`��W/i�#�tx�*�y4�R���B�)��f�gk{1�Q{�* 8�0���e���ʜ��X��e��,է��B��e)�>]�{�5�Z|������{7�)�����4���C���<�,�ȃ
w��(��I|��myV��)8#�;�oІ����``:$�������g������:�B��j���\���T�L�AvU�Qp������j�-���b���T���P��*p�����ù97�߅���]�J�L�0C$���r
��>,0k��W�)|�w][8��&���Q�2a���&�N��5+q����EĤX�P0�('bݧ�=F��/H|G|;t�p�Q�
K�<�����9�J���T ��8��(1�%b��}�p��d�G2�ӳ&8��[�������	����_���H!^�|pݲ���jit��u�E�W�c�����:ޙ||s�f���\T��	F�$����l�
V$���G���]���J sV�)��օ�r���n%�X�������ص�}�(��X���T�C�R����J�|�|��^�B��`��R��������*�q@����&�905]�����F��u{��[�=Ь���R�=ǯ�^�}��|L �E#]5��p�F���
+�$��/��p�6�px�O>&�vOE��81��9>��q����1&/�����>'1@����/oЍ�$������o�{�X�,c!�'����0b��uf�����CD��h�l�K�$돲̠��!���?��Yp��PC,��i�ح���d6��\����g��"|(����4G9��	j�hw��&��PPR�[����ԿV�y��,Us�
�������4����@�
pl36#u�����s�����!���9�9�b	�g:Á�N�h���Z����[��f=� �y�h�g*.T�ۣ����]��ۍT�6��)g��Ki=��b�M�F��3Q 5HP���  �u�x���L���爔�`���!�T�Ȟ��i8��ڌ
��(���i\�$R�(E?E��k
=��)[��QR�X�3�ń$�}���w������_�?��?����E���$ʮ��m;�\w��H�c�'/{ ��������(�0,:w��$-U�d`OD��fxD!�N=������h�3�;t�
�z� `�lQ�F�Eie�F�O"3	�e��^f�7M����E�Fc�9L�HRu�t(�8
2^e[�q��]� ��Ds�ڨ��w3�B痛8��ͩ+�'7u�p�i�:�{�(IV�L��4��D�@M����0���%?@����z�y@yk ���0!��������^rnx����"�}�*��y���!2C)�pvec��?G+��a?�$�Zδ�:Z���A[q��#=�qY�L���]4���
S"&E�,I�A�MI=tPN}wB�I�y�"���yXhw ٱ��Q��8��	q
��ZP�G��f])'_Ѿb�����Jˊ���IK���&]!&����>rޅ�L�(]C�T��$[HN3�������"����"t,҆�ܨ;����
��������'�e�����a��a���t��x�`yv
%�@-����,QEzU��w[A2&�.fR�喷
P����q�4�΍�����b��.�N.������jwh�Zk$�5��j,Q=�r��?���g�g�X�녊��/W T���]�M�8�rFF����� ���R����ğ����dː��_�O�#.�N:L��6[Pw��F�z�f�T%�o�6�-(���N��Y�&yO/
�3
S��3iT�M���E �Gf�2N���y!��d�O1������a
=WA�j4�ݔ�&�OW;yWהe�s����Ws�������
���j���lXltc�nh��frt_\Ry{ U�{'�l/��zKS:�R��(zid��� g7��I ����j$��%����D�$B�@Q+���'z� �v�'e\�(�7t2�	���@�nVPA��~�p�����g��NeK��=5o-R�N�sU�wAl�b6h0�}���b�:�M�p��fM�K[�(�S�*pv�w=��V=N��6ʅ�&b�Co�A祠*�X���6X�#N�wߗ�̀>�
�[�+=��alIK�2*'���<��)�3%:21�<�䕬2_5����'o� �a١+��\�g�9��:D��C!Q��8���� j�1	�ǽv*�ys>;n�0Π+�S%�ߡuT�N3(�I�Dw5�(�"w ����B�a$����)�冩/]
�)[y/�'�̀�X�4:����C�I�ȅ-�)w����b����lw��-��($O½!�#xV�G����9�A��D$�Pq9�������X���`�[��k����(8�+�#����c���Ƚ�&��(� R3�Ҿu[7��!k�.�%L7u�q"�] �~Kba_
��'����ˡ��̸_�~7��e����4y6�"� �毎7}����LY4w������ �/���z�|SYC�@U6���IBB4�Irh�L0�O�~��ȥ$_@Q��:0��C���J��P����qK�-=؄7�� 78�q�w"7(2�q�z�� P�M!�_�^��Sث�<(��gl�����7r��VӜ���O:d�e��ʾ�uH"/�eK��Ce]�>W��T*$u{�Uo,Lu#nt�W3�9�Q�5)l���)���׫Y��~U�X�'t �C�c����z�%�Yno���ԑ~��O��5����o�5NR�����c^uW}[P7D��c��;Vj�S0-5/m�n���}�j��R��m�QDΦ�bTv��*��d>26\�1���Ì-�	��"�D�aЭ/`5?'B.M��ſPҜ)�x�EXϠZCEI�z�����"��>c6�M�� [�˿��or�W��)E��3��4����u6���'���K��������S�V<>�a�sI&��V��JU�,/E蜳RM%7�W֦C��W/��B@������S�j=ϒ�S��s��T`���"�=��4M�@�+�G{5�H�U��@�Mw(��TE����z+������%�$wu[�
(�Em;�mj:�n�q����"��Յ�3�mצb�{����hN���z����*P���ԈQ<�T�cO��[�V5�*�+[��2�WX��6���ӳ���8�jl�d����:{{�B�~REAU�6 Z���8R��*������A�� ~`wQ����"�+����2�b�A��W_�����cTI�� %^>q䘶ud����dɧ���+��N{�(�:eA��d�ɬ�6h{9uPP�+�Jr��� nR�]J�bM�.["�:���ܩ�m����4d�s�.3��ɵ�EW����<#�����>��-��I�l�R������/=����\5�?ۉx�Yd�0�n��I�I�WzD�`+������b�2�ur�OKǗj�ʽu����( ���qJ���B������,�1�S�T�s�V�G��F�@���E%.�(
�?H�]F��������g�hP"��{�d����-�iK���Zr;Au�w���I6}f�Z�\���.��($v
��6	�����K
P��}C[�I=��m'��ල���������u9�v�8eX]��rk�yn�Z,ˮ#^���AљN���˷�&�v��v����u�_-R���(�«��]뙢��&����4�_��p񺟺���*>����^��$E�����`�R`_JX�&D�mP�"��� x-�wG�VT&���7b�oa���zYqU�m��8U)I%O/��˾�Vj�}2�5M����Kq�z�$M�y�+H�K�2Q�:H$5��h��[�Z�����Uo��+�k�)���Fm�@��G���CK���^X�%H0��T��1��� �f�����x-(�f�1��� �͟뵩�{���}Tg5U�*wMl�T��O�n���Q��� ꔃ)0y�>�[��]�N�K�����-������N٪z�b��1���y��P����^�g��H��_U��̯WǶ1�r��1
����o��'��s�ҵ2��#N�������y�	�_��~���^����1���L���ggＭ�_�d���p)�Jt��\�8`Q 0PI!Գ^�qt�	�q��>��gr7;���_j&�7��:���wQP�q�ȏw�.ft������H�ff/��3`����M板lz��&W_b�I���a��Ŷ�Ü���?�f���y���y�y����09�㝥+�2��N�/��N@��^&f��4�R#'J���T�|�R�[Q�������N뮫:��׻� ���V�ru�'�F;?5��?=�B*�dLTۥ�&m���~������g�TU=�b8��Ec(��j�ھ�Xxqu��r����������XO!%��4U����9^���c�A�iH��d�P���$�d7'ש)ی�5�APV7��T�+Ы 0��hD�N�Aag�]d��<�hT������$N�0����	��&rMEC���tǛ���@ʟ!��F����5��ޥ����zm�U���W��ߡ�a��WnP� j`5|I3N�7�2�Q�[��� ��r!U�LX�"�^���º�%!�c��jߢ��[4�R��U,��&o���z�#c�U����u���?}�'���CWY�����W�c���3��Y5�}�$��uI��g�oo�k#�������K��g�MS�t)�`���tu3�?;�[M�T}�R? t�ڤ,��j�C��.��}�GեvX 1�����jyZ=�g�Y�ŉ�*�kJ:JhKa�>�@^�A�Hu]l���m���U��F)�絈�3�k����p��s��Bx.�C���?�L1��xb!��.��8�ZQ��؃�<��U7�}cF����b/��T?�nR�k��ϩ1�^XCp����*� ږZ���z�34�Ԅ�5���إ�2B�{Q������}(�W1CY=nN��+�U*�ep����!�p�����Gh�IUF��Q�I���?[l
:���ň%!���4��Vn�
�*-����2g*>*V�Y�j��d%�{vӀ�dm5��{�vP� �X>2㖔}�p*c�]|�݂Η�N��h$�X�V-c�jðoK�W�j&zťK�nW;OK�ͫ��e"��bsY*B�z���\���ġ�|v����z���_��i`ks]��N�w7_�:>_� M�0�ϱ̦U]�u��m��u��(��U��\Ԓ�)�ɹ�<�ع�D����D&�Fa�a,Y�ld�e�e���[�i�^����N:����������*��?Y��0������A�:?g����R�Q�K;�P�"�܈�Yu�1t�f�ѐ.T������꒩p7)�����=�u�&��Yҫ����k8�^"2��UG����{������q��ƶ�����i�kGC�l���Ӫ������1T<c��ܞ&��e��x�YC�������$���n�4��>�By�&�ְk��i�f�qb��c��l�lY��3�R�&�g^����")��fR\�s�J��:����.���gR0��d� �@i��y��R#g�J�	b��7�m*U�(WB��<OZ�TU5�%�Si,�g���r�5徾.z��53���ô����V �H	5S�7A��բ�@��J&�R���+�jU������l�^����Ǣ����-s75��;�g�I�2�m�u��J`�E��F���Rg�a:Dh�k�VQ�� }4��z,N_@w�����dI��%�HP����rjS���D�'[�ͻ^���M|��������!U �?O%o�:[�J�R��u�طx��m�Zܚ���2�N��wi�ʉ^�������9��MYh�n�G�6��J`��zB%��0��sj���I��g��H�JHR������?�l�sկҎ�d�]JNc˄��ɽ�+ﻡ_�,@U��M=�T�{M;�{b�~J�Mc(ɢC5���6g�{w�F
o>��+������Oг��c��q�M��܌��`�e(6s �{�����0����B۶ȶ1ڗSUQ�V�!^�N�Z
#�)ex�`�����2�Ԁ�'yT��ʾr��<$�1Qv��5ZE6!07�Ռr%V��
R1������
�{m`��T@՟�I}륭�[��������K�~]Q��iJ�q���s/��~�ֻ�*����t��.��������?���0��,�y����� ���f�n� ��;��l�k���׺����F��
�m��U�u��j�d���-t����.�U��Q�{@$I�Ѯ��BhZ�(4\�k}1�_��]%0e���a�2{b]�&���<���@5^<@��wh��t���x �\��nז�-}7	X��%)�YCQ��T����һ7�H���Uf|���JNe������X��r��!V.P�Ê� q���@[� L��fկ�S����Ӷ﷨R�����x@��\ݤ,�3�c~z&�G��/Xۯm2�^�S�NΊ���<��.��{G�q�S������S1�N�~�m�:t�Jj�-�gG}���/s��;���W�h��)*��mL�0��%e�s�j�8��-��������,�S�C�("��ɕ���N͠6Pl��C�3������f8�TS�c���7Ӆ�sϦ���攋����k��|,�mt�,Ց��Ew�\�b�mc�,�H������4��m��w���(�����CR*�kRI���\��;.}K_�U��	"�r+W���Kd��*��t41/�����UXmx[��sU�eR�E�F\�)kU�5@�_��4�UQ7��.��n�������X��WQ��y����]O�7v�Y�"E�93��ۇAk�:�����zJ\� T���6h�]���[]�y]�F��R�F���������m7Q�`96V W�F�MgZ=���,���1v�c�rd�b�}�4�1��K�����K���X	U*>bv��)�_�|ޘWl�F�6�B�n�m���C�W�V�vk�N����=�U�?.�t�g��:��v���7h9�[�����jV_߰e�}p���2���?|�Hҙ���ae���ۦ�N�E���'�'�__[8���}
�J�u
�|���L�M�ɛC�Z�	P�GT�B�WG�����{�ݢެ_/P���'�s2�5Ҟ�=�ju/�i�����\G�f���d���h?k��,���8s��^O�,�kU�R$�H0����|au���͕2@�����^���ٵ:^|s�t�|�Ǹ�dWTUȸg�P5�ް8�z̗]�B�1�Y�5��4��n8��T��.���FSF��d�$ �s����{�Gw�֬����Ϟ �G+��w���ύN�X�|n��V$��8Z�"E,����<�K���R:��cRݫ�*��tNyKV�5��"��{,Jo7��5u0�؞o��ȼAf�f�TM����X�S6���B��8��E���&[�Z�߽����+	3�2�鸞T�{|�cB�U{�-�mc��8;L70ٟs���͏���
�+�l���)�����2W|>�ν�?��y� �3� L7���7`���<K� i\�[tk]������� jG!�V%n��+�1��z�	g�g���<@Aš׈��Cnit�G���T���)j �MY�[��.�;�Eɉ5�w�"�i�궝�t ���ݶ�����ˬ�	�'�e���q\���mEo��ں�(犱��s/�_ד|W{�q�e�Ʈj����]ؿL]zZvX�M�Ϙ��ֶ�w����&�x���*����2��]��rv���Ç��G�	[��,�o�q�lƌ'љBp��\/�M�5��.��*��]�]�.�X���A�t?ϫƫׯëW�MT�K��<�M1�Ta���1�%s*�̌�mb�-�e�i�k(+��Fub�<�O,���V��:vX����I.(Q��0�z:QO����:oCYI�Ju,t؟�6��vxQ��m_ұ9��� !���a�@l�V���ܹϸZL��D�(��|fkzO�Nq�HwX�qQcr�&7���R>��p����L?|�0FU+0�\�q��W���1�+�1��k���u[��[��qa�Gg�����Śi����8�2�}*�}[�_�� �Et��;��-u�*"�4�T<�-*��)�𮃵N�0X���u2�[��=]PT��_S6����\�� 8�7A!�eBy�ej�M��.�}(=�k�+����ӴF5�U\=����Gt'ϥ�x���+��5��|㪢�{kq�`�[���;�s�4�W���^w'�U�䤫�1@��`�V��,O�8�	�Ș��֟PO�<ۡ7��N}���+p����nxZ��R���/�!Ȁ*�����P�3��GrM��1X�_�YZ�b���i�Z-��`oY��ܾ{<`»�-�|x6�:{мھ�N�?�d�V]\W������Ť�Z�VL�߱�W�V=�'�j�����Lq��oϹ�r=���Cڕ����}� 0笌n ՘$�SMT+b[�X�M��j���v�ݘ�g}n)Pw�R,)��\n�T��!�rM
�U��͞��f����������|�6W��nFւp�֨���D��P�z'�ϡx+�ya���k?5�^�Њ�- �D��:�:��ĵ�Gkox�([�Uu�������_([ ׄҡ�K+W�ؐ�Ы�a�F^FJj^R�9�$b[;w���gd��U�a�n�7�8�� p���ϊ�P����ir�]�"���+��Q�:�y�H�m��)�E_�Y�� �9������j���{hK��x��V�"�x��By��o)n�{�����P��s�D�W�-�'�{f�+�	��x����k�Sʿ� 9	u}��06�c��&���^ R��d`rƞP�.n�ru�Lk�Ɩ���'�C[�JVB{��H� ������0Pݢs1#��L*�*��}&��N�Q&e�MK�����[*6��b��[�_Ltj��fC9����uW_��s�$�g�3���\����Jv��)���QyX5���ݣ4�U�P��n��r�r����@o���I�܁j���"N��ګ�_�v����E��mפ Ã����|>D�6?�Ut��̒Z����P��&��r���p7qJ74+������*`��S��R2ޒ�-:T�r���ɑCQ��M���������Wr@Z�ğ�>�v
�����y��֗\.P/�cjȇ^�j��֨��DA�Jd�Z�T������$����ؤ�A����щ�vw��5hb��To���Q-T�L����&�-�=w.��Y�h$
��:�- ����2�(����C8���{�f8��[�v(k�r,iN��������$� �;��WT����&�a��Ƽ�7q8��4l�ϸ~t����~���a2	ZQ���m�7�}ω�w~_|cs�>�vP�1�CY�z��ae�S��I�@����Ŷ�.�s������� �}k���T����b������>xW�2��lR��$i?i�++����`���#�z�GdE��!v�X����J˒q�X��j�,P�
o=���;늘J���[!C��e�~,/�Q�����\���oN�n�GLv��QbT1�����e�W��ڭ:���V�+%�^�QNq�[�hĵ3�-� ��k�{T�S@�-�
������qwU�}�5X���ƅ���P�v��+��[KahU<�^<ӥ��bT��0iͪ.�0YU5��!H��Վ��b�'���-��[��_�U���e��{�J���qQ��XH�c���+�մ�:|1' ���r��TQ��y3i�	�"՜���7���2������e=)Np�]��tѩ���z�%�K�C�WD�ڥ��y,���\O�&'�n�N1`t��X�3T*����Pg�D�9�u+l-bLU���-w�a@4�Gb��[O��"ǵi�M��(UTھU�-�7���������g�.���ݦ�1уF����5��N1k!���Zx��_B�~D6�}h�=ѹ��HS(���	��qw�9�ڞk�%^%Cu�r��0э�DJVʋ���;�"���
nn�4Z`���
�Mʪ�Q|�^����bl�oE���CS��M��|Ҭ�᥀��Z�Tk[��Z��E��� 9�]�]��Y*��}O��P7D��?�~�zВ�f�v(��|ة�a������8W@�t�2ed'Lu����j=��K�ޠ\����R���25(��T�2��&��C-�FÔ*�էBzb�o����mk��I�2�I��#d_����ϊ�V���}�53H��/<pq�{������^���+�`/��nQ�h����(`��j�Bɡj�|~�r��v����k{q��e���]��8t�h�׷+<��g�W_'��=鯣vs��m��5�m�~]M����-(H�|�����]�+w�)7
�*�V��� ],�L���8���x+�+(�{�m���U�������}w�_n��v��f����@񚦡Z��]��ޕP��n[�������P\mM��x7�w��ͬ<�^�z�1��ݘ��������ٖ�7x�m]M�ʥ��b��>ʼ��E��[�w�10�����6���Q����(W��x�͋��c�7QD�p7�.���"f�&8������נ#Hs���,ݕ^�"��r�"�������2����z'ʵ�@� ��j�[WnN俍�$�I�_A�p�D�;��]�+w�)7Tl�KC��]�+w宼�� ��J�K�Q�p��/1JXj��R��{ڳ�jxj�,�t�~f~��dr��'^��y
J���ͧ��1k�*O��$pns����#,�09c�zd�����w[�����+�Ҿ�wir:�6�2�&�4[nWyS�߬��&�I�:�����7��/1��Ų�+D���4e�lT�7�68��+�q0
 ؖ�5*ڦ�!@�s�O�u�.|^�Ua�CR�83�������ҹ�;�+�������~�ٙ��n�T�N�:M�A3��)����k��I�'I�^��(R���k� �%e;$~�&R�}�m�ٌ���L��M�+B�[)��&�����:7�Q��)ny��5|�\��k��N7L�1��J$U�sћ�Ɩ%���gܖyr�:�9E�Q.íb_�;]��[T�?Wt#ȫ.=:I�޿R�w1�U����=�nv�@mD��.� 0�ģ����=-��swD��0�d�Nt]�pc}v�]_��������h�E�e(ٞl�͐�Yg��)��u}�m�j���c��>sǝ�.����X�`��޿���@��ǀWTV�� Ce��&��oy��e�4��)�*��I���ӡ]���+�zJC�+��ݏo3Y}� ���	魘o� S˧fv��|w�v�x#��	�`8W`�M������:�!I��[�e�2Ӊ����Y3����ci�Y��3��Ԥ��:H���R;� �쀶�;���x<l��E���-`�R��z��F�
��W@	��U��C�v�i������pn�׾�۾��ޅ����~�Y�*��]��]�ߕw��B?���{r~�Q6�t�Xu���o ��]_o��0��{����+�Z��̻�Eu���� L�w��o����`�r+ u"v�A���1��R�������{��u�9����Tu����<������jEKk��1� f�;����'�=�u���8�?�����Qj��T�TU�G�u2��� �=;+n#f�u�׳�1��:�7)�A7�~pMni�܅�%61�%}�1$��:�@$O�~�}Ռ��[?u�R�T��Ck�D&���H-�-1Z�YΟ�{��'N�~]���%V߫��7)ǠA>%A
����pq��F��Ň��H�B�Z�dǉ��43L&�՘Uu~�èC䙤�a�g���x5U��lذ�� ��乽�t۳��y��2��7߭��_�i���Y��n9�in��$���L��\x�do�<y���75'x�摛o�)��涕@��ܢ"c(�������]9�D�);�%���8�(�X�P�>�N��"�s+]����O{�ls��ˀ�uu�m��g���s��2� _��v;��)9�.��ͩ�?w�ui�ׅ�%��
)h��k-7�5��l�`�����%*�Tn�2�]�� ��Md��vn+pW��;^T��TM�قjU��S�W��[v�L�`�r�ϋ�ܱ~�]<մ�Pv��������������c���(�S�O���,'�$R�>B*ʋ(��ZG�_q��i����(�NW��+-�k>Zi��]�ۇ�7�6���D�\�~�j}/�S�wc�@�/'9=lt��ѣh�j���ݜ��[��I���M5kg�L׳�Pn�j�T?-j�JUդ8(.���˟�Q�g[�������{�=e�2�S��>UZ��?�T&vI�7QnP�n's���3�����'S���K-H��tA��_�3{G�xѽ�t��{[�/�j�X��^��z��� �0�9��Jt־-nȍ(б���b�����jە���MG?���Bxʜך�
���.��V���ηuYx�c	N��P|#�j���8����9�ҭݽ��TW�z�ө��3�X ���V�8��� x�+��]ٯ��D���PQ�hcaf��T��ސV�Oow�{�^.Ƿs�C��P�����A��u�R�k:+�+�X�4���u�M-�u���k�����*Ó��g�.&4���*�Ҟ �v�u����~�X��]T��$25�_��n�y"�Ξn[o�&�+�w(������MJ��,�h� �3>i���E�s�gkr�+ԏܘc�/CB�,�����S�z���B3U�T>���4J������Ӽ>U��.;��RA�;�%���\�-�nۼ�Vf�8�Ք�XnϠ��'�;;jT�7褪Mc�X���F�}��#鰙�nc���tK�Tm5��b�mϝ2ʭ�;�$7�2��3G)ʜ�#gk+t��ԯg�*��-��og�Ҏ����{��ԅ��P������z�����T�)�߮R��= Z��Ǌ��K;*z�Ns����m��E����b���>ZR{ǽ��%Ӽ��jS��F�]�+��h8xl�li�]�ݛ�7f�ߗ��^&���ܕw�ش�8O�!$X�٣�y�ʍ2T�-�z�:����]��2SОR��~n6n�Ӳ����=���F_p];�\E��H)V�֢B��v-+oѹ�:SY���y~y[��]��e�H�g�ںe�ؘ �jڗ?����鷱�\�T��R�#�k�� J+�h9�^2��z���}��b cx�x�-���&��������kc��wP�r	���:z���>��+�p���z��L_��r�<2��F�"��*�񵽊���w��-������1����s���N���49��,7�i�ȯ�c�mn�rWޡ��fu�>f�9�[�wuF�z?�x�%�ܕ�r酁0�l���E�m ���P˞Q��\(e���v5�]}��7�Q��A;�%��[����?rg��'�)Hmt�>Kȴ���S�(���|�þc��w]��W�X�!@-�GK�-��=P,�h�T�/��֯�3�5' �c9��6%?����{�������ɌRɫ��M�;��C1ٟ���;�iݺ�!�^A5���x�0w���=�?;nѳ{�s�� �;�t,�˯+�]��f���'�䯩Q�J6��&m���t��,��Ǵ�9����]hh�\��I���<�C�����8���d��~c~���
��c�1p�n�i����W�E��m�U���TjD$I�Sѵ�j1�M��p9�����߬��9��S�	]���3z}[&ʎ�U�֒ɴ	6Y,)L���<��#,�m�`��&Cl��&&&�X	�L�,2�W�v�&�$��ԩ���E0��ﴽ��iU���ru�Q�?;4���~��4qB���<�K���v�v.uύ��Y�5A���DG�����Q}b-%#U(=u��L`����{��V���U�M�~��Vv������b.�3 �c\�q�`�)m��jB�PrL�N�5���YX��	K���TB'Nr�bS�󧓱:/�pQ�j���X����A���?��͢[j�|���1R������b�֙��b9o��&����X-*ժF~s�?�=�_���=ԭW�	��wC��ۿh
�R��p�W{&�
�&�������AT ���>��+����vb�����=������}7�~Uiب��HG�゛�ᛞ�V�Fcl����IiD����N5�J�lb�sw-����(�>�
Xv��`��2����ɓB����^��D�}��tM���wy���XU�+*�T~��/�1�|�hUw�lB����}^S������p,��xWq\؍���W�8��CV�\'��ݜ_�(e��Q���+��{\�����{��u�wPM���	5��!U���ͨ�����f)���M�;�����δ����WWby�"ѩX�vi3�kI��5(�t����:ѳ[�ՖB�k���ם-k�lpAQ]o[�j!��/��yw�~�}'O�,����j
?�&Ų�dѓ;pRj��V�S�cAN����x�@}��4��54�Tvg�7��>7ޓm:�U�	��f�VZ5P%f��u��3���;��MF'�� �J�k���c|Y�gXR��_��2��N�n)��8�w.��WW�9CKꔼ��y��$d@:�o��m�a�u��Ȗ�i��S�o�T��|��2p��J!K��W����;�j��R��{Ů	�)��b�Ϟ;�4F̡�q:�+W/e|]�#MQ4T�b�0t�f�
4�Ӵ���0<��̴�2K���g��Rέ�	��

Oi^[G,N�[�Q"�Y/�=�nִu��;�{��|���"�du���Un1�B������J]m��Y�	[@��;�V<9�RGo��A�����G434���b]�(���S��2��"�'Rs�K=9[z�O9��F�M��$UgGj��M�s�O�>wǠ���TD~y�y�i�Fb4bj��ɫ���j'��c��5�*�ރcs�ͩ8Ħ?[����H̶�[eH�E��+�4������X�ߜm��/ħR-n���Ks�
4�g�|t�<�Zo8��Dă}˖PR9�����_
f�jݦ�]���u��"��o��M���~�|N����I��9�W�1�
�z!�d�T~Ӿ�w���'7vk�]�s>2Fӕ��d���������e�i@E�SvZ��#?m��9��%�z�5�I����^.��v�D�nA��2��)�Z�4�2|��O�U��xl���==�������|�)K��s�wܷ\4N:}�݁�{˹�[�ں&�][�"P3a[T��+C�qK�8:Q_�Z�U��T%C�T�{>��܆������i���޷�����ԎT82S���ܤM�,�v�)�c}ʶ�J63�b����DA2� o��kw�{�Wi�W��;��Q_��.�����p��u���&��o:��$c�`˶�߅�:��H��R�_�g{M�P5�7X�WCy�h����++���������ڗ�B�>�Ԛҫ�9)Ճ4��
;)a�[K�9-�����s�X����X���P������y���>"�~J�b���Y�S����D�>c��?�'�cX��-�ڂ�k:��qP�J;�o����;�I�_ԩ���dMNMAYaꂣ����m�+�H&zNy�S)����,�#(l��g�w��Sׁ����jkj0�6N'-R^�8�ά���鵠Xn\f��X;t�kI��`�w�	�{�*�Z|���J��#��?��^���S�0P�UX�g8E�6�]�@W[��umݻh;��R�5��4w>e��*�LMS_Ljc"���$0����}�b��)��P�s����I�X�aZ���@U�L�g��A����9F=>H��''H�?qp�9��,]s�.�k��Ğ���cE�0��k 6�xu��4@�չeڇ��,5U��O[�V�,��S>��ɽ},MF�Q�a�o\�zO��~�g��AW�+�f������[����������7/[�c�ڞC�����eM�)6�b�b��k�N�µ��W��+1
P$�h*�^O��
tS��:V8�~�+9]�������x�>�2C�yÍժ�w�r��n�g�i
ݦ�caپ�^a���+Gpz�V���u�xw���P���j�z�ĸE,��Ȏ��gZ��VSd)Z[XWm�N�
�E'�c��?{o��ȍ,�U$���}�3������9�x���RK"Y����H�(���{��e�%q-�Dfdd�-YaK�.C����?Y	������7��A��=rG�ۭO���dgT�ٻ�]���>�6�ǂ�����^P��',�����"uX����"���mϿ��B>��n.����G���(o~F����G�w��Em���8m�q�A�'ݚ���'>��6��uD��(��.�ޣ�����Qny�Π6�D��x����v7B��Φ��3�o{��Wo6�N������nyݟy�0ѡWz�}7�U�筧(�ǧ{�mP���.���Q���������蟂�E����o�L��/z	~h �?�f�����8�4-��L��YC~�j̉�)�o���O��#��#������j"�{[4|��������'Nؽ�LSj�tYB�>k`�ˏj�WF�fV�{U.¸����p����Y��6cz�|���g�HޞҡF��_|�������O��۠�rf�o�HR�u�{zx�b�R����R�����|���ڧ��I���U�����xysC�|�aTrG��=��֤T�J_zz�{�)i��ԃ#8��;oN���ۼ�����3��&ͷ>��W�}����:/s�A�n1��X�RnY��w,�]�)���/º�x���nE6T����#��Sm!��g��cڛ����~�mP��7����l��+=�o���ɞ6��sn?���5�Վ8۟Z9xM����ݎ۽ѻC��n4��w<��mQS������E�����z/�b䛶#�>;d�F"�|m�_v��-��mJO�Y��C]�Ӽ�o���4����R�x��V0������������];�<�c�4�K;賨�������
;�?��,���7���<��-�A<-T'n=�ÓhI�|����]砋�?��9�4��fq�F�'�9i��*��d�tP�}X��E)�������O��V����v7lr�%��w��Z֣��zCؽ�T\�~�i��~�O��������j���y�X�z\�����irU��z������OA�ǳ�zj��V�u��u� ����{꼉�����}s�� �r��'���w���h��\.��uI�w=|zi�g>�*=�缜��al�����}����~_�V�{��:ͦs��q���uH��V<����⒩N><c�·��;�<榁!è������{aTm�����R�浪X�#/[��gr�/��C<G'���"ǿʤ�5S�ˡ��ǁA�+fM��E��vœz�GL�C|�nA跘2��6�+����XpO}�4Ǯ��n�b2���s�U5�X$0���Jj>6O;;�uN�O��-b�Ms�?EdlgJ�Jᾡ�9M��r���L��0�Y�ڗ�Н�ͽ&�&u��G7$>,IC�8���`b�ٳ\�ˆw���U�[*)���m�oit�fa」��C��Q�s �����F�a�|�<�uH�sf�� >>�����\��3I	�3��3�C�"��5�w�F��6ϧ�͵B'�<��A�F��NL'Σy��N����I�?">7�i�y[/T��1�ں�������d�y�����u��)\�������E;�>�z�Ooͼ��`�IZ�MS��Q\�z�գ�T�s�x?.�����vK���2���f���uZ���8?O���|ͦ�wtt��M,��5O�z��r��f7�����9�Z�@��^A��۝�_8���ɭ�{Sg%�|��%�t�f���cs5$|�����~�Y�P�}�Ӟc���Ҷ�vuw5b����������T�F�_�b�7�}S�{�����v۴��Y�+4sx�v[��n���j4��������5Q��㺬ߓ󯾆�uM���&����e�ut�(�O3�)��� 5cO,oΒ�����P�pF퐷>���zsaLo�b��^��M;��X��'3,�"�0��q�]_]�@�ie����>���������'O�e}��{������1C?�
?�3��jpͨ��2*��txΝq�Kݮ�����IN����VG[X�]�c���wzp��F�B=��̺��n�z�yF^;�6«:n��R���k������#n�8��\�QޯE 3_�������KIO�H����|8������~Z�\�e%8(�g�^��Z�k�ƣ�T��~ S�~��g�����L��Π��g�徻ͬ��=��,꭯�(�~��pi�0�{�-�{�&��F��u�8q���3�����e���]]^՟��ɬ�06GIڐ�'�����]ox�g�}��Q}������圦�jl��6GVx�a��/F,nX�k��/�Rx��*�:4w]��~�r׽����Ӝ�G�i�C��#:�M���S������Uz��E���7�u������_|�1���X7TFm��3}_��gϞ���/�#l�0��f����߻?=�����7�C��)��}S�g3p�g�������J��8�{�1��^�����"�����	���.�f�a�]^í�-�m����y��Y��m��c������=����lI�.�T8s^����^�{���c��)�%z�o�׼��?<o�����"�����NO����sA��Ϟv�ԓ�z��I�yT�o�������F�ޫwV���fޛ{��`[�#��Q�q��;�C���?�rS�}�us&�����?��ܢH�y��MNn�`�x�����@a�^�9���+/s���6u�=>>��uʿ9��|�ͰN�{�8��^�_0�!�4z2��W�?��G�=�h�����tT7�f\��q�w#�;��T��G�z���J��P�j��U��dR�h�k�bP07�����9U��rݮ�M���������;c�L�bW��7o�1'_P���g��A��87<�NLjS��FϡNp�3qк��߻O�X��ׯiD��.L�c���rr:�B�����>��C@Ux*�R��A�W?�{�7
��Lt��2��a	�~�Ds3n������rq��\���A͋��m�(c��^?a<Y�5<���_��������F�~dn������<¦Vmf��DC�yq}}E,u���ؼ�����3����3z���jd>|H��>�s	�.���yT�+�6!���z�!�%)
tp*�λ���9�&{���_8?p�_��r��,����G�}2)V�]W�t ��g	��!τ���.�e�L4��G�E�E��ull['=qRܷ��㘼��gi8�3ī��v5��-T<�W��O?������D-���I���<#,f�	���=�^�g��^���y�4�Qz�4�y���xc
�A��pl�E-nn� �B�����;��vުr�-@�-r��]�?a�h@�����3Du���%\c�Z=S��H�K��c�+cl��}��"��:'\�g0��Z9fH��)�����A���ߧ������J'5�'��hk6�}����AR���֡"^⻢y�|��y�B�{ϧg�,?��������F�,;��f0F�m0	��4����G��b�_M���)�oFf℆G�&���ʰV�� "���z���3z	�W|�{]�|z�Ր���ӳ��,� �1>cf���Гe�8{��!�zhH쯾�����[�=����k[������z���,w]��iH���7�pۤ{# x�KUY/�L}���[?8�ǵ�GDR��v��1Q/0b�G�\DfH\SA+�S�x-j�����)Dcs��|���å{�{�;�����0C�٣��� �U�΍b�(+�X�w��Kҕ�`���m�夛�x>��|��$����N,.�^W��}���ȋ�E�`A!r�&,i/[[D�=a���!6:�WQ��KOLM�W�����G�^�����s�=�~�����o���w�v�x�~~^1��k�f���X<x?f�����z�8_���a�Ӟ�(�J�ȡ�rn^[����k�m�܎��xSb�,���r�U�ł�)�ю�a����y�������7�\}���Wn��%n;�'k��Ɂ�V�;��*
�&����������`�T�@ct����~�HXT��'�I՛���#��?������~cb�˯�L�~�m���/ҪV�\���,M��G���Ѣ�C+yäf=�y#�Uk�
�zo,}��#0����ҟ�������n8��;zV�d�a��,97T�, ,�}5~�Q1���p��ta�P��Ͽ��~��Gz20d��'f��D��;�;=�z^����� qXsQcq�p���9ɘ� �W�S|_��z8���y���(���]�tc����c�7!E���nQ�����v�M��n~������igd|�,�����hQJX�&5�1����߽P�竗�hH��㦓��ZW��7ǆ�qE"���,����wڒ�jF��.0����>���������?�����_�[�MծA�e��[�sw�9_r��0I��df�&u�1�m@�L�����??>�z�����!����em����?�dx('��Ƈ�?d�O,��߸�\Px�+3���A��J�Sx�{�f_�|�dhT�� �蠞�8���P�{����(�İ�i;��\s����ǘ^o�ـH�IV�����L�KX�ϧ�"Gn�)�H\�m�V�I��nL4�u�ɤ�jɥ��
���Ƙ��zݼ~D8ú������F#؈�b��8�� ���#�DA��a��
��>>�n�?b���_���P�;�ϗA�< �����Ϟ���;]�X�s�u�Bp�|E:v�{JT�MXc(�Vf7}ds�0�B�R�H��t�>�oY70���'��B�����D��^7��Ճ'r=��y�Ϟ>K��?�K�4$$�)Żc�Ǫ�	�"�))�$&��D���&3&0eNiQ�-/��씆��?������ﰽ2s�'\�oa�e�`�������I<Ԟ�]I8�Y��cc`�ױ8�m�Cn�s�EU�;���X���-�Y>�G~bP����
�k��$z\#�[R	�玕j6�`h 6�79��\�{]ǙI�q��-�\�$�msDX���iئ�9���?��������Y�~���
�'Qx�����������` ��c�0��x�ѯƀ1�_��(�����1��h�E��&c�W܄4x�aϛ�gPs�ᔬauY��j��`��啛F���?��s୩�^:��`�v�eZm�L������l���~����eڑ��%=�� ] L��2}^w�髯�C�]Y�9[�!����O��'O�pa� V �'N��"S"��bc���jؚ��xOL~,��u�]�p��c�k?��sR���>xh�=[�/��@Ba���]6\�8�n�-���l��h	K�����NQǛ���_Rm���w���\��!�C#K��ե,\S�<C|O<����9��y�����=����#�{g��9ܸ��u�T<Gl�q;ZYi}J����|	$�K�� !`�U� ����	�5x��&�=ǀ{�� ���=�
����1����_չ��v�y���`�F��\"�!
95�Y�A�j�$�W���Cg+o���7mش`N����j�w��?K�[vN\����zɭ�/t���8����gj-i��L\����_XU�&�,&]��W"���_~�%���)(p+P�~���:i��=�yUB!<��A�I���9���X��0��������������T���q��4�;������=�0�eK����$^���yY"m���@�-��/>oz��O���_��P;"a}�6V�/���H�����5ƍ	 �О�?�����'�j%\z����_D 0�0XJ4a��q�0Ѩ����׫����� #���"��c���rS�c�q�\�y�&��>7YQ��]x�8��:��,�M�0����?�0�-9\�)I�׿��B)��VX�&Bd���v�Yo�^��B��;Z��ciB��c���Vӆ*/�e�A9��ӖIf�I3:�D�a��_������äC������8}��W���G\�=8��K|��9aKL5�Cu���X*k��X`�d���jᅧ*B8�Ғi0���0����\��J2R��u\V^'�c�R����|%���Y9��c���m��Řk����f�Ɓ�a�L_�2j=S�$�aԨ��d%��lcv~nb8�`<���S`��/�x�^j���0Ѹ�DUK�̼��3@(���%B�hK���x�	���0�L2�7�d��ܼs�����,����py���˚+�ȖPG)clJM����ךQ�o�mx7KO������[֜B�e���h���o87��O-��Z��T�bb)��+��!��&\u����p/�5'9I���+�׳i���p�y���^�BQ�>�±pyv�6[`􌧦���98�rx-�yM�j��aW#n&�|�ᳰ�.�W#t��L!��둊�k�[c �]���?{������1X��R��P�z��D$\"X������Բ�^�Q�4�0T�����\���@&���܀(θC*6ʕ-O3�9
+�n�(Xh?]
E�����s��0ϺF���s�3�TMᵛՆ��7�'<�z�(�������z�<|`	��c'�츪_��wk1��Y���W����w���� ��2h��>=�q�lj��[^�%S�Q�����0��a�WB�I|^�߱�T>��sz3�X�Gs�&LD�j;z>%���-ѫ�^�����2���L�4��-|�����{z���
�
��}	>�}~�%'y������C%�����y�ej�m����?<ߣ_�
Y3�=��v�؁������48V����I!�M��mYŰiK����5+�.�9�4V�_~���6�'����?���*A��oA�Qhs����"��9fJ,*�+&X�cl�*�&�*#�Ǽ� St��5o�@A����^��Zu��	,'�udF�폃����ti�?���y�o��E�!�;Sy`h�9��K0�L{�l��%�܏�h�<0 ���f�'��h�@��6*����Ù�Jj����]�+BÅ-����B�P5lQ��4�[�F�I�k�[K���`��.� -�^)����ҋ�=A�A=Y7�����c��K�����K�xg�u���,���LB��~���}P����k ����㹣I)��I�KVnz�ST�6��M#U���_�A&���f2/T���6H1�v���iqf�9_&���ʩ	��Gi�{�z_��;��-����X2�W��L�������uz�t�~"�GU��^2UX^�j��k�߻���M�I5�ww��?e��s�^��&�7=[F�m3�t��Bj���� �#��0{ݺ�sX0�h�u��sd=��g"��c�h���ł�|^*����:�8��h���YE��p/�Ax���
甇jB���)xh
/-��^49�9�-���QX��q[/]�XR����?5��!c!�/b�<��QL�1��qn1��+��1�l.'�d��
ùu�*�Hlʗ�v�`��Jx���+�&�6pN�:b
�ձp� �#��!��>�u��.J��e�=J��:y� ��|||7`�j�A�w`1C5�F��&T��jt�t��/Q�!0���N���滢VY��l���S�a�-�2B�[�Zۤ��GY����%�������ѯ�a��)Iٛ��<B��ָ��]�a���w��S\ST���c6O�;1c?��<��2�T��=l���F(�K���e���k�_>'���E��G(#��c�L�ƽ)W�@n2��`���rS��U��	�uy�+�׼�Ss����^�~�P�hL똁�ilې�u&���@X��a���c�q}G)�c��'w�B��uI�`B9]��m�X�ţ�7�+6E�cD�	��P����i��c|�k
�\s\1�8V{ƣ%��:���&C��?�`,<{���L����o�1����m˓��"w�w��X��/)u��S"�yv�@�r��ۭn{ngLU�4YF[}� �D}`QXL4X{˪��S�)G؂y�?��?���;&��e�7Gkð�xpt�"���e�3�0|,QD�~��k�jE4z���ᅡeߡ����������U�:�B֏UQ��'�/G����A�_���X��JzM�+�
�`��i�'���c�����aQn$m�o|?d��A�k�Z��<|h�5��q�HO��q\��3W/Y|�p�<~�.�5�ѹS��F1��z����QB��/�(~��VfjFW�_l�ڰ����+T���Z�`LqfH<�����ƽn���Fԅ��rl|'l�=~���G��\*�.�������<�"�Շ�'��pؼh�i���4���\�9�:�ՏH���'��!��*C|ϊ__^��9�e��b'���aF�J<��x�"���?��~��Ɨ\H�Q�w��p�2�L�L=qa^�5'�UI�+����)mcL�_PU��S�w��NW��ΐ6y�Y>�d���D̗A}�8��M�ӈ��!�]ֹ��������Gt1Kss�7m��H�2DrN������(���k�4��`5X��X����dq a�����ՠ^9���̘��8X�����%S�8�}O��Ә��������㨀y��@9`�2�>��fr$��F�.�#�Ӧ��'/!�#B�65l#���2����7m�ھ���{8>�Am!K�<��)����i��f��0��'�D� ���X0J�^� 4�����Q��']p+e�-;������뀙�=۩����3�w����B��D�hU�Sv��Z	�d*Si��hl��Mň�|�4/mZ�^Snp������+�W����01�r|<�pT�	!$� KL��T��־�/?nZԤ�6]j����.��b��~V�M���X�6�����)�y�J�`,������_T�z���Ye�G�p
Ci��a�,,������ɼ�✬�t�$�%�ګ)��K���=���wf�SQ]2COm��]^V�?��F��b������3$�6���R�@�.~/aX9M�n��>�� �_r�S[��=�8B�;h��cz�;]�K)3����n�/%Z�rB֝���=x�_~�=d2���?�^���u7R��D\��Q~h��S���5�Ƴ:юhx��r
�!&�y�V������k����j1S�=��Ő`���e�װa��l�6UW/#�����<��C�u[��)ϋ����dښ����	OL�:()-��H������qN����E�gu<���D|���?2�"ã�F��o�!�FU8�q2�����%��V��/��9 ���6O.�`Cx{xp�a��r���;��h� �O�<��o���@K,��"uo���xs䚺��v��:/�y�y��VJNf��^�Zb^j�)Yٕ��{�vB�������w�I��^lCU?�i�`-P�����|ݵ�)S���TR���u����V4���Kvޘ�x���~K?��_�i��������2�����/>�q=��L��&w�����e� �X%����)�d��}2Y�������;�b�b�q;v+,�s��z����i��8ۜ1�0���x��Yҳ�=޿G��<)|=�y}�BQ,�/���%}�h;X�����(W�jK�tl��x^2�ta}x��S�j�xt��s����؇�A8�ͩ3v��P���ā�M��Dc:�1=��0�;�W̚�p{y��U���'4����6��g���%ꀝ&��_���3�sK]܁�ð�Gׇ�ދ�]� �W�e_'��[z����i�O���[:Z�9��7�x�F�b�R�//������Xˊk����a�:v�PU�{T�4U���hY�L�,�~�P.�� &: ���}CmW����S	m��e ���>�ٷ�#�+�Ŭ�L�c!~�ヅ�����3�Y`t�u�^��F��mY~?���u�rI.�`��8��9@�◟~J��h�D���s���a<��	
%H�}��W�ޙMH|6 zx��d�N�i��|$���4�s�Y*̎J�j�k�aҟ�;cu����7�'O���T,��aXׯ��уtV���l cs�vOc�IM�`ax��_�����{>_Ђ`x��l�\�7x]�U�AA�F��_�W_~���z��at�VݸhLK����RY��J���//�Q�cl�,��b�hy��y5�?�s���Ͼ�A%��R0��_�����u���dҋ���/�-*�͛���`� ��ōцJH��iQҴ�`��"yz��G� �P0���*�j/�D��5��LD���1��q.1���=�ˋ�.u~-XW���cu..�����g��չ�)���K�"p�^��̩qg�(��U���_�ǳ���:�j�w��%XЎP�����dPs`Xm)��%���Nc���<��◹a�u��ӏ�_��?� ��l��% �d���&?G�S �S��5���=�k���w���),����1h2C���������Q��S���?t1����㓓��&ݘ���2N�N��B�//_Z�Mz\�u�d����/�\���zy�0ԒS�v�yy�ka�XH/��#�|�勨Ȳ�/6�YI�n��v@m�w��M��hwu���ю��M�ߝگ�(�Q��{S�S,��W�=gB���º,������������[���ٌ�YD3��;x�e�),T8�哒j�(��yV2Өw��F�{\=kT��`��8zV�[�#V�Q9*�(`�g�����'��c�q����`a��t�<ej`ۀ�����i�	%0��ުK����,��|`,�}���3���Tm��o��|�O��*��A]Ȩ��p墏?������aЩ	L
8W�XW�����=��{ϑx��C��k��;¸����b|�՗��;*M"I�/���l�WsN�d���z~� @H�٥��k�E�� ��e�[M�,�!y���v�R���V�C\gL{��w�x*ᘺ��`E�{�����Ԝ..�K=G��f������aCٹ�H�"�C��ί���:cU3(*���e�����e�2�ڄ�}T�L��V�J6x�S���X��a�T��/�;�k)g�|,R��N{��\��Kd���vk�mЙ"ƙ��vg�Ux���#�I{@��9�����; ������ow��1=����-������T%��(D�
2�����?�Vp_�u�Q�h8�)�crҳqI4k�'!��Vn1q��hR�ĔZEC��;0+@LF�J��FWܧ�p] W� y��)�mqRE�R֘p�, ��T䵾�r����H�q,d|΃0�܄dp�`��Hz0�W=ug�$)i��M�>2�=���Vtǁ��}�{�������j���:Y>K����5ϓA='��m���Ȏo�C*S�d�3l�����j�a��1e�owaр�kO�����/`�Әl��{�����5y�H&}��~�d�����Rl������l�V�[n�k(��1$7�[BлO�k�!yEW�VX�`��9W��b*XVܠ��{��YMɩU>�-���<T�o���n�v�bn6d;�JS�߻ʸ�U{��9��{n�pō�3ϒ���V'�v���IYn�{�΄�����ghl;�����ڗe�%��ٽj��Ym<x�x^�E�1:��"�#��U/0���x�ꝷ8�"&���Ȉ�]�$����◄�KT��j�HAO<�'������Zi�=1�G��W�Q��uS���!c�1����ppt�vV��=�z����lhC=wP�gV����˦ %���Қ��d�y��C(YὍ����cc��q=|� ���צ��T^����:X��0Γ'�'*�369`�,A�a\�\�f��m����Z\��1��^Ub��vHȋުs��&<M
U:M7���
树��!(%����f,f��"���!�bP�0�����û�-� U5��p��T/31Jv�א�����ֆ�������>�ۙ�@�	�B��pD5�S)�,%�WL>�����bY���D)�1�-N&�<y�p�4fR�����B�'/��:A	�]!�ra�$Ε��J`������o\��(~��\��{��coܧ*mZ}R��Z�=V����̠a�ej��+�� ���RGM�X+�Vj�,���&��bb�WM8ƥ��"�P��8JT�y�4�̬�ܛ��2�-�:��|l�.�훈6-$�pM�|	���^�6]��1�;:���@nr��Oη.n��^�a+��&��i?9�P���+�?⣞�_f�]?��5�C�@ʆI��{���ѦҊP$�n���hשKP��:ƻ�hcƷ�zO�M��},)Ռj
#I����]���ɝ�s��{�\��^b�|�����ce��:���b��6x�����KR���?l�Z�Jo�&��ݴ��������������*���p��$����C��P��n�Ņ0��Fa= ����y蝭�b�K�`PqQ;�Z�6��F�_����yBp��Ņ�Azfz�mq$[2J����G	������FBJl
�@9�v��4N!ai�k���no��1oe�o��rx�}_����J�I�J��Ӭݢ�5��"�`�ޣcoN��fm�WW��r���7�{5��v�q�ҍ䞺�%f��� �a�
�^����ƅyڪ��xN�.�K]mN�5q��}9��!|v���;W�o/-GLחo�d[��`\?lO�[���i2�&��f��\�[<�B��*��`]=5!N�g6�h$���fٱذ�c�-I%X���CcǷp����RO$�>Z]+�0»��:Kpx���ɒ���Ơ��=�R��+l �H�� %���Fѱ4|xhX�ye���if&�S�y�̕�q�9r�s&�����ٮ�P�Ia��bs��эtP94��	�K��
0��6�60I������L��<���<-��d�K(껪~�u:�6�<G�)�З�ð�<�n�[��KS�R��<���Tb������`�D�
�L �'Cʹ�rYB��Ґ�[F-�Kһ�ǘ�QXi*ڷZ���lv��ٶ'y��{ߴl��vڼ�y��E�:>l���94���;~W�p򄌅@%���idm+��]m6iK)hE�)EX�5��iL����N��-t��ӄ8����Ƞ��n���sṺ���^��^�)çE���3���$ķM���:� �i2���B�kq���UC���Sd��1uI/n��\��o�ss]Q��R���C�sygN�U�$y�K#�Pʌǿ�	�E�!�G�3u����߱�險��%q�+Fl��N�ӡ�GԠ�!B{ݜ
�0D҇U��0^8�>��+
�lCi�X�l���)Z���؛��ϭG��i�SҧpX�Ds`X7�0������o����E��ϛ=d�Xtє�t^7��5�ud`��,�SY��Vݿ��i�G9��9,�������fY���S�-�c�zC�:�։�u�!�����P�0�T�N������}I^jx*q����d6â�A=�JL�Ͱn�qk�^�ȫ�	?�!����@#��}��.�)ş��L-uK6��^Y�%��Z7VA��ܱW��؁����'�}, P���<A�����3X�:�L�77���Ux�0N
��Z��n4����dI�ŵ���{��(���>���M��Cv�z��w�� ��J��9�Z@�:Cg ���)7�:�j�>>>�e��x�~Y��!�i}�\35����Q�[�u/X�ڼSa��ԕ&Y��qhÏ�K���G�c�D�su�~���21�r�j�Z4�P�639vmZŚ��<(
(�m.ESn��$`'�ɓ�%���{|X�T>����P�[t
?f���)�xȼw����i`�#1����E�B����|++\y�悲��u�X5j!OT۷+v���g8�І��.@�6(a�wH�EIJN��ʍ)�db�O���wjj�/�ha�7kk&�w�D&m��������~��Q��o�}���oz��q:���cz�2��c��0hC���[�"?���'�E����ƴ̗�I�GۨI��O�׫���VF:��`bq�"�r�+�=P�(54�FI֌l����Ҁ�M��Fl�J5�R&����IW�hOf(�!\M������ުA[��0��h-�I}%����_��'{���ug0�.Z�� �E�'D���1썦]�NT��]Ģ0�=[ԏ��z�C��M㺸'���y�J�H�L���>ΚcbT�T/�xfJ�!헇�!E�;:�D���1���I5�Sݵ�J�I�{�Q{
�3G߽	��.��k�.EZ�j%�T�rd3��8��?3�!��o<!��H<w��P�b0,qE��x�XX����I5�/�����M������]o�DU��=����jY)t���_���a�}C@#_ޓ�؆a��|S��$���˵���1S"�3��H���ySfD�����6Pݯ�Bn͋�"�e	3ۨ%2�"����{	b�Q��N�	��"��Mn�S��`�f�LB�/��X�Se������פG!��g��"m���N��g�,[�4u֕8�����f��*�����e}�n0�8�x��i���( ����1Jȅجl������_핹x��EY	�H�ǐ�����Ƕ�������ݞ��tDx������	�%�O��μ�$�R^PK�9=��հ\��=���(2�Me�)ݺu������X��r/W�W>�e�������'���I��"s���7a��p���n��%�0�li�5��5��_}�T�
���5��]<��'~��ֱ?�Ɏ��{_wc2db��#�=�Z���j�i�."_P��l\[�0[�O�� ���~nZ�֒m�Q�sa/U�P�4zE��'e�@v�}T�)[/�-���Pr�Z���7Y5B���'2MVr����XR�I�V]�҈���ɳ>>��k��'�;�o���� L��lp������&�Y]��K�㫵]���u,��VR�(��]�㡍l����SDtL��(�t�RyO�{�m��mc׿���ν���B��z�~9�͕e�"?���-�KC55|����rpA���B�0 |���yzZB4�������$nUc�)$qx�E_��4-�1y 8�*S#1je�#	�Z��	��<��� f���`1C�P]\ס�9�����Rj1�EKj�/�c����d�ϯX�{���$�#���(�X�U��˙[�Q%���lf�s:��YĀm�H�x(�0���^��c�W�w]��2u�ۺ1ϱ!2$wc��17�c���3ePq��DQc����Ӕ�$��n,�g����j�������0�d�f�3`Z�u��^SLi�M"1?W�b��rOW���2h`pn�%`'��sN-��Rf�I5�!,VY-_��s3�	(�F�P%Z?'�i1a���#�e`��=���ƍ*���rɼT�%cQ��[C[Ϧ��*gz��g�Aw�q��<S$2Vο�N��y�1pF��?{�%<�����EV��M7v�9p^t)�ƨ��o�ؕ�o��o�ۦ�4N�lN�L�&,<kL�c����F,Ta`���V�L,{]�K���� ����� F�c�><"I������~�S
4���$�t��x��6o���6��I�J�G;V��~S=mz�G�������{��'0�8�GT�$;)Ck��M��sPsr\�L����1��i^'͓��o>��S2Jl16�gK JD:x Cm����	\I�a~��9��0��@a�qhדE^��j�,�<g+�\0K`��w��O��(*�7�Ӿ��At ti�4*/R3X�l���H*^f��:��\ Ye����0�ĉ��H|/���jMC���HCtv�����zv֊ow�����n�WfLGL*�l��IN#� ��@m�Ou#<M�?��P����$v�s�n��+��2� F�!-O�Ce-�`F�X�'�s?���Kb�P�BH�Ey��VgR��t��xˏ�>�Is�q-J��3՜�c�Y�Gc7�9�o�6M���K<q���*��F�����J��:����.�=7��a`vL92��宛�h|���I+*�*���!]��m��7���r��N2��Aul���T�JN�a>���0�E����q���(³2X�N�)`�G���ث�(���w�Ԏ�S*�-w=��޼�KtȰj��KqzL���/�/er�� �j��h��s��8�Q5k�L�䔡��jp~�����]X`�ɯZvz.N��1-�)2�2� ӹ�뇮S�\Z�ů����LA͒7��P�4�%F8���z�_�����D�cQ»���n��9igX`�!erK���+4$�k{�LC�sx�2�9�������^�������d�g���|H6nw���CiqZf��\ul��=��T��#`�kOD*4��^��m��H�*~O��c^�fLo���Z�R8?�|Wv�G�eH]?�6!�z�IH�H^�p]nHN%�1��U���׍��I����z|8����� T&ү��U�D/Nᏼ&*C������u�.�ɳ��ؐ�wĉ����b�j����C\,�(W��ʘ����Ư �Li)�1oKB��
�S��-�-^��� 5�_��6��S���#E2
	8��ٳzo��M�����Ɣ��� c
o�����i�徘��9�0�3��skF'�;�fKˁQ�qtx����h�%C�Ҷ�q�0
����7���X�&S3y=�U4��!�h�Z�&y�s�եl��Mx �x�Ba�[�j�l���� ͞aO%6�my��'D9+��jq��Ql���~�[���/�u
�x�nu�VY7�x�NY��%����9n$�8��X��)��$�o��ۨ48d`J�[7S�%�:qP�@8<?���]m-T��Y\~���b4�b�&������C��$�[2�l�*R����5t�I")^�\�\��{�����]�veZM���.±2�w�����K���y|􂯣�
��eM��3�������C�q�V��xn�k�)��s��ޙ����LP�]�!Ef�t����4��,� �1���Z�X��||a�J/!���"���e�Mg���������"�[��h�h��������0O��0{^ +3�r�J�a�J��������ئ�k-\l�E;��c�V��m�1����T1C��-!�>��:C{X���vDN���J���E }ܽ���JZI-��J9v�ɭ�-�dFŲ�r��z�quf		'�_�t�d��/��w}'��r@�k�g���&~���3��=%�Cx^�
0�y�P������F9u���"����<� L���	����[%%�3�����<QЦ����J܏�L �J*%ON�Gn�E�e���w�X��[R�,0�P]�j�k^vNf�����x_���������fu�l����}q��X��.����qC�����
S'�n����)��IA�'қ���1zYID%�0ඳ%k�-�bٵ�ν�����8SG/&�2Ĉp}���������y����Q�G���*�K�{w%��[Mwn�4EF89:�-��Di�c&`��#��g7dj1�����u��D�UYM@2V��k��i��I���M�2�ϲO�ʳ˿��R~�!�X1��S��z庬�������k~`�}�
x���c�=O!��:��o���/��~��jV0@�nL�,�/Kh��+zV�w�FQK�F�vU�<O]r�]ѩTZ
�r�j ���Y)(6
$����!�����`<��Jt<U��Ū�>%6;���R[�!�KP��&B>+��p[��]Ɔ�_�q����،/����
QFO�aSA��cks����vЍf�͆�כ�g��&�SW̑Գ5��Y�hB���6)�i�/B�r�[ݑ��}�1�����X�Ȃ��!Ns��i�A]���D%�gϢ.������Ⱥ}��^o]�ޒ[0����R�׀C���rHyV��	����y�����5,Q��ϳJ�*�/��m�.�Q_���M�{#qǢײ�w��5�}�s��a��ӧ̔��\r�oB���F�h�^A|+)�SU���~�)Q�M���м�(E���)�<q�Y��ݚ1���N�!�n�k�K�X؎q�������yB9V:�G*vH\��	r �f�!���9H�*�X�*��b��ۀ�w�f˦��>����q�1O���� ��0�l��<٦�����i*�L��o^ɖ��V�i��e�WYuaG��vҾkcќ�T�j���p٧�|uƘL�Ą���#<���.��%�T/�R��՘��su���d�*<����ExjJ��S�����	
��e����<C�J�Q�����k�*��:��D,Յ4`X=z�.��G���yV=�Ǐ3�3�&���mh�:ˁ���˶��+�������y�nLSK�L2���Kd� ���;�G���mF��_&zp��Q��9���2|.ǥ�g5�33V��9�*�@�nOt.� -�fΐ��������sn�}'i���G�3#(V���d� ?�d^�e�EA���W$&�<�C�׎�S�/�F��H��$�o)�7<G�7K�ۢ�eLEYi����2�����Yݦ9�x��l�d(�G����>��F\�䋃��j��%�ϋZӳU�>!�h9���짦u���)���F#���R��?ϙ�3��i��`�R��R�_!Lw��)S�BtM�@#ڬ�J
ڱ�� ����z��Y���M��u�"yny�m���?�΢{@Zn�s_�SJ�~���Q�+J���I��9��O��7�;�\���.�;�tc+���0�x�57m]��L�HZJ�������ͣW�Z2E)���*%
X�z���7��+G�v)C%$��O����ĺ]=+��Q�k�@s�=�;a�|���ߛ��H��*�S���ƹ|�ﲞ�H�݋��pW�ǘ�*" X��w���d!��Ah�"c����O��g�����w/�p�����}�b�����?#ކ�ޡ�0���Ķ*Û��A�}��:�6y��L�j�3X��2�k�dF��I�Q����	r ���YuCɻ��jH�alè�__�L/�� /C��jt��:�%��(Uw����;k��"O2�-'��e.*9ԤYF!Q�8䀏z6�
���d�G��J�E�bI���Ȼ�q���Hv�?+|�j ����N'~��摧�L����)r���F\]��D�ֽ�9~Y�9��W����I��!|�N�
%�!�V�f�yl ʁ�4��V��9�JDC���+���0?����ߡ�6$À��6���'��dǎђcy+`�7�K��@ļ`�\ph@�RY���A}sv.�°���Y ����c�6�W�L��R;�]�4w�i�1yPCN���{�����嵵%��2�$Lcҽ�d %��Yy�o=����O�s�"l���pȗ/���'O��\Hr��	�/�0�ae&}��S�w�~R��C(����)�7�(m���(��N�CbF"j�ih,d���6-HB��r�s�C)ј�N��Ӏ�ؒ��n�Fq8�-�6$C��1���%_�%y]m��n.�k�x����엋�>�ב��1�^8�����JTq�8��B�x}^_W�?i.&�S����k��>}�Į{5�(aUC�k���{�X�6iܮ��$v�ZEI�w�8�T��vrM�c�������z�����AQ�a���H#�8� ���z����������}@�zAg s�G����D<広�""Z�PM�֤Ri�J"sۅ��%����X��n�%�~������~!���X��*p���t����b�2+�a	�`��UA|�ѪX֙s,Rx/��8��\]-u�(!������>wa�_��XBcb��>]�X!�&�H�}����M�`Pa��8��h�;�G��
��8�{O�`a�mYj9�wl�c#z3��g
����&������~���r4�Sh���b���őc#5U���G��v޸�ղ�}j0�0F7^)7��`N�59�Ʋ+&��:�h{O�U�mo�7������N���zf��VԘfp.c�Ę {ǆ�β�R�8>�$^�i�nPw:+�q@�3	%�p G�u��Y	;�#��54�c���c�0�;���+��J����g�fw�0'��)��hD�=��f�Qda��|!��R��U<[Y���jod?���Ը�X��ü��e�8��
1"\�7�Z��� cLP���ϡ�����ie�!���o�R�S�x�ko��	zU��N}J<n�./7��J\CjF�[iL��:�$Et���ʵ7>[;E��<9��m����{���{xX�ۼ5�#[a�a�����#F����ae-S�'�L_�U�y� �0�1��u]x%�6�P�V����']ڷ��  u�IDAT�mY�o���K^�u��k��'kkJGLy���9gr�T��}�5T�i	���J�qt�p��6��D���9%�u��}���^�5�sk�b%E^�7��6P���6a�Ѫ�����n���%07¹�gƆ����R��M0�ޱ�[4�fN�W��S�"Ӆه�\���QM�/�uh����1���(K쇭�.1�%�]9��n���1z&IAi��j'�%m�5��Ϟ-�:��[O)�a�� �	'(�����K-!a��UEȞ����m�ZOsQ�����!��E}���}��
g��h��8��QQ[ �6.����,q�-�b��rN�e5.��fD7޽u���T�䏦�N���~/�E/�=�D�����Xvp�s���3�en�����#����$W��w��6�K�!�pɧ�s3<;��MT�tU�!�;�J�u��rcqX��3��K�=��0y�ɡ�����_|�%���dl��m�mj�|��.�E+�"�tq��W�q����b〱D�j��FwS����7�>L�]!�./0D$�X9���e����y����E�1�2���T�%.z�v�����.t[�T�#�N�3ǋ��UkEl�L&I��n`�V�'N&�D!3����7�K���l�c��?f���w}��M��=�[]�S�Ғ��|�����$/f�6g.Nqf�^转��U�LadI�)������זD����=�}��w\K#��"�L����xڡ�Kd |�/b��I�S�e��|Z����CR"�������[�:���evHu�1%�=E䂤���|�����?<���_,ǵVݫ�� r�ģn�Nɓ�1��m�Cr����,lH�B�s�>x�0�d���9��}��l]�1̓������g\^���ǕS�t����H�wڊRH!rsq�X��al%���U�R54=}��&��+�a���q|2�J�qc�ia�A-|T�Ju�b�S��@�:>9J�n"0������lB��3�k�aW%?^&4R
/�	/�Q�_����
��z�-�޻������(�')q
}G&�<,�R�����'��ʦ���DWTӼ�J0,6���]�NJQ�r���v2;]�a��y|p�X�6a_vu�R����.ø�Tm�}�ҿ���T3`��W��i�u��_*P�����v����g�>K���?�����E	.B���<NW+�L$��7l��a��=8�T�o�n�g�~y��^�y96;�����pup����ztie�`%T���ܒ�����;�x.�Ga��9����kKJa~�S�>SS�����A-���q�����bg�`ebnT�w=b�������1��n���-��m�C��� �E����;f^g��'����ⲳ�ȍ <N,H�Ѡ"�c��\�C�yժ�f�l1�SiF�j��J��6&h!����"�f�W�:,�|޹-�}��7�SRk ����%�L�`�.�a�,���7o��^
�F&xx�9X=��c�릑�����og׭M�sW�&�u�9ځ���[K	.r��c�x�:�m���!q�u�8�ǖV�A*���B�~IC�D����N����~���K����O��)�c��:�U17�a�)���M��YWn���1d���ȵY�񁎥�w(`S�V/�/��y�������ŭx4�s��;wa�t�u]��sD&pV(R��M\�a���?��$j�>C���dE���+�"�]"���a���_�_,B�n���qgJC�C��ݚT�:1O�����w��ێ��� �+T���P�uU��a��*NX?�
�|Z'�#�u��ȣ#�!^\Z���ΰ]d���pY���{�
��v�j�*F���?YV꺝;�lyRcsD�`�X�ֆ��1�w�wZx����x��zh<5�w������ߨ�[7�S�J�
��P�J0���R`-?ʐǱmt�O����1U
c���z/[Eqý3�ĩ�3���+7x����EQ��0B�����y��O�)�qP��)p,
��/.:���qx�J(i|a��Qn�0<�:>�i��*���O�䚒T��@Kc�-� ���"�C��R�2�����8�t�$W����5���IT\WZ~�,�n{�zWp�3�Ɇ�=�1}��j���o�!B�ao���3ǲ���/�=�1��Ļdz��!�{w�s$�����yP\Ҥ#Mil�E�ڣB($�e��?qF&1��e�,X�y��K��X0���#�V�]�~1"�b������e���v�3WAwṡ�^݉����?���{�A�E1}㝶k�F^3^�[ꆑ�0v�?G�jI��`��^�m���gw]7�����Y�Icؔ������Z��cC�a6H��3�Ք��I"��s������7��\���O��Yy1�nm�ܼvË��#���_1����c6�$4�a���a���*9Ĕoi",�ڢ���M����GMކ'�$s�)�PV���8�@IԹ�ǃ��b�D��^��]��#uc����_||2u�����; mhQ9���$���i=���CR	�ї�_��]-���J
��<s!��.Mm��	�X�]��H�",��93Ϯ:���4��U�X�j�Ke�P���?�Y��\�^��W���W�<��D���<~��]d�'d�'f���	s�5������{�m�Į��h9GG'4R(��u=C�Y=4.px����bj���7~�iP���h*�kh{*7�QEf�}�ZD،^"�Fc��q�26���]7���S�m�S_WJ��_Uo>��9�x[�^I�������ù��ECG-$��8Ys�~�����ϿDe柕���([�36�5Bq
Qb��Z����qQn��wx���Ob�x� �@~�^�d;���W^��]M��'/����S�v���a�)T
\z7��T�.ޫtF�/>>�Z��Het�e���-+�E�W^.&/k�!��6}���ߏ�2L�Y{+k[eS�G����d�V�V�-y=�	J�P�)�V=���5���M�ަ��j��ڽ�S{�ㆷ�P	�*��;��<cѱ�o&`U1�/y�Ź�������۪�ۺt�M�jvpr���x�ɹ1�OaD�-�3��(6�.�؏S?��[��.��c�cb��e(��8��sqW^�i����3��^["Ί1�C5�q��:~9���-���B���&�w�9�Wt�!0�]�&�/����WUn5�?��on�8o\���:�	�Q����pڋ��_u-
�Z��5��Ki�R/,񈹂s|V=d�?5>6�r�.�y���+W�W4]M�C�;k������Q��g�������Ŝ���c��P�Bo�=T���Eb?����M�����-���u�H�xHF@����ڥ�^�� �y;��T�]`_X Z����K921,�����S��b�n����;7FlO1x�� ���k�}�Z3�� ���f۠�`:m��ګ$�XK=��3�ȣ&L�P@T�̅a�zc��V�Wz�&�gL��8
|�U?+_X2��T;�,�U!��bF�ߟHj�b�LM�^X(z��ۃQC�¤�y�(�m:�X���۰h�ph�}���#�CF�T���D�+��6�j��񔉬�f��䑅�
�cEDc�U��Z1N����y����\��ʐa81�p��g����M�{==�e@A�/������r8����$ab�5,Ugޠ���Ko4ǺV�%��ֳ�TO�f�����������a��s(��t_s'��_�T�¤��d��>���A�����堓m<�b!���ρ�!��n��N2�~�H��
��*\�k�k�^J�u�]qIYai&0��عOOΌ�rte���{8)�R����>�yW|=8�_�5=x&�}�  �+��^F��	ҮD�8��$�ܳ�"���[�����,���`ԇ�<N���+�q� JB�n�F� �>*����d�uLe�六ʫ�<��n0H[t6>%z-��q�Q�9&n�+������*��&�2N���sv��Zv��k��>�o0��4h�^�R�+ֶ]��T�f����ai���)X�Gy�������ֹ���]p=f��c+�H�;xg�q�_�J�dW�\���'�ކ��k�X�c-6��D�Y��9���(Rɭ]��%��>rRKD)(Y����8a�o�c9������M��8�/j��p����a<����2��/2��&㫲%��B	'7��������JI/��;�0�\�$���\��t�x�� ��z��٦���ԛ�|��hܤ�
�g�O���ɓ �t\ptL�3��P�hԖW�!���+���k��o2`��0pX'#{dm�lT����`в�H��|�`S���V<� xM�LI�G���L���!x��Gy�1������b㾌�J@@:�k�r����8F�A\�������� ���K��BO�C�ժq0a�؛�n@8L��� �J���96m�de����E�Tr�s�(�M��S��8�|F�Q?���Gi��57���\ .
�U��$[Hml�.��Z���cl�>U�)���(�_�.F^�^ҒP�^'>��oʍm��SG���Go:��;}�(��1iX9��_�~Z*]�����,%�}�w�����0�R'<���fP�DC��2�Ԍw��W�3ݸ�=�o��B����\3����zut�Mҍ���㯣y <!�d����xu��`���Ħ�Cfć���f0�X�3���3k�I�r��ex�{6�9��8�Q��Bg�)3�G�[GM��K��j�lR�Jf,�KܴM!;2ÁaӼX`��!��o�	�@7vg���筪�*},1�s&�U��ݻ�a���~@*�ސ�8�+�A�<\�%먔򨤾�,���:Ȳ���FL��%��}���:���sS��7�^|�5�����&�C�ȫ���țd�2�{���Źy'ؕ�jWQ��c�)�5��!>/�1:�z�����A�!��7��v��_"�b�&���%u{zM�a5�6�Ff�>x=V��B�y�.l�'U�jx.�t-JH�=$9!*M�����S��sO��� Bhx��:#mI�C��^{��X�	7�����y�h �l��"��&��8����
#
���{m<�����l#�s�k�V��s�5���nY�Iy9�L���z�~8ۇ{����4��ԣG�.�C�`�#��U?o�-#'O1T�`��Mk�����we�<DT��b��1|Fd��*)<O&�<$gAȋ�$�kF/U^qc6=�GaC�;�����]D#�K�]��Lt�U'#����ykj�Rx|���b=��r��Xl@yr�T�Ul:� �xhc�G(I�fi����q ����q�d��A��y�0 �,N-|�y�^�.΋2�jTO/N�㶽���e�U���(�0A�+��*����J��O!t���}�p@�v��b���q�_1� �r��".4�����l���ɱ`,�k�;�J�cu/��τ�ޅD���ܠ5�3~�)3�N���*���W݂1��u5�D���	O6��6Zh@��]H�̱�#U�-�S`{^�̏������K�E_Z6;k��������++����Ɣ���V��񑉱�|�6��}"!Ai��2e��Fc��®���{E/�(����2���m�̴T��� �}�^�*?�Wɡ��
�^LcL�H;���� �r��U^m���(�@�`9^Q�z4��DT��L���A�I>�0ٔ���)<��u��/�e*��CB"�N�X��N��S��[MY�<A��F�����x�z��y(���IJQC}�-��O�~�K
ϋʙ��DL�_�/KI6L��c��fU�0f�l!����-�xΓ���"|��q�N�0��������z�=�FFD'���w�~=_z����\�[IO^bp�J���+���^�we?��ǒ{��>����).�\ޮp�P��X�)ެq�Cv�:\Su�=���x������w2¾���K��νX���|��"�禓�J�B�{�^�'����$$����.�ub���S�
=У������svͰۍb��n\�چ��j~Ҥ�֞�� �l�/�5���M��F�ע`�����4�e`?��0���k���9�Q[�Z�j��mt\�j��H¡^=+��`ܻ��o��J׾��]�iZ��<;�r���IZ�F%��`�G �!�U�}��}�͔/8�f'X���3Hz�\[����	����902Q��F}�����ƪ$v7YR��5	�a���6�{��?>�h�}��G�C�E��8�9��ql����ϝgS骃ɠ��re�6c���<Ӣ�sN��t���������v*x �2�l��Q��Ǽݰ��[2�*���[]�B?Bj\K�<N�����U��8�9�`<���~�š�ϢoOz�`n�]�#������s����l���!&R�� Pay`�*�EF�Ԫ%|��D$��sE��;/6ەws`����ӂ�C4w�~��'aPq(䋐Pi|-��@�g"�<5"�{������Z?��0�TD�]Kq�IS{�]�O����[���p�6T������ ����I��5�n������#�}�a	6�l�j���l��v��U4_������C"��.�kx�p�{���d�����Ttk�S������1�y4aDs7�%�t`$�p��l�;Mͅ��$�=Q��Y�<iP�u�m���g�Z%O����i|D��<k���GB6�NK��&��>~yl�=5y��D���(E��a�սO��к�bs]�ˢ��e˓k/��|�#!|�kcfI&���Z�x���6�Q�H�m9��7f�� ���M�����e��>|Տκ~2����L�})p�¹R��Y��r���ν&9��%v��(�&�s`�l�|�5�G��?��e=��62��Վ��K+Jǁ���θ��'���QCS�WKe�X�����-k��Bf����EDE*���ʓ'�1�x>a$=���t���j�B{�LJFD�C筈#�d\[	��wY�ҩҭ���QnbC��D_�'��-��ʆs��sV�g��s�;t.+�@�
?Gy�����;��l��u��GP����̔܊��j���T:�������߃A݅.���~g��4�{���{�I8086d|�w�hn�;'
Ĭ���ڄ�����#���;�#'�V��G}��C^l���5}�nj�#9>-�څ#]T�|�qݤ�D�Z'�~�oe�|��S�Z��%�Gi�rg��5����8��j*�ٽUw\yr4��l�.�0���zx�!5u���UՉ��/�G��C��p㸁�#�%*�
��Ӳ^#k�q�
�By���R�5��ıɃ�nH#�`x�B�l7��Gح��e'Y�ep~�X����V:��TAR�˞O�l$��O��}�ز�~.�AF)`zԍ��7�����6A�QT4O�'���=r�,�@ˉ%x�eA�|j����]�G�(��/�md<9�ʅSt�A��ì��R�Mt�i.qpE�/��t�Ԋ26\6_�	��p!��̍$¾�c�h�}%@D�Gj�K�܈.M@�}l�iJ�����;��	t5U�w�>�l�w���%��2���Ȓg!	���&x�&D�)4L��@��1���4f�ܚ�U��Ty�p�h1T��ٻ|Nֻ����w��hdj�,�T�:X.��á��6`���$šl6Z@�oI������/5Y6��K���K�}����Q���H*Kc�����G�N�6��rj�hc�����<<_ն��)��\��D^�B9��lz��5Γ��lFr�����MyW��\F��"���"����l��ޙ�cG{��rS���>P;�
��^� �D��
��׬m�ױ�F�B)��g�+ˣK��a�ᴷ��Ey�����0���ʟ�|my�ؚwjJT4���V�?4'�ϋܺ����OƠ.��rn��v�a��[���	2+�Q�H$)�w���IT�=�4E����
�j
G�kGAv� ������@�+#������%��H�P΍��!L��:u�<��tE�W�I�HpqH��=�g�~�2�6��y� �T�Q�N�xe{m,��=������駲X?}8�~L�"4��}�!���6!n5�Ҁ����Af����"�<� ��x��a�ƩnN`U��4qC/�Lb	8]M�=�s�1>�@o)�g�z��#&q�+/ع�8����� ��zU�~��}�.��ՐD�"�PLMl�mɩ%�J@5���9i>��EMs�K�U��Y�X����E��[���Z�0=�����k�jP������B
}������I��xo��`���m�=,��2�O(;�wQ��,��I���הI�� a_���{7y7H&�'|��Ԡ���SRK�������S��<<W��8s��B�٩\�<'*�Sk��Α���z��2�c�f/%�n){����6�ka��Qac��ƚ�U�dS��ug3��5!t��5{ge�,�{�~i 5�G�K�`�-�g����q���!6�w��;�4]�mn�P����y}i�
J"RHĄB8ր���݈ԥ٠��P�0���-d�M��R��F[n
�A���^���%�K�Y`�Yy��!b��W�]�&75�F���z�V��
(
�9�0xuĒb⬃m�6��[e?j1'%���U����"�0vo�8��F��G5%_8�j�d��DZŝ��Δ�[�Aj���7׿4�S���t8��Fև�Ss<����-1���KÉ]u7р�85x�G�|���j�cKT��Z�!�������4l�2QS5��I�R��

�d.�����ў�R�l)��񺐜��Ǝw�}rу�Ҧ%�ӖL�O�XD�\'�tou��W�bE}ކƖm�W��
�pEo�Ǎ�;Xe7�u4kk�\ťڼ�ja��M��Q��Ҧ��+�&ו�̠���3�������(È���1��o~��*�6G���Ş����m�[��y,A�v�{f�ٙ���og���׸ �d�NǱ�*�N%�u�x9<���\?<8H5����#u'����|M[����l5�����\��M���_���f��iΰ[��K%�*�����$����-Vh�R�[d5��b1>�E[D}���t�j `lQ��U��ށ�KNX����S�7A��$����	:nt�--2�ޫ<����!%0�O��s�ͺ����vj�=Y���m�"�KE�D�*�P�t��L����"�O�JO;l:�^�x�3���2Y���S�e�=��̰���3C�l5� �d������^�1O����04�8ozB�����_�	���4�
�	�)S��^�X�g��"��r	���.�������8��L�(E��&	��~���k�.� �t��i�i�#����Q��I�#��M_-�O���b�$�x���r��;����
��͐Fl3�1C�VL<�.��G��{�Su�u�^"�䟶ۉK��d.S�틿4�<m���[�a��c&��t>@���x� ��	7�*���}%��>�L������w���T$WPqmJ����A��N4q�W��B0��VkQ�s(���&4��uGl���zx��Y|�2�#<O�l� d�#�BgK,&�;�w���_�C,��q��'��$��5��Z�w�I��6$�z0�iF-8Z�:u�V�v����R�*�<�&��)$�W-�⢴����⟡/����6ʋ��wyW�f�Tc�b Ǜ3vU�hnn��1E\�,�	���60����Y���cf�`w�xpB�@���g@�,0����6���B�i$�9�9�F�X�����U��ŀX����0:ɯ%*�?�E�ڸ��Q�Vd���ǈǛ-)� '�'ASv{�`ߐ$a<6��RL���$V�$�?\~�� �n�0T����}��B_;$yB�f�2%����s�����G����Z���S�j�8P4Ip^f�si��E�Kq��PƩ	�d��I�tB�kA���uŲ4öՕ��^�+�.�lau��Z�WT�u?�b�e��4Y&e՘p��~�ѧ��dV
�Z)��f�_�06���\价(a�ű��(/ �w��w�|j�f$�ۙ�z>���O�`wz�m��{p�!�'��؟������ח��r꫐�4��5EU���($�N�m�ئ����xN�ĪVg�t��_�f�z�sp�j-v�M�4��m"*�9�'���*��D��I&�Qo����aoyd},�^�$�	�u��U(�[��ȁ^V���,r>17l'�탅<�)���dWg���!�lHWX��" ����z���+홹pNw�i�&� .k��.�Ƀ�D�710hX>�f��,�bA?]�lS ˏmS-&��r�,5Nx	Ls���X��E8��)�g�4mgLJ�eV^h5{��.0��>:$LU����Pw�1�����g��m����-v�HhF��f�O��ʂ�p[.g���qr��U_I����w����ձX� �(7�:���+��鴖-üh4b�,���(�^����V3J��dŗk��&b��!��kFYiuw:/���!�狏�k0H�ML�<(���<N�J�A}�����!.c�4��Q������Y�̖_q9*>�ePUr�f�A*����[x�x���G:�/����4`��<�%6��[�+�j�_�9��ߏ-���_��	 �-����~
0C�A���f�A�d���WSrϛ�K+���T1����)�H�{`�m�qCvn\��Vo�yŞp�D��y��b���I�=� � Y��]l��{a=�HH$���S�1��b k���mk)X9��E=���e�l�t�2���H��Tӿ2C��R�䯲 &bd�v�ߜ�U���`��dÃ�}#�;�*���2�������T͢�P�ֹ.ѕLx�Jn�|f���3C��j����P:��M֬�l�j%�ݎmEe��ƕKٷ=�ῩF�Ӽ�dos�[8����])�v;�����
������d���aAd��R�x���j�?Ҟc_����v�S��k�ò����Q�7�Ef��4|;�0��n{sW��_""��@L�ӛ����tp��f���n����B?\��k�.,�Am5�`!Z�h7�N� �M�cv�Ϝ�_N߳7\�t3Gxopq�j"���?���|J 
�9�da>1�݂�L����I�+�(�������e!�ǌu�u����},�N<A^44c+цYO���̓�wF�ب·�TG�o�����]SI=�uⓖ�2T�7�ek	r�i!O_hb>�� �N3P�}�O�V�ک��^���֎+� z��;X+��XgƁ�g��ǝ��2Ў{�f�zZ������bQWs}���<������<�����]ξm�ǘ"jLV���#Dz�F����#��:Yw�+�J�3�(��{
0�M�wh���[Ш��K%�)�FM���x`��	�k�d���|��1ѳ�f�yuc'/*��斂Q��ٓ� �*�Θ�ϛ:T"9zg�LB0'�c�`=�
0U/��X��S u�q�Ԩz0c������LY�T�~ɥ-梧��)���B�u1$K9������Yvp����c%�p���?k�\�@�^�=W0�4�a�uߛN;���q�F���*��` ���A���� � �b��P5`:��� u�8�<^�Ytu�wd��"�ۻ'6��[SQ`{�$m2�N������?����H�uc����3��Z�8?�^U��ș��Cz1��J�9Rq�Z��@�KE���OF���X�m&���F��&$�O�Ќ���I)��q��Y!#�4����?������Xʿ�X=F�e�ǰY�_/َ�7V�"�[��Tc��j��B��/O/� `˔\�N��'@��\�ĝ,,&Yp;����� �ܗ�!�dĢ:Sݧo�{M�.�%�Cd0��+�-���z�<f�>���s[�!��������v�E)��\�
d^��MR�2?v[$ql��9��-�U G>'Յ��8�H� ,�;�+�۽��ǀ��X`ޝ�4R]��Ì���Wb�U�W��ˍ�{D%�]�ٮ�^U�̀}#ޡ)	.d{3�E��ߕD\}��ʰ���XT��CC�� ��6$L>^Lwf'B�j;�f	/��Sr+�􀾡d�5�Y�}��o/ [r���b �Ҧ���٬��n�NY����� m��r���O���NxY>Gb1$�!&���֗:�l��>�YƇ�j'ڛx/?�d���Jemx� J��jL�8�U���SjRzU���qvk�` �'���\�)j0���}ɍ-�Gs&�C7Y�;�Q�jD��&3�pY�Z̚����z�Rk�};CĤAO̐7�@����\f�}y�]2/�1 ;dД���;E�*��!�o6�w^����[��ۙJ 9j0�Ơv0��U�AU�"3�y ؘAI����OLNҒ����r�� ��U6km�j#�d�8�p� n�д��gQ�GT��;��x�Ru	0�9��{���ns�]��[�� \5c��߹�~�O�((b�`�������[�f�m�yF��l���q��&Te 0�Pe���:�ج�{�7� �+�E�Ɖ�$�E�3>��O��-����E�2������W#�S���Źjz�7�$�A�<yP
�c���G�L�*M՚�f�����(��l��{G�"F4g�co���{���@դ�.��Yx��G��!�#".�ȑ�ESj!�U�5�9�-��{g��nj��`�$��?��z�0܏��֊�W**sb��|���at9X��(� ��4||1���'GE_�&��o�}�x
 |�����v�c/����]݉Z��n3V�0�	Y/
0�l\9�b�˗3O"���Y�������,��1���A�j����;��۱�\tʗK�LX
q�nfl,�Rku�kf���!�����,b��H�4E�K�Np�E6@���kr\��4.�՘�.ތE��"n5�����Q�P�JͣI�^X벘���b�u�`�����dg9�_^^�\�9��lC%O���A����r��l���� �(޶��$�C�Ӎ�a�>rY�o��n��b�������G���_�A����Y��,��6�������<}�I���/s���uz�W�[�C{�6G�u�(�ኄ�} u����}��X\�b۞�o��>�/�Z޻�U���!����֣�>3S�/H
��d��!UY�T��0 <e���\U1Jw:�b������1TŻ� ��F�s�U.n�!?U�d�)k�P@UPL��|{��n*��\%p�2�_� "�.rA����{����y���xX��E�X�-Vhe�oY'��� e����5?�!�������K��YE6kwnD�½�Ō����n9u�ɡm�30��0;��ڒA/����޴�8�G�-dU�]�|o&~.P�^H��96K� �c� �X\c�z���v	��׿|+��#�+2Q��D�W�Оm��m�����%��Aj��ҕKikqN�[\�]�P�خm`����Ь�{��%[������s��\$���"6��:!|��:��Ӏ�1u��S��-��S�D��~��T�ln1�?�͍ ��X��z�zU!�=�?�Y+�L�8�t��ۊ̮RpO��A�M��~�a@w��e��l��T�)�E����L�mh�W"�����E�c�ڤX;���,�����=�=
��L˶[Rk��G�j�A@`	�<�np@�d;Ih]���Z�%nnֱZꔬ_Ƴ��.b�]"rT#�oF�2~� �h9�+��{�?�3�ܠ��x�Hc�FB�ga����O�c����P-5��;�Fױ�������+����|eU�X�vB���uj)�E�r,f��I�8�\$LB�\�<�A�M19�Ų��)��O0L�HE�7�K�����%����p��dx������,��"�[n
�=X5Z���S����08�0��ѩ��y;z?��ҚwFk��Z�=L�]$�+cq����V�2��Mnu�ķT�=E�W�q�l���	����,d�ns�B:���,/�b�7K}x{q���&˶ ��ٸ�{t.YLw�ܰ��VS~����Le�����4�q)���c��j��'t�#�/�\�X��"��5D��WT|:a�$ˆI��,��M����H��u��xb1��*��ѦΡ�k��!�*���~���(�Z��s��RLu�wBJ	�1]��bC���ښ�0���������Y�;Á՚��iP�|���z�$m�c�{>R'��!��<{;��8]T�+������9�����{>�fXDE����u6�'��kI-���0(��i�S	�㩽�U}� �"\�bA_#��T%D����l�n6��  5�Ֆ\�?g)}X�u�Cm%D2���?�9"-5�=����
�����~���:Se� �)ta��x �gS���u�\�XFVæ���B<���{ ʒo4F�l���}D[��9����4�Ё�:�>`(:=jjk5�7E~>��a��^w?��n��Ȇ7��G�E��'�KIQ���b2�B��K���j��������E-�UE͂�(k5���	S���,�|C#���k�[y�(�i�L��]�$'������ܠ�~�$�������L����J��FU����Ã������5U��E,C>"u�i�%�SҠYJ�*0 S�u'2�֖N�Vl���(L4��Fjb�<N���Μ޹�}%r���Z���
FԠ]�1ս�0��,L�J⃤�������Y�>�n|H���U4����QWx��D��0P�� 2��?_�S���dY�K�%�g��-ʐ�MV�����5��`6� �s_���>@97 �~�h`�D���F���|*��]��' bZ�k�\�UR�o�����T�!:�y�6�AaclQ0�{O�oY��k6q�uFi��l��҉f���f��}�d�P[X��.X�eҁݒ���sd���х�K"Y0Q�g�]R�o�>m'���9ϓ3�QW�~�{ �s����Ѭ= �8��� �v|��%�1�<��aq�p����7�L�t�19��ۛ.��[���^;���h{��'l�Hf�Ѝ��:oU+G<ߒ���[���iM"�Xͬ�Z`�
i->bh���s����Jk u��nY�O�~1&I��K�@ߝkϷ)�_$�$t?%��'U�X��7�hFGܓ8�WK�+���j�"I������ox��v�z/-�d�V��H�̥~v�p[��+��,3�	:�������*��n��Mk	R�����O+���*K��F������A�Eފ�!h��'�T�ݴ�JL��.?�H��}T[�mR��OX��O�h ?�k��6
���H"g3v9�zZ�ɷ� � ��H�m�O0b׹NC�F���G:ïQ~m@-ɲ�_�{J1�Q���E�K��)Y(=���	T�[��DΨ�8Y�J�%�ݫ[;]'�wH	�����D��H;w �����jz-(1(X�MyVIe:�	ѩ ����ڔ�۹����X.��M����z<Y*�[�TO�Vr�_�����%��t��7H'�9Ö T����ƣuu�͢��	*��g	� AAn�&�P�v�K��q:��p�d�LAO�C��5?�7�,8|EїJ.�(Ā(]]���jv��v� L��J�n��J6���!�l��r�%��ݕ�H����'>����T�LJ�Cg,v�u�U]�jS].�������Ez臷����r��/*G{���R �!���A~��4NN�0��Jf��u��&��ug=��>u��;�j�=/������x��~T�Z�F��*˞ ˿nȡuQvUM��N� ���E����y]��z�͇g�g��9�Cc_���v��B���9WG�b�u�o���6���V��q�V��̫��3CGF�CG�Dׅɐ@�E#��
����6Ɏ��Mѿ�΂b���"a��D���F���S7z�`��}[<$�Tl�Q��ѿ����db��rdv�M]�{(�T����32#�7)0�$0�,��%��fJ�Ek��U%�N�ۦ�[s2�$!��#�����ܧ|m�V���ΟΏ��-�UUOhc08,�`��X(�C?� Ms�=�/���^��.��p%�	م,�;r��H�@0,��wb��t�C˗1�\e�J7��Y��̙���8x�]�m~Q6�� �ј؊VF'�NW�i��e:�8t�`S� �Ha�K��l���fu�h�'=�#g�(T�z�Ƒ`��Y(	�~,��Z��~\|G�X�l1ӻ����ġPo��s���p1�)��h�]J_�ģ�y[�wO�[�]��~�v���q����4//n�K�,�M��DxE�`�غ>���!	��J�w!ڣ�"������>�ʑ#*Y��S�q��BH�6�;��
0�\m�^�1x� GJ�3��T��;o��=t9���Y��0��~�gK���k��lT��w�铦�������x�Yc�$���sعC�l�z}{����QZ�L�r ���ە��|J������{tK(صAFn��h�'s���I(MVʉ�,��n>�tSn�>E�@ީ��|�q@������l�l����4@�j���*���uꟗc�V3r�͖׷���[�-�H�"��@GNb4�\0X u����nLxPk��ml).�����;�g1�bǔ/�:�d:غ���#�g"�RH��ޮDp��r��^�_�%IcA$J~����3�5��0mgNn�&b"�TF5@V::���Z���k��Klf���܀d" E�d�3ؔ0I�Z�@`wΏ�����,�� �(1��!���F�spI�:!J���<y�XOA�D��^��ܗ�oW\2�������_:���3�,�5����:T�'<�l�!@�h����DrV�D�?c��o��ژiX��u�b�����J���/���ڴ�#qp��K>to`q�y,z��ګ�J�F�T�
߁)��By��/.��)�`����Z��Y��E���F� )��[��|�&;3M�&��� 0�\��Vb���ٳ8-�gjq ]lv�>�,i f�@i�A��"��a?�`�8���Q-�vbsVzt �[�"b=yY-������2� ��1K�\��s��fR�&�[d���ϮtOxH���V����ڻ�X�~w�Q��Tk<Ìk�ހ��}k��x��
ʞ	�Tn�o���z�ӁiX�F+7��'���g��G]��d��Kr�
�h���6�eB@������( ��ʾ���In�;�j��,2[&�Llt\�T�2 I�b���τ������U���q]���q�$�T)�⦩~��ӶqS/�t����N-���.Õm=�&���c�J츗�Zԫk�[�=��U�U�J��L��P# \���v��w<6���wS��<Z�[���㯶ɯ���2��.x�y辫��0��&��`*]4���ZF�3��'w��X�ͥ�ں?Eq�?HE75X;Ia��r�]��RR��T��5?1I�fzp�S��?2ԩs֏@�.m���Ń���;��֝����7����K�2�p� .
tD���>�01�Z&��+a������y�,�ӧT�9M�l�ce��uP�C�:�1�-�M���x��C�O#�z���O/�/�X�'���
OR��!�{�n��dC������>�����͸7�e��D��^�t�c�D@�^X�C7�b���-��3t�C6�Mf�#�c 5�-���'�n��ɐl��v�*����; � ���!k`���?���*X��N���d@�	�@ߏC���').g�0�.��H�wU��W�m��i��0V�l��[p-[WF��z�G��;��'=h�������:�r_�2�/F?��z`��⭬��*>����6��^ :�� *V� �m��?���{��� ��~�V���r �N������f�j��֯�����T	Sq��i��ǧ�fF�Ty`h�;`�H�|'���=��l�f�+�$��I�ߚ�?�^*�`�@7����2<If����+k`���p/�,�ۼJ,m����,��B2$��0\������߸�>1��ET��x���u�Ym����>���||�~:Q`��SJ��:��*�f��8�Б�|7z8RH�S{&l`����ը��JA>-ub[��4�#�R����6W����e/�hX�F�3�ݱ�}�@3	4��ڦ����E�+�D!��IC���Ӝ-�Y�g(�+t���a(�n䆺3��y�I��n局�(�=mМ���Y��I`R2:2��qHqqn�t��p�U�^�k5_�Swi���8�����םc�c� ��B�p0�s���l�����������P&��`������}�ܪ���-@2�+KiQsv���}���"����liy�6��Ę�>.��~��<u��5s��T��*yE��н�������s<����(����>���Z�A*��`9u���LQ�wX8� ����8ܻ���6�su�χ�C;�/�y?���i���T7D��!���gl� �\/� ��%���'���ž�e���w
6Pm]}\�����R�P�V��ޙ���f�����big 57 V�j�w�W*��v\fVşG#q׭n�I,�`k��]���w��������>�n���K���OP���,�r,�w���$��:�)�'|Q}�6��kcx4(F%l�v���<&ƭ�x��E<�`ց�9P��t�o��,�1���5�؂�⧎]*�`q��45Dr�o)j�|�HO��±=��Ż�۬U�������/������� ���&Ȳ�@̆��$��^�dS�a������1�M��F���&���Ѓ�%�g����g��_�a$i�Yy[�Yw�����kiz��J��/��/����!�h[���P�~�n�4�ca]=���kT,��A����S�JS=i��^����a�6���y1<P��գk6�=�n嘾�O�c��Y��1mz*|vy��X�����S��w��q��s��hWg��}�&�N��I�l�b�,�m�`ѭ� ���kL�8�B�E5�83u@-q��R;�CWJj;`�Fl���F�e4ZI[�m�6|Q7�d�wݖ�+`e�l W�Z.1*cy`d~��35<�\]Xa�����t�t�W>*�H�W���
� ��嶌J�����S�<Գ���h�WH��Y}�yR��w��.(X?߻<����� b�Ev]R|<1�y6�TUI�W������:M#^-�GH������ٽ3�1��n��.���h��,�2����;�uɥl����R�>��v����X��+����ccP��eZc��F�����$3Fy���S�~���^�i ��A%N�Yi�lX�����/�J��LR�AI
��S�-�Q����y~ j�bBtr{G����f_)�����w'S>ֱL�����2�g��=6(�Y��t�+��E�Ygq[=�69�� ���<��Μ�=���q�r���xPտ�y��@�C����ѦVx�!�}��eKi��(A ���A�bT�4�q�U1��d�r���-�K����}d�\fz=�'�K��`F\"Q��Y�{��i<F�S���`0�x�� �V��\��	3�8�����G�_L�og��R�A��fU��/:��|C�X��;����+��g�|~����|D���ҩ���>�<�(uv� S\9p��Z��T�[q�Vx럄M[�m�� }�_���q�.e�䄣7�"��擘�:4cʬ�Ⱦ�=[M*��	��\��� <�[�8�d�+����yh��F�d�PԘv�=��]s~��@?�߹ �5�%z����ùd	 �믕�p������:�]l�.R�p}�(
�j��.Զ��W��鬻��K���j�0�8�eY<�3�!>�ﲲ�b�i��7 ��F�\;�/28�}�ى.�}8&�m8��C�����'V�]ǆ� ��[�+�����{܆���y������5 ���ݝ��z�.��w��R[�!�r�otc����p���@��:���J���S�_g�L@���=�?�/O��p0�e�"9r��Ψ�/�>B��8�%i��/_�@�ئ�Lq�Zҽ	��,�Jr�zO�� ��F�<�{��Lee��ރ�k�tӱ���O��>+�ɒP���6t�m�^6?�����A��ꁁ�����]rS�,7����$�,aD~�;�΃�M�Ck��Ű��k� ՘�h.'����VM�ʠ�zN	�V ��c(�QI�dK���I -Ѳ�� �ky���Do���^֟慨��v�&h~�yn|��� E�J�[z=h.k_��"?�c��kz�´�}M'W )�ں��U �����q��� cSto�_�]��� )������6����a2�(�{�\CF�e�Ӽ���GI��T��<Qf��[� �@e���G�D��o])�e�N�� &��8'7��[�3ܣ��Q��1�E'���n��&ؖ���o���ư��#���Р���6������8��n}����{���x&������V�W��P�������5�>=	ew%��9 3�9�X�O�8�-8p�(�T~3�	Z�v��wI�L� ���Ћz��=}�s�����休�n]��\c����]������Dt.*���(��yq?T_X�l�o���X{���	�s�P��ڒ���XVX�����;��r+��S�
�-��?�u���*�0n�qӎ�6�8���h͒7��`���W�6�}��X��N�6q�w�W��x~��իǎĤ��ş�Y'�@Po$�Tn�hT�\��e9�ֿ��Z9������W�=�T �ʺ`�7c��gV�:��ZW@q>����ά��ߙi�e���T��~�[%�m`|W+l�%��h�=o�t?��7 ��2��_���݁>�T�p7Β2�R�!^{�ۨ����^x �.��蛼Q��cq�����׃�{g�܍W=,��4d�����>�㻡_�����cp�yky��b�#N#
�nj:h4�3����"�ͬ�d���)}p1Z��?��4�����t���#D-߭E؄��1�Y'k��9�z��ze�x���Mn�w���΁�c`>c��e�,�˘�4�ߑ��2
�������n�\�%fhC�o\LK��96n��X��ne/\�YKW^��S�(�y���o����kW�I:6n���ȼ�4Ie�"B�i��o�ݯ�$[Pǘǣ���ÌR�)��Z�'����,±�[m�}�������Io��ߥ� ��*{���a ��Sߡ�[%�r�[�4(�5_;p�c�禜�G'6��K�Fπ�6���=r8@�3����z�ܧ������R(�p��o]o-YgO�d֧\�}��^�)v���X����2���Ѧ(�&��8Q������ƂC����~�d'���)��B_���Ѻ=�%T�J��;��]��_K_=�4З��Q��g�=�����e�!U]8w����.:$�1j�L5�#��ιN�V}g�`T� 5��`T���o�*ق�Z8?��2E�W�VcM6��PM<֋��i	l y�P�[�
�wN)�!�C�����|~q#!����!S��|��n��ǡ�����[��R�D�N'A�-�K�Y��t��M��%`-�ɟW�r�����'����j2�V����ʦ[~���rI\�����6��W���}p�2��}��/*6wZ�����%[�o��nZ\H���"���R��m*�p�l��ˍ�޺����,9��'�R�Dr�԰�g]�F����؁��5Fq�!i6���i`}�t,�z��ì�m��\�%��jL(��1�:�cI���z@}V]8�3L���#���هzܨ����
x,�B	����Qs�-,+���`e{�鿩K�%��[Oe>�$+�{���Jᜡ�Y�]G\����׈fƆ��- �u�lQJ�w�`*�.w(��r���n���D���l�����j8�'g�΂���v�*�2��~7r`d7&������h�o7��V�m���@'��X,���Z��mj[�k J%�9	X��D
w����ʕW&�y���o�";�gÚ����w��X/&�߻�
��º�@u��8-���ه�����p9�]n����	�vŷ�7z��Jo�7��a�(P$�RV�6~�}}�oIE0ia��Vb�������v9������c�ނ��(�̠�ߢhq�e�z��o��ZaL��o��9����<h��*0�r	��p?췣6�>_��T��|N��Ƨ�*�ߠ<,�~w�H(�t��Y]��
�ӿ���~���^�^U����,�3[�E��A�$�/' �x�o��(�����\�PS$O��@���鋅���^����^�<3�:�k�(B�ڱ�!
���������Q4�RZ3��������o��v�Ks�NZ%pB����z������7����@�9�+T��6/y3Z�Ae� UϺ8x��p�r?T ��{m�
@�
��=�Et%�%��u�s4�i�D��k��	dw������w[�ÿ�Fy�c�pG~#���H�^�A ���u��R�dw���m�DV��Ce�|}�!�ѩ�S�fP%	Cݑ7������F��̡�xf�6�3�R,�q��d��K�'����D�wQ�Bs��`����N~g��\����.F���~��f4dA��{f����d��b�U��8�����E�(
Ĝ����{��L���	�q}b�8�g� *�'fKS7@9d�g_����>�6'� xw����o��@�I0lX�-�'��=o���쩌g\8�%/�ݱK��k��:/�/u������s�7�,�v���1�_�"��z��#"{����M��t���H毚3�-�������)�D�<-}בE�Z�T�F@��<#�L>e��N��b>_Æ*>���rt�b ��P���jTc��վ%���: i�
�	���V���}�Oe`W�5�V���ڏl�:;�[���p�\�c�I��8�s��ˁ�ߨ�5�M/\h�O,�r��9���7�WY	>[��?�}o3���4�jn�t�;�)'DnQW���Q�s�5a�CF`|�z�$�"��~�z~&mS������c��������^@�J��΂j�|MxZb ,�&�oGө5^꬀�r<��~.�ӳ��z,-�M
o���6���>P�Ľ��D�^)4��{��X�Xg���c���{�N �m@(��b����/�ז� Բ���n
0�[sh\^I�'@=A���b�N!�$�����?55\1{=�O z��%��e�)��f�*"1����z���G�~�Y~LZ�<�ew�e���߬t	&I�:�=k+��h�����=WF�)�Qe��t��O/��so"p��j��6�L"�yw+�8Hh��߯pJݟX$��j���f	,~Ǆ���ܨ���Зφ���[%��14ꪁ�fe�ʀ�l�ŎMS�s�@5��F*)R�;:��I�l���j�U����l���ն�<Ի�Ȣ)V���-ِ�4�u�P�O)��tK��n�!m�S	*v�3����3���y���GJ)׿G-���2����P#ɇ��*�nN�آL	7,��R����Z'�ָ^=�Bqխ1 ��ԇj�SZ�?Y�16�IBL�@�&���lTU|ہ��N��CvR1��Ӈ�,z�{3������a/u�Ջy#��Ξ�L����{�
��ܕΩ��)اӵ�3uF�.���2�v�����������`*��ߨ�u��l��-��l �`;��o�l�绥���T��{��f�ԙ�BM4I��2��b��%66�����%Q�
Ñ+܋��׽�b@�/�lUe�G���{ey��^�C�A�/��yت���]_�x�+�[>�_�F���xf2�ϴ#�1�]�5eE��d�RJ�5�P��o�q�N}�	pW�$�B����L7���c�'��-�>�r��>�<��_�q����\!������t�ب�),�Gjn��tG[�5Q_q�*��F�~Q~^O��u< �+��֊����O�n���jj��U C�Ѐ�n8�-��Fq|@T�':F�������Qt��K��f��>7���%A`�n�=��<���:��x�Zj�����d	���{��˰�j]�<�R���<P��	F��}.ZW��Юu]01�eJt~�aճ]���Wv(�p.� TI}M�^/
p/�~���v�A���5�Y�u�W���u�)@9�Up��>d0e�U���X���/sC}��P��<���WZ5K^��s7�0O�r�XLL��x��Ub|^�+�?�����\u
&1��w�_%ӊ�//a�wW[�kUO�סH�����F�1a`����|�X4�=iAO�^�Q����Yr-�|Ր�fN��3בv`3�`�`}&�1��r<�9 ��P��[��m��g?�p|Б#J�|�:���N�Ux{Q(�(��u��u�ۋ�~͝Љ��=�&e�#�#��{PM�V�	�8�7��HTd`�4���sp�
�nl[��`������2t3;͏��:����8)�)Y7�Z��O��t��w���B}Dh�ߑ��u��ӕ��'/2��6��`��1��w���fO��;���������������L��:�ћ��V�5�ۃ����:t��$��(���H�Z���F����UEP"¿�j�m[�-�pϲM��X��X%�4hh�����v8��{pT�GO��\�`67����z��y�u7��C�̰�ϫ����9����ifxd�@~�?��G������g��h�s;�bn���W��	�`�<��9�z��
��i/�+�Ղ$$�Q'�q��V����
���`5���G��3��@��
^Z�f��b���N1�LS3T	��"J��-J��(�����qzf�7� ��ʹ��?����g��3��j�9٠
�ᚆ�/���U�X;aU�3��b��ts�|��g�>������V�%����ӂ�#��^ۭeu�y���j�qq*1���祡�.�N��W�b����v{fKs����z��P���o�>��|����"���s��~�Q�����h�f"ӱrǏ&�5"B�������ig��N��[���'џw���i�T쒢z�"��dw֣߳<c�t)E;����U, 5Kr��`�-^�[��?��i�
��_Ӥ��D�+[]��Ka6�i�=�wc���7�n�9���]%���=L{ ����Ҫ.�o���}q����
i@�e&��Fã��}��D�S��o����"����Ӣ�e<b�J�L=�����~~���r�N�16R���XT�Gb?�H����zx��m�났o%�;ϭ�*<���Y���c�S��3vц�A���n�� u����Yw�N"Z�sa{����P� �8�� ���6HKl��,��3�Q$����y�)������I� �MS �n�d��w[���*��Սt��u�0l����s�>���WL?�`Դ�ft9�|2�Z]d�d�ͻ��`�h��oZ�!h�JoÑ�]!JK�=�F�:��ꟾ�7��o3�
M��-å��{��2�4:�S��Uۋ|��@{x�]bI^/�W-KZp�@�؅��P�;��� m��|�-��#s@JF���L�dAW��w[����1ԁ_wl5��udB�K��B��C�v3٨��O��%L�(!��T�����m'���$+�B.��-�u*~]]��C�D�Xd˾� y=�F-�?����tC3*;��&Mx�dfg� ��pʳ��M�� v� �%��*�Jk]��u �f`ZOma���ӫ�K��ľ��kd��u��ޡ���0�u�.~ﮯ�z+�	�s�¤k�����3L��i��7�ˠ��&x/���q��l]���Ii���v��Kg���P{�=��!�]-���r�tC��h�5'j�j���7����K7Dd%&Ͷ���y��ƚ<����f/e�ǧ��<0����Id(���������t����Y�<j���_ ��<�PwU���n
U�U^Uז G�[�BΉ}1"t[�������QҔK���μY������ ���?Ix�x�=?��v�>���~m�_Q��*����Mn���%V��o��A���Od0����;���%ݥG�UkV;g3fD�ڡN�7�xZ��q�p,�)�����$)�s������J.3,O�1�څ��i�����o�\B��$��u��$ak�<��J��j'�`��� ���ȸ3"y��+��02��B��T׉�W�J�	L�!܎�2�@e�Y�ud��%=�I=Q[��75�Y�&؎�ǲ� ���K��2�b�� t�p��ʒ��j-� Ҥ�����^π�����|�+���*3{�1���m36��q�����P��������xX�~���*����gHo�z�m��B��	��G���D��6���C�������%�.۵��������x_�5�|���� ���9����*?GN5�vV!����Kj^t�g����D1I�z39<��'��/����v�ݣ������o��E�_L'J�Xl;*��Rf�^��/V��*�)n�c��	$1Q0i�>��'��cM���G�p��2���sh��:���Y�\�GK󎟹Xϝ�
�P;����Mq�� ���Ys\�ȯ#Oʈwsv�t��F&����"=Q�P����6j?QǴ�^ǭ�x��hA%���lil�z*֮��F�m�XZ��3���[��ז�2T��V�9�g�d/iF4�[�Tk[R��Y� 5?"���vA����ύ���Ϙp�� ��:Vt4f%�`Ө�� 6T�`N���.,A�՟3`�OSu0���	|m6� �Q���[\�R�:⃱�J��N,�E<k���j���q��
 ��O�U���`O�PѦl��������u�Y�k`�9b~|�$��G$����=�j�i߹n��^GT;�~,լ���3|�4���:,�Н۽O_�>������^X8���5�0ϱ)ht"УN��$0��<�<L��a�vG�<��i� �<i&��q���3��6�9�R�O.uZD��ϣ�H��]�HE5BKz��0�U���M�5�j@o������ju��^��d�����s�䅀lҵtj�̢7��$*�^k[p�Q�;	@�hZU�3�OF��Xg�O.ԏ��9~u��Sl��>�e�t�V�������.�b�������YP���w�j��� ܮ�m���4�p�
e�+���+[�Û��-���FW�<4k�X5�F���b�Xn)ПV?nج�a��{U��7�AHA����~�n��K_s0C�Dx,>OK:�(��a
J�Y �u�):������:J߲
���欄�y���a;��]��8��NV�U�g�^��bɦA\s"��}�b�Q����,-/C(��y!Ȋ?g��I5 ��O3�OE�n�BWȳ����@;Xb n�#���ق�rYR6�P��X����#;���n�
�p�H�uR_��1�6|�����ڕ�|�bl��K��K�3�>:�MR�v�@��`\ʙ��h�IZ��c~���X��&n�K��g,4���?vbTt�J�˽��3����x����hi�"��1����":�d�&�M
f�M���^q)�-�����^�<��F��:3!}���x=�30�,���B1���5��H����H��������*p ,E#Ȕ�S������(N�[�Θ[	�e>y��:Z�Y}l��S�`q��C�Y[,�k7�h%<���J*CR:;���6 �Jǚ�O�Xs_m�B���}���T[0�0LƝ�3}�E���]r�E�;��,�`�w)�Np���[�f���*f�j�;1���p$^��.�7�ҥ���~F����"�X�ॻYNPC�dlJ�B������-���߻�����]��ի�ATfs��u$����G&0�h�0�	���hI�j�v�������5h+������\���s�ݖP��kP���8��J�
z���T��f�K6\����}�1H8(o�K~�G��0t�����e,s]��w�[�k�̺��a��u���u��?M�]ө%�ȴ8�}���Oq�\���A��2F��1���K���c���>�N�>:�wX*�����_t84������¿D@��F�/N�F�4́���㖺�tQ��<�~7�Ȯ�`�HKJsbz(O]k��Ƅkq�d��J⽶T@����t:�B�5$@)�n5����[�sw�~�VH	�Ԏ{�Z��y¢�"���-�ܿ/0pŽԓC����Y�M|�S�����0i�7�#�}}�9���C�u�=e�bYdG�}��X��c�Z��c�fĚ��ñ�vY���}F�x���^�G��ӵ�9�-[\E-H ���J_�\�g�J,e�<#�;iC�Nfi�:�lR֭^�u��nr� "V/��T|�.�����:��Y��zݥc�W7���(�� �t~g�$,�}��z6Gμ��^i�wLɥ���I-�X�O�=M�=�� ��$Jͳը�nr�eۍ��6'�6���o�&��}�gW[%
V����A�����]~�U%7��q@�5��[��s?����1��u�n��|O��󌠊*�q&��B���==�Q��xoh�����㧗�]ESl��i�����kʕ���/�������R��o�n~� �����J�o�G�k�M���w�3p���U_�6匕BBe`*g��߿ ��g��"������tӧ�����(�"n����ޱ��$����������~����Ӊ|V2�:co��d��%��~��f߹���2TH��~���ݖ׳g�A�g�__�?��V�_��-�ώ���|�$�c�'��R�]'��������+������VuOK'���<��סn��.��޳!�*b�Ź���%�{�GI?�,_2��G��������{�v�^��%�2s�E�au��K/V>��K�񳗒���������xQ�	��O��9�}P{2�B�L{�b�.��><I�U��Sӹ����O\Z�X�|����Uz���| n��}M;���ձ\x����蟗Oԭ5�ry�|ß~��z�K�����Y��(�oy��L�-�w+����R~q+����. ��Ģ��qe?|�Y�������ӷ��|bmw}Ї�㱓��"������B�B��dں�+b���ָS�o����{t�<P�J��WO_�v�~�|���#�Vל�/�ț�+�%�'y�O��ϖ�ǅ�=I����+��}QG����K�'._��lbC��E9s��y�/3��,���~�|Y3}����+��V����?*���廜)�X��O���=߀�]��w�.�T���|���]>�|�w�.��|R����]��w����~�]�#Mi    IEND�B`�PK
     #{dZ��S�  S�  /   images/e5551f5a-2fb7-4493-9527-57db21faeaae.png�PNG

   IHDR   d  �   ��'  0�iCCPICC Profile  x��||eE���Vx�*�g\�$�{�R�f�IvC�]�%�lv7��l��U����E�4��)"ME��   �4AiR��=sg��E?����d�y�3��)�s$���_�`Ψj�̝�h�{���{�U�J2:�T�͒/�,\���Ց�'�~��ǒz}���J��~֝1�p I�W,��K���- �~��g?G?K�0��g9z�J�'�7q<�ݭ�S�d`���>Iƭ�?�ha��������sA/=a`ͻ����;c�I�*$�̚�x��ch̹���A��$c�\�?<+I���g�\�FЭ�m�Ϥ�%�����2���L�Ve)cͩlf���:�����y��C�4MR2M��4�1�5�kʴ\����Ӕغxx�ඝ�{Y��"��t%,I��ݒ*��,iƫĿ,1h�HZ�Ix�:��&��;�%�6I�8S�ׄQ�u ���M��{���K�<@u�ǵ�1c�%m[��&���_��^[�/X:<4k��j4m��>o��Dғ�,�6�~{��ǆ/<�����,��qA��m�b��(I�x0I־<�m��d���䶶H<os
?>Y/�*����������\�\�ܖ<�<���|аJ���a׆}�5��pm�C��Z}T6jڨCF]6�ѕ�;���ţ�����1��yb�cg��b�?��qG�{`�F����J��x��V�b���X�UN���ʌU��j�w�ֲ�-��կZc�5�Zs�5���'k��k/[g�:����7�׽�+����p�m�y�6Zg��7�k�1�\���6���͏��~1��m��~�u�J~��[l��V�m}�6�}y�/���EM��w��W{�+I�ͮc����r��[O7]v�v]_����w�񀝎���-�M����I��y��[���>���w���η�n�պ���K{��6a��ݯ�c�^S�q�7���侳�~c��N���L6����۸�����l��O����[,9���.?x�e�|w�CN>l��O=r���>z�1W�k�=z�~'�;�SZO}��#N��ߞ5����\r^������{~��ŏ_z��G^���Z��p�'�=u�/n��/�~�˭�ܾ�����;���{ο��yp���,�����ɦ�����y~ʋ�_������ޘ��No�w�����?���-�D�X���3�0
�]�ɇ�׍�`�a��='���W�4n�q7���Ru��W��r�*Ǯz�j��~��׼`��׾}����z����kn��F;l��&�7=u��o~����K_�дE˖Ӷ����m����^�ts�ǿ�B�f�o+�5�zzc��m�n�f�o���;v����>���']�v�ΏM~i�w�>v�M:d�nS�N=������~�w�i[M�e��{�����7��+�Zѷ��[�o�ϔ��s�<`�wf3��}/���9��}h޳��\���*7^Դx�%��ׁCK�t��g,��;7}��C�=���W9�z�8j���8z�1��=��?8�ǟw��?���kO���מrթ�/������'��s�g�z�~t��G�sȹ�w�����'����-��܋g^���/���h��+߿꣟���r�:�nv�6��׷��q��7��r�慿Zv�Q��x�Y�_t�տ��o����w>����z��w���������?���{���{��?�������?v��?|��?��§�yzڟ۟��/��m�����?���^�����m�+����߫�h~m�ק�1��ҷN��eo���s�~���><��?��֏�[1Ɲ��ɿvo�a�&������/��5�ͱ���t�����J�\���%��������k���kݼ�=�<���������������	�]���'��֗�M�p��-w�j��{o��ˇn{rӏ�^��+���gϱW���ߪA�7��5�[���o��rǖ��|��-�'�z��]��o'?������Z��b�W��N]�u�n�u���Ҵ1ӷ�}�{�y�^˿q�7��?}�����o�O6�6c�`�̡Y�g9tھ�w����>5����ko��-j[����t�qK�9誃o[��w���|�f��#ڎ�����;�裎9��s��q��	w����>鹓�?�S_]��io�����=�3�?�}x��|p��}t��?^q�xQr�'?}��]�Ko����O���+�ꨟ��S�>����~q�����ȍO���/_���z��nk��r�:���7[�6�s�ߵ��{���u���ܿ�s~?�����8��=鏧>���S�8�O��?=����L�ˮ���\�����~a������}������m�^������.~��7.y󊷮���8�����{o�k�k}8���Ώg|BH�#�Q�Zä�s>����G�ї�i�_{Ӹ�ƽ=�ܕ����ʯV~�ʕ���ڙ�����k^�ֵk߶���>����_��FS6^���Mo����/nո˗fN8|�s��q���~y���]�i�扵ݿ�o�,;���/W�[�=�Q���v�n?f�uv�b'�������:鲶_����o����&����;�N���[���ݳE�iӏ���=~��s{����ߒߞ�7k�C�O�犁�g<8��̧g�0�͡O�[mΦs���8�kA����p����r������J^{ل���~���C�v��q������Ǭ{���Z��<a��8���'|ʲS����ӎ��Q�}�1gsֱ?:���9����;��������p���s�~�����K{��.?��<��~v�Ϗ���kN����~�ˮ����n����~y�����<s��r�w������ѿwW��U�Y��U�w������s����`����������cW?~�����'�}j������g��������=��#^�ދǿt������W��ο?������k���[;����}�9����]��߿�?~��_�譏��ɇ+���,/n�$����]�b�No'�Ӯ<��wW�x���a��R���k�L�R�H`�k��$[�̱j�Ks����#u�l�)y`��������%�Z�Љs���־w�N}'���ڤ��������8-I�w/3������u]�N�������x�ۿ?���x�̞l�����񊜡�!�*n�Ff�����+x�O@����D���W���������M��Fo�����/�����o��*_��'���c��㎡�m�W��#g �N��޷S��a�! �~ ���C�B��9x�-��|K�_��	�v7����x��k>�b�|�x٘.;�LaaB���}�A�U�����߭+Aֱ4�m�'�lP���T�jK�$�����o��ȍ�7"����T>ukjA>����AYƀ[ǀ�	��ݴ��P7�N7W/z� ���!�)U���a��&��u~����X�~��,w�����\Ɠ˰i�
�>w%Mu2hQ�IԞ�m2�N�Q���c���\��ȌdD��q���C�&���Az���>$d����fh�Z�'���t|
�RY�,��b��O�!�/��Mg�5��d�!e�l4�W�1���,��6n������>��m>�b��;��bNV䝽�Z�V*��zZ�ۻz�vW[�g-�3���?gh���EC��U{��g.���^T�7s������2��}r����]g-\0<�?��������6���ӿ��ٿ��L5��I��d�:Ј�������v���T'��tu���X�i�2���oR{g_Oo[�$1��ή���m{m�sZGo{c���jc��}�Í�ޖ��m�}�Szz��u�M�6���=�h�:�U'a�s��v�o��Ο3�s���B3V����wϮ6��sw[�.��)S?�-=m}��o�X����jk��n�ȻuL�Ԧ`�X\_�NVm����̘�jmMp�XZ�R[˔��4V�L��l�h߫mR_�Ծ=��4�6����X��>�mj_Ǵ޾V0L�n�m�:��kjOO�Ď6�T�؆�����胈����Lo{*�K���Ϯ6��T�[���ՁP��U[q��gTZ4;H�Ty��l�W��ͨ�'���Se����͝8�����6eR�ܕ�{ں��A2˳>�4HqbGK��B;�G��6����o����l��Z�X٥��7��x��}_�Wml���tN�ڻ������]�z�v�ֆc�6N��m�{_8a��5u
��}��V�L���݇�����1�����'�����L��[�i���pJA�������u5ɾ=ܿ{��rB�{�=m�=�L�sT2�v����Z&4�#�dk�Sa%�Z�״jT-���U5�Së�ո0�����|��OV���g�"X�E�1+MZQUvSߏՌPR`M5��Q�)SVWtU���/c5�,SUY��pK�	&S!*&J��%3�GGX8��S��ظ��~R�D&9��(-m�*��J��t,�,u�gBXj��GF+�⺒�И�?v4�yVe�k�a�c��d#T��Q�Qe5w��"�i�0��2��T^�b���Yn���2)-��M���(;��1���"���L1[5�$�}d��������יѴ���(Q�T�1�����*V(3E��A�d��8F�4V�Ɍ�c��:�d��wj܎>K@����u^� �h���F,˔��g	�	�&B2�II)�
���DZF����f������D�љ�)��ĖZwdҰ����X��L�-�z6)T�Å[�)�Q��pH���� �ɌT�&d��Y-���:S#�z��!�&�f��c��3���VO` �rͱZ�o�Z�yjmN!�0jR�z�՘4�\b��6�*�ak�����$U�,�*+p��aF�jR��	N��\#�q� �V*���he���5�2)�r#`��=PY����	I�]O��X�m	��b�ؗ�}a	Ο�贄PX2�P9U#�ġk�R�
[�X6�hN;�#�feʉ�ڹcq�O>�s��#��I����N>'��N*h��,�B=��$�!�Ԓ|)�Nji��n�c&ͬ'���(�p�b�Y��*�5o�uDF��Wd��֑��d4#����� mWp�ďȝ
Rc��0h������ؘ�QW3�0PZ���P�
���{������V0v�c���P�GW�4��)X6l�,��.�9X��
�!�
�9�[G����9~��;l�(HѺ�f�S-S�e�)!x p�
6.!j�T����(��?����g�(�����"��U���6U�TBR�
�#�g�k�C�GX�)q�>@9�(^{^G�PEi���p��A3�6��[=� �i�������a��hH��K"�:�+���疤
5�)Ed@%@�f�0�Ԃ��@�pĄ�2�+8#�j�FZF`|!Nj{���6�8Z���7VuA��BpO%N�W�)��J���F��* M(��JI��p\���mf��RZ�@�H�X�V+1�_G��Y/!��R2L�,ڈ
,E���u�$G��¬�z8;�pxX�2�����$M#,�(nY�$����q1����% �T��qdX���i�F(%�:��f@V
SK:@& {��ZJG�CiZB?&9��ٚD�68����#��B���Bt *��U-
K�YOh�m�f�U'U�ۑ�`�F�wrHaL�>��@dX*2-�aF
VO�&a���dH�Ҍt�֎��0Π��a�a�{p+`W�ϑX=��4�גpp��wX�EE���!&: u�"$\�%,��(]�5D�����ı S�c� ��)����W2�>��E$geK2��[��4�I��L�ɠD�ӒL��H~�4�L
���<p0L�_�+Dֈdڥ~��5���e{���*e����8t�đ�U4���u�b2M^�B9%��W-�=:��Q��:H�'���j*��b�����H�#+ ��'C2���U}GA����#�t�^
�uI���(B�(��(��g��z�-�'�X*2�|]8aC���
$\챾#�#<�Qsʩ0�Ó|3b��%eq UC�AHڎ�,EŔ�q�9��!�������{8VSVȉ'�����J���LX*/Q�(.8C�����<�BF�E�!GqQ���cF�f$�.Z芑%E��! ]�<���QM��|ᨒ�#� �t��
�����[�*d�xc=�g >H�E���H�tMZ,Ք�1�����Fy�&B�V1��Y��%�֨\J���nIu'�i=��u D�����Uj5:f%�@�`�P=red.��paι���� eU�:p���:��d��/�� `d��i�@x6+�XZA��?F$Y\80��2b��T���9e��UB�����P=^���c\*��8xPޒY!]� �V��Ǒ
��"�{��b��2:S��& �!�:�hH�(�� V�-q�EGAZ�H�sN
7I�V�Ҳ�S4��"'g�z
"�U�Ҭ�g\,"��J���L��|�
I�GV�Z?�MK�F�\�5�r���K|kT�T��|�����@��%�5�pF�.��\��\GU����\�l8;CU$��'\zH�=���EO���\Ru&���qFs�U���%�=����� ST=�j�EONY���*ydEU ��1Z�-�:~��6p�)%��r�YL�d���b��e������9a�Գ��{6v������M���'+�& 08���34�=y��D	Q��a�������K(=E��B\Flir���irƥ�lG֔�{"IǏ�'�Hwa��o�T%�&@oq��q��ʼ8_M��%3�ۃ�b��V�9��&S�l*+�AظO��lJ�3��L=��9mI��R�|"	@LU"CY)���be
0@CN�ƔH��
��²��b�p����"�p�1V�5�e*` -�s��6N�SF5錕=��� ߗRM2/��:`=\`��g$�p<B9-U�Ud�J��%^3�SQ��rߔjT��D�r�J�f�d�v-�Ne�ڒ1]�5�JPq�lؐl54����֔@ˢ'U2*i#OE?
��dX����k�U02.:OH�Q�N%�IoyiS�l��xIFu[x�n�>H\�����)*�k*�"�PO%��J�Iт�)�r5Fኍ�)�`ٜ�)z!*N�*�@aX)=yL鑘(�&QBS�Pw���fS������ğ��fya3��ss"��<y�����%'8Nk�uC@���� Jz�����?���\����l6��T�'�/����^II��i��lѓ�}�]	XC@N���e./����?9˔�G:Lm1���\A�	T>���y�U�'�,�����9HZB`,�r)I��5	5԰�
���5��ꎰ.W��*�ɍ��e)|�I��)0r I=%�������V�5�
�R9^I��=� uTCr��X0C���2Ms��}Cڢ��R�l�}�O�Ӕ���27�M����C��
[�oG����U�YQ�Ӑ��e�5�Q��<5ݏ �q�!���[f%�6��R�EO�$=p��D��IVҳ �
�vT� �ߑP)�[�K�m�	T�b�S�`gy����S�[��(�
hKF�`��=�Td��~����]ʧI����Jz��39��T_�G����2Y��>i�,/=��J�?�GOS�ocO*`[Jv32q����0�Q��I�  F�ψ9=n��JCB�4u,.Уz"C��j��V�a�L�F����B�\3�S�+�g�%��
�8��È��`�);��)^��O{��y�f��H�4^�%D�J;��pY��H�M�,�a ��E*3����jUYRU�kK�\:w��9���.U�����n``�0���m��}���7R 0x�D����C�C_�!e�BX�	˥{% R���(��2Oغ� �]�/��'�YHH�С��p?Tc��VL*���0����H?�!��j#�I�:�r?�8!������TN�tY�4ܕ�'�7-J�1�r{� �	��T==�AX��7�DQAf�f�,.�U�&��݁�4�dh`�SWa{�/�_����{����IlXn��ɪ��ϭ6/r�a��q{�6ς��6�̈��-��Y�y �K�U���dPt1D4�;`����DO�讑�HXmރ��5{�������?wh��>&��x|�������}F^���*K.I��K�t��������4�:dP����H���H�#T ��{�JIǫ�S~%y������ h�/��\+]��ܓ\�Z�R��x)���"���D��c�����U�hϵ*:u�I���"x#^�������i(�ʽ���v{c:��C�-F��Z�I�����YF����7C�ܓP>'(�6�KK��V���rNbk������(�V	hH�ؙ�� xG���'vҩ'3����>�@J�xuJ��]�ͰObe~9�N<W�M�|6hDrR�r#����f�5�(=i��$N �t�HQ�o���M^�j�#�*_��õc/�A��)����O.(���� H3?��t�x���4�<	8�G���+�$\���f�̌_�R���r�p�9�?BA�7�F�T9^�2g�)��'�Hs��HL���8A�� ��ۚ零,גe䋤��61��taF伂�3g�������ʜ��o�z��V�F�7+�n��.3s���K��]�|�J��Ѝ�8�;��q�/RYDG�QE/�u*�Z5L�g��t�Ϗ ���,7͜���'��Z�x����r�.+`�ĩ�n��Q� !�UH&o<��7'�4�U�+��kԊ���@�T��eF�����^+h5�!�;^���{�X�C��C��� 9�ίݑ���@�4��u��Y�9��+H/�&�nq�2�	�ȯu�d1��+9�M�l=7�)xh�T8��M���>a
E*���b����
�IhWn�E��j$S���o�.�K�+��X�R��
 ��"e4���ר���?�"��I8O��+DՉ�Aa��'�:�zI%d����ݞ�ys��[--���^ؓ�Y�\�D/H�DR������b?~0I�ϓ����C�k%���Q��y)�z^���!E�Γ�%�$t�xYD+oR�@f�P{�y�!?�%��t{*'c��%g�[�t ��n e�������O�I�dA�G�xe~A�Z�~0Lt�H�����ێpL���T��*��y��`B~9V�`�y|b���<�E�k/��כ�je.�y�Yo���qs��j��
I3�I���y������g��z}`)=%�y�������R��/a�[-��� )� S���]�k�>�_/�f�	@f��Y�0T�5�T��@�ԯA���,�K�t�5�<���;o��̸�6��Ht��r��Z�]�Ԇn�3^s(�Z�(Ȭhu�s^�_���w� Y���cO��10	�)�[�)�7r~0�% D ������A-��)��L=��0��n\x���@�5�)>µ$bk �6d��Y0�	r�y8R�\�<bFK�ޜ�U�[`F�@:�8�!����pR{�����GÌ���	�H�<o�a�h8X�d�4>��aA��y���*����!�����F6�*�y�0ٗ�cH���Z���a�n�$O�g1�����P�D�j����Ѓ��7���"��{$a����6b��-0���2�;fȨr����cz��@fao@�1M+��9�[�V+�z#��6��b����O���0ئ��	2�L�4�g���0�KY��GHNI��[�0o/�p��yxeP6La�#$���pł#��@	£�z1��}��ȴ��ĆxН�a8%�~�Ȕñ 'h?n�0nһ�i�:Sx�2��@r;�!R#�a8��c */I�a=o�a����Mʤ�k�ƹ����0�),�f���խ�Kg޽�.����<��X�v�#� o&<o�a�~�
��o=)�q#���r  ����E�"<�'2����rވa�kK�Dz?)�=��@Hʻ
J�6-��T�⁴<�J�x,"�p�Ap
>fa�J�q#�4Ͳ�aCʺ=�ټ|#�����D��*#�F{���2�w
 U87Z�_o�0�|����7S�,�mHD5U<�Z�CNJ���a���y^)����SE�04���
�~�>:�y��a�=�,�l�y��H�b�<����d�tg�������^��0��>���a��� ��ԍ+-�����މ	XH�T ��ވa�+B7��@B�r9Ȉa�o� �ӤB�����g�ܬ�,t���(1t@z�����Ւ
��>Ȉa��ZRp�*S���1�D����o��/��LF��5`p�������`��JŞ�м"��T;��rO���@d�0�����
#�u�[`	�*�*�I+�<VFC�-�@��W�,�Sd{��^s�C9o�a0�I�$G�y��?��a(���i�f� ��a$!.H�2�|<>��H�_A�*0�1�:���'Dw��"�A���R��{�,#���)yH+�a>���H�.���9I�L��"b��0.`uX}�Ï1ZC�����=�����:tCLR��T~àU��
�WF��v1�A5`�q%|R�HJ��,��4-�v�y3r
8���W�o�a��PI�,ر�F��e�I�:S)���Ak���2:�"��-0Z�<�D�g��sSà�����������yC�}_cR��>���|MAE��>H(`�i�k*b���_Ae�O�gY�&�"��O��@���1���BE��)x�R��ރS�������x��OY�:ӾN�"�Q���p�W�l<o�aEw/>D@�;�U��8*bEy��K�t1�x#�Q��^ri�~�=o�a,(���8��vz=�F�~�!�T��G��y��Tg����0
��?'��Ǩ�6#��v��/����/߈aa]0�B���X1�,0hHj�*b���^��@�P�R�`��0h܊���a�~�O��\�n��>1��9��t9�y��(k���7S*6{���е��`�' ���#��pm~o`��`0�sH1�Ί���{Aj�uRGC��Ҥޤ1��8UGC����T�����a4}7U`p1'��up1r���K�ky����g:b�|*��^$�uC~� /1Lx�����g:b�qo�#�q)�;�h�>^5�i�b�3���a�^�Oa)�
$�g�7bL!y �GP�i��-bL�|��y� H���1�PޭhE�<I�sވah
xU��Q��c1C�FS�ɏ��w�1�~R�TC�1KG�)����ݐ�r���a�<��C87#��/t�0T����i±y��#��!�j��?��M�wL�0�>���[�U�L�0hUAa(��Wf�^J��0huO�2Q��U��(B𴆊$���+ӷ�x]7�P�wx����t'�-0�zC7��0��y1�f��>��I+<^7�P��;�$�{�D��"��V$���SP�e1�c�Fp�H��&b�
�4�
�M�P���-b�J_7d��|�Dcx�쀀����j=~�à5�����p ��^'M�0��K����㐉*lP�d��&b�߇�TW�����>U�ݕ�a��W.�u���;��F�1 ���&b0J�@NH��xC���� �I��}��Dc�{����k�����DCu�`8�Ӡ}�a�
*�=�F�c|��D���zhv:�q�0����w����R�ve#�!��^+��QXl�-0dX:�V�[�AFxc�1e�!y T�9[��)|�l҄q��ue1��/��l�O����xa#�J�>�b���EK�Ҭ�-0�ʐgY��#?�Kp���06sϸs�4�4��h#���4l��C�|l������\�#97�y��A$�BH�y��t���җ���s�P?e>^f���}/,�y?��S��>Y��
Q����-0��Jc�P��;��[l�0�A�0�^�2��8��X�ҍ��B��7�I1��YAH#U�Fj#���c���.Hӕ�-0�h��?�q���ECu��7v�����ك�MgA|���6b��p���0N*�-bk�2=�N8Һ�Q�[`K���y+?�Y6��.Z���k��պ�3^�N��� WuQ���   	pHYs  %  %IR$�   �eXIfII*     (           >       F   i�    N       %     %      �    T  �    p  ��    x       ASCII   Screenshot(/��  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:exif="http://ns.adobe.com/exif/1.0/">
         <exif:PixelYDimension>1392</exif:PixelYDimension>
         <exif:PixelXDimension>340</exif:PixelXDimension>
         <exif:UserComment>Screenshot</exif:UserComment>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
����  ǸIDATx���$Iv�<"2�ή���ٹvg�b��hF�J&��Lf�*�>���>���H`���ٝ{�ﮮ3��p��;�=�2��fz�SSY������{�7]�E���s4�O�7���A�h?8B�>^�HkY<
�w��G�_��}�� H8�:��ȓW�x�g8�9�>��ÓB��El҄ z��Y��;�[bϧ0gP�^A�hLQ�5Uv�\��nru�@_;����9��O~���]���w]O�ŜNNNh>�Q�u���3�Ni>�1��J�
B����x¿Gc��Q�?L��ф&���J��z�o0A����oi:;����� ��ތ'|Ѷ2����9::���}�p�&�ի�hē^U���d̄�CM�L���m��ݣ]�=ij��f�|#	�&Т[��Ǐ�	O��l΄��ʟ)!�u۵���*T�߅O�>�G�1�z�|�c�'�an��],��e�4��ss����6����b¼|����7M�,������ղ:`�xzx�Y�)s�t6e"t�!3!��/���%������d���q��mnn�(�Hk�3@|O��?�}ʢp��N�:{��{�0|(�E��F��bd����E��1����&ƂuH+Z��T��pV38�.�(�A?3~o�?��)_�����f�Ҍ��ڢ��ѽ���ÜRQ���oq
�Y�a�ȑꂕ���)�9�6v��1���ų�zs�0,��YO���	��n sY�u]	���P��������<T�ގ�p�Q�� +��9�<��?4V�)d�H��T|��mml��/��J�a��
��K�;;ۢ����D�=d�r��]�L\�6s����X_�|�����TP�u��o6A���Eʓ��+���=���+��W��KL������{�f<�@N8�By��'"�	rt|$bp�����Ç��`������}c�i�#�5�O5�*sk���+���.ݼz�a�X8F�ȩ��$�1yc2��fE}��u�tbӴ<�?�?��?�����;����p��o���GTc\Pӫ/�B/ݺM5�+v�����L�Rxܧ���!����A�<������(\���Zs`B��U��oP�E��P�v���VxN���9�_e΃�`� ��"�����7� �'*���Zt$�c1�g;9V���U�#���ǢpcB�|���l�l3��Q��~K���$�rU7`�*�1=!��`L�t�#�_�儰5���-r2;��!�z[����E�Jꩅ�� � ��*ӓ���X�#�m���>���d�t����9���3�y���ٔ-�y����.�>��	D����Gc�(�&����.�{�ŵH�1�<Χ�1}!���2q����	����>��cz�����^�I�s�y*�Ť�?FT_ܿG|��k�6K#�*7���A�G{e°��7�������?��7nJ�̑"�@��(�/�_����4���ǂP�P�q� U�������+$.�2.���M*c��K�m������������[w��?w�n��5�W.�X$E�;��&�q>_��ֶ�#�⏂���	�0�����0tq�ZM�X�O����
#>���|e�Ŷ}z�`�����L���v&����b��{ e�2aqs�ݽK���ّx��,6:�d||Mx�Ă����c���b�����,	PݼyK�w8gE�w��B�i��ϙ,&>�/�t~w\�f���x�3-d�Fu��K��N=�_��h�z/�(���#}~.l	(�$ܺ}����Т��9u<�LD q����G��FB�-$^a���FL�_~�^~�U68���rΌ��a_x�ga*�\9AVX�xO��U���e���?+	s|zBs�j�`һh��&�3:�XT�!�}��T���	��F���ߘ'n����Bxiu���l�!V�Xt�1(��R4O.�jT' 4cV�x�k/�4L����(�$ $4l�P��Q�͈.s�����tFǰV�9����R������Hl���3/:ԏd�I���I4&F����[k�	��>�>1k>JЩN\))��#N����ʘ(�<[�a�reHb�r��ǡ3`sd\j��"�ܢ����(u&����:% ¡��b٘ �r�-��Gq�yP)7�o�: ���KB��r���0
��Y�&bq-�K ��Sх�M�:��z�4����ct���ϫ��\	��U�y4sI[B�/K�ѐ��a�C�R W`�c%���5�AH#yv�9���f?������U2įdfm��wo"� �O��y��#-h{kK��V�DW��$^b�-���r[�9�7�}�'�)x�[x=
<��{t�c5AxP��N�Nh�ga�6xh�(P��d*C�Zro�� �lY�KsX%�T]��X��\���d�0e�������'�W�������M����K����������� �P&MƄ���𺣖&�?�;}q��N�@~��rP�жQ�%'�C�\�4:ɑ�� �d�yR�Lt�]b��-��bF"�@�d0�c�����|��xT�J����O�Ν�d�5��J<���)L����f�h�b�Kg�>�V�!z�����&B��#�:�	�_i�!XS�k��R+r�i���>��666��W_�����CU���H��JuKWB�>����$����H�Iq��-h�sg�
==xJ�!M�J���1_��	�D����E)p�尞HC𢩪�c�恣Ưf�x��ұ�Oy�AD\��K��4���.s?�%uE��J����9����"��{��	�Z��,u��R6 �cU�h���,�3�&�[�1�pQQ��Z����x7X�x���Ǵ����z ��8!��s��+Yf�x
��&�1`��HT�W*f]��nȗ)��"��.�F�WI�{n�b��I�n��٢s='�8Ӊ.�ϕ+WD�!J_�qCN��R�$O��C���1�nHDȋE�Y�p��,�7!2���I�'�2�7X41�r�*qA�p����.��p�FY醫	���zC8�$/��SLi >1���rY^`��ݢ'�.�h@M_'B2�B��@Q�Ϩ5�F�Vɹ�EsIYe�j�e8�9d���ɣ��@!����W�Ĳ�JX��U��r�ؗי*C8��A5 UAg�$nY��&MP2TWf�+�9�y%b��Գ\���,#�L5��	������Od��� �k��'(d�g]~�4y&��7 �{�zU�A}Sn����>m�h�ِ����>�������}��(���M���qO�&HWD�(�=>9�����ޡ�W�"�ϲr��֓1cr�����"��t����`+Ox������ӢKˉ�AFP�FIN���|�k�Q���C]�ɟ�JBE��P�3���B�]6<���}65� Āa��c[O�g�*9���*����pD^��y]%���j��?���|�,)�����4�����mߓ$��d7�5r���q��Q��8�)Q�'��ұV�Sz�J�y�����zkkC�+=L�ɜ-d��a�lln�R=|�T��Z�z}��� �����"������ə�B���������r6޵|.�#�m��+vʥ�9�q-�
��'cqa��y�"�F�M��G�.I�5�������+���(�&����܋�wC*��C��CD�1���Vc����> -���2�߰�aԁ����~��)��H��K=����� "������+1whq���l*��|�pz|D'����,��+爡.�b��\T��Y�2��0�uX-9�t�mmo)f��W &��p(������J0r ��&��X
�`ۻ;T�c�+�+�n"C[�][�#O�<���C���T~f(Cూ��PЃX�[��(��c|��U�.�[��ń1��
G�1��L����3�1y,���Z4��V;j-���ȃbՁ(X�""�Dd�9(9��ꫢ3�P(<�X�{{Wikg[&�\��K�0:;������}�tX�O��������c���`Ԟ0!��, |�T"f���ի���_�^ ;�7
M!�I��GV%�*�@�@{"�(s��s�ITȨַF�0yw���ϱ���#���Ipk.���)���xX�;L &f�t��^�f+�SWM�א���*���Z 5�����C���������O���;�����]��A��[	<b�=~�^�s�^z�e�q�,&����]�F�PW	��	|q1TƵ�(��~CƢn|�ɾpr�0��<��I��#�|�(���G̖;q��@<��۷�&?p�"��	�x���g���E�� �yҎ�<�O>��~�_�o~����L(���ߣ�B�)s;)p�����\��c;x��N��B����z����W�\a�>���+V��~�L���ļr������V7����7V6V#^?z��޽G�<���B��~�7�HP�E��M�����������d�H(����I��=�Zv�7p.������k��O����޽�Ro�_�����L�I<����t��=A�o�񦈹��{_��.���>f�vI?5�͢�⋲�J.'W'_ٹ�bʅ'���WT;&`@<����C���E<@q޸~�����M�{e��rU��i�_�<���ҟ|�1����-=dN��;�0���c����I'�B|E���8�U)	� "���O��#�޷^���wK��,��?~��P�h��Eses�~��~@?���D��g���'#)��ؘȂ����$���ʒ�s���	C�xˬH2���\��>sB���O>��>��S!��^�W^yE"f��)]i�D����ݱ8
�88B���@��/>O�Xo�����?U�2�OFX�%�&z@�/>����/���C	���#��1� �{�!f16��ڵkr= ���(O���/g�S0~\�	D��jĨ�},;V�X�����B��Պ�fu(A�	��?ؿ������w�cA�[:s��@.S�߃8�W`����ŗ^y���'�|"Hv�
��bbϘ����_����i~ʜ���=z��!�`p�A��b�����8���7�8�}�&^���p=��
��d��t��f�;��2o}ᠤ�C���:���ON�ʂ+0��ypX�x�	�	i{��6�`�#�T�� �b=p�u̽�w5w��	t�)O�w��]Y���|�+qc�ĸ�G[&���n)q~F�/�����E'�o\��vö��77oܐ �'�X����a���Ct!�;`���r���|��y,���( (������G].[�"Ab�� �@�۱�Yy�ޯ~ŨE{��^9a�|��_����tN��) Lu��WĜ�k(k������$�u�5z�����?W�΍k9o�_�<yN�t)���>��^�U�!+���pL����5o i��a^h�x��[�fx*��_bpp����<~��������S����x.�}׺���I]��Ѡ���H)�ho��!�0�;lW	F��z��u��}��Ǻ�q���Ao޾�,r�o���^~���������WR�4�x�2��\c������b,<�n����g,j`�� <@t����PY��}4���`��8�~[3�>�ЗDY��C�ʋ���≸��L�'���3�dU�uֹI�}E�>�:��� �e�z? +qƱ<Ɗ�����ؚl���҂Wrz�e.&J�l��W����X�w�z�-����N��Sq��L��(}A����Z&
���@�<�ڬF�8��a[l���LL�L4,} z�w�b�O����ͯ-�q�<~�evF����I���}�a�O�ܲ1l��BN�{�{��������"��_���y" �o3���/~�D��av������f)�P���S0Y�*T��f�,AC�Ufb�n�ꄛ���N��k4�Y��u��)�)ԗpjP�Po���,,x~A,ɨ��]���>#)�^��\n�/_�#a�L�j����y��'���'S�Lq[�`QN�a�hl�`؈�-�M��^���$�.&m�>��3�Bh�d��=�}�����l��9jS�:Ei�(�>16xR�����LI3j�P1U-4A��O����Zý@D�ۛB$)�K�g��DJ��ڌvKی�m���_���o�N��(�����ՊT��4�^���8fq�ڌ>g�E����ӎ��=�ʈ����x���s�5��X��3J����Tf�XYA��ύE��6��g��m�G�V0�+<�G@5��Ome�S��H�L�t�ސ��ٞA�*�ߖ8~-�>V�c����
�ؒSVr�jI4@��M6���;�)�'�����n ����ߡ�_�5Wz��n�}j��>��b����X��O\���hEac|��;2�O�}�Iu|n��r���}��GP?7�(��,� {�}�Tϋ +�t��Cf6&�eR�=`t� �F�t1�x�gG�(2Zy�7İ���g_�O��oX�?�*��}�{�j�� !<$�yf��oj����3|o���~�0􅱩1��x�5[?Z��T��D' �q��%\����N���m� �X�����[�!{.	��Cؒ�A��9�)"	��3���W� �
ԅoAΦP*?�_��>����k,.����w��TU���$MX��1�rT)n(a�^�1 ���8$9�n�G���[Ҟ�n��6x���K�Ӆ�23�?�VX�Y��b��J% �B��Zy�R�~%�~e�H�I�,�^B���$�X8"	��0UjG�D���T�&1�-���&O�|!py����{t��)�?�������o�K������Y+U8��خx@�H�e��'�`g����؎�h��7b����CD�0W`��|,�ƒ2���0�nr�b����M^`*b�a�ci�)��n4g@����#X��W6����LV��#�����M?��OduI�a�ڪ���G�lmo�_a�y^υpG��� 2����}[�_���d�a�v[Z]�&
q}�����q�!�^�c�'�g!� 7���<�c�� C�J̠���'J��⅀ژ���b=~�̮^��P��A�=gS�.s������?���`����������>�7�z[2Fn�D�5�����槴�l�@�A8:�;��?�w�N�X��MQ�����˯�B/0�x~V)	4� r�a���w��\�3::=��-�ܞm��_I�B�@�XD��7�^�-�p.$�B}�Y ����W_�#6��M���M������r�:�'`���K�gFW����J�ӄՄ��3���������o�@���>���[f<����D�Jp�[̅/����v8"յ�[��L[��]���/��~������?	A���񓁊��Ap�/#D�7��D���L�;����`|���bh���H��6���Ap��Q�� y�s����=�^KJJK@��m'�����}���������C&�(XV�s�X3�j�E X�+	���߫� ��KUB��I�������������D��i���P����ċ�˟�\�B?<��6��D�A�b!�$�ϻ6�)����G��;[t���P.�����LH�GN�[�[v�P��J��	?R-
~��?��M�����|��D������s`}��w���Ġ!�g����7^g#�����<���{�Ͼ��d  ^ʅ��v��֑�� 0�/�տ�{���1��m�#*��oݠ�c�C�}����5�� ���g���2�T����w��o���gn���-�RX�M�$A�
���u��{V0�&UC��H���^`�o�)+��u��WX>���_�k7��ہ'�֋��ã{��­�����/
Zdz�n�y<-)�"�*a��������/�����^�Qz`���7/<���0T�����>}��\{����?��pߋ��l%���\�9�����q.A��ue�	b�z�k����A��w��bE��?�Gz�_��@��@�7�}9�2nؒ�[��������$���������B�eL���[U^���`��hr���,2��B���G����O�#{̡���gn��(]�- �>�HԸ�G�o�F?��w�����/��:R{��$�TȨzE���%ɼ�J	�ߐG7��mO�>�������?f��%��?���� D�泩X��$ �N���N���������N�r��$e5#):��e6.��Z����ٍ۷��-��_��x����?�1Қj�-�? @$�!!��<���">�dD	��sb�H��R�x�/x$��.�F.�:�+_���͉��|T��Rƃ���?�_����|�Մ6����6�Q���.b��5��M���=ԞG/G��c�y_H��b�be��ٛo�E���=����JB��|�$��g�\�1|��7��̥�� g�+��E�r/Җ9Mʏ��~?�CB
�g��J'eY@Q�s�޽k���86�����*�����s��ce"!0�߾���&@T�7��k������[�Z��\w�މ8+���tX��~�;�o�����a����Aa��G^~�eI��v�m��M�؍&�F�}�(���P� � �~I�8����T8�r_W�����N��ѽ��Lv
�[o����@F�SP�#��������#$��w�O��-��Eٵǲ��Q����2��(�f1�}�;���;.��#+D�k�m��]��">�RW wU³a��<������������ڝ�paY�	0�6��H�6t˶�N#�5�D���:�4�
�Ţ��i%k�o��B鲇����ؼ��>� ��r_CH��\���:��^Wh� �$Ҳ����[8��e�ेT�n�+n�Y�.�U�  Ψ���e��k�D��A%�	+��ioew�F7�2��+ԥts��X��H,���[�)��Wg`oL�E��U�,�֬�����;֢,���D��v�o�X����U���e�2��[ۢ�և.d�L�Ք{�`V��Y��u��Q��c&�-�'�锽sV�eo���)������w���YC~�}������E(䖀_� �j�k~�>������U�<��D�^�T4t�+�w�&�+����r&y�t+2����uq����<�%)�A�1!���?T%HO�ABZ�Q[�4-��(��EN��$}ˋY�`�_� �(Q{��]�#��z+[B�Zc���#{������±��*:��6]GA��C�I-��e��t��ظ���H%��V�lib�SŔZ{�g�S�~'��_]d�{���C���)W�i�25��I����J�%��D���1�3ܓC�V]��r����=Nj�䟅�8!�X+����o�X���R�DU,����9��{>b�&RF�h��^����dj����+��	鰕M5�I�����yw��
�	������W6�uA��;��r\�mց4\��G�*I[jP��ˢi�y+�H%����`[ �<������
4��řn�����C�Mn�`};i,+��o^ޣ<�a��s�w^(��W�Q�(��=)��瘣���P:QS^=�*u2�i�S�t��:�~Mz#��??��ׄh�b8A��N��1�χ��6���j���/3	��!t`�ڊR�2�o��Yk��ET$嚑S*Qv��)����<��M��,�x�����>2��t�`��E��G���2��ϋ�K��^+~)���W	���Y���YUt���A�[Ɋ��1ĳ��pE'�ťP��%����#o��� �OZ}��� g��}���_#�[�DRR8e�$���v���t��Q��Z}�u���@�\����*�9(�_�l7!��-���t��!�M�IG������ϼ�2��h�|?駸�����j3���y���[��s����� ���a&�*d�ǹ�.�!�?s�$�}<���]b�=.2ₔ��ʥ|��t��gM�B_�{���7�xn�2�[�MT������eb+_ױ>�J��D���ɸHg��]ĥW�ԗ���и~�N�e��n�++wώ����c9�0J~v�!�^���%���x��n����#[X�AC��]5���p��]�W)�"p����YA�@�f��{H$�G����|f���g*�����:<���Y��o�B�������}�sˢ/�)#������]8gb�۫�SH Cq�x�e�9��a�������q�\�M:���%�?+
�V��|B��
�LI��Y������tDg���g����6ID��s�c}к.Ëg.�^�����7�lQ?�Y�y��.ow,����N������.s�{��岾ş'���E��aq@���8����9Xɫ�]���_u��i)��Ķ���znyK���9%m�OKڢ��C���Zo�0s�?�m�R����#b�/VF��]t�r��O����.��c���Y\�x��z�@۸|~��>5��Ĳ:��]'�BJ�;#V��9s#�o�8'�zh�����2�xdL&�}��AO����l�h�K�Ń��зH��������Iٚ�qY}��<c��0Px�2˯д�d����i<�C�O�il��_�������-�pF^Vq�!E
�Ͼ}I�<Cd�U�:߁�ş���ϲH;.!�pH�OHu�ϊI����r6ܸ�м�8tT.�,R(>S2��3[���Y�c&���I����yw,\$�~$$�k����-]9hh���J�%��@fյJ�}P ��]�r2\N��l�f�i1�"-W+�jh{�;�3Uw��V~���2i�>K!Lq�'��d/��6͉�-��Uֵ9�6��2x�ٽNV�y0��zXz�4_�����6��5��(<�̶Jƥ���O7J�i��K6��b��Q#��R-�ͭ���	��sj����{ai6��q�w�@�[EV	9:r��4{����r����䇳r��IRr��3b1!����r9[��9}f�<���w�v�B�/��S����I�&�A~g�b�s|�����+����$^���~��a��̔�Pv/+�s��dm�ѐ��I#8���B�9Y�t�Ϝ��}ͳ���&p��y�i���RiA�0��w9��vw-y�zo��OX�5�gՀ �:'�n�Թ�*�B���s��,7F��)WG	��l�T��UH;�{���i;��_�+D���	O/�ՋY�}�2�k�,�ӂnE+��]$<r��ד�{k�-z�����(�����{^�T�38��� ��.���0P��Q�_ł�tD-�������l�߾����[��ER�wu�D�uι_������m4��x�AdX��TPm�R3[�,Ψ�.)��[+։^�;L0F%�t0���pM��}K� b����ґ��W*����h�^��votc���UQ�鏎�ڪ����LD�g�����&�;q�n�޶��y����j���t��m�f�1��]���'�r?D�C~������E��w��mp�ŷ��M�����K�RJ�BK4��?P҅n�*"�vC�G�� �W碆���{��"ֹk�t����Si�!��G�%�t����(S�h��ߨ�G�H��*�jk��;��@����I��믿&פX	�5�Π����F���r��zJ���r�1�����1m^�J�3����dF���-OS;x�L՛�o��u?©m�����.�x�)�����^[P��ڡ=��/D�m�(wB�!��:��*�zhT�"�\?>y"��\�����JŽ�����Ûo�\I��q���wy]=��{�Ԋp�Ź��۷^���Ѥ��TfK�}#+���CQ�~��v��؞2q>��s���|��u��sE���A���}�x|@-+��1��������՛W�f��������������ͥR�6C����X�&Z��d���Fړߌ7ebd�;^/�������t��N,Pa��.��2+6����v�e��iׅ��ފ�BE8�1���������4���%��&�\&}ww�9q��=x�s�\TO}z��$�n�o�AT�v<�tr�m�H�-Ni�=�'��������H8�ڵ��V+�yU]��l�C���K/�@���ZQqh.;�$^:Cs�mG������>�������.�C��r�c�(1m|�V�A�tM��j�w4�������}Aw�=b�tf�/���]�3���k,�1�<�Fs��	�lT�-�t�s)�D6C���vI̝�+Bu�(���tK�H�GҎ�weo�&hj߷��Cad9!�U�*��^�"��K����H'��,��'{�O����G���B76�j���>��c�W���+���b*�. \�s�QE�vJ��Sِ�ʮ6���-_�X��ye��G'�窝3G��L�?x�7�,b4t���m�W�	�r�b���ū'��+ t��u�2nA�ob,��Ë�V{�o0����iGF�o�cL"��e���h�t�Џ�X<��O����H�.��[&�tz��
�nD���=�-�����]e����O�0r9��т��m�(A��cFs&��
�;�mn�HK��m���;�U33���e^�^DS���pG��r妉676d�����#�gW?Q(��N��\c������G�0�?��um ��4��\�/4
��-��C8Yy�!�g2���f�|�Mǰ�W�T�l��AQ(�@	5Ccl�-�sZ���O�y�u�X;�������AQ\�$�lpZ���ъqJ��J�-E����������r<�h <�v6����~���߻+���YFj7�#p?m�6����T�a�9�HB���\}�U����}�!�0vw��b������#�˖�dd#i�i�ؿ��{z���o�(_�ER�i�*�A)���H��ޖ*�Ѿ��Н�f�9�>l𷷞\U=O4�����W����
q�b��-;)��b�޽����]���x�m3&��l؈��bH{�/F��������EH�����)� ��uM�ܿ+��mb A�,Ʋ��DV�CA�6�]kH��DU�E��I�֖��c�=�;�|����G�����d�Ȉ�&�旓]������p}$wP��j�6�Ld%������j��ڶ��R���G��g���6���0�$�%��h�{����+$��P��F3�q:(7 ��|g2ސ��z�_(! E�.���o�9p���g:����x��dSǊ=�f�m�<�}��v�Z�
�k��V{s��H���Zl����!�H`g&�G���<����{���V=2�/m�:�B�Mnc5a�8����PWI�b"*k��M��j��%��@�e���d�����CF4/'U�c��6Y�C7���=*���K%������H_��;!o#6Gٍ�V$�[��6��*�˶N�/�)�����)���ĕ�m������d��Jj�4�v��d���,O�
�dW�Z�!�C��d8�����["u�>Pp��b�g`��Đ��W�ҫ�T�t�W
�^�p������Ψnd��@Owx�]�q�J�ʔ�"M�d��6�#O< ZQ�cSv�Q�)Ȁ�1 ���@p�p��eߘ�H��,Fl{���k%z� �>.��/���z�-le6��1��C;�IY0���T���8V:��5���a ������'�%�Om����-���5?����)b�U�X&i�WOu5�g�[�`��T�?�p8��L�@g%
�jl�:pވ�ȸ�N��Q�.E]�a���<�P\�T< .�����6�nc�'EF��3yyp����H	��0�vc��yb���U��9*�]���f[�J��^�L�m�����	��o�W��c{�Tf��uѫ��O��`a�o:��e ���mX?��K�V�P�>��	Z���̀y7O�Q�х,u5�h�8��?�˓�ӭ^=7��w�@_�c��7�m�v=::�A�t�5�5V#<��v�t)�"!��ģ�Z<�����8;��TBi����;����Qg�I�I���ݷQW��4���gp�x��y¥2��ql��L�y�܉�(˛�$���9���*�X�ط	�zg{��-�aU9�p�9�͍�1j�'GW�K�lK:�O�_�Ŧ#���2$�X3do5��b� �l.����o�����[�l��ZDܢ��c�U��֎n�Luwk��u�8�H��	b>��2��P�cV��҃�+���ϱlT�6o�`%��/�N��4���.V��3�011c햻ay	E�i�5ڇ�'2_��h��_��A'%����=�e�2<m�20)ň �X�Q��b���=b]�1駧3�y����������'],��.�C4�+�>7�Px��Q�¼��K�HvS���b�kyR�*�>�1-eEF���܃\%@p����R��;��͐w-P�Ge�C�:&��̐�;�W���-��!:������l�K�k���Z�ksc[�ۗ����GʢjT�b���E2;w�@G^��&�Y��ãC�zz�l-���>#jG���8��
x�����nI_��1�0�X��Q;�m�>�Ő�$�egJ߼�řl�'�F���]���wc�7u����ͮ�%���%._�LJ��e�!8�����A���:���vK��)��r�6Gb#rK�(63��bt�^Uw�d�l^;gzl���e�¥bPAenV��_f�hK�WKO�pg��ed�Y^0X��Ƃ�2��8n	�a*��AʀØpз��(�i���+�
��'#�7/�lt]٣��m�pVA�7����5PR=�+lG�d)[�5�J��5w�M�(��vz�������������DJv/��%�=7��ut%�m&����mf��3���ʍn��[��g$��GPt>e�*��Q������6$6��V��������U$; `��� .�m]7'OZSn���t�?�CI�59�M��f��G�7Ţrq�{B��G,�W��z�����(�m�1nl�h���I�%��y�ߛ[�	ek�Ⱥ�"�Cv+�]��沽����wY��H
��$1�?�r���U1	�d���w��l��gœ��0����!���R��H��7&�����EZ7f��h "UHa74aTV]k�!�C�g	��*)1�l�Ӳ��Ԇ˝ �ņ<�û<��ֽ���LYF��!�
�'^���?�`"�b_���?���h���,��H�()o��6�����P���S�b�g���{��+>�)�{	�e�*�mѠ��97`0dpW'\k�m��d�V��?i�� sҵ������
)C�?@�-L�~P�!#D.	���a�bro����`��7��i.{~�O㐑������]�8��y��5)�-|�H�q���½��鋭���˹�y���s�Z��y�Z�Fq�3�&�[E��^~��u��G@uZ0~�O�[������_�k@���:�8��Y��±�_��ڶM�����{��0��X�u�R��'l�^�h�;���х����ҵ�=�o���__����X�PY1o�g�E+��q���.�ʀ�3-B;֦�����S���9�==��|nѴ�"1�EN�7	���cik�|Aq�dQUܐ�@D���y�&å�S���=+#�Z��HQG�B$�#��u:Vf.�L�Kqu�+����,�RD�	.�z�J]�+��l@s�=�&�$fP����]�2ǭ$B�99���;[O.W�1��bR�]�C����S�X�)�Qz/���w0nA�p>_������m�Ήc��IVu}�0o}-�PO��٥�e}��e�L�x�l��ގ�#.����I���2�#Q�M����9K�\`�5vX+�o��(ɘ#�#�f�o��g��]�i;��q�\�(���^!}V�����4y�]$��*��s7+W���#f�!�!;2W�wu�NP��rJ�!�!���".��Qo��M���L��D�����
�V��tK�.�%BN�+z�%����� �W�]��f��ԙ����x��Zaz��:=@�Q�dx
N)����4��dD�pV&��Fhf��>��c�Eb��m/���y����2�H�*�g:xTM�̱s�'�ȍIu�6*�ڋ+	sֹh�v�*Z�MU)�b/���PCZ!]G9ju�JW�_�8��b���]��Pם�z��lW�m݀���Fѫ��#+�&.���9�����dz\�8@�N���%�G��"���e�EGT+�]��ι��`�8���p�u/w���XK�leD�� �C�-�lAH&�/�Ե�U�ΪnB	g���*̂�������=Y-{G�=31�� �-����`��9v؝D�E9K�Q�=@R�
8�h�m�%����)xY�x�������5��ؤA)�h�<X�l��\c�?=�&%)Y&�{���TI�L�9�+�Wk��r�ui�H��n|V�<�d2_8db��3��3�0aF�����
�+Q� ��H	���=��8=��b��G)���s������*|^Z����p@'3�3�NA��{-Y���L�/���9W�q8̴�ʘx&PFK�	�n{d����H�I?�9s�(�C��x��		�\Pda��c�w�\٤�{��4�(f���\�3S:}u��{���NTw������g_Թ�,]#v�Ɇ���=.O��
��K�P���m%Gy�Hyc�$R���!~nk��Z5�.n!���"�1��jP>�3g�au��&»7�ct#Y.qhݯZ]C�d�`3M�C�SU���V�]Ht��57����l��a�0�}"�K�^��g�Rﵴ �tA�Y���.)���!v�m�E�?`�/_K{ )%�Ī][��ZN���!A�7.�X��lp.�=�/Ti��}���6���k��آ�^a�_���m� ����jT�dH�|�D�W���}(�a�Bu
Q�����4��8����G�MV���>��=|���+�������Q*.x
�����]wf���c���EQ �K�՝MR���>HO]��I���c��Ƙ����nOQ���r#�5�[r���y��;�l2��m��=�4����
�S�A_Z�ꮷ&8��!Q��B@��I����\I^�Bj��8��J�AA��>Xs�HR��Q!��tf��F�C^�Z�Lw��IG9�By�h�Y̢���&���g��z	��1f'bL"�av����"7&�������ɹ̜U����
WAH~�!��[R��#���J�X5<S���|b�=F� Q�%��|�	qH+ñ�=_��eٖ)}Yrm�=O,�G��j>����|��R��N>�c+��Mr�d���ڹ>e��}����\����C삳�p���3�L��+O溭���ͥ�hϮ�<*�R�vȉ�n����Uf�{i��Y�.�{�J#P����.7�$��zI�S��a�+ev)��T �B߈�`��M�P	/
��2dNpc�Aa�����MϦ��aP�+Mg\_��:��U.�g�~.�BY8���'D[��(
.�ͺ5�JcyK��<]nq�b%���J��n��bN���@\��Rb]\��1'*�T�Ø��5�<�4���+4E!+�G���-��G�g�OxX������#�T�Z�țx��fa�z�����R�R"F)ˋ��Г�V�P��^&B��^�ԥ���jQ�����J���@��F�q����9O�K3^�H��>_�	㫎�M0M�yU*�����w6h��fS�*�$����%hw!eϋ6+DU�R�%���8�'e�t��	^���+{�H��K%w�˟!t���VL4��S�0x%���r7q�0�|��)?�"q�C��_� F
��XD��N����k>��fDG��$�2"b(� �N���6F3ea��fªc�_"L�g$C^�^�*{�]HVr40�(l,�TcS
�����9�C�~U!�x0:�U\�m�IHWkj6���oT��H�؍y��苲�]l?� Q�s�}h��A*�b1���#:A�%�Ç��=X)rm��9�g#�|HU��o%��^ߐ���SZ����s�e���mob�<�֍!�8Qʭ]/	1,s>XR��?W�����*h�F�$����?��৒��Tc����%V�.�.���K���0�^T�0q�Jk���c� "�6��'7�$�3Ag����'0����۬XAj�[��XJ(b4nk���l2�r���sO^P
8�X��]�R��X��[��l����0;�������"k�&�2��ʚ��OQ�L��:�ʩ�*<�������U\��8+w.�)I��>rC��gV�����	�I|iYC�DK�"B˂EY$T�q]�`�s$$����Nf��x�>�
(G��y#߱�(d����h��,��Y�Y�E� ��"B<D۵.���b?|��>8~BO�<�I�_WQ��G3�&c�Q��BJ���j����ȚsEY_�=O�sJ�ER��ԉ>!�����B�Q3�#���Ѧ0X �H�W#.n�,��״���J�U;�j��.z��m���3�b��1�&��Hx&ABFE�j5���%���'�bz�e]<0X�Pb����jP�+�(�g�͘����srY(::<aҥY�Babk�@&��F������I�s�ͨC9��;p����h���:�m��-JP���[(Q���r>�����"�ƩsD+�Dtr|��0�z�YdB��(�:�������\~B�X�>������&�vĞ��0=(<�I?9QH�"I�]kU����� 7�V�
��Co��xq��/�)��m /�Fa���V����h^Fa���{i���Z��8�L�gjm��R�kb
c��ٖ�׮]����'X*��_5nt1�ҵݭ��.{��T�_C1ml�⁏Y)�Є���J��E��^����}z��q�.�#��Q�;V�I��#+�� Z
wk;�ɱ���Q�A���WA{��E���7���/zs6�������Fe*�P��\LB<aqI#F�����p������^x�Ez��ԏW�Z�)�5���s��y�£��Q�,!�O�lR͊mc�M�͂��ڹ�r|�H���߿/r����&�&�9++��M�w�"9�أCQ�.]�V>͜1�TiU�o�Ҍ�_�$���f֛r���5��	�"D�d=���[��N�f\)�֜�xH���O���H�	�����9���xE�۝�e��v��넖�ѿ|҈B�^V�罗l��ׯ�8�I�����QZ����m6��-��Br���s�t�F�C�1�G�Dי�1�U(-��\3G7��ǜ��AK��7&��z,u���Z��S�Y��},�����v)�q�ĝu����hi�tڜ2Aަ�L�rj��Y�n��t$*�Ty���ϭ]��i�[��J��2[�^]dm�ð�R$/FJE�����
yÖ��v�b��=DQ���:qnH�D>�`��bw����5l�/dNz:=i}����m��ND�Zb	���<*�t��$K[�i5(��	�> |C���F��h��,~1�yee֪`�L�1���d��u*��F���M��27�+Q;��f�f�9E��I#��_oea�Zapt&㫄�iL�"�_�(|�X��%����J�R,�w�!T�6���*	�ɟL&)���{ ���}318:Q:)A�y2�6�Wr��l�w�:K��Zܷh�ZU�����Q��T�Vy'QY���X]1�p��si�R=�UR����_x_��C�8No4
ҚusuІp&M�\�P:W]
�[EK֔�ή����r4M�(%���t�ȈTq��r����;�m�ށԓ�jM`�Ȫ4+Z��mۑfI��6�ӊ����t:1����.��s�>�`Ī6�<Y�A��j_�(���h��$�n:F�ag(�u�:5����)Q�^%�A[[lm;���8t�mS$-��~��`jmm�܇�	ж�B�L�BЙY�
mq��t��Wf��Ĉ���|b\g�!���љ�q}��5H�W��?쳨�zؚ��'$8ed��ec��ڪ��_p��t�c��8Q�J�͍-U��ne> H��\�������D�ܼ~��<z��	��	oMay�,������i�TWS���-�Ҡ��@�?O �?�o���K��u��$�G�l�{`��A\A,�p��#�$J~2N�Ĺ	�[��"WI���!�/F�-��o�/�9�`�ш\�sg������0\�=|AY�Sy8�-��B�bÉ'�Lo�	8商�3��f'kB�V�v��qp���.�1��>�̀�	�U/�Ƀ�nr4�n���B��T���$F#����Wj�Q�ig i(]W�6S ��"�����mۻ;�c��9q1��Q�@Lm2����5���1=�*ry!����9�E���WKW!\C�8>��N� �7�&�:GN�:�\�2�d�"s6�<�m��o#F�����,�@EzC���X��
_Vj�	PQ7B$w\V�ֶ�u��Q�Md�bBQh0*Z�K����U�xYI3��o�;���U)� h����Jx�I��g§EA�� �ܕ��Au��h�j�ʜ�zN-m�tK�&���ģA���E�T��c9�&�2G*�L_����v��[p@?�X�����3�u��sm�$i�	��fn"B5)d}4d��.P����� �,=�G���Ї���T!��c��J��?I�fe����^3[̣$'��I}ukK+�Z�7_�kG������q-Ҏp��r��3,����i��lK�i��V���!D�`���܃9K��Ԭ�]��.bk��D�4���ͱ�teB ýc����������
v��t�&M�s��W�L�1�Gs�!�;Hdh���&��o^:MW�����j[=�� ��ʓŋ�1���)+�6�b��"Q1�}���d/�{$��!5�����������C��_�C��z��ڠ�޸C�?<�vvJ���%�<��	:1�Q�v�ӭ����"�AW�2b-3(���?�{�hT�I+XSh��=^Y��C�2yu��=f�"��!��I�	�[b2�F	���$���'E-���gm
k�%����J{�j��Kq�(M�ѓQE/^C{?�~%��%����^,j������(�[�)/�7�����5�#�ɤ�����+��	ʝ�r.���b�R�6	!�s������VV� �>��U�R6�ު^�d�'U���0�15g��������0��"��֜>��7���{4�b+�iL_�N�I��m�</V��b#�k��{OM�s�OU�dq�R/91�)f�q���b	
��Io���z��]T��"͛r?j˝�C򕩧Am��V>�8hJP-Vle�ϓ����v7�.�!��
-�$�?��_���ϦY1����݆�2�����O�N��e�e��N5!i]x�J�Kp��:z�ʝ�� ���N�b�Q�W��PLܵ��t������8Q'Nu.p$�yRO?iT�N�w���-��$���	1�M�%�գ�܈�v��n �d؀rN���}b�JY'2I��������5]d՞�c��o�B~�rR��bYt���^7�q��$�шW�S�坸]�( 0����Ur�{�LN�4ڳ�}u�Oͩ�8ް1/���MP<&���]�c(	�r���y�V|�Lɔ�O�'���ԣ.!�}.J�Ğs��E�F�)���fZ��1�"��-q'h���g4z�D
���͘�ؐq�jr�S�[���TD���Q�n"�L�Ę�(���&�+d�����7�\A}"`��|zh5x4^a.�d�Q����$�T̐�.@�B$�(e��ܴ-9M��}O��ő�mv�X�=�AM �ij2�z�p�Q*���>"�f�O {0y�']q12��_�)	A``�G(#*M@hs��K�sC_��uhr�תX��o��#M� S�9�N�;�r$�c�=h�ۆ�b��s�������y<3�ԕ"��p\M���WW�%���䩯���K����yVk^��&O��M�)s޼�-v�1�K&�5V�'�9�탑m@���vE,�1Uj�"��Q��_�h��mO���=l�o�,4Z҅D�n�'�5q�U#�?�f��� jz@WW�5�^%��CA/�\�Q噸1��!���iux1MJ�{*�F��������5�q谜���r�y�	� !��֊L3��m�][���zG[d�⸂"��3���AY�ت�L�޳����֐��9=ᠷ����/]�l��"UnMQY-�\��Ý��h�۶�@�x���ڜr*�є��#�0A��e�D)(m�Qiv<�5(�ܴ�����!��X��ܳı���l������ż�P.S�ԞNې&����#��e�#(���3'dE�r+zwSt�Fq���<�G����4�#e�Jƥ������1�l!�;dT�a�A�JPM+�֛~�E"@%�~51����4�s�,G�JNf��9%�2.�e"ߓ?s_{���eg�[���Z�q�諶���9!��^+h�;�s����܉ ��J�J6i�n�R���Ĵ��RC4J�(RW
&.)�Aco��[[\��Ot���R��Kq�F�&������.���RcO�7m���{|,�iMk�4�@��3;>�/>�BW���>$vWVG\�V��V{e�ݛ[%�����;�'���M,�z�)����,nߋ��蹲\ �1�-R�/&������A���>V9ggg���ZZė"�7]��|�j�е���ޞ�)t��]�T�t7]��J����{�z�?y"F�6��[����d-��&�|b\?$��s��6.Mʦ�6�uRV G�%�9
S�%-a�<}*�ԯ����V����?����x�]ǈY��m�\��G���1��H�"�/C�_��d�궗M�%9��V�f+���.BB]X�ya�(h����Oऴ�-�<�Ao��
{d��Pjk�&搉O�"��힔��C��"R��E$�z�	���P6���A��Ƙظ%ֺ�;j_�;��Q�õĽ�D)�dAĐ0+�4�G�A'�I& ���kS�����l�AF2WD	J{�PK��R�X�~���n$�5�H���ȶ
&P!��M��N�l �@&���.�@�c}J�KyQ�ve/���T��>oic���/�P[��ZZ'J$�*�n�d�����7�sE�>Fȴ�/�!m��S�Ѡ�6&nާd蔇eJ�t�y��`�n�����K�4���l����ȣ���P�
�Jt?�p�<!��+��f�;|N�/�n#���dz�-l�}WR��,�S+� cF�!癉�"J�A���i.�_<�;����yGd2r�~,�N?J�.����}R*�˸�ox�U�%��?�kf
�3d������ח����\��b��dY(�('�Q�h1y���b�`{�����H�_����qC[>����p:�LGx�Mko_� ��`�����0 Ro'�ۣ�W{��:K��IѸsm�{�mI9q��\�`+�7�D؅��N��8�c9W����X�jj:�'K�8��\�8ս��%������28���EJ!m/spD���N�]9�#�h��B �XR�B�6z ���Tө��]i/\� ���H���Ju�yKQ��Z�>[LU�z��ww��B����܍c���<p�]�~OY�PZ��t^%5դ>Awp����ھ��_#��DQ�(�*%�m���K�i0d��NR���:�6����E�޷=��A��5��$b�d�:�i���Qb�e»�a��Fck���v;���G�,�C���������ߍU��q(K^�zj��ݧlE�l��V�!�X��D���Ŕ�r�%�q��[�>���Aԁu��F���iL�:�J_Kϯ+��e��c�p��o�Y�&kVz~Xٔ~6�{b��9�e�*� ��$F�*��c�ɾL�B��j�Ud�B Mf�P��,�������T s^���gz�";�PW]��ݭF��:wa�&���L+��byz�:��-A�8��4�����fH�3���8E�.���Vּ���.���P���G�Z�-�T�UFun�&�)X��ib\Z����&M0��V��+Qc��zCS��^�Fix�vI���Z�����_� ��cR��p6s�պ�X&P��n;b 6&�0�j�`��ֽ����Y��4LŲuw��G诠���D}O�Y���3=P�<�>�D9�o=;���]�w
�Bɭ�g�a��Ů��|m�^ mT$���M��`���B+$�y�Z��N����8�Ӣ�D���
��+ە���ʲ�cZ-P�Bt�?!�c��~��_�Ri�g�x,C3;}x�|q�v1E4C�D�))]I��]m�w�龜���ճ9x�[r%Dj��+�<%�������g�Q�� �!�\EW bh�)���'�3�0���s�%5�&u��8�X$�3��&��a����ڹ�5B"���!��bL��n��JH��µI�UѼ�
:�@i���IkI�W�]���-�vۇ(/���̺EkT���7EH��E	"�kϭ�%�.�1ݩ&统�.�"��<w�6��dq�J�P�t0R���B��&G&]�PjE�i��uE�U�.q���Ȣ�-U���d�:i���"�)v��"�N���r��R�ۗP�u�~�B%��!^&J�m�D�kϑ*5��AHE4���EۢA+���壮rZS��;ӵ�6�!���X'"*zpY���N�Y]��E
�4RsNZ�@s�%/��V�e��D�금���2XDSa���V,K��4�F�:,�pb�*g�Q�:s�;�����)Rwq���A����hH���X�,�BH��sZ�!�9+͆��Y�:1��EY�#�IP.	f��|u�{��Y��sW�:�F0�h��\�D��"m�l�kkZ����޷���ˊ0�������o�E k+�h�<�o-�Ҥ%�Ɯ�J��DR՚TMEYE����	�r���%E	4����	V(j�F᦬�@)�CR�C�^j�~���r*ְo�͌�+�t��\'�;�V]Y���
 �o���e�?��u��u}��ƞC��SC�ucr�9G�^3�J]S��9ZB�hI�k���+Y��R����	)�b��&���8�*�{�6�)���Z�"�%�d/PZ�z/(UI����}Q�Y��F����%�Rnׄx��0���>�&F�%���#�Zعףxx�o�����4[�������b�k��˜ๅ�Ooݾ<At+�6�yK��Ѓ�ǒt�
£�pND!��pl���#�{�!e�ܒ\�75�c�o�,D�$	���	��	TF�#��T'n���ҾYA]�]�+�<��`�L,$�#�)�S�vXBGy/�d�TlL�̭�1���[�_� ��/��%�
A�*���a��9��SFC.�o� �fxT����)V����M1=�Q{<zR[�5qd"�]�{ac��	�ݶ)�$;�a�|`�fO)�Do���&z���+�E�H#��2��DG���4�3��{ޱ��1O���1��N�5
g�S)�|��Wu5Y/��t����"��Ӟu�aMU�#3�<����J�Y�Ŗ(�m���Z$�KX��u��� ⱞ/���dƩ{"����S-�46�l�����F�X������:K͊��?��Y<h���;;;҇�L�[���x{������L���S&���y��k�R�Z!��ʔ��T��V�'�sKtS����2���  \&3��pauċe����R�5R�<%	=V��a޻5�4���ab\!%�d�
/C,�o)���Y�&���{���tG�B�oy�/���iT���}
.9a��Nis{�|>���j ��ZY�S?�}^��hm[DRz��A;݉�B��iV�,�!�mq��Zx�2�M���
��)�*��M5�55�Wj���b=QE�&x��0������4�p>�f @lQ�Y]� `F�!����i�³:#d�{lܳn��h�$m+��b���˓�i���zKn��=�+ :�v��Xb�GD�"����ln,��(����~X�D�*
D<@%�	Ć���z̍JO�跘�"�V��-a��֬����97�wl����J���O�I�=�x֎ħ}/vs�td5(U�|T�:���7<�x�+Dɟm���#m����<!�C�50�Ѧ���c���\�9 I���r�f�;%q�i���md��p8G��O ($�{������Q{1�)3u�yy��+�Bj|��n*Vs� ��#%�{��8E�+�R��3Z�=�&UC�Q2b����XB�M��wE�2�����C���B�]V꒽���.��,r�ֹңt#U�p�횑%L�ַ�Rb��?g#R�tsW�.%IW��S� ٛ��U#N���ĸ�5�>V�z�,�����5S�¿�an�{=&Q��y�׀����L�E
�6f���0xl
P���IoK;8
B,��a�;�;��F�Κg:Ry�������Y0s���[X��Q��=5��$���Bx�nAY��h����6"������|�O�TS�R)g i�歕$�;���g�g��A�:	!�-RMz�-L�'k�d�P�;��n�[ y������eg��碞��a��(�#[��3���z�[���(�	����\�*�S�����M�[`V1�*����*X		 �G%)���ZiU�BV"j^�%3����� ���'dc~�+v��s*�1�PT��S�򹕻^z�%Y@ ,�ޕ+��q�[u�M���^����MiZ����Қ;d���5��7&I�/�~�9dSڧ�X�t��Y�hQ�իW����Ф��}$s��ڂKW��u�����MV0��4�	⎑|0�!E��Z8�a��w�ޕ4"��]�C���D�lܹsG~o1DwX_�ښ�\���W��&_#ZL��]�4 �9::1A	�(1ܓ����F�ͭmz�[w�.�{M-=M�=�ٱ4��saB��s��*�@~���aR��N#}⚩��8/{ݚ(�i+W��1 L�������roND׉e�Q���r@k�s[�@�i"b��6U&B]W?� @6]T�Y|Q "��WJʹ�XY报�K�*�^��>
����ll1A*1'��Ʒ� �Q�G�>�=��%�LФu,�����Q���fUkO�ʈ��81{E� L��T\�F,���F�>_��{c�j�U���I�j��i7��s-u�P#hJ��,�b��"ؒ�V!�䁻l�W�#,Y�!ؖ|��(]IZ��w/�5Opt��M�6��1s��:H��^R�
#�%�l���摹��X.�[TH*�\ �����1��R�s'nח9��Mqz��
�>c��fE��FY�<���p,.�i�X�"g�;�3�I�\���!'��1G&����V���/�W�V�x�NV����N���w��ڜl��==~�>�ͯy�3M��:F�K�O��t�S��(絖�����,x���ɜ���d��_�|X F��@����da�?k=Ax�hj���c:>�j|��ĸ�(ocD�-ɝګn�y�JTs�`%�8��j4������Л��Z��1�������1x��!ȍ[�Y�n�/~��4�oK62���]J��cB�nW]������{�����a��J�`����E'h�ՙ�C�Ûm�^��sV�s�� ~��[.̭lM]�~����gƧ@�L�rH+���R���2M�r�)s�w^�~�?��?�#^4=/�/ܠ�����+���GW@,Z+����M:9:�V��MD�>����;�ߝ���P[�6���ɢK����7����Dod�� Ip'�}II�v��v[���7o�O�f��{��ݞv˶lY�d�I��I�b%P��]""U@r���� ��2##���~Ϣ�h�9ي59��e�g�&��wb�u�Qh�� �Zq�J
xN+"� �1��8��*��H!�%�D��r�R���>z�d��NS/\8��|2�+���������hp�0��E���/ƹO>�r�z�(��������	���ŋ�����a�eL�*�r#��Y��hPٖaG��0�G��֓���~�7kqq�&L����y�]g��.-�M���{ڤ�rUY.�߯�����z��h�ĆjF�S�4?����0��!���>�jr�x�9��8Lw�_�^�PB /��������҆Ԭ�����s	WS(W  ���9Ym1���5,��~&��FP��C�XpJ"��nq�uZ��Y��i6��o��>��'���'z��NVi���L�|�p������&?qs�`N3�;���E�����γ��ѣI��=�	�s�h~i�f�<���E#� \`��B��OQ/��@��^�B��B���dA"��%���Erњ�},��)-�j�0Ƹ�����2�=CI�J��.�@���.��G�%X�R�2��3'���>+]��6�������瞣�c��ڻv�'�S^~\����g�j)k榘��x�Q�C��a�#884��93;�N��J,��%�xtW�F�4a4�Nk�����N�k#�V�i�Տ6뎚�+�5����O��?��{A�����4�x��d�����w��{��?��v��M=�=�e�ڵ����^�}Ė��{��1�Ŷ�*=�ߙ���܀i��C}�Ƨ�-f�d5�U�������N�+�����#_��e�a���(y�k��\yWD_�+�����-��cw���AÚ�f�"Z���������n�"%l�B3$Y����1{XR�#Ti�}�jt��Y�M����g��ChFj�� ��8��$���I�F����`�B������]|�dyd
��Œr�uf�o햆a��y���(�3̼�\������O?��'�rI�GDu������B85&V�U�/+�3�W�
U�5I��/i��( �T+�����] �\A��ikg���K�M.)�pD��˨���U��8�\=�q��K�B���Zʢ��*�t|��8!�n�S�ɐ�rj������5�G�����ac��څ���R�$�U�$ɫe�		S�).*P#�4��VT��KF��N�����-kM�eq�)����%ԡʑ�|�D9����QHM�A�€�2m�)�~���8��$<X<��U6��͝��9�F���z���Ӷa�i�'��45H,�|�i0��E-q=���D�D�"0���ՂOl�B�u(	l�|�8�@�
���nG��&�y��;_XwlԦ\��]X��9&�o`��7od��]V��^��'B�C�P�2R-�����Y�L��˚��q���B�j�[d!݈]9�KW�*,���Oa;`E�ޱ_L��
�^5>,�֞߀sp�H�g�=�,Jk�W��Р��D-�lzw��!E!WPB5�ؾ�*/��!\�5Y���w�?��U��������X;���&�ѡ�A
�gee�������]�d�X8]��֦�����9���6=-���,���B���ڂ�i:��2��u�1�Z^$�P�,V �"|���G��:�y"�Q�����������Ӭ�"��	nȗE]��خ3G�mt��q�	
#U[V���ұGkBj��vy��#�~�$N�x��q�����Yj���/��E%oW�!ֽ��H���H+�iLt�N̳h���
!����3�E��G6ӆ�P,���i�I�j9�8��~p|E&  m����]!CG��[���m���8�p�L�4�����Or� G�����Z�
i�j4�!�hx�Ɉ���$l]'��/���0�԰k�ڻ��j1�a4��`��|_P2���`Hh6&�9�ɒ���R�7�˒��A~�:ߞ+LW�t.���1s������� fI�c���YB1�_v��{���Ώn$9 �%Ӣ�ܮi� �i{ؽ핶��HY���
et�I��dD�N�q�A�qن��'-���@S�"�K�yM�͛EU��������0���+-N|/sI����53i]���]�"����j��b
��*�lLV~��2	�ARu%��b)�Ȭ�è���d�Zk�l���5/GB��!9d���� Qo��BhC:��}k���EӞ�P��EDa�A8=hQ�_��)g0f�� E=!�ܹ ��=C\A��<�N	��"]�+���T$%��(�`o������(����_�e��9m\Vj�5��z$N�,F|�>��<,�E�����6��K�,ءiY j/��ժ9���KJ��;uXgg����B`���ϑ����'&fH���3���փd��tw{��K/yN��]@۲$k>�R݊�"Cl���%����?�Y�q��.�#`Ω��+������!�w�f��Y�wU5�,�/qQ��������^��,���B��̕�/Š�=t@�3�n +���\5?�S�r+�^B.S��ly�ZU��D�U���D�
�v���$���p��k��$Ysj��SE��;:�������	���H���&
&����m�S?a.���$�W��}��zS��� ���c.��Z�ȝ�,���l�l��/�\7l��dA���)��#�����9�\���o��cϖn��])��:p��������(H�	:�e��?s���\K�k����Τdu������K1{Q_v�ݿ�rB�����*#�t��%:x� ����)�UKi~`�n2�|Q��{N�i���`�+yv���h�)ԙU�'�&���\��W�<?>������Ú�/_��cw����49��f��x�qP�Z�+�*���db��.]po3z���t��޸Q!a��C[u;�<���S�������JKʮl!�$��Ƭ,Z����wY�v�b̦����J5�in/Nu��տ�_H�ur��T;�%�h���XN�*4���dOE1`$k|����^zd��*�֘7�Ѹ��P��|��ͱ�n�ɯ�W���,g�QL9�4Ѣ����WWo7o�+�H�Ǭ�D'�p�`l4-���*�kK:h�G׆��]Ix6rǥ��f�ן\$�?�u~�x���]d�[t��(
=���J��	2d-j/1�X�����^�(?Xb�7:�+��j`�l`SaK'�ͺ<�QLY��v��+�OE�߅��z�����n2/hz���2������$ѕ�L�k�(q>�]�vK�%y�V.V�u���kl,��&W���PC�!*_W�Dj���LU���0�|4�1���>�)*	Ts��$Kp��1Y֜�H@�&+��� �W��9��06;�,��#��C��mvx�"�'��Uo)T5Δ��˘�r���H�ʣin�~�ˬmKKO��=t)�-���]��2���B��=iЬ�]�s�$8�R�^J��a�a�(k<�v��]o�.����-_ n.{&�Jz3 Y���A
�&�����6�mYS��꽆I���<�d1�E%�BR[4�I����j2�Obc�Ʈ��IJ�?���Ү]�X�=,��϶{�µw��c��u�6�;>�������lָ�#y��)��	�L?����6=�xě6�7�x�����Iڰq�3.a6`)v��M[�l!k8��X�eE2� &ߛ�%�#�q�u�Q[�	6� gϞ�������jt;#�>u���۷o��~�;��������� ձ����>�cǎѩӧ衷�~�o��_z�/�z���xG��/~Ovz���T �‒��>��#��p�GE���g����g��K/�Gę������'�ҙ^�-#[�f�<�M{P��Y]ج�z��V��+t��Y�=-hh�v���IZn�pj0��,Mqq�N348D?��9���͛��G�������#���i�t=�8額6Ѿ�=t��k��χ|@�=ݴo�(gȿ�⋌�s���i��Z���U�|��YY?�b�JI�P.6SEYs����֘��-�z����?�W_{�����wߥ����F6aFK ��Ѣ�g���@���ԃ�T������s��;H��G'���_
r�2��v����C~�o�E�ԁXv�����=t�0�4n{�u�[��w��o��QƟ���̿%��ѧ�|�.��J�ڱ�)Nm�f7gERUQJ�4��ϕv�b�az������5�I��/~֡!ř����/��N,�چ��t$�S����S�Am�����͡�Ǐ'=O�J�7o�}��ѹs�h˶m�9�
vp��	�_�����s���m��U"{���
2
�
�s��K7T�r�l�yA[�B���2e������C� �����v��S�"m����NP�8�ȭ����०UIEp�����)�}��y���L;��e~NOO���,uuwyj�OW�\�l'-h�z{�����H��z��,F.n0�j	m����{о�@짻��2x 6]w�TQU(�I�yA�Ø���^REU�I�sne��`���Oa�
U.Ɯ���m^{2�N$�=s�$���w���@� ��{���'�-��4�*P�����m.|E{=uإ� �E���K]��/�uw����ίpם�y�ꏟ7n�'O�<ݻ{�nݺɔ���ghӦ��y��1ݢd�$��cF�p�Y�E=G,8���� dǃ���K���{��q�}�՗4t�_�#/�!c�絓K�.z��)匌lf�ו��8��٪����6JFS3~_+�9�3�3�5���C۽B�8�Ů=�,KX�+�"yEa�<k�����_�~�~��_��A�bR������;hl�6k-7o����!���OyF���-����s��~̀16Iy�\-#]#�rQfE���Ā�)ܭ� M�5�s!>���A{��e�%�!��KS���q�T'Gs�,{4��Яi)�P�
!Z$����6od����:~��xj �m�Zǩӧ���mT���~ސ&_��?����S 	��OU]�8��!Y��w�f)�lĵS�"�q�JTE�D�V��e��e�P��j �%���H��\���0�km� 
}�����-QĬ�JS"(v�\k2�n��d�r�_�4���(B9uF7�ȃ��@�+�!|�"/����2�'�h�p/�2@#[T�ꈦ�;{�e4Z�~!.�S��Z-</�����O��;f���7m����f�lg�j5�6I�_|����C��� �d��h)�y�;yW�M�����s�L�ݝZ2�$'�&��@�����U�K�s��J��8�T/q�0�)ҋ*���Z�\�H䚈�~��>4ˆ!�h��x��}.\���7䰷��r��?��&;D&@�|9��T�&�!�>$�E�a]�+�����/�c��v��;�Ax�F����qn��jav������0���[YX�����*�nݾ}����;\o���G���c~��U�(r���o:e5���$
M!����C^N";���lsMM]c2�5�RƵX�XWGIVEEC�)bgψu�k����I����N����4���<ݹ3Fw����~@;�����"�7�o�|���Af;_�݆ɇ���E����	��_���ݹK;��.�/�{^u��^�4z̅b{�A,�t$�w�����F�O�*�qȽ.oc8x����7K�$o���H	/fњ���"kjŬ�,pӌ���P�E�������5�|���S";�ɠ��?�ȿ>d���>���:w��x����k^Ki�w��)������ϝ=�Nǟ��=���df�~��3o�@��<2���������`LQ��c�'�ې���͛7Fcr�c���u1�B���"���ƍ�&��V��@��BhW��qFY�[���gS�7~�3j����;���K��ֵt�����~��nڲ��4��s��z���)���7o��m������B�0��/�B7�^��[�r��4$g[��u_�n�$�М m�BH뾧�`�����h��^�L������7�]����Jp��I���)L�d2J�����%l��o���xgw=E��Ӧ��ğ9y���Qֆ]�k�N�qld\D˿��2����ǏӡÇ�>��~�6n���wn�	
|(/?Qd���QCq�DƂ�ͧ������6C;	�`���cw�!�X3O�9Wmd�f&2k�!�/[zMC��%��su�@8�u�W[^�.����e�\�]/�g�|8A���
�\Ԃ}`]�7o�Bol{C<�^�?��~H6�t����ܽ^�E���I6L��{8��i(�F�jO�ր�ooϨ>L�p��f�\��QTl�|���B���ڮ klJ�?a��4�~fz�o
`�U踷��n����[�Վ��IZ����z�5�9W+��/9v���&�"�&*��V�Lu��Zxc� �y5qK|嵭+^�9z��ܿwOZ�utg��"J��*$����>���P+�4k�k84�T�SX���}�)�.��X	���������m0��X�1WC65i�����'�����"�,MXH�<$YC���-�W_�~�h�6S�����T�nV�2T�{Z�X�o�x���2&*���2�g8=�?�\��������޽k��%M#�K&[9���0�̇��5��q@	�t>˂�[OK���v����o��4=�����o��6!�Vh�Z�l�k#4���~�nr"	���G�a��\c"��R�+�6��I/�^�Nz� ��#P���*�u����1�'tP˭Qvg��i�JA�<�%8q>p�Uo�/�F�&q�"q�5��������O~��Ң��z]}�&B�N� ��<<4��ŉ{B�?�e��W_sh�TjWݠ�%uG����ʵ���o�����O����],V�v�`�uh�mރ5-�.Dp��Q%G�/Ӥ����o�O
jA&�
8��ޞ��D�~���f��_�e�������}�����u��2�A|��ȞG�yr�̗vHi{�d��)��ڗ��:��4k`�C{Z!�ր����K��gg=�Eܦ��ݻK�w��_@�Z������Qa�[�N�Zq☳�q�� H��Y��+WYӲ�+�
�:�8ǎ����}v��������χ��*c�ט�&�[�eg_�ܢ�/0�D�zZM"����)΃%�����w�~1ޜ;��\�B05����;�,�1L�ƍ�L�'���M�݊��J�%�{�Ȥ�	����9�-�L���|_$��ݣ�鋳�Ӆ�.��M#t��!Am����[��{2�����=}��m���9�?:J�����D�B���	�Sݾ��裿|@����y��W5�����m�m^��0�3�\�����\�o�h���JR]D;{�m�@37�Г�'M��^e{�W>�}�$c@^�����NÛ�Y;4ӣ�rע,:���xt�Y|�K5u�J��!�g�}ڳ�?��O��u�[�p�M{=��o�a��^�}��1:��__�|�;)��?�OI!�|��/��2�9s��{���w�66>μ�it���%S���k���V�~C�O.��R�X�X��}�嗂ܱ�ܡA]���9��j�� �iO�&�ݪjoPI�Xi�q�ׂk��@����cGyr���8�Y��{{z����{�( �0�� 0�H�54���2�P�� ���2{C(��_�/�en�%����]l�Fc�QЗj�����a��Q)Q�ӊ���#_��gZY�Z߂��mᨸ�%-&�D����sž8��3�h���t��ֹ�9�%C�<o�ĚϲjC�>����Ň����O�c{yY���f� v�����kfZ(J�Q�dq���i�J� '�bea�fc�Z	�Z�Â$�kշ�����m�
��(A@G���B=�)�:Ǣ	@+N�y���� ��]�K������bæZ���7�J����!�;&vg!Ӿ���e�0���������D�,(XW΅g��=R�c��*�̓�N|V��~Nm���%Y�/��.�99ět�7\�32yw�k:�8����dJ�cc�MH��N
�@��P��g����T��Ɓ_i�[����jKag��J��H7��hra���3�k�>��m'Mb(/��,���^Z���eE�gŞ�U��G&�M7�J�X�K9W�Z,�-�ھT㴧9\lBw¢j�~Vxr]�|��J.)������);)��3��+ �K��)�8��'�^c����#���;c��M�D �ˎgAG�-}2-��Y'F�a��ԭ��֦��Ԗz�6&v������m�����HpU�A�,�u�����=^�d���y��"��=ӡ�}��@+M�Ak����H��a�p�>�%�Op ����[t���R棰�*�o��oi~n�)�c�s������eUAyxN�x�y�������Bej���.f]0�bᚻNTe���`����ʍVt��Q*�в����~�������B����^�j*$(C@~��g��1v/�cX�09r�8����|��e��Oz�	/��\�,���C����F:w�K?�3�Oڹ����u!s^@���Ů\��.�_�����ի��}���?�|9�ة'Sls�ٯ^��ss��-ڻ{/U�# ZЪ�b�8KkYgn�`���QXNo�l��e���jb�E:0�@��XE& ��������1��[�h�Ν422�I�G���v4���/x[����L�X���N1�!�*�%:XfU����\��E�hHSy��6��-[����,C^z�ea��`Ŀ��ijz���'G����dq��)Oy78�6�1@��%�'��5���jY�@QW6�IL>c��9��������l�tQEz��w����Z�|��n�'����E��.��o���2x�_ë��4�{��5Us]p���$�0��ǎq�-v�qOa����IW���#���~�o�����~���M����7������l�\�|��8@��s	�����~�c<e�L��"/+�F���'��`O�Zx��YKi���{Y�<�Z�~r�߱�qx��򀅸�')���&W0vɵ�$��W�6u=u�BA�H����Պ
�LUk��*�=�R^=��/�SX)�9r�nx*x����a�ݼy��ul4���:��i���rd]����P[��XU����,�J䩋ř�C�%�u2�P5.�����-[�2+飮B��EvgC�ƮDY\���[��١R		��{��7LMX��?��'�Y�XU���b[`,H��OP�YƑ_ⱌ���q�U�s!�po$�W�������\�%a�R��fk 3��j��� M sa���(��t�P��70�g�y��>�<����ܫ�+//�x���y�+��������� ��];w��/β|8v�hJN:�U�J�5�����Ԧ-Q���"3�Z/_���d����:�j������6m����g?�g�z��������,�0�S4����p��֭�ͫeB����K��u�Y1z�����Jc-����CL��<߇�?7;�ٍ��|oݶ5� "lZ�d�?�݌�2�;��< 7Ck��y<<.H��I��7�������_�С�L-X����Zӧ�}��xP2����� \�$��Rn�c{~�b�=£܃��SQT�� ��;����0?oV�.p+h#��u��	��燠 I���B-b��j�Z�+8%��\�f��VW%�\xhnu���g�xr&yd���߈���Ѕ+"+.Ĳ��H�~��Ƶ�t��>.��>w�4��w�`���=}��� �x3撤�wߨW��cd4K[�GGf#Bi�Jj6L@�A_Y v*�X�]r؋I�������3�p�pO�0q��?Y��Y�p���=qf���"����i��!���k�\j�Sɪ�?���e)��#[6o0���X�ͣ��&��G��"I�J���o� 	itV��T���X����Tė���֖kI���,[w�s��o���i.q���ơTP��-����iE'3h�cnS��?��U�}��^ظꇫ(�^OjOk
!s���W掗�@%K������.����!��#
�sp�(C5o���ũ)~��͒m#-ԅ�]iޗ!q�S3L~��#3x)����s��.��cv�4�������Vm%ѩi��5�u��G�]w�LY\0��-![R�q!�~Nn����hKH�a&;;��6xȐND��\��/=_2����`K-�Poi\���"�o�lJ��;�
�����!��T����6N�F~i�v�J��e^m�\o�]a�"�O���񺍎"쨕.}�'\�3D���ua��B[���7k��B~��R��^���n�V2����7X�
{a!>����ߥ�Ϟf�B�·��sg�l2�3$���[L�K-

���N7�����!�/��3�;C?�Ꮘ��d�MC&
V`ݢ49�V��4@`f7�b�_��hc��Sc����.�&¬��Os�|�����{���\QhEo���(���%�r�@�-�oE�m�Y.=zC�K'���s��L��8���\�;t�Bb{	`�Nٞ���T�$eR&K
��As�d�����cm���N˟��U�z�Cf<]~�5���%r�%Ub��5	�����������G�A����j�4�\Zf���pI�u���v��o�ݻ}�ݟ`�ڱ�S�����?�E�8::Jސ��W�3|�W3H�޼�a��uղ'&�֭[��I������1���t#��ꭄ92�fV�+�.\�C�}�;�BV.�:}R����X�Uo-�Z��[�S���
e*�#��JN~ږq�L?5=C~�O��5��d��f߁����&����nߺ�^���;|�#w�:�|�k�͚^���_~��=̮��µrg|�~����k�����PN�'��Dj*�Nׯ^����M��ũwZ0Id"�j�֩����q*<e;�Я!���xTR��B�.yæ���	����,HB)Ɵ�����@���i���/�,����}�u��r�gtI���Ob�!�g��B�A�5�駟���A
�"T@m��<�T4L|]m�v���Л}�Ν���|L���d��@�1j�&-Ɯ�����nݸI;�m�>��j�3�X&��g���'��S��_ˡg�$w#���A��~�,�*���V0��Wj�7m����B[�|o� R����h��[��՛�X������{@��>�A�L�T�o��o�;<̊e�uT�>$$���; ,]<XT�^�z�:���S���
=r���6蛒QO/|F?��/���ѿ��_���@L�
ˇB��/~�Kz���-}�c����B�(C���ߢ��^��S������t��U�$��i�s� �Ξ[�j�������*�r�S��3�Qg�j���zA̢�E��{xdM�W��PW'u��^�����U[�h�����EޑHzˊ"hQp�c��9�8�E�
o��`��.����&���K������H�<�<7�Tշ��p o�Hp�#�`�ܙ�w�ʹ\���&'����`�9UL����K���S�rÿ/��r��3�G�l��%JG�M����5-Q�`Y�=���v�8F�"=�°�����	7p4o/�␥�H�4�f߾��E}-����cw蓏?�O<{X
b��m�z�}�9)�l	^^8-9�N�kז�WS�1\�Y��I���6�,\��XOEdb�S�����*���Y��@gY�F����Y��2JJG��7r�w��Ӳk>�.#߰����/�ݝ���Ǟ�_�"~�
fP����?O��ߡU�������/=��^S��إ�g�(OҩS'�_�.,�sq��=p�*	��z�]�tQUu�c
@k�E���HN�g�7~�����G�ywpXMQ�%!3G��~����"�������H*�$�%�/�R�Iq^��� ��A��S}-3�
2g�q��	MH�������5U:zh��CԷuͣ�tq��<�k��%\���.�����z�嗘� U��4?���h����-���z������=���rΟ����2������6 ��ǎr��G���<(��S��� ?���Ƚʾ��~���� k������K��8%ɿ9���Ȗ��������]{uM�t��I�_QC4�׈�$.vB/�P.`vպ����4t��q����A}��	Id �������
=w�Y��<��~z��W��z��	pW�v` I�Ѽ�o�៨��L��Y��i�&����W���#�T\��;�C�G�'v�������=�M�F����RZl&��>*�7�6
j06ѕ���O��Sߙ�0��в��4�Ή1�7�PJ��P�R�r�7��4"~rQ�Ɯ���,���jh���~�#���Ѯ�հ�2�LLK�����fc��4l���$�B�J XK���F�"Sj��M���
rF��Y�xR׍�s�Aj���L�U�^�rx��Aj�d=(��8﷢����:5�k��X��U���J��x7IN��LPwc1kd��������,ߦEv�\�|p"����ŉIFB��	^i7C.E+��(��ؕ��m��}���Y�3ۊ�i�~��M�Fq%����C͚��S�IŸ�>����s�Ʉ��?��st�����vhoCk {&�1q��Z����LYD�P�g�Peն��av�
f/&~��Xk'Rg��ou��m,KW��d�\b�:x�T�H�*��/�%k-�Ү�B�I��hWJ�y͢�y؍�-/�UL	�nᕭ�T[\��$��J����J���������-�^�s���nb���p���)�-H�eDC�2~KJp
t�>fl�+Xۼp��mK��4�����$�w���d�b�\"K����8N�{6���|��K�����,�SG��d��t���"L���X��x��g0y���@:�� �d-
H�J���c\� �VFꊕ�ڬ��X��wJ��5��&�T��hbG� �L����vgdg����8Ν�\&)'jJ���!�y)m�?�n��
�ڜE[!��
�p�N]�1���~���K>c���T�N��K	k2�UT�-8�J��3�c�Cy"�&!}ؒ�6�B(��D0/n0�E��6�c����łv��.m<q���j� 4��i�X�9�R~/�U?��]��(��0D�-ZB�󳼀�S�8L��XM^�
��@[1�#��ΉI�J�(�"&�5�dQ"��S�UJs�Z���pD�V����N�<����T�&#�6�?�� U6v�j�͡5Hj��U=���_w��eq;��69��n�!Ι�!�9�/-d-/5:q�&b�����i	�ik$�f)߇i&����-���Q���4%�s�5^[;��n���p�G
G���f u�wv�S>��o���D�j"�]��
yHI�bE'4��&�M��6�AbM%,Q>����"�h`�i�Ѫ�P^B��e�Qɂ�A~~�JI��lٜب�xp��W9#�3���>���a��m���|�h���!��QC2�U�f�:Z�T:Q�#����N�+6Pr]�9
��c�\uf,'l�ɭZ�E'7��79�r�!�^*��"��Z�E�L�#e�_��s�]��i��u R�9-%g�\v�]�&��cEk�(��-K#+̹TV`�$N�5Y&6
:�ӝ�j��A�6^���Pm�B�,��,AR]��4[YJM+X�y(h�+�A�CN��(˛D/��I<�haSu����*�� ��N�1;�?�$����S:����?_��=Vequ?�r�-�������7s�u��49��z��u�s�V��b�����3늇���e�Y�:xJ�b�ֆX��Ɣ��!R}�X� �ǵr�B�f��ԛ�jz��9�V��|���Lf�f������i�j�ֶ �
ʋ�� B���n2��XŦ�ӭ`%��~�#RwQ�d���]����N�J���QH+m$0(U�[/ɷ�ڮI�i�vO�-�n�Q�N����N��o4�i�M�"��(�ޕ�����|�W!�u/Hr{�Iȴ̝�p���5R?��Q�JVA�%����&P���<��E8/�;�N.�k�!h�в΍�rsԭ8c� ����.R˛̈ҿ�m��Vy(�L�HR�0��N���Uۺ���Ӣ�3���m0L쯡`����.��U��Hɔgf�����gŘ�$L�_�h�cZ���)9���\�c�-�L���x�־�p��n�Őƕ��RP(iH��?Z��E�z"ף~��)	�u�S��E^�a(���ҪΝ�Q���SIv�Y���ť&�i4��5����}���b�4n�Fw*ݧɇk�A�j)�$!s.��E�����{�v΋b�S�����6��'�S�j|����
'l:q�( ّ��:������X��^Du��~�zv�ד#��G��[��RN*�wd��X�b�	�[� E�w\݂�m���G�R�JY��,K�	V��cmϾv�b:c �.Q&Δ���jr��-�-Fa;���,���6�����LTέ�06nC\�VC<2�<*7�΃�a����"� �$�[ӚG<��[4�5 [ˊ���3kç�W���a3k��*�̓<z�8��
��07{L��!�lĆE)�Ar;G!摖mފ)&�}'�"��&�Uȧ�;��o�om��k�Fa�?�R'���wc�D؊B=%I`��=3K@�$6���^��yHI��ՙ��@͵�tK���z�jV��b�N��m�ූ��a��zHD���ʣ�3Q������	��dP�yv�T�M?���%�G�0������6����QL�0�Z8��1�{���o�T?[�+w]��:��*�*\P]K*��WX�A���>#}HvZ����H�K�\�JklsI�Q��.�o]���k��x��,�~n�d���@:�M&��D	s��V�)8U�<PQ�e��Y�(�R�M�$jY���꾓F�5��ߦ�d���Z��R=Q��5�A�$��.\0�
�d��Z������eH²���Vy�i��X���u�0f+zMM�I�Ǻ����`�T��A�֔x��Y��(k��x�6��vG(���F�F-���E���:� ��Ag�0����uj
]��p����{�ɑ��ٙ!�S�2'�E0�jR��yh��'��P��� m>�oc�A���G�;�2��	�F���BYLN��B穠�T=8��{r�1ת�C�3v�6n`�ށ~�R�iWV~P�s��ȵ��ay�gp�����
����ѣ���������--,���0�!���{2��rZ!�%��Ѽ1�z;��cw��2���RP���;O�f�3'?Q�	ۇ�id�F���o��/�BP�=8����8F[�m\���@���%y�-8XQآ���T4q	3Iw`-�P��>� ,�L��g�qy6�pQ��c�.F#b6��Ď%�s.�se��y��ˊqf�E����ׅ�S�����皾��>?Fg�����Ο;��0�pP@��Lp
4�G�(�O���`��K\�qp0�oE��M<x�`�������8��8�h����wfj��͇7n�[�oч�ŏ�,�y����!GA!A%Z���ku�����B�e?���k�-�'O�`W@�h��^:u�U�n����4����`��]�˾�ט|��Y�>�?qo�F�졮�^���v(��%Y1~�7`�1 ՠ{��}t�������mz�]���E�փ*�ȿ�������
�����^y�Uz��3|���F1�z�"��)-����L�
�j��`�ܴ��+���;��Z����j�D��̝j��W����s����� 
��e��0�(������Dn��� @�uPpO Fp��%����Mbj�'�ט�l2`v�D{p�����������&���������0t�%F�
w�i�t�g�[Q���!��-J$��N�\�wa~���߸q��Z�q�� ]�t��:�u��Kw�*m![��S��%A�����ڕ��������366�]FF6�=���넙�.�ĵ�1�r
��_`�@":�Y�_�{������@�&�����vڳ/�z9��Ǟ������&@یL7X�&a���k]�NT��e^�)�.?=�`�߾9Ʋ%\�`��6�lt<,XX��rg|�*�H���橢�Q<���#�<Tp���G�R]o�׏<�I��勗����ڶbq�?{����w u���ԓiOM���+�(�Yi���VN�~y��<���G�n-�"��f��;�;.���р�azy���)@] Z����kO���b���w�.����l�����=����ԦM���_�����^}�5������k��n���&�˵"ԁ�R7�r�f�ܼz�j5�������t��uuv0�D�l��NVB�3�aPo�U).���5�-�4��H;���E����M~A:�����3?�w��aO��X����Ȓ�L��e����釬�c��
���]�L{FGQ�����y��b�H�z�c���k���o�}M>~�؈��?�b����Nf3����?��^=�����P�^D�1k�~" "P��M[���$w��|��l���v���Dz�t��]��1^��J��G,����_P��L0����q��Ӕ�O�0��m����1��&�6��c�:���7 =5�� 	(�%O���'H�	��	#��4<<����~�@��[��-?�c��0�	�Z''����]��;ζ�*{�rS�f�8��PVg�Mi��<P&�T�]�
H��6(��@�h��T[��kv�W�o���|�kzݬ���@ol<�Yjж����\�ԹjUe�kV{)a|d�Z�7��A�zp�>?Z=<��3�|��6"��a�`��?:F	�����pL����
|�-g(�^x�;�|��Ǭ	�����]%�s��d7�W�=�A��=�F)�+T�./�&�-Pk�@�X�-R��@-�� π�����=sP-�aSU�sA+쁁K�s�S$y��4��"�Ф8u����@q'�e����	�=L��ݧ��ׇ|�Ͳ�ْ��Y�2�;v f�8h�h�=�Gِ<r���h�� m�8���M������~����;6�Xo5}�f�P(Paq&���DP�{=�V4:<(�{ Rl
 ��.��+X����lP�q>�V�A]��|zb"�U�d�xYE���ĝ6���C>�V���\h3
����؁`Uv-C VD�c��Y��O�����v@���2�d��I1������"yM��c�>�S�������A����^�*i���r��>4f1D����î�:���񋰸$(v�G�~���:�Y�t彁��Ѝn%_�T���(��Tݵ��"��XV��;���� ����>�1�r`M�(( �����۹Q�]�K�^!�x�O�4�ۿ�SI?��_��R5���P|�]�3�D�e�P!���V�O_��Nx�㚗a�<�lP�����gՊ`+�5==���]��ĳ�<�I7Ri��EhNi=Z�ֺ fQ��a��7���� ����nO�PC��i«���Җ��x�w{{j��~.�$	�� ��N�����'���7fh��m��~��_ѠW�a|�c��-5��Z����\����-���<��Ը��S�T`�� ���Xx�:�?�����<c���,�7&�]� �Y�.��'����yԒXV�*[&��YGN��9 �xk�r�˒[^f ��ĉ��fp���2U�6q���|+~������2o�^,��̔�����=��۳a�qv%^��߽O�K;��|�G[��G�i�N�n��d�	���`M�~�OO1�&y��~U]=]�-����C�5�� c�A	/pM�pekW�_���]���Y���-8���,��G6Ӹ��!@/_�L�~��ݿ�w6�U�mصೋ�{��	���E�����gOpU<Y���c�,,+���$��ħ�4�
8�v�
�5y�������mݶ��}�9��[o�W���$��q���`
�Z� �w���=˪7Tn�%�>/�7P<(���;�Y�	\��4��/Hr�Y��]'�c��]�ʞ�s���o���;�-����������� Gh�[��<���I�Ȃu`��)pG�nc �$��\@W!�ѣ���]N��׹G=���W����^mF����?p�
��/��u�=���_ee�7F!�aM��A)��J:�`�q/��*#I�k.EMjY5�+Q�"�P4�Kj��L�����t��s~'-x���wӹϿ�ݽ}��t���bڳ`��z!��'�p?C�1�l���l������.ܺc'��K^մM�Ij�
�
Kl��_�p�S�j��]��9ׯ]g,�-ޮ������}�?4�<��M0�	o'!�������HP,Ӫp���������o­��x��:����s���{dh�0�>��)|Z���:��Y�?F�lea���N��72����(��a)wV=O�Aj��-�p��Q�4��:=B�\7�<dA�&YfHW
�y~��ȃ\:x�}��gt���^��o�ځ��T]�,���K�8/�����l�"�^˗��~Q�zJC_Gg;�[�����
n�6�(N��Q��W-����=���P&�i�8�'r`�l����vE��y�0_~�p�#�_e�����$�g�-�*�8�����7� �{�b�l��w쐟�N/s��\�c�!R�l\�vY���1A����%/&i�ˈ{���}=������t�S�j����s�<���	�q���E_���h ��!��c��%A|w;$9bh���;�n���$��^/KF��g �ە6�� mdiq�n>��w��# �؞�<xP��A������mF�_�C?�w��t�b�
0�XVX'�p)��0I�5`�m�~����r�+p������/�8�x�G��ܾq�Qc�ܴ����m���]@�|8,w����]A5䚸�\��,��Jg7�T���ϣ��=48LK;���=4�_����lᇎ'A?��^�#�)^V�^?q���EU����lgW~V���FX��q���2�������wqם� ��Q�M]Q�k�S^�aQ�a���J��{������D�������v��v��F�����(�)@b����F�	i:U�mY�/���'���1;	��@לo�!e�=v��GxbA5�=<9�Q!ɡTj��莃�����������Dlĸ8"C:x�繟�<���f�,в��sO�3lz*,�G�Zˢ�� ��]��Ӂb���U^���9x��u�W
��ɚ
vRV��Ѕ�n�̶$UfI])Y�,
"s�^G���v��_��2n���5������O�"��� b�Da\6V�h���eԓ�*,-��"򤽍툁���� `Q����q����lȘV� ���n��<ec�శ�a�J�[�XP�&u��hL�36p|���<,���p,DGO�'�o�O�"�5�z�����|��-SW�6��YE՞�p������~��� Vѝ��װ��ׁ��
kX^`s#��Bv`*P�=�m���H$��pl�ވ�rd8�K��2l
�)lBll�Я�iQ�J~��,˚��*�H�I�CfY|���#�U��݈��8ǲd�YV�^P�1���B�eg��?Ь��< ۰���O���=b�Mh`pC��������kI����d>�����,\����͔֡��l��e�мi�~�XR��dʚ.N�����0œ5�_E�z�/k-��������݊ICpd��Y�v5������q�*ٔ�9I�����nP���|�-�� o83��Axs�OP&��-/זⰡ��	P���PSbzy�:�K���뚼�c]��M��i}q��� �=l\���~��rA��q��Y����Ⱡ�P�Q���D����2�1���&+�L�
c�DP��m{L8�rq��j�!��(�+����v9/ת+Z�̨?V�:!�ׅp�m�"�]�Z�f��m�vpÀ~�L)�5M279_5�J�[	!����������#Ƌm�-W>��%k�W�,�Q��0b=��Dw��0LA�KXJ��ĸ�����7W��W��2mՑi�bE�^�T��-��Z�|\
�N7h.��p�O.:>'2kƣ��%d��������E�C�j��/T���̩��T(���1�X�Κf�;�<��ܢ�U����ֺ�mw��$)�+�����$'*0n�&@ƕ�_^R| �j�j*E���\�����x��4�F/�-'�&I�9�Xw��O��)�.�
QQ�_&�/�����5���Թ�Lz�c�a�&k�\�+�[Q� |ε�E}�:*ժm<!	��4}�T6��F)u������&�����ygU���b��z����� oI�]��۠�O���X�B��.nv�h_�]��8�����}:OZ��le#b����Ws_�''k�b��8~p���LvgK˜��b�`���$m-����NŅ�pB'9ˬ�(����9DVp(�@�I�m��k_}x��P�$�\S���E0�¨��Bh1�]�U�����QќZI-J������h���L6�ǯ㢁��E�Mg��f(,���r-%K7�z�<S^G'���ː�e]��%g�"<�xeY��b��]m��f��.t����Ƈ�Q.G���(�^��Rt+nDE!��48cG������!έ�i�u\s�h��nWp�xM�EP�;'��$�=��'$$���g��.hN�y��E�4�"�4�����J�i`�� &F@iva��+��b�3����u�����#�2X�jG�3�Tcrs�Hh/�0t�UQ����H�Zc�\�QG=��Aǜz}��$J��	�t|�2i�lx��H5Q�4m���Wctk���`�|U._�
���l��YW���(\�w�Q��;�(o�X�hlL������A�(y0xX�߫o���X��5ːT�;�/g�{v�d7���6�0�n
�奧�y[Qe����$�i�P���O>x|cJ�-J�Qk��cu;D5���-���m��\,�@��|e�Ч�,��G����0j�V�\I>[�����6�� �˵ؙ�H�3�g6f�<�R�Q�/KǓ�A���b��μ,�Er��)�5��T��֠jy�̡�r�� �N+i-��< 6��l�D#K�Z�%���9+�W�J%K�S�bzݕ*oLf�y�R_]V�.��WP��2>�^�,��xHq;Pj&�y����`Y%:��+4/�+NH�����2�D�����'m瞋~*#-+3��e�6�E��RO�:$��x���Z����Cxk��I�vv��B[g[nm^�zU�֬�R��"�� q��:K�4-R���$&��r��%-��2/~�����$��^���J�BNo�C���fN��v�	����8y�����kxR: #|+����@�'AN�VT�K*����a�;Q�MvvQ��@����a�R&系FUl���K�k��P�0tQ�P���.HGG�D�_Qг�E�v�s�@���i�i�uƘY-�]h�]H������~�-�jg��&���,����0.S͸�{�\2���3��Bn���p�M/.�Ȍ[�����5a��6�y�tf+�8C-9����-*`O�����Q��\�L��"���^[��[]!���W�O���-$��Oh����M2�@�"h]�L�.����V�2d�[)y�X�c��m���Y`�\�)�e���K2�/�Eܻ0���ιv�4څ��?�_Yc/Y�œ�K(�YR0�
˒���	N�U-D�qc��b��Xb��md�V�KfoFh�л0����-L�W���)� �Pkaj�3���������g{�w$�@Sv*t3�yY)��Ei<Īz�-�i�pQP(V4-���p����K�FZ�U���k�	�IpM�(��ge����FG��
����m>���l%�[}w������s�8�"r8�n�B�4S���&�7G��[�e���6�����p��he��0FMWYE�k\Ҷ�t�|�%��Q|�����*crk�4+/,��r�Dҫ~�ʻ����q�N�7��l�G�Q�.np��t_���K��vvI�6��wF�����Z��v�5���1�^��2    IEND�B`�PK
     #{dZ?�>�oH  oH  /   images/a038ca8d-f9eb-4e93-ad0b-b831193aa106.png�PNG

   IHDR   �  c   ��T   	pHYs  �  ��+   tEXtSoftware Adobe ImageReadyq�e<  G�IDATx��{�W}篌�-͐�_�K<aF�	�!���2��,�v��?vON<J��s��X!�c�l��q�g7ɑΆ�eA4�+a$LV^�0Y4��H`$�&X�H[�����.UU���n�����>��3�]Su?������BCi
C�
C�
C�
C��Da^���|y�!�3���̙�D_L�0�h�\�}�)!
(!
(!
(!
��,_�<|R����G�4%���wB��Ȉq+!��!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!DAi�Y����s���fj�H�U����?�[�I"���ĉfd�n�u�CH��R0::j-H��V�q�&���!YQJa֬2;w�2���aj�UnHV�R�͛7�� �f�����*�rH�A�ƍ͞={!�RJa�=j�l�b����W<�	@H+�R����wlxx8hÌ��mڴ1xmY�c3��QJa4�w��t4|pl��J��۷oG�t ���B�����n2�c3��BH3�^�c�vs�u�����B�t�0�f�،t �-344� ��#�v ��7m��o��1� � ���:�>��]��F�(a����%1��u�������k���Q�[��aZ��ߐ����pWؽ��{fH�t�0 ]�2���h�Ha ��H �!�:V���AL�gi��T�fvQ�0-F����{��F(�0(�)4��1Eƾ}�3�I�����ne�(���<�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�((�0X�k,W�����`���^n�����tQ٧�F��w�����4<e3��Hye��A
�ym�U�STJ��H�&�^�ϲm�h�wM��a�>\d���Y̝����-C4��`����300h6l.|�TXap�$�t�fɒ�ٯKj^?|���׉��ƾ�X���ā ���U@rn��ǎ�cǏ��V�j������{�k$����WD
'
����cEY�x�Y�r�Y��>Od�G�O��2�'&̾}����7���`����6.�b��P��K���ua�}����̓�
��Zs�e����|�>�!H��#x@lzU��z#�<�DB-e��s�����n[{!��j��A��c����G��`���_ֽep^e�i�װ�D�8P��<�,`������W�B�4�f����3\!�A���\u^���ݾH� ���3\\��S���}�RfwI1G%�jխ�E��s�h$2�Z�H�;|��L�~�����T>U�*#$���'N��wܑ�v� �=�]��c�\ǲh����e������Nmq>Q��(6"F\[�R�����Ê�DqTFG�N������ka�dA-�SSS�,aڶh�yx��c�1Y��󊨂��L��N��hHm���5\��=掠2�h��lz�f�#����]ԏ��������@�{�/����mՂdK���
����Ƶ_ B���$�o��!���c�S��p^}�Ka$��M�o�H�v���ip�����J�mHIҰ�)�4��u�/��v� K��Eژ	���8��V�/������эtD�A��}�N4 �Z*�o?d��A:pq1��{ר���~9�_nQ�?��9eօo)�W��X��4�ѮJW ��,�!M\\���Eͽ|�oS3���WT��^�z�w�=���
�<I}���+a��H~����P���g�\�z� �G׮�^\H_�\��z�m�4���Z �!*�����Ho�MvqjY "Ktl'N��SB R'�<�I헃&N��Ge
�{lڴ���aO�@Z�G��YY�5��]m�`ִoQ�>�(�Y�׸�KҨ�H- ���}� �B�b/DC�Z�E����pa}�Վ.��^���g�~�Ad�y�{�(�����=yD��d8�mAZ&m�jC���Θ�LT�m�$��i���0h� ��!��B�))dyQ��R�+5qq}Ǝ.�o�8�$�_*�aZm'-���@>e�4ۍ'�̥c���
� �'"�T������~Y�Q\$A�A{n�-�\�[�� �@~
cL��r��f #e��c��,@jTI�PP�=1���X�����~�o-���e�޶c��EeAdA�1�,e�~��0�yͪ I�D���~ �=��k��|�J�ŋg��"ұ��SY��+$¤�3�v����&E������JԾ�ㅱW�5a^��+���RX�2�Ğ��}:v~���t�f��2&s��I�n�.�+�d]([�6rg��ƶ_&�m�vE499a�Mۅ�/lVS6�]�w�4_��d9�(����Ʈ�a�9�^�ViT|��:@��I�%��0�Iۅ��x��W+�M=Y0QRd�ws�'����t���va��*=:ǎ�&�,�'n��"ei���K�=d�^��.LV ��Ŭ,>w�,��v�,�]X;r��"�Mj��2��G�����`������e� n�k#��x�!�/�r���#wV2ǵ_��Ο���=W}���m��������c��Ap�ȑ�s�=�n����č�n�0�D��,B�j�i�"��ݗ#�2�B���l��}���Oaj
ױ�{,ɷ}�EF��l&�n��*#� ��mYM��>nDL�3.���}��0>�R��}��v�l'��L���r�Q\�%���QЙ ,�d�/��""̾���u��-Q|�ȝ� ���
��t�&���[�va��kn������|�ap�"n���j���w��s�tl`��NpÕ�u�s���pR�%���6�����1^�����>�{�y��b��pK�������\T�>�hZ�cmf�\R���t~�>�>�i)x!���"j3H �iB�S|�ܫ!��o����$@t�l�$ĥ^����yEe���;ʠ���|��e��"~ ������Hw�6�D3V���~q4�����0 ��ls�s�P��&�g�9668��-[��ۇ T@v�n�����t~�ϫW &A�*�5�*&q�c�7��U�%
�Vx��<��-Z�PaOJ�\L��u���z%�IB�t3c�%�d��RD��I`����a� ��w_C�/.�r1FvO�%��y�N�g�C�櫸�(�󃋊�ݲD/*z����jj�Wl�d��z�1���Q��^�}�>�08a�D�b�'����7AVYV�qϞ=��T,
j�;�W{��&n�%���r�y�yD/�C����t�2��,0����pe��!ݕ�Hصkׇ��D�4q�,��K�`����y�V���b�-�Dp�R�1M(�,�Ȯ��pO�I����Ep�~�t8�v_�0_�%�0@�A��=���V�8눃����]s��)M�e�-��Kz���E�[�֮�]<n�Xk����-(R%�0 '�СC�^��5��h�ɚ�-��8I� �f�.P��H�Еo�Z������A���Ks��ej�=�QY�r^!�F6��� Bf,�8����k�gw�=Ԭq���'��~��,(����G��h@΅�̬v:?�+"���DJ�C�蒷)�0
.v,F��l�k��,:�#���f�E���k�����W�Ư(�������]���?�h8��^�Y�xͶǎUV�YT�I m�miw�b�F��x^'���nwق8����ֆ�۞Q 
ҕ�f����|8�����Һ�'챴�o�K�S7��PHa��(0.9��R\l�^"((x���+A��U�|`�<��%�k��X�^����*���ސk�&Ƀ���.�wc���'��k��G�:��w�[����Oi��""����X��XB\@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ�fdd$|҉0�����@-�[o6o�m����y�^`.��#����W<^y�<s�ET�y�K��x\p�)��y��k����r�gf�9=sּ4sμt�\�\g����_<sּ8y|��f��>��a0����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������8��_=h=?P�����I#���xײ�߿��K���/�2׿�/|� x�淾͐l�0J���o�S�N�'�9i��ߟ<i���Q�T�Ț�@ڟ����1W��'���@��]����u��g�q(L(�O�����
��ȃ��c��ϝ�sH���;�fKC����sr>/Dx�[�"�?�o�_�QX1�Q<����
� ��P7�{�y�[ V��d:N�/���"H�H<�����=�kQ�:-�Z�5 EU�ٚ�4O�D�����2G��	��/|���R:<��?������i�Dᅩ�V����%�#*R�_[��P����]Ha$�<����@/"�L���u�}
!�"���_�<�"h��kY��mo��%�; �ߞO��� ������x'ҭ�|��(I�k.�}�o}�*�Ox!�����t� �<����w��E�Aۄ�;�-�;I�N��a��?F���4.wa�r�fAź��	�:��䝲�"�������O���>FBZE�;�4��C1�y��W_y���u*��?<j�T(!.@Թ���>�կ�ܶ�w�/����>ω0��O��?���{�����/~>|,��uf��������4�rA����0?{���g����/�ϞgOiǟ����;~�\:���ο7�>�!��5Wg��-s�GO��O~�<��݆�xṓ����>�[���C��4-�S�|�L}�3��2��΁�*|�aɻ���l4���w6�>ja~:�������O|�R4�s�����}�4���?P��Z��=b):ߛ�Z�x���N/���.~��)��SBPBPBP�6���g�������qC��i��˗�_������o�>�&2��.9z������~?99iN�89�|�z��O�� FE��\����>9	���hU*F�t(L@o/
[o����5�lD��$JA&<�X�N�	���fY�nCt"S\�B�<xLLT�v�F��W<�)�>8���(A��KT*aD��c#GNH�444T}���Z�vQ���A�ש��OZ?��J��fI�x���URήԿq�\$�+�_my��
%���"�Zz��\.�]��B_s��;V��my�W����\,����@��;�b
�0�pk�'{0�^+��V�|-��k[�����V�Z�(�
�k�cػwoC��/����� ��Ep!$U�X��@���\7|U�f:V�wh������By�Nx6��0R�Tҭ�R-�8�7��( O�#�?���1-\{�G�{llo�Y>\϶	cK"��Q¥�Rr����(�x�"I��20��P;�N�p�GGG��m���]I��.�4��Q�.�NB�L��'�i�ҳ����ۃ�\�ٹs�ɓ\�Am2<<�Pý���9O"l����D�-[��m�m�Fs)+΄�����^�C��Zu6RaJ���-�����
v�G�n׮]��Q���B7pR!P>�~��!�1T��<ߺuK��4.��3�l޼���K��+��c�����IB����I�A�C��U�iI�M���i���h"��>u���@(�sӥ*!�l�|W(z�Z)�M	��B4��.�Y8�l��vR���Um!MC���4RV��qU	ca*���7���Q���t"���T�����y�f\�Q�҈����V���R4��G:�S��� �a<$�"B\cw �@�zѦ�0l��N@���Ëɗ�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�������==���p��b"�
��-���54%LWWw��E�1�������ܭ������ �Չ�"�k�N��4%B���)�֢����n�c�Z
C����"� �X�Cmt�dB|Gv�n�����+��7B4`�fQ�.A���h�0�h`#c�.ύ���J��Bh�暄�����]S�A->��I,z�()
vW26�Ey��TV�00v�vC��`8��%ۍ��59JS�8 9�F�� �v����G A�Ҳ��x��W���M���2Dm>HH^`�err�����`S�Ӵ0gv����G�����e����.�.9N�!>c��m��\:Z��s�0-#~�T��h��ݒ0L�H�ӱf�^lZ�E�i�{*L��}�ea����2-M���pL�x�=���td�j���!�Q�����1��0�|i�e�[F| :X��$�L���-�A"U#���Jhe��&����/_V�Ȇ0�UeH���/�ʂ̄A~(�p�0��L����L��)� �ĖE��gAf ���F�1I����,��t1r�!>`��c�#+2�e�^&��{tRY�y�ؽLڅ����e9U+��ae��2
C�v:Lv��\D[�f�&�Yj�٥c��0&b�'�_�]3/sa$g�4�\u'N����ɰC������Cڂ��pa{z5!.A�n���l	3
�p^���)����0 �Hx����0�9v6�����L.��+o[&�q��΄�g;��]�\��:M��PF\�v2�B�A�E00�K�N\��L`�c(qI�p*��S�٩�-v�慎8�R��[�7=:]}�r�yJ&������e�܄���\��d����Y��
�d�ե��3A����������)qI^��!��M�gOqA�R2��{���$_��twwU��]�dE^����0�{c���\��:pNq���t�yJ�c�)��MBZ%a\��0蹐�v-�,ɳK�"�=�t��ICHV䝱�Ԇ��)���0�dE��/�%�6��C�Ln�d�bH�Ԏ��:���#�b�+�X�+aqA;�(r]�]FٵLZ%�)1Bn k��qE^7&2%#DAn��.{�)i{�q����	�{��K\ߚ,�&%[�f��'h�oܸ����b�5�<�܄�����-;yϟ�����!~�s/e���5R��l�y楋��'gf�ks&������~�%(�0ga�\t�!~23/�ESx�#��a|�)ǵ)�03/3�cfΕ�ڴe���dg���҅�(e$lÔ�\G��Lg���K�㢔�3%�4�I�΢�m~o����+���/�0�F���䪔Fπ0�0�Ba<�dg苷�aJ�3���4�W(�g��~�R����VsIׂ����j�䕯}�y��_/|�%�kg~���ُ~l~����k��H�_�5�VvsQ~�mo1^wM��������k�1�����%�b�Ht��w�SG`�z�k��~`|f��/�yn�
jǙs��>���_}����_�|���x�y���9��%*"]���_c����ɿ���3��aLn�����]9�0�(�gg���ް���k�����}��_3?�淪���~�\yCE��_�]r��ξ/a�Qbo|�b��vg�"$pYS^u�s9d�������n����0�gN=g��w���o=a�>��\Ȃ����w�O��o�hôc��df���|�ܹ�\}ƅ�\l�y�M��@���1/<��y�D9���~ȼ��~8�~���g~�;��8m|�E�i�6*%&h_8z�6��ϸ��Ef�ŗ��3���9��3�-~w�_7׾��{t�u�'�e�~�y�{+�� �+���\��M��W���<h=3�=��c������d�Qi�8J��6L�]}�k��,����	�����o���n���G�f�UW��=�������P m���w���,1�^��_}��˩S�3��H�y����Ϧd�>�+���������M����di����p��N���%�a;��?7?���B1^�`����7�?� H	�[��L|����;K�Z�<7a��\�RFGQ���K��3^1A��_8y���8��g̥�_^y� E�}��T�X�z�㗿lΜ��A4{��;|~��_����0��.nJ�#7a�F��U
ݶa�
���X�`N�炚������� C�^=nt$��t�6z��Ϙg����WU�4H�~��S&k��y�qհ#��s�aw[#�l�3Ά)��{�}�y:H�N������0��fƸ���W�:�,r��#�L�a�����>�l��F�����[�ϳ��sI[�0..�6�9ㄚ6����IP���/��˛����޳����ӗ��3�����8��=۱�}[R2{򬨤dn�S&�1�/���ʠ-3?(��~�/\uUx�?�=m����Nzߙ��h� �q-Q�R2GƮ�]}����=�~���L��W�m�dy�ŗ��y<�ۗf#�\�8�x�g����8��![��%��1mI�\�S.#����N�q��41i�{[%U}��%(��U��/�gi��ib�)��N�0��^+�:oy�e��%;�np�}��l�Sϝ2���?�׿�M�� ���7����#��;���
�/8����g�_���;����ߌ���J��'`�"��AKPi����3ƚ|��3��G�+���\|�Ŧ�oR���c�ߜN����K�M���\}����;}�����G��x�:nD��c��'��sN�G�q�5yO��E���jk5��d�u��l�3nR�W͎�?�7��W���������_0��bsE �o|�*�ԓO����*�.�9��,WC�@�p=�O��sҚ=�c?c�^ZoZ+��6v���qM��Epچ1V���ߠK�5W�6
ҩ�}�S�]+V����_4�}��G8��?|:�,��B	3�q�������<�5n�]��4f����w�g�9�0�q�f�F@����φQ��o�3�"M��{��ߘ�Og�c�7ckQ�a��E��a�B���A����z����(O"<=+ë�F=�/�6�O�lC���i��{���C�p����z��(m�0ُ�sa�֔�g��/���8�6�H���0E�eOY�0n��Q����"��Rt$�0��1�����0�0g)���8��P�d�%*���g��\{��10S����Z\oE�\{=2Wc0���%i�)�}祽��S������9k���Mooo����bJ���e�k\Vf==��
YM����!%��>w�O����@�l�q|i��H�<11Y\a�J�a��u��WO�Sa�J�@���YW3�H���._.'a:��}�6aa|e�qef�/�sʜ
c�c�&]
������w�'�6V�������>ʝ���Ka������0��n��g���)�G�ʘ3>~�X�ز 4��R���k17�'��7g�Ԯ���ڕ08��\�q���yl�F�)�Ν��~�}���w1�KJ�G���b/���<��#��:44���;f�5�O�M!��\���$O��f�ìp"Lm:��B�#�+Y����
�a`��,ˉ���٥L�	*�9a����������t6ftt4|��`v���>g:F�A���x����i/�c��^�T���_�~!�!ڎ�R��{k�1�_H�@C_�1{����۳y�L���1��R���k+=�Y�gaƪ��~!�M)���0�,X��SbH���ٛ���̄aw2��f5M&3a������!��`���^k��,ap@vw2����e�e^c�DY�O�Y3Tӽ�*�c�_��"����[�A�V*�����c�0�/Ц�(�ʽ��D�1��߰g/�:�߲0Lǈ�HE.����e-	�t�"�P+iYK�0#E�)���e-	�k�-�1�/�Х�i�n3c2MK�� �%��������A̦��m��B�':�)�������FR����[��)a��pv2)
CCk���FB۶����M	�������L����v�/�0ب�^�@HQ��{�r�ja��h��Y���A%��-��p��H��2Z��c/�����Se44-���!�����*���`Lƾ߿Q�c/y�WX��糽��C�)��|d�n�n��,ܔ0)�tB���6 n��4��]�	)#���ja0���IY�v5%L����s*!��!D�!D�!D�!D�!DA�������ׯ<��!�0����������������������������������������������������������������������������4�ѣG�������4'N���Yoo����1}}}M��%'N��1��(P�A�3{��5������5k��7����l�����ٺu�!��0u�(t���Kb3=}4�[< 
f�{��ڵ����Ea�¤���q㦦D��ъ7����}�v�i�޽c�������uhhȐt(L�ׯ7;w�r��(�������8M����6���_)L}(L.eP�#ڸ�����0:2�YA��0��5R�ИG[��.��1C�����"��ԑ��3tP$wR��m�(�2u�0(�h���H�mc�
kl�P�	iV��5�4Y������;������P�bil޼9x����!�A�ݶ�V�J��!j��n��4���:"i6��CafAAI�Qڱc{�	���C�̍7ޘ��DYԤ� ҿ8a ��P�Y��!Z-D(�{��17�pc��!z�*�\k$�������qQ���t(����$��(d�4,R�uIr���*L�؋�ޘy�e��O�J!K�%�������׫�i#�vG���`�0l�'CaLzAEM�%�7�3��nVP�m��sF&�ƥel�'CaL�0(P.ry�o�g� 7;��<	�cQ��26���xa��M�|.p5�,m�)X�kI°�O���#i�����D���j�cd@�IJ���?������T��r3؉��.�"���D��]��L�0l��O�c#c��W��I�h���/	D�w��Carm���k��h(�i�6� %E(6�k�0932rw�Ϛ�.�m:	�]�N�0l��Bar�ޔ�F
w洱���1������R����(��L�I�.�q$Țtk�sP��شiS�lh�1k���w4��I����&P�Һ}]�)�i�F��=��Ѥ�6�+P�@�u��oL�Mf͐]��^�H�*��
��z�`���ޱ��~�T�z �$	���0�@j�{�Ӑ��!m�����I�d8��q@#i
g+_ԛ
�,iSe���0�����Y�hK���R�%-K�^����0����������:.m�L�7�)LF�V���Y���ې��-$M�Nn�S�hdi٬dA�6���-ՈPiSe:��OaZ@�z��aQV���i�(��yZ_Lǚ$���ŒPE��4I��xU��$P��Y��[���� i!�!�c,����$��E��Y�U�*��F	�i���{�<��iK���۲Z�(P����w��ÒH[`�] -�0�<dK�F���ŷ��\�(P�:hz����j<m�=�ۆ�U����0)���8�z��~�3{�6����;�i�
�@��@��^tq]X��֤vgwR���Ш,.z��%��!���㐛ђ��;��OabhD=aq$m�*4s�X3�M���?�����z���	�#�w4���M�t����0�%덳��ץ���A^����6!�S�f\�z�(�)�'o܊�.A�?m/�Nh�S�Y6nܘ:O��K��\�v[�0����0�20���@�
�.��	�g:&�m�:��OaL��X�dr�I#Ȩ}�]� �tL�Z�i�a����� �L��2�lUn�#3�"R���1���eo�w�0���oim��}��Q!lZ�D��/LZM�.�$����I�~2�̍��F���z�z�>�7U�̍���7ꥈ�L�l�Şv�em�w�0��hi��C:&��'����ha�X%2O|:V��A�'N&����$�)H+��IP�`��N���!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!DA.���K_2/��!E'Sa.��&��c������0�d*����b��k?{�!��[o5��L�yE ��?��/�Ħ�~�J���V����=��[^��[��/�>�������L��`�s�u�;bif�z������"�y��l0��_gO����s����g�
�HFHQ�\����g?�ۉ�3��Sa��`����n2��zs�M��|^�]}��qccc5�-_�,6e�?�����{roo����ٕ{���_�^2��)���w񾲕]�} 6{�~*��]�{�;!c�!�7�ծm�I:N��!A��?��[�@B�3�Y����?�ש�·q��}Q@w��^-��ׯ?o��N��7o��^�́V��5qoG����O׼�֭[����5�罹����eݺ���I���Z�
����/�Ǯ?�~cZg�0Ҹ?�Gw'�g͂ha0D�J^��W�Zȩ��v�-� �]�!]WWw�s�6n��f�����wx߸����'�0�9�\B�f�4Y^�����s�"�G�BNjv�8Y���F�Gt���5��}aAJ��Ie�ɓ'OT?�ZTD��۷i�t���Q	!Q�褽8�0�����q��>�-l���]��0"��{,ڠ�K����0�.��m��s�����D�h4���e˖��qR��m.���_�r�n�X��n�jZ���_�}\�	Q+��� ����K�ӏ=�j�6/}�	s�j�\�@��6��3���P���u�N�v�	��u�ְ# e%�lՍ��?�6[�4�if�
��S(�Rp���eO���55m�E����-��T�+{ll�i�-�?�*xm08�����蓦N�L_*��rz?�((�x\wݢ��#E�4�÷�_�.d�m�q�_FG���F���̍	��dL'k��O��� fGoR��A���C��'I�0�챒F>c;҆�`�WSB����Ԟ=��;���ς�
I��{aP��9��y����R� Ht�u�7Ҁ߼�2��!C�=�HWo�z"e���{qĽ?��Dà��o�{���0��6{]��C����ٵkg����V@Ã�K)�I�tH[��G@�ÂJ��� ���-�fH��B�>h�t��5�uJ/�4h�'���(!!YAaQ@aQ�S�9�F�ʳ�0}�sҩ0%#D�!D�!D�!D�Z��Ţ�����k2�C-�4�)�,�b��Z�d�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�aN�8a&''����ݦ�����t�@��������W������1˗/)��G���sz��H%dW@��]������˗�?+�f׮]f�޽�cL�w��x��A���A�að���1�����hU�$*��x�{�@�5k����`)�g�����?�eg��,��?v�;~<�w�>($x �l�|W���@�322��9��۸qS�(��,�0i����ҥ�1�/6�-
�.�}���92e�LM�Ç����9j�+���c�vS��SOT8K�,	����!�*�c�*���c��቉����糨�N���֭�I.��2s�m�;���������W)��շ�������}�@���g]wݢ�"o/tو;��-+�T>K�
(����������5�8�����,R;�P� 7^�~}���nݺ�fepQ@��H�v���{���j�A틋�g�C�,�YD�KvǈT@�EDh���O�;��B��������t�F\XԂ6��D��c�a�֬0�{߿d[(̽��Wm�@�o��P9	T>;w�y��P+�ā���;���J3z��Ո��oŊ��֭[��А�B���qP[�WjFH��n�͂�x���a��Q.����V��sz߽�dr���g����_��	 �Ie�4���m_ذ���3�e���
O:j.m�2Y]|&|����"U��,8���n�ϼX���f�{�cn�v���@����Z�^X�qQF^G�3��B�?[�U�V�C��M��jx��\e�z�{�}��tuu����#�
#��B\-Q F4�$��Qi���Zuki|PT��Ϗ��k׮��!uo����[aP�H�$�KΎ�D���E���J��������r����-���zo�~��L�4�?~���� ��DI��hR�p���a7r(G�����Tj_ϊJ���jG ��1���M��X* �����Jp�}����h(|"DZ�]|pw���p�^���荓T����R1{P2�j'2������}���Ɩ%�l :�[�6��p���Oz=+��LjEJ<|��b�bHU]w�*HdR	�<l߾���W� �؍R����e�"^w!���2# i������b�b���v!�xǝ�Gy��$_��W�l�6Z}����O�&h�q�9b���,	?��\����\`�c	��1���^[	�e��������&v�Y9;]W�D���T�v��w2�8�1;��ܲre�|��ز�c]���b��n�&ȁ�G^�:��
}�!�ΩLJ-B���m����1/f x#�݋�����q�D
	���NQ��[��or�#:OP�d�(�A�����$U��ؤ�w�R[��,q��Ť�(�\`�	�O;���2X��H��<x0��Q
#��9$J�ٮ`f�#�i�/��Wt��(�����i�.���0�A�]�D�ζ� Fԫ_1�Mu� P�5�Y /�GF�}��^c�"'���� Pca����T
&��~�V�s*�BD��()&�d�셊H��vo�o(���]چ8��T�_�,j��(�&w���GeL�h"�W,lh�6~�(,=i�T>Z(�������2 ��apN�=��a��iM��e�ymד2}�}aQ�q�"E��7�jA��X��j�F���#7~ͭ��$�q����/�^イ6�˩�@z�@;sn�pU�S.�,�(.}��H����3��k;�mw��&�gl��EŅjά���+��Fv���Lk[�F�*��w�J�{O�^:ہPJ+H�2�'e�L��l�����*�XM=�$}��,R���R�e�&kf���Voo��$�P��(�}}��}����Y�����������dQ�h��4̈�N�iY��2�yE�)�}]Lc���2��$�����RB��)`��v�0v��>AY��(..R��2�'���pO�^"�5ӆ�6��z�@�E���RBy?,;+����v�0�"A��Ǜi�ed9)�>�v�DVsN��2it�	�H��^ ;%L{?�3�]�pҲ^)i�%��vtl��4�h�ɗSG�8�[ t]����R����Ik�ǽ���m>��^�';�Y�IQ&n��Y�P���+63���]bw7��@2ݦQ����rn��R�A��Z��(�դL�R2;��=���r�:0;�3N���}Г���'D���|���b\��j��ko�v��;�TҲ}��´�~��@���d�X�xqux�r?�I�F�kR敹TL�U�Q��fw�,��&O�Aa�m�耧-������7� �?"K�ZO,n���I��e��5��'�i�ǃ):8>��hg�-�a){z���J4,S����E�I�oeR�=����b@䕕c\.�%�4vti�xQ�'G�2(ԭ�G�(�Y�����b-��n�"�����`�%A�����(��+2��^8)��r�hdCM���v�i�9ǃ�JQ&�{W�������u@�ٲek��
�l*�}�e4�2!3�5��c��tU�h%�9t��7d�R@z�ܳ����D�]��j\�hQ��T��}����Y��d��`eF_�.Q����j_�� "�T@8������Ka N����nf�L�fY���%K����hw-�|�yT@8Ni���1P�K' �o* o����N��GRz�P�g)M�\��I�QYP}X�p��M!����~��Ѻ�ݲ�p˾&�`&�[��Y�n��X�}u69N�8���`dD�Ǵ!9��4G�iK�K*A;�`�w��;�y-�Jp�1��f���A�ҝA�`w�qu{�nI��&\�mj*׍�Q�6�,�W@��AZ��iZ]8.�Ȫ'H�EnÅݲeK�d����rL���2E� �m��y���B ��ԑp�b�Ռ��Z�rK�ڦ{�D�w�Y)�g�` ���)C��4�6m�nb%i'mo�|&�
i[P�Qǁ��/Ӊ�Qa�\dL�Ao�DԎ���[Xx[;0g�X���0�2���ر���v�H����`��w��D�me�1��`\�-
(�9-�0jx�p�^�[���#����/�⊚��lp1���h����Vq
>ϧ�LYS <Rm��E�}���M��Ѐ?.�tb"��s�U�H]Ha �|�v�i����Ǭ�_-����0U(j[E�D���Y�s��;7!"G#k1�(hw��VA�A#�Ta��!�En�B���8�k���-����ϕ�����L�d*�4+[�0G�N�,v]�#�&x��D�V�8�h0� [��\�{�D�u�sY�i�̔)B�F�(�M/2�Ǯ�{#�N9ץ���cy�UJ��������������α�������[L(ĭЄD)�0Qp�?ne�m�pR\J-��X�n=�ɌR�j��N��dKi�A*&9`	!�����Y��V���ު4HͰ�YQ'�RZa z�$�H � �PZa�ZLt�:t <��!CH��VYZ	��ɲ�X��˼�%qKi�d�kD�����i�����2�bF�ٸqc��!Z:B�)2+VTVlĸ�Y΅����rD�f:ı��c�X��i:�-��l�D򣣄9�`��3����  ���'<� ��pÍ�s���@�#���^b`lf�~
C�ӑ� 4����V7J�$��c�A�e˖�fժU���2�ԣc��݃�W#$���	�����' ���zt�0����@H/@��];kv[&$�R	��bY!F;���@����t���]}��q��G��!�5��������������jap+/o�%�
#!
(!
(!
(!
(!
���9�����!�
#!
(!
(!
(!
�?2�p7�O��    IEND�B`�PK
     #{dZ-s;�.@  .@  /   images/3e0a96b2-ef1c-4fb2-8b57-d71cbe1f3744.png�PNG

   IHDR   d  �   {㓊   	pHYs  �  ��+   tEXtSoftware Adobe ImageReadyq�e<  ?�IDATx��]|T�����%Xpww�P��k�-VhKi�����-E��+$� �5	��~s�p$'�rw����~	ɻ�}�������8�����8:J^Ԁ��(�g�A\�ŕM\1$��8&�{�F�gq�$��$��� �u�ƨ�����'4BU8&�iBBb��ŅZ�jEY�f��)�l	��>|��\����D3�J��&LO%K�$	��o�~��D?7(�0K���I�~��5,y���Bc� $!*�$De�����A�2؝��w�ҙ3g�L�Ҕ/_��~F��B�<�`��$���رC,��R�:ui׮���!00�Z�jM�ƍ�#F�D2׀F�Hǎ�y��ӠA���h(uj7rr��S��Dttyxd�-Z����e�R<�@�����ݻm۶�F�M���I�0�N��P�4v��ׯ���P�֭I"1�MxGD`��f=��w�Q�X��s�|�H6B�=vpp�3�S�z��_fҀ�I�m$�yS�n]��>}:ϒ̙3�Y���7G�E[��C3g�fojI�R��ܹs?����K�#2���QQQ�h@��[��W�rw��NH�ҥiȐ!�+�?}�4�=;U�X�$��;!ժU��J�*E�'�7��[e�����A�2$!AAAt��-�q�:=~����r�|��S���(}�����������u��={�?C�r���k'Dt�v%d����h�":r�(ݾ}K����+����p�"Ըqcvϗ+W�R�/_��+WҶm�����P^��}<�Ҧ��v6�.]�P���������K�}7R��Vʘ1#ըQ����M9rx�������/�ӝ;w� �?�����eǏGy�����駟~�A��Ǿ��}x-C�t��)�+�ءC{��`!M�4�~��W�޽;���<sl��x�b<x��LM�4�lٲ�v-�u+vU�X�>jӚnݺM�6o�e˖��ݻ鯿���ў8t���ً�h���}���@�������=��瘹9s�	����;w.mݺ����O���6m�M	��p�СT�l91CFq�I��Q�b
����t�K/���3}�Q[&�]�vd�_��:w�L��Yi��S�*�y�`�����6��_��ݺ�Lz���ԩ�[�u�֡�&N�-ZВ%��cǎ6k�����f2jT��b'���P�����$��m�<y*��f͚�W_⫫�A�DgU![��Ǉ�v��bq����5<��v����Ey��Ϟ;����͍�T����7��7ԣGOV�5kִI�lB�8��V�Ǐz"��Y��ɉ�h��ԪeKjժ%?~�BBCQ�Կ� :x��ͬ��O�
�eȐ��M�,:2W"2 ���W�R���Y^��G��c�39r�)S&Q���g���8�3g���6!dܸ����+���o�������2uծ]�ڶ�����;�:d0=|����bp��Ѷh&�R����/?�,�����o�!�o� O��q�7��:�k1:����K#�h<do�M����m����=Mk֬�N�GŽ����[4����j�P�<u�څE	�����K<�p��T�Vm�3g��)��0���ݣ߅���]�f�dDFFҍ�שv�b`<DD
1g��}�)իWcd޼yb��K�i)�&dݺ�<�?���[#�p����S���^z��.��q�G�^V�'B�9p m߾�MMk�a���������o �ѣ�!Hə#�EG(��iӦI4�a1�Y�v�H{���0�X�N��E�����F��Ȝ<e�0%�%�(-Q��P��h�xQk	A;===��x�1`�B��+t���?+Z���xVQ��bE��[�rC�YS�d�6%�@F،?{??��эɘo� ��A��^�'���ׯ)M�4Ij'b�ѱ�*Ud��9w��5*R�0�����~�ڵ5:��N��x��l��M�%KJ*�"�ɓ@�(�lM�֑1m�1�ܙ�'N
2���G�B�8z>888Ʉ�8�s�v^��a���`uqq�6�~��ܽ{�X�<H9B�={*�leʔ�h�dl<��~A��>M?�g�Xɛ"p#�Ӛ��}$BȜ%3�c@[=zD�K�;w����Ư?�msww�؁/^�5����c�/�����5~�k��3e�Q�
�M��x�MB��<�#  ���,����Z�"S�<!:}�!ka!X`���b�z��d�ΝG�wS�xf��݋jժ����b��CёT@o���%戽*�X�hz���D�9c��XXf8Z�u�5���`�\�Jߔ�}?g�\z)�ߍ����3f�WJ:�<�7�d�LI"^���/f�)@�ݺu��6i",� �(���J^H
�2`Z��K��;}�+wLy�<�#fF��KB���ʕ�C #b�S�No����T��Bw��xV�N� �"��m��G���֣���sXW�߅(���öm�Ұa_�YY^�G o��B4r���D ����1�ϨM�.��6m��gϲ#0����Q�]�Qۏ̊+|�.�'ξX�	�Y�ɓ'ӊ��lٲ��Jnܸqcً�20�^�x��*S�,թS��f�����jժ<���b^��L~!fw�B7����byx�`稵���-XOp �3�9f�h�ǧN�n1 ����K��7h���lvZ��A	(��V��0�6��C蹦͚�>H�l�L��]]]韭[Y�M�8�j`o�A��8�$�C�֮fk&�d�����K���獟O>��l��7�ԩ�ٓ'&�}u��Lٳ��]�ٺ2��0��+�g$[�&����v&�8O�<���©k�.T�F^,)^3d�=F��r4k�,�%@���Au�֣aÿ�ӧ�k����X�A�\�F�z�4�?@���aÿa}�g�M��&m�َ!�x~A
Bh�4m̾ 4�ޘ,��b|��%-�k)�W��dt��Q�X1Z�r��}�����i���5f� *U�$o���Ĳ��Oډ�ALaf��6lX�֕�`�=ulm�ݻ�w�0�7o�"�VG��eX#�A�Gu
;�ǎ#o�t�Z �oߞfϞ͇D��C;���K��=���C:v��.\�@y��a��ډ�=8t�f�-� lu���ݻx���Ů��e*(�z,$�I��3ׄ��Ɉ}�ҥ�RVЧ�v�� �I����a=�fͦ'O��f�c���]B�`V?~��^�Ц�7�ŝ�8t��Ĕ>����<t��޽�ܹSL��X8�?���}�5klhٲ%կ_�]$�	�=��)�D�M����{t��eڱc'��	��7�B�qn{�^�F.b��U6.L��u:/���h��q!�X}�P�\6	`P�d�X&��7' �p�R~xJ�I�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2$��֜�0C��D�����h:q��S*I(#a	4�>af��9�А��,a_*ӑ�'(��䚚j�Gy�􎱔�Ցһ8PZ�W�=�z��| y��ء�	���
�����X
���h�>D�=�g���݉HIL����#�.K�K��,α���I\��Q|�$��n�h��]�_�.���o���M��aA�:<�^��Ux4��K|Itb�J��0jeEGEPTd8E�GG:ES�PB����E�Nv D�~"	�"B)fID��CqE��#�1v�O��*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2HBTI�������g�}�u9a��ط���/6��ߨ�!�N��������5P V�nTd��Q��S���Q��g'��t�H������rvr$�
�#1_���1���X���b� �F�8* �yt4QDX8����Ӡ z��=z���<���'�48X|}L���'�S4�+z����L�lL Hrtr"w�l���FY�d�L���5[v�r��K3f"WWJ��J��vhI2�y��HBD�9h4\3��IC����WH��ҍk�����tC����`
W��h�����f�qpp$W�T�*eɚ�����*X�.��W�(M�4�N=�I��̢d�Iv#D�#�فЧ/�?�;�oҹ�'��9q����01�o�u�&��m"FXX(����Ā��;�TLH*Y����Q�
�(O����Ip)�e,d/1gӷ�Ғ�����t��m:s�8?z���{�n�w]��U���x���;�tz����<f1y���,u��<��W�JUkԦ
��R���)uj�7�ǆ����Q,䵳E�^���%:rp/=��Ο��Œ�΀�0�!)6&���YB�/��k���Y裲�+R����zͺT�H1J��-��(�gN�Aw2	B��Eҵ+~�s�f:�{;�?w�+�h���)ou`of��6:��`��{�rK��ʔ�H���FM[R�B����L��LNR���ظ:��
�đ?�G�����	�C����pHV��`��y���
q|��_���"�iˏ�^���3WN%�a�����x���dX&���t��c�o�:ڽ}3ݹ�_\C�_L��I�����K�'[��ФEjҺ�*�]Hd��˼�h��XJ�$��K:tt��Mg�VJ��C$����@]4g&-�c>U�V���J%�6 �ԙ�!*\kK��utv���t`�:�cݺ���%���,b}��`�RT�u*U�9gέ]�@��h�������t'�?"���W.Ѝi�R��S�V�)��S��1\X2<�����K"l]?=�M�L ''geuupPo|J�Zk�X[��S]�[��x���Q��R�r��iӊUqjJ�.�X�8�W]�zxx�{\�r1���w�~��ի�A/_��ׯq�����ה#HVBu~�t�c�f�B�s����gAʓ'eɒ%�����3!nnn�M8)Aȋ/9�(D,Z�>}Jw�ޥ7nP@�5�DO�<�gϞ%x��#�\�+!�������E���%KR���(�����.�j����+_�Yƀ�Ȥܾ}�Μ9C�Ν��ׯ���'~�w��h�g[���he����#�+F�+W�:uꐗW1ʙ3'�x%�%T��q__��Q�R,�L���������,��Tb��
\ho�ƍ���;�I ���Ct��a���癤��}sV�/���]�\�rT�fjР�*U����g�����Ǐ����G���{����w��}�� ���#����9�
DFF��U��VD�&M&G��E|MKٳg�#�ʕ[��\�-[vq�����l�K�OOO�@ܭ[��t��A��������$[�$�?�@ܴiS*]�T|G� 1 9��v�j����(���<�3�7ns%�$ 3��Rb��M���Vƌ�@�LD�bE�P�B���k�Y��jժ�___ڱc�޽�N�>MϟkuPRg�r�b,^R��_�j�ZԦMjݺ7\X8����ʕ�,�/^�?y@��3��a�����$#�\���>��*��2eJ�[\|_�ʖ-�׈#x�m޼����o:v�X�̱��=�/� _۶mK�:u�W�\!ooo:y�$�:�/ݼy��P��F�}����$��:w�,-[��j���RŊ�J��L̗_~�����
Z�n]�|�8�B�H3^�;�B��mݺ5�P�j��>>�h�ܹt���T�4}�b����!� �ѣ�|;�C�g�x��FK�:��^�zԫWO2d0?~�V�\ɳG�W�-�D�h� ʛ7�k׎��oN�8I'��: 88H���!�W�k���ߏ�ϟO�2e&~AP]j߾=u�֍�m���@�	���n_8o޼T�Z5^�ݹsWL����ߘ���n�
	;f.�+��*U�r>��9r�%���'z��ŕ;�СC�z�j��wA���A�]�~�/��#��\\\ؓ�#%��a�C\�R�����P�=|��C?�!�ِ�ε���D�B�2HBTI�� 	Q$!*�$De������(!��s��}uBZ�7�V�p�dʔ�␛���ۨ�)��<T�D� 6 a�$��ڵk������# ���c����S���7n,�o߁�Z
��?�K�|�	{y�:u�oF�HR�(��ٳ{��G�$~��w�8���8�6m����pJ���7t��I"m�/�6��D�`Zb�_�Я_?钷!����۷ؠB\�Y��Q��?�!b��ٳT�B���,YBE�᨝u��&[E�s��"�-I�m�Р}��Ӱa_	�e88� !��ݠA}Z�z�92Q<���@�#��:t�@���7x��ub`ԣG��jժEI�tŊT�JU*]����Q�722�5j$|ڲ�I��@P���g觟~���@�=��«#�B&��hp�����LB�-L�gb	��B��A�R�'6�����hS0�Ӏ��uȾ}�$!I�X> ��\��YB
.�G�����_���8~��J�7oa�^����Z�jӟ��Q���������)^��콊͚ܰ5�3�ӹs�$!3�ĉT�R%ʐ!������pB�ଈ�r�$"�G��A����I!,f�9��FEP
�*C���(�9�^����L>��sʰw�^6u��+)&+�q���	*I�2��/�P�p���:ń.\��8q��6mB�q��-�L?�����(&�qv=%��ƍ����)]�PL�#�T9z�(��0�;DB$Ȝ9'P
��A*V�@k׮�����~��i���+U),"3S�Ν;�3�~,R�y�T
��;�.\�H6$	�x��1�i�Ʋ��E���}\�|�$L)�?~D^^��W���d�)׮]'	Ӏ� �,��1����~HH��Dd"����,�ń,X����'	1�۷��73f[�	�O&88�	���0��3f̠�宏$����)a��u����ń �$�l6��5�Iq�ZL\&PV8pb�m��7Q'4dn;^^=���bBt���<1OJ�eVFm��|�7�P��YPڽ�lY#���і�bB㋀���FdL���N��7e礚
8Z
g���7���{������#�
IIqe1!�h�����qr������!\l�ݥC�Q���E�df�����w,�6�})�@�G
qO+�ĕK}7�,^8,"B���콺B NN�d),&���-u\*X�ЈFE;����'�	� �����������(g葰�pR��:i�yw�x
s��}H%9ոr�%�@g��Q�:qE�����tkȖ�c��G�@�� y�x�G%3D˄�с+@kMe�2[X6ptu�'E���i���u��#f��J	�&Pp�r�Y�j�&?K���S��M���C���}&�,��B<߽tir/S�\�wK������Yzv�F��u�S!�DV�[�A�g1CBŢ��ԛ�.I��J��磨�n
�cnDBt::�g����t)zt�=�p��g�,@۷�;>����7"6�
�.����`��p�螋�����T��#GE��}X\=uS/ι���FDF�&����X����\�JRfAƹ����7��o�^�\�Q���������r�("4�\�:�	��{D���UN�жp�����mRY�$YY�Af~\��1Y �����H1����~����](k��t�?ݾrU��7f)2I���LE�Q�R���Ejצ��7)[���6�<}F�v����h��6\���
�ϓ�'�bB�	��+�V:�ݤ
��1Q��3D;��ߏ����F�3��s�@G�@d���P̌�ŊQ�X;���N�D������LӦ��j:�i��F��h��f	25X
�	�'�� R����aq	������?'!��ԢW¢��Mx��%/� G����� tJ��;��LW(K�\)~mr��3DW���;#uHAz*Ka1!�z��y{R	@HXl���#1��{tp��>T\�&�gZ��H�LrME��s	��(L�Tnb�M�#"���bvG�8VXu�QBDƊ�iu������
�']����-�3J��z͗�h���Xmݚ�X����+"+�3�&;@t��

�L�����o��:N�Ly�ғ�O�uxE����1ڿAڿǄĚ�h��,*�]�v��H\�`1!�i�+���t�:/kVdň{R���h/���A�"�:���sT�I��U���]"�n-Q�e̞��=��\\]㞭�hf�n�ĘY��-Ju����E�K"O,&ǳPgDi�5DV8��X�3$�S#1fpL���%E�F
��w��R��@�e����{�����=^��̗�r��q���)����E1�� :,F�����	�k����#,��A�"�` ە�7�c��4�B�C��I� �8B�߼u�^@΋1���rL����y��%���s�ݾ{���,EK��>��o����"#=��9!�������g���Ř�kKE��_�|a�b��������+�/����c��&��mڰ>.����:�i�-9����p�������>,�l�)f�A����ַ%��s��z�kL�����ܹ��W\��R$���N�$+'����XR�v��	��ELsGh��u0p�F���z�X�*pq`��|G'K�̼4�@K`!��(�ӬY3şa���]o�aӂk��(0�P\?�����)�i���Cf�!����� ���s�%�����%�+������b1�o2�w�gI�L���鯿���!BV�9{�#�1-%@8LΜ��S�NB+�CQ+P��a�R�xU�"(�:e�d.�j'B�1J���q׮���ɑbb�]F����䘷�*ų�f������8��bB��Eh�-T����'O���U�һ�`צW����F8�ܳgE�QL��q�W��J?�E��~���������s�G�Q�X�!��(!e�����VLȥK��.*F+�0�׹��>��Ϗƍo��B��)S��订��	9x��h��,D� � �������-���ș2mF:���G(��B&Z��!���=�ݻOтZ!�������ߏ$	� ��˫W�V�G���aa�,%,G��Mh	�u�Ș����������� �>,M�����>L5j԰�D���Y�[�n��ݻ���,!Ȉv��-�:u
I$	BM�ݻwQpp�Ɉ����RjT�^�$��v���_-��45i���}F	����;vr�E��%��ʕ+���"9 Ę7�(!p��9s��
��=IX�ȅ�ڹsǵYTXR��@+W��L�2S���I�zt�ؑ֯_�����?4H؃3�\�4iB�s�&	�Q�^]���^���i�ABi��7oޤY�f��m �o�-i���F�Gqe��G,�����ЩSGZ�x1���HD��ϟ?�`��{4��oÚ,ʔ)#���K�»�%KV���N��!���{R)T�j))	t�Q�=�3!�`�����E����n��E�����sĈw{�Б�0X������f)[p��]����U��YY�&M"�=��ȋ�3�~������2:C��o=b��Ya���el�`qbD�:���YS�Z�0@�ҥK���#�cDCyu���l�=��������0Zk	�!*ʰ�Qu"��ظڭggJ�P��y���{�y�|r�P�$�ea@O�P��[LHlxI��D|�_�h���3�/K�2HBTI�� 	Q$!*�$De�����A�2���B0�����ӯƀ����v��Ln��E'N������|H��踬Y�Rɒ%�]���n�:N ��o�~|�����|T����&����E0���Dg�����4g�\j޼9M�6��Ɣ����v횷~���]�vU\|>9�
BP���҅��b��م��!.,,,����X�u�?t��yڴi#�Q��+W�W������\�xQ�|�	VR��~�>{��.]����B�
����,���Z��3w���$���5�!!��Ι/_^:y�!cɒ�$!�X�j��=V��;i�D!�F�u�.���Y��?@��(f�9&)��	�����'�}���h��C��0%T-����x{{�W�5j��l���ۗO.]��Æ�i�С\��0׮]��ڬYS>|y��5�]�v���)J���gH�7�OeyT0��/_�$^�z��1�,���q���ըQ#V�u��fB <x�*�{����f팥ԩ��IYb��ٳq�+RV` ��1B֬Y�	1��ib�}���x�^� ,T-�=E	)Q��;wV��L���� ���d�f)u0:�A6��[��ϡ[�fMNr��E�?�_|��`��7.K�}���PW��3V�d׮]�:`q�x�v������[�h΄���wC�_�ݲ�:�F�+uK��S��+H�wp��X��5k�A�2eʳ����g͚�A�Z�F(�����N�ӫC�~EϞA�h�H�g��3x/�-���W�	KiW�P��>>G���W��}p�*�w�8a�8�?n�M_|�ѕ�ƍ�C��V�Z&�>�O>��	�3��8Ȣ,��N�2���+WƓQ�~;v���!���B�X�R�*�*U��͛7���ǳ��{����� �\$0_ud`q�4ƒq?~����1�+�ڵk��)w�;�mR�&�p�n�9i�2*��{Sg�̑�@�`��M�s��q�hX���)��UK��]�vc������kЪU+M�]y��	m۶-�ڳ��ƍ3z��F�ƌ�В�s�(M�kK��$L���:�:2Z�nMK�,1[&k��7��+y�ლ.4�7u��+2x#%�X$7TG�o��F_��}@����>�O��:ӨQk�h��J��qߛ�]��`��a���2i��d7:租&�7�|���/_�	  �3{��Im۶�lԦ��D�S�N�cǎ���o��g����P!:2�g�c(C��4g����ʓ0#Ջϙ�T�����?��+*���gϘ��Y�>��� �?��ȓ'/;�,ɳ��ʆ�{<�]P���5�#GN�f �^���ɩ�S�T��[lJiϴ,�)F��3�BT�?�g��8���4h@˗/�� �[r+�'d̘1�T}�b.��0J��k-#�����sҦM��Nl��c& �+V��pA�N�h�����.���}�H���+\� �V��\%�P�^=*R�(]��R�^�$�rOQB�u�J���'�ٳۢg�⏷w>�Ӊ+d Mj"��6mZs��<(wÆ%�rO1B`��:�/oM��W�^q�n�
.��Z�6Ĉ͘�s|��ՋP�t��;,��B
���[�:\��ׂ�U��A�JŌ�*�S��=�^�я?N 59'�HL	���%�6$!*�$De�����A�2HBTI�� 	Q�@�L`fO(#$. �!��+�W./�����7����$��"BR5jD�W�"��#�^��\*U$�Z�݇���}� c߾}�Iչs*Uʲ�&j�"B\��#�jU)���S��/(ݗ���G�c�l�2���-a��q,�#��	�"#���!�r�Õ�m\C�X�j����d���{O�FtJ��~���=)
�b�=���&Ы�ȹ�9�OOi[�&���xK5m�4t��mފ�z5����9�Bt���G���Ç8��ѣ���;X�!Czʚ՝�����9<<��W_}���ABu5p��\�oذ�����i���{����@�����g@��P@�T�b��V���~�V���e^�'=5��}|�e�<��{�(6,�\ �\��f Β� �̙3i޼yԽ{�Dl�6oނ�=�����ׯsڌ��~����K�ʕ�R��Ǐ�|'gΜ� 8��S� o��tT����y   !��Az9ciR.��io1���r��i���=!�s��e�7�n�B!k�Q��e�y����Bՙ8�0P�� J�a�1�8|��p޻!���A��ܹs83��e?>a�T��=G��9�G�l���ĉ���-ƚ�lD��[�vD�^�v%�x�b$u��)���(����u�gH�"E(X��c�ե����q�F�㮈���Q�5cƌ�?6��(�<PHt�m�V�%:r��o8�Q�Ç��ѣy� ѡ��ڡe��$���a�c���b�G	�U^yj����ŋ9��˗��Qc�i�3Z��abԎ��ݯ__��}��	�G�+��b *���1U��W�jժ��ݻ9,G����у 1�x>���¢jŊ�2��3�h�b����,�aS�Iv:q�x��1zq�J
������ � 芄7:�g����������Ʈ];��Brc'q�5�ݗ�fq�U�F}��a��>�6m����Q:2 C�>�Ϡ�p�/0Q�����o���C���5Ya�4�� ���<"�z��0�[�55 �k*C'�����@�;	{Bc���Q� fcE�%�,CC��`C���-[�+c�A$l�rtm�u����d�4x�����F���ޕP�#�-�2HBTI�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De����N�p|ge�jb؝��/_r^�����G�q�|d%͖͝���a�:u(cƌ�R�I/TF8y�$8E;q ��)��W���${�n���2��-X���v�O��
�����f�ʧh�hٲ�4k�,ʗ/?�@5]y�� �d#�ĪU���/ڙ+gN��8`z�ߟ���GS�N!�|,ǻA�=`B0����џ�͍�L^Ŋ�k*>Ά�c�?G"�/҆��AѥK���MM�6%{Ჿ�>�F�%f�+jР>���[�iF�9f0�6b����;i����F�;%5��1؜�s�۷�x�4��/y4�#E�J�.%�UX��8��9sf&�V͚,.f���hђ�� N��H�e˸z���Q11Xte���_{���,�VV�(��ƨ�6W�|d��y���qn[���lڴ�>��3W&�|@�nݢ&���I��`#N��^����Ƒ�q�'РA��� �[g�{��� ���C�{��c�螮���W1�1}-Y�����1c���R�r���r}�H��4u�$.ō��k}����B�"AL����M\Jw��c����èQ��A�u�ֵU3iܸ�L��!C�k�.L�%�(uIp�>�Ř���1��MAg���'�dX&!!��X̌���*�w0�8�3g5iҘG�����$�����ԻO?<xת�E�`T�A}�V�Z��܉;7)g(u�a;�gܺy��@������	!۶m��,C��Ž� �|T�ӓv��I�:v�U:rԇ�5m³��9s�AB����{	����D��pw���TWU���a����Q�c��5��=NnB�̙C�=XG藨C��_f�J͛5�Y�4����1�!k�Q��U����O�����BI���4�1r��,Gb�HB�CM9r�.]:��?��)����V�r@(]ԺUK^_�0�~���&O�ܜ	%�ׯ���jԨ_��@��V-[�T!|}�sꦤb=gr���麀uL�����8˲Y��\_̌�q�'����ϸ���Bf/\��5jȲv��T�J����ʔ-#LOW!�'���#��PaQa�q��)�
�j�^y(P�ʔ.�bR�3��A���Ãʕ+˙�@�5�>�&eﰐB�fC���h�"��=�ݻ���Fa_�t��%�N��es��%�*��:7�������А	��Y[��i�S���G��B\�|9�[��*&L�%��O��M�#&� C�O3��o#W�HL*�&/��XٚMM�4�5LH�F��6W��C~���w�
���j��t��9J�&�贼< J/N�j���ă��8}���?�ݷ��	�d�|"&�S�x9:��5w���w��(E	�´e�Y���A¡Ç��[f($��YP��x�BX-�g`%��t��΋��ժV��\�.���BY�L�E�U�re0s�n�3�2�rݺ�1SF�,X�ʔ)�3I�����{����jB��7e��v�V�J�z��U�V�aEn�<��u�MI5)u��a�a=]y�Q}��U������u��nڰAj�Q�w!� ���5kų�)��1��!���Aw�|`I�Մ`�?S/�e��,A�_(�F���h��3gN�:{'x�����d��t
�0a�#�l̊���(����ؑxM̠?�\�톨�^)S��k�N,S1m�m>ǎ��3F?�WR`5!eʔeg^ &�1`� �k���i��-TU�X&�v�>}z$�/H�+'��E'�m�BT%0h�>A0 �{����	�Hw��$�)Q����v�<�:u�;�ˢ�XMHYa���Ģ�a�&���F�?��C�N���4a�A����9v\,S	����P�Xܽ{��l�j��+k Vfp�ڵ��h�+W�O�/�,ĳ
���x�&M�Z�j5!�έ[��E���SҞF�u�Y��Ӷ�;h�Q�ѳ����>yK!r1Gam����̊)lU;۷�@��2�W�={�P\���{�g��~+��=�wv�"������տvG/]�\t�踺�Ɲ�XD���b��F�9c�v��;a^�^����_|au�U������+����OJ>}��F�sbq�D,xkȇo)lB,�����ɓ٬��J߅��K��o��HcF��\p��UnK!��T�(�J�k�n���Z`��7VtZm�5�7?~�Ɂc:_���~g���ߓ-`���t��j?�
�J��,��0fIժUh�[X�_�`�"��@
Տ=�}M�&M�Uِ@�elx�޽z�,���20;
1�}�v~&6�l�ЪU+�>iC��Q��g7;�H(�"�+�#H7��7_�R�.�����^���j�%!���֭��F��ϰє�դ�SЁ�^�M��[�w�΄�
6��`˖�Աc'A�h^o���-�ַ`�TQf+w��m۶��c�qrH/aN"�R��ST@�����ѥ����/�`��v���S�cp�w��y__���9t��i�@@�-��l�7o^ڽ{��������l�ԫW����7^.T����5�B^��c�_�~\֌���7o.�ֿ�n��݇jլAͅ�՗�=9�83�i<���k�u�6@�,aQ�����m�K:�Uz���S{�����斚Wƺ� u?�E4i҄f��3[C������ΝK���BD$���Enž���)@M��8	4/��強%������q�t8��#�u����ਃK;o),�&L�@Ç�ӧO�ѣ>\���1�K�.C�J�U�X^���d�텘�J�Z����Y��2HBTI�� 	Q$!*C��e����?��@k֬�J;�\�Б,��×/_Ƈc�.���!��%�Ē�d"9,�֬YÑ�����WB�5�d"D�n��.�o�����H�dS��9�vA |�
��HB�5���r��|(2Yނ
�
�i�h��p�>�V�XA�}7�v��A�Gaz[!Y�!�%��b[�yN�#��Rdaح[7>�>v�8�嗟����"=�2e�d�W�>�\��*�j-Rlhb���qG$�H�u��0�������{#��]��YQHB����A�t��]����&�H&BL���G�ϻ
iި��A�2HBTI��`�����I%LØ�(�OArH>V�@~�G�%,�3�pUCHDn����cǐ�}���=��'�T�,1t����D��!���p��ɇx��OΝ�F)
&$:��������h�\l    IEND�B`�PK
     #{dZ3��C� � /   images/cff7cff8-0125-49f3-ae91-9e6ccc0a4cc7.png�PNG

   IHDR  R  ~   �,  0�iCCPICC Profile  x��||eE���6�ѫt�q�"�����ٰD�ݐd�b	!��l#[`a�.  m�"M�(E�HS�. � MP����ܙ;�w�������w��L;s���;�%ɾc�,�3��$s�-�<��Ǟ{UWz%���K6Jt���-]]	~���{,i��G�i����g����a~���a����_:`���'�}�s��Dc���!z��G��xrzS����
:�jKf����d�:�Ë&ɪ]�i�=<�2���м����3�Θ�$�A"ɬ9���>�Ɯ;����I2��E�ó�dm����}F�5k���6)�L\R��~��.Ӻ���nU�2֜�ff����[��78<4�M�$%Ӵ)KӁsY���L�M�M=Mف����n�ٻG�e�'+�iIW��d��-��N�˒f�J���֎�5��׭�Y�`2���P2�l�4�]�3�M�^�����gI�Ԯ�� T'~{\ˁs1�Y�ѶE{oR,���g�����u����C�f/��@����jM$=	�Bos��;}l���-!����b�$I�`�!������d��c��$k��$��@�y�S��������������)�9�%ɵ�m�ɓɫ��6l� vmاaY���6<��ڨ5Fe���:d�e��]����G_<��1��sژ'�n6v��+��s�wĸV�x�y+�v�MV^��C�LX�;�<Va�+�:c�?�ֹ�]���~�z����rͳ�Zk��������:����i�m����w����~a�/\�aۆ�耍����M��ț�n6c�7p�c��_L�x[�_j����O8cˁ���국��f�/o�����iv��k�}�/��u�|~�8X�Q{���Nݮ�ӷ��C;���_;�岉��>:�;�<y�]���~���t����ԍ�Zw[�}i����O���5{��k�7���ߞ�w��o���)3���f>��}���y��_����^�xs�p���]v�w�:����>��#78���s���vܣ'�w⸓.8����O;��	g����g�t�%�u���Oν���]���W^~�{������|r�S�����r�W�ܺ�����o��󮻮����N|��<<���?^���lz��g|n�秼8��^���]_�ፉo���x�����^�тO��_�?����ڕ\�|���pݨG6��3p�{�ye�A��w�J3W����*7W�^���[��5�Ys�Z�}�:����z^��>�p��&l��&{l�x�S7���W_nL���MZ���լ��ns���������=���7�x�XY���כ�-l�v[5�~�vޱ{����������^8麶;w~l�K������n�!;w�2w�q]��vo�+�+O�j�.����=��/���7_�֊���޺�}��͘3�p���3����{�~WϹ}�C���O�W]�ɢ���/����Z���c>c�%߹��������#�Q����ѳ�Y|�����q?<��.��U'^{�/N����N�|�����?9��3�8�Գ~�c�>�C�=��_��?�`���h�O�^<��/�x�֗�}E�\��U�|�Օkֽv������冎w����C7/�ղ[�����κ��;����~s�o���߽|�w�{���������~�؃?t��w���G��g���������'>�������̎��n������^���F�<�o+�����������vx}�o.}��^����<��'�����>��Ã����n���c��_���a��Fm:�Q���Yc�{����ݱ҂��]����U�d��V;~���8u��ֺb�׹g���{q���0z��7�z�6�}��7;a�K�������Ҹ�Mh�r���n��6�|�'7����[�ro�x�{��-���JfU��v|u���A�زӔ�}�e��C[O���kv���Gwy���]+_���ީ�N���{^�6f���'�����W~����ӷ��{l�&�dm3�����x��C��{�~�Ϲ{�S�^_����٢�Ż/�}�A�����:��e���{�*�m~8;���ݏ����>�S�=���w��p�9�铞;��S^:��察���>��3�;���>�чgp��~x�G���@�%}���.��%���ν��+��򰫎��q??��3����+���w\�����M�����o�ආ�+w����~��o�;w�]�]�w��Y�ιo���>0�����!��c9�ѓ�x�c�?������'yj��s����������em|~�ƾ����x�ٗ��ݯ������?.{���/~�7�x�ތ��ݿ��ƿV|�����m>��x�'�$:�%�5Lj8���Q{��{�}��1?��7��m��+����U6Z����V�r��V?s���<�K׾v��ֽ�����+�_�x�&6]��M�?S�ŭw����O8g��zh뗷�x����m�X��+��˲�ٙ�"q��Uݣ5�ؿm���cvXw�	;�u�̘����I���z�?M~�}��7��t�޹tʏ����\��	���L?b���͞��⛛|K~{J߬��?}�+n����3�����7�>�o�9��m��������?|���.^��%���_?(9x�e㿣���C�]r�I�_r��G>~�kG7�ޱ�/�k9��=~0p�ܓ�|�)�N���CO;�G�~�ǜy�Y��踳O<�sO?����~r��_x�E����G.��e?���+����ّ??���9�ڳ���/.���n��������7��WO��̭�����o���?�͊;G�n�]��W�g�{W�o�}�����������w<rˣ7���]���O\���<���O�磟9�/�?{�s�����x�{/��i/���K_���;���?����o���Vo���޷�}��w��w�n|������~壷>��'� rX8��< �8!I&�+�jŊ��N��]e��X��I�J�s�I�����I2�KI"�a��g�ly0�j9.͹�g�G��1����Ã���צ�L?h�C'�Y<���Z�ޕv�8IF`��'�utT=`M�?���iI2p�{�14��V��@���u�5x� ��������������v`�dc����ߍW��U!pS�0�0{��_�+p|zT/^'����gԅx����xm��7z{�~o�~��ܿ�~��W�zF?�W�3&w�ok��9�v2�@���z�3��i/VJ������hq�>�[�P�Bp�OH%8�����/���� \�������p�e
Ҝ.p�j���|��n]	��Š�o��?If�����W[2%iǘ���|�|�En����&��[S�p,D�2�:�L8�=Ȁ�Au��z�c8���!O��e���7�} �s�;�5-�:��g��?�?�2�\�M#V���+i��A��"N��tm�Aw���$%30����@f$#:W������S�7i�D�� ����?�!� s?�4�@;��J�8�-��SX����e��|�I|�?o:��1� $�)sd���2���K���gA�qs������l��g��A�s�"��m��j�R��������;����2<k�9���9C��/�?���?<kpQu`v���м����������ۧ���:ch�������޶I�ƞ�E����Uf���N��$sՁFL=�����������8�����e��JO���m}��;�zzۺ�'��vv�M�n۳h� ��:z��;�v�u�uU�'O�n���tOn��k����=��mJo�q���E�ա�:	K�ӿ�kx~S�u���Ý���7���|]}�{v�aܝ��zv�6N����Ll�i�k�~��J�(�[OW[kowKGޭcZ'�6;���Z'u�j�5�eƤUkk�k��j��Z��e��2ejwgKG�^m��z���ٗ�i�q϶�����ImS�:�����abwKo��)}]S{z�'v�y���6�TİgGGD��=ugz�Si^Rm�v�����܊ί��D�ڊ�\48�z�Т�A"���k�fk��?oF5?��Ξ*�e5�Xm��a�����)�J�L����=���Y���H�A�;ZZw��!?:��)=nW~3��sw7d�������.�8�����3��z �jc3���s���]F0u������Ӷ۴6K�qjWo{'���	c���S�4�T�2eZ�Ķ�>ld����I=U�E<����og:��JOKgW�S
��n��d���I������������#��i��fZ����A?�c��V�2���'[�F�
+a�ҽ�U�jt�W���^U�ƅIU�����~�������8���R-2�YiҊ�����~�f��k�q����O�����2��~�	f��ʚf�[�O0�
Q1Qz��8(���8:���'%�JM��=����&2�9�Ei)h�V)�T���c�e�k<�R��<2Z�Hוl�����AGͳ*�]��(4�M%�2����*�)�s]iMs�Y4�q����u�r+5�`�Iiy5n�E�م�Y-�)�@g�٪�%�#�%�_������Ό��Ԡ<F�J�J��X�05e��T�B�)����U%�%�1rנ�*Nf$3T/�i%C8ľS�v�Y��̬#�J�F�-6bY�܎>K�MX�6�1�HJ�H�U��&�2l�p�4[��M-5�$*���NA�� �Ժ#��e�F���ƪ�fRn����I�2G.�R�H��
<P�C�G%�Lf��5!�$��j�x�י��5��56��@���0�)l�8�z�k��~��R�Sk+p
��Q�:��Ƥ�ր�{� ��)�T�[��^G0��$��e�TY�#f��p0ZV��dXOp�T�9��@H7�R)�F+s�u���I)@�����r�
$�tMH:�z��mKx��ž�K@�p�D�G�%���ʩ�%]C��T�
ǲ�Gs�Q6+SN�����~*���L���p�8w�9iwRA#�5f��	%�AX���K�uRKK�uk3if=�Fa���K��*\U��y��#2���"�'����&�q4�xMl�i���'~D�T���@+G�$ͬ'������ ���B�%�ZU8|,ܣ%ͬ'�/����;�m��>�"���N���a�dA�t����,U�YUX�ι�:�^��#��0�	`��FA�֕�0�j�:~(+L	��CU�q	Q��u�Dq,����p���?CGQ�h������?�>�����=PH�?C�_�?�*L���ʩE��;�:��*J���+58��Iޖ��	�LC�d/n6�FC��� \��_1�?�$U��N)"�(�4����@���#&��I]�)U�6�2�)p
P{سդ�������z��� ��
�C����{*qR�JM1�T�� �42�U�hB�TJ*t��b5,���h;0�\��Z�F���*p�Z�!�:�t�jx		,��a�`�FT`)��| �#$9bFhf���Q�ë�R��%ͬ'$ia9Eq˒$�TFp\W��a�_G�,Q��$�#�Ru怈�HS5�@)���76�R�Zҹ 2�,�R:J����4��pE���$"��(���p�_G���r��>��P����j�PX��zB�n�w��0#�8y���(�؎$�'�0��C
cB�"�R�iA3R�z�0	�o� $CZ�f̠�p�v�u�!p}�5�#݃[� �Z(|���	x�a�����G��j ,*J�d1����%!�B,a9�8�]E钬!Be��'&���2� h�LI�gD`E��Q����.8 9�([����
�Ԡ�O"e*O%� ��d:EG��e:PFX�i�s�a
���X!�F$�.}0�P�9e,��c}G�U!(kd�FƁ�C&������ܭ�#�i��)�%�j���QĎ��8 ��A�=9X�/ WS���wD<Eg9X�?	��=�ȭ�;

� ,���{���P �K��x�@*�@� Dq��<+֋l�>Y�R�g�C���	r�W �b���A`��SN���D૘+��()���@�vd)*�������� ��)���BN<YuT�Рd�Ry��Dq�jd8��)2��(J9��*3*�0#I�p�BW�,�(���)�T�j2�3G�tQ ��W��(�G,U��bV!����?C �A"�/�-wE�k�b��d�qF p�d�>0� 5����%�*V(��F�RR�wK�;�O��g� "wnX4�T��R��1+���[0��+#sQ��+p���W�@(�"ׁsd��Y�G&+��x�(@ #C^N³!X��
�W��3"��yXE�3tP��U��)����������TE���U%�R)�g�	�����
�е��=�T ,�ܣL��(��q��5 aԹGC�F���pl�{,:
�r�F�s:P�I�-�J������Pmi8a8��Sa���f%=�bIU��gR���TH�>����mZ�6��"���'��DO^�[���"�g�[����� ��(q�Q�3
v�%��(��:��eU�b`���� 	E>��C��YVG.z"�d 䒪3���u�3����w�(���Ѯ~(]-����YVK.zr��T�#+�����jmy�񫥴�CH)ὔs͚`z%+-'�@��`(�%���%�	;��e��ؓ���M�@�=m��=Y�(4�� �1�p�䝡�����KL$J�����մ(u^2@��)�T���2r`K���fN�3.d;��\�I:~$=��@�{�~��*�5z��t�S�V��9�jڧ.q�q���s��"�	U6��eSY���}�eS��)�f�)0�iKzFϔR�I �`��J�+S���@ rZ6�D�ŠU~8��L#��� -���/!o�ی��-[Pi�ϴq��2�Ig��D\���j�yY��y ���%=#A���i��Ǩ"CePڧ,�q�������T3��%
�SOU�5�& ����kAu*�Жt���U���dÆd��	dwH�H��Z=�Z�QIy*�Q0�&+���%^3���q�yBR��w*qpNz�KӘ��`S���K2��Pt��A�����OQ�_S�q�z�(iNV�M�$&H	��1
WlDO	� ��L�Qqr�Ty
��H���cJ��D�7��(�J�¸K�0�0�
=Ed�?'���4��\������`t�L%(9�qZ˭��P�3���� �!����U�'�g��g��=�}�f�P���L�H�EO[�f�����J�r���0�(sy�@���Y�t<�aj�9EV�

M��)���r=YfiNF�G�A�c��KI���I����U�HV��q�Tw�u�J'WyOn4��(K�cOzPĀ%H��H�)a��\�,���B֨W��j��J
o���Y���+�g�łzl��i�S�`���p�����e��}Ҝ��g�'��	�h
���.
�V�;r�p�6��fȊ���,3��	�
���~��C����2+�QT��/zR%�S>'Ҹ~H�����V ��* ����J	�J^�o�O���(��;�×t�R��ۢ'E�T@[2*S�(�I�"�0���#f�̸���P>MZ=DOU�3n�����:=Z�甔��2?�Isfy��V���<�8z�{R�R����K�?�ׄ��ZP}Or 1:F��q�TR��cq����A*0��W�e`��SGeR5��%�z䚹�^=�.iĞP�Y�F��SN�9�O�}~ڛ }̃7K]D�H}��J���(!��P�	 ń�"]D"l�dIt��Đg�(Rq�Q\d�V�ʒ�BfX[
���1����)\�t�����vȅQ.H�o�,�Ӕ��� ���'J�����)[�
MȨX.�#(�ڼgF�L�9�x��=�|�t=��BBz�������&�bR���a��F��q��PyM
�i��!�	I��F����pʤ���<O=	�iQr�q�����N(���)�)���Y&�
27�dqѮB7?���%C���
۳����ڭ�O�[��Mb�rÕMVm�n�y��Ӽ��c�y�u�yfF�~�mD�Ȫ��]:���EP� ���!������&z�Dw�4E�j�������.�=�o���Cs��1���s�.l�6��3�r�VYrIR�\�����$��uH����!��-�G:^�g\DR���ݓWJ:^M7��+i�Ƚ礥��@�x���8�Z�*����ע��b6�K��缔���$2c�tňx��G{�UѩOZ�	��2�-����Ll�HCT�=�����jEh1:��N�|T��2�EhE`t��������9�@��9^ZB��rFO�s[�/�uG��J@�@��Μ��;��?1��N=���%u��RbǫSzt�Zm�]x+��At����n��A� �����,�W�7;���D�I��'qX��E��}+��n
�:W#�V�zU~��x��|H�HԎ�~rAѵM/�@��٬���Đo�n�1�I�9?��x^�$�Z�6�df�r��B�疛�k�I�
z��0������9�L�d<�D��Gb�\�	"o58='��|7�e���,#_$] �����ߦ�3"�d�9��7$��V�$�~�5Г%��*52�Y�u�6�p����,_B� ���U�nЄn��x�Q䭈�~��":Jߍ*z9�SIתa�<�$��|~!��f�i�Pf<)����s��]�kuY�$N%t�����Bb�0y�I-�9�)�r^�?^�V���Ҧ*��X.3�^��`��ZA�����r�_�s��z�Z��yu~������a�s]�ru��_A�xA7a�v�㕩7H�D~�#'�)4]��ym�g��iH�Ck��Y�n2o��o��S(RɜW��H|84�TOB�r��(Z�V#�
$g~�ty]z^�_�r��MV� 	�)��&�F�DM�9'�nN�y�5�\!�N�<
��<	��K* 3HV&��|Λ�f�ji	��6���r�Z%z�@ʠ%�J���7����I
���`o�\+�_�� �K����V1(�w��/�$�c��"ZAx�J2+F��+ϋ�٠.ጵ��S9�k=/9k�j�)�u� (�t�d^��N&2?B�+���
}��a��;F:Mu���v�c�tN�:��PQ&���E� �˱��@������q/�\x���>P+saϓ�z�D��܏�è�U3��PH��IN�]�[\�g��=L��K�)q��0�g�,�"��|	�X�j��_I����\�X�\+�i�z�5{O 2�^�"��­	�2V��~��� �e�_:�˯��7�y�,d�ݵ��D��e�C���r�*@�6tC����C9�*0DAfE�������'����ޠ�{2]|��I�HH��
�L���{��/�� p Y�ܤ�j�N!�d�y��t��n2��0L���u [ɘ�![|΂yO����������0Z"���D��x��0�W��đ����0p�և[�ڛ4'o�<bfl���OhE��yC�@��Z�'��1�GC�8
��{.FW��-0�7�HN�7��Uy_�#��Ⱦ�C:������EuӬ yȬ8��a8D�'��&�V�}��d�0}7�9��1�#	���p~ǰ�=o�a�՟0���1CF��/���{�2{�~܈ahZ�Ρ�2�Z��1��7&�T|���6�WO��er�Y<���_ʲ0��>BrJB��"��xx���ӄ���[`(��a
S!i���+)��H�׳�a���%G���$6ă�D�)Y�D��8A�q#��p�ޭ�L�ԑ���[`��F�{؁��WD�i$�QyI�g�y��g>nR&�]7�����Na96+��n=o�0X:��v�]<� 恷�0Xm�r��y3�yC��T�%|�IY�1t�� �t�6�,b��=�a��>��F�\[�#$��I��ﱧ�BR�UP���h���-0��2��T��c1��[r�S�1kU1�i��R��I���1}އ$��U�5���ɽS �¹�"�z#����,���eIoC"b����Z:pR���E#$���J��] x�*"��y=�T������[`,'�E�	gA7e3�[`,�ER#汧�F�'D �O�;�֟E�0��4��U����ED�� w�n\i)�-0]m�NL�B��)��F��X��_*��AF#�_xCY�&z��-0�>�f�e����GɈa����̼��TH��AF��2���T�j_ޗȈa$2'�}���|��g2b$����&�t����0HWT*�$���1��a\��x�g�"#������0U���x��H�UэPYNbX��2b�n�R�Rg���0�"������K
�y�)�O�%9J����YDC�\�NC7�9D#	q�@j���F��
�xT��XЇ�a��yX$\E8!����1"w�- m�:�ce1��Oɛ@Zx�9��FRu1LL���I�fàՆq�����~܈a�¸D���G����d�0hաbZ�:ݤ�k��R�nP�2�𵷋�a0��A Ï(�㐊FR���`��i�3�[`��S���5ؼJ�x����JB��`��U�0��/sOʀ�1�J��-0ZC�H���С�i=o�a��m`���%�>��������-�'��W�u(�[`�����w�i�k
*bŘ�ABk��MK_�P�(�Wo�
*�}*=��511}ZW�����*b�L�+�����n��T�0���+}���	0��uZ1�E�U�;���>`�y�(�{�!z݁��>�Q�(�[�ިXx����1���?�ʐK��k�y�`AA� |�Qt���Y�0��3�a�*t=bEwȳ� |ȧ:��Q�F�9}(�=F�1�k}~���xo�ȭx�F�3�!X��Ǫ�a�e!��A�@�P�V� �����҆ڕ��ޗ�A�p��V|mEG�+}D媠}p+��a���ح�礦˙��FY�@א��R��ۦ���D�=�?71��k�{���)�C�atV$m��R+��:b
�,�&�&���ǩ:bڭwx��T���WG�黩�s�9i����a�d�^B^�C�<>��h�SAPT��"���k�x���`��l��?�À�{��X�Ky݉F#��O�#���5D�"|2K�T 9=�p��`
�Y<��O�Hn�`
��%@g��@執�a0��nE+���Iz^��FCS���B�J��a�
5��M~M��sވa0E𓚤Zu�Y:bLa}�Hw��,��5DC_�ࡄ�¹�}~�#�q�گ�(N����y7T3<���lz�c"���)'?�:���8d"�A�

Co�2C�R¸�Ak�{����5�bW�G��5T$	�E]��-�뺉�Z�Ã��89o�a���!�׀��͛�a�5���-OZ���Z=ޡ'����%��1�� a�n����/��a{5�C��X@Z_G4��W���W0o"���~oàU�:�!�/H�k�&bËg�=4T������pև(�:i"�!��^ʇ�� �L�0`Pa�z� ^7à5�>�X�¸:�L�0��Z�;��ri��Ɛ����4�<7À�P�pB*?,�[`����-��GHz��kL&b��3���6X<��g&b�{Á��C��x�D�PP!'�q5�k�&b0dv�CӰc��#�1�e� ��]<\��+11��Z!���b#o�a� ���z�J2��[`C�)�Y��z��o�0�M�c f�&�k��+ۈa,}Q^�fC}�����1P�!��.Z��f=o�a�V�<�����]�����{Ɲ3�!7����E1��a�p��`0�c�����Bɹ��l�0"!B
̛��/����0����o����(��2�����xa	��q��_o�0��*�W�����<o�a,U�Āj^�ع�b#���)��R�y%���җn�7@��Oڈa0��
2@*��5R1��uK��wA��<o�a�G%����K�d��-b�3��ᰃ�4�x�-0����n:⃔<&���%�;pt�͇qrPao�XCߐ�I�t֕�r��Xz�x���[��Iϲ��w�Z,]��֥��Rw�$�_�Q���d   	pHYs  %  %IR$�   �eXIfII*     (           >       F   i�    N       %     %      �    R  �    ~  ��    x       ASCII   Screenshot�lK  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:exif="http://ns.adobe.com/exif/1.0/">
         <exif:PixelYDimension>1662</exif:PixelYDimension>
         <exif:PixelXDimension>338</exif:PixelXDimension>
         <exif:UserComment>Screenshot</exif:UserComment>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
���%  ��IDATx����b+Kn$����r���f�����f�i�m��,�(���@ �)��3�ͦ�D��2#�@ h�駹,�y���Ҷ��N�T��/�0���Q^���g]���yL�O���g��>�~��?_z����~��{�z�=�vl���/����>&��]����c�g��K��>��)8�+��ֵ���?ȱ8�y�����t]��+o^녟����k@�;=�<�{UV���Q~�Uf�)�;���������b��8w1浭��k�\������1��F�n��ֳ�ɦI�D/��+��4�a��M����M�,��g꺱��up|�5~�{�9��ƞ������>.k�k�;/�x�n�-ϝ�<��a�	��z./�I���k������^>�/�k'��/��<!.0��%`�.8��|�ȟ]�g)/���V }�m\�W^����<���B�nB�
���(�~˵�X�\�i�r��m�g{�׮�*�n��"Hl�s�z���-� Pci�3�$���P��j�Y������`��Y�� �uRl��
��s^���k[}����4�5��s^���|H�����Y��=��'?7{���WS���1��%��ǩ��nD�{��n�=ޫ�x��!��s�����L{yPy����ܗ�lUf��q@[v�i�޴*��S�vv8�oi��_�j��K ß����(����d�~˹��(�z��1�d˖�k��h�5?����//h�����! �8����R�;���ႁR�K� ?������G
58m��B�Z��n�<�	���j��MWe�8�U)�R��4,L��?��)��)����T��� N�$��(���ܸ��
���p����}�����s�+����m#���i�Z8[���D�lw������{ �ֲ����"'@^[d�,�#���^;޷��k�{���k�/���6�y�<.�ւ�З�g{��w�{C|&���u��o��ۿ���?������o|ӞgS3H����c�'��� �`F���Y7&|��X��
H7�NVo�q~��<[ V�Tޜ,��z�d85_߹�r�s/�c��1	��^u�Y��έ�iD5~|������aT+y��O�ʺ���f�ǹh��GL�Ȧ�2�j��\^ݨ�����|۵���i���T��=�k�齯��kǺd�_�K���l7��wm-�kV������6�|���]������w�����8��rk�-0�vn�sE[S�ப�V�b\-��z��߬�K�Z��>�=j=�����_�O�Q�����p��{yi#�s�����5��%���r�Sv�l��i�s���n���X�u����j�v�a���	Hi�ft��K q�Z�7%>�X��ސ��e��}\������?_z���fs�����=�@4.s�y�f�����js�ڶ�o������Эq�;�kc~�ҹ��o���S��֓p{+�.[�d[�������,�:,Q���9ߗ �K`�?%9=��6m�eե���[���2��XK�{N�w	L�g�ݗ�+(��qG�� �k�*�V�z}�k_�Z��Ā����D�@ʓ"�:�����۽�1�����*͏k`�?�__{ϥ_��㵽�;��ݯ=�Yp2��+V������U��k鋅��V������g��va_s���[���}�r���}S �_Ӽ�0s�>����`�ãi�E[5@ҕU��LJ�!��9^WWB,؊!�J��$�t\��	�?��.�g�_j�����Vhy����w�z�cE�����ϥ�9N5�.���Zq\~�	ەh�r<�N���<??�?������j�� ��Y�����_]x�I�M���Z�[�Nke9]�ޮ����]�?�o�&9�,�8�8��{/}�{�_�}�Vvv��h��r׬.\>�}k!^;��{��9,@*`*^SD�4P��"Ȗ���z��=��ɭ��&��ʏY� j`����Z�[�����P���p��5���⸎��7�n����Rz]�ȑ()9T}q�/?�ŵM�T��۵�aU�Vr�ĭ���o�z�~H�<�	,�e��+@���ɟ��ׯ�Ŀ�z#z7��U�eS>,sp�[��53>_߻5���o�����߽���O����um���)7�-E���^s��0�f�^�k\[>��Z�Ǿt< �C����kns�3S���]�K_h�o�Q� bx`�������
8���K�~e����k���������3�%���#t�M��ſ����Ks0oa�V0��B3
 ������?|/���hQ|�߾�ͫ�h\�5���M��M�$-O�(�_�|)����<��wy��ϟ?�u����o�1�y�d�f{[ �fM��[^7/���������-��g����}�s�&l������|	���T����9]Q��D%]�����߷�l�� U�iT��`�}�/��z�ƾ�t���J~��wN���[��Lpk�*p���פOЅR� o��c�y.�7�YH��+�R�V��D�=��:���� 8��������[����������bm�������f�P�������{&����i��N���@1���|������O�������/����xL���% �����e����v�̟�<�/��[�,�j}~�g.�|�k���5k��ud�k�.�5������\�k�5�c���cѵ��5�f���Tt�/9�)}��
��k}������I���3(��j<m#H(r�Z��h�E:��� +�\W�A28��]���փ�Au����9�6����[�
��������A@���S9,�#����l�jL߻��6�µ�7�W��'L�.;\wX��<� 
`�k����(�v�ǀ�[`�.���|�^r3.Y�|�%���?�|�f�~˱��sڂҵ�o��K����K����t�����k�@�;[K��wl5�[�즶l"��,hM�8�9Rr��A�O��r���c�f�͓Y]�����9 �C���[. �KPŵ�v��7��V� �H�8��0���1���XO���vӸ���Y���Ҹĸ`�������lN?~��\��sMA}����X?,�mr�����=$x��Iw��' V(�F %��g^(/&�y������3@�w��@���U��G����k��%0�f�^����~.�k����/�_�^�����2���ZxϷA�Ks�7�ɬ�������۱��K�!;���1�L�4�8�2�b]?�%0EVT���V�1S�U�i,���(�L5G^%jIgQ�֖}���΁����<W��(O� S���\�E���>N���_�"�����W-�YzNr}�l�%uu�E�oR� r�t��{��xps�h��.X�E]r��m���3~�[�@���\��luw�k����ϳ�a[+����e����.Y��6�Kחݳ��l��K�|�\��˟����f�G�:�Ų-�Cω��I���E��<�܀^�����q�	Ƹw�.��s�k JnځT�$���V�<�H3-�� ;��W�w�1QtH��Z�d����F@
�	��p���*��_�B����Q�����v��`��	���^�e{�(,�X�kq�\Z#�<��i��Vf��&���Z0�I. ���������w�iN�j!x1h��H�AVYH�5�E�W!ݴ1�y4�^}�U��)"����rIULT'�� �9i+�]-�q���Ť��}��|��)i��-������@�q��Q�"���@I���>��ܶ��������ww�]�A^"c6�[�q�����"���:��"o܌�F�ە5��3����'rs�3�<��%���(�n�%�F]�xv]XB�-���� �tVeV+�9��t�_ɽ.UTh��'���yۦ�u1����Q��K��R4��߻�b>v��J�s��R9`QzTl#�Q�}�s�d>��+׬Z�h�~�]O���HYxD�⨹���0�vlU)�q}W�[�ꅠj�s��r.S���㳸��>�ݻ����$� V���-��$�;�QO'n{6ĵOT�]3D�,����iA�_����?���_��%2R)��^�L�����տsʕ�P��/^�t��I���r�粓ส8�g͚��D��A`o	>Zk���B%�3G�H�����xE$.�m\,����q2�.���;�Z|X�zUD6�:�:�����\^�@��S�}/;/������tNހ.�t�G\�|�`��r���r�q����=Z�L���x��2,ݻUw6�1�]��l�J�4q&�%DW��@�/7鵋��%F���B�a�X4���{Q�h�6_p�8�����=�\����3q�x�"=с��5�+xb�XH�gb��J4������&��f@������9�x-�_ �����'z�Ј��p�;1d��s���/<q휏s�N<��l��x��������������OY�쨁Ù�����7�r4
�՟̒�*�֪]�cȾd@�	�믿���������?�ub�,`a04��ˢu�{^�"��dd�_&[?�F��P��@�������V|=,��U���t�67��|��y�Eۗ�2��ʀsX�mc;�����gV��1&&wV��cnn���]������J�����p����\�h�X�&��.����bjOgD&o����r^8���Q@��'ۜ��agr��r\��g�P�ƣ���SY�B��p+����mX5��,��QT����y(��Ţ˙sZ�M%,��\�ae��Ƚ:��D�X�@��u�ߍW������
u�U����\��w�H�7-&��������Եt�k�b#S���5��#�)�4ʆEQ���(*B�����ƌ�ȓW���o<�5�������h��6q�
�
��F�2.�����'�F9����
N���{��y�0?���8��~o��A�Ԯ�V3�k�|���N��_�o�k8 �+����H��E:{=l(��)�� �H.�T�Z��A ��ڐ\ x��鯿�Z�d���.�!7S&=n�IM��tu>����d֠�v�q�`��ЬĐ��ݻ������?���u�1i�]'v��w��n�I ����K@�/׵���r�K>'�N8̱=���q}�D����r��)�NE&%\��[ )&�k-�EKւPm�ܲ��j=ʎ�'��\����T�`�y�����ή|��w�qM��NT���R�\�2隶�c�~<?�eAcǵ �︻�),��;��[���C�V�.tq\Xj1	O��H��Z��4 j.�i��ԂýQ<x9f�,�Zh��$D*��`��[�7�Oq�Zʹэ�	�?,dl0��5}�t�X3�6{ә�8�}�^��A
�XE��s�}�W��a�Yօ�����4W2Ns��}�!�A �[�Ê"8�U��w;y���{\�����9�fe Tc9)k<�6�c���e�vK4h����*�B��������������1�$�f�	zN���`��/�8�1��fhM�em�:==�el';�nj�<k�-6�v��*7\���' ���x����_@�m�5 ��?/�ݾ�	�Xz���2�9����Ų�vbk)�_IA�	����c�����0 ���Í�V&�y���E�3�(x*���\�-�p7����,��I.���ݸ�������r	d�zvz�.x�w��	��q�������]�ܟ�T�!u�.��t��sc̰h�Uf�HĶRwJt�8�Y>����y�Bw�y9�mo��.s���nnj����:X%s�0�]���F�C/��kx�t�ټ�'��~T��*�� �eRY�zϭ�W�{��4��{d_��{j
�1&������\��,�N��Y��܃e�/ks$s���z��4���� ���NU��G�	�t����|1�a����ʼ��}	>3|+��5fh���)�0�u��ū p�:��y\�r1ޚ/��*��Dj󎻾[6�[�4�����˸��&���.[�!�9i�+���7ޡ��>Λ@z&�~�,�������ٹ;l�.�|���I
Z��n7L..���ﰨ0��� �#��d|)^��;n ]*LG¹i��,�O �e2"�@�V3���l�o�-_�.���pN�Tª�
�T�����Od.��Y�j�+ ~]6'<�g�Q���_��X�ߗ�~E�د��u!������2x>�_����<?;�M�O-�
��/^ �Y�j��g��C8_|?����tX��YqP3J��8W���M�Z<�i0~\i	 ����<qH	���])�+[�'x6���GKQ��,�έ�v�W��R��)f=�}��bƼ�XBM}�J�:��;c�bQ�{���㒫��������X���|��B������&�� oB��s�w����ߋ���7�W7u���Ÿ�g ��`G�VL�e�T����ͪ��w�2H�vIj�����h-͋�1���.@{g�����)f���'�y�c�(Ć�sU֤]O��\�Jw������c�� �".�^n��;e�H�h�%u��0H�X���.��eq���-���?L<�@�w7�X�}�w�Ggّ73K؂(�5a�
w�E�+��d����.��k�b 7��������f�Ҭ�����(���f�H!4l_4ݪ0���p��Z��w���������o2qZ��1I�;��^8��U)��1�O�X��S�@1�!�%J��ˤÄS>\-/	&}��8��i��y���� VX܍�	�; އs�Jٰ����+?����+X���0/H�)�����W����{�y� �r�O��86��x����������<����\	�3fH�h�������|^Y� ܤ�(��ȇ��#��ViL`0O <}���픑m�/=@ ��oI��u�t���4������p�ܴ��R i�<�	�"�~XE�{:٘H[�"��tTSb��>W���Ov}��'Z��8u�Z�輺�?���J��-C��zh4a͐�ˢ�l�2'�f���D?�{���_S���$��w���VwQ��W%E �j�H�뱝ޅ�EwSXn��oL(��N&���4��l���jQ����yH
�� �ާJvsq�d�܈E2��]�'��؝l�0�p��ss?��t*!�k 5��1+B΄��8l��y��˧f� ƞ�w������P �Nґ��t�צ�h���PЍ�@똠{��7��M:��P�샎�͝���"R�ND$Q[s[=�t�Kc�, �QW?b#� �	��̡��ks��J���������X r�đD������V�S�餯M�@��2�m�K��z�R�Dc�6�D������D�ʊs �5��\<��븩wb�1��ʔ86O��-��w�۝ݍ��k�!��[!�y�@�Ojk5q��x ���U���Y�,\@����NoQ�������Q��Z�x�4w
��rW|�"�������"U�Ckx]�E� ����_�R>�~��@���(�0wZ��p~P�B�9�p�����?�M�HA-r�EQYvS���%��K�r^X�p�>��I�ߋ���I:$8&��fh�������&��^�9��WKe9�r�ɸ��� ��N�Q�*��5�a���ir��%�`L9Nuc���z��|j�=sqޝV�0�Mp���H�1��-�b7kʠϢ���Y�lŮ��&�N�,!\�Ԙ0kJ^��n�s���s��@�p}#z7*�!��W@j�'�Ż��&bR:��+7V���`� �2�b ��� p� ��R����\e��J�R�pKq�l¤�X� p�V�%�v��~ۤ����u�z>0T��`o<�h u���4���H�����eó]����A��ė�n�77E�[��l�٢�����q�w:���%.?aA�E�I�T4�J4�	|�#��6+��j�u� 1��]'\�G\�&�� ���Y8IR	ʙ��2 ��7}X\W�Q�����~L�]�a��G$�Tk`����hgsC�I����*�����{��r���e!VP-�Mڗ�Ȣ��y�I��E�� �y><(?��a��4�9�ɤ����M<4Тꁮ]��l�,� ��W����Veeҥɬ�N�Wr����e]��ﵕ2@G9���c�,�we����ǯ��È�9<9�A�-�&)׃~�<W"|��8x	�ڂ$ͨ���N`�;?('~R����o��:��jZ����ѧi�8P�#��g�;}	��Nܵ�C�_%�P����7i���k��=��\�5���Oi�5)H��g�����5jr���Xy��,�l�V>�z�:�2�h��B���f�7����Z�;���v�ɢ���EJ^�r�;#�%�4���g&��]�8X�@�4�K��3J��߼VZ���4I�~c�s���� ��]����ν�t�8(�bz6�J�gJ���ANº�>BS�6��dt�ܢ�~����g���4��$�d4��>�7��Xu%����<M��u�����vu�޲X�%o��ZW$a��X�hx���m�7>C�oZi�l(8�<�Ώ��,�#�nl8bɎ�G�u�v6����GS���r�B�D���+Ξ����u�(t�A��g�<����m����p�SA�Q�LK:W��%)1�j�{Hml��:�je�ǖY1�"}����ϕ��=�W���u�q�5"w@Ć'�lq�������r�Gq�(�厫)��v8h:'O�|�=̚�����ãg#�f��%&�,��)R�XuG���s�ӈI��8Bja=�ƀ����>�DA�G�9�S!]bn~%�3�טe;�({�E{6KB9���D��e��� � �����Ь"U��U�����&���h�Hnj�,��63+؛��(]�n��F����>XY��,��`)ugy��V�����5�4��yn�腄��C�D��4�Y1��3N.��$P��k�ܯ�=X�'w���u��믿-��,���1"��U�a<�s6�X��{��� #�2 m�����Y����p^�� 7
�s���x|f�0S�*�nE�)��poSp��*7{��y���{�(9�9��֍S���h�u�p=�-2,�T3�|��W�)Ċ�f�Lĺ?{���ʴ����;�M����&y*���#���EJ0}#j�rP��/��E&ԕ���s��Ee)��f=..�ނK��� S�KD�6�1uy��}��ew]���&@�I�dL�[\��;�t%��I,5F�w��gia!Φ�"�"Év/��4��d��2^s��E �IWn�gW�ke�G�7)6�tA���Z������}����(�=��g#��L�o�{#V=lt�I@|�0�W>:8�
?�����bs.80Xb�E�u,)���ҹ��A��{s
�5^w����g�\��o|>0�R�����-WK�����RF�����{Cr��7t��.o�s핣5�^@ײ���������s�^��H��1D T�#2����i���G�}]�s��B8l��v���=׬�,*5��JhQ+A�Z���v>���j��4%��ܑ�c^��5 \��i,BO��+źtci��w��Bg�5�@�A��n��ViH��{�ʟ5�?V���X@��ʭ�j���b}q0}�"U�xp��w�Y,mT���(���WΛc�&��E:��"w��Y@ԄԚF��p*���T��2A�1 �U<,�2ɊEtլHD�L�T�s��'+%*X`��������H�ĸ�HI	��]F��F��V�2���`I����Y�Q-��@01q�,RKR1qݪ�8�4\B���3��RY�p����D��o(����΂߳-������΢���n2g�:)ťX�)�<؂�v8�BaU t��7�)�j�ߙT�\�2�R����?��P�v�@?K"�U0�ň��i���;���H{I�T�F�饸vl����;d<�77cX�C�s颟����W�d�$b����hWXM�����P�:���)�F�>�j���N�A������3��h������z[ߐB�kB�3�S9�弻z5��G��'�c
dAUּ��0֞:��d&�nm��`2�u�tm��M�����7���|C&^gS�N����.�*������_?���V3o��o��T �D��CuTy���J�;���$�fՈKb�[�ƩК��s!�[dTS���x4�B'����h!��u!����K��+~G� d�$t����W+iΓ�	,sG�=E��T��VC�����g�	PGը�V�	�6��F���k�T����,,)�;�Ɠ�.Fd}��-F��XdC�J���R�=6�\�LK���Xq\�I�;C���E��z�M���g��v�`�Y2�&qh����j�����`��s@j��N��R*�u�NI��#��0J��V��7n�3Uz�l ��,�-ad������Vb�^e�W��mSWHH�A'�@�.0=�X$F���%QX�7��,.?Y��˭���4EJ��uT2�[\�r��7<2G���Ez	L]G���)\=�|	�t��b�Q�"KK�E��Rɓ�Q�!���E�o�trkV��a�ź,�nq���pm$U�`�MѸU�b ��Ȃ���H[*���!�q���"G�v��q/V�B ԕ�|'�,�K8����T�F�����������82����(�H��:0p��9�F�;<�1a��/��Z�`�z$9D^�2y���?	� ��F�Ct��]s9\�\���Wǆ��@��WV��v�B���Ϝ\�	��@$g�c��3��͛��T�v�sg�cP�E�=��<{K/1XUZ"n�+W�o;�!Q#g���*/��w���w,�䆍{�h�ws��\�D�l |�9X����1���XO�҈�M��97�т�b�@\�����h�'\dۄqg +X�4�ߎ�Ȣb��H��t���*�p���{4��V���ݔ�u��ؕ��e^!�l��KV��1�?��o(�,n��0�+�!��	�­�<��5�0x�L�^ ���}��u�7�������s�ZN�P��W�|�Ny
�a)��u҉X�@A�IGwe3Hc���\���,�M��f�9\�b��@�,���ieV��&f��r�9F7[P�rB-������W��|�ʻ�;�wf�<���r����.���ad>"���2�(��)M�8�Jk�剎�^N�iLo|��]�|�jY������\�4�0��4�Ҽ�^u�X49�7��������)�����fM��ߤ�TH7���h��Tk�=6�O=��Ѭؓ���=�N2�\��9���~���d�q0MY ����2y��B��lƣy6)�P����Ò$�B+��Xs��qTl��\��-GJ�"k��k��A(肷d�#{%t����{�#N����D
��kuR�à!��Q��Ē^�Js@���I������Ѓ��o+p�Bxp	U2�9I�*��e}`�a���R
xYt�TaM�X,�&?�v��12L	P�2��-]�:�QW�N=X�yN��WR�B�Yt����3�i�3�Xr���O9'�v�)G�׋d��Z��ӓ
/Ƣ����̽�H}�ua%�S��[���M eAV�R7y(ůW�?�hI��qZQ:��Y��`Jc%�%��@��݈��q�S-QKv��&����F��/�-�_[�杏/�W�~ P�����\��3�r���%;�[
�,���K l�C�u�i�b1gw�=[�>�{I�U\ŢT阧�I`ρg���Uҧ�P-6"���[]#Q�F���h`��1�RH�[��i���p��m�&� �3��<��{���:�u���<�+#<=�d���~ٵ_�O6Xu����lN�7լ����Eц�%C�v+�>8]�� $f�<�kf`��뗯�9F�]�ٶ �)%�
��U֊�u�n^G��J�U>�&�t$����N�>���8cӤ�!� c�͗A��GP�)[1�l1M�ù`q�w>)2���/,D�d>�$��jVR*L#��U$֤D��Ľ�h����^����wi�p�yNV�lE/z�=,>�G�Y	���|@c���be=y��3��{\/�@j�&��l��>R�Qi�t`����l!�)rO�{�fM��3�MJ	"�Q��m�iu�3����5hG�ȍj��J��w���-竅N膻++�r�EPh��C�`̯�A�Μ�`R6S�U,A�Ӻ��������
ߘR��u���)m�e��K�u��Tk��������v��^��d�Egu���r��g�1Z|��-l�W��Mמ(Xj��쓆@jBw�529NP��5���u(��M�b'ǂg��87t�1PR@bpb��+���=V��o�0�Vid��pcΟ�,@�,��dգ�:D��\�]�.Ό��k�{g��8v���1��d�E�e!-�딲U�2�H����'Y��~PW�$ORXD���� �[Oo�9��]��6�k��q�|�&�ʹ�4Zh��0o�	u���(0��)o���u��;6Nl�qM���� @o�l�p�nM�U.�@��1Ƈa�Q����Qa}��[��e�H���y#c�>xU�W8wՌ>ʆF��vjQa��z=�\�['d���jU����$t˜[*үM��)�ԅf>����cLG-�"��Nl�7M�T��s��^z��I�N����aD�u�InJ�d�<.+{�n����ϊI���d��ΛrW��e%�z����8��A�z�ld�H��N�:�6"��8[a�~�1K�k��h����U~��]W=
��!���]��wM�S'Wg�`�9u���z�(�h��^um��8gr~¶ksT,�k.�˷�h��;���i��*7��c�B]�H�+V������do�z)`k�uUu�1� �� �ǣ�8�Jj���"
��x�.�)�A�J��<�Kmջ��?�Y�CZy�< �?� �B����	�zGL�z��廏ߋ����</�S1`�nS�o&Q�1_;M�|R��5fa!Dq�,JN��<y��}�(�w�ڒ�� C����|�.k���cI@z0Z��Q^k�3�$�ۃ��a6y7u�%��4�FU��,�X�A���"�4C*��+W�T�v%�,RD�ihy�H~�z��Z������r�L�	
��U�ȸι_�`�Hg�71��zQG��~5�ֻ����8^D]7.�e��јt�[�.� �'.�I�-���{���:����6.Ց� bGС6m��b-g��)���ּl��PLN����b�ձ�����=���E�^FUE'��l-Oȥ��dO�擻kl`G+OK�=�UK��2zͥnl���4�����h��ڂۉM��A�� 0)����`���Ǧ[E���q%n�zL 6h�s��G�\:��;1���3���𜬯 T�<[:S �|Z+l�!�c7�S��hp�qa�EZ�
ƵG�w{&�d��C�ylNz'V5+E�j��pݣQM�)�qI`��1��#jo\*-��5� Qjk���i%#X�ˁQlL�9-��Ѳ���jG5ـ�h��$F��^��3�7*R��jgJ�� m���޺|̰`�8��dԉNv�0�v�e�?��� �,��}+#�+`����+�|��3���[�GѺ��/J@�&-L~K�QHY@E�"�D�.����e)3N��TR��,:���oZ�q8x�s�����I-��zq���4��uU����$y�*��-C�u+%�nk��d p��<�� 0k��cD?������H=X݁[[�fF~�Q ��9ϱhzM& hb`y�K�Y���+/Ӧr���Q�jj5.'����b�aQLN���,���lW�|:z�F"݁{�1
%���$�ι\ݤ"[k��&�Qm��hiC�0���$dHu�G��3M)+ҷ~�O�*�L�A+6�76�T�rȰ48vS�[�bxo���

��k���4%K�ܻ��͔�A�{��=^ǵ�������WY9H|v��=ߝک�"�~)֗5mU���oi�j����d|z� �ƃI�Kو���3zpNL�Y��q��Z��˒%�h���!\��5UO��]H5�;}��En̓e�0XE7��(����q����P)q:8��ߛ[�L����Y>9w(E������ߍ��)�	���P���dV-?�yb_l	�,�,vw�DkYw��R�2���Q�1'O2z��}��t�GK	�Vt6���F&�&V�;4�Y
N/@�q�~�J���-uQH���;<@�Q�x�����W�`���]������������1S��mL��HaT�ܺy�g�$��8F��AwS���0�J=�1��2uS������,X�n��V��ƀ����
��b�bĸ��ܨlɖ�[�9�Eԟ-0f����-/����<aHV�g����q�(��Z�Z����r��
L�.�*ӱ/aP/��Y|G�H��=�B*ы�B�D(58�=*�$y�0$�<��W݄w����G�E le�f�h��9vF���:5�%yb���&I��f�>�&�����R��n>�%��S7��AK�ꝵ+p�xN�o��c�N���k��XA8w����P[-yGk˅ģ�:�Jkͭ���Vm�B���g��7�l1�YE?y!�;N�$������cX\���ꏻeUp���k��A��� ��nR�{�4γ��6� �s��xc�U���y�X�s��j]�ʶ�u��A�k�4�9s�+Yފ�� |�q)M�ͪ�ַ��Df��Z����A}�b����c�ƆŢ+���f]��RF�J�,2��f�'��FY������l���Y�ō1$j��0Ƣb�����^RF:f�S���U�Z�h$1+�����̳d�5��8��Tۚ���VH��Q��-0 N��d�W�@qk+�/���0t6���� �\{J8L#�.��Z9$�彰T�O�r7�VM?��a������2kA��/J��J�Kv�s	��{KM��� �1�Ѣ���/���՝a�5ъ���X����;=�E�e����X�|�.��qZ��� i�d�3H�*g&n�l�뽽���Ƥ�5	��I�{��0
�Un��L(�? ���8GX����w�z� ԭ14�U��c��/���&<(j�Gԛ�F��ei����2�E�95�7�T]h�)=˜N�(�\��������:
��y\vև*m���}�0�D��2>��Z�{���v(�(�B��EjD�`4���~�����[��� i�31ù�q�B����N��7� �;K)�x�q]U���p�YmI�NZ0�����z� �~jBWT�˼lB� �����`��:����gԞ�Y=�3�|.${t�W<���+ �&��nQ��ݬ�6n�r��ɕ;�B�q ��	����C&Z��n7{��%Z���,��[6��ƪ��zDo�H<>}Vyʤ��rJ����}^����k~�O�/3�0W�y�k��	ԭ@��Z O�#o-$����1�;�;kJDV��X�+�DZl�C�Zڤ�e�"+��à�.�g԰
>+Qy�q#�����h����x<�z�t����T�T�� �D�����_ʓ��x?�4{1,���RWUH�,��VJ�'%>�7��;knҥW~�%�� �ȝ5sd���<mEì.���f�^dk�{a��{���;��"	cd�	��A6.�@��U�vο�c L��e� ]��b;��,�<���Q��NXJc��n�	�Z��d�vֱ�Fj�A�0K��:����jӞ[л*N����M��r]�K �� �y���f=5���װ�eY/�c�����k�6|�\�U9)�l)tQU&�)�KV�v
e��f���Y�r�K0�)�����Z�z�H����D�/�������4S�m I�x ا�Hy��
g��eAU�]Ŋ�R��@��w���K��VO�����9�k� )�SJ��Z�J"��Y�T�7&����Bp��E�gY3��tk�QX��ts%G�ւ-�ъ~,��_�_��/�?��?�/?�R���ߗ�֪���{F[��sDe'�����|�/_�3�j�Q̀S�i��G�g̀(5no�zƀ��)�Am�`J��`��q/03Mn�)�]���{&�Yu�Sa�I�j�"�lC�tV�[�]��9l�W��3i֝|'�+t,@��֊_���l�2ԊSy��McL^��S��<��Ϫ��(L��ܛ[O����h.aOT�m��"JRL����lY�B�9;�2}��D3��Y��g�B���'��XmaT�!K:�.�f�f�.��
�L.L��z�|��^���~K�K7� ���
?X�6�#��h�.�H�l�f��P#(n�Is�5	 �`��T�B�;˂'���'�,�n��̈;��i�I�`N�W���fϓV��� .�7(wi���Vζ�J7��.��9��N�L�G@��v��㣧�>=j�nB �,�R��tc�10:�{s�q2le#R!���TV:��π�dӉ̩�6��-Zn�H�Rq��*=��
��|��]�kp}����Ze�U���q�+�Y܋�0��b)Rg`yb�b3Op!�נj�ɏL���%��0���8{��������%n=�nz����N1����֨�+"�>ͣ{�DşE�f�2�ڸ��.��ծ�����}^�D3ff����E�֤�������4�5c�.�Z��Kr�I^�<W����D�����Lg
�/n�8?���0xAj����U0z�Q�Hd�<.�xy�^*g#-���NNO�J=�Fϥ8����T�j���P��Z2��1d�
���/,N�F!�3�&n���#a!ª}�,.�`Z.�Si�ڒ[d��62��STC/v^��d֎���h����|�H٤���A����6�q��ĵ|����ճ���H91��j����¢��]V=װ&=e7)�;][G8��Ӑ:������ާ���1�T�l�,�ϙ�a��$6�\�����ؐ����C���*u�,n��_�^cl���`�֑Qd8.��֩��G�Q��9:3�^�he@:,ލ��d��9f��-�
d��r��O�0��&�4�7)�����t��ǟk�M�2��^c���Qi�:�*J�i���L�7��AUf��	=s���6.�4D3}`�ǀ˚X%0�W�_|��R��~�W�b�u�'w���]Z���lwf?��}�:��Mz���.P+óT�r����Uf�7-��ohU���цc��5Y�Lc�U�m��&�`���O�N�f������?�`����i
���M�q�B.���m,m��(�L�nj �a��:��Lw�^���dAS廿���g��o�����U�f y��/�$���%�j�U�u2|P��epP����#�f̖
L��,8�w��+ 5����J�����\48�O?�, 
.����HE��s��A"2*I�T״L}��!o�ns�@R�Dv�H��to���d-3��ʸ��M�.#�b��rՠ�@!t�I�Z��C��y]�y��B��x^�esր��M���~��8�Y�P�����`�E(O+���z�s��u4s�X��Y��	�x4�k����,�UZm��E8�h�ؔ�TК�u��Q$(@�4�nj�8��-���"�G�������0L�

���g���嶀�cN�7�~[�ԮZWB�P�)��t�q���lLr����Z��fK����8M�*��1�i��za�������W�v��u1z��N���0V�ųq����hG�c-Ց�~&�#um�:���S�@-�.�bF��8k����[?��借O��#���X�X�5��k�E�g���53�q,�=��,�Lk}+�ք��DjsX���d�)�!�{t�p�4d4�^X����Y�.ߩ5���>�N���T�a�W=�I����5�9��U���,KĜ��#�ߞ���.-�� ܨL?mr������Q���m+kI�k3S]
l���
��XV�{/	���ݟ�(wH��9콤|���xD�Z��\b��Qj��s�7@*��z0I�M_�~r)B�j�[U1h�iDfu=�v��Uu���b͕/~�e+����񇳻h�s���qe��(��A�c��t�f���'�8x�(�@F�%ɓF��J���8���I�����˄�F�(Y��e����X?���D���&s1���A�@�g��_j�f���Q2�f��ꃖ��&R��� �Cr�U�f]��z,`A�m��u��бӂ�8W\�ϰ���u�m�*^Z���tŕ�iV���D�ժ$q|��И��#�ުE�Z���'jJb��o`Ѿ{��GX�����
��8&b�Z���D~o[*�;كbO��O�R8&�[��ip��*�SA�\X%l�é�N�`CňeԅEF���I��#�yK�,�"�>A�@��>s�Z*����'(#�ͽO�i���։w!����pe�&�0ŕ`�>o+�8���<��aH�@V�d5�q/��-���+������9'�YM��k�(2�Ze+�$k�nb��53n�B��
Ms���`Br��1�T�}ZU�Е���6-�'E�z���R�(e�D�jn.�w���0儤���,׶5*}����h,�§VU���^R��`I���n���,X�kSb�B��,��RU��#��/�
�Q(���7�����\�����//� �K��%*4$��,����2�S+X��7����/���T"����I9�k?�6���!���߂��
LG��3K����H߿��)8�ުJ1���\*�X�u���A���-��l�Z�ٽ�\������%$��9W&sW���Qfy�d��*�j;/�Wl��g��/�57\׺ �I[����g�4Cm2�����I Q��䛼t���0̩ R�Z�&�?������+�UvΝG�c-g�U3�M��Ґu8q)L?��{����
A]U��$��ie�
��.|��2��V�@���w��5�
P���^p��1��߇�#�D1�s�QvlX2�|��m��!��i���FN�_�-���y#��Ux�Uޙ��\o�]����V��BP�����+����Q�:�dp-bLD'�闉���S�^h��*�ٜ��ֽjmյU��9�?J�S�pm:���dp��f�7wB�@�`�+
*cӑ�I� �	lN�e�V�ѽU[r��	���~,�BE -R���"�5�DG�������/�������
C�?G
l��Ŏ���,�y.�<v �M���V��'��E��J~s�}�r��vQ}�Zе�k���v{��3P�uD�i�jO'si�
_ZY�i�	�XU&�RU�V��k] ij�X�ww�N���;Z@�-�iE+ú�9�L�TË]�e�R����I:,`^WQx}^=W>�d}Lۙ�|e����W�?���s]�d���Y�\����u���j�P �Q�����o@h�������Ug<����m5�V���p��%4�&��}�}�r��Ҵ�OG+�i�����e�P	� 8,�&����&CK���y3��;y�ܓK_�-�f<r�V�{���#_��a�nY�8��"���I�b�,��%��~!�Xu�s� �ј�[S"!�8Ǖ:�Z�ɴd�R�O���=+Uͅ��p��R#ʂ.����F2\o�eWҞ�Q����nnҷ�f֒���M�"�Qu�D��*U���J$�?Y�G7����:q��E������1�w���&OLtP��F~�*�?�e��{�˵b!j��N���+����i����{�R��d�B=��U���7�H��ju���E�G�r�Խ2���6~�|�\�Y�U�aډ��e��#��<�)d<7Ԉ�:�kZ�zs��y.U��Tw�դ"�(��+��cʂ�1�� �E
�ZJ,ڊe��9,����l˛V3R"�7��t6e�hJ�`�Yp�E�,<�
"��A�O�H���݈�"�-Tmf��a�����0����ɭE���wnA=��m�j�@6��	���X�6y+
���!V���/�>tڳ�ru���l�ɩLv3��n][T�A ��L�0�j�)�V�g�!�ՙ%��<'����o�2H� ׫�'�5�1��k���5�=�ԥ��Vyp��b�����:��B5b]&0�*6�۹wŤ�,�W�cq0�x���*<5�)�k���i�JMѲ.������1�;u�m�t�X�khr��:Vk�*�5�G�@W��� �a����P��8�����!����Xz�ss/���H�z/k�q��œ�h"� ���*��8	�h��¶�2(Js�P~�XQ���:�t��}��xx� �H+dI��Q[���h@cwc���<�U�#��MC Ъ	=������R*Q�~'(��p��hP[�"�VZ�V������h�7{�v%7?	��[�Q^�lhў�>(�:R!�),��:^j}�Vst�<�$��`%{o)A����¥+���wI���ɳa����[����M^�])�x��K���C�N@�q>?�����/�N��S�D���P,h�nB6�D��nH�`��2*>n٪ԅ��bv��w�;��r�W�0~c`�9��e��HCɒ,R�Y��ŭ�u��2GƜr᦯�<kk�k]x��p��|p�y||��8����K��h4�E�[x)~c��=�ִ��Yf<�n!�n7&���q�W/SD�9��c�W��7Q�y�>��9/`����]��-�t�e��9u-���)���rvCȩ���;V���xHa�be,�5�CZ[��d1���t�[D�p1WMx+����1�p�N��)��&�6A<e�p㓔9�9�O?W|��u{����cU�(����"i+�4G���Y��(-�!����I܊&��[�J�{h��@�̡�f��of�ϗ$6��Ra��֥��X�a`cD��}�PG�,�GNX,Q�s�G]ʺ9��Y���8H���+ei�P�E�Iq�t^���'��h[u[���ͳ���Γk��	{���d�םɆl�s�P �l���x�)�.�͓�#��A��Q���0m�˿G"�jSXA�zJ��*��eN~��.�_��]y $�&��5�U˲[+֧"�:U
:ywO��a��xqE�^E]j�Uhdp��&a�7I����,u����>��C�����>�A�Fˠi%��|�XI�C�3XXҟJgsۦqW`��{=���;�֢�t�d\�A�B܋؛Y;�7N�2���Xe��2x�.��C��:2��Ff��l���/GQF�Xx|��`��xr�*�֦~Zh瀯 �9��i�.�cb��, ��3�hyԤ�,��"ܨfQ$hKj�Ӻ�={F�Fn�(�.����A
�U-`�|�Ȳp�;��Z�&D�FD�@	dIё;�nխN�9�l]�Ǩ���U:�
�p�.
���l@�<��	��FtZǲ��&C����E�b3��э)Zѻ9�$���ԅ�Gv�ޖ�xOS t�:��z=�T��鰪E���`�����o��&���տ��^�~���@4���{��k�o͉�C껜�]��e�,�\��#�h~T������*� L�>�m���kL`	�����2������,���:Og<.�ֈ�<@p�
>�z25:^�|����-�qL����+�|�؎*���g�Ï?x��Y�^37��vnN^�gK1 P��^���Or�pY?�?H�i�����I-Z&04�-m\�]�G��h�Q��U0p��7��/��p?@�:�i��*1��|8�WQ�-'T�p�9�3
��3s?��IY[\��NsE�|��(w��\ub?-M�@p�Χ��`���2��ë\��9u����Bk�>\Z�4�bU��"%�H��(�{˺�;18�ef6Z9#F�uהh	��qY���R��b�vsW�E��b���jD����qF�KK>�g�0��誅��F��&TJ�H�d˗���4�Qǆ>����os�ݵ�aZ�9pts�ɓINzue���'������0A�h���4�� ����Qg\ ���8�k�v�Ĺ�@P��2�plT����O�����@@�2�p�C/�N ��h�tb����H!�X 	�/�H?K3�L��u'��6�L��Z��QM&����O� [QG������*T�,���� ���yC��O?IU!���ڪM� ��i�2g2iͽ�U:�I��ڑ�XTV3v״��N�-�쓼J�Ś^[���,�.�, `�J:g1���o���^�H#�z F~77jϖ���"�lI2T���"&"����u�E{lԭ�A�"���5��ɁV��}2#+�!��h"��p�(��Z�3���wF=�FE���I6�\E�Y�q�Zc���	��Y�N�̖��[��]�7�w�PR���	�4��3c�T�y��ֻD�/hY�7@�iXU?�@�}NM+M?;��)�x�&��c���亀�
x�Ѓ�ʀـ�.��j�v��tV+�5N"�/�BB$-[	g��,"'�����U�����w��l�ȑ�~Sۻ	���v���zʧTR����G�q	�h>m�h�O�� �r|��7�+
u` D(@��`a"��h&7�%�����L�/�`�Q��{#U��PK�l��Z��.u���%��\����	]	��G�Dp�qM���n	�x���ԉYp�G���8y����K���{� ��
,�_�Ż��|�l���]�Af���=H�����廏��&=I����vvoXUɯ�v���{:�$%�x�������9���w�Ǔu������n��&\�X1���>O�\�CJ����
�J��3�xn(��Y-�z[n��ճ��x�nmv�?C��6ɓp��;�B$��N,�y����}�ׅ�I0�C��H=-R;�4��a�:�:zH���C��]a�M-���ֳ��bra�m��0��r!��:�NL�¢��άOrx����O̪b�G)��xS-�܈��_~v] �Ѓ�R{�Rp�DD_�<U���Dtwv;�k�����E�y�h ��"����? � <�djd��k���,����e}-�ը]ʀ
?�RX�O�ZP+~�\`�bsf`u����~\�U�� Rђ��t��#P�}���} %,;p�8g�����4 �n�%	)c!��j��Υ��[kwV���L��������}c�b$����g�M��F����-v���Ng?�d��a����<�@�|�;��Ki����Z���:�K�֚�5�|Rg 5�TE��b�.e��	q�j/���h���3Zؠԃ�V)ӴRAhp��rE5XrU�M7�y$A�4@�,�c����4�,q��=�A���*�M>���b�±��V�<PX�8�u�9���b��Q���$j}�N�7�5�&�D�uJ�%�F�t?���$� �O
-7}��������̇@�ߩ�UkV08,Bd���X��&�~^@;�I������Q�K�פbύ
�"�-F�B���_��W��뽀($6�{��g�FD���6L��i�5�b�<�4�)��+� �p��#�c�i��P3�f����R�p�)��D��֪w�����Y�&b�~V�h�[�2!����.:��C�R�t�b4��0��|�˿�M�������3�7@�·y�l]�.&顡��:�X�ݘ'�{�g����ʻ5�R��R���� �w�w���0���ØP~��:���`��>��*���	^���Q��T�Q���Z�оBiG��b�.���ޔ�	!<�j5_���F�d>���Tp��"��͍j��kVE���'+����]*iI,���OKR�pcЍ|o���Ւqm���"�>q�K�2!���E���R�쮑q��v�K�o2IKi-W!�X�Y�NԬ/<��S��V�9��S����ϣrdg r�]~��JME�t+�p�Ά�Aq�p30�qs1�-��5�8���̗;�]$�mǯL� `�+v[�*���]>�9����6Њ���R�8����UF��m�`�sZ�f�N(�޳W>�2��ƅaQcB�c���
��N6B[�@�rp���kĽ!7.2m���-h�M���`	|�Jy����$pz�1w�i��<+E�2/�9�s��h�wP��.���\�K,D�����A�,���B�Y,�Ӳ�� ���&�4�:�^���}�ڼc�ޞ���ƚm��oG�K��׺1�f�)����}�'� i��=�������#b����m����Y]m���쾦f�5����Rd<���>&�R|٨m�U�b/aqk��8Rw�$i�d��*au�q���DW/������!�b���U0N��,���E\�w�����E����]��������wޤ_ˑdM;�Kuc釻X@��<���֞�Y�e�b��(nם��p�*�6�*D?X�#�,�O��cY����Z�$��ϼ�7�XȍU��\��NN��!@f�\&V�^'8\0<<3�h��Η)�6���dd�*���e�A�܂YD��>���-�L�k�p~b/s�C�1�E�=ͳ�Qg��&n�a3#���Ζ�v�x�=H����4-M�7�?$j�xG���:d���2W1��yRۤw�I�`�\e@���+bqE����xܰp�q� RC75���ܔ4��h�Ԝoy�ng���^�y�Tk��Gs>��ɼ�aEG��IAɛ��'�Z���p�Ck��dј�9*��,��V��}2��&~t���xl�6��`*��k�T�A
W#i\.�A�dň[_Q�;Z:��<Օ��9���4 ��
]�;͘�ϝX�YXJ�^Ӕ����+˽���+[��.������2]��n=��w�� �<��"���#Hoﴄ��.^k>4��B�+]ױXI�y��~�Nݿ�=(~+�o����y/�}�n,Isi�bU��j�=�d%YQ�hc���p�q�n�����L6ĠF�gPy��$3�"]��	 �a���\)��՟�j�����?��F�s�XUQNN�\u��ffɄw�^����%|}�"Jd;�>���޺�j�r�bsu�{K�"�f���h��g,����mndS��wV��J��Kֱ��σU���Gi�RŃ�h�GZ�5�C�+`���zb\���X���a��˘8��R@�ڼG���jy	>V������(�X��:�ǳ�rKxs���,)�Xa�*iE�0Y���}�s��װ��½̀j��k��6�B��L���0Lf�Х"��Z��}�!y_�동%z�ψ�/`ڞ}biq����j'�(6��6��o=�Y�*�W e�r)���[��Av{���}��|�o��&`��o��`!ii=8m���]_��	�������ಖ�5D�Lj���I����௿�*���_�&էif;d)@�|��I9�`�3�3�PUt�U�A���d���c��Xf	Dq����"���E�,<�VЧ�^7!��o�MAՊA���叿k�ҏˆ���X��ِ�xa�q��R�z��r���x»�}�=e��?
��f�4��Sa�d�R[����R��^Ưb�QՀy%r$X���z ?e�lo9��K)���1k�>X'�I� ��Nb9�
`��,��~\/��ϋ��{��M��f���:�2��FO��F���"`�7��3ZS��e^Z��{��8����5�,K�2��Ԥ��Ȧ�F�d`�cd��`��F��c�R�B��ˀZ����3�E�5Ϻ�Ӧ�v#�,T���"^��Nƅ��0�JY������`�>���j�<��j�P7��b��%j��b�e�NV���p�]vL , �g�|zN�8�d¡{�˿2G6j����Vy]��C77���H���]g�w\��;vo�M��߫��N���0b���+��������ɤ<X�\�HɒZB�<�mϋ)~�i��\��|���d��BP�a#��Y��)YM+�ͪ�l�u�S-У[��4�E�����St1�/�KeQ�ײ�2�Gk�J"���_�1�qy:>zYA�)%N,��H+>k˛��(M�R�;t�˾ؘ�(~P���e���.HHY�y6�F��`�eЊ%����&�R�\�U�V1�wL�%���,O�=�����}�_o���|c��Y�6@�_��6�ɩZ�x�Jg]^?�{���*��lj��N�#j:^X��ǫ����֟�h��6S:�s1�Y@�:k�#��E��U&�7��b������gӊ�f�D����ȿ��7
�:�%��k��gI�V�������U }2@,e��"�`j�V84�+�O�ĞGI �=�Ϊ��Z&�^�N��ں`z�@�Pf� 0y�3\,�����z� RXKHՄ�@J
����m����ZvR��U�?��k�r�6�b��H<!۱��b�9�h6���'��v�¼q.*����������}R�b6����o�L<zDNI:rh+��E��<��rlyz<�<���3���/�)	ܠ�
6�O�d�$��9���l����7@�g+�[��$)�''I�/Q�v&?],ӰV�K�=�(�Ǔ<�nn���M!#��<�1V@�j���oZ(5m�\�<�:�H����v�k��t�9���5��Å�J�x�/p׬Y��v�e�	�L�/����m�	GUe�oP�l���v0���}X����N�*�{=�Ț}W6�*�òz3=4�FMND�z5�a!�ߛ%y��m׺����#�
7�V�]�E��Ӣ�l�w/���oJk�����8i��p�O�Hv�|���5���� �k0K¬u���d����y���C�����?>.���$\�dUŊ5�=i@%jQ(�=\���h�YEs�(&�4x;��;õ�l�,��~0O �:��L/�C��Uӱ)hK�*����9x-h|t�+αiZ�i�z��ì�:"�nX/ԁ��ZV��&N��!u½��a3�c]ב�&�"Sy�O�\���C q㥼 <&u���sN�yQL7���w.F�X�E
P����kCN"P}��@kؤ����m-���^ܤ5xne���Fp�`�*E��}Cb/�!u��U��I����Tq���(;�h XU��o����K������U�U���:G��s�ǹ���e�K�<�i�h-2A+�)�mJ]��5��Y�q�S4�u��yʩsy����D���u��w<��Z�uU�8.?�"�9�%7[2V4��3�sD憖J��BO��N�@F�6�f���Ho'�*[ �s�e��%�j�S�I*��|��GѼ�vek����՘;L13����6`c!o�5NwBH*a���d�Y:�j*+�[����N� hXĄ�@�8��nj,2ȸL"�@	��*(wC[�*J u�y���WB����Cΐ�J9����x������1Z��Xm�6�&��rR%v�^[4�G��eN͖�X���V=i ��/d�-o�T|���y���ۘMO��u"LΧLF��ٌ�h���?����U����ִ������T�iT7�--�Y��Ά�d��ڤ�jY���"����9 ����zi�굽�F�|@������RU������,��i���n��BR����q����(��`�0�sC�L��2LO�W���11!~����n�j@�+f�s�z�t�XF��I���Vf��je,������h�p,&��1��,����"��."��&!�o�>������'�}Y,&X��rJ��Bd�I1�$[�,|�MuSrէɀn(6��>�jB*O�g<�/��r]�H���ʳr��u@�Qg��C���b�}q�eO�i����V������SaOx��YyU5�g���d
P:Ʒ��Ⱦ�cm!1�#�����Srg�w��F���<+R+R��D����1ڜ��c�>�1�4��6�3���uf-u��o
�֨2Qp�n6�:��fEYy{�����u����щϾQ�Pa��xhj:5����+��mj�*;G"&��2���!�Ɯƕ��Ճ���ӷ>Z�(�i�o�A�������U_��k�z�]H^�����u(�8���=Z;�:�<�L�B���&^h���!X���q!e�U������'�rÒ�SS�m��X b��|��&]��!;�<{ƌ�ܢ���Q^���r˃EZ$z,"��w� `�A2C.�AlO���I��\Q,row�i���y:*��,-��
Pj��E��d!���#����xJd���eH�r��)�-��d:'>���;����`��̠ U�V���mE�04k� �uT��4M�� w �f<��F�������d�9m�l�GkU��0���	d�z�5ǌ:��V�l�g"�C�(>�&Dm$7ٝ���?l?2;�a�b>���~�f�V�������%S�v,�@X�k7�D�b�cށsv�L��Hq������}0ts#��0��e��ӆ,��S�;G��֛K��y��ۻ�=�Ju(�V��2}��� �ǣ�(c~P���ޢR����@���ft���Y�F�Z}
R�$cP�|}�\]e���y��|'�����Q��JA���R,%����OU-��źā��*5�E���ɲ7����{ʁX�]A���\�l�C �e�He0��k�w�b� ��,-���,O$��i��V�¹���1���,<�i�o�-�����I�Fǡ'��Ⴠ�6���2��n�,&��kC3��B�0���6M�e7$ = Ǯ*�<�$ޫ�`S��J��IrD��ZXf�{ �ů��" 
ks��\xxH].U4h�^X��>�����r.¿[�����g�,��8���l�|�N6�/�ƚ��gSOX.���⫝̸�`R�J$�̡��A��Yͫ�*���k~Dm�㳼�VlG:+i��A��4est
�F都5���59���,E��]��Ȅ����r����H�E:9mPI�6�v4��cQK����%ܜ���+��Q{|�{�Uq��E�� p� �{��Q��i�Ө�R�SI�Ԗ��G�Z���w�mč�N �#u�]ds�h�"�W����,4惣en��9jiD0�`-݉&�����|���2v����Q���\��`�x��
m�z;�Iw_;�N�#�[��%����{'�9珬�c��l:r�Lb�¼2���5N�2��EB�����>Z�� ��w�x(=�\?���Jz\[�Vlg�b�TJ��E�4d��b�!��wH#�J�[׈&�f��p`�fFf�6��ڍ@�����w�{X;����XT���(�x��N~+:T���:��	�
Ny�^�%Vn>����1�$,N	,8�"�N��| �|�:Kj`2Yj%���t��F�"3z�U���ͱ��&",���8c�%M��{36�;�h�j�UW�#�s*Ni-& �0O6��-{��nQ�F[�w�P���e3��b� �R��-s}*��0��B
*�2�ޫq�&w�ש�`�;yW����jR)UPx�!8�AL��v0p�E�j.ގa6�z�G9�F�A����Ң��b�ܝ$R+u?M�'���x�"����I��e9�U����ֱ�O���_K���kv�M`z�����?-��r���í�uF�t�����wk�Ɣ�dY�J�c�1�yp�TZ�ًwP�P�fB+��U���H�{.葽W!b{���ƂMʱ�w*#��HA�,�ld�@*������ʤ���UIU��1.y�=�F(��Q>p�NX�8�gQ�ה��1�ai��A��0,�\xy�l�l�<�2��/U;P��S�}�R������<{�U>����C�@�պH�QG���K�o\�(�H�\�&�#�\��	X��V�V�͘E~kYO��>]�s��_7Y_����t,]s��z}	��kJ�5X�M-lm������]�\Ǒ�-3�zC@�C�/:z�����:3g$��譖\byann�7��M�R�U�D�ů�����#� ��rրٔ&!����X��hbrڕ�x���]I��+׽0������d|	�4��Wm�<!�S�?\������{�^RB_�t������;o�a�=� �葪Ur&��	,�x^Ҡ�]�!5j��9N ��=0;��X�l&&�Euj+��l��بxl�zVj&���U�~e� m$>������U�nt�mLz�RRY)�_<��i�<R�'�ў�M$6xRi1#j�}'v��ÿ��^��-\��������x�0�',�-�������xSN�Jm�Q�p.�#��������=�0��`-��xN%��L�4���)3��41`�#��&<��^1:�BoA��2����DI@$���\��o�-ś+�*F�`fm�x��r�"!$�,ym�z Ytb��y��y*�c���;��wh�����b�(z�{�Q�[�����D!:!`ͅ��^lY���bc=���M����9�'�R�\t��y�j�Õ�HfMb�x��m��b��u'p�KHoBi�~w��,�}$T�8������exXą[aO�L~R��ٿfy��w���O��#U�T-r�9
�ڨ�uR>��T���>�����W���Aԩ��?%�7J��YL,$x]�a���y�87�iEuR_"b\J���V6T$h��ԟb2��SP}��:�Z�Á�'��f_ �\�3$���d'��6X�O ����a�'��.~�s�C�.� �<I�e���(�['8'�='o��G�vq]$Z�q��X��K���s�)�a�x��&m��=�j�:��5��7"&��!k��{B��t��{�
&�ޫ��ދ�jb��{���tC����BnҮd��rΚzP�h!�J�\ͼ��.�"�T��cN�^�n�Y�v!�/�\)m�܀IV��]��WF�ɓ0��t&����z��א��K̸�H���*����6���/��͊9��yW-��eF��QB	��h@�$�WKD�u@���]j��������d���Ζ4��,AO~'#1K�t1\b�D��@윺���r]L�јY��ML��=k���v��m|�:��Q=?)#�����&iR��c����Z�۪�7�6!�F�$�'�q��(]'p�¤~�.J�D����hS��~»C���_����~?:u��*��2��COvDh5�3��Kv�6Yx�+ �g;Ο%C,��$��~j��.�qŠG{��J��>�����y��Cv�8�t�d��~�I�,
����&��^r��ѕ@CӜcm/ա��0LQG��W�ܸag�L�%U���*C�h��;��=Dm��؏�e��cV����3 �%	���G������G[O;{l�;��m�EO��}��?������0~V+�#�dE�ɾ�t�S�o[B��0�U�V�Q��Ѽγ�Q���/Rü&���%�����^[�#��8�B�J��:1�D�7�ʆ���A8��c�,�`@���_�YV����C��Nk�;��1&���8Ąѐ�V'�'Z��Ε!|��!�ѽ��j�:�9V6Z�ic<�lf��g��G��9B��k�q!����<�U��2�I�E�AY�,�GVڙcd���Y=2�ΠP��tj�QY����ƻL:O�I]H�:d��E>�:Db��)6�H�*��nL���������:���,Fe{�ƵQ(q_��Rm'���U���H���*����zD}����������E����YQ�'�"��jG����x�Ӕ8��m�c�7ŝ�KQ���&������~�-Ϻ��*'�18�$��H��LS�S�;3��\���ȳ�,����x}w׽���x���b:/�/>n}l"�F���'R��5�E.Ae��Q���H��֠ׄohE��u�i�$I���Ʊ��
�5/������v	�ur�L��9xE�A�F"-����Dw��z��V+ؾ:�e�,|
C���E�Z4�����{�F����P����P���!����N����1`tL0�Sy���0��|���o�GPӨ"��e���"x���h\���Ԑ\'�#øj1[�F�u�uV�t�Р��mdb{T�g��H|�����!u1��Zw��8�����9�oܠ��O���|y.��0�qD[~�.�(A�k�f�h1b�,'���1��Tm�/�,�G�j"5�SK�ļ�U�d LSUW�ռmw��H!K����pA���o�!ݹ\bx��W�P䗨�XU�e��,7a���&���vvj�'�bm4f�����V�����2��v�urm�GSvTм��6G�N�q��n.�n�֐>��
�R�v�4��Y'���������^8[x�E^!6�S��Ͱ0���駟�+�LY���8c1�qN hN-y�4�r.C�2�@6�B�y�&xE��q���E��e�^��7/�h�V��5hZ�;T�((�(��ׄj�ucb�T��^�{� ��w�f�U��86�Ň�p;4�r\zx�a�[}ڨ꫅�%�4����.�b	�՘���3o�Īʺe��?�C;zh\�9|������0O�!�&�^�:�K\�H�E�:�;*�g��ĴP�a���Yޭ���zx� R���k���g���&�-(A��=����p}4�3�{V#]\�� �?e�w;�#Rf0+�XյdR���klb<t���}`�	+�Z�jiyT�-��<�'�b�\I'�e�"�����q�[;�ｙ�8��6�/b��"�KB[ު����|~�������ܣ6��8�������5U�]�g�g�^ӧ�	j�L[�|�9E��"�؏A���*�!�a�H��h2H�0�lPw��&F���Bc4� �j����y�ڜ�l�u�
�'V�D6����5S,�̹��9���0B��%<��3���3C+lr�a�x�<y�F��Q^_�M���f���Ä�_��1c6���~Rub[ԙ��L�a����B8��4��Xlx�y�&���VB�c��/�BcX�z�Þ�[N��p�b�{�����5ʒ���O�����f�L��CHu������Kld}����`Ʌ	?7��S�a@���!&sp��Dխ~���eyȉk)~�y�N�7�������*�a�OJLL�ǆ�}vu�l>�Et~-H��X��&�CLQ�M��Vp�����t�f�?��T�O�s
��*���NC*�#�P�h�H�s��S����������Z������ap���>b�M�\!�ӷ�H��u��joTɚyJC��y�m�Y?9	b�^��3j�S�a�>XK\��� 
s1����y�p?ۂ2�$�F�ܱ��C��V9�p2�h�f�I�o�:��J�q�ZiL{`fɤ�ׅ'��C��'ǌN���X�0Qᢼ'z��H_X�Q,���v=�΃������!�8�%_��ҙ��^z)�Ѽ֫H�J)Q�(CȪ�=&�ư՚��Y��;5�"E1u!�&�
Go�l^&��Ki�F��%�/k(�d�#]X���)x���5T��Gj�ӔUnHƿ��ѣ�ѓ0�.�O�9�v!��e����l�؇Hs��a��?/CO��� ��v^=�q.�T�F��[�e�?�qM���z��7Zĺs'�q#n���k����3xR����kO��7�g70Z�鮒�sC��$/Űϕ�O��F{���SײTc�z2����=o;��\�p�)��[��o4,絥l6����8�ʂ-����}��8�pih��գ�ˌ�RJ$X G�j���s�%�w,-�q�C$ar�HE�=���|a"�O������YX넻�O�9������~�(�I/��bJ�����Mx�
���'mS_��̜�d-Q^�ۈ_���Nx�mRA�Fs�4Q�x�5��;O����q4�=ʚ+,�����G~8�87����$^�d��[�ko:^(i9�gQ��lrgU,��Pˁ���8JE���ǽ�R^�Fx[���%�Ue�Iq�j?@="̣��1���=ǌzu%�m>��>5������q��:��ļ̾�V�&\mQV��'S���e`cF/:����Դ9��.�zݠ�}
Q�������^�+cT�
�J|���M��еp���۳�N*eyh���9�4ȕ��o`���{��Pڈ���]��Dn�˵�!���y�۵�*���|�X��`"�������6�c�K�%z�%������J/�T�e��jG�T�fo�oebf����Xě�}r�S.��4Ҡ�i�{��`���jD�(;#Լ�0�x�]Jrp����� K甴m9o?��Y�"��/r��� �}9��'�"ђ1�Xm�˘�tƟ[�0��prN�ic�'����B{f�S��,ܹ*hpQ��0�����x�m�Y�	�0Y���[&k�x���81>Q�X��:�z)�s�)Ts�a3٩"�V���$�����;+�H>G�l^�������]�޽�L�P������LF��6"��C����sw�v��Z��9����>D|����Գ2d�bS�_TU�E���k�HPS���}j�*�ѕ�k��ũ@%
��FK��_{�_�R��}ꛊ�y��N�X?n�u�p�W���[c��%�WSM��j�	�+��{*�8f������������M�l�)	i4L:0V��l"�}���;��%W�n�k��G*�K�2(R����[΅-&v��b�]#��ő�u�Nh���g��_أ�K��1�s2��if=510��7�7���0/�Bc&X�k��܌~?GV~v�p
�Y�*O�)��
�8yr�lvC���������pb�y��z�B&��1�?��d��+V�*�F=���aT/��d{���+�4��F�޻��$=��% ;�D�i�O���0���]�=E[�@r>������bc-�d!D�W�K�|����PL�0���³��2��Gt��,�e�f~���A9.A�R��T��Y��־����Bw�����d[t�%�|�S����'F]F��/�׀��<��_��_~�8�|Mh_��ֿ���pÖ�8gG�}��6H<���bۺQڅ�&d�t�/!h��z&�zE��y�\�0d�0�kV#���Z�UY��q
�<2���pu�]��� ~�(Y�)NpyP���1/Z=��7|1�d�`���AӠ�Ӳ�&h�����.\��X������%怂�Ml��/��=R�9��L���ǸisTa���<�#-1���L,�`St�s�:l7�fP�hs5q������ߚdX�g�&)�M�����YZe����9[�DG�06<R$�f:;�Ƴ_�{aD��ߕ��T����z���}�v'~� ��1]���.l�r8̞@e���˙sH�U�p^�����T�'�Z<I�CX��mo˾c4���I=�[�杩J�uh�$��r���e�>�����������:��(�^J��x����M��.x�ʵ0B��1����:y`c��C�Y,�<c`-[X��d�)WCeH����:����6��������;''���%���I[��j�[W�Q��H��pJ*��=�ND��#eѦ�f49/�5�N�W( �?+k��P���P\����a��kum�PD|O�[{
�_��k��6:=�ţ��Z�p?b JH�dp~�j��hԉS��W�ę*G���q�T�S~)k��*���:��Z7A�(��
�6��e5��<+�x,?���Ex?�
�CC�F���Z{
�b��9`,��e�rث�	��D��v��6�$11�W/<6�5��4m�[�;e�hC�kQ	�A��XlC���.�Ö�L@����[�Q�SJƉ#Ne�^�Y�M�<BnV0����84:7ICD��r�K���Q�w"�O�}gc��������kXM%�`�,J�]e�u�@u�S���:e%˟	�Q��*,�1}��!����+����/�#*l��]�a$n�/T���M��Kq��:I;ym��
g��~��*R�������R�nW�\I<T����KPEwo��j�l���8�*4@>�T�W�YaPA�j|Iaq=V�k��mʀ^���`[�����-��K⻗�14bVTU?*]f)�,E���6T��;I�0Z��t�2,��^ᘕOa-�gpu�u�!J=���Q�n-���$zA���M�88������a�⌆���+z�4�T����}0J�"q)5v{=�*��UҒf�<��j�tt�V�����`.����ګ5��A]�00��k<rB%�@5G�9Z�!;��0N�)[�d+�*��]� �<�M1���~���%��v٦?-�;-�r��.7�j-R9�%��*��-O�j��{��S�U0�L�u>�>.��(#'{v8�wz�e�
�����Z"��7����?-Uh�lߢW]�ʰ��d�l��ڽ�`Cr��g��c�A�Q�3�rq�_x��U�[c1Z��Y��#0"$cA`�C���33YmjiR
������j4�]�Fx��%�1��*oSkc�5��A�Fqlhp�T��*T}Q#<�����D]�r@��/����gB���96��%�C�ɴ)��>UX4�x?�i�i�
������>60<旸D;J�(6����֒{�М}��r�4(��}Q���Xm+�E�+ͽs��v���#}��Ƙ �?pAq������=�����	ii����9ۄp��ke��������eV�^�%�.��M��U���H2�{O�8�{��y{3�{W�W�fZ=��&	a�X7�Y�7�P�n����>��bÇ����QӁ���y�8F�d]�e�����̚��&��B7�5�HQ��1"`�V.c�D�̐���j���7:�u_yֈ~֨^�Hݻ�|�j�3�����RtJ)#:5�{p��y��zK�d�4��I�ZxOYD�J�����㧨�)nr
r��z��Q�1�)��B;�ir��l1� OmH8���:K�H������/u͉<����ph��X�ա��&�ar~.7:\��p�?������Q�X9D��ũVY�<>� b�Ȉ*�=�w�!S�wG/FJU� �k�D��>�
WG������6��Cn�ݱ�27�˲���W��D�V��VO��]�
�����_\���»#EG-�����߱���U`���a=�橞� /��C��������f��x�/�cOZ2��E-�Y !j��^J����)BK��@���q��^�!3�P��0��#ᲄ�t���b�R֤����,�ōxmrF����6��/<�3���S�{�~��6�[��Ux�8�
Ee�m0��3�>x�ų��B&��8��3����ԃ�%Ԝ��I�,�d>�O�t�F�:,F�:a������6��C5R�i����^V�Vɬ#~iz��þ$���-���` ���w����m�|M[8.��{��"|w�D��gñ����sh%�V���x�B���$�y�Z�����vUE�,��0H�����B,�ˬ:�O�����7ՠp�(��^��ƌF(�Yv�;�w}x���g�6'����Z�ŷy����y�z�р<d��5�Nj'��ҳ7�c��e�C��iC�Ϥ��ͫ�:��J��r�V:�Jzw��<*/����n��c��x���H����1�J�l����tfƙ��1hs��	,(�jE4��hE����`�h0��<U�9C�֡�5����t�w<�Ns���G+���y�N��}�2稒S��%#��=��ĺ&�ٔ'���J%_�^�!;'6J^(��";C}�|q*��{��$[+3�S��V��ճlLXM}�֥:��{�Y�^>�p���S�� �]'�?Pڷ߻G�ifu�ɐNSbZ0�M)a|EybR��>T���:q�֬/(%��3�3`�O��K��R�p��c� �E9-�=(W�Q5�_<�H.�O�1�>gӄ�؄��җ��E	���,�x,j��ɵc����xn�_���X��U�$EBT��A��ۅ3��Fc�n�%�|9����#'z��z��r�Y�E�(*H9$r�j��=E|��zP5^P`&7�y��1���|IE`*�g�p�Q����.���q�m�#��;.�lXJ����S8?������'��`�L`�+�v������k��,��z�P�������y�L0�p�0{���]�qza������Տ��s�#AW��ɓ�r��;�/�oSk��j�57�H����u���[{�/���*��S}��(oD�H�p�L�.�)�2R�U]�^)OzQ�`\���1�}X����0Jd�atL�h�3l���8��:a��AM�v�O�-!�o[�M,�z>G�[�]YS1x��G��,�EC&O����՚��yj���Q��������}�]p���?y������e�F�޺��Φ߸G
�"y1T������C������&f5:\��ۇol|��po�V=t��g]�e�;X�Zb�� %BzU�-�mR#ֻ��c��a����s�,{����E|�x�Gw�l��
/�/���;CW�؄=q����"��q&��H�5;�dG����#�I���j�8�G\�WD'�u���?�P���d�0�'���oT3;3Q����א�X��OB���X���N]\ Ƌ"��L��P!�cL���	j� �A�Ę;#������6�B�sX��P���S��3<��jc��&���g��T���V� �7�1�1��H�H�`�Obn?:q�?�.�H�2��i8�%2��9y^�gF���~c��/��4��u3��׿n09e��]Q�(����L��E�ߌ����1�R�Z�٩��Y�K�y󚟻,��d��{S)}̼��;�� ��
)�E���0��66.�;]���f�����I┲��n���N���&p��Ơ�K�����f��.�e��'_�A�!��5D;����D�a%'����om�gf������A�xyk��P46/��Ͽ�l��9P!ø�7j��3���b�/�P�3��2����Ӓ�[�����+���5K��mq�s`�[MV&�|ѐ���1N/�B��14Ou��D�Ԟ�~ �����e���i��{��A�R"eT*w��1����5�H���W�Q&�?�:	ѐ����=�X"�Q#��`��yd�b'n�T�5��}��U����iHk״�~.i@􅢌�d`y+FQYo�9֛���+����y�0�*0L�ѹ_'ǽ��)S�d��~g!��:��	�{\<��wʴ	��N�]x)�`���Y�ƅN/����Z=��!�r����|�M�!u� �|�#C��M�<8����^�mX�z������NbO�ؽ;^���D��0�6
�aE����7yph����L�5Ż'.��\S���Z�'�2[��uS��s�Mc~�1w�2.�yIKIm�Kx]0*=Og?���VS�������o����1[H�m3s���b�EG��Ѡ
�s^���~˒ԤNe����I:7q�>C�:)����m��TX֏�N�6��~�a�Qm���jG&*�J�����Oj2�K˽�0ܼ�6��*�&���aZ����E{g&��(;U�-jYmO����NU#̰�Ru�����dlaGa����>^{��aP?��r�6/zƘ�@�y��<������Q�Ð�y��<e�=��M��dOr7�Íp�^4�������-$�͒�m<�� =�ʾ�ln�ML�r���Dm,F����Y��DLa5:�g����d��8��_ܠ
8�D�zS�t��Qy���K��>�/����/-���A
u��x�*N'1�l!�0���˛�c��S	C*�S�k��r���G�F��{��&Bz���/lC��bob���`�7��W|���e-_<Ǎ��(B�D��=�9O��D��z����LTc�{�R�r����������P�b��8���+�g\ǎB-��z����d	A�S�����Y	��5�'�Kx�C��a\$Wi	��D��8l�	����ޫ���%�UF*lB���䀩v��w{�|�z�3��;�O�@���5��й�s1g�̉#t|�`�`���zmH�K,���Jks�o�?��\�>�����T�L��40���(1�4xt�w��7<Oa���PWHe��wVJ�״�f
5��ryW�V0��!	0I��8՛��a6#�J1�p��Yܣ�! �hL2!z�E-:�@/Nc-�,#
���/�����3��N��U�m.��i�J`��	�:8��)���r�6��2�T<,S��^6�'�p������Fx�֮'����[1,�tB����:sC��%�����O*X*wduZ�^��Eo,S�9[���j4�m��6_Cd�J$���dD��_b�K�F�7�zC��!f�I���Ŝ$���� :DjfHu����U)yA@��1��jh/���)T��Ս,�܀ޯy�M���/�ϥ(pɾ�:u� JoT"�5Kf��+Ѧ����dᎈ���ɚ��SZ����T��Q�f�?/Z��PJXy<�0�� kM)\\Q�X�}��//��7N"d�1p Q�alY�o�c���/y�O/�5���tTJ7��{��Q�(b��7o��]���׾�'�F)԰��[g���P��d0��E��ް�H�'o�P���=�.3�u8ӵ��K'�*8p�cп����\~����l[<���1�2�C��%�Wj[]bC	�z������.��F�jh9�%� jR��
Π����R���5�𭋵�܃qҚ��E�J ��ߥ80i:���ƒ��|��Y&z)j�Rx�f<'�2.F��F/�<[�Cu�(�`�G�!3�<fe�go)]T��3��D�����3�e:��5<P��@���ָ3)��̣��sd�	���	�'(���I�D�A�����6��)�f�XUvtƲ%3�W��%
�֖��̳�5�I����z�Z����*�+��C��Y�����fϦ�xj-2G�����S���B�O�f�0P���.�;$JI�a�ؕh-BvIؖ��VC>���ۄ!������ :���0�2HN,P�#�G�\��FDF<�h{3��������`��B@?��`���kEbc�l7�}l�;)��6�wVf�ɾ����Ӑ*a�'��Gw�*�@�^)y�X!�kA8uK�,s�~O���&)[�;\J�nӒWUAF _���xYhPsF��/7Zk4>��9����tP�RO�����l����p������$�C�J�l.�*�����hU��Kx�T@�v1CJ�sDe�"od�UAm|�_�ͣ�c���E�5˦�iɲl#�7,��A�[0`4_���^�5���Mi���%��1���&�7�zEk���65;�V�1<oi����u�7��o߆��9�&�O!,W	�����P�5&G7����J:��e�S�T��@�kr-G�5Q���/�G�Q`Ѐ���?�:�ym����
X�FG�E�8R���k�*6)�h�&I4�F�*>���]#�������ų�<�aP���%���9�_�Y���7�|c}h`�@���{����}�"l�A�+1��hkR�j�ӝe�]�Lџ��c`�)'���J��ᆆ前P���e�}����K)W�_��T�\KI�)d y�ڈRG#1}�e��ݣahmۅB��f��.>���#{s�����A�sw��8Gr���P @�#=�w�ޗ?���������?���s]߳-ek��&�]�+��1b7H�b��g��MGB^gaD`olŐ�n0\ޓ�>/kؕ����������?�S�{��ŗ/)b�8��Ƹ�B?c^�="�RL��YNV"�_�P�9��b��W<VL��J%�H@�~��N%��~vo���(cu	y�y�S۷]�M��(_a�� tʕ�D�V�N� Y��U�H�N�!�Iv���6��r["��.����9���M[lEb�xRJ�/߮���o����?������u���6�0E�-u��x�����iؗ��>��("�k�.(�J2�7�2y����� �p�6 :�F��߯�~5o�.²G� ���}K���(���7r.6�j6� �dR�~뉦R�� aК#���~�UUh?{��Z�섑;)��(��FΦСA��j��3%%�:�q��� �,����Be�;�ڎ��5�Ю�39�X������eRy&6�;+ay�����簔�G�i"�/<�r��[�FKf��e��^���Z^,�?3���Ǯj�����}�{z�g=gh�����Si��R�rb���ـ���j������S����H Ó'���8��kJ��b��Q�D�+�a�4��Y��2���7�����u2!<M�8y��2����n�y��N�!$����0xƭ�
"U+)���J�������H`�~��5����yx����0����iT�D��\��t���R��nz�j�a��Rj�dl��F%V[�%1J�1VݾȖ��K���V@Y l���ٌ ��yA��b�fl��������h�0
|]N�J��z��V�vC*o*�E����2ň��%�tx�T�O�{4�k���L�JZ�QZhT�C�LQi�eF���fE$V	�Ⴭ�c�h��!�AN���\3�A��;��&�����>���*�i��WUr����?k^�v:?�8?ɲY� �#�!�?�o,d[H-�,V�h���!
\$q�̮�0:���x����TگD�œ��H8H���L8�ơ�O��9Ws�ugbV���`��^n-DEp$�NbR���Ya��PQk��9)Ǟ��jD��s�4��Z�n4�ީ7f8���(eE�����T$)�ͦ�jUR�#E(���?��_=Q(-���������,�����}�wkx�/�`�#=>E6�d��s1zzФ���\���MV�'��Ï�P��P�0%���~�nQ)��5ԻI�ʊG
u���+�Wo	��ݻ��~���l�Ta�a=��E��>����%S���?�`�����qoOV���^�z��������qfV{x4B�4����59-�T���Qk��jۧ(��|燽�w^���Q�0�a���(���0LTfS��d�1�f�5�Jl6���GG������k���m)�Ah\���6��*� �e�&|�a��䆅	\�W�ְE /��[;` {<Z��2��#(&��p�����B�{O�R���j�R�V`SE��#��R]��s#��7J.q�g�-t���_Z_����\C1�ʔʉ$������դk���p�5
?B�Ԩ/~
�	Q+5e�M���d���G��'2=)�&�:Ϥ9Y�k2Au�S�#0RfY�8���EU*��N�_���=9��0ޓ���C��K��̋���k��~�K�ʹ^QHt�T���{��|�l�� �����_*{'���E�1�K���axjH��"�Uޕ7j�U<�\S^�M�<y���
�a���"��}�O;�f�>�F����&�g#1g�c��J6��V���s�����n=��.m��d����4O�����]P���\w���g���5��5�}��C�\��Uh�^_�0^m`�dWIM�	"��$g��8�P�.���j�*�?y�T��.U>z}P�E��C\Պ�*57�xԼ�j�?���=���ڗ�o���l����A2�B�D:�^�^��/��g�:#�Ā����xo'%]TՄ�`f�\�p�����������]+����/�j�'�P�����K;��;;�%�E)U��G-���<Qy���\���q��	���sZ���A��o�?&�両QoVO��z/��"�i��RR�,i��8cIƐr�=HW<��M����s��P��<|�ȲN[�^���Q��!%�4j��9�i8F�s���XY��T��yD*���Qk��.��6�p^8pj}��k�ki=����Wo�h��2g�����AE�d�F�����N�U��gS6�-��ڐ2A+1�M}l��}��x8O��ٵc���զ>C%��(�9��C9���w�/25_�����p]уڱ�\bǃ�������>���d��̀b.�$cy^f/�X,����H�6�X�j�[�(� HFi�E��$m�4��3� ��?�33�F!ZԿ�ۿ%Bэj��$u�1���CM�T�d�j���o��mA,F�Q�r��tل�x���=z�iЃpo��l�:f>�Gy�u��W������g�y�ӺDH�<�4�U�Q�~�`Y6��>�+m]�k�l�k����56�u�F�F5�l���/S��M[ym2��dK���-R�ғOYH��z,�%n<���f˵���t���t�.4���,{�Ui˒P� ,���lE���C*	J��{��9�S&3�����M�Ç(��UF
xH�{a��Qs�J�,����ֺ���b��!O��f�ȸ*/�WF�$�g�����J�~Y�W��N�Pxs�^Ix/�p�҈j��̬� X��ݦs�H���htSyGm\A䕔&d|���?��&����Y>��C�����aSm5�'���]P���8�<0��γ�N��VZ�X-
�A.�k'�D��EZ6����������~�۸x_��-�1%W������$�zԡ����*�qK��[��!e��5���}��os���x�����o?��%����ŀM���_E��8��#�����*R3g��:3�]x�˒xp۶��ԃ,�8�5���I���7r5[�V�Ϫ�g~~)��z.��,��b0j����1A�	b�0���Gz�p���̵���wV��"T�*Au\��1pYǉ9E��"�ݶE��������z�=W�@�W���,_�T��yђ�y:g�T_21YfT���>�u�\u��m�`�cc�<�&<�*6�����a��g�ЛT�q�FM.�D�6��jp��;MJ���,�|Ө�����Iy��CS�g
U{y���w�)�A���u��A&��[;`LL���,��t��d�Tߓ�|�����qRx�&E*�N�0�Vds��"[�TRx����ʛ��Sj�k��-*�u),y���CYV8��{��c�	L6���k|���$�4��ήC�9��9�/�Wɪ�4������o���{e�����@[uq�-�EU3o[B)����|�ј
�m=�a�)��m�EV�Qk�<�}��O� �"�X�%�_��ˎ��ͳn$���^g�/�<@Uuw�������[F���6�+%7ږ��(Ө���S�K���^v�5��.�w���H��b�mS���]��5���%�QTs3��m���R=uTR�i��~�'b�D�ׁe�Y����L��)ڡ�ЬJ��RR�Ι��	������>�^�ad��O��t����g�=�0}&�K����k��u����~��(�w,EU4Ž�4���W ��{;������8����ѡSP|�m<¦$�n�6�������<�K�\zf�Ϭ��޳�uN����w��Ѳ5O5���e��f܅���>������y~�uO��_�N������9X�񴰼0���>z���S�]�s!o�`�Bk���)Zc�'x�ƍ�:�')\ͳd	�ͻ,��(I<���H��d<�ǭ��Ә�f�I.Y��
�dD��J�Y���=f/g�KN�|�g! y��n쬍��Ƚ@���\�����w�?2\i[�|zAQ��9Y��}uF56Pf��l���2�c�q�QRK�{_��x�0� ݁/�0���]���S{�I z��f����.<��m��jj��։��k!Λo�N����1�gAx�΀㺻�ǣG�hj̵���C*��@;�ܠ�%{�,�i� �\g��?�5U/�,��#����:�������mq�/����G�),�ijH`)��[��g$� ����_��z��D����F0���H����a�f�=�a-A5Ed�	�����9��;Ab  ��m۠�,�N�`jT�D%���:���e���,ڲ3�`�/���<�hH3�F���:ǿ*!�(�to���GUx��n�`:�2���9�:��&h�����춢�z���X���� [タɾ��(5����zM/��g��
���}P�z�Kl�����T�I� �yb���l2�]��|���A�������3)��~�'r�՜��E��$z(�l
1���t0j�rS֛�ґ��/���:��Eh�R�G�Yz�2_�D&�\�;CƮP紤q�P���fk�6������^��ɇ߿d�4�ߗk���<��Ry>���"$�?��5�N|鿯�v�Yt���p�嫗���K+��]3U*O׏��bSֹ�&�!Q�GIFZ�d����^G��=f���������ޟ{�v��_P�߽��b��9]�`H7Ft{�ͧ0^��*L�s�����۶�I�>��$�������(�p�!��=�H����	�6�U�q!lD����F�Q���L�.?=�-7^rz�^T.e�I��=�.�B�]�=ʠ��5��C#v=��ڄ<��9�U]cnO�jK$~�����o�_����B��}�*�a�ݨ0#��J67�y�!�Ӌ6�|�e�.C�.<��������@�Y�˦�\T���)a)\�2����S�Mc]o��M=I�J�\��2����#D`|�47}����9w{MX�8Ȼ���}{����Du\[�y�y�m��*�2�����^)u)%�w�ړ�[Qa}��t����ڎ׼�� ¯2�q-	i9(PJe@����'�!~
o�E��Y���z �j9�f�S\�=��%&���K�Y]�/2�$a�	̒_�.�
�����x�'~��m*9��`#-�ё& ��������߿3E&^w�JTzbݰ�ML�w] �g
Pj��!=k����g��2�z�ԙ��)h��&4ɍ zN�Tj2܆�	%w�\�mUR�
��p۹h0�ὥ�w�+��Z�� �r!<2QrQ�jC��p���~& �q��Zy,v�F��:k��?�j�����=�K�qO��~�Y����_#=Ϭ�W?��1��-���`�>~�3#zO1���\�2�� �:
��Ȉ�5l���Si�d�+W��M�>S&:�����ob/TPP��_��'�imD�ƴn�7�����T��8��������s������Z��[aR���t�q�φ�zj�I��ٓ\M���N�n����D�n � #�k�ɸ۳-Bk��l��Ҥ� �#�Ab�a5}��m�+�	]��Cx���l;��7p�~�����ӵ0�ކuMɹ^�k�����t�`�4��L�Z?��1vk�:�~kH���L�xf?�N���\�7���6"��+�� N n������E��5v��f����x�:@I�����EFpI�6wy)|ގ��}�w��j��g~΋�����>�Mua�{�YdH�#�������nE����o�9�l�h9���>DThw�c[U׉J��Մ�EFC�)���,ah��{��e���)�k��\Gj[�?{�~��p���B\[,�ox���Ǉ1��u��K��6�_?�ݶ�Z�6{
�Xb�0���tlX��i�:/^�0$�@�Os�>"�C��%�-���j7�Z��T	��E�D*S���\@&2`���3��|P	��q��h1!�	�R�=I��8��߀�d���2�{�H��⎈�ެ��2C��� �º�
�\d^���Xn����|�Q���ŸBHd_I��k�k.�x�}ˌ��-�h���U��x���G����^*���;/N��2O�g�9+���𪖆j[c�Qᥳ����S�j�#61J�?4��9|�Cl�S���	��'��z5��k�������Qׁ�뷭����gHf�����rx~���xi3�$lR<�F�	>�yB�2�ʢ.�@l#"���ʺ遂��2�Q]Ԕ�<R��7����c��S҉����S�uR{�)x��QJ�I5_l�/A`�n�y��E�j��k#k�ƴUx�8(�~����N�L:y�3/�!��.=�E���}����32/�g�Hޝ�m�Z�2�rc\)���ы����~�'Զ�%�6�Ѯ���g7��;��( �0�x`C����5�ľw���b�Ra���4�d� #����YE2���i�s���6�k������ݳg���>�_�w^���C��u, &b]>n������hS�ή���h*e��	*���	��A�`[7*+���}�����zzn�9�'eT�u������Fg�C��K0$U��<N�����	֙r��k�^�r"� �����k"���;���~�zޗ�h$�����q�ޤ�6�x��iv��h�v�����~�}�5K�� ��7	��d�it�j�ثطx�u�=��U�e����i/��B��8k5���G�7�F��6�^����$�\#Ֆ�fX���6ɤU𛡽Nؔ|�z�����#@@��:���i��n#Y�~��O�`�Ïߗ��?��cB h|>�?=�0�0�777�q�GIVGI��B	
��x�*6��z}=d�.���!<ٛ�ߕ��D�}����DS|aY���;���w��tvR�1c8�3�q׽�F�r�EN����g'{/�+�wN�i�r#5˲��Ն^}U��BC�WLM��+�~�N5�P��E���f���v�ۭ��t@����h��H�n��F!���Cքc�]F���)ڜ%0��~Jc�ؽ�6S&�����WC��+�����rv�����6�밐�)3�M��w�N�X2
�yh�E��Ӿ�0\ڲw�'(��8����E��0��=`�T꬧<�ө����7߼1�{�N����l��,�����!�B��MW����RaǙ�O�[g��,��6�+O���3K��L2��P�o�H�V��F�q/�*>�>�¥/"쒘N�Ŋk�*W��	���I!6����%���)<4�C������k$�,���w�J<����ь�鴷�%������wc�����	���-���,� _6��ڍ��ڪq���R8�a�=-�z0İ1����G���D�B�V^��p���]���g[ǯ�R[�p�u�|����ՑD��a��x���i�kFG���B���WzU��[ٸ��D��]�n\V<��{	��Rm���lLl�)�#2���Zu�K��������*: �Ǭ[pϋx�҇`��<x���Ѫ�umŪ1�X�GI���C[m�-F�Y����~����Z����UKl���`�K����_~|ޘn&��7��!u<G�I�|<F�H��j�n�%q��i�S��R������l�א�F������x:F�a.ZH)B{�,������o*+�0Xʶ��=I�<O��?V�&�������������?0��TyHV�HKF�s��?���~.�%��.��nO~˘
.�gD��.{�[c�}6��˦����w��:��Z?�-{��3���x_0��0��#x��޿3�K��`늻���e�N	<h
�
|w���q����Z�N��]NB�fztE����|��&��S�M�T3���'��CH*�#��&�0�L���S��ĺ�G�L+ `����0J�:H'�5��gc�Y������_�m��K"�l�s��5�z��%�V|��wM��+���襂5.O��ZR2���QkV����M?�?kH9���	�|p$��K�g�9Jʨ߄���'M�ݝ��AkI�!��в��JZ�!&��W<D�<����vv-0��;�J۾�a����j_\T�Uow<�$~�����(
����W�\4�OL@�z�"-Vi�I�eIuv���|ҧ�����i�~iq��m�s5�j�=VM4P�Ҿ�\��Q�YT��g:�yȃ!o�k���
�y��[�&���a��㽵��|i�#�v�@$��ʏ�+C��_�>M���?���[����D��S�Ph��q�}4��L��H�@������]�h��j��k�T��x�&��F��
��+���+�z[�D�ΨOԣ���{B,�E�S��B�m)5�=�{�/>����C���({&<���
z �%�ǣ֊s���|���_V6[h/l�	��8+��W2@ p�(iX�q�e�I��{�+7�G"<g|���ntU�{�����+xv��xdHS�x��Ű�X�a��P`�]E�z��N%�b��ՅNA������WqA�'�p-<Ykr���^m�8��]�x{2�2���x~��8���<�*i�;@�K���,%��k��¹Y��ģ$��;�T!��W��dּ�bg���v�l?��'"���}��	����%�ty���9F���.�5%� �O��&	VOz�F�J���N}mbB��r���*�n��F�i>5���)���&�(3*m�'Ƒ��K�\�S���QF~ㄵ}�����]�ѽ<Gӈ-�l�v>^����{{/��T�@�G��F��!I�hB�a�N-u�4�M~������m��<cH=y�y��� �	�,�a�I	'�H)�
��Y����8����;��kh�ɺi�$߄A���\8$q0��}��ou��?�P��O��X�� ���io*�mk�,��{[/��\�>�ԑ)0���:a���`-�����j+l!���1����}W�X���&��Z�z�2<�R-C%k�R�o9�©r��$�ԙ�O�1r!�uk:�/�c����j��Q9����?~��ĸ���>��C'1h���F7�C�eI|L��T���G�?��PQ�a���2p#ƥu�c�E;��jc��gi�+FI����u��$��1 �|�ڛ]�6/Fܻ�2ECΗ10~�(
�`��T�}�(��ꥺ��TSI�q?b-�ɅF\
��~q�e$��E�^K�	B�q�U�ᯚwQ0q!]���1�k����J��`z�7m�F�f��a�˕u���My!ie���n�H�m��.:�H$h����X \��.G���;V������)������B�}q@wMلL��5ǯ>酵 ��$�����'�FM����B��<�9}a	2�ܻr�2����@�� .��
W1�tro]���[���G�~פ��&y���!�q �]^q����b�}dI�6�,/`pzp�* B���|c����r:3��}�m��~}o�u7}4^�%��6��L#&���u����:ϴ�fJl���z�,��&�h�\�o2ۙ�e��6<�h��Oc�H�!a���!���ܰE��U�u��a�1��3�����@d5�d�ԇ��j�N���s���!��Q��	`�F?K)�{�&�_ّxY��@���Z�3�g��9��M�}��k���'��5���-�4��R�B�q��'��B����]}3�v����������=/^�*/_�`�����1�>��74hP�G��1Kltz�7~Z�{�!ԅ���t{�4��u���<'�5AL�K}�C�����fg���:{��PxX�'�pqC�!�H��Ґ>�w@9�o��,סni3X����.T�|�,(�IpN�0����c��zT�xU��m.H��~[4�CT��e��}���2K��a5պ�,!��,Y-���2ySA+�`��r9/�SX�y�U'�,O��?�����W�S�8&8[Sf�ü,�T��vC�gC�I���������z�1up��%>\���͕�vN�e��$�ޯI�y�돲���6�����|��Fa��7��L%�]�Ԙ�oݙ���ƞ	�&�W�.	�W���M�t&J}���7����po���2ʵQc�_��~�j�ƴ�W�2zҜl�Z��`c!Iȷ����s�kC<1�h��vOH�y���0t�G�νRS�V޽s`�@�Tk���<;�35����Ƶ�c�7��)\H�^�8��"�q��Ę��{��.��Zg[8U����Y]��U��_�����5[�:�b�V���A����ǹX�e9;�6�W^D��6�H8�-.��FK{x��0��a$^y��Ǹ��ޕ�>ءz�y\P����#��u�{e�^ǈ�θa�,�Y6�	��>j���a���l�jm��so
f482���:�I���$y�6V�'�sa ���]���y�FW�?[��S=���\�����������~oUf�G6[�Z.ꟄϬ�~���!�����Yu*�h��r�oy�dc��0�{�tB��+ê��-Z�p�+���4�_멖���:=RW㩫D��M���X��`����#4���)$W��fg���^E��
�6��=����ً7Jv8=+r�D�T�,��K*�*Aөj����~��u���wi��B�~ 	��z�[�[`���^�@��t O����e3�u��TF/cMf��:����V�$=�9�>S�A��i�ݷ���ܳjj���I�ѓ���6�I�hK���Ƅ!
4^�^�[&Z0v0� m�����u^'㪹����Q�`�p@�L %������nn�M��:U #�C�,���]Q��Mv��23�J��[#����Z��ֿw����K���*�bQ����2�|��}�*��}�=C�y}ݯ�k���,듪f��}/�={2���@�������o�i�uE��� @�r1|;�߬wG�g���qaT��V���N��+�q�S=�9�s��[ҵ׏�6�%�|储�+�N�m����8�V�<K�uR�)�l��m�8_�3#ƞL�s��wx[^�zm'�4e���Ι�e=��Lw�]��`Sb1՜��0ػ04š_�"�b9��2�SQ����ߛ�ђ�xK����g��K�W�(�Kũ&CW��6k�b��mxV�ѸAgJ��O�ir�����_�x� �S�|�� }��˅�	�`'��N�^)�C�t�L�������׿��OѺT
�Z�#��SF�nm�1�%յhL�͉`�zt�|	�-i�E5��s2"���}���~�N$���cv�JcOyE�ED���?���$�l���8�^�p��d��`�`�T��'���?��V�v��d<�������h�[Mp�I[�}펵!����*#;,���D�"�T����'M����u!2�6���4��E��{�Gy�����I�))P�;���>�x�ڄ�)}�))aצ*/sw�0�y�3d���m��3�h��@9�t*�|�@�/k���@,(7�~_a��H�:ƺ��B��'6��ݧ�l��dz+�"��gI[��ڂ^����7N��y��c��4������B6����M]����ˁUsF���v��Ѥ�=C�ٰ0�
W����8 ��9����Eb�a54�}����s�XcqN�:�,����a�	��:�2�0����Z;77�9[�+��?E�z�P�\�
�K�5h��OV?Ǧ�]z�W!}R�+���8
1�l�������6����_�Ay1���(���+
��I9M�Q���A ���������oj<��{��lq�H)[�}�x��{ͥ���Mh߇��p��@��ZKM�Ab��a[��(�"��$F�p��nq�Z{1)�������h-��!�㞛�~v-�_�ק%W�J�C����;p#����#�(k�;�7�yYͱ�ǀPw�BU��L?Oo�m��,|}�<9Ί �"2�g_\�#P#��'�t�dEދ��p�R��0�d�����V����3���Ɍ��j���:T:vˤ�h$N�hۨ+��C�g�s�0�ҧd��Us�s����i��c�j�W��T �zx�{�j��:��0/J]xh�V���`7X��v5��*r�=���=l��bks�.�������A�c�غ�P+�1����4���C'�O<���=���1�Z�'7WS%�,ٺ�"V+lD��&�l|o���b����ԅ�I��*cx5��fj9Ep]��;:�eb�S}yK���V��۷���z�1AH-��~^���z�l߮��#Z#?�x�0H���ץH�s99�S�v�(>^�mj�<�q9��Me)_�EI��?%
��	)z��;�'��Vwb��	���t&֔�S_ͯU��k����C�iT��{����)����򾖪�o`��bX�E�zz뺤;ǌ�8T����S�0�%��B��4~){�6��H�Ń�?%�|�1JO��(�［��fkƗ^�����=��~����N!I&H ��x�U���f������O�Y�tJӃ��_*�<����� m4�D�ǟ�:5��/)K�z��n�o��'�� 6Bx�Lj�������2���6�r|�<�u������U^"���Bo����'�莆��*�0�5�Æ|L�bd	e&mz����y*iHc��4��sat�s�3���E�-;�*��k��5���,8�h��;����d�_�_�P��~���{��|�͛��Ո~�z�߽�f5�k�#���%/W���yU���1���桰c��p�d�^S,�X�i�*�{�ƣ/^
WjM
;��KTN��qq'�Y((>����g;���*�{XXC[�u���J-���%^�CB���*n`c�-�L%�����
����z�P�!�<R�-�sÈ���z��S����#H=��V����灯�m�|;�V�h��M}S<�&Xݙ��nnrI���.**��~�:C}�ϫ���?����𾝱h���?���'I��t�pn���Z�5V%�;�R�a9��l�c2���?�d	e~��/�xv��0/�~4�=P����9ߠ�$	_�
YB�<q;L��U��7��}[~��7�>-a����00'�7)�ū7���+3��6�/����7���
�M��[5�"g슀�*(ı�%<@?(п�]�m��F����Ê�W	�[�4[�`�Gn��#�󪽊M�TpM��<������O׻XvQ�𙱽m�@��Y�h��s���0�	��)�-��3��u��}�!�HN������fh��#��l��(~�rs����Eg�KTm��@��cS�7�}0��50o�#��x!eP	a�5Zb!~\k{�A�܉���3���gN��ԸmdG7Q_�
#o�ﯢ?����X� (|�#9qϬ2a����k�F���+�)(B7�����Ƀ�I>M�eS�l5�2C5$�(U��g��0�%�)x?BU,�l��/A	qҌ/
|o5�	���dg;��{�<���pn��@��9DeW�eo��ɓg�xhL�B�j&�R������4U�F��һ�߫��ՈvٗI"��>�@���b�v��u�+�<ކ-�1F�e0��}�6!�[��s�r�BfPD�Е�p������٫�nn_���!Ex�Ǳ�Ͱ,�}�ߌgeH7-�}-�&w�큃�do\<<���0��1�B�n�ub�/kh8S�z�0=�^�ڽe���n�a?Z�`<�Z�4o'&
�Sk��!����؂�lk��:�UvzNU��z`s�f�0����.��uYzz�翷�-*����!�m&�I��tj:�`�-�j
u7�g����U:�	iU��3��~E�]G��]=��־�
�TZQH_y�T�P,捌���U?�.��
��gi��t�T�MlmHEC"	�&&���N{���D�=Vs�C��Y_���v�ʫ����Pv�d���XI�z1���`q�z�g�Oمp�ทԨ>�~<�:l�:��'�F����ͬ�uM�ai\�d�S)�Dq�)8�x�`�z��<yޖ5���g���:f��	��K��V�|�{7��J�(���8���ɑ-�q�6&=���Oo?���J��I����<�j7߫x�γ�G$C���臜
(�z.}�m)��P������[� ����^ �'�(Z�P>�_���/�%zI��y����BScks��`��~۱5L�fr"��S�A�����p)���%v(hj�#��ΓWJΩ����5��h�Q%���^��B�j����W'����2zM���IUjj.d/-7�짱��i��r�(�����}�-K+!�#�z|��G��"Q����r����a���QO�L⚦�;<ѽg���-�G�N�V����S��5�+�=>ϸ��V�p܇a�R;�Lh�C�����n𺢍�] �����)_��\"�$�u��a�U�*�c�Њx�~/���W���p�Enc���{�)�0�]�]�*�������I����j	G��[�,{��K��D�����q؄��f�ø-����{�
���q�-9?�9�'�J�k�G����tj��"���ǣ;�h�~�$��a�8�?|�p7��=ڤù���|��5ح�^��ic �n�R&��P����>~�dk���g���h����(O^����4�KU��oڐ�Đ1�<?u�1h;\�O_����ԟ�GS�o"�%3�x�ˣ�I��i��~�¸��D6l��C�<�Y:)�6z-��R�v��WC�ܬ�~���Jg[�OOHS���H��5{]�x��-	���:mvUO#���u᠑!}��r�'�W��6�M��1G�7�_YH�k����M�Y+C����1�,	t�Н%ެL�6����d"o'��Xx����l�O�0ɑF_�����]�`˒����[�1��w^5t|���F�N%g7V�3n�]\����3������Õ� 
`�EC�:�BƧ<�An����EA��L�P���7�q�@k$)HKZl�&yX۽�=`����0	���XԹ��9��}�.d;�ѽV��m�2�UkZf���K=IO�����x|֐jQ��U�o�:]�Le��+��ԍ�"pe�8��:Fj�������$G?�I�8�n��V��V����[�X֛��Ӟ�"$+���%n��@�fPu[􏶈���������Gx��|s �SEH�?x	_c<�I#�P���2]�T�q~Fx<���T�øš3���{I��lً�)}��N������6��i�f��v;zU���m�,4���S_"�SF�a��ɉ�VZ�zZw�Uc��VY�aW�d�Mbn�k��F��g��Q�C�C�x�7xH��1����r*lS���e�H���w��Q�4>�2K$Xk�Ѣ��:�*����Ō���p7�����w��h�<Z��Ǭޓ'G�	-�Z�[����՘밆���Y�嘱���Ko�����v�.��=��ߧD�`,U1���X���kS����:z�7���]D�G�ߒ�R� *���;�u.�<M�S4��:.�&1�a�U�ʙ���S��I�\H�8:���U+��z�B�e,� 3�a�R�ur��1�W�1���x���O����@�J��+:tpm�3>��TWd����YA�Ax#@�1�����A���U�T�eF�ZN��|k�%Յ��YRĿ����{���F�FzL�ǥ��5�扸���W׀n�����DJ�̧��@���{+�w�r�n�%�ߥ��P!jI���U���K��6�v�{<�~ps���7���-]�`��˭�z*9��^����J1�M��õu�>OA_b{`��3YǇ�z���t�~��mU+ڡ����^�W�b��L�g��rн���b^7��w�Вp���6j��Im%��|t��IqҺ�k3B�"�
{��G����hb9K�7+}��<�GZ ���VGk����v%[���Ґ>�MS�c�[�M��bbY�Kc��E�-��h��I\U����p�N��F��BY*��;�(Hn^h�#���1�N�����3�xH����P��\�KQ3T%ImM�"
��?�!m���\փ���[dT׹}%�ߵ�!�R�Fo'q�h�#��n0�[3o��kO��c��o$�V��٣A,�t�ħ�,϶��#Bz7�%<����1�41�zZ�,��.��a��%����dK��١��I0���ς�/��&A�<^`���}]��ɬ��z��#;3�Q[g�%�B���rI�Q�?�&��H���(.>�w�5���ZAd�%K�gF���=�Ti�Y��.V���hI-�����B/w�=Rwȼ��?��E��Y7Xx��P�	PZe_Kt��D}�i����U�(D�gb�aR��A��3ި�Ɂ�&�o�������=;��v�<�L�R�%�#��mSxN��ncd�qS<q�y|!�r-�?|�
��R�BHxt�Ulʳe�3�ә��dۚ�):�ȓ�$M[��a|�ε�RL�C����˹�� �e�!�2��^�Ņͩe�]D۰0���M��?סE����W�5B!�/J�F��S[�+�-n_��x�H��Ŋ�J�^#�}�0l��Z�D�!���6�mb���#(�g��KR�z/>��G<ؖ����1 ���z�;�j|�a8s��g�m����KU�X�/Z�M�}Œ�h��P׬��Ɠ�S�A<,Ό�=	�(�&`��iCpO�@����â��<97�q���4O����CKDrqp�y��#aH�p��՞NxK�'O<�� �[x?;݈YA�p�ԇ!�\!��$8'VIN'i6(EX��&��5Ga�E��ﱘnt{k+94��#u[%�'���&X��<�a���mTZ�C� ��=����c=[o}Q�q`/I�^�#m������AE!��O^���}L��s�-2�&p�y-�q�guk�D,���qL�.�<Ѧ,�	��Y_�j��7��v̓�7T�<`Fu _�1�4֣i�5������L���+z2G$���M�9�D8ӷ%��R%:JR�k����Uy�vJ�~#�S�z����j>y5\�D]+\/��p�%��G��ݝ�	�-�v�EL��P:9˽��K

����M�`�=�FtF����AuC��vgǋa�ޗc�:l)�9�ʃ�rB5\+;~G���L��x�B�.W������k�0�?���о^<����K��5�&	���0�S�N�BY�pwwon=x���AR��Çμ�RDG΁%���]mW�*Rk�߽3�Gx1�>����w�h!T��xd�|�zM��^X)�+���w�ɯ�Ŏ1�h�p�_Q�)?;���#�K)YC��T'!70l��Sk F%Ų�Q9i��X�}�3"y�A)�8&�"q��Z�|��[X��JO҈ձ\���!��;���kg@�ˤ�l�f��¸��0�:�>���$<rZ�)	�f�Ή��W�zZ�u�\Q§���4�Ȉ�q(m9�5�����Xs�&~��U<#�Ak�� �7yѮ�e��f�VF��f�A���
�F0-:�a����@w�P5�Q_�e�O���h��9�=U�G7�5�b
g��L��,��z��c�Ԕ<yĥڷfG�ߗ�JnV����oF�ia�����_���K��*Eo�$�:T����M�ӳ_{�ɸ	������XH{�P�Q/�K��{��?:�������877�P0� ��F#��bg����Gv!�{��ޅD���AaD���k=����@�WtIˉv��X���i^8��g���l;*F�_�l�V3d��ʛ0v���.�k��P��M+�H*� ��w����TF���+`p//_������8 ѿ��_����:%<"X"�Fp�8�������3zrI�yY��<2�϶BCu�%�����!�|�%JK9�s�-&�������sd��{�0��C{$?aws@Q�1P��pD;���ߟ��<-����V7�Vy�l�wrQ�U����}�zDI�B������]E����{V���L.����G=1�AT?c�d��١�?��˥��"���c%�n����:�{d��Y)<�R��(�~�F�l�u�h�8��V���4�tl�=E,�gc���ΛgY��XX�I<�N��`�����7o߮^�k�p��G�c�#��1�AV�����G���7�"��Q��II�=x�Yc\?����<A���K�����c�i�nd�x�ך>�+Z��ٔ(����!��^eL��Z��4���1k����!����`j@�fLCX%����������~��{�P9��r�޹���߰Ė!����SON�W+�	��,9Zs3��*ˌ�^�y�ۦ���:�:PT696p�7m|.�O&�|��2W>>���v �M���D��R� [���d�� $u`a�\�Q�����3�����jp�����X����,����u6�?qo�`�q$	F�* E�%�L�η�����B���֪%$�:ޕ���f� ��mi�u�
�ޑ��nnfW�$D����>Ӵ�6�_���3ez�>H�8$c�)��qmV�Z��Su{B@4�6���RJ3��d��usV�5 X��z��R�[�!����G<~�G�/X��W��u�39�����dAU��s0Mio"�8����3/b�����t� ��3�0�ҧ���;rG�-N<�#n����\���7���~�C,�S"%ā���?���ca"�ÿ!x���1(��<壖yC*��C�M[��ΫZfk�����<�r4A3�������7��F% ����ِ��3�r� ��R�����;�Ϡی@��o�-�}��5#�_<���O�}����������Ⱥ��}A�(�vk�n����<�Iu��,j.�J����L��z� �~~ޘ2_�VXq�o+��\�MW9&,�Ƙ�ƿ}@[p@��mZ+�a��xL���ѡٶ>�]T/ʯ~�uz�Z�}�����g��!��I�
���B醜{v'�s'��A��q!�-f���X��&S>r�Ћ�X���j��2���PR�`�-�5�9�*�";���y�c�����<�Hۓ����D�j����&/�O��Hc�7i0'́vCߐ��B���4���v�.M�j��i/�-K�B�����
�<��Cn4"�s��m�~ ����\����?�Ok����+��S��T��� ��^3R@
������Vi�I���8T��_dg���x~>�hJ!�^�~]6�K�=���*��]L��F�}��5mO錴����h��=r�C��պp?��_���oH��2s����on�)�b=��S�|o޽��v��A=��a�3�`0�̋�_��h������Q�}Rz<G(�����16�h�aȒ�\e��p���>R<<w�k�]�8xD�s@B�G����V�mh^��{��6���#�Z����H����DSt�ƾ^����I�iӠ<Ƙ���GV�VFcr�l��qm��{���6=h�Ur:'�U���/�9����[4���LU&'�d��+˳Y#z6y��^�':����{dF�`�I,�~�?�$N}�04����?�H�J����1j>�?�;q�T�iF"*c<R�+Oާb����J�T;��(>�[�6�0`n�[eA(;��SՎ�X�U�ˎ)67���O��~Ɵ� �����9<n�4�&�A9(��E��Z9�x�������]ܧ��R{�,�&��z��q#�b���A�ԗ��h<̽x~�>]~����� @I��+lp�w��!����:�����c�]��l�����#�P)�x�N�$��J��4=ʹ��t�
?�U�z�d���L���2%���7�9�r��ߦ��kt��,�D	�]�H"G�P<J/df��(k�A�CA�W�|y���k��Dq\��Bk�Sd�A��8���!1/�=�1����6�]YVOd��I��"��r]2z���HXce��[�n-y���g����M�뻪�Bv��9�K6z��d��{	,��ڗ���3e�u6�E2W��NcTQ��&��'J��{^�����k�Ë����Vz�������=�#*bF�Z~�Ġ:�!�;����{�]�,����O�߿[3џ#���詍4_��H�#�m�R�T���n�OK3
°�Tg���b/��Mm�<ސnR�Qa�l"�XX��Mg5|z^s's�93?h�g�{�lIM	�rd��U�~��?ň��Ե�/�^�nDk�`���T;��∐/��������nt��Q
:���v�w\�3���)*Ԭ�}��{�W�$1�)$��b�Z�\���lc\�ZFnΛrA���Ȫ��[��2f��O�>����J>�m^�R������m]�E*�S6�kmȇ�2�Á���ټ���"�W@p�D�6ڤ�l �1���_|�5�X�{R,"�k;D����=��,�H<x���O����}v��THQ}7�i>tR��T��l�~(�j3�NzuqGM�Iy���l{
�N�ysǸ�J�>�x@�6/>���HւƆ��+}]d�o#�Ywy�ҲG�Bs��WkI����n�_���@�GRe6���9����"=s�v�i�r�5��A�h���k�S*>$�&LĔ�n�کn�P�\��Y�SZ�Ţ�����.�+)�23�t�����(7�8������O?�_?+��M���`f=!(�[��Ys_I��DY� fp�����4�"�9 ��L��pm�i��o6YJ7^2H�� �@���]�<E�34�2��:��$����q,�|� �Y��/����f�G���dS�IcX�7T�8�c�4	�-m/^��}���!+�h�3�q��p%B'�!�K��"�ĵ��7{����տH؁�"Kƃ�S�JY#�@�m^n@(;��e�<DH��Z�r���y�U��Ӈ3"�~�a��M5��kVJ��\�_�U�[���6�OR
�=;;�+�7�=���z#xj�Ԯ�R��!'�2΢̘����p-�����܇��>NN�]���De	-�Bi���6&�/__3ꩮ�j�M˥���-Wn/��^e�H}xG\��~���f���^�y�i���>�UDj���|d�#��uO���A��>�Qܟ�l%=��(����0ZFU����/�J!��g+���B����kX�p㹹��m��b��4��ī�p�����xnѷ��-�4��;����OB\nH�@�g[��d���~����:e��S�̹����!�A-ڷ��� �fveo�3ek��z's��3��)�JZ��ޖ��<�We�,�7ia����{Nՠ�7�/����'��M�i�4�U	v�!� �����x|H����8o7�k}�s�kԅ�'�v���� �C���\�gi���24�pq���7)Kکv�w����{B�����-��s�n�s�b1"�b�F*r�A���ިI��;6�M��@�Nϙ�:����ʘ�.2\�P�| 5�"�4j9�2�T�n
GY���mW�YAH)լ�n�	�I�,�}t�*�;��M�����{j������{�π&�N������q�O��12����=B�x�0�Tσ��^�0}�=jvl$�{=:>%��{]e��Sl�l0]S��k�����fecY�����61Q7i>�0H5�p���QRٱ��!���4���-�6����?�4�ޮk=L��sBi����.ޫ'��9�NM��c���{T�x�!�Y2֭�E��Ԟ����6�¥t2�>�}�{��r3��q����QS|(t]�R56b0��k�w���$����46��$x�"��0������@�ߜ�=��Y��"�DT�x�x���V�̦�S�9�
������z~�3�JPl���s�& #�N�(����;�N�h�Zr]�[M �ϻ>�(�;�}�V���w�:(�bL�ʙ��u"thăA�Yd����Ԕ�վ�'������4\�ƹ=_����n1Nd���6�&v��.x��&6�9�/փ�Z|���f����7kP���^���F#E8W��4��/C)����@�`&��������^�F$��L0��L����I�n��O�Z�T�]^�[n������7d��,�7���=�{	�&2�����ʩ�6x�P+ݤ;���8,4߼}0	g�sE����d|�v'M���m� �Pj�Y�Z�)������T�_�q�";��O8�"�����[[�����i��GA���*�g���n9�{�� �03 n��������c������{>���ށ4UH�(]�d�.� ���i�L�Q'���9ڃ�Mdf󼨣ΠlФdX� ���k�nx-}H�q� ��,�2�c��ڌ������.J���hl����7G3�xed�k��x�i������@�f���gE���1�GF*l��S��x힟��xT �Q�E�ꪂGTm�4aG
�ǟ�Ok�#�c��Ypx�k���W/��,ܦ&h��^7ҫ�)������/����Ӱ�&6��}Nv����f�Ζpwv�d ��Br����K~��G�Ƈ���W�E�����H<��e��f�i4>����);����c���Ư^
��E��E���i?������J�����	_��%f�[�_gg�tI	��#�;4�( �lo��25G��~������x-�.R2z��F� p�#��,��^�qP �?���7>{�|%jE+�L�"��F4�~�k��y�'#c�y����׏�bK����F9N2�9(	���)�j��p'�P��\z��J�\m�,<�CX�<�[>>�bz�C������v�W�� ~��.�lnY�x����_D����W�رP5��+l�H����M��q,f��,�ܑ[vV�WX��Q���  ��IDAT�j\A��4�އ���Ɋ�e��N*�^�:SL(���%�C�����놎 �n����Q���b�g����(-���Y�?c@۰!�S���������*�����t�qܬ��2ޛ�A�t��=�Y8��Iy�RX�2� ֖��G��#�����Z��<�>��sj�FB�Q�acX���5#��6L����Z:IUT(�x�Y;uW0q�l2�a�9�X��0ݒ�~�b������B�lKX۸gw��b�G��w���� ;�z!%�=28崊�[&2���H^��?��u��y�?�?��7�H�\��d�X@rd܉�*�q��2Iź&C��S�t5��s���ٵ�iP�'�n�M�A�9��dx���t&�]�`d��F�nr��Rg���� ��iP�"�̬йMdȝ��b�b1ὁC&(��S7�pQɢL,��nt-�hL1}�A����_)KJ8I�Y���yfv��o�	���@�>�6�cV�ҩL�'*��k��d��ë�laa�y�QC3Ts��p���娍'�	B�iʱ#��+@̀k�C�R��ɕ:�'���޺q�+���& J�	D�=�,{^+�=�����5�=��j2Ξ�R+~����-2���JG�F:<`�<��������{˹X��:���x�JSA�w�6�̾�h���ޮ���@�0�A���y� �HX���x��l���2[4�}��^�W�f#G�f"�L�ȶ0A"����IO�� Ð��!�H>&�S#<AK�.	��iq��=��zʳ{�Ѝ�\OW�)\��V�r�י�e�����]e�I%q>^�,����r���A$|wB�����h '�cR\�  {J�ܼ޺�<a���%���鋛|7�%>˕�Xt�Jd���үsP�:|5L���@�cd�S�)v�{�`H�Sj>�3}�Դ�_����}i�IT����	��@�>�lO|��͛7�0�� (�I\Vttt�)�u��pREBJU,#��9
:yQ�H��	i��yI�f�,��f\�\0�1���I���=��׍���w�Z2��������_��:�D9��%��c��0[��X,1�����x悢�����cU�^��2\�r���=O��Ll^�N"���fʦo�����̠�{�f�� |�7�s�P�IN�fu�E��̓<fUT�G;/�E�q-ll�����G��Á����o�M����ʾE��k�T���������3X�TwyEC黪p��V�)��1������N%;��B����	l�H�T=Mq����L��u!�y�:���<4��9Kݍ:��蒖EEE�~��E*���I���+PR`.t�q@0�d�J\ǀ:��̦���r��55�bZG�����ΨF��/���#< �����4�JƲ�.�-�Pd���Ȯ^3�wo)t�
 &� F�X*�Fd��׬�L.AZ/Q�u6P`��N)v����sZ-��c�m\����-���9�2L�qe�&�A#���ƳUH`�3�S���F�Ȓ�5<P�ny��L���n��_��:F����H�@6�7o�C�m@Ev���� �Uȧh<t���2j�s:��u�|МT&S�,g($*Ӄ#����.��p<���xh���<e���o�7VM���k5*�����!���5�����1���L�����Xz���61'O��_�;���S���̮&��N�^��@��$p�)�inZ����?//��9G6��	CZ9��������kje��0h�5f�Kn�]\������eE�4/^�����8U�4��ct��5�i���|����=��̑m>�'��=Ć��).R� C��Uû����pi����-ltE�Ҹ�!;�|P^�麉�E��8<��� �v��y?@� �TI�˒S�*5�Tv�+�M�
�q���^Җ:e��v�ll�f9��8�{�#�s�y�6]t��i���9�wg1�j���e�of6V��b�����!�1y��������D�C�v~����;���ohrML�L�%��G�<������/)?���z���l��'vr����sv�c̎��`=�u��0����qD�;Fs*+���ދ�CW�I������{ �Un1^�Y4Ҟ%4����vIw�s�q�l߃$i��TT��1�����%��U0mzBei�W���]���Y �򣒃�Y�t��TA���e�Y�,�m��9ƣ���v����9�#Q�pOO��>�^�R*O���i <7��.�Z�#���u���?�����G�Z��y��D���n�AN\��B�_<Oo��u��������)3u��~<t����pٜU�^B����[�.#�B�v���-7@:}^�����ݞ��δ�|&tXq���g]����5�.��΢��}���C܊�n�܈T�B��y*�����8��2=iNW����=x�?���v���R�|�EzM@ ����N������t#͎ME{LZZ׊�n�!@�ݰ��n�W/"���a���^��'��=�=9-G��$��)��,��|i����(�p��_��)l��Ie�N׌G��1="����dS\Ĩ@�H��o����߱�T�Wѐ+�C'?��0�������῀Q �J,]�"Z�/Q1`�R�!� ~H�gڮ�磃�/S�������{���δ����n6iO�QX��>'z�u��@270�} �C�$����(U&�Aa�G���$�c��͌4��m=OD��*���S� d" ���¥���w�}�"n"�Nx�?���j�[6�v�������ᵂ�h -(P2ƍ������1�mf�Sz[�.3�As�4�2��ͨ t�XB�0]� �d�;�ht�� W�?с��N�J���K�A�seQ,��k}��!��\x�UX/�ی@��mN�%�[q�Dr�{�(��D�?����T��D��ξK��<�!���ᷱ>�p��e]�U���ݻx��9���md�w�M$:^\_�}�bx6��ț������F���Z�>��;q��q>�]_3�ب�z)2�g��l�7�B�'M�6zf�gcȄ����DD�14W�BS���1M	FҴ���e8���
� ׆����g-Ł���5��H|��E��gbq�O�Y��/g��J�ַ�`
�����ũ@��j�E��:����j��l�4��倬I���g�	�IX��'66&2�m������{A�;,�v��
�������'M3�i��ٙ��(�PN�T�	�l�4��͛M,�ql�M�>pj�̃����5�.9�&p���΋� n�QV.�m��O�w�]R��{bgL9���[�ݖh�LC��������Le��0]_�aNp��
/����i�f�e�g,��4޻�nyz�z	�*��%�2siJzu�u��^S�ȸ�G���IB�$U�%�3.x����=�)Ԡ{�aX���0\�j�{�iQ	�w٬��w��~���Zd����oޕ�ݻ8���Տ�K?�����0�ǚ$��u���U��.eV��^=�3��5����<���:�������t%��J�ٛ$�8��,����s���Q��YKa����H����VR���5�<}�0�$�yw��7>�����O�0Dn��X��,nT(k<����rgӘƬ�4�_��MsS�,����ѿp����o�$bI��4#��.�PV�>�CZD�h����t��l�޽{_ǎt���6[�"�_��3�!�'F\��<FF�&��.���Pe����`m<�O�M(��g}V�dWz�ᘐ��\�l��t!C+X��/}�˹�"�w֜�P��4����Am��f�v�G���57���5��x�,�3=f�Z����+ �\7��þ>�g�lL�`l��P4����?����6�LLn�9�N�1"�$�� ��K0;�-F���x �	���0�9��M�C��a�A@CdȌAg������r�vڧ��d�K�䢝1��"�dr��؇�ˬ��Ԇ�BR�W�0���^l�����x�
ѕ��v�	�,�#\��q�A����4�)s�w�}�����F�q��"��v�������^������*��Β� �B8����E�e8�q@ ~��u����ct:�'~� �����s��N���!�Í��{k Mw ͕�@��cd�n�-�r������u�
���8;�8cB&�{z%2��I���Gn�x�:^�מ�ާ���E��Ѹ����3�������x�$V'���y��c-�Z�.����Q��6+����7�>$���웛8�Lg�'-�;}�%��K�S}ςr�"���J���Sx��]|�]��P����)�KxP�`�����p�1u��l���O�
��1��%G�<�5мz�����&^� ;;{��=�"ϟ��fS1�9o���Y@���˸��a7��rl�4U��O��ʊ@��e��C4./�Ĩ�y� �iۦZ��w<S�٧2�Hz6��Jj�:#�z:���{����G<~1����gU�J��y����
�>3T�j�,��z؛�Ƚ�=.ǘ�0�cVOu���Cuֱ��ٜy�5#�Uٔ�8�)Y��9]R�L����|�4�UB\t���)q�C�a�QUʧ���S�¨�}r�X�ȷ�>�@�j���P�H�T�4vh�PH5�Qj�1)>��JF���r�,Kds��4����bZ�N��(�;,M��< 7�m�I%d~��_�o��Ɯ��<�\��Z�����l��Ag3�)�h}����aVs
;��Q�T�C��Qg?���^r�
�P�B@o�9�Pv�!%~��C����I�C�ּg��z�hT^Z��$����&���@w��8(X(�;���7$v�*�%�sY�eLU�M�n/�_�u��E�k��pS*�(����~N���(���^��H����繦=y�l;�5t�ٜ˘�n7J�S�i�ɥB��|>�<��Ct�7����C��4[J�y¿��㫤� (��a[l64�Ѩs��9dN7���?r��ɖ�"[ec�PKב�K_��(bQ�ݦ\0�J)�I�L�����NA�pCe��y�'����%;5J&�8��ѭ0K=�Z�ob[E��P��(�����)�C�7|(٫�dj�t�.v�5�j=�c�_�j|~���ˀ{yO��30�[�ۮU�^>�PKD�/����eo���/��O6� � �x-�����B�_\c)m�4�Nj�D��իxo_}�yK���Z��rj-�/m\�B���F��1/u�iW����l��2xnwヰ���ݨu���FP)K3]�(�euQ�b��"�ʱԁ��,��8�zS�W��(�>��oo�z:��0yϢ��=d��L�ޏJ��0��[��F���DU�����������<[��&�%X&��s�Hm�՛�R� ����f-����#��w�%�mf����`p����F��w��3�m��/6b>��_�Fq����i�,\�r�
m����9�{c#+]εy�����K�P������s�A).�exaFCO��9;�x0�1�8�F7���szeE�#�l�q��Z�J�1wn�����M`�+\�S.i��k�G���������#���U�ڂ.�GIl׎a̦��+t�] �0�I0 ���d��	RB/Ѵ�B-�!��Ϯ�gt�c=?�:�������X�Vv�o�^{!�8Yf�H�'L൙�r�`Ȯ\���L�}�w�s�Ჾ&��zB�0�e��ե6�t�XQ��H�N�aB��%�Y���s�{�`�T܋���1�\��>J?o��g��_��j��ZB�\�i��{U����Ѽa��>�{�1�'4�g���|N;$�2>gdU�s.Ve`#��2c%�Z��a�%��\S�����7��ￏ1�(�r�[3�_46y
��4}]0B���>=A���ӳ�s-�Z���3�N�����aހπ{��@6�+��/�uV��R6p(��]������|?��2�*��ޠ�,���3�G��of��~U��IHA7��}���bd�'�X��(��p�;+�>iu5(��fD�7]����m��Qy3����=�������c/K
VU'x~�x�'f����嬩�;5˶�����G�:{�9���O�t0+����l��Q)��1
���t�q��G��s�N�S�A��B��%2f^@c[�3jk������F�P��e���{��{��QSh�X�����{������2�~e UF�~�ϊF���SV��HB�a��H|B��ף���a��R��1��w��t��m�T��S�ĝK��(�������RBͱ_B�B:5A���Ҙ�&7!o0��}N����Q�\��#����GuB�Pلr�E�g��%�C��8�B�s9�ij%�&~?��͔�c����z�b�Pe�<�<��TY�L������3&8��H4G�Sږ��Ĭmּ"��S_����1�|^|E��cx�yFv�q�w�cq�[R|��,� ��A�eZ�3*��hpr� X����c��=�mTmc%�p�5���������x�8\��#��# ߼�5qWvp�:��`�%#�J:��#.H� _(��a�e�{䁊;5��_v0D�nB�}��(w�=fۣ�ݔ�{r~����8\pPڐ�b��<i���X>N�\e9cpUCx+����9�me(�Q�p�;��t��:�u�r�ZV����c]&-��ԾϿ�1~.��#���l����A8-Ё�ۘ'�7SNs!?��%g:��s}J0���tȠ��6[�����R�TJ�����1/(�VU��S6d�
쫗H�-��d�I�8M(Qʳj����1nX-h,��1,�y�*0·�徳����o�#��]�FaZqO�H�����W)�c�������r�#tE���MP�ύ;�y�ҁJ��Ԕ�݆��5`v��4������T�и���$4�n�v��/Bݑ�q��UUZ���b�ڼ�ݜ\J��&��=�x�<:����x�~�ז�����LX�g�ꐥT�7�԰.�׽gO4�&Py��Ô��N=���}b��	�����nH�C&VE���z�׳��OB?�G:@� ?iƔa�pӇ���ZL��� ��*@e_A��TL�F)7e�T�'�NQ}!	��W�������8��"�MiL-��1�tQ������˥�UFZ��O�!��kd����b����垀�nwN�;�]��_���]d����*>
�r�\5���V��� ?H�N\�F�z;6�塵�(�l(�σ#�Hi�6E���-��-�#>o�q� �	v�E(G@�w��&�,j�=i�Tjꮃ3wf��m�%�NM0�����|%�p/��qp��%�������e�Ǎf����
)c�P 9P��js�Q�)j��%�S4q�ި��8���j��8d<6`眗��
�>�A�n�ڇ`Vȋ���L�m����&��7(OXs���(#?�����\p6M�A2�J������r�=wG��!�]�b2�� ޳M?��>W�XBi���Y�L� ��x09�0C�DNgһ�����!�7~�Y|с�=�=�,y9�2
*$9�!]�S����:�szC@bK��W�qV�H��
-��B���pdF��w�	�����k�ee�/��RO�y��V�:����x���M�bFK.�%7N8���� �XZ��0TR5���{m�Pf��?u�!p��"@�{�K�P�����h]q�,a#����3Iܱˎ:��o�(v��ZP6��j�b�4���0>�B���Xz�(n(�3#�n�����@66)l�'�����rB/jf�MCI���0\�Ѻ��t|I,�jQx�5�L��Z�u{I��t9�D~����t�4]�q����[v;�!e�Y׉6�8o���3)a&�#��_J�����=6����q���i"�i;^���]�3�����Urͮ�����CE$u
Kxm!j���BH�א���$�e{��i���ʄ���
a��;V7���J|�~��E}�/S�ZN$���E�Z�h�^s���>隆��8��o_
���h�$>ϗL���	5�X��p�J���Ѡ��-e1d �D��|�2�0���!�	�Y*ۘ��r4��BX�G��?_�_����E��!�3�<S��?�zU��(?��Ͻ	��P�!L�"�gGXM,���u���Ը����� r��������(s��zf�t&h_#8t=e��m�OFz_��D����W�	��F�Pcj�G~1���7�ƃ֤*#���r\��?��)1�]u��1ѝ�N\>��|ݲ�ܘrhc�b�Y��S��@��iN�I��	q�"31�]`uU)V��#������c�}�˄Y3�N�΂�#v��B�?����Db� (:Ճ�E�\L.�&0$�w�%-'6��jz�]�%e���+ߚ�C±�6��-�um�罕)�������<WM��x���3A
��eɑ!�B:O՗8̱gK�y��)�%���%wG�������|bZr�3м����%ٔ�Bt+E���qX��F��Ŝ۴��B
�c(��7"c;�?��z���Q�韙�t���mb�������������O���Wm[�j%��0�gR�m�M�X]��42«��
��>�9~�r��N�:�����������x8�Āc���Tp!�g+�rB�%�w�l��R��R:�BL��a��U�O���Lل�Bi�Lk/���O�!Fq	tIg�����MY"5Jc�����]��a��廏�1���ȶ1Y�-HP>�j�I
ZM���4�5t%�w}O�AI��ˠ��4�1��i��ω�{<�
�,)�<��b���+]�$Ss��l�Z��^�� �i�a���a���.q�U�8	 �x����Շ�,����ZJ�7q`��J���(�փ��o�%���{�@N�T$7�������|^�y!;�6&/9a��p������ns��BQVGu����g��Z�/П���S�|��l�'��Ǽ�Y́o��[�9$CdFzmc��,�MdtpQ���sm /������s*��De��!�x2?[��Q����_԰����됐��]W�J9���Va�s����g��8Qj\�
M��W?����bX�ǂ���#�ۧC��uh$�/�{h���]��54�Y����9!�g��.0�^N��
��E&wr��%���l<���ku�=�)�;��.Sy�J�<CC4�,�9����ơZ����C�ČRC�vG3����c�[�şqoBEt���A�b����p
Afe!Ǣk�(7,��تa�3��Rg�[���Dȧw(��w�N��͕�^k]!�ڿ�� ��!(����:�`#f��}�ǚ�ʏ�gE�J��,�7�����m�݄�������y�0|�V|`������)ب\���x}��K���Z�c�Q��"�#�;񍱗<`��{�HkR�_yt��/�t�G��5�Yا�x���췴8I_,]���r��$U��L3Z���F�;NSv�q!�Q�l�����Y͟j����E�,E���D������˿�K���')*J�6�lO������&X�y� �GC	c��o��>�(`��؜1�qsT�rLuFˋĩl����)�܃�sQ��}����bea։�첝��v�� 6�~a�8r����r��F��������-�{����x�F$�`{��{|�>4��&O�"{��)ǛZ�.�{ġ ؘ4{�!lp��gNk���oU�k��I�KWK���tY�� `�����n�"�k��Q�{ś����x
fs�oD�ǃ㖗�4¸�g��P�օ��C�	�����z#�\մ��g:��{�]^��#���a���5Fx�i�Q�u��z���ě#�jz�{8<� �դTX���cr�}@_�3@
��Р�ܢ�J/��2qH縠b����}p����}5_����	��<�Z����MYr�D�/��Gi���EnB��3V�b??>xdk/�'��\���V~�8�D�Y�����p4���������% k�S7y��d9.�6@j �F�T5�O�� e����Mt���Q�Ar\l4�ؔ�pѱ�
���AM��0 �ѭ��(���mw[���V�O��	|Q�f�tq8�\zPM�\�WHk��i����N�6��ME6�k�.?6�[�s`����׈�͑�!��B����.�~�B�4��R���D-�J17�"�N�܉[������q�w��ۻ��N8H���=�|j m�|���:�_��9������ب�7F*,��ڢ ��{$
8t.�SAv�A��m��� �ݚ���eɃ߭��{v�L�0a�X����N6á�i9���1���"��Qm��^r���������k�~%�T,��7`��#�l������������s.i�]R$fO`�~���8xZ�:��U Ŭs�z���K�!���6��ޏ����o�G���F�/Α��+�ÿ�¤��m�t�V��}ē�r��`t��,�3;�$���D��ɕ��(SW� ��]WUD�J�E�O��|j���I�<��Cᢌ��Ǹ�^	Q<z�عJS��D��7�؂���wmv��.�ki���8ib%�<n�W��p���3i�i��j��s2cVaw|���|�����ׯ����C��;"-�u�k�Om�$�c*P����&����	�x�`��P𡑶�MvU	5^�W|�m)�����Q�L�g��G��*����y�؊�X!���4�{漮��!��/�7:\Nɚ���.tB)�<��멼}����w�����a��c���Dbw����\G�8��#(i�d��s�R6n�U�M���ʳd���s��Z�S�EG�~����H/��-{��koL����#7��}c����7j�I_M��f͝���p'i���#��K���E~�ˋ70o�N��3����� �}�@�m��S|w �"ri?�ޱ��4̼��:qxi*ۺ�Fe��x+z�e�u��R�}��yMR�8Иa��M}iT,6�%�sNvE�2�3��XI�JM��q�kz�~r��9,���I�:��33}ln4�����T����TM�cvq�5�	O��bTg?~N�Lx^d�}牭�ܤx1>�����p[L�Z���$�s��e6�U��7f9��q��Q7DL`ϟ���[� ��g���5��E#�Xg����r�Gq������2{<��h(��7�_�M֢�g��rZh<���Z��٘��5�zU�3�N#��X��Y�ƕn�JKW���BW��o��/�F���v�L�Z��_f���k����=8[1�[$�V�ܦ�	$KI�l�#4��P�ؽ(;�]ՉO1˽\�z�N)M,���C$��')���0�қ�t���4�c�C��M�F��1ƣ����AP��*Ӈ���T���ث�H����ϟT��i��[>٘}��y��,�/�G�	����w��֔G�g��P�������4[��AAC�a#f3!Lg
�R����do�]��Q�G_�&�d$�q+��Xw'݃�$�08�s5Pњ���D�E�7 �M}x�>>�|t�#K���DI�uWk��H��`7��S/Ϛ,̹�b�&���k�T���P���)���ߧ�?��Pi��W�ք)
gOzX����k_�KӨ=-$�ϵ82e���n	pM8��`A7�iߌ4��:�=��C6{��)�L ��߻�@�C"t��!�.�PCo������!ƢT6� �_6-�L���4;�CU�d ŉ��<�v;�9{ub��)O�HIk���"�C�,ߦʁc���y������e�N	)D��4<�@J��8�Q�z�����r�V?o���n��?�ø����(h�`,	>K��2(2P��� F~�N�i����+LR�B_��L�75ɳ��6�L=�����C���O)����N���U)���C����$�^�xx �4d���(G�pFGF�@
���f�C�Ӝ�p���u�R���eP��yJ�y�do�)�ǰ�[����^�Q.A��n�`�R��X�R�B���F�z�gk7��������E�Ǫ�������f@�����s�׿�i��瑀��ϣ`:r�H�&�A���.�=t�'1�ݡ�N�T	���i���jrժ\j�4���Q��Ժ��!����U�:�*�0��G�Z���9$v�2�)�5��u~�)�G����G��b0��iɧ�0'�R�ύd���F��9{"[��%3�&ѢM������ba��&�13dΌYRX�%�����2�X4C���8��1���:�����^~��+�Q��.�bq^�H��"1�����Y�Y��_~�K����ğA	�m��e��D�F�&3��b��K���pֺ����ׁ��L�`<ݥ�;�Q���LK!OtLΤ����)),-���3L�w"-�n�5�����f�SP���gKS�ݞ��+��9y��bc���=�/iE��Lb�jB�0<I�c��)5�x�����C�͖ţL�E��w�ςA�Q8��
��_eé Cu�L���f�v���A�l��;�4����0�9J��ի7���]��v��Y\9�Fօ�&B��#;�χB�ar��`�$hʎOnz�y6����)�yl��oX�WVF�͹�20	"ͅb�ɩ�.���^�����id�S&���5��At��������С)u]�58�<���i�����������ߟ�)�쥧tiB8V�h)KC	*�d�E�Zӣ�[�պ�*쀅��>6�Q��(7���L(}4���#�z����nD���	�}�"�T xo�X<�`/�%��*��({�u�(�9K����!Eg;LN6I���=��'e�������f����qU�%��@K��UD=[���w�&~��jr(�F�$B��(3r[ٍy=��j�209�6��t���nw�TI�,oa��`G?P������3�M0����=F����Q��̨ܔu6ۇ��p`�2iO{�%#`T�Q0$� �eA�+h�Bh��e�}��jK8(�,�<M	�:����F�HpY�1Cޕo��:G��w�:2	[��.�4���}��hw7U���,��'2�o
Z�R���=�t��Ǣ|����o �g0�M⢥\�@6�`�W�:e�i` \�"-��H�V���u#����Pv�K�T�Ð�Sz��E�C&�Ax��A�1(Rab�����Z�bEc���6�u�;̞�]ދy�O�(�H�q!Q��.�ٻ��#(>�{�.)��N�-���m�I�jfaC���cf�n�~fj��cc­�.�q����3�7}���Ӡ��H�91Zl<6�ٓ��o������2�,G�ɩ��a�X3��6��z���	�ݚ8���M�떪�G?K�1�q� �ߨ)�,��}`�E��r��Ma�?GJ�T�M,g�{$*c�w%I�����HI��1u\�#G3���ڬsG��>�~�f:��2O9t�Q�,T����˹�#Q�E��[�\ީ�|*��KdȋꦮƠE���o��{笌�J��L�B|i���xz%��_+9�7��N3v�6�°d$��W��ZA���6Ҕ��3h�@jl՚�O�@y4�%3RP�`�L5ԟ�ׂ��SZ��ցy�]P�"���e<�}�����8x�_�|Y^~�R�Y}�YF*h�����S�zr�J�����^H�5��\P��{Һƫƚ��:�F��6j��s��{;�.�x��:"x)�O��tH;1��aq����k&���&��{i��4¸-�)��R���������೸��LG+��(U�8Q!��I��ԽF`�D�&�B`��,hj�q<hz�e����{��̢�s�3�Ѹ�T����*��$n��YM>�Uͺ}�0k'�*]qM�M�����9f�Ul�6-8��%OA[�^��e$>�yrQҲ����6�9�i3z��$~S���?���ˀ�{}�T�F4}��:�r~�E���/��긶/C5%��>�)��4��a�;~n�"���Q���gb���X���dUyp���M�yH[��a@��`�pD0M��ha��~�L�$���\�7oh�w9�=`��nG�~�\<72��*��d�4��t�s���l��xz�vI�����S;ez�k�ZZՅ���U����&` Wu�4 ��d��^�L��;�GSi8#Y�OY��qh� �
&�w�ְ���Q���@���'�V�P��"e���ɝ���.S�}��S$�i_���ma���<��e���I�gM5�����q�OfdC��ݣ@�<
���8��+��6��PP@�M�����J&��(�Ϝ����A;~Gzx㎜gE��E-��;7�5��s��9X!���`���Њ���P���Xe��	t^�~��`\�(?`ܣHf�J��������@M�&���(��%f��c�T�\�_���i��$��|J��b+2eO�R׼tT�	�1&x����t�� ���E�.�Y0���X����1�;.~�O�I��1�tC&�����3@*?<�����a�N����E�n#J��6!��jp��5a�!e��еi���:����2mU�����X����в�E�_��h��uF���_}c��f��ݻ�A��{��dp���Wk�r4$�~n�z	���.4�E���L,0K2�pVc�u�~�������}#����z�02&�߽KF �iQ+A���.���y��9���� i�}���O�l��oބj�Y���e�/�����|�T�cT3��ٷ���'�9��:u��\oBz-^~3����ԭ��V��k�I"�^��HT=9C��$��jBWnA[��y��:��nX���]����Q����/=W�>8�h��yW�y>/<F�����������)�Kk�r2jb�������*6_y�5x�M� ��e�jM{5��䘾�-߮����F͎��4N����zc׭��.��{�9G0%�T���/�L4��	����N9.�A4n�h/Tނ Η%J��Z]�8��C$���T.;ϙ��O�cf�X�W�eq�s�l���I�;�	�M��:[����{�����~-0�x��AP�j]�_��}͊������s��gr
��RC�1�(�ޒ�d������k�]sR�T-�u*���!�C���zf��ob���Q����&v�����Y��~�J���V��ր�xV��l�O�p��l���`
��hT��I�!p�B�|=����ൢ�h�?��<`'8��/�������
=��<�-x �O,�dӗ�ɣG�)�W�P2]R�Ŧy��yHG��O����!9D���"��T��ap����t�_�P���´q)�,���,U" ��^���S5F�dH��{��b��^W�ѶYlĢyN�)������b	5>���cӓ�ڟ	�G�6�\�	���b���<,�ƴ��]J�d�E�>2?�/&�#��	���e⡎-n ������D�v�n��X�c�N|?�8�����Nޘ>z	�v\�
��;�krΠ��vѥFP��B�rXb���C6"*��K�6O�5��*��ꌶ&"K��gͤ!.��F�-���8U^>{I�����0y/�w`����3���my*��k��yX�.��U]$L����hY�y�$��1��4���b������ߝi�����%�Fa��o����B۟42��9��>�kd�5�	��2�sJ�Sp	튏����VyE��(cܰ�M��(�Ү��(�������KR�ĩšV���N�l��9�����kD��ֿ��`̭�4d1����#��\f��M�8��Q陮
��93�(�������lr�%H������<�.��?tE�8�}��i���icȦeD���̹�~��ۯ�����^d���u�tW����5�h[��U���`� ����St�O������oٵ7vbɰ(���$ۄ`�Y� �eh^�'�޳��;n>6~N5��l`a�ൠ�ƅ����p���8ت_0��y+��bd��u�F��Nh�(Wy�E�-nt��iקf�x��6T:Dm��Fd�oww!��q�q-��Π��}A����OGL/�YDq2�<l��޼~CK@2��~�Ҙ�Q��W?{٤@ ��N���SX5��"34_e7P)�}��Uu��M�z�Aݰ$�n��ǎt��anbm�����gF���;���{�+d�����ee�9	�1� N�6ȅ��&��	�����#�:���`��N�L��X�//Od�p���3�C�0�:<�<h3��$=�7��x�K�q�{=���u��D�	�~H7�οW(%a�c/�ى�D4��-c=��N����0����cݜ/WI����e����9.��\��`��|g� �1�X��Q���}5^����k�\�'�Q: z�4�!ι �ǽ�y�ۃ83w�RG��P���^<_nt`}݇Q���$�j���'(�1+H��1:zs��G�5�y.[�M����T��� ںe�@q����c@��M�8k��J��l�3��D�i�i4���%���[xM=������\Ap�a|��2��=�lU��?G{�z ��7�Kғplnh}������%�B�l��ETdڵ�3'����q -���^oQ��t ������S�/�X+Qr2���`}Y]��bH�х��D�sC�9��Cڽ.��O�������7�+�â��/hj��b׷��NՃ��.J��m�"�/�||�]D1�ؘ}$a�,S�lOlP�̃�`���;b��m%4(j�у�%�v�	�x�{k�q�1Lu3�&x��m:�?�~8����_�"���OJ�{O�I�,�A��뱔a�k��|J2N�	L`l���sK��,��"�h��?���6�q�I)=n�w��@��2�#f1�s��4����*�?�O����\���m�gԔ�^��|�ds��U~J>���]�6��zrm��}(��Y�s[�-�4��U�^6�4;8lhA8�\޼}�Q{��7�|�	�'���L���GtP�M��/��|�k5}#������HsJ�а#l�o2R�Z�!������t���
��dD�M��N��2#��%O�c���ۓ �1�ۻ;f��#I�XS(ɷ��H�`�lKgc�c�nY��
(�?��� ��`���t?���#E������w�>�Y[��$Ɩ���S����*N�}.j��T��}�q���e�g��pRj =�S�@쒝�eI�'�e�s��2�T<��$v�]= �������z8��[v�C�+�DP��DgTƋ{eU�M����	�Nn���|t���PZcg=m�I8f�Ј$6obn8��}^[[b�o�8#0e��+
�Pg�R'���;(w�)�<^�;4��0��2&��ÔX�	f+���N4�1^�?�&Cʦl#OluLS�=Ԇ��Y$xR����q�)@�_�I|ɒ9���;�� �mܛ s8��/1/(:�}j�M��J%v������]HRw� ��l�����4�!S�hP,C�6鐟�Ri#����C����>ǛT�Q�p����-r��)�l�1�,���Sc���x^J/��yxZ4�JQ�d���d�}=���	���5�NE��~?�3�ɦ�u�99���̢��8V�2���2�1�q�^7m�`19]A�����
G�u���z�~��8/M�#$�rU)6�!M�s��fa��/�6h�$�9أ�h_~q����V���2��۵����Q2�}Z�7�gw�?�<�����MK����V���������hAW��p����X�7��8VsYq'1�`Q*}��12g�V!xpvc��774�؈l�j���R�q����Ŭ��'捌}�an�n�^a�M-�Ge�|]��j�3�M����O8��=yp�����x��������m�d')�Ț/�9u��Y��נ�t�}17�gR�Iɬ�$ek|�~��\�����������cuB�ы�`W|�%�4�b�kGl�jՃ3�����RG��s�Kof��۪M�8�y��.KTA!;@|Ƌ��p_�t�F6in�y��9�Q���!�	4�R�R�,k�#�Q9�ψ�4��f�DU�K�V�}�!�G#�t��D���e�r/���W[!-��}@Y���:�
D����U�a-���|��$����J6ע��xq�!p`�v#�NS_��zK)y`�튰C�Uȭ��B��ӱ�4�PyR&��d\5Y�i��_�O����c�ϙa�ţ�h��|����Ң�)��Y�|�ߔq7f�՚�0nw�fUW(���P$N̹���9�@�AP��as��_�%�hO�!�Z�,@��WLU�D�pn
�v�� �_����(�F�d�L�U��Qw�T�ǧ�[��^��hnXmЫ�Y����H�!@�M���1>�t�~�+�	����a�~����JdcX�Muc/n��������wa���ȝ� z^S��is�d�>��4:�ض��颬p��eI�/d���)��Lǥ�T�Ȧ4a����4�=�χ��V�2�Nc��gK��h�xl�骢sw�ِ3N�{�I��@�D2�V�H�H�@�n7���@������a�̾U�Ͳ����4�[ȋ~�4�麇 h�ܺb�����,�&-��@z�h�^6���=�g�,�ڇ*T�����8���:J.I%uR�Im��Sgm�ߤD��D����ʐ�T�Q\��N���%�k�}e����+�Ď��K�����)���;fn�k=�9&0=��?��(��m;g��� ����q������Ғ��P�A��]�;�=�a >��C0f���e={)~n�j&o_�=ຄaI�����G���O<����i�1�Z��*礃�R2�������Ç.��	�w�]���C�~���6����m�'�ɬF֌ps'��ĉﳩcX�%�+"��!b�l�*��G@_�v&��ϩ�$�o�=�T��3�-��NC��G
3"�Dŵ����#��(6J���9��4���*����
h-[��݁�Ҕ��	?���B���o'KwC2m�pC_�ޚ������Iσb
H��Ǔ����y��ɢ����
����b��������IQ���C���������w�Y�'ŽW� �_�4�'P�م%"��a襠	��.3���D\�;�� [QHJf�� �Lj�s�S����f�Әת&��������b�j=�5D�nޞ������r����}�i9�L��3d)vxږS�F�7�cf�!67����g����d�cOK? !����z���Q�^΀mI�S���n�l4�v)v��{Z�	�	�׼䢏Fƍ<�\~#�bT�o8����Ⱦ��2��x�~0	*�PʯJȀ�����od���f���zS�����ڷ�
��f��L]SH��?��$��'����2b>~�D�ᡏ�������f��p�~���Ͳ>9�X7�6	�o�S�̰fei6)NC�`]W�5PG��/�*�_5��'��w�<�&S��5e��$֎=v���L��Lj���:�����?������A'3�N����@֎��L�S�A�qe��c5ʐ�Z��i|�B|l�jWq�&]�^u�L[�cvGy�*ބE��Ԏ>tr�k�5A�2�cf[�n�"��$lȣ�'u�oB�w�qg"6����äFK�!�GYtW'^`'2/�6fj�A҆����q-��]D� f4}�q"��ָ�g�S�C���� կ�A���p�.�iL|N�L�����u��~I+,H�I�������5�cf\+eb�q�Ry�i��)z�mU�~��������P��ry:I-�Ϻ=n��F�M+w�o2��x��5��]t���]�n�@�?��{���͊���"�c��Ʀ�����^m��^��x�?���;�r�ɖ^�#���e��0~�����4��i�x�R�E���'�_�	�i�y߫��2Cl!���+m�u*�<�N�0���U-�+���9qddHo����`�򺝓A�r�M`5����7��:�}�{b�hMJ��+8���N�k�c�_H'CB��C��u�ĭ��߫�j�T�2jlk���6|���_yt������ĉ�<M����"U�xn惹����[κ��d�k�Ig�y{F�@NoP`�x]K
���et�=��y��ެ����Bd�,WM�	+D\4K�H� y��c�{�M�Ft,|8���y��7��1d|�l:��}ǟ9�cs����	����%�:�����~Ō���~p=0Q�w��}Ѕ�;���s��0����b��xu�F9��DS�04������1W���XL����`�,
��pAd��5�j��>�<�q��h��I8�!D	KP�L��<�]I'��n)v����>֐q^�>��r̪� ����v]O�@I�˗����-��yT������c*����)����Z���zƛ$�c}�A�&����6����Kݍ�$E�"ke���k�'ܻ�ς�A�1���%|�{\�����d5�aW�Ql�L���ȁ{[N��q�0��T /{�؄ډJ��{I�Ac��x߸Hc-�>d�S�b�:t�X���Q�R�h�`Z��+�xZ��;�w� ��s�K|���٩_7���M�K��fbG���$��%Zכ�WH���y�yC?Jb]>��ǩ|fp�N�0��g�N��{И6�J�EΙ0������6��
f�����3�#U4���Ej��%I5�I��I�zC�g����b<͆ґ����i5�����
no�'4nt�I�#��c��n���q���΋��~xJ1���Fc^.�>�@Ut����-�K�n��Ls��?��u�Yl8-KfBf�C���	��)�:���F:0�jCK��/8�[n��*��5�b�Jm��߻�9q�+��d�d�4'
�d�s_�i���?��жu�}�P{�̫������:�R�9�$gu������|�T�u�7��"��)����ڵ����]�8���p]9u�:��x��)�[�Mb����j�9>z}�?���3ړc��Ì��#m�<;���A?�]�5��Q?1nJ7E�L�֬!Y3�;������p��}�TcfC�q�M�k>у��\<l�-�p�b6��S�pn��I	rI��C6~lm�p3��w����۵|{el�w���y�	Z�������&����z� 
b�hA��Zv%��x�'��1��g߮�'�5�������&�G�`]x��z�U@Θ@/CF��&�d�17/N/20a=�y�������5��i8���%��m�=�t�6��І�դ�s�g�'V��۔ٶ���;P�S�۠8m�?<g�?������,L��Sa�/(��0{*�4��9����o٬�5�6ܸ�����[y=�u�/j����e)R�����+�MP�nh �e�t��Z&M�2 <��gwZ#/�9��?�#{�"�g�V�f6Ec?�����>� �h�������s1�t7TW��IHh��
A��E�Ǎ&+��$�;ޜT-l�p��O��̮�d���_��P�I���~q���n/ӅA��$ͷ�.� KzΝ.:A�mI}B3� J��FI��%KMs={����H�`8g����06r���'������K\�~��r��.X�S���z1���{Z�y�3�"*��}�J����*�N�P)�/��pRИ��n�����`ia���������"Rג�ݺ�(�{�� �Ƞ��d�嬿�R�����#������,)�K�fڟ��z=6���'��x�_�H?��D��� ���9sN#(�q7q�)P��R�j���r�t�l#6��
��?�ic�Sv�����F>��A�����<����O9.Ǡ8�Ğ�q/<D�F���1Մ��f�x=��Y��c�_̑H�8�p��L��VY{1S`���0���׿.?���HV>���]�����O���]���(B�P8���t/R���|}Oyp��߱S�5��e�jReݨ@q���5Pq����J����M�F��C�U|�?����͎^Yi*����k~'$X�Y���U��b�sl��=�;nйf�����b���h�Ah�E�	;��p�7�4��M��G~�_�����-:���Mo�1"�σxy�!�)c�����Ft:z��R��	W�K���M���}�LÞ��̓Iu�P����ӲMe��V,!�I㊙���f���l��#�]�NFI�\ܼ*Y�]_n��؉�z8��4W���M�-��im��uQ�px��1[�0;d�شl�<�o��J��]��ON�8�� �vC9rc23l���<ظv��[��a�G��*�`���vbִW��cx\��������&N���s4x;�Hǆ�E�����Ԯ�a��*����N��~O�t���3��UFZ�jkg��RHc��%��`b���T�E�"(����ep��z	*�|X�0�>��ϸK��?��2A�4�!�a�/5�~9�~J�+��1�~���UJj��/g�&�	�F=�(�s���tw'�0+��ԉ���7�f�],rl�ʸ)C��/�����l�s�[��c_3N�K�(Ȁ~��#79�s�+�և�e�b�"����73k����të��7�1�U�˚U��J)���$���ުcn��Gx����ļ��z����v�0�y,�g
M���.𙱴N�qQY{+l�@�G���oF��]�� +d�`��3�Y�f���g�;�˘�e��Aj�����>��ݦa�V� ���ӣ�蝘(sZF����c�)�}���� j�y�5T *�;av�}�]���� �u�&�Yt�cTJ4�O ��(�V���{/F0Y(]�k����4=ŵ(�):�����JY��{~�쇅P۲���˗q���!�Հ.:X*�M��7�|ݾ�&ҫ�^����(ZwJ*�u}�O���փo�O���f,/u6��X$
8�^��:֓μ����y�t]���oS�l
u#U��?���7�ѫud��ε1�E��,0�&R��q+�#�"=ǅ��=;�kw���釬'8}@{������
��7��;n^/&��Hy2KW�Ɩ���J{�����coϔ��po2��WGx<�����υf���R�\O'Y�.:�<R��y
�	��-7Gfpb08�GP�Y�~Fl^7��G�"�i�fT4��U��x�Z��aҼ�sc�SHS�r�(�s:��l���ٱ3�Td
�y��aFRt]B�+�T�6ҩ�B��J��7�,�7bH��n]XO�@�{��5U�9���"v�em؂��B�Q�i,��*��	��2�R��>�h'1z�dvMҁ����S��w�H�����q�pH�v����σ���ˬ3 ����!��n�:�ヽ�7�~~�s��t"`~NU_��T/=E ��]���+��&=�Cŧ��<u��v�71��+"vm��j6�f���K�q�y,�,�I�7g�i�ZJ��+�Ĳ��m\���r���'��G���s����|>�1�l�(/�,7?��#��|[�[�	G$���j��"�ۦ�dqy:�"��yM���{Q����x�w��則�F(aK-u.�؎.��1���� �t����V!R��.�WP�G�����������y�1Y��Ae���PnE0צ̌tK�kRC��j�z�T=���2���7����yv��*��W4�Oq�D�Ce3�fM|dc{�j����ml����^�U&���;��9�|7�T������=���ZA���G����L���2�_�m����w��"�{~UV�
d}/;���tN*?�c��xl�b�x/�9�7���P�8X�ܠ�}���	� ��{����3�-Zf�c��N2�mzf<>����C�AX�C�N>�:�g<��}PU��w�ƞA�����?M���@���]��Ȧ����� �K���'>?D5O5��O�a$���E���?������Q�6�6������8ii�p���ό���$����s�3�JwO`ye:�P�e�V����c����RHPZN� X���4Q�������uRf?�N4m����$���2ȃ�O'O�4�b��%�g�
H��{2G�(3�E4�QM8&�v�,{�����"�&�E���ڲ�V�k0>܍�.�.7&���mO�c��Y�R(�KA{�mG��3�Ci>G5Y�%a�j�5c),j`�]���}�>�7�,0��>���~=��o�`��
?p��cl��b�l�����,�v�H{s���t%���ٜ.�����%:�/��B���/8�h��8�wn���Mv�r��'%1� ���4�&i�b�H�#�z<����dD7s,0���Su'C�9\�񲗪���>���� '�"��>*�8�!hI�A�%�����(tJD�Z����U�����^��g��s���(kW���ݺ�;�������3K��fw�I�es��1B7�=�aSrv<��A�;+��A6�)�CU�+������7k�p�yo�@�:9�ce�C8�[���~~~�:NU����G#*Ǧ�r8��>�⼪<�l�S6�↊N2,��2 ��f�1�r��<��$�9�S4�P�,���E�L����su�CTJ������a��NX�g�{4�iJu�i��9�M����H� ��]t����$Í���>�r��Vr�B\�+��f^hփ�^�=�GmBNv�AJ&(��������yv�	A��b��ce����B(����.�i��\x�������Х�PGL-%+�(qO�hm:c,��"�R+�iʪ���h0��
�dѧ�����;H���kr��S┡份�k�.b�R�H�s��!��.0Y�e¾o�:{M[>�G46�̢�=�=˦�؃}s?�=�����1�����FS����z��b��%���
P^�(���*�n�) 9�g���
]=(���{I֞��¦f��9G0��8�e�L8�Kn�kY���t�;�(����O�$��ϯ����"K�1Mģ8��x���e����3|�קQ�aK�K	]קYt���i-5�Y\ü��/mo�%ɑ$��G]@����!�-g������a�4n�*���X5��z�o7��BWeFx���������s�[��*P���^clO���
#��3�e.���$�[��1�U��<7��wZF$�i�����s��B͉�x�(�E�R%��2x>�ª��������$��k�R��:xѯSPO���EĜ�dY�V`E�C)+j��WI�y�':텣��M]rf�b����!o�$��_��2j��b�x�k�](]�NC�=�^԰�f�=+�(��@	�� ������ |��±lbj�s?�h6
�q���6�	-=	�e�N;��H\<��sS5��$6T5a�Ƞ��Nec���`�H�mܵi�H�C��N�� �l��Bo%`$Y�������������`��5���ϱ|zlbZfpCQ�i!u�EF m�o7
A뫯�7�~�6,�(���4M,�/cQԾ�xl�'u߽;F�og��n�Rd�AM��ei�k'ꮌ��;+P�<�
Q�|3�Q�y��i�T�~,�K#^y,��w�5i�^+A6+6 ���0���D�T@�e�{��Y���Z�����4Q'�}8�5mf�b���$w��
W�LEL@���}��V�ؘ"�����q�(SO�ȘIQ��@�n�x�Q�#����m�q=�F��
�v�4=oə/GT��6�����/,��r$	>�(ψ=��_?���h�� �A� ��W_�����,����C�V��@gB��1�ĳF��0�:�d��z!����P��o�f#��Y���R0��l�`������ɵ�&�m�E@9�� {	<ԃb��<Hf���u��Ҥ�	6L�K�{&A����Hܹ�R'.�qդ���))���m6�i�^~n�L�Σ��r`P�I�]d�V:�)����h��%}ǩ�`y�xn�gk���̱��#p~�����߾����6�$<���"����t�
*lh;�i�2�m�b��z��K?��w9�����r��_�Fy�����+��߾��0�B(?�r��0�qʖ�C��{��ٮ����g�)����q��I�'A&��B�:�]]�D��ҽ�����>(��D����G���5w��Ð��N���b�"	'�*����O���YoNl���G���>)P9C���ޔ��u&���]X7�	��*�t9�4X�n��/&�~����/|<�R�����"��k.f4m��N?Cs�ۀ`p�[js��\���ƴS�٬��$մ��RT�Q�P��q�!㎲~|�2��l�@��f�H�=d��Hn*�Pۚj�%���^�ЀQ�T���C@{9��!�0�<[/�Q�WQ�!��_�`�F ��]���e�
֘��f�=C��;][z9(��Ǎ���bŉ&�gw��Ͻzyn��*N@����:����x{vqF�a�Xl��V�=O�<Z�>.ґ{��(f&��W�H��6�~�>�#H�?|���[����_b�=`:���c�f̀z�E����z�˱j��g�yMk9?l����&�I&8`:c�w��F�(��X����l��bs�;�#�����l�m*K��w{mJ,�q=�y\Jg�,�p���}�Ld�fJ�Y{V=����4N'2j��� ������Έ�yhF�y���X�̀ץғ�J�<�e
�iL�m�<@��x����3��5�}���yx��8i�W���X��kς�N���Y��áʺY�������^���7����^�{�V��ƻ��$t��xS����Z��RQ�w{K�P��r�Jχ��bܧ�ѱ�����!Uy�6��#�1����E�n��,qlT<䛕��I1��L����r,��<1l�뛄���|��z�ƛ�����.&Nc�P.[�DF:*#����]����ﾓ�{R7{�	��,��!Q �'w>#/�����9�}H���?k��c#��F���������n��׿2C92����E�.2J�u�BN�4 �u��ʦ-�A��tp{w[��Ue�v��C��R�O�U'	!FlXa����^3�K�V? �B�F���E5 �[�aVm��'|��[�Mg�9�K[|�_|�(�dҺ�Oy�.��q`L:��+0�a��<�k���ӟ�k�ￋg^���8���l|���E4T��|��j�@��eUPj�:��z/l�n��9���v�x��X���%��5|��;+������������%��A�XO�7T��Wg�\6��d��5��{|�*CG��
� |����u�q`�3 ��Ž����z:�`���@l���z0�i��V�4�d���.�h&l�©[orl�3f��t[8�7�x�W�l u��
��h�T k�i~rH��I���y��DX���N$:FL��e|y��?1K�)�����v��^�pЄ���t�I=F�yL�
۞E���f�s�p��v?a �����������E�U�9%�~�l�����m�X�R<i;a�{U#��x�; 1X��[Da,�U'��b��*�rF=�a�}{i��B��D����*�^�e�Q�8n\�Q,�;�Ԝ�Ⱥ�sނ;�∺����#(a�%
��:�˼$_��Ui�F��wӚδ�e,�b�Y�o)���/�U0X������4q$��a�I˕I�fB�S�
ĵ��S�ߖ��t��"�]�;
�=�^�Qdh]<,+���Lx{��fa�b��2)tӐp@���_��yVmAPu=��.�,�t�~���=�����,��i�T�[�O��'BR���T�r�|��k��8	�� ٭ȸ�I��'k�,�"���:7���Y���,��'���t�R2FC?����Ć��hb�5�q����C���Q�MN(��^̄q2�b:�J�^��=�u+����:�8Q���qt�c���di+V�x!�I��}d�8���pJ3�l�4M)��������Zό�)~���Ked-���&��s��R�%��T^.P�W\�����"�R5��e���-����t�"Zp[��L�i�=��[Sy6����ZF��u����DB���0��|��C���Zl�&���L��?�#[�鬑%/^+�7�3�~���pJ��0�wI��GzD6�$ӍIc� L�̽��62�4曦@mK�FJ#�������of5F��W���޾�Hy�� �7Ym��{�,�{vH���j?�!�.8���/�|�ow#�\#�_)��.�Yb2��$}��l#*�`BL�J=��لrR�I���!�K[�2�|)�hv�������UȏC��U,1W{�6���������D�$~�(gwi�J�u=vzG���κ��a|�@����GT������b��Cq2Yrƍ� ���$G~�d\4vv����q-������|�X���nh:@����+H�Cl�3l��<�rn˼*|r���������M�و�
YFf��!�M2��S�\��&ס�L�eO�rpw��b�lE��TtO�˒� *p�����~�g��w�E�A�^6z갻�剘)!����ݝޫn��}|<�fюI'4gm;��NVb�6���xֽ�`T���f�^2�j]ྛ~�^A��z�R[���*��@IH
A�>�R��f䴈PSi�Zha2��H$��1&[�5`!�<�i<�b;��Nr��W����k�e�X9��H���y��T�������Źew�Q�i�3c�$Hͦ�@i*\S���43M���f�WA�E�y�|����aT��e/G���ₙcY[���$'F4JE�r�E�� ��䚑��Q
�D�.���ӘW4*����|�M��G�W9K��*�ӹQ��Ԍ�i��,�9�Å
��X?��ctd�	�������j�6��Dq�<�.&�6m�Aq	���N]m��ً�S�@S�[�\��o���[�̬�X�!����ُ�\���
^$P�X���I30���$΋�@|^��_� �y8�q����gqρ��+��r2�qm�t#J̾�No�jH^&~��v�lǇuT[�Wu�kgE������6���1�����nHo��)۬�t:Qm��OT���!f+x���b*�Mœ9�Q�3�[5����Tw�7�/���Z��JJcG��b�9�qh�k�PPT�:����28yև�^�m�I�33P���r�٧��R2R��9E�3�L���Nh�.+�v.�K'�m�T�}�f�L(6g;V���}r_�Jg|��;��J�(�҅��M�/���:'`r�;��o,f�fp4/4R@�D�e�#�
���ݖ�qq�w��1�$��R�i�H�Ji@�Gf?�����l�sI�R�=gY�FE����d���X;.��Ǣ��b˰����2�1ć�C�lCeYO�1?�k��m�ב�"�ޠ���w�\c���ƥo�mf�8p�3c��D�+��d�ēRMr��Y"P"S�ӟ���˿�Kd��m���.O�.D�&�=N�%�#>�ς�NX�af]��⾓4?&�j�[��@����C4v.9n��f� �0M��z��{�m�aJ͊�~�f�FجĨ���tO��Q�k��4O�(�����){�F��<��;g��sv��	�'fJq@��P�JF_� ��oD��NA��KN��!ݲpݞ�6���uY	Ն�N�������2�.�ͯ����Z�M݀.�k߻�gb��NknJ��`[����Mۖ~�_��e)?�t�T�ҡ1�����ڽ����kx	�*}ee�l�󘭢�*nD�GH;��޿��D9�nJ�%i�^����I���3��,��@����+��3o?OW�}j��O9,KC��S�L��96�KJ���Jn�Y���xA/|D!����FfQ7��h���SH?F��I��H�(1�j+�q/̑�E�vaI�qNp���m���Ds�h��pH��I����n��_�5,�br���=:�RY�f��C&�r��.������ ��H���%j	w��aAVɜFɸoab�N�o��L�7{q_� *�B��24�jC�Mr}�lA�Rs.�/_c�ف��[4�1��CL�4͹v�j�yW=��gc%�V-S��ZP�8@LHf@��{�u̺��;���I���%�nfB���y����Gp��+xw�3d��{���%��+^sf&�R��oT?�ҥ/��Wa�q>-���0Y�,�##uB]�ir��]��3*�����4���ë>�8� �|M�2��� q�4m 9��_*<ћ���m���UI�j�s�s�+#5-L���8�d�MbHX��[���"�1��/��es�5N��<+96� M2wpF��-4։^�N�+f:]��a-�4�6z��z�@Kd�������������K����W�J
N��=7є�M�y=�T�՜��>���d�m�7�(W`}�������xV ���P�<����w�4M�tHCeu[y0p��R�H���0&DA����k9@���9�N�e�@CF����J\Qz%o�LW�w���ްm��Ѡk?����e�z7�2) F�&�C�� �5�']T��V���&���IH҅vW������T Պ�倸�����%�k���!_�J���_|)��C<7T !�>rM��%�^�c42��|M4��8� ��<�#�1ӗ�@�r����x*���� tVYǸ^�3͈��"���Wd����3!�JJפ���������*���(H�r�����e����n#kG��7� �W+N΢��I=[}�����M4t�Mn,���v��w�������S/p�PoL��.��3x���:�F�V`Ҳ�42�$b�g�pa-�%7�f1T$xQ�ص���7L���� �cVxש��9I�M��ߏ��[@=ׁTʝ�$�/�d�xϿ��/������őƏٔ�Fu 3���@���SaXn�ҀƎU�E�/��s̉��Uކ�2,ݶ����g��#G��ݣ$�V9�:���ζ7��}�2oպn����A�e\Ot�qH��"x݋PV�͊=�z�gB���%2�+Ǧ�tWդu���̎#�G�i�(>�h;1q��Y~�e<�A����|X�C��D6I����_��w]�Xz�걼_ġ�Mz�l�y_LMv�eyv���x*3��b�cmWUn�&��q��V����v�U�;�kd��>� ��T��Q�������Sڹ�h���LS`�;��J��)����.�Η꿥��א*l����ԫ��>N#Л����=��z����gƍ�f�n���S��7?m%�c�z�$�ԝ�&��(E	dc="�~|`�?��u&��� |�]�_c����TL�X8X�p��R8!m��ak���Y��P��X`PK=�i?�Q������`D5��;�\�H����(^��#o������l�n��/i����+g \���iRb�L8�'^��ɍ1\K41�m�h�^ [��*��48^���C��9�E�� d/ �= ����(l;3�rmωi2�Sz1<>=�&$���\Q)�hޑ�iB:�?�<KV3>���uJLv�n��(�a�̭�����D<&֋�x9��&�R6eO��BvyxN(G	{0�8���(�O+�h.q�5_���d�ltbo��E�t�\f�i�zn&YYׁC�s҆y���FO�v����wU�0%���s�rh�ݤ�v�'�6+�o�wLI��)�eR�E����B�mRƚ.�&h�[.�ϱp�f��l�P(h2�g��y�DBw�t����ܝ���t��άH����Ԛ��`�a�����)Xp���4�">�C?)�]W0�QC�p���%�&)����q̬�e�4�-+2�t�r^i�pT��fe���Yphs�h=��v��$wR��o�J=�)���햍"F`s�<�n���'kʣ��d����
�U3����A�F�A+�B�0�F��lm'Cq@�s����ʃ�MfǨ ß�͙�sֆ_ �}�"�ДLO���r�����1ߩ��h��j�2ˣU7m�b����n�[������P��4�V=a���̊3;��2������i�pJ.��S�
m��'ǐ,�)ް��Y~���;枳�O���V�v����m(c��!Kg�fk�Yp@�EK����*���7����wS�S���П��1C@�8����`���1@[:T%�Y�ˆs.��	3#��8����97�OxS�U�3�wJ�J/�2��KN����.5G��('F���z�'m&�g������\�<7���68�Ҋ���>2��T:�'u;#�u�F)�y���0�X����"�D*�kh�=Y�%$0��&A�뮨GyL��Sc��r�(Z�$��@��}f`��̴� �4pZ5n.9\�^�? `�ؠ��"f�>>�������2q��������X-�5�1����~U�7~��%�k���jp[6�i`rQC�n���slXVFR��EIKD��Y�3��N��qO�%;�k���|WF�D6׀5PH�0�6���/6H>s?{F�K}�{�v��Z�e~���w.�B�w�RPPs4ɜ U���M��koa)͹Y�|��59��Y??�ǌ�;d�]6�@S��,J�J�>U�������r�m�`�KF�R�&�K�3g'![cP����S�����?c���tb7�K��S.��Q�Y�62���4��c�1~�H�X�m[H�{M��E؉�_c�X�6�����<�5n#�nU��̥�G��8]^zzfdx�0E^9���3	�����玁'�I�*�!切���;O�8P
aL�9�����s�2̂��X�-�Q������D���� �88�02x�ψL�R�M���:Kj���`��[L4�����Q��q�q�Y.�|��:$��|uô|{#� ��Ө	+L����ಪbj�Ͼ�l)�:]8(�����4	quHx��Q	M���A沖��]Q3����\�A��?��;%8����\��:Q*%?��%��@���E�t��K6��k���DcpV���[�r�+�V�d��{kM����Ep����p��G�ԕG�j�)�֯� [J���7yA�a1�~�@�`j3| ��	T+�����N�,+yZ���2��Ix��z<����6q|�����ȑ�ƹ��pG.S{=�B�m����`锞�)�<z͓?As]D���he����"��w)_{N��� �I�[�1�qd�n9}��� �gc�jE!qY���(c��N� ��-4|Oݣd��7#�n��g@�q�Q�4�=��d��>X����|`^�.�q끁r��f�\�͉�svs�U6G.t�w���W�o9r^���"[%�=CWi���w�=�0�FM��#���^��$��K� /�B���m*��������6��4�1_zH!��.�_~�eN���8d�us���,���,JIn_�Q��T���#����g��G�_������;b��cjH[V<
��.wͫ��f����\���E�&fZ=+x��6��+OˋL���Ձ4Ae�*���ɂ�ê8�q�:��-����N���^8��Ŗ+2m��)��ۣ!����Ҹ.�EZh��Q+>�5�5u�]}g,(&�T���1�?��!�� ��8T�l��u�m����*l����Y?�M�،����K�8*��נ<0��X��ٚ�m,�'��Xg����%��{w�?~|l�_�}X]��añ������a� 4�(���q�����ǟ�xp��Sf��.Ql����d?ٰ���_g�沺J�N��>U��n�%~�'9[a�̼��SJ�s���no���(q�-����F����.l�ĝ�/����s�)3�h���З�����J�$���9G�3fb�����Ҍag	G,��]w�t��bmc���0L��X�bu�iT�lx��4�ȴ�ݴ�����I������W_4�)����)��~��.pX��x{m�}6$�R���	�iҫ��t㰩����7&�<�F�}x W���
��]���v�|�)�c�+3G �%��7��г�C:����@�,iȌ�;�/��t׍eH9,�jsT�ms�Р��K�,���[�}���
&o�N]�y;)���o�=��+��t�i�̨m��[ß�a�z����{�V�lxJ,i4���g&�Ɗ3�e��V}Fv�R�6}Rsa!�/�7*ooڰ��Ȫ�`np/�$�cr��|���>e��M�e�� �*����܀<�\c���3����a��������Į,�F� �؟bM�x����י`���q��
@��Ph:����և��u	��z��q_�6y��&*5�rT�%����ͻ�-c~���wKc��ujI��ޟ��;�K�{�-�%4���`�/�M�b _�p����՞t%ܑ}Y��=)�w�ްq�>�u��EXm���l�:�������,e�(2P�z^$;�O�p��(�t�4��q#�����N���p��&�����>FT�4��|Q���j��P�M�sc�����1�1�"�M�moZ{�DK�}_�ї*�7�>T��+�eSloQ׵����B�97��z�a�@=�{���mT�س�NZ�����ѯW�s( &0CU����&��-���8n��0�o�,\�䱰ەl�[��`�S��R9�Ҽ���|�j�͍��f�sSSB��vr%��nJ����5{���~W�{ˮ36�4Wt���i�lx��A���������g������Zw�(s��T�:Q���1�ʠD�����i'8����l1i_�/��,���j&�!��|#9��5�ak���*Yn[�)Z��֓�x� �	�M4��'A{s��C$��_�^��=�S�%��Զ�RhC�������ld	n�(;D �2R���r�6���	�f���DB#�����`؊	q������4.8Ci��ҐX�uĀq��wl�7����RT�_����GfT�������P�)��kz٠���C�s�y�|��R�_��;=R�{%��6�uƀ�/������+��`�1K�����Gm��{�L<s��:�{�DV1�3Ͱm��f�"�dT,���22Wx��kUҽ|#k�@�á�%B��A9gn�
[,
-X�1�'#� >���u_�70Py��D~�R��8>�,�X��.���0�d��m���-�$�>aR.�C�Te�ӳ:��8]� �:�%��<�>�}7�J��͈0�ޔ&sm}�D}S,$q�M�2��C�A��}��2���|PvU�j���&3P|1#�l��(���ܼ����<�������]J�J�Ru���L7�C����b�:Z��~
 ͓�ޏp}�����Fu|an���x������@�.�up����1�~ l�:6ö�!��0�0~c�"GZ�Tj�U&5�pJ��涌��i�B]�D6:�`��N���q��_2�H[��?{���-�󂾗��L�삞����O��cÍO�\�Ӑ�52Ͽ�}`y��ϐ��<?W�0���(��}YqOCࠒ7�ޗ8p@c�2P�p�����ͻ���D�S!|����p��qzo�d�nS5<'O��z��D �O�/�M確��&�~��b!vWv������5�1R��{̸��{=(3��(8��?Sz,a����+������>j�wK2yΠ>$��1*��:�����Z��'{�:ؔy\�+��;�����jLm5�[e{-�d�.��u2D�}tW���ܧb����Y}���r��y�&�4M9��%���[��
�j0�������b�n���ԙ�L�0rs	/b�,��б(��`� ۴ 8Acc���p^��ƫp.J��W��
͊�R�M�a��AϽ�A��G�뉛��B�F���,_���u�����L56�v-�N���-�4�<4���{��,�sS��:��)��0��e)2��� ˒2TK��9p�M�q�҅G��>>�K� $���P<��y��2ݗE���E��!���D7ő_���2��܈'q\a�;�^��93�������Vٜ�d��
���>��XT|�������[�-˳�A1�(���r�6¬#���TLpxcnf��Ţ1"8,�o���b%ם<)&��;)�)o���=�zu"��d�{9��Zk8�U]�GK�F6�j��(��WY&�R�Ӆ�Y,˹�8�u�s��徃�C��޴R������ٓ��(�d�kS�&:��lBf���_5e�������'���2�Ln��F*L9k�	X�(#�,��ǌ�v���ƬZ��,~�4�8������F���$wbww��>Ǉ\J�	���=0By��)�m7���#��걳P̓�u� �W ���5���a1�����*��Ә؛ڭ��M]2�L��Ӷ ���:��^�.�<� �N/7>7��l̋ڦ�A��4Gw��@�86uOef5yѮ��0�f���C2,�C��+0���߯g'Y���n��"Sb��#����d����5���ϨƦqMlh^30<�A�>p���X�1��FlPC`�"*3;5z�>mL\��)=u}�v�i��㙙�@��!�_#o^�r�4"�/�41�纕�{��` ��BL�f�7�^���U�YU�]��A}�ϰID���䁽�SB�u�9�nNA�iz�R��:����L��06=	�ROO;�@�	��%}�?���A<c�91�zo��e4E����5%SmMm����H�ԚGF��8�"+@ E���	�p����O,��������_8��&=�}}��ߒ-}�x������6�^���0Ͻ��fm�7�-��F���$�_M�5�]nv�ƽ�=Q�ƍn��i�\`[�7�h��1�d����?���m,k2�*w�Ѭؑ/Y4J/N�8;����8���_ŵ9#9�M\��ک���;ós���!g�tS�f]S��r� �����ր���Cʺ,� :�\�dM\ {��'��(������?���x�~�1~�� �V̆ɚOWј���>W���H,81���3c2�׸�ڷ7t#��6G�)4%52�b]���R�nu��X��3�1�X�?�+�6f��,y�3z���=����F��
�E������N{1,N�bA�@G�g<�Y���GAp���^��p��z���Ax�JE�����U�������|�!�v�c�y��8�XK�0=E������´ƕ]gUΧ9t���+��P���yvٙ6�T����u���%VL�~&N�(���H�ǆ�/N*yZѽ��C;��RWd���r���NI���1��E/������'g��ˉd��X9����4	����4-[�a����z'�Y���:��e�ъ�]5�JJ�]~L�k� �!�]���m�Nnȵ��M�t�r�i�~#`i���A��bq8e/|>�)i�U�&ԃ}L�->_�͵�T��J�'|Q�J�a��,(X��MX�}�k�4��ڰ�^�Td�;gI��n����T/�M�y,r�e�Y|j��Wj���-$����#Fȇ���_��p�x1���g���{b����~�d��P�lb�i���Yn��]i�n�H��ɺ�7L��$��.N@5Um���&qfS�z�~~Nt||VkR���0
��p <)k�,�"-�T�;6��M���T�1��)��aQ��#�ǌh��):5m&����ߨ����5(�����/�Y�ϛ����s�����A�����Cxo���w���8E��Ą�S�r�Y�]fk[�>ϓ�� L��`nY�*�S�������Ʀ'�Xa�pfԛxp��a�	T���*ɁcE:aeG)����>F.��~�/e+J�[e�&�r��Kq~wr���8f�Nd��������D)��uQ��ܬ9u��v���Pe�3��4�Ep�qo��FCI�`jf+&S���;V�q�T��>/mn3
^���������ʺ�kr�~u��ָ���5�VKf'�UN���,���BZ��X��oOm�)x��!��ao�S�Ϊ�F˖D�[��L<�����2J��4�;�s���98�7����X��TT��FD����U|0��ج	��|����$+�S�eC7�i3����I�7{1kl���xP��I�T$�sJ��9m�񰽖�ּ�O�گ��x��4u�Q����rڞ����Y0X'�pX�ᦛ������b��@�}�}`���؂&"tG�S�f��lY��pI4�.�Kb7�xQ0��J�oH��@̊
R�l�\�'�"�p* �OLM��k�gPF>>>G ��6���t�o޼M�2�~~������M+�nw��]���{��K?<�:�#"�h�[2���;�Yc	�>}-��'� ���_4� ��{`�LIg�^[�%`݅	�=9���98āՐbi,)�Q67�3e�y
����"�{�����R<2� j�b6P�T�é;%f��n�d��F�d�T�\�}�ad�^�i�����.����UY���&�|AәŪ�L�1�t��o������Q>M��r���I٨������PJG����!i�3Gw��!�S���kAL�i%*q5P'gnBN�ԊK��Wq`������3���m�at)��|]��� J�X��nڼ����.UinP/�y(qJ���nt[Gp�i���h��,{>�a��}�9�T�0�d0�9~ߘ�%t�B&�ō����`�E��)�~Y8�� x.~3���5y�y�9�|x6fYȓ�c�%o��ˢ<����?��|�Aux�g'���)J�Yۆy&y4�@0�TJ�����{�9@�,��Feea�f$�R��ᛵd��V	�1C2!,C佚��{�n*��mw��ù��g	�$�������([�!�X��9�-��kڙ�i��51��oZ̝e���g����gLh�8��E��c�,�ָ��4B�y��tU:e6��tj��A05�c^4�`
Y蹂]w��P��%��x�$z�%��巌��y���DP�l��Pr�0�=�J_F�d@Ul5Q\Vb����,6���1^sQ��:�����A���eucp5l���iu̓���H�oZ���<�H�ba1v� >?��F�w�)���%� ��C��h�ݦ���>���]�H��)_����=b�&Jh^�I1j�a
��'�N�o��~j<�&��ܯN��4��h�=~�p�8�<��?�1L=�Y�a#8�,�;���y���]wײ���I%�����^��D�iZ+���H��I�.�M*\�(�=ӕ��3��Z{*���.����ŴLX>�
�,	�2���	��EdPZr�k0��� ��:n�MZ�������au������1�n�{%��w��<��{i��d.�3��`J�V�gѦ*'�_U/m�\�yT������R˹��]��πR
 nץdf��W�L�W��3���)��7�:j�GT[��B\۪_p��ppHu耯ej�ِ���⩮\P��7k�1��� w@s�H쬷mϴ��4��]36� 2�@>CH��Q�y ]��"6��;��m������:!��Q8]�KEO�Dn�M�d�Gv�Tq2���a��"c܂��0#q �pG?���6*ֳ,�z�:X������������K�����N� �i5tش& ���d���aP0�,�&%��\�Ў�/6>(�����j��┼�F��7�X����G��O?�������ⱽ}�/�z\�>(�ѥ�����A��%�~�̂"�+����G(?j|G,�˰��#�/� �>+d_fk�P��������)j2��r0y���<>>�̚���U��i%�~O���C��!'�YY�	���s~�o�Pז15I�V�_gY��d>�$a�9�]�'�,,�u���S;���A֒.�|EYT���D��9J�k��Or��V8A\���E�/�st�=�k�;��=g��f�i�-wrXZ�����3x��eBc��c&H|���A��@�З�wa����Nji2���^
�1�CH��"=���h"�s�̋�>��
�w �h�������xsQ��}�>)�@���cD�qB����~<�g�
Q�	K���x~���ũ����nB`�D �F��ہ�!��"���y�5-=��׎����������Ο~"��2ԛ�U�+g�}���q�=�o#�n��<�n��|�IG���ȝ�-�e��o�&��}��7�Ձ� ��$[6\�R���2�&�fTW5r�?g��y����sVW}�3R�0�T�y�l�cd��0�e,Ψ��5��M.OJ�N&0I��̣R��B��G�\d�,�=+9N�k�P��N\�6�[1Ľ��� ��o����$Nko��*�2~�TA.�w�t�Wȴ�Xq���&�v�z&N�C�I{���)�ؤ��wf׬�� ��:�RY���N�꽫��T�2��⻚/��U_M>�%�+Dg���Vu���49#� �:#-1��LF�@ڔ����
ݎ��БG�T�ߍ-����VG���B/�ޙCKG�_?b+U|1�n��F���W�X��$!I���J�b������u������x��aC�}�۝�1L�0`�$��pP8fX�vYo%+��D]��,�?�d���J�5^������Q�"��Bڭ���H佨b��'m�/�S��3�< ���/��N�/ۆ����,Ɠ֤��|�1)[x&����5%'���������+g��(K�u"��F�q��5���|Nbd � g�Ee$��;��im����̦*���D+;��E$���l#��y���I/2���D���hn.A��9��ZΑ��]��9�YI��x?ާ�m�*�y����m���'fK	fיJ��=:��r#C��!7D��}G�*3�i��w܃�T�1��s�#ڶ�/��U�����zN�I
�?ǽW�|.���u)�u�n�^� j�>I�0<� �Ĭ��K2< ���I/�u���/��.�#8�)vk|��N�qN��eе
��4s�J���/�
�r�����H}ّ������7���E/����駟�x��<8i�Mß�=��P2���E=�6H����Wo�����n�P�=G����S�O`%�� Es ׎נ��)� #펍������*c4/����F��b�� �Os���ŉ� �v>gC��Y���x&���L��M8��$�A3��Z�� ��H�?oA����;���D������1 ��}0��'���--�>;!�3�E	��t�#P�@	Li_���H��SR����Ħ%�ƦN��=��`�۪��{Ѻ��m��~'���)��,$��1���[y<p�Oߍ�����l�B	��T��n�u���!
�ag����\S��o'd�ϱq���<���^A�G�W�}�5��0g�4<\?�md;�2�^��|�����J����yev<?_q[���^� 21�t휥��o���d)�2��A#�q�$��
�����p �7VQ��&�7H�	�X�%����M���HX�H�h�C�w�2 /
��������Y`Q�K�["�k�{��ft®��JWS�����a����.r1����.6���p�D>���[��D�;��@�׻��n�~7��d��Ɗ>n7�*�, ���ؠ��NGI]P����;L��.]���x���N�q�+�)DzR��\t��^�>,NF�5�0g����(���p�0E��Rk@���I�m���ta��ȥ��ÓuC�����`����[0�@�uT��^dYr���j��ˢ�޷�J�Ms�c��M#Ck��ڀ{�!�?ws8p� �� ߿���7���6���/?��������ݑ�Fl���(���f+���-dk�M!HrNzN��<�x�@p��/�}�|����~O�7]$F6/dN�z���a��@;Ӿc ŚG��s�o���=F���Ҭ���7p�9�9p�4����f�f億��|���~;>ӽ��Q{���{�͟��&l�f+�O�۵D����眢d�1�`]5�'�%�L�FK���}��7��8���@�q��6�b�L��y|d�q�(��5'K��=W�Mq�*b�Re�:�<�	�onL�_���g�l3�L��t�)m��F��̛>"x��lyҖ��iX0,�E�^�X(� ݨ��iO�����?b��|q$�I3~|�t�6jb�KwR��s}8Vc
��)p9�{�.�X-��ԚF�;o�Ԏ3r�����(�E���P�0V�z��yFZO�$��IC(��%��L�cPf�)ʦs �`�й�/�TwUZ�ع��XfyM����u�{�1Ӫ��\0he�(�o�SG��x�z'Ïm0���嶆c愆�l�ز��b���hH���.q�e�rNyl&5c��j�e\G|�ܦ�:2�(�#���!+6���g�X���S�+e,�=+2n���=B�*+�	��!dm|���(Y��fI���LƳ0�N�F�d?멘|֢1g�x�8�&�L����XmIƮ�kM�+�֪,.x�K�h��s���X+}���]?F�����JW��_�is������--�'���%|%�t����_w����B�n�7�yYx�'��^�R݊Bc�.w=;�zk�,O| �Z�T�1�AJ��KĦ�M��4�?+zp��09�6��%\c�vuIղ�x�v�t(DMµ��o�׊����)ʖV��9� ��o�gv��k�tcbv�9��Hd��,���[��������oqx��͙3���@�y:����:� �N2�54����y��V��M�o۹,F�1�]ݥ�S8��,���أgڶ�� ��aHޯ?���־��}�yL:����`>{I`=�q��ro����q/A�3aj�b?*����M"|��_"X�M�G���NH�5���<�zә
���<�Ij@�g�C��#���_a�"���I�׀o���u�ָKޯ�=�>���U��iK>үb΁A�c��,M��5�rI��{;1�@)�1��yl����ۃ$�Or��l��ķ�`�k�Y�wG�%Mmm
VZ��?�G�2��"�^�Ц�Qzh�@��$;b��ֵ��u�� r�b�f�x��ڮK�Q8׬�t�1��q��.�!D��L7%�p�j.[�W��v�q�|6.nD�D��.�%mſ�C��RG��<[׹c�I�\��ÿX:�ylL�/��+�*���&3�V��օ�]����a��Y3�,R���F��N��ۆ#sM�>����U�/AɄ,�ǭĆ��?� �-�Y���f�`��r�՝hHX#�7�=m�I_鰲
-�O�({��b4��3�l�b��(3/���9>�YA�����M�H�'�=�)*#���3z.�E�P�=�2�ԝ����d���:��Z��1�Q��rfFM�7��0a�I�(�T���=�ۚ�I2����k`6B64͞%�5���;�a95�����I���/<�b�{J{���B2�]'��c�b�Pp�'�)�C��(�	fC�f���T/i�����;�g7��^��j��ŋ������T-�I­2��-K�J��XO��,m��=�nyN��>ưm�\��:&�x�,�Zc�������j5]öa�|����/i���?G@���m����5y*K�VB�� ���P�s�J3���A&�k�K�FiEcj�Ņ�(��В9�^�l/��I��69�wH����"�����G6�os�a�>h;e�ͮI�cL˒��x�d��T.�T����{dg�q#[�����?��i��
�"�rh�GC���nnL=���D+�pHI����Nb�ΰ���~Tkm����l�N��xm�*2�ݠ9a]2Gf�0��º�tд�,��/g�O��@�,
g^5��q?q���1>ײ��ʡɔ\h[�uZ?��������hY.�g89� �jÉ��ɋp�sB��uK'6�;ChC�j6�j��2�!���*�z�Y�Ћ_�*#�"�q�4�~'#m���5��?R�Q���n���q�	�M��2(���y� v�悫\�U�)�p�_������^ȸ&s��k[��{)��"a�"�b���!�>��
�qʽ�3O�#O�M��  Q���v�,��@`�:�0y���,�f�9��-���Jn��3E��	���N:`Κk�9=�����ޤr�c|˜�Ix�����Y�̳�"CG�f����	�*��t�7
�t4Q���*?C��� cMT����6�u��A�ʵ���Z��:8�,�!� �� ����/#��J�׀_���	��v�M��k��NW)�y���Q2SNкS�25�-�](�.E)'����T���J�S$��w���pf9'UR��|`�9��N	��қ�Ik�<��'�9��Mr9+ZT��mIJ�߸'�$���s}���A���:}I���@eZWl�LM8j܄U4xk�|�+��$��h�|�{�;ߺ��5m�E�R���w;��A:��u�)�F>7��7Sb>�؁�q/G~݉���1�<�\o�"�ax�S�6�0�ȲbH�a�s��Ϣ�Pl��I��$�"��T�-6M���}p������,�����
���͑��p���>%l:f�_���tN�f��&y^�*��3=-��F�-b���2\n��@RM���OM#�)�|ʶe&��K�θ,5V�HRI��׹a" ^��&mS�x�0�"�~_e���C�t�?Ŵ����j���f�&u������8c�fj����wsS��<��4��7�gl�s��m�� :��9h�om2�Izo�c�1JЅ��A�mmoWfs����5(�YG��X����-K����KBqe����l�Uc����`Z��1���VAx}���z�����?�6�T��%�$W��j�Ӓ�f����(G3�X$�/��9�iu�_ ���P�͑PCIg��B�D��$�o�0Ң�iub�
Oϻ|�,J u��@�a�(#XV�j����s�lx<������.`¶�r�K�_`��2]s�c^37�>�3V�"礟�"�l�fε��ޱ���|�,�c<[��R6��s���]y��E@��_��u��+�#4��bY|�ή���$|tl�ؔ}�U"��o`|�!🃓����n@�y����=w6�H��#]͓9٘f����"���_�mp9)�El7D����*��,�U��(�×a\3y�X����<)#�Y�B<�p�K��^8{dG��,'�d��]4m�B���V�6��4;�[mSd�1��5�"��t�)ẫYMn
{�#x\�y}����J@3���b�����������_�o���Rx� �۴c[���=�&1�>��f�N����"˙��QQt�Nr��g)vm*�Z��w�&~Cn�bYݵ�H�C:;����3~�,��u�ڬ�Уr���%�������~i5hJG8�C��of����jzj9d�2��-���;���V|�S�lR���]r�S��0�����͍��K�YT(jq3�t:$���~�&q��Ab9_,g\R��g+�*�Nh��נ��1<�.M�Xm5�iG�����8�p��+�Qj�x�᫮�<J�������ܗH�g��.���su+iO�h����`�"��if�ߋ-��;����l��ƥ�hx+�c��{�`d3�L ��~l󹄓�4�~�V<�U�H(�m��k�%�l�ϼN�+�BU�nwJz+�U����m6���X?YǱ&Va���!��B�S5�K��~P?��*�����/VϪ��
�i��UÆ�t�Y�T����cP����ܸ�Յ����Ok��MRVa�ȳD�|㬓�%��d��$��;������D��"���[�c��/��=���p= δ#d�m�V��U�Z�~/����yJŗif�0ծ{�Y9'Y�9�����&��<�!殶��v^����P9<�<�i4��RӾ�����	��z��U	۪�߫l7f�/Kf�cG=����P;DӤ�	E�͒�*+b�#6�F�x@b�YS��>r�{Q|V=��R	;n/muh_x�j�b��3 �9���.�b.9$ig�hvSVD������b"��g�-�-�94��ac!ʓ��Sf�f�Օ+L�<���T�4|��?&ō����t�g(&%�C&Y\�i���͉�\�y�OSʭ�@`}a]��+9eYXWwu)��G�^����]:W)�^c��W�����z,�'Y���d������0�Zƌ���>h^������&%�����2�t�yr�F�A�9�ķ;��?4:Ѭ���ǝXnl<�).�.���"0��,-���ŉWFR�዁tH\�Q=��َ'gR�p�&`=z#����I�ڙ�e�ă?f�
�a`Xˬ�F-�P�|��Y�Ɉ +�^��b-jz���C�
U�I�xַ7T���R�z�C�u�Y��^���vi�m2|/��PVm�)�tx\�����6�X�!�M�N�n�:�K��B�!�
֭a.d��5�a�*y�5�:�]���%��9�nI�:~�gfuP$��R*<����ɽLz��>:����w6}��j9	�A�=�
���ʒ=�ص_�N<�4�Q��Q�8���KY.����'�y2�Y�	+���y���a��?�`��R��1�H����ddĜp��+7�.2]� ��W�Vu:yFэd��-u��*BqY�P9.��׵�01���4G�ϟ~��)�<��$q�(s�&�ӓ<I�H!M#o`~��2cf���M%�8�-3���<��(���h�ݽ��Ha�dV�4#mx��)��=�5*�V�iF��F�4�逫�h(q���ҡBd6r�r��.w��+?1֋�幡M���H�%��Y�0���d0�Ф8�>�d����^�^g����\��HY�D%�lR6K���g�Ua}��)�X��I8 ���F�ޞ�>��C�,�1�Y���8м6����cn����.�5<�sg�l@��!v�fH�����ƣ�{M��p�w�s�ؘ��8��v�n"�N���=	�1���(��u���T&P�)|Iθg�a?n���*~�!���U'ALh֝wW;�=�'ko�G�3R��LFZ���H׵�F�(��61-gFy���߸]�w����N��i+��T֮9��1�S����3��KGW��b,�v��\ۈ^Q@�Q�A�|��7GF��R�cH.��X�%)%48�qY4�b�U��1)��%����ʱ�4i �V4�LkuQ����̾>���xg֗�w7�l�|>�$TA�ԉ�����h(�~�:!����@]��MU�A�]��i�^�t.�쯊�������p=�O(�}ݿzhrw��[:��~p�fW��5qQ�bB7�1��P�g�{�p���ϋ�Di��E��ڐ괬��5A��H#�T���Z�Z�h�?Fè����9L\�xM�o�g�����r"�	"���0ݖ�k��Xi8'_T#�y?y�5��v��|�z��`�{J�E!�]i���ԡn���7��@Azl��'�[j��a,��2V���h	���L�烬J���Hݵ��r��t�@�H�f4.M��W�&�]���z��N���7y��&�͛�G�t���.E��kS����Q��:�TSQ-�t`�h$����ȚsF92/J�zZ�����o2h��ذy��3��9"��@�S�Ȇ�D^b�V�pZg�x�Q��|8c���E�YT�#�7?'��C�h�\^󠮳��w_�`�at'y"���# źa����B	�^0>� �?᱊ �V�/r������J�q�8��ZB$mǉ���4f0S@6�p�s�7{A@�j��p�f��w�4ظ~#
/�=�Q��7�����b;Q��wM�~�#h�n��й)��A�~~����43��:�#��%6����g��,��0K>s�ߢ�vDw���'7��m�-��\q�C}��ۦI�ʢ
�6[$�m2P��6,a,��$Ţg��jf�i�����5��~�?}^��ry��PQC�I�ۋl�I��WY�$l������(�(���5|/ܫȿ���UWC����F4����(�'�t�w9L���f&E�$������ѸG�i���� �����EG]��;)5`,�sSc�膇��+#�����И�ؤm��8�CO-&pw<i,&�����9y�,1	���<�
3S��s������?|����C�8�1o��Ls�Q��1�#�:�$�%�mG�����<���k�߾�1�����q�@#nEU9�]	9�"��C	=��l&����^����;�D�����2e52W�}Urj��)3_�!d��u�ּ��ٸ!b�c���z1R&G���<�rݷ5�N���u��3�j�e���9�$^���l�XJ�U{ъ5�xcf�n0�ss��.��\s۵\J3��Ø�<����@�89����m���q�}����z�������#-s.������S��6
�%��.F�y�n�ǡ�瞢dyN*1��2�Y�k���~?���.O�S��`��U�!6[����[@�
1N��_�x�\Nqŉ\��є2hgvΡ��T�s��}�gp�Ol��]���	�/�ɻ�)֘���Y
�4~Xd��/F`c�@��#�w�ϧ���hr,��P��̚��0�ǁ%�NF���ڥ�g�m�J� �~�9F5;$��]��ҥ�WL76��:\p?(�z[�<���6�a{]��Z��Q��j�b7�X�]���5Ny�;���(�L�k�q��E�2����Y�S��8ֽ�z����J.([}�TݔP��"�RᲚ��g0�T|RE����	���@'��|����a��0f%���TS��YE���$��:�4��$�Fت�Q��_QDbC|߾A��m�N|Xd0�h8�l�MǇ���%�K�����kܰ?��@4U�:%��F+M�R�0y��%q���\��?�>�B���V����>�n���1ҏ�=@ևR+��{n�eN܇#ug��paE�)�U(�D��(�?������{�ͽ��6�7�>Sȸ�t�[��!J��?����/��~�Y�8��,ИXzf�?1��S��	(������P�|O�u]��l�x6V��KV5'���
�_Q�1K�f�mbd=bH�3��:��STcy<�߹�U��NIu׾@5Vi.(8��:�R���D21���m�c��T�����T���-Y��<���Z�W��488.�3�|A8׈ς�2Z��\l��B>�!ACZ����r$HV��*ύRq�Y �??۵���w��e������|����ϥy�ল?��.QZ��I�g��.�ܜ�\jM=8�
�ߠ���J}p�Y�E�8��F�x6_�7��<7=��p������
�� �!���A��g�+Ӡ�X����������}�n���Ǳ���ia{�w�Y���_b��z�@�&��f�w��u���<s|��¹�g��
���r�u���!��o��cR+��ѐ ���>�(�n�ϰ*�=�ߕ���~����O�3+W�a���D���լ�!�����L	�1����g�J��>]���wE��k��xFs�Rlr�L�����X��@R|=�y����X�'�\씕�j�fIO�Ľ��1��hj��C����/	�Ovmܳ���tM*���!���?�k�F�,;����KQGէ�6a�j�J$��_'�y�,c���6R�Ikz�9��`�w$�՛X�.2��n$E Ս��Ba�	0W�� ����G�U�zzv���6e�VH���)êo��!3fw��6�RЖs�8���9e�x]g�����=��x���"c@ Ģx��}\�߾��j��F-7~/ot�줢BP����Ok�EA�d�`������
��qEc��C��b"f��ms������8��S�l��A�8����x,�?��?5?��8$0K甍�c�+B�2�Y�S�N�k����jҽM*�TÍUB �zwc�@.�| ��_B�7��_�n��'^}��h:֕�qy}ג/MV�H��akwwl| ��7���g�����YwI5���|��3�T�;�7[u�EW����%S�,F0�.6���c������W��F��~G�aQ�*F0,ĳDe��#�q�G��{�
�P�M&��X4k#���t�5�d��Ȅ����T�����l��2�G�pH+��*y�D�n��pp�H
��+g9�dGv;�O�@I�����C��Tc�i��yCyHFGUx譺w�ZcSgr����r:���X(8�%}knd������75GL����|Y�`T�z�46~X�_BF,�zTm�6Q۷3/*X��0B�bx�4΋(c,�m��,�!��3��[פRF��	ev�ۙv�=�s�����3�ڬ`ڒmj�2<�#�nW|f���Ʃ���y������9@LA=_�3=H�k�g����wYJ�I��.2�.���GY�iD�F^�����>&�`N\�
�*�d��4}/,�� $�1iQc6��<U�*��N�L9r{Q��� �t��v�g� �S�fH��x����� �ٿ�Z��]��@������ � �a�w�A��̛�q�<G妜�I��h�]�Ls� �W�z����� �2�^�A���w�lZI�i����:���u�>��R:�>,�ǐbC|�ݷ�-`�����L���bEF��Rς-�L�Mՙ;whw��Y6�o���8���� �g��� ��mt��f��u`��S�휵�Q�3��=;��� ��1�9cZ<ὐ��0�A��il�G/6��,==���������o���)�KM-㋱��=|9r��*7#�w��V�D�aq�h����2�����ō	��>|fo��vʵ�o�u�2�1u|ſ;�O1�`�ܜ,�8�3?g��lM����7o"Ƿﵫ&߷���\8\��p*0��u���A��ˑ�t��F��_�=r)o33<W���Y�#���K��&�ۦ�����+B�sc�Z3'���r�eʝ!$�3D:��D�����n FQ�!'>H���=�'=k�ׁ_���cNXH+ɮ�l�\ }�w��H�iE�)|��8#�Ƞ�/�axw`]��UY���Ͷ$�S7qcQ�"+�����w�'���`'*9������q��}R�h��!�Nio���ܺ|E;1�0pZQ|#�DF��tr?�,�Xl�J����3o�m~���tDv�Mh�����ɺ�vlaG��@zHɨ1%c���EC�xe�����Y��T&xw�9��SP�s��R�X|��j����u�:������m\H!��}?��J��>E�,���;S�8���ӡk�/P�G���� Ɵ�����US��A����h<� YA̕��c|�6ȱ�l��]ST~K:�S������{xwwUQ�s^�����d��O�T`9�fُ����v�~��<�,i�9�ye��_��J4�<zP���j?XS�V��tc�
L����>臡���F��w��$���,��H7���o`��Du6��o4&�])�t[�U�%��â�K��̍��B�(�}���\O�@U6�y�����O��D^�=�jŕ�si;��M~��J=Q�ʼ��\���ܘp��t
��Ȧ- ��tJ��R-cD��U�|]<ɰda(�BJ)=3�I�؞2�K�����PAi���Q�$Ϲ���\�>�N8��c�5��g�A�j�t*�YӖ�Q��!���a����>d����+�Cs����쇾��׼g�fY�e�V�a Ҵ)v-R_6��5�q�l�-�N6�I�2�9�
I��iԉ���ƥ3��W�tv�g�5g����Su����*����[���d��u�����a�书�e�H�}EoE�G��]��"9���n�d��4��T5ú[�~3A�U�k-�������k=������i@�������WKҷOvܰ59o���kf;���Rqh�!�Ӝi9=/ݍ��v�Qvb��?��f��L��x�k>�5GU�z� ��ӟ�����.���̔N�ũx<U%�>�;�\�/)ر��o�ʐq�]��1�qId����P�	��.dʖql䜒���c�7�y�>�s8���P��@s�B��]d�Qht��מ�x�6e�)��Ý��WS���
��H�AI�T���qlu�+`����@!��)��ԂL*\�|?:��t�2��R�5�o�<����*<��h\�{�t�9���]1&4�6�+V�>g�Lt0��ᚇB��%��V�fPQֵ%��I�s�Xm`=`�(^f�����V~�3TK}�~t��b��T��R�	����vx[��T�R�b௸ok�D�3Q�u�}���}ԕa��pFZU����w�������pY�N�:�^K���B��M��ۦ����W�ZP1��Ï�@Z��$��� �R��21f5�Ƅ�|��V��7`p�j�Xo�ԸIdB��;�s������ �	av�kL�x�%�4���Eg�����x��x���p�Y_e����f�H7�\��!�G� �30���Y `T���}<�_P�>r�ߗV�eΖ���2��+��3Zn�$�[���^l��n�������}��铍��<Ϗ1����9���ڄ�h ����:u��؄�QΗR���`,�ğ=<Ce�D���	��^���7<����ZW�#6OQ̀1�v�)�Oy�~��9d����|��6*��&�s��c>;|�y�+2��S�K��Wed���h��ˌ��t�@�y��	�\S|���'TQ�M�C޸x8t�qH_&�%qcO� \0�<7�+�����_���0݆�p�{{�N�R�h��w��}�|����m�d,�����sL<I�6�&ڄ��+�uu��H�.��R��̉��o`�?�̙0�r�rY�H8O��s<�i:'�}fz���>&>��T��+`!�(�t�3i�����?څ�e��Kצ�q*+@w��E�C6�Ω��������g؂�g	-K1�5����W�u��/��v�	�AO#+6#T4OO*�Kw�\q�\t�o3 x�0#=�ZLoH|R�=�dZ�!�Δ��"���˹y�ԩ�>�z:K=p�!d�p�tq��V�C�|��93`�Q4"�8\nb���Yd���L����V��B����ߩUx��VP�f5y=��$Ok\�m)�L�z8'+`�/�}<��X�̀�sc�Z���єH?$t�f�]����+0H��\��Y}��@�ۍ�l��Ou8p#�D����s��6%!�M��w�����yF��BJ�J+��n	��5�a���fa~8a4��~֞e���o�~-��&��ɇD6Qxg,_��ùEGv�A��e�xmQCN8)��d��A�9۽�x�A���e hL1��aF��?S�f�\X����:ȸkZ�	��׍��o�s#�7 �gQh��# �Ok\A�Ԯ��39)�k�[����s���1$FxR̌�s�|`X�@�6?s����u`yt�31o����߿�~\d�lqx��������w�b�1l�B�R��,�%1}�ZS}:�wUc��y��&�AⰚ'�A���\7��૔�%_ԍf	����yj�ck����vc��g!ue��vcj|M��%vs�gA͊���4A���k��Dg�<�o�z����$��}��,�ss������͔ں�,u�:��՘p����/�>m6�14����i\�EL�E0���9j06$p"�*�����#��8�+��M������ت�ى��*��+�ill��h���Mtp�w�aL��3������������7�va3�)��s�`����lW���A������[����.�����@���gq������쎂P��z�f|��?��YOfCs���]\=O'P)�N��"��>��؀�ϹY�*(���E��D񷡞����9-#���QLV��@����k�����ϒ�sR�2ci����v�@yZ�vئ��`�2���^|�z�����N4�@K����GO� ��b�����̍g���K� �ذ�Gs���@;WTaN\��)J�IJ*�d�
��~6��
��T#]��zV��A�%���4)a��{�sM:������.Sa4�:���@�+�O��]���`Q��$�<op�����*�	A���'g�2�B(�pb�᫯�d.����aY�k-����B�2�3�xs!)�$�櫚0�΋ȼBN.��C�� ��?D6���,��/�����Y����^�)NamU�z,46Z=���:���>U%�
�s���E%�Ͷp_7_n��a��_~�%��o%ǃ�G,�������h9����Ad�ܩ�r��6N�a m�,�`Қ?/׼JV.�O�|e�L�����Q��Q��F�+���
��o�����k��~���u�^xvo��A�!����U?�j�<U��Z�,zg�a�jm����-�a:~M���)�i�����\6�D�M�*��I��Y�ml޼~��k�����؁��J/��|)M˄a*>){
�VK�iJ���=a�s�����X�'P̙�8Su.�Ԍ��.�/|��_��nV�Q#*�k��Z��d��/�����7_!��{���5ӥ�I��Pu#���o��vZ�G�%g�%�O��4���^w"_6R�:��������j��ʇ2����*�N��]Z����Y
z$ç�}1���,!)�]Ӕ�u���86�L��������#�n��q�Z��k��g�so�Q ���]<��3��nP��Sg�vI*��k��P�����3�M<��1�3��[��9����7�x�2�f�!,Z�-��,�a�}�ЉCF����lVaTU�􊢴��;�Q��\͜��Y�^�u 0��X8��YS�j��ЄG�v!��Y}ч�~\�2����F'ϴ"nU?U��ke�0yv�X���?^ދ��q�T���?�5�C�T�Y���&��JYf%��q��mq��_�޴M��H�<��F7^"�������3ϼ��F�D�諮��273��@Q��T	@wUVfd�����9�*I��2�����3��+=h�,�tf��qx9�
ㆌ�TT����d���\������AjT�(/u�����������s�繜43E˴�&C���1C�{�@���`lE3e�5�Q$l�a3�OY����y�3Tz��CD�� aT��3R�"f �U�lQ�7+1±��J^�_����H�Ya^����e���snTm'{V�QJ�,����q�ㅍ�g|9��^�����ބ���(K��Tx������v����q�_�Y��c����Ȟ=�
��Ғ�2�/,���)�-|�C�y~�Sx�D�D{���-%�F/�3X�@0Wp�7/n�3���d(�s3h�vS�ʼ���Ȼ���f��x����ja�	" 'ϛ��e�fn6�����ȫf~:�����������Q�uqq]S^���$��ݷe�xëP;��=aMk:(S^:�Z$t�a��<�a�\��^��)q4\��^D�
���_օ�<�<��<1��d�ڙ�u]8�������Y����@q.,���&�J��:�+�-yu�w����FF�&ԳHazF��iCp{�Y�$9��-شBB48k��	��ث�1������9�Z<�vb���uB47�ڰj�;t���
5�10��D	5.nvVe:o���O�A�YȤd��& ��!�|!{*�Q�]��9��/̗���Z%�R-�k��N)�,$#�[u�)(��������9���U��l��$��>!w��W���x*�j�XOF!d�f��\�����TI�J���B+k�*��N��a��C��V�9{�.���P;�����-ͧ���kl]jcI&�b���QlӔ�x�=��[;W-{Ѧ������=��ԥ�|枚��T��4���_�ƅa��H�n�f�e�rF�#[V�������u.4�֡�58����W�aX��p��2�N4��jz�1�o�S�����&%��ū�l+�QL	p���˙���غ�m��C���+o��
O���W�%����f⬲���#d �ք�+�!6M�h���?��fC�[ukdOx�!Rr��Fd�*��!
��b�c�����&�����3ϗɱm|v�尗�
�\:��KY���g˭6�[�%����|������ oG�S�|�Mк��{���'���٦�<���z��˄����!ڥ�Y���>�:�A��!E"'���&0n1����! ��9�0�u6�mϋ7�.:ֵV)`�����û�w3��}S�xP#>2G�C�
�zX$ɗ�p����.�(ŵ]���4+�����.��@̮�\�,f߸p�VL�{�B�!p��)C�z�4�MV����X%��WiR2V���N��:l&R�"鴰�[��v Ī�ڵ�0�� �sb!aA���|G�k�3�e6/��aN��;Uuj�	�w��!)lx���L�	z8��^��gс�k�9�*l	��y��c8��L\�?t���úby�H+d\�:6��	�_PJ�~���uL�2�F�$��X��`��`�34Eql
W�g���Gs�:���h.'\6ROg��ս��R��}z����+�4Ա?X��M�愦H֖�X ��s����ً�'�9p%1�Cx�1���ڪk-6lz/����yn�'A�;��{�L��F��ȶ(BN��nY2D��$�hs��*dS9jf�Y�9��S�s��>!�C�S�l]1)�,�1�:>˔`�)Q�B��m���
�۾,�:��sn �<���8�-nv�8�V'.��zuba�4��X��~�Kc��i���x�����~�E	�ޮ�U�xF�m�E/��$u�Cb��1ZHAn�(l-������}Rg��!&bC��V�!0O�|�3ͪa_�'ɏ�%P���sk_��*�c�Q���>tHI�~������'K�O���u,�ZE��?�׺iʧ����ں��&�i8�z�s
���h;�e�6�"�ҖUG�q�N61L{�c͒E�'�$��t�+k�Rv��'&ux6�� �wֆNf��A�~z�}0 r~��ދ��>M�8f��^����6����������F=0<0�o����n�1���P���]SWT��o(�O/RH��m&�ʒcgE��o}�Ǐ�Vp4J�j?&d;1N�a����)y�I�2�@��vR��J6N�����t����Om�5 V#�q���%�g|��2��	�?�^��9�J]BDz����e霱6�)��M�4v��(|�x���3�X=�6��G�ԩ�'�`�5��i�5�����w{`���z��Y���og��E�푾 JP?��˯�� jQ'��<=�PӋt����#B���U~�!��$	x�����TIA*4�����5�{���0�tg��M�R&��m`�~eY��ҫ�
',Rb�wz���Ԁ�:�f8Al�^]*iy(V��B��ob?���x����P����;�c0�-ϗ�I�N�2s[�eNM��d|��n�ǡ�)�@s����t�ӫ�Gj��E��9��l!f��D�h+�{(C=F��C�/��ۤ犱0���?ܪ)E�y��HY�
�Q��!4��p��F�w�#��O�j�ٿ�	;W�A}f��_�:��js>x}�>�97���I�O��u�"|�L�G"m^B�0�s~����tō
/h0�q���懓M]9�a�Xc;IM�y����<��{���$|{��"�Oڙ����ϡ܉-A6�?|��r����|v��M�!b�N�%<����"����C8�rᛱ.����#N�����@R�!��:=;����h�dIP~��
K	)w	�c%[�opPWrԶsz&.�m��2���0;����uL��Ͳ���d��BV�E�7`���t�m�׺�^��!�'���:�Z�+k��q�QR��7\�y0M�[�
a���a�꦳�7��\�Q�M���B��ѥ�Y����c7
c�M��� <y+R��~�ǵ�,��}N>m�5qJČڶ17���y]$��6vsN���B��
�x}��Y�
q#��?�v,]IC5���|x�� �#�?�y`<�n&�;�cͷ�
��hH�r��ܤp��3��p��=�xƙ�l��]��C�-·9ڭx�Z�i(Ð��i,ٕ�6��]��&��4����"'s��*���gA㨶�j̆D��B����*S��U� �VR�5?�<= '%�Y���k��"���TDb�]\�!�c36y��/v$׉[��b3I�wV� �k�F������z",\��:*W�ǒ����{I�$^�I(�H�_���%f'R�ŭ�t#��� �Whª'�0�����7���ز�ay\��-'�BS��c{���p�,�Ɇ�zI���q٘o�$"! &B�[W�jQ��阚��!��a�0t��N�lܣ�֯_�$�4��T�Z��&�B����9�9���}y���|���/J���Fϡ�e��&dU9�S�qE(}�"#~?w:���\�qu�M����?�K	�Y��
lv�VЂ،9�T��⊠F�CN�E�6'�Ӽ�$.�؈�F�a'�¨��Έ����D��F��	��+�=f�Ž��j�qAGؠ,�hŬ�bf�^D��[��d,?��~��?P_�#�\/����CR����{P�}� <���������F��u���1J�v���}�8!w+x�]f����C+��qg���l���>k�h�����j�48ie#��=�~�����x��
�ii/~9��$N61�m! ��F�o"�����������ڐb1�ر��m6������;D�z)����Ƭ(�}҆��{s�p��@�Os�ڑ&MG6�y���l�J�'�����C�=�C��>���X$��Lzα������4�����GxH���`�+���z7�k��O�G|6�~6��Mr�!��.�����U[�V|�8��J��hI�X����am�)���!��3oŶ����K@�}L��F^3��P?�j#��H�w��{�_ڈ^4�!Ǹ�*���! �>���1"�\WL�cӗ���<�Ļazx̸&~<˓ۋ��
�ssK*��E��k��ٷ����F/y��B�R*��7��$CO���$Ey'&�f��ʁ[I�s����",hA*�.��;������G�p{��/{ʘf4湧�}xq0"�e�)� J	�8IԮu��
�E�"��7A�Z:�=�����=���?�9��KB�4���R��4�r+%a<iH���U�8���������ur-<Ү������(o�xF�Bf=��|L�',p�0��RD¸�����a�J�'��,-���ƽW칅g�(;�l���(��MY�{悥�u��c�㧸6<���{��FLx ����󰷇�����K.x�8��M�]r:q_$g6̻�[��4#e��8lwF�%�Gy��H9o�p���ԵC�Z�����^%eɞ�<7�B鵄pD�_^�/�{�x�~��X�Dt�����`%{�}_�\�\��ց��g�������-�c��V��M�\�]�D�z���(�����:|ZjE��^p�{ka����`���t|�}ӟ~ǉ�Y���fV4��H�����<��3~tƬ�_4��b۳͒?%~����P+#�����bW}|���J���I_���}�u��lw�����/����p����Bn0\0NAΎʭ��2n�&W��Q@�#U��� ���_�3�Q��^�w��1�w�U�կr���$ak��x���K�tH���f��;5�;�~'��j�#���}nL�|[舙hOp&�h��ś�S\��^[��:�}��p�Z�^�z�s��8�Ɇu��3�#�����B0��tD�z��q�F��g0�Pu�H�s���|nx��y$,�|���"�����6���
��3[���s��3�p��i��y�}�)kM�ڜ6��Y��J�Ig�C~�xPB����N��M��s�7>�v}�	�(�ё��
�	�k����L���>Wb��p�]��ui�)�gt�DD!X�
\�������ipNx���e��?����S��#K���#)+
�u$����0t��.�,��Y'_�^Pi<]%^L
��T�~l�l��0�_[\X��=��H1���� ��+g���Y]�oC�Y��<PS� �{d4�
��5ٸ~,60��޿̾;���8�}r*��y��Y�ܧ �cr���w�V�_U�����ۑWiO�"�̺�MR�p8:��!e�z�6H.�Ov��s��(�8��A<c\?�@�p�0�Ѹ��N�7������p��y��qk&��>�u�y��q��[7:��pٔ��*Mo9-\t���L(vjW��}��=�e����?f���-E\��m�k$A�
�s7�{c����7�>��t�X��S�xb���Z# ǋkJ�1��O*� ��x���d��T&#�����i;ȟ�j�<��>X8�29zҜ���f���t��t�L�C�S8�O�F߽��Y
0��xi��_�5��B��iH?�%�YW�ᬋ�iR�"2d�@�n�ޛ��^0�l�J��.�/�6���|6T�م���7����ɥ�!�ǈ�@�ʿ�뿖����H��w�zo
���燞'<�*B<�mh`HY�|��(-���v&�s7��s�/�8����?���.�c�,���Yp<k�V��[���Þ�O�
�>EΞې:�7�a-Bǚ���!5P�hV&�;��	�)6��ۘ0>�0���q#ևMx���_"�v�Fa�����T
������%ädU!�^�0��-���0h�!�|c���D��o�(JR�~�m��w4����`٬�x�k�k� �������>K5#d.E])������ex֧Iz���	����B-Cl�Y0�;fy�N�u��W������J��Y�4f�;�:�3��%E���Z�Z�d F�O���gF�Q�J�+q��ݻERSus�h}�,��.g�iHO�4���{�<�_�C�����f�M�n���-3e�wp	+u�Z��풡��n���G5��\m]�=���:P����r���,�v�+���XE�q%S��ј?==�'�ٛ��!1����.R�rxd�'�����>����@!�R4�L��g�o%�8Vs��9�������+����ů��'s�g�R�H*	����4�e���.���R&�o�#~�"�lV8�^�}lf,~X%���a<
qPZ�6ϕ��)u$��γZY�5=�،ѓ���j�0ޞZ���)�'��ߵd��T)�����k$s�@�EGu��n��.�&�w3��Y�kVߊRAd�*�]b��	!W��eC�r��9�ÛH��9�ZxO9��C���$������ؑ=ĂB���f�Y�]���k��?:�i�t}�M���j��bs��wŨ�_[����Z�̒K���ͼ5_G�9w؍A��Kd4���J��^�?���p�����N�VIQbjOV�ƌ8�V7�<��BɢPY��k��Hz��~{#�T��>����#�2�O��p�mL$�S1T��Xôf�9Fx^��k�n+��6GiJ�Au��7��U�8��]>�r�x�m�6�΂�"���-���ׯc��0��.���`H��ѕYg\�FtYx����]�04�p��GUU��&�����#��E.��Ԧa�ƀ�Vv ���[���Y��Uy�6�}�i�pe�BS��1>_�1Ⱦv��N�\�Qt���Oɓ���AB��C�z���8>j�����<��HkC
j`(��Q�Wz3e_�57G9�O�xZ�Kb[N�I-s��u�Jgx���6�I�`�x#�dk�:�(R ������{�Y��Y�4���y��]�Ǉ��E��zld���b���8��8���0}Av߻��a���'�hX����� w�=3��)C��<9\�C�׀�~�؄3�!X�]:	���Cx�H
�8ؔh�q^x��_�ބ�|���Kb�y�E(O����>>�H�\�K:>M�؋D)+6( a��wxn�;�㐆Tp�F�W��s���j=���W=�y��Pa����*:�J���uL)��18��G��w��}��> �"[m���3���9������x$^ѽ��e�>��"TuB0���
�Ϛxl�L�n�x�^	ZYe�?W3�V��s⩧�����UHC�7�j1�5�������b� Opb�ھߗ,�h�7ʀ��#9%6��3��-Pw��4'%�R����;ʐҋ��#�P�@ϯ�J�ׂ�V븁Dq�iD�}n�Q ��ĵ�(���������}��Ҩ�U_����v�	�Z����qK<���ڒ�S	M�!����/�M�{L.jY2tv��:7sy$^Ȱ�C�,�y���ق�����G������TF�u�ᑞ���'�`cpx���pzw�H��[� %�u�S�1�������S��IM���)[�Pq�}�F�^��|E��L.\����j�	:��A�<Ր������%��?i�U��'9�,��i��+�f��5i:�� lT�/��^���:��e�L��ފ�{wR��O���u��M��{x�a�T����I��XZU�Y"��ͺV5��4w�E�vA�W��a���6��m���ʢ:�1�K�Q�|��v=p|���H̬�1�����u�n�HbEj����0y�� �
�M�Q����k���%%�,W�W-��s�7��N�NԿ��8^v�G�4e���e�S��吶I�6�?�V���Ϥ?�hN2�j��R��(\[�vN���ߊ�K!Ȕ#����5$�vl�l�+��K�$�f�h�BayQ���6���~�m����j����
s0�Za@۫�e��9�'MP1p��1���'���vL��(��+��r���4���3�X�5����&�N'�mc!	�
a�j�&(����:���MlŽ��v-mB��O������_��Q��S$jH��(Q������e�&���$ի:�43�}&����8�C2"K
��-K�u�'�H΁alLp>$��+��	�Q|S^'�w=����!��Ƙq��gG���g{ޘ��Jؠ7�����7��>_�/1n���u�#�j�={�A�R+h�=���G����>$w�7obְfD���&�_���Y�	B��S�#��;e���Ny��qp��jdwS� �����UHy�=ϸҰ6�i�觎�H�Z�̈������J�h'�C��^)xB�|Y�*/��Q��Jmy�څ�$i;F��N���	��N�=����Q�6V!����ݜ����.��@�p&q�O/��M��t)��O���ł�F��� cf��D���|N�uqia/��j�R��k��ժ�)��������*�ɞE������Sd�7�,ܐ�^���8w4������ ��b!�e���MUו	�ƻ	��H�&,̱�@ϋ�4�)a��rx��^1O��٫2성b�8z���%��(|<G<�,��L��v�+�]0|�bH<ֲ�0�6��D*Y�غ�8��"�l�Ĩ|h^8��0�N���0P#A��Y�F�ȣ��(����{�a��Ο�q�7Y[�����W��P%����%��!�����Y�f�Q����vS�U���D���))N�M0Ֆ6A���D�f���"�vYj{��!����i�@b:V#ڥ�l�#&�� ��{���-L	��m��T��+_d���Ζ�,�"cy���9]�y���6����I�QwJw�ă =ɭ]�W�M��l\��r;Ff4�qېz��l��������0�`Hc-K�S*���;>�	��K������m��SLث�N
N�!������|�<����:�(��F=�ߖ_�%ƚe��u��jH��}80ׯ��*
~��m<;?��6&�~R����n�
�0O��������"׻G+�ǧ�.tF�z��H�ʻ�:�+�(,}�ถu��3�1�eI��G]�e�x~�N��W݋���T���W�?'x�_��B'y�e�G74
��MF�A�M�����Z�;�%1v�"#�S�1�*\�  ��IDAT�#|T��4<+��_[\y͒W�p:�N����b-����<��y�'���>i>c,\�����,K�d(c#:/<R�����#e�ܗ��Q�z
OUw��F/��=�0��6�ւZ�T��E���h��܁�	�� 5a�6�E�uYc$X���{��M��d��<�m�����2[�!�!��UM�.N�6��S��(Ʉ�r�I�;d�6��������$���;6�,)�+ZI82�Y{_��t�fi��@���O���W}�v�Gy�6J~lb1Z�!����̎�S� _�W���X����e�xƥK�<�ua�Ӱ�D�t�!b�W5�h�cx�������^�&�$�l1��$yF
>�+�p�.ѨP���7Z/j��0rY�=�<iE�w��/�������j,n��띗ZU��Zk~�*��ߍ�&5�2���.K^�8r��u��$����2*�kDv=_�[Fc@�i��s��49��x�Mh�MᬌL�S�S�ޙ�Ec�h�k����kz���.�e���~�;�kQ�ep�Â�@����1�s�ȝff�fo��Y.�;.P�������Z�ϐ/kh*���g���Վn:�:/U@b����+F�/mc7L(B��ɲd��j�9�ٓG����>Cu|tY-�=w�u����{��<��1�n
��?x롶1������I�	Oq���
*G�!rB2����>F�ޠ9��6.fɍ�Z��V������ўm1���Ќ�������h1���K��kR;�Y��'{G$m��ɶ������C@�w���ï�c��9�Q��"�/�|Y^�=A$�0�U��$���R=$'���ê�>�~�8�LC8�n���p�y^���? �d�����"�^��<e	�F����'�	N��?�ujS@d��׫���"�Y�]UeƭV�Xg;m��h!���N8�N�U��.�=	�*/�5g6r#{3�'G����������6�ɡ�fxN�,�4Fq<VQ�")8��b����}_�wm�ZN�)<J�'��W������r��ަ`�_�5��N!���Jf��6~k����NaP۲L{eX4nǲ>f�Y�x��^��rEQ���n�ʄZ	
T����~'�VÐF�z�a!�rȅن�T���И�ziT��K-`܎����lWV���}��!�B5����,~<��s39-�aoƙ����)r��֙@���1��S��o8DS^F;����+�j��",3�Ė�w�%�x��1���M���/���u�3;9����S���1��x�==H���JT/)�s��ج߫·y���D�������1����؜8�NX�y��}��J�eͱv1�O�vjn9;V|-j�E ��P�vP�L�(�e����?��Y�ȕ�7�ƈ�����[��:[Q��(f�	6�k��߅��O�'�������x�wu���E8n6�����bń^��\�J>��x<{ gån����M���A|����㨕9��[q��V��D��i�;"��W���&j��m�b���A0�[P�־S���=���&���pʼ[O ^M��+t�(ٻT�
�.p�_~��E�$4"L�G�ؐ.)H-֛0�7���m��1��q�&f���y� T�m���&ww�d��*�
/g���OE��H��X8�
x�G7_S՛���[8����o���÷�r7���Y��::���g���S>�AIU+tv�,�����^��l�����p6�>���2��S��-�=��p�����M���^�Zwj��SSAl�ߤ 8˯{)��>c�\�s��T��Gm��h��LVA	�9v�H0�P�������V
b�E��'�qH��W���Ԉ�j�@��8��b��\��F�0����g����1����1�=Y���0�cN��y��>�hJ �|GNx#n�Pq�)@_,ĖZ���[����𐱣�/]RS��D��#
I	5�3�������~�L`�r�Ȉ��	���Q���̥g�Z�Q�h�{o��7gbI��FK؄]{y��.��,� �e���Xi�`�1����0�-�߯r�p�sxH��{Q��$�QY%��Js�Df�|�~�8������u��m���!?��[wq.|�5^�h��E�j�K��C̛��l|�W��z{6�f8D��Se��Ð�yo޼JJY��n�L�M��Bf�	�E��:ot��P�A�,�8J�f9����q�ដb�w�6������&������^��Ý�ga�9���K�2ꤡ�7�$�I�9�b?6b@(+o��r +9,�� ����D"|m�}h����� \8��_c����-�$�+:4N���L�j#��1m����G{H$�爨�R���ܠ��!���]\�J�W��h�Ti���{���x)���vN|����G��jw���]mGڄ�b��Е�����/�oc�-ὓ��k���z� �-ͅ���ED�$�����(&�[	lDE�L�4{ۭb��H�fޞ��� �H�F=z,�f%xf�+3<]�ӖI��^7
ZS�5([��zm����$�&oj�D{��5�n�xL�%UM�ON��tX�(�Uxn��'6¡�K��c	R�3� �ީ�5�C��v{��aH7*���}O�lH������ta7g�Y;ǂ�^l��4)=���׆��g�T[����������^eE9B�c�R�ׅ��wGO��:�+�z]d�#k}w/j[~�gI��MR�T��T�੧c�
�Oz��ӄ9t:f�,�n43=ϣt}O�a�G͕ʕ���#�y�N���>��]kA3�� 1�Y�)ְ)bv H�B��ӺT"Rς���<�rD������{���e�nb����=#�V��<��}l +m�ﶎ��͢��=�Ih��Z��q�/�⬽���ih	J�/xqWal����� <H��\f���I ���7�D�s�2h�oq�K>�e��<��φ�ݯ��#J'��]����/�F�t�Z�ͷ���(�S�7x7m��:�xO������x{}6lq���!l�Hx��=�p��Ja6��؞����&<I&WN�}p������[��0�!*�wՉ��L�mE��B
C
oH����I���c��?��H]�����
�N8^�_"�q>���/I�:A�b#|?|lc��p���U3= �$y�;$����O�^�Rj�`�5<�ׯh\#4�R�}΁��6��B	b����1�����J��z!��	9����H�T�q�k���k�:= ���w2js<P�&%�NMa=!yd��KL�t��q���HO߷Y�@��������Y&����]Ipg,)�ͅg�n�8��Xv1��agC���iO�<�k*ʕ��֨�9�!#\+���{�}b�޾
|�p��eAh�Y�G�𮧽).���3�Y�"����s���;���_6�'c�a�N,w[z��W,BX�*�4��׻�w����p ���~�79gX:��^���N���9CTa"v�l�p��j�M���Q!z��W���A}�3�����5�>V�������B��ߵ��ko��ʹ�$�G/�/K�\1U��g�)p�&�Imp-�+��
����J��I����X�T��0�I���TQ�Q��UO�}��ە�*[�Ӡ
1^;9ʆ̿$�Uk�-�����^+�K�6¹��	JV0U,7*b���{z����<`-+���ی��}3W_]�x�A�7����s�>�a�s�)GS:5���I�%7Y������W�{z�-���h^9,V��^4w�\ys�s���!�m�mg'�mEe8&M0�R�J&�;���Z^S4zJH��˸�g�o;U����F�S�=j��3�ȯJ:W/�΢�T2~c��x!��˗��N�"��<�����}����QC�i�\r��0Z__�4^���Z��AF�����9L���S��D�MC��4�ßib]��9�w6�Q�¹i���W2����%JH�<�$��A*0�̬�+��$�a�	0��+U'�����)��l4f_�/���g5�vJX��2�A�JB���$������N��ǆa����> xmG��z����E�J���b�����]�o»��E�OlN�1�Saˉ����]�C�1h�T�I��]�U}��<�	Qa��[K��V�3���kh�[\��1��+��.>gXƟ�3`, ����9.�ʫ��fo�j��9���ڃ��=�����%�c����t� �.�l����yc��oazw�]�����,xbE���H:ME�5��s�,�_�ò�������Z��??�g�c|,�ec�z�ܪ\2f����H@�E�&oq/�����^�Տ�t�y�}���
z0�hP%A�]y�E�p�IJ
�[]E2��UTX#��K%=��m��ڿw%���������s�*%�5�\4R��{��2�L�u�����Y!��
��]��=dE��_����taHݣ�5��Ɏ����=����z����n��>�b� �y��U�����	È�8^I	��,���s%6�V���N,�jo,�R�viǟ�^�~�&�^?�Ա˞R��=Hպ�������G)�՚}y����{B=���)�C�f��Y�,�xА��'��b���7�!;EL�̆x,"�'r]�e62�W�*�h"�S�	���I8;me"�JO�nDd[F0�Nb����ؗJ_�N�#)�7:�'��W�O/Z#�c4�ѧ!�bsws�h�x�}��A_{6�d�-X)�u8gN�9:y���[�����ː޲]A���4������ ��#= Jˁ�y�1OO����r"���|
=��ߩmn����q��2��D���gA	��r��Ԣ�����?M$�pf�C�˪�Z���+��n+o��*�)�u`򀒴��m(���7a\p�H�g↳�� ��W��*V�f�:�?{�meӤ�k�ժ�|.7ě�)iR�Ԯ�.�mȽņ����/�f��,�<KB�3q��Nm���y���]�fs������Ɯ�@�Ø���@�����G@d��e��.��wL<�,�gJ#���v���G4��׫vQ%�6G5�c��5�wV=6�ۆ'��8QG֟qT6T6~2cf�ɘ�z#-[&�!�RXB4�Ԟ�'=������F�B
�l4��4�Ϲ�srq�ui��-\��x���)a.b�N�	H	��t_�r^��-X&�G�A��������֘~�0\�w|�gS�f#|iփ7Qgv�;��xK�2<웋�␺ �t�:똸%���~�	��AA��\Ðx��hO`���)�����Fa�v�s���2���x�i2&y���+u�r^�eNo���W�\�%��ߩ��	��{U�P��2h�%VJ��c�	�_�8	*3�P&n*�m��7&�2��D�seuǈ���R�k���c���;q�8���?�
Uj]
�HC^�y`P���?������a�&n�o��{l��D��\��\�׬E�WBԪ���흈��D#a��k,�A����3���ae�6g��z���n�����*�@(̽�J~߾ߧGm��k��5�B�)�xR�P��6�V\r,�[ZJ��3L��t��q�Z'�`�n�)"����L�a��[m:q��~���Ԉ�o2W�k����Y�]�Q�F�+A����z�X�]�(v�x��)ۆ�Nb0�̲�^�� ٢�"�PsS]�!��V3�Q�p�J�V�yjTV������Y;sW}m��))�6��n�㞽����:ra��j����J1�~���^�8V�g��僾lU�Tg\e��DlS�[��u�a���Uj�����a�w�Y2�$�R�����t.>�d*r8�S��Fh��:ذq�#�~ ?rTr�%���X�U�K��?�;$?��x��AX�A&I��~��&����-a�Pܯ����1|h^D��[I�H,{� ��z(��+$6��1�BX�[� ��j,�f%�v����h�`�vsu��Ҩ���T�����е�u�����u%J[x��ǅ׾<tKB`�w�� ��$�А���Q��^�e�x)�f��{^=e�)oSHi-=�9�	C Q�)� �����u�^��FR�,?�~ʈ�}������1�?aF/iQ��L�Pۍ�wq8d�8为�J��!�f5%R����6pV� ����CL�t�� �uJ�]�*�G|��`!`�ms6��B�ºU�i���h����܃�=��Jڟ�I�9WV�?�����08�X\ ���:�����7�������J�"�u�Q����OC�L=VnJ����i����\��v�(�q��U�=7���!u���aCꌆւ�H���{�Q9�og���r'P���00���"<F���$�*�Y<?%�`,�%x߻��v���nH�}�M	O;.��66ni!��n�#"%u�E��iO�s�߁���O?�����(\������u9��G۞�6����raQC9Idz ��E|ǩ#%u�Z��5o�6,���w���ĵ���u)�l��{-6�1DV�q=+�T=O��q�wmD�ɺ���?�So����PȿTL�G8�1���b�ن,2p�"MD���1)�N˹��M=E���bu ÏʲZ�
�xH��O�^Xd.���je �xw]���iǝ�u���#���ޒrR��j�Љ�B�7����
���1靭v���!��4�C}�
y<��%&(�D�~S�94^'���cq�PЧ�(=�`91�g"�Ԫ�4A*^���p�JDo��ÆP���(O,td�^p�����	�M��=��-7s[C�ß�:#N��xA/���+���=#F:0�����@j�����T"jQ��u��"W�ƀ���y�߅��5w������2��z��?�JYt��?��tkAN�4<Zܳj�h�3/1T�)
W�>�1�����3���T�N�j�\Ga[:u
h��}N��s�G�"����!����ɠ�aχ�b�*Aw^o��4UN���{aJu��.��W_h~�"1�������� 	�2e�2��+«����ċ����i������K4e���a�%��jA�+x@��}��mϵڬ{�_Lrx1�$r&t6X?|�cx~~��d�Ub|���㝌�cY߹b;���=&D#���UJ�n�����	���%B-C�1�uC ���X���Rc�M�O�8rGV�=7��mFW�����3?��S�ن�F�P#K~�Q��B��P
�!H�iι�bR>
4���J�>i_gX���]_��"��A�w���lz�����>Y��lr�69 
��2��)��R��gEa�L��d�萅0��@☞�U
��;C�T�P�;�[�؅Wy<d�u`�á��7U�s�c�Q�BB3���x��X\,�chì\jU{��~p��cG�m+I-%��1�����O��S�~~���M��`�4DU���ou�"+Cٖk�Þ�[2`���}Ho����#TB��X 0L/ϓ��o�_��/!�*�_�=��۳�6U���D�;y��^�̰�*8G�D0i>d����\jH����s�� ��U*���8�7j�^B�d_���sx�_��Z~�����/�J�X|�8����h*�T��[��ܪ^�ի7g��FE��e��!��Qy��N8D5�X<l �7�$Q�f=��'�&N���f��sa7X�	��z��eN]�ˉo=Tl,���Y|S��=�y#�i����x2�D��/�=�Â����'6�����0�0��}WWM&d�,"�X��h�(m���\=|>��ꈾ�Q��g�09&W�B�rr�qu�_@�p�I���A��f�ͪߚ{��xV�?=��:UN�Z9�(ȗ�)^��=�G�J�L��z�k�Π4��.����|���"����:6���f,�?� hs4ϓM������-��Y�Fk�掰��vc<4�٪{;���8� �-��&כ���ӟ������(�q����&��	���R�wP���*!O�
(�_˜'*u�қ��Ğ�)O�J�h��SU��y������˯�~p�,�J���?�!�=�V|]X�6�!�U�lo�=��{�����P�w�(j/'�����.��v�%�^��p��,�wYj��j8��j(H���kzb�a�����⋒�����Bs�	c�^��*3��*QF�P�е�^�'�S���Jd���#\�(J��}?�ǚ�o��N��y������%����}`�����Od���&�r��7�����@�UĢ��ŒS�hJt5V|��I�����0k���
��êO�B�xHƁ:���XK'hq;d��H����e����PW`�	�8b����6����n��#*/:\at.9z��Kבk �6ڧ-���u��co��������1��ͻ˒ڤ��E&�S��+���#v�S���tl��G		D���0Qs��΂+�a �dT�C�)x��6��p]�_\�3���:H�xR�zj2J2���Ҁk)S���F�jN!4�ݑ;/{R���)N�P�7���(���%<=SU�{��.R���N�X�>K�I�̳�o��g������gV��$v��/+}x�x^�.x�~/%=Y��F(�D���+���B�8n2�>Ӷ-1$�W=C-ЪV-˒���P	���Jn�}@�����}�z�i�ʠZl���g����k3LЋd�g4��u=|@<�k�WH�`�㑡1��OU<�fp��=��K�H|�h
R���O��3�����ؿ��)�n�8!�t:RM?��?f% �hb�Ɋ�	���z��;�*:��d�^��wj�'��&XC:R�-�<U��G��ڕ,,
oX	U�x����?{t�	}�1ӵ��}��rQ�խaY>�^9R���,w\��%�յ�{���t>��8��˕BAh?�?2��8E��{�i�1��B"��)�c&Ƌ��*5K,$�p�4���7�R�)�a��ٮ7i��Y���"S�'�W|p�)~�\�gQ	*���0K���>�Y�0��*(��b��҆�<������`D�k5�^�Crc�Ɉ�k�%�h�⅊4RwWXH=�p���~�-Zͱ��%_�z#��?��+y��>�0�]b���Aߒ�6��wL����dV�ͺ.�fw��køU���+җ=Sc����(rs�P�=�a��?U|��~W;9Z�*��ȕR�GzL��j�&��{SݘD;%�MK�g-J�zw���:�%(������J7�D��f&�"��:f��v�vPu���:�� ѐ���8|ɋ�<�,��x��
�����طj��ğ��E���A�v��S��}����4�Y� ����AȐ�/i����Q�<R�BaJ8�I�_r��.CZJ��孄��nČ{��~�wUm>��¨Vj}%��C&T��6'aH;?X�tSb�6���	q���A'��D��uŤ��B�^6�d�A�k�"n�!����% ���	�LM��j�.Ѥ��O<t��C�a$6��i� ���ÏaHq�֗�^�jl�	ho/�=�[@М�+ M�U������!�`;Q�6���:<��Xy��z�QJ*�)l��:�[X��LR����DH?�.�Wm�Z�JR�Ϫ��z����mt����z���gjUFG��#���9���_5,�h��jۍ �Kb���lq�h�B��b.����u3B%-��V�V�U�}:;l�qG."���yL�u͛�Yۋ;��bq���)�#��52�g_���sU�|iغdYl�ѻ�Y����8��r>�ի��\Ҡ.<��7@ՖU��J3�N���>e�(tb259��IV'W���@��M�l�YB��Wz�MB$��WמRo� �ը���cw�'x�I^{!����wl���;j��IƦ@�`q��jm��T�$R���ך��mP\�	l�ݴ,�k��/Ta�W�E��H�D�<�����.i�f*'��������Э� ��8Z��Y�V �dXUi+m�'5js�N�"ʉ��&N�1v�O�Ns��i����4pc�5�gO�m4���.u>c��[k��qs�LY������_-�go޲W��{�r��U8VQ��{瘙RD��j j�4_�0�!V���R�T?U5,G�lO稗A��?�@;�<+��OT��ss��E��f�	�2��B<��wh��>3�%�j)õR1m-v����/��˄�?����_��$T�M�d�n��-i�����b�|���͝����lY��fi��c��P��+��`����	�?pX�$ȓ��"0��f���RK�ξ� �튻.�)�{v�^�-t���	cm]4/���wV(c����>G�����fN��]`�F�7�o@2���< j����^����ȋd#�	B�	�N��1��mx�䫂�c�d�����Z�w��܆���n��nj���ޟ�E/��ۓ������Ǭ����]���}��#F�<U<]s�2~nx7J���+��]�MH�/9.������@ev�3�ctr�5��hP�������J7Jn������0�!C��P�T"f�ip�u�
Ǿ�q��09�}�37�=ΆÀ�}R�0A�k����e�_����g+�b�c���3��]�麓q����/�ѕ:��x��:?��s�5���������S��<	*^x$ލ����d�(#4�z��O=�uKf�X$�F_��X,*Ró)���!�g��mkHC}�<���ؔ'-�Nٵ1&ZYJ��);�+_~�%��KV�����Ґ��aR;�9H�Z�>�$& D�q��)�r�>J7af���k��6ɡulf�o�S���t2`�?��s�����!�� j�	,Ӝ0aM�!f�<�Bڮ�w�F�D�p� ��1Rh�H�<�)0ޢyG�@ߧ1u/=��_�^L�����
V,�vXLL�z\d��ac������%���ۮ���2�hpna4����+AmB�S؞�����L��C�Y�ǭ�p�w������P+�0�'�`�u<�6*�(ƛ�=K\�%nCR�b�T���2��X��H�F���� �m����ƕ]YG��Q�yP[��i��&��X��a9ϓ�z�n.�(9������s���c�JT��{��$���G*�k�.քqL&�٩<�I/~���d�&��b��	�F�u���8v�ISJ���W�r������Z�*��+�J�i�P/6���L�y��P��k�M���Ťps��o0\��=>��8��wY��hQ<*Q�!u?�Y�?����] ޸e[�mo���!�p�&�.�-���p����5�۵�=�>)>��������8C\�l�V
Y�&N�&���u�
���5����k�]�9�%������a�c^`�Y+)HZ�-:�̚��1w��b� '���v&0��]p�b��̚^��j��/Ƅ7e����ɪ��˵�QX1Z���bݸnY�����:�~���7���qxNm�9D��I�,4j�B��{�ӄ�vZ��O�c��F-�T��1�%�z|�z��(۞M8b<{ZϷ�/M5��]S��Ŧ�n����-|������ր������%v�נ��ؗ�q�2 ��^ ��{69�Â}{^�V��FWȌ+���g�6�&8��i�,�((I�~�^<�c$>����q=��2��p�e�ɐI��L,d�
����b�k�^���F=�4� 2�0��n�|h1�j�aD<�]��K��G�7q &�t_�a��9�ڂ��n�.юE���]���3�^هl�WڊB(�m���]��`6l����	I�~h��Z&�{TLysa ��e�e��"x��䢂S<�h�|������
g���a��?W�@���unzl��.=� q~g���ܨͧ��;i&t�^�d�A-�Ik�,�����veу�:0��/l���@ ���J@T�¡S!������8��D^8�� J���{]zf!6��D���*b��X.�Z��T-mq��V�]���Z�*��f��+5��>�]&}Qn]*�9�Կ7^�9|鑦�O-�m.���"�&���^�]���ʣL�|C�6�!&1fCWJ���?��5�/��>�iý�!}�6�W�'���rt��#*>6��1�`̉_|�D��	I.������$�*M�υ`�����:͒�P�u^_3��%���F��ޑ����&��	�����<)`Ha\.�р��]a��$f��dޥ1�i}�K	���A��u�s��:%��V��Q��SŊIzw
�&.���� �S�����w�}�{y��:H|��h���"Ď��ń�Qz��7��ECU������:��3Q�U����<!�׵������v
�Ǳv�!_��b*�.=�w.�鬀��٫4� ���\I��l�,�(��z��N�̂Ȩ��OCJ~rm����(�r�z�Pdg3Q��sB�]QݰnJX.��.7�e��H��la�y�3���\b���Y�*�j�>��(�����@h�؝����DH����yW~���^F�/�?���"�K�6b?���!(C�O�%"GB�mf�¨���(�0G��:��\{o��U�H��aD�6PM��W	���a�!��]�=���U��<��8����=��u�^�������<f��a����9�C`c-^\]䤋���"NLxӬ5ˮ�c�̗���w�V4��v�1&�8n�=�QO���0;#��ڱ�~��ʟ����/�����ߟ����%j�D��-��ya._ebf�9��687�mO��W���7�kH~Y�X�9'<��:T�B��X�qj�Ԑ窱�6i�(+ׇ��?yУ��E�k�cw"�Џ_��C�ψ&X߿.�Qg�#K3K|�N�-Rji�Q� ���!�?h�j�QUB{̜��-�5�;��X��s����pi�z�v�@�ȱ��'�~˘ڑĿ��xn�iHm,kVIF�|��c��Y80j�;y�s�9I�ng>(5YN<kTH?K���_��؋��]�.�;ӫux:��P���,l~�
6�-��p8
;�'d̀�锕@�-��Φ���c�x1�l[H��|�S11܀����*<������ۼ�mtZ#\�ï=)-��q�>�GW1&�z�6��R[cL�x>��&�&��Z��;�9�$u�T������ ޤKR׫J-�r�qx\#6��~$mM��FԼM#w��w�1g7�u���d�1`��lI��S&jB�wm���Z���0��0dnC~{�u>��1�����8gx[� �4���5d���DQ'��T���rׄ�t\��a9�+
B�e���i�ޚ����z���\�0iL�3g�m��cj(16��ѝ7ݒƽ��I�����fz�u��j�����9#<m���w�G���I7�X ����Tt�Ĝ�9,UV�J��MOJ �Yx����Z;��$�-��`�Vg\I5�e��x`7L'�Ԗē���ڄF����]0Bal�^QG�l;��C��<�NG�2���6t��á&S<Y\mj�CM��Q���>�cA#���~��5���9�4P-�����<`D��@��Ľ*�XŜ�.<_z�OO�������!q&uJW����d��5n؊WT����&y���2$��>>=�����My�S.F㌭�8�}�L�ʬ�7ShlD)&��U���û���%���@��Rb���MR�t_7��s���)N-�cQJn
�Tɏ���V�Hr��c���� kh�荺?(�D��]#����\F�tvl�F�,ʹ�R�L��
z�u�5�^�,�3Ų�Z��5v�1�=���Ο-�8���G�Cy�������/�!59��@o��3��%�kV�`p\�B����c*t�}I���䬊0L�G�H�7łR��4R��؈�	�,4Z;�p��c��Oj�<w��s�-ʱ�l|đGz��&�צ⚵�o����S!���s$[�\���}
�.�"��s�q�΍�]AYx6P��Y>0�	d~�"얆Ø���hS8��|�a�e�M�m�}�0�51����cR}���"	ջXO�L6���P���.� �'�yK�!h��ύ)�Cͥ��(LI��x�M���v%��N��`�IX�4m�Kr�������P�W[�͈��&>g�P�H���4E�Պad���3��K���N�l��f׆��MF7�w�JG*��<���:[�x�Ш^�~��+���B��g쀾���{[��)C�)c��7�l>J6�*'[��R��8ln�U���n��s	����Q;4��м�p�T
� Y�\x�7��c}������ L�$)/�ΞH2���#�0�q�P��Li"p���^�d�eV�t��Ŀwݓ@C���>~�@ӱ�cK�7O0�)�{1��az}��0�I�P;�O|�S�k�,�j�%�[��wݳ!o�mi\К����5n�w�Ħ'Po���eN�]9[>�P���8�����P)�g�89�[_TY�8��·M�B3��)�}�=��s.~|���cvZp�i�Cw*�e�͹u3���$˨IۧQ�<h�]��߻���a��������yΖ���jIcc��I����N�#�m�`Za�Jw��h���f�KfP˚�gZ�;\��0`.i��
8MtL'�tݳ��L��kD�Aȏ����S������E>���t����槉�����b�NY���+�H^wC�X\'�����Ʈa��[ɼ�㸻{�J�&�d��V(0NXP�
�7��Nl��#�d�S'n��WL$��A+j���h-�����k��n>����g!�$�9<�q]�����*���>���������RJ����k%%#���<�ΕB9c���'�ŕ)4�g�>U~��3���B����	*� �dfx�l}vYq��8�S�\؄����8Ϥ��s�w��{��c�=�K'�~�)!"�NDW�n��!�A��rb�������>NI;k���^�!�!�k[�Do��N�� s�4!\4Hv��!�ә���^�6l�1�`r�EM��ԧ`UݦX��etNl6J�	m�Ĉ��ƚ[��]UI$��!!3��֟�%;���jO�y���[�:~a�筗�b��1��.x��9�&)`:�'v�����U�Y:�!r��u����d��T<:�E�?��hMA��jCi0��B��u�y��� ��"t/�Eą������cx.m�����5АSOs�x�v�
����XO����U��%�����i8�%�V��[�Tȷpnbbh[|6��AõP�������4�NT7�;ȣ��$�T����(W%��)$�,TL�k-����C�c`ڛ�=�>cc��<6�s��Mm��h�Rv��gV�{��\���抱a�����w)F�4�ږ�C�[�����6�e��.V���5�W;��	={{�^S6��v-�c��?��� ��:����R�xļ&�3�)ӐVV����ۂLUK��e�JW1kϝ`H��m?�Dx�R�7���B:�$ �?ƒ�+a�}��R0Ț�Mɧ��Z�2���EP&wO4�p`x?}&�ξ4�S&���e}iħ*7�܀�8�7�6��QF߆���
�l���l��4j�B���q	�7EX�hO�!<x`z�-��f2��`�1����>�w���x	�&w:L(���G��̷��F]�_�믬��f	jx�3CkÚ���c��j����hX��&,L|�>�)h7xe��U[i�N�8�s�_�����ĳ|��#�������4&,$4.����g��C\� �
��Uo�?߮(�a��8� 	,!L\D���i e�4��6�g��B",s�w�i�Gj�%�N��W�9 �Պ��d�E���P�(����F�����՗���<>?�\ņ�{�Gj���0�/>%�I������=:{�Չ�^�;�:i�*//Jl�P���Y��d�a�h���[�pVՖf�������C�.��J�7iY�S@��_��+�P(�lOl�����s��K83�A��X��>f��J�R-����=6Et}���<�\d$9)��D�&�K,�&%1u��~5�4њi�-��O�i#Y�S·v��d�1�g4Tъ�v"᳢�\x�np5��y�Þ��o\q-ò��Wp+�Ns��8��Yn$tb�ܞ�c�&�`�/&�"��n7Ys^/�哕F�^Zks�UL��J�dZ��Eo-���W%��s� ڸL�����5Uy9f������ɞDr���I���	1���Z�.=agB�0%���z�V(CB�ٙ"Y�H�I����}[����X�)�I�<�?׉n��,�,���l�k�4^����}ɤԣ���ƍW�NDm��Rlڰ�1=ρZ�nj]���R;@��!p�=2����2�OZWmrG������^�|6���5�(I�E�\��o'��'͋��	��oRs26=�ٰƔ��
q�V��ܐ�F�sc�i�%��r$PΝaH�)bϳ��#�O�KD��H6�՞��+��B�+=�������f�:�Jt(Y_��XZ�]Q�!�t�~�͵X#����'j��*�%��o7ۜ������#C�٤Ҹ7��9<G�w��E��J����g��]���$T��pت��T[��<ܠ|�kj#�q���Q��u��8:|�A�C��-�*=�넦��&;�z�r(gwj2���]���8�G�r]n��C���������'�D�����A��V�L`{��m��K�>P�̂=����d��@S���OY��d	�x'�j�)��ߺ�ƔF�%�W#�$�d��/�z�+��.	Wd�>?�iJL��6G����z8�$,6ɞ�-���ܐ����!���}ØE6�6�Q��+��j���0��n�ס�V�����@bh�oklS�P����>a�`�`}�3?G��}�6�2�s�jU4
�M����?{4��K��v�Ն1]X1��7a�5�޵��c8�"t��[�ͽ�1	Ri;��zюꅷO�x��Hg2��Fa9�QԦ�3��7EX�������s�2�ky����)D�Z=e"L�V�?�%ӊK'�*��h7�k�V���aJ�'�3���x���?�|p���>1�.�k�ö�=�����9�����|����0`�J�kӤ��E��p��}��Y>��>�_m�c����zn��-5�GT�ŔΟ�S��7{��Is��:No����cR����0w���"4��N�e�A�3I�U�qt���⇀��;�Ic��
ٸ�	��&���V�a�Y��L�+�vx���8�?X���E��so�Rc��}-63����h�2�u����l���vO���xu�D4]��_l )��2���#�ǧn-	'�?Ҹ��%�r"��+��Y[��4�V����L�;\\I�Ek�/w��X����vCM�[����Y���R2���i�;�K�R��4��&�ۉ�� Wٚj���P\ؒ�aJ�I���j��,�o퍆!�Q{偍���5��ԭC��m��fL[O����D2/�_�sLd�]�f�d��će��cۆ�ٳKx��>Ss8G.���6	��Y��j���T�ۛ�?�b�"����ʉ2\<B`�B�ŭ}+�~^��z��G��:4�K󻶅t�w'8�@~у�J-]^.֌3�����5>/�4�udϽR�H9�I�vw��R�d���G*�
	�h���@z�6"#�`NA�,9���a��ب_8���1������.ʴ�?���c���w�����r�bH�͍?;>��3�X�Bkh�%EI$g��
���|��>4q�O�Ĩ�'�-(�c�^e�'}'�7�{��P�ڬ�m��~�:�K�����B%*��/�]t�k�>)�:7�j�� ��[3���h��ᢗ={q�䡚�`|�����¼�m�8�z� ~�I�a�n�-�a�KY2n��{i�\H�G02�*+�0�KÉ�=}��;s�	�}�̀d�6�u��vW��s{b'C�?$�`�����-�^��?U�����e�}�wr5����=c�E��X*]K��^V��	�Y�:-��&�:-B���0�J�yCB�m�L� �]�Aޗde�����%ǒ��ߚ9	'u����JnE�.��c�\�Y��1�#��t�A�zڦ��Sn�|pT"��1J"�R��_~M��9C�<��t:V'iY�ʬu"�?�_��\X�&�R��zm6��<4&��O����P$��j968�z�L�;�'UR����oO�أ]*Qג���~PT��d��X*4M��<<�L��>�+X�O���5)��mJR�K<W�7��{��v*�@g��+!_���p�VV�>_��\G��r:���$0�.!��ʢ$��I=��JQ�mfg�G,P��!�>��(�C�I
я�̭t����:�Df-8ˌ�8Cq��&	\��L0͙h �p�@�ԟ1OO�}-͹9�}�p�c�䕽GG��D��9���ËԢ��rb}�"�&O;���1��]k�>�Xd�l*o�!� ȋ�Έd���P;8D�4�jϿi>;$�!j���xմ�a�\�u�."lօu�֮[�L'��^9�꣇(�èdߨ��Rۍks��,�[T*>=�w�4�+���b8K����v:VC�?y���3.�7���'�WL$Њ�`�2���c���1����g><�Ա.�*]f`S��U�A%��_P����<�p�׵\�a.���~��ߣ���؏,,��}z�Y8=R�+�ӄ����6�*��6��f�~�u���Q��Ami0Lt�rG��rU�ɩ����V��8�K$��i��Z� }H���s������t/�k���#U�����H�EZW�/p���00��Ə�i�ᑺxW*-�<�j��d(0�Yu!�Z�5z�M��TKm��T).Di����4���҈�5���KE��'v���c����oYN0��YRh/,}8�*���v�굧Ę3RS}{&���x$q�9
&y�Ĵ�x	
5�P�Sl0%��p��[��Ð���0���^�y.xܜge�}o��>`�ḧ���������|�*��pS�/(��Q�P��M�ki���z�ckG���kr߄�"��v��z���;+_��kl�wY  J	�ZԠ������;@kZSM�$��ةK뼛�Ђ�ɨۖ0B$�NS���=�����XrQSL�A��}~6��=���<�j�;��N��C�X{������b��n�PIlR�\M�Y�NgƝ�6���#���r<ڶ��>f,ϛ�#
}�9p-���(��ņ�zv6���y��l�l��>6Q��zM�p��7z��ڴqGd
�y`�2��<€�\��ax��x�!;qa{!�]U]Q]�Q|`g+��1O�������D�=g������ M��]T"���&��<���q�P`d���hq��Z�;td���MǴ��W�lQ���g�NI�Fx�}���S���9�	<߹ψ�s8��ߢ<�������;��R�Yf)E�>�J������lU$(��"z������0 �dzg��X��(%��+)Ҙ��dM�fWĘ{�_2����Ō��v�m�v���j��>wk��ɂkA�;*���'1�5��@G��k�SI���c��A�o1�9���6#��9�B��:z��Hx��׏1@&��26LiIC�$O���"�� 1ZQ��Cp�����3M-���O�9�_��*d͔ͬ\�W{e!�!/�c���LI�����%���C���rzOcN�<�1���>ƀ�dW���4M�dO,�[�����\�<đE�_��y$�d@]d`ʞY)U��C�z�Z���Y��\�Viar��!��9����z��I��0Be�XG�+�\&\� 9E׉����u`ua�Sץ��1������Y�^����%��߻�',��L]��-OaHƧ�+'\��	cI9, �D]�8�{c��b���	��Ѵ���PY�|TJ������S��VMG�=Z��b�-���h��>5�Ƞ��!��9��	o�c�8�g�����&v�H1v/T:
��ٞ2Ѳ�Z���v+Tq���P*�*�˓F�l�M�a@��a0�n�N�}Ub�m�M�ǽf�xb���<�"�k�ǡcL�q̍�] �d���5À",Cś[�X�����4�T�YCF���r��-O���m�m�s������Z�,b*=������ʐ�f�^�xޥT� �j>{t�Ӷ�B�W���IZ8s)��)ф�tٮY4��k��Z}�&��i�l?��uz��Ǥ�!"�<il��SW���d������F~���'1iH/5��n�Z5��z��8a��2I�Ĥ�aD�׍�I=ۡ�����^�o%���6���t"�|�U���T!"��At�ͮ�u�8�^�>e%�e"ϭ�t� n3,�����"�;��h-��	�SS��Dɾ�P���x��Č��=t�W�1���?�����J@OY��ɓD��5}9�Y�g�92أs�k�b�Xe><2H��lD�}M-,a�7�b�R����'�
 �5#��PiZ�~�<�3u�����=Z7��
�-1
&�g��Uc����&X���1�*T����S
U�2l��n���^��mH��)�>���"#� �x\YV���OqXN6B����L��}^��c�p�.�����h!ɸ�jZ�Y1l�^Vn<�w�غࢤr�RrZ�+p��E����׶
���P�ŷd"�X��ڪ��̅bG���Ӑ°G�c�$1nBx�������n	9dc�F��~�����?�=C��8��X�!����u�Jb�@��oܺ�֢,��8���c�H�{�G��f�6JM��vZ�yڱ���]����(�P���f����W/㦂�DI��I�"dΎ���"��E�M{0���o���5����b�b�vʕ>O+�[�] ld��M�P�x�K(%�օ�c�g�&s��(���u6q����`��#��w�WQm[�T����eJ\���՘�cV�g��Y�o�T��'�Z�ܐ쀷}�g��{�{��a��<�B�*>R
1eg�����!���5 �8e*��B��vR��:���"����$Wi9N�y>H"�x_5���=�}EU��.�	jm.-�fѼ?H����UM��_�/��KۛhIn$I�f ���L&�LU�]=�o���d�fgg����x�yD��-TUDU�Ar��:_0"#�p�z��H� c�-�Y,^�-P'ఙ<�9n���
�C��!��F0���F�2gY�;���
őI�'�^���ŠtL�8�;�1fC�0/d�-<'x���%�g�ὲ�����0���3AVÓ. [Ԋ5'��#��'��qf&���,+�X�u{�%9/)V�6�;�����`{��J���7,taJN�s���9�F�b�K��XyD`j[��~�V��ƲN�%�W,+=�~,檎����*��ǇE(�� ��$���Eƺr3�;�x�l�p�v##����c�z6M݆��HU�۷�csZ�M�	��h�\�?<��9���h�~��{��s�J���-��� #A��~���EAC��l���h	��2�s�..0��/A���JLWc����|taʲaos̰z`����PL(6C�r�VU�áB���'�5� ����.s)!H�HQh`�iX0BA*p�Px��� ��o�����gx���$s���P���]�;;��O>��F0Ut�������X�V�$��h��jޝ{A��`���\�HJkݿ[�L�k'݀���e5��e3�%�"e�ʜ{�T?{�[�����Ơ��5���&z��4���� M%w2{j�6k�K�
#`�H\ͤ�['���	�j���#?���wa���"H�$�kI�`ֵ3�����V��;}�����7>����=Hh��z$dD�a+��β� ��<���{���Ԣ�|�}v�ms�VɫW����:OG�� �,w�N�˒�Ŵʴ��z���J�������_����FC������=�w�X�������2Z[Dh��#w�$ԇ�Bo�#�'�9,OW�k�N�Z��B��������[�����%!!�w�>z�_>;B'$��FV�ћ���ͪ��Y$Ĉp��b�G���)>˵'�}�F:-��JH�<Ú��D�u��yB���/�
x������3@ѺS<Ql�=�����r_2�T�FQHO�X��)��8S�&B������	�l�f;�ҙ�M&G,�� 38C�����VI���K͸�����U�?���O�U��L��z ��֨���4�,�,@��c���.��Z�����r4F�2Ff��KN�ΏYЖM~�n(/�%~�����F�q��"��Υ�q�k�U\/<n���{���ƌ��N���rdǒ�ws#�.��i�'d[Wv�G` N�1n��ͅ}�_���U���ug���Q)�I�uBbg�{k���ap����A�Q��{��`�!\(���z�����a�L�@2�& L�,�^��ك�y�0���ғk_�Z��o��@5�>Y��iã�u3��`b}2���!�k&�!�ҲX�Iaq�`��8�dT�߰9j�>d>ڂs�Pĥ!|e^�2GͿvG������G(о�A��aߊ8�o6�r�L2�)}B������-{_�8T*�b(����%��U!y��k�s��r������K�|��>d�:{�ó�;$Z2�_}��
G	�u�q����[L�L����n��a$����,��j�I�����m��b��p��l��
{�Jz%[G��+b�&���ȧ5� ������wB�?�����v����*����MkBF�v$n<�u'���h��{=��Q ����][��h�&h�5��Tm���M�_eװ����2O����R��o֗������HY���-GKDЛ+�ݬ���M"&I-��o犕	5q�"a��H��=v�,x�*=F����}��o#�`T��Y�Mt�#�g�I%9����^R,��3���ֿ֢:�{�2���<T�jJ^<6)����|�����VJU{^�*�Ɖ�:y�p�G�l ����`b��ڸF�� B�ģ���<���`�rl��4�TCG�A�����L��Y����_��omS�˿ڗ�-�;m���{26���;]��DK�S����
Ɵ~�IaK���ɻ!�tg��[�7߁2�Ww�\����˟��'=t"�=p?~4�$XP�7F`�\��FID�̢�?�`���{��PJz>�}L�,��q'I����T,P��m^\�i�R�;�B	g��=�A7�T���#�R��1hJC0�:MH�D\Pvu�J�p��DC������d#ʆ�t������sI"L{1I�-�"�N�eiĜПK?�� G'a�A��%�hF.#.��g��ޒRl�3�|դ�,�s��;�
���(��]wy�������^�'�<����e�=!��n}������0��(˴rYvL��4�����h��dY�h7�ϞA��k5 ��T2lA�<���t�9��@�X"�}�R��K4�<"6:��ϓ��^�J�a���z6�M��4OΔ����}���^z|0�ިxi���&c���X��ͣE���A�Ma*F��A���?�Q���o��\�A!Qf���G��z�>�`�WK�mS&�l�M��f�nZZ	��9���zXXz�0f具�֬�����`1���7�}����}#��\��,5}�Aҫh������0��\c�C���#ɫ�z�s��}@��Sr�f6�0�LN\�;+�T���,�rO9�����&/#��xm�	26\��Br��tĳ�=��*���^���̫O�w�UA4G������g�B=؋�{��;iZ+�{MY���T�H҉0
P�p�;kX�����Q�?��N�&V�0�5�UE_T!Þv;4 �v#�����{���׹�W���{Of0)ֽ�-Kj�\3�?�O->Z
ɷ-�`�y��YA�|97�1� [�x6�z��}�	b����L��A����ȧ�$W�џ~�E�����[9�!
c[Xzk���հAo]A'��Īo@|����Ĭ�g�&�н��#�l����m��~�
���:B�b�ko��h1*d��q�&>hC�TV6�h�����Ou�K6�%0n=�C���va�Z��.�n�a�-x.����wj���^�a@}�$�8	�+>����H�P����9x�^G�"�T3�u��+M��b�R��dB��W�l֧Ÿb�G�	T��`�rH��8�F���O6Y\�쭐-����R9 ��x�$�b)E�������xWX�c^j��~U|��Q졋!�yh_��B��B`��X��L��zz�L;�����?֊�8A>���D
�RBI����;�c_���*qL�2~��qo��!K�:i����C1e�o�p!��ք��(]���B�h�̵�a�H�AE�W���y���G�;m--�Co��M���'5��SΌA��Z�b���,�#p>�.O8��&�5����y��b��č  =����4X�D�+G��G7��?]{X�� �{�������VɑJ�լ���+��ēy�X��Ԣ����1O�G�4Zyƅ���������}<��0"�	F�]����:ks�V�Κ�����/�Ю]=A� B� dURBZu�{��$D"ݑ�3�,�l�(Y\�sl���hTp���mJ�����i����ŉ�p���������ʶ����,����$H�ZEVE3�@�;ͯ36�Xu^�<F�56i��+�(��8y��9ؽ�w�Dr�7��m&hX���U)9[<����/q�3̆�֖�y�Z�'���5� Ʉ�Q� �H*6�L eKY&�r?�A?�axI)��<{
�ц�#��%+�����$L�wc�j2d�<,#�<3�� *�s�-҈�.>v��Bc\Yh3���dq�������'����軛u�ǩ�.&T	��^/�/���f�>K�sQ����k�/bŶ_o�p[���C���\s-��.��� eN �S����7a��Y�����f�}	GځK] &A:�t���lG�����1���2|��b��'R���~��>�J#���#F%���%����b���_~�I���\��Ɲ�I���(JDE��_����ʵ�|��33ky�]��Pq��g��!�EW�Jل�`$�T����Ųn��c|�j[��JP�:������϶����;�� �Q��p����CD+9ן��؆��ƚ5.E��z��2���7H.E��XEUѼ쵶C�3Y��=|| ����4�=�L�ޢ���F����\��2r�l��$��d�K \^*xau�Ⱦ+��*jd���Y�f��)R'���<��E�X�gO.��U6�"�	[q,�(�Fu�u�_-�����@Q�k�zP�#�c0�ת�ޡ��G�i�Y���N�{ؙUJ�m����5����q�a�5+\����5?u��y�_�{V��uO?�9�	e/��u��V��yX��{cθ��k�s�m�t+0����^S�4eڡIݔ����*D��f؅u2�3�{����O�i��*��T6���"�Q�Niٱn��TLQ:
�l6�h�����s���a`��V?<Z�MBs���D�YZY�h�*��^jP��z Ѳq+�7�r����d=jp���v2����dC}��ԧ&Z���r��NYZV��Fgj� ��ϫ���̀m˒V�h+�����$Ðl}r�������D,�x�\Y7m�}CaC8EH@�ȋ�~� ~�Љ�� ��ג�	#0����,�*jJ{^ѹMH���BZ8�.9���#F��n����������[aa(c^ܘ���!�n��'�N~�[�P�g�v?�e��(*��u�}Tc� %��� �c탊�+���R��D��9�W�@8�2e�O=�dY%��Ic!-���Xn�Sĳ�C=Px��d{��V��kr�4�	��H1QE��J=	�Ń�:u����6���ѳk,��t��^���KT��`ت��|τN�dd#�� .�|���V�L��(�(`q�<��3ar����V2g�$&~�j#�_���"O����8�|����h�G����ߠb
�A2>&��g��g!���b^;�v�do$@�P����9�a}��Y�Bd�p���UŨ0�b7Uh�{���%�L��n(��zh��N���y5��L��Y�ރ��t��g�,��dGʓZ;����:���0�F6�d�!zDwzUTd��3��}V�H��uJ��hYt�b���ո?��O�;�u�rR�EH������9~vog��U^Z�Ғ|���e�/���1]&���i�_��%/�ڔd܇��f��<>N6�#��2����a�G n�D�s�uB��>���G���q�ބ�I[�?3,�������C-��>�3Y��io2ϰk+�B5��Jrj3v��R-'/���E��dC������oz����/	H�o̥�fr�-�j$���v"�R&+fꃈ$��-h�j���b��
s�BaV����������w��6�']\Zf*��� �\�)a��~��Z�O�X\;R��p�X��-��D���?�Y�+�"�=x���(_���	;
RyI�K��[L������������Obo��j��!+����*��1�L3V��rv�5���ʄ��B�_Ą2��*�Z���T� �-BT�	�8�%���4Y/'=;pi����B�#I���c��ڊ:c�Ζ�4�EQ:��w�*!�Eq�B&���H+_n��Ð����y�D�[���{��2�B<���`�=�.�O�GZ
	D~6����,�:@ߙώ�t�.h ��9;��)d����)�BTz�W�&\����]��y��	�R'�k������;8J�g���]VM,Y��	�͹J�@���9�{�����}�|~��K�{'@��Dh�UKMZ�~DUC���V��������z��[�ݠF�w�����U9Y���G�H׸B�4�XI��tm>�@�bq���BDsߑ��1z,�ӕ<{E��p�G��ev&5�7P�����I
T&q���"T�V�%�,,8��ꮣ��������+�Й}���mtv����[��ǜ%ƚy\u��p:���	,O��Q�����U5q���Y�Bܨ�Ž+V�ӳ�ʏ.�8�ږ��*��� �A4>�`κGX�̛7/T��P��[y�X��R�L�TP��s�	K��KaR��	Y3g��`_.��Zb�D���Z�S��ꨒR��������1�8�I�m~�3�j��=�V�9y¨�.����8N�+������@�hr6v+S�K�Z9�t��SŅ�|�4@��l�{l�W>Rr��P�~���&[f�o���j�=�~�L�d�Q��/V�=������v��r�e��0 �&3+k,������%��F�6M-�Z ��0�ota�W�|m����" �ĢءJ렚ٛ���t˾�A���&��y��*�`/=�ֱܯ���Ջ���׊H�l<�\/�YL00�d�ф�+�lo�oQ�
�u<��d�@Zf�-j�F]5����#�������h�v���
-�+;�Cc;#29h�[�n��݌�5#И�b��r����,0qr�������#�uPP(���a���F��y�0g@<�P�FT�=�b��� �k�$bł4�����TXQF�1#��� _,�-�]��I���E���V��N�:�T[9Xυ�J{�c�6ﲍK��Vj�7S�D_����49/�)g��Z{6k�B|�`���zP�=�1w�p��Ͳx[���So��s�53�ß��̣R75C�:(��! �⺪�t&�z����r�<Y�!?��YJ�P�$"�ƀTY
w�����䬭l0y�|��ni��je~��7�!&��\���a�,�ʺ�*H_i�_>O�z� �,�-��%�G�9yTK�Y}R��䕺'J�/�O?���̬(�^ܘаB��������Zg�)KE��l x)Z��Zo	-H)�@�~\	�M��F����ϕ<F�/yN��",��`�Q�m��I�=�f�%���ă쓧u��Tx����0��{��V�K���
�'��ܡ�� ����\��l����E�p�b��2��k��=���*Z�N�T����a$_A$��}�oad����=,'���!%�� d�҄��"��1���3�� 2�p*�Koeί���4�[��b�&VPr�����u�0��`E���C��ߏZ�vꬿ�������SBBܫR�lT�V�,�V�ٹL��
(�wN�#��,֐����B^�D_���4��p4V�q,S>�!L�{YҋT;@�(d@��
ȝW qR�]�;3����>�e%3-'	�=�����O�@���'�x�,���Y��I�j��߿�b����OWJ�Arz����j�K���nIW��Y�֞��H����9e(g�˗�l�WNֲ�>(���~T+�ɓ=�8ِ���Ma�)1�j��'���YX�E���jUӢ������i�����E��۷�0}����fX-�G�"=ƪ��ԪF
�M�.�5CZ�+�iu��;�Z�"HE�$�!�@%��Qh� }\��*�,YW��}"��X�tDa� � +M�Cg�I�Ғ|7F���+l��	V����
G��<��'�b�,���	�b�7�<ҫ2��}1����xNƮ�� 觰�̼�?zW�մ�;K���!�yr�;�a�P��bg�l���L`} ��Z��g/	�5*1n���,�]b�������$� Hz�G�ĬSnb��gX����Bm���Ls2�^���</����Z^Y�f�t@@{[������vU�Cb��.Td?#(L��j��yLP]�eh�8i��Z(�{Pk���}��$]o�K���7� {��8�O#CpL�Y"��"�#��m��Q��8�I+�}��tj�p�O������Ζ�V�p8���'�*Y��� ����4kN��=���%�U�rL��F��9|ڷ�%�c	����``���_�E��ב���3[�<��m-F�Ԡ��a��i<�Eݫ������v�	$�Da@j��#� Q0�	h� 3����/�0�Ue����P���y�����5�^'���Ei�RN�����T?�3찎��Aޤ̫x�浡>�L����hY|�`�,��	,�e�;K޶��q|S���V'�0���d����'���YĲ�Tϯ{�!{��wu�aE�r#Hj�J�AY�xv�ʼ�ⶵ�Dn2x� ų��R5�����v>��I��C���T�*d^�p'$0Sfo#ǳ��cL�*s�IY�'�5`aU�>6"/mK�5k�K�gf�\p�O`���2Q�q�y��Y��|B\m�Z��R�/�b�3�7fuSU�[���2�2nc7yFLʨ���?�5E��(����i�
�VWQ�b�C���^�ҽ[4�cƕ��.�:G��R �[�B�M�Ig#�xB����=����Ě����O��8Ҋ;v��B*��u=�TY�ü��<��K��#s%����=<�X}B5#���@h�X������ƦwTD{��4��̯̏(�Br���}����i�H/&�� #�Z�׍		��e�o?[���?���?�����{��aU�& wч��:;�g(��mL�і�=ښ����Y��#���Iy�hunULmI`��� ,�:��b�
D"m����u�v�<�=��F�\�
�����޹��/>��(���YX�p	�c�1|)��m�M[2�m��sYae��Hr�����w�)��&H��d*�I6����w��.��{R!	�������r �-��7��_-hV�ui�-a�
IDb�.�nr ����2��8�7�{��в��wr��A>[�3�~���K����JY,�LK2��g'�s1����h�n`�J|�]�41j��$)/�*QXr`�M=���*�����zP���,y���@nTÈZ�+�Ti���Y�����*Y�>8�R�$$�˅>�8�~���Y.w�{S�6O:�fn֤�Lw��%`S���,�����5L�����>��?�L����ɞ��`�4��T+��	�C�%������k�����_�����r��.������V!+�+灠R�A%H��l�qk2�ZMBjP2�xn��kѳ]9|Eɼ~���L���:�d8č��MdV�	�u��~���F���,��!�$>%�5Y{Ih���ū�k���s�������-�����E/}��QRN"v1Dd��^?G�Os|��ެU���O	�1xٌ�ς�7�Fzݵ6W�*H7@��Ҋ�+E�7��e���Ԁm<8#Q�[�	-Ж���ߔ:�T�8 �vk<�2�ĉQKE����'h
FuG�8���~���\R��Z)���:�@j������-���@�>, ���u��p�(�3���H�4�����B��~>c��Gk�_��J޲d��K
 ̥	���3�l�!2�����Tb�POS���;Kܦf�W�Z�J��R]�f�ǌw�K1������Dc8�rn�sT&�ׂ:�����'��L�O_��R�:@�@[�ir{X^śj��sb�O;*_�~��$��&�Z�l����4C<��'������\�6��6�v.Ժ;F��%��)��`�C4��U�]��uO���/�?T�QJh��.��0�]0?-��Hq���f/n�������� �	�/~�Dd����5Tv�C�Q	U�+	uXTB!�c��]�*�$}�T�<���m� t��f�	�2 M�,v�,�ͬ�Z`�^	⎃7�B�$�_�l,Y kdqX����)�sAO��l�=��O`��R_�$2CD;-���Gj�e#Y<l�k%�|V�ǳe����+���	�m�������B#T�ЂXH�Y�G�:����T3di�v��N��\�ܯp�� �=����~��!!J\Q����	K^��������	������'�s��|��0�*��߁��	i�十��%�� �HƪɅ�fzJ�i��?x�19������ot>>��F���^���	�,*5|%Ș��tv<�6j\����V�8cYzP/@�6��0�����'3\����YY�X�j=�s��A�70�{��L�f��gI�Y��6��e,D�����Q�B��:%z/��x��hB��9�b��#�<�Y4�b�k�(!��|��z��.Y��>�:6��"��qc��%-$b2.�L+Ӻ"�9ۂ2&$�'tm���?���,�n�k���y�E"e���AFh���ZcM"<?)�K���Q;�/����`��̢�H�;�0+%k8$�����h�T��[two��n"����O}�w��S U"|<����/�.��U�BT��|SǷ4_
*E7��h�_�i����1�f-'���<���b�/c��a�Y�V[� ^�ĉo?H��$xW�&\Ɋ��%���Vw�|�4o��V�gз�k���6�%�Oel�dԟ~jk����_vȎpI-̰��.��`@*0�`)����nҘ���#PR�*��3�ǲ��5	N���ʆ� ���d�B�UΌ�Gl��]q�*�o��O��s+r�Xt�g�E��B�,�d�d��:�]<�PJW��'~Y��R
�{�3�;W���A&�<����Q7.���2�����i�El��ؼT�tD��ܦr)�1d���pݙPe>��£���Vv�^f�ס�����	�at8�U	X��y�k�rK�ļ��-������TC���w��bN��8��h�=bb" Ξ�4��)#;&&�����CJ���_�V޼7*5��5�� ����t�g8��^�
�Q�<�1�fQr�:$�Xt#[PT�p��<�G0؛er���-TH�0��n*�����n{?htS4�PͲ�q��?�O^�Ę%�I���V2N�3#oE	��Q�(�Gt��"�0�{����!]3K��"��y6�x�������~��s�b��z���X�ۃ2~U��3Q���c���؅Ejkw�J&�/"�IS";��Q�`�[���U@�:�+lƨ��ep�ek�9�f����jz�ʂB���l���H��ݒ���Mv���+i���]V�T�d��W.Ku�;�k�0�"5A����i��,�_�%�x
�8a� #��s�~Ql+��
���0����"9�"��I�y�t����a�{�D�ڣ!�ջ��u��K�J�En9����K�2����!�晾R��g�ɉ�#As2ws���G ���Ѧ�V?J1��oTK� h����Ы��H,�w��s�AeJP��5tPGY�J�Ȩ����rZ�Pn��-Qc*���n@%�>]�X6�^�&��HΜ��B5�O�q/և� ��~��X��{���%%�;����(� ga�%xX3��?��0��G(���Ǆ���n��دG���f�XU�q��9�*�h�F&-��Y��c�]����̏�d��X��FR�	q�\٦�؋D�|2��u%/��q�&�)��&�d��I>�X�ռ�[/B�	#+ ֻM�.u8��*s�Ks\%ٛ̽�s���ѽ�x(*�����b�}s�nq����a��rGh%�	��HV_,�^^s�3�W�Ԁ��f�𴴕�]1,j�4:π�=���H����A1��@����wr�&���z��>h�ݽ!T��hH´$�1�sri�V��Jez@B���<P����o���3覑��/���b�2��n
�^��xĦ�/f]_ί��Մ��#�XX8L?��o����ަ%.�nX82&[}sZpY����(0"�Ț��)h����V�q�֬|��C ��D,K:�T�o��]f�XQ��)^Ԫ�ȶ.Q�Y2���Q�-���us[���:/��{���R�) �6��[ēiQU���./��ƣ�qߢwc��}qq��N	�_ {^fk;R�
�;��	���ppK��<��t�>�2���݋�η��d�I�v�U���Q!����x����$��L��=c��X�u���*a��O��MY�PuD�zf�Y����݁�������Tt�QK��n��pH�(�_�zR�c�Ϸ�(o5д��\/g썶=�ƒrv�rxBo-�[����N�<��~Y��5))�����'�=0��ރB�����I�D�0�~/ D������e��N�+x�dmIkB4�F�s�k�~�g���{���6���5�@5	-P��h�e��E�7�̜��X*ndҵtV�u�|W~Y��L����J[�9��[ڌ�{�0Fς�ӎ�(,L@A���Eq�倸c;z�`KR��u�m���&5�ӣ�)���o}C�yH�X�B|��a�,!.�x�՛����^�������>��G�Ӓ���?�����J�L�Z�J�;lljd9x�b���7t���Tw\�3O�@E�[;�OWwZ�i�� BF�(�%��Z(h�lɪ�;�j,h���3/�R0���&L&+�e����#�_�.H�2\�/��$l�쫯��À=o�����A���{u)պ/�5|�u4;J�S�Y�L��9c��="/�e-��ZC�{�ҠK��#`�чޚ�ɗ�#nQ�eBX�*V��s���,ހ��Q��p�F����w�6e��`1��#>�24"�^0L�<��ܵ�>DX�����N{�YL$�w@�<�6R��()�.����}$�l�d���ߕ,�,i�3�H�O�"���^�Ze�n��T��tBك��� �HA�l�b]����$A&@��I� ��KҊ��F�p��ks;��Ć���A7!S|s��*�H�`n$N"p�Z=p�p �E�m"F�D6�d#��>M0ka�
!X$҃PL���Q���V�s�
���T<�B����B������u��
����ߛ�#�M�x"`b�[�l��|-��Z��Nk�͵�����0K�m����/é�B�x���7f�����S(��6�Ξ��݁��%�{��;�{��>���J��R%Hx�\��B$x�9{6�S��������~V5�,8ם�*�;C�6����Ř��"Q:{�	�/-h⻙@��~ډA[�<X>�@x�۝{g�V�����}G�6��k��9�;m����v���3�P�s&Z�a�h�nR�����e���U�P��=DxĔId֥��g�|�;7?ڮ��!2�-
�J�&�9�ɠ 5�^�*d#p!�Y�uT�2->A/�MPA�Y����
�D��b����~7k=�Z��߾��K��%q�.�N���ɿ�WȑXdgQ0Э1��Z�w��Z jѭ�P���=?w�ś�'��VC<X��U/��%�#����|x���r��
5٬2/��ن�H��a� 2�Jx��� B�gi8&ց�1�*��bm��X-�#*�e%Ze��pԄ��,/%
�FxaB���gp���`�:����,�/
��Y;��!
�n����KWe���uʹX`�s�11�J�	g��hئ^�7���Jf0��֬�q� ��1���o4d4N�̤��R���Y(�Z᪒�%��ueB�!�?W��D�S���>R� ����X�e���+k��!�@o�֘�J�E����[\Y�42�3�ع w2ժ*a;E�!/
��d��PK$��uc��V��g��]��zx͠�[�\��8s6�GFB�hWK��2� �!Ft*V��4*.+/C�-YM8��C&��b��:��|VX^��f�t�m#���c�a�~_�q%�75CvP+��<�`"�Q6��* >>x�D&S�c$��z���5�b�ˢ)�=��XC<�[v��
&!uw�I���8ʃk�YI��3�.����+�H�M1)��/�(���Y4��ޟd�ZW���؈��m�ЋIY,LPB�Ï?�@�a���ʦ�X1yB^���X�ujfS:;(J���Ϻ1Ņ��RF��:B&yn�	U��x$�r�$q�?@I�|� d&�ӳ�^�5}�̲|'�XP֗)\q��Fd�e�h��:+~M�ݼI�X�;!��&yi��f�JI���?"�y��8۳F�����v�� ��H GA�%����gX�zn�������L�3���Q��Έ�����ep���Ef��`)c~B�U����(��i.HY�nݰ���\
s�����[����W3�c��&o'KYI�Y�&�ѱԕIS7h�f���D����#b�̑h���qP?�KI�T�!9^ٞ�rk�'��(]5Y�4g�]������j��k �5�tY�L����ĳ�`ƀm����RR'=eԊ��������W_~��̤��������/��(]��j������L�Ӄ�׿�M�.�=�tvS������$��V�b���1��b>\���,�2��ɘ����
������Y"tۊ��h3d��[�ʸnJ@�u�S������ʿ��O�?��/�T!q>A��S(� �Y�պ,�����^2G{�CZ|�	�`�;-��Ib��W�N񒂘�$k�����-R�'�T��B2�q��{k8�X�倾�KRaK`�r�y^]�]�nqxi5�ݯ�v�V�|�"�����g����|�ͭ	Pُ����ٱm�ģe\Qef �\�wo�`���F�#k:!�&n�4���x\��L�����c�n��Yc��Q=��l��r��۷V�W���Y���'?�T�'X��l�H~ =���P�|T�閛�rB��5<d�ŋOTl< ��1��˺���k ϳP���V��s/2_�'SjR��ȭR}D�7�u���:T�SJ�%����$H��-ʈ���y��2KC�eA��L�Q=Cn�l�$XŐŕFџ�M�͝������Z{�ŗ_@�[�P2��5�:��b� wИ�!O �%��1H���/�P��.`�HR�y�]�ip��6zɬ���n�7Գ�V6!���*Dr�A[�5�;�99�Y#��X�>�^��>�����:/_�%B��=(�2�L��/���)�D��:ˬ���(�kl98_fbb�-ɀ��M��T��|B[B,V;�ʜHi�h�<f��8��v��i�Ͼ�[�@��2a��C�ϻV~�|���$���A��/�|�o� T���;g&;�;:��Ԭ�s��Y'W���d��6a���M���`��{�:Y�܃0<9�3�?����=��?Q<�|�}E�턎�X��H��lu������p͊Qp�_`0��k�[mgJN��ϫ�)��P,�=VG4�����{nb�<��<�X�����v83��G��#k5��������ɧ^��D:ˣ/�q�P$����d;b��,h�¸O�������fF�ENH9Ϭ�%�:.+P���)��j9�#n��4ެB���Q7����]`)b7k�`:7f-k��BP�U���C�P�^7���i�#dn���CӮ�̍H ��W����X��v&I�.v��4�̹2� ��J��^5%%�o�ӯ������Z�(P'�7Y���MM�(�@VQc����O 濽A;�Ul�Eߧ�{�>��+,�q�)���f��&E����{�[�MJ���H3���+��z=����]�^������+3�k��M���5����bu	W.TB|���A��13�Vf<˂˿٘P1�ɝg,p������p�^��ɕ��%V����L�	����4P~���5B�=�j��PX��lց��+�ȹ���e��
�a�]f���XJ�|c�'{��r\�Pv�J�S�O�2�|�
e�K.J�����K��p�Vi�28���*H���"����K�s]J_ɇA���V�uN��x)6E#$�?���Ad ��]�X���q�e��ز���1��V��*n�T~�5���X]��U�I㹗�����k��u)�1�ԤҒ�N	�w�)~T;2Ni�F���{��_b7hLL��6{\S�y�9\��8���?��������V��<����7��'맘?D�o��)���������o:G����Z��NNj�hx��H�w;�CM{�rI{��3�+��h.�o5+y ?�HA�����@�cW��u�1>��T��l
㔌C���}��^���߮n��k���ȟ�^а�szx2rn�ɲ�b�ҢȢ֬R�I(B���^��XV-�F�^�ú�>i�I��|#b~�g�]cB��ʿU��X���²�`��݄ɽ��XF�o4_�~R�	0�UxJ�JHX�u~BՓ�{Բ�������i!{R�u����;;J��3BK
�q�Ӯg��@���,K��w֕W�{��u��h�x���d_
��
A�h.@8���|�'$��h᪌o��"�وW4�2Vv�e�����l|2⤔��aXs:m���	�H�&a�L�V�ŉR�����j�+>�F��>/�;ь�6w�%EZ�h|���A�`%k,qeVRƧ5��8e�������a�M��1����|$�5�}���F���`~XF+��)-ԮƤ�Zm[��٨���
���Z�e0��-���Y[r؍hמI	DX�� �9�UG̈u��gnƦYcp�@{����l��Ү��b��0/%�X,ƽ�5�"IC@��'*�Bv�@��u��H��mHƴ���|6-�X��2�X����-����Ck�΃���(��=��흹+�6�v�i�a�'�K�C���9�T�TN	|nM�3��H�w#��G������x�u�P,S���@'�cU��aT!)�f�OfE8�F�W(��s�=C�rR�����=E��90(Yk���>w�Y�hPˌca 2J���v��ن��Ͻ�	�hx�����i�`+�>���/>)�[�Wu��.������N�dec�Ĉ�! �
a)v�h5�(�=��S�Y��4���������Q��e|�);���/�d��D���]�B�gްYd�|�bR�8Fu%�;�� ��(0�/��F��M�q�G�G�M�����H�����"dw�=�=Íň�p���a< (oqM�-���.��j�g�S/�&����x*�=�ɗ�!@�� �!_�%��\-Huɠa�k�jX������B{��
�bG�\oΙ@ԇvŚ��̩�R��
�|��<G��x����&�Ș��ڼ�L~��k����; �5�	��;�����َΈRlbJ�b�A�4˜[`p.��p�+��S�����f�E����-�蕊�[-k���n��|�ֻ�b���rU�B���`���npV�M2�J�qL^�T�l�L&4�q���ͭ���kr��n
��-DC�!
&�),)�2�#�����O�9�V]\����&$S�L�X7R	"�d�z+H���s�V�~�ړ~o�]\�6��apl2g����O� ̪�����b7�X�V��Dٛ|)�e�E��*
��:�{Vc�`�v����:�z���&��]%��6eqx�'-�nn��G��������������cJ�.{c�gu��m�pб<M�W��M�����a͚r⊩ U0j\K�Ssw�ղ��?dϕ�\�Z�D`�ߧ�OP�nJ�3�%�*G4�[p�>��m� 6���R�p��AF�9���� -�����(��-d�'�Rn�krAK��.��m-���k�k�d�y;��b2w�3R�l�*q�iVAO�AA+��K<=	�#�h��"��;��E�F��Y���4
�_V򢰅���Ln�OaDb��^1�BMa�(2k?C�	�����h4��"P�����w;XG�@/��P��}�yfAJ+�?�Ӑ:6�r�b�K�7����� hAZݞ���\U�#�L��A3>+�$vz T�,3,�܊��lu`i(��}�Vc{F�yA���R�=�z��V*�B�z/�w}��F�4]�	��R��E�����_��#���Wak[��J\42�'lOM+w�~��J�I8��*�3����T��dr��2�K�at�dg5��0�����WR��z1��
Kĭ� �f\O��,��l��ϣ����?�l{8)Y�D��Β�dvz��@"G[A#���-^�3G�UM&�M�1�"���3i��؇u,����jB��T\�Y���u?5';'֓�������1�.�2֛��9I�e�
q��M� ��yr��B4Z.۹d�s�ZIǎ��� `\����F����3B;3�6GY�� �2Έ���8K�	60$��G��G����ix��IJ*-���$0a�ig��û8���2�u�[a��lxI
bR���x�j�ea"�Y�(����)���pH�>���� ������j�*�d�n�zD��Es<=X�e���0�97Mm\�����6!kD��3���T�
�|E
��:w���+��� �̩\�P��.!Lf�D�ԟc�zpi�����,lP��ն+;w�8h��i�]����`O��Il3z��%�4�+8�ꦡ��Yc�6�m.�j�*�uk��3ѨE�޲Ҽ���5��8�}�QgG�O�b� vw;�#A'�X��?/5N�A�ȏ�/��6����b����5.�+</�+��п�~�Z��h��]W�H)��+��Y!�<�d��2g�� �l-ޘݨ	,��K2Y�/�8%
<kOm���hk�*d9�)�#�RJF���p���z.�%5�R�L���f�F0�O>�T0!8���S#��V�e-�� �!�l�2��}��'�q�53�A{�Da����$��d����s��(�/`ot{��Xˑ��xU�,�Z�'�,��D�''���G�8�]���#�꤄�L {�Lo���v ���;+f&%�@L�2몙M�adeiʨh�!,�
x�w[\~��2�O@�"�ǧ�j#|6+��|���9e�A�\��b�wt��h&�D�#-V*�n������ŐH:�D�8[Hh4H��|v�e�kل*�[�ė�mA�)��Q��!*�ܵ���N��gzH����g��.=�ù�\�=*�&E������,Hgߗq����*������{2�c�/���;�؆A��N�2<�3����IA*<���G��E�,H8��p�I�X��	�l!������X�ZD�'~c򑷠5M�;�G�W�D�s��%�m%����{�Z� 5��/R��
ϟ4Q�Є�4�:?��['YkA
�%����͑Z��8�D(53�̒3I���(�f��jGs���BMۍ��� �b2Q�u����>x�|T.�p{��d�hѼ7�E+�<
����U�����gW6&����ǋ
�B ���պ��vv�f�I,�k�ĄEa�m7�#���-�����D���3���q��vc��AK�k]J(��Z��J:+�0א���Ikb������K�ٳ�(��/m9���uM�z��Ƀ�!_�gX��V��a̝3��?�!��et+D����=w|͡��1�Ӫ�j����H�>	Z/1#Db��iK��\h�D���r�LF�I�m��-��[+܀VΖ�����{<!F:$4�52<���݃�l�x�c�]k�&
���f;'p��S�)F,H��� Z��(]��ap@���!��-�Z��+��Al�@�7�%�6�`[��!��%�Yנ�g�b��*�:�o�`4<���Ye揙����$��4i���R��pB�b�
B�YZZ����	��jь�bt��B{#�C�������#�L>ǜ��Pc��Y/&�'$:HPc���x�!AN����u�Y��?�bY�%�W((hMRIx�
��05k8�l�@��߶\&/��T����.pS����"��P^���y��:��p8y'Z�k荒Q;z���{_�������Y2�Q!�[�5A�ѣ���.&l��ͳ�빓� k����M�z�i�l����`��~��5��b(�:�6!��F}�s#��#�?<��x�-qyэ�%ҚTeo�d�1ob�O��2b�����1}����/��/�/�������?�q�%����Ҝ�����`���"%��ڣ��8����Ԫ��C�ԯ.�6�jmM�x��]G`��v-�j�6�ט���#K*�0��\59�)��4f
E-��i�&�^�&@)�(���s����y�gGV���U��1�΋�-	��B�P7=CZ;Ʒ��!���e&���`a�h���n�������>R�{H�Z���n{�.XTqH͵���MFG�bm�;a�:ަ���d�	�.|��ܽV�����z"�##�l$|6�Ґ�ɞ$�sVg=d�b���U�%.�v1
�7��bVii��f�<����sT�Q�f�Ʌ���~����W�G)�%���oj`���u6�4�7�XlE1����|�����GŘ6�����5D�i������M���	3�T����+qϿ����e�-��ߴ$Q(Ȟ�M.6)O-�xV��'ب?`q8�f���n?��9"Nf���%7�-ښv�����R�u���-l�/܂�poL0�e�n���t ��_�\[��O�⬚t���"!B!���P�DC(�f%!�V����9�=y�Ň�2�[�OK��z����Z���(p�������R��7X�YM�hk��S�B!sֺx+&�x�}�R�?�� �h��&�U�3�Ë�x�Y��tA������g*��)S�����ka�4����`��Vl���[�q#@=��� υ�l��gB�-ƭ��E���B�*�k B����n���D��K�4��8G� l�Ҥ4��Έ�z{p��,�s(D�o�[��A�4���
�mH�����S��5���j�Jl����QZ	����������)}��	X^^d�і�s��W#�˪��pA3�	c����ƴp(0;׋^"p.�D�Iv��t����P6�M7a/�K7Y�C䥿�� �[]�^M�������h�%ǋ¤���/i�y�
C�����BEh7\����ܨ��5��h��ka腡fԏs��K*j&�5�c�\��'���ҽ�<>� L��a�H
S�JE,s�T4H3�Q#:�����'�d�<Ȱ��$iaR x|��1N*9�NJ(osvrl�0�I����;����߆?�kL2lB!��łZ8��>"��j4B��$	����]H�E�\���d�u8��/�a�DW�a8P��^U�HuN�E��e4�İB�G�D_��U^��/����"�C�Di��7��m����,ز ���������Qa�8^q�il��W���]�KƋ�TgP�g.ġ���+]�E�����E��G:+�Rh���F0o�뉣+
�� �x����������BL+.�����������j	��wZ��
o�����zR��K�"ׂC���w�[8�����Au_C\^���Y��H��p�	h��M����mU��}�"ͅ��9����� �6�S�2f���g>7�е�� �Qa	$�GuIC齿��_�65�����<o��3B]����<Z�˳�zM9���䜼��^,²n�&�S
'[��A�-��u��M�vmDW͡<����$M�WL���]{��v����55���"P�A���pp�āV�c(���b���@�q�ԝ���͵qLTS?'Q�����ʵ!]����ڞ�ϼ�<�|��5z���&r���{C:0�����t���a��°� ��j���L���*"�=���mT�Đk�����_/���}w{���e,�n��h���:b-��-:Go��\��xN���Fk�kT�FW�3y���e)1������Z6cʹ'�9��M�J53�\YNjw}f�*��5`�[W�p,~r���औ���VpvV��o~G�����k{��['u�#�3�"F����� A�?����,�(L����m�ľ��I��LK )�I�;]��e΃��_���o�����7���0����$z{*�M�D|�po�˻�j ��F�лu��~�������^�r�V�P�����Y������!�������G����E���h*�qAZ	=Bɥx�"u��Cd\6)���M���:�k�C<��{�ֱ�}�ѯ)��TP:�C�U��%<�8C&��IǓ%� �)2�f���iaqt����
��l'D���*P/H�@|On}2,���n��ˤ���W^����U\wZ�����ji��a'�,y��͡OkB���~�ן�J�R�l��p���u�1ǪS&)t�ަ�јy\�$�b�9�^���g|iKR$��P�"ݷ���d�;��o��V]i�_�\����r��fp�
d���#�:o� z��
FU\K�+��JRD����^.#Ӟ�*�n?����O�Y
�\����{^S�l`wE�	��zb&(�|�������b�"�&�-�0d��Pf�$���Y7�[Ʉo�q����f�?g!���	���`!<+��exV��u)i3$I}խw+�����{ŚY����Ą��F|-7�	�-m�9��,08�W��vG�u;C�e���ee�wo���k�?y�� �T�ҽ����a��
k��ΊϞGKmB)�E�-��O ���<���o�}8۝!�>#?K���(�;Oo���z�� �g���	F{�q�8��n��z�M�u~\zCC�b�i�u_ ��\_;��"l������2�}��% ڹ�c� �3��V�0�(��Yr�Gx�G� �%�n��$�P���W3��=W�E��� ̖B�����Z|����ul+��#*�w9�85��i�n%=+H[w��?Y�n:?�BT���p���c��q�YP�|r�㙻���0/����6���愡���n��k�[�Ʈ��
�Y���������]���Bp�{W����#�E���<g�!A��I�V���f5�;�h�Z�=���%�P�.+2f�ՓJ��m��n�!P-m�4�U���wo���7�J���{��䁻2n y*�&���k#�~�U:�F���V)�(KT�X%�M�}�6��#�@��(��ý��{1���L;�4	Y���n��K����Իn�������=��q��(ka�tx����o$�[Z�e�K~�Ί+�~![��}��#&i�e����Xi�����-��<���Q���F |�{*�th�ƹ+�����7[+�&w7)�k���[��8�# ļ���F��ϰ�d�1��_n!�u�`=��&Ɓq�ｵI�C��M�����}�Br�i}����s����"aI�_�<��A�Y�n�XN��m����PX��`hK�0kz�v!7��5��]����]���Ш����6��@��ȉ(c4ɣvw��R�.p�Hs nH�<km���jz>_0
Q�3Iݜ|��S�!�Zߵ��%ָ�[Q�}%[�I�*�t���z�C�L��m�	#į�qRu��%�$	0fηI���~1X#��6����cw�@	K�>�Pά[��8JaX�ST��/e�����""`��17sۖ���Os�U؛���8H���x���5���[B9��֩uQA�=#=�O����τ�6��=��E�dM��"?��VJ���S�?a�]����S�
�{�r�[\ؽ�����-���%�a��n�(�)�bѼ�P%Ƭ���m�r��e�[g v�}p�:S(o,���[�|���TZ1-��t3���eK._h�^�V��*绤�8�K���߿u�ʏ�ٸ�	�Ą_�/J����,��O���F�iK���ª)�[KDh����,&6��|v<��I԰�<�g;[Q��Ԓ��[I �bU�����u�(�+��oXLi_z��a����h��}������JV[Δ�}͐���J"%IJ���!�yj<Zu�&[�4��^<�<�`L��q7ɽ��'��y�>�S�Ҧ��8%Y�Ș���9TNK�}�6QP�y��Ԓ��	������ٜ�Eʉ(%V%=@~%�l'b~��Á��bf����7[�=�$���!Y����S�|�3+�kWX�y ^ؼ:˙�[�@��C����^� ����:��"�_1|@���}ٝ�ˇ�-R$4p�D�u�cx��T�	*)G���=殭�ln��N
��#yF���������=���������S;u+�a�t���1�e�?��.l[2*Z���g����a8��K֥�k[��E"A�V�R��wI�v���מ�?F>(��+V�!����+�钖�7|��R��
�Y�N Ş�O���5<�~�f�%1�_tw��Bcm��?�nO�^��Atޯ���x���>]�a�,����B�٦,\�k��8]']�nB�6��V�w�bz.҅�9�6�-n}S��aUl�� ���y"í����?'��"�ԆVNZ��v�1�!���'��Ei��FK_~�4��B4�-d�f��[�Y��s�c�v{���SR����ׯiX�����b+Lu���^���B����<j��z+��_�kӴ�au4�t��Z���g�S5�h�j��$�`@ޘ��/q������B��"��-]�Y���O�vV��պ�Z�r�jٔ�f��%�uV1�!oȬ��X�^r9����v\!����O�����rfrc��E[��v��n�������X�k����twsś,�3YM:�3\�\Vm�tqQ�܃cI��\�4(�K��X?>��m�D
��|~��X�$Q�G�ĵ�v.�W�Q�aV�PH����y,�_�D+=)u[GVp���\;s���1P�w�PW*�0�J兩����;�i�H�Uu�8�qi'���&Bi��ȃUR��8��LI��d�1$�~��Ы��<,f���)9��C�O���l�h��V��w�����R���5��p�ݚ��fhy�b����`�)��S��lx�A�K�C��h�{Av�����/�ä���w*�du������-	(ZE)��Y��~�qZ^<������6�@ݘ��ܧuǓ�r��_�=�!�脸o~]��h��w*��F��6�qʘ�s�Dh��fܤ.����;�|=�|qo`�0)h-���K��LI�۹��5����)����S��u´��u�qEjr���td��K�6�y�R��Ya$��kSh������o��#������կNBw����3N�gW�����!�qmV��8��U'm��SJ�t��@�M�qA:�c$�'�E�Ԫ�'�$B:�-٦פ��/-S^ޯM��UhӺ�+�!ֱ?9���~��`�'�����r��N�qi����͊y0\��*��?S�4a���t?Gۧ��	RdZ�ɂLe��pBh��+.?hf���A����;�(0�4B�ҿ��cU���|{Jr��ݔ>e�<�R�'j�=�\(�)�)�f�m��jnEWO
Ty�`M�K���&���l͛ݙ3����?V/��f�NA��ʳ?�rvk��W ����p�@�,\��[P6ٞt�8PZ�<��[<�Y�w
��5�Y�!԰��T8Q�otK�o�=]"���-�޾��пek<�X����-���ow%C�sI�PI�%K�VV2�x��!���Y�u�.���4(�m���_->���|�=��Ŗ�B4�Ҟ�V�u�ֲ���I��H�z9��ݷ��l��Y=�E�� ���/-n�g�c�����ڸ�u�x��Z��w^�k1�xM�n�����~�N�EK�ژ�4���}���ܧ��\�(!D)H��u���2�����u����Iy�������2����5&�F��I~MB���[z�J�	V4[?D9���qP�K����u���kSS/>��(!{L��(M�J��3�sZ�nusZL8l��U�����a���"5��� w���'�\����qa��Ǫq��İ>1#��I�m{w�����CQ��7���I�n_&�m�<��pqm��vi�a�Cދy��l�$v%T������ۥRF�Yq��˽�<�e���U��NqУO<��3��[��D�*(���t�vm����u��ͬ�|�� wQ�Cw��p�M�pZɋ',�����:����Rx�\��sa�Z�E���+��e!�E���smQg��Ù�M��r�/j���b��	���A�ܒ�$�/[,mޥ��g��O�H��,S��"�����E�J$���,{�j��5�9�DFE�"��ܵo�l^T|�����%%[m/DC��c07�ZaI�R2�2B`�����L>6>;溃m�٦c�L�ﳡ0�S�������\,��j���i����I`�DKqX�������z;Dꎉ7�bF��n�-%<n����;���c2���e�!-������N���u�?�W^���;~Q�O��ȷ�����c���,�z�=�ikN���:K"[ afY,���A�qE$Tx�)ȓl����r9�ܷ���}��ձ$�b�f��k�7N`�q;�<a�,���K=r��;��K���++y\<\�����i��|mEN�)>���~ug����}�B�_���k	�Z�1�lV���k�0�||�n	���!I`Z���gi�2]�[��pkj�xfH�NM�ckbg��,T��R:>k��6r���I��~���}��ڟ���C?&]�ӅRz��1�X9��38[v�N��\�h��y�#�J��m�,��ǥ��L��-�<�W�f����]9��w>kkݒTH����,�Ycc�VS�'�5&���b�].:7
��vM�-h*���+yM�^�i��qc��e�Q�ogE��r���>Y�or<�s3c�Q��V��b�箬8,�Du�^��Ỿ��R�ӗџ��I��{�ſE���C}������;})W�������DQ"u%���Ȑ�d�*)tIl��tV�v`�1��	v�K!z�:ޮ�ż���0�v���9��z�R�O���qq.S�T�f�Iıq�X;w�2$@��#FW_aq|���%�����������"m����,/�l�/���[���+�\�Z?�5</((��:�F@��Յ�t�zi�1����`Y�X�pH´nƷ�Ʀ�J�҃��u!ƹn` ��ir��]���q���:���j,Z�1��㷛��jZU���tm���L%K4�-I��:TXyqk��B���Ic��ֹ��0�Y��Ć���p�A}:(;Ko�lg�m�}�N��&�u��u_�X����Ւ5��3˗,�N�]�<������v���j≬}�3�V��~c�C%w���~����i[v��d���0�/w��0�	�,L��	�NX�$H7{�ZLۓ:i�n-Ү��!�^���u1�����__���V�W���4Ǽ��˂8�B� '�(~��%�����E�}m�[o�ør��r8�^�m�)��|����|Y�&��J����
��kI{B�:ۈhr�P
�cI-ea)�bK	�5KEL����r-�Х��Wo�_�o[��IB�2S\p
��j��[q~W*EQ�ll�^�0>3�Eg��Ǳ�
������h����+[&&ٺ�eC���a��s31���o��k���M�����Z��&�j�Lŷ�zX��m:� �����}��6��Xp�I����k���T̽��b/Ș5Q�J��J,e�[��[Ӆg����!>���!9��2��[oT��Uf�E�>ځ3[�I�of�?'���a�9��L�����J������g����k�:1� ���{6��q��\yI�1^r�;L\QfIK�Mփ��65^��ݮ��~x"�����f����zw+���?�彳`��P�za/D�s�s����������!�_�����VO]�G��ʢ�m�P��j�+��H]�B�v���*�!����6��5����^l��i����ic$��^v]���t��\Q���V�@ɦ�%7İ���v[�XZ�8]@�9�GJ�A˓k��](�˳���Y��ޜ�팴M(D�H�Y-�r!L��U�q.�3y�r��a��M����^�	<h��B}���5I�����{�dAJ!�f~����r���B��P��O�����f����6�m��b�C�ܪ`�J����.6$�z��ݿ�m��{�x��т���'g(�7F�6����6?��__�6B�ʥF��S>9և&
�L(�p'�3�_ 䨿/[�����̷d���u+H�)��x�n�%k����Y-��%�&��a��ܤt)DH�+E-e���*n�&�`�:�	>9��D�5V0�D�Ō������N~?��0�s5�\p�D�/&z��ox�Ͻ<��~���O.[%�s�I�/m�p��t���+�l����[����Ȓ��;�8�����ZZ��/�ŵ�ۡ���3�L
p�H
���7Xt�j	\��M�ʍ��Au!J�(���\���.!_C�ۜfM�{�N��R���B�Sم��-ǔ9�[!��$��nt'hZqNLޏV\ý�P{�Y'^������P�;&pMh�a��9W�ׁ�K������3Յv����9�4�y��B0Ϸ�Gz6��?k��<Oc��t��p����A���ds�^&t�T��
�笵2(���/�D7��Ğ�9�'�}�5h������4�k-��59���g���|ie���v#`�5o�w}��R��H^�� �n陂�2u:A	��������/{��¼�ul������][�t#w7d�C����.m�.f�l% ��\���� <����۹�J0Lm-8�ݵ��F��8:���*Y��r�����y�e"b�C�R�_�I� S\�;��3t- `}n��z�����s��P6��gb~��K_W��X%�z����♙�c�_����Tz���.ν�b��m���ykj���6@����q�S}��M@���Ak=��W�aN���8�s���E���k��:�{�:�\��,̻�l�B����ac�O1�R����|?�Q�1�yp}?P1˾� ex�|��b�4������RP��Li̍�F�׌)i/HC����aQhL*L����M��i��?
jZ�҈���$�пG����7�~㤂a*s=�r6��$��k��GO�kL�iO�%�qު:%u�N�Q��T�&�{K&���-�S�z#�
J�^K_=H��/-�x1(�& 0}�L��p��X�9�u*�bB�2���'߭@]||o�bW��/�W�9�fA{�.Zy��k�� R�%!��讏��<�_!X��L�(�f�\���w]g����i��#t�����wm)���7�Y;�0,X�hlX�ǔc����|D�C����ެ�|��]�~^������M��Ú�$���6B�Z��?��F��l�~�*�����1Hդ��b�q�)݈���-j����4{;z��˽��m���,Rlt��"�ԛ���H�J�i�0�p�p����&>�K��<iF԰F���0��w�a��#�:l�j�X3�~�E��q7M�KyN[*ڣa��ɉox��p[bc�U7-*��l<9�#���a]��"�`�iU�8.b09Ⓗw�BR���^�k���7>)�R��:/w� ]g���ѐ�Б�ϫR�8j-	r������}�DV
�iA���	���=� �j�Ε��>-��=t��B+>�\ׂ��i��ZW��т%����<;l~>�]�=��^����%������b�&<0�����P��g0�C�W-Q0b�t8g|�E�'����9�=���ޑϟU	��w���2�U�2�Ie��1=��ߛ���!� �4��f2��Q��b�L���B3��H��dS�����v.���P$X��6�bjrs=c\JG.l+�����@�T7�Xn�P Bi%+�DN��o��IK��،/X�� ZH�T�,���N�����, q��g�5Y�ys�o���b{�G���f=)4�dt�U&nּ5j��<�)3 3�����g(��roʩ���q��Ly�r̹��J�A�����x~U������rx��xx�?��
� �B�;�I
O�cd��{�����l��@��)��֝��!|�J�s��R����y,N�>S���6��(I�3iz�nQ6D '�g��d�*�΄��k��ܢ��9�H�WV�n�|ћ��a����N����-��$*,&"Jb��0���C��j��0�S��$�ݗe��bN�d|�d����~��|pC����Ĥ�6b�ɡ����#�N�IU:��QK�W��)�%*�B���!⳨�ƹ�{�J��a>�Ε;��ٞx��ђ�1�T�q�m�����[i�!�m�dj~0��W��V�rN�>�sţ���[e�9��zc�J�/vó�o�,�.g�k�F���Q�a/ip7sR|�B!�1G5a���YvM�خ�@���اW<�{���
 ���|�!Lq���M�6��p���+�a�u�v?\�����V+y4�FK֫�u������y���n,����is$I�,h�GD�̣���fEFd������ٞ�#�q��=W 
��YU=-��"�p�(
s������R���hǞø���up�^�&Q�f�+y#��а���l1��W�I������@�{���!���Y�x��O��&v�Wl�h���t�3-����FŒI�dz�\�az�p�Ս5��j�j��*��5��h�޲������έ�w�z��E�.<Vz�������7C��rO�Ets���{}�l�Q�t���5^<M����\?_`{�w��_�����r[:.���K��X���6,�&Ԑ�;�Զ��/2oM5���<�ͨ���
=�>����hܣ��m0�j��u\{�`]����P��)8���'��=�
�U����h��T����`�r�u���}����mY�xT���P������M~�d>�rD�v
i�)oO�6�����Qjr�c3%���b�������x��;C��G�e�X[?��'�>[ܛ�j�稗�IXH�̇��k���-	W�s��^fw ��`ה�M�t��+���"��"a��"灇[bY|���I�=��A����8���o].�d���Ȳ��iƷ�T�w�U��U����[���9�y�{�ĿG��Z���o�q��t#eߝVV,�X�r.n�w�%��-�L�?2�����}*}�L�m%���Ɗ�s�Դg�0���l�IR{�m�=Ri��KG�&j��{����3Ȩj�������$_8�������2E����"Ch�N��	��NM�Ƙ���o�N�k՛�	%0ѥ�S��x��I��J�c.�j	�V� �]����Rx�p�k������gb[O�h0>��ǛP�׼ 	_���'�y�Wc8�s�j�)�*���p�z8Fp_Ǐ�"��6a>����^W��C���W0�Ϻ�҄�a��f�L���u��1�����H~����㗚9��nz#��p�<.����4��a����_�r9�y��dcd��ƺ}����H�u3���Ҽ/��dQ�0��
�
`I�hF�!���k�<��g6n���`���:Qa����9��~��x�)`:y�I��}d>��J��wb�;���=1Û��W'0���9iHڦ0��H�R�Vq3LLd�5�[�h;{g����Bǎ����݆�'#'��t�jo��x��N�f4�5]���7�X����P��U#�d�q͎V����J���z�FF���������Ch� �f����ލ��s^,�c;��Z>�yN{�S��mc��ĴZC���C����#��5t�V�(�H"Ft���0O��(����Gnj��θe����U9�y<�'?������a��~�scw�A-��㭅cza�l��Q�=�ŝ'�e��&�cz�;iZ���,_kJ~�-��U'���ϓRH�ǁd{�n;��;[��R�U�8�>�|�v^k�4����u��ۊ�>M������27?%Swm��!*�5	��E����K?A~�����\'~g�����������V�<�G3<pH�_�d])ah(�~dѭj��� ִ�J�����'�<�f`;3���/å�y�`l����-zb���f�O�|pѦо�WSk�M�ළ��ɆԎ �Ӝ1֪�o�y���\�T�c28#"��ݫ�mi��ܰ���C5~���>�a>�k��<�H+���t�3e��Q�i�	��d��
�ǐ���y�@Ư����T���׶j����T��dL����� 
�j��>�86˜�Q{X�^�b�"�z4U� ��K�����N���qW�g�R��ww�+0���kyy=ˀ�ܮ5��;��2�pBj���x*����+����/(��x:V��8�����/2�([	q��yNѲ�m�=�&cYo�p���Y��q�^��&UCf]�8ݝ�����;o��D�-n���Pŋ�����k��R�R5�=Y`��h�݈��߹S��VPQYXaT��ZhW������bE���t�z)w�q�'���{���}ib)�Y�^��I�M�;~l��^�/c��`�D�#0{�`	0�f;�y�H+�i-���F�v�z$�ء�m%A��N�ӂ�8������+9'�����<��Ś7�k�j2�y�Ѡ;c�h�Afw����G:p��b�1�Q��Y�[9�/���7Y�>�� ���C��V_|�v�]��P�f�����,ľw�׭1�䍲e���1)݀صv�8MX�ًI\�z1JТ�{0��N��ha�$7���=P߽�̣,o�j)^J��>r_0��a����� ϯ��i��#è�(h���P��`n��(�x_�x�~͌B6;t�w�Ig�E�+Ƕ���=�\ڗ�������&�TcX� '��6km�[x�o�����0��}y�}1�SZ���8���%ъ��;�����ی�~��z���%:hMG�=�5��_ܰ��D�ƙ��\�<L~/kw���d�~f��ܯ��<�"p�A�;��`�yBRP���3-�<�����|>�o����v��E�ԐN>e11�RJ���>��j��^� ����H���G*���A��d�Rո�ܒ�qf|GU��X��q��}�N�&)m�!��R�E>on�#�@)���f���Is��*=�|�;Ν�H�!�]T!:6��M�573�BV�?�#,�a�E��+���7D���;K7�7�a	o"��z��nz�/o�LM��ae�5�B?>�4Σy�摒�>K��������tާT���~���2��1���.�F�օ�lcU:�?������#8hr8��^.�r�^�7Y�R�m����d��ì	�:{gL$Ҹ�"~�c�(��Z�i���Bb��lD��&����GzΓ%s8�z�~&�+7Ӄ��g���4<�ͽc<��nv��1��@���p+A����nz��HI^71g޽��%rc�Q��/ylQ���?^�]R�~`���4�ؼ����uP�X���Y�-Y�dh�d!����2�֒w�)����1y��a8�[d/���ƞ�9����%R��wx�ك�7�ȳ�q�J󱩴,<He3��4ݓ�WR`����y��Y��&*?����g4��8���Lj��� @7.\��#s�BN��\S�zDX�V�o�2)<X��H���?��J<yJ+��Y}C/�������aWLN�{�Ѓ$�	�p���=�E<�)�@�=Zۛ����Mi����l�� �k-���P��2Y�{�����B�h'/@�ƛ�]�����5�����Ʊ;��o�L�E.o=��PLp���=.r��sՊ��T�--<���z��5G4>��9�98I���7��d��H���pU%���"c�wo:P:1��O�ӜS&C��j��Ox@�9��{
�Ժ$�[�&u�kl�L�Q�J�u��*rĈl��d6ݘ�1��W␠A��ܢH#<��g��z+Xn�b����8/j�K��,���Ui��kڄ�>߀7��:o����o�7s��z��Jr�Vh3�B�K���fQ�x���l޶�������	�P�}K��������c�헭+̹}��߅8u�����[T��[C�F�����.�g(�n��5�nHØ��F�V�7u��`}G��A�8Yt�	�)wS*3uO�C]D[5����ڝ>�~6u,��"'B�6X�`�.�A}�8H�	��ͷ�8���v/�U%q�0��ǘ�'��F���`0 �e�6VH�q�ym���p'̪�����$�3����H�\���%iJd��Qb%�H:�:E�&�6�HhrR%djHk6�QeC�ϷЫ5�k�Ʉƹ��t馓R���D��rc��1]k7��!�0�о��q����m��r��xj��Λt��zc�9��go�d��6�����{Cnr�
$�Z�ļ�AE����N�Tɭf���qJ4ɁND�����1�s�kU+�v~�G(��7r��t%ɵ�`�R��"��L��V�1->�tq�JO�'��:,� �1���ry�څ�#=J�Җ6���?}�W�T�l���&]��<���n%�u�|���H6��sTC�
�&�������'�	�L�=8�c
�~��-p�tU�1XU1�|O�w1`������q
;Bi���wg�5�wa�m�4
�$�u��j��,���&�N����W9P�6�.SF�x3.d
�=3�Z6���lC�|�1�H+���f�Z�c����hq3��M/�jl=������Glt�v5N���i2B_5�I�%���ޛ��ȇd������'�e����~}�X�C;�;ʪp�;Ҷ�gq��"���%�b{!{eY�P�'�-"��X8����J��ݵ� _��:3vH$Cl�L��ր��<0���E&�浓~r����E@3�wS����C����\�"��h�7n��0�dd���Y�<���(�Z[tb�b7Ő��'4�ܦ���`�@�I^��p]���ɯI��YP��I�Z
3�h�����1(�
��*2&5�8��HqAf-6c��bx*����Q޴�ދ�{x�)t�����
�7x����5���}�Z����m~��qv�e޷{�o�¿%OH�1U=�n=��u4�3%Ⴑ0r=�OR9�5C��ᑾY��+퓌"b\�=��9�g�L���ҭ:*�J_�����x	cB�f�9�!�AU��u��t)��bʊ���%��@�b�c5왏kp��X�)´�K\�i.|>�0�q�17Cr�a��e$�S� h�[�t��.P=�U,Pή6)�G��!�U�Q�U�v��z"s�<5.��,�u������[EGe����z�P�м�����4�w%�?��z��k�HxKf�0jY��OI$E�3�PaHn�m�s%����PNB�^��ol����c��u�rX'*)$j,7�<O��o�	�j�9?���w�'�/|�Ͻ����2���[_��8vy��n�)B��2T�4h 6���!L�p���p��dl�|j܂M�_s�g�1[��|��}O���Z1�01p��5AHE��"2���['�4n��B�x��[��>�rO��C�����#�7�P��*�o&>Ұ�%@]��!��Uj�등��KBGX�i�y���<RN$���$�w��>כ�Иxn �J�/xx(���؉Q~4�\��4����)C,�T�hf���8@SO"�1�vJE�ND�(�-4� ����c9���u.7�\g��F���,��c�O�I8-(��\M�K��j	��O�b�y����m.n>>�Jݿ��8�{P�1N� 6���o<]0�Zx�#�DSa���z�>�{��*{�\�������8�`�Y�R|ml��.c9�a��������1������e�I��k��g-�%�G�=o��b��7��A���p
�TC�M�z9_��`��PU,P�~=�-��i!s2����pf�X�m��u�{��5��)m�����*��^������g�qX�|=E`�6G^D��S\S����,EEџ�n��7}ǐ�Ɣ:I6�VȻ�����i����M���!17�P
3}��I�_|v���Q|j��Z:������	5i��a�/������V�� �}�n�T�W'�y�X��C!_�)����*k��yo#���m%yڴ7��2��޸nK�;CԦ���jrЉ:�ag3�H�Z��c��m��i�R���i+�ޗ=����!������[���|�3���ւd���Wu����e��T�l�E+h*-�{4��C��.����������x�#����Z:`���*c�E�q��1���"048��L&��9��C�ܟ>����$7��'0~��s�ڝl�٠m����G��\�Ԯ�Q�Tf-����0������y���m>���!�C?E�i��(	MM)��	B>�OR(b���۶D�/���S�T�eqT�	�t32Ђy��#�n}L���l^��M����	�V��O+���$�4q�����j-�:F������'�}�|����kzH�0J�Zk3����ń�n:Q����Jx�@6�:�]���W�Y�p�$	G};m��(�MC:��9��S��}=uV.>���iM���X[�Y;�l��M6o���Ynn�B�B-ئE'�q�)�5醻�"!|-[�:r.�2HZ�wj����e%���B���	�s8L�U[��][���F�����W�qwh`�B�dd^����Z�F������{/f�E��eI{���Ң#��\]BѬ��w�6�j��uɞ��.�I��f����:�mҍs6��i�	c��������g�c�ݔpIg��p������mT6�]k�!p���&M<��~������s<���h�F�"�(A�H�s.}!�P"d��+���[�ߘ �o��Q��#W��,c)�m��u�F
[��a4V鸯��Y�1�Q��״H�����h�g��G
��u�ʵ.Q�UM�l����-=oFFEľ�7#���Fm�)��v]�aY1���L �[��7�%/�<�:��c�Qϖ�=�X3��q�m���O�y�6���\�l�ч:0�0��!��O^dA���k�YBWx���?=<�ǇG1�Z�t���ÿ֋z�X�K��'*�N���71��Ċ�~�������)j]��6�)Y�k�&���"���1撠�� ������u������T��Q���/p����Y]M7us�I��~]���z_��Mx(R����o�4�sS�����W�@)yD�}�A_�<(��W%qrh\�)�e�w�V솊Ey*�h��U'�
��S![%s~S�D�>�w�<t�����V�o~A��N�DR�Ę��o��v��l ���"�h�d]���'Ch �s�pz-50g���j2l�8���(y�׽�͍�!����(̀I������ox5�7E5d��։&��1��\9��Pq�Y��C�����LOQ�n1�-`�*e�V�����9f���\�4n-y�=v�]�l3r#�������y>���nH�$�G��g��.9���t:����EئhS<�ٸ7�?w|Y:�}׭0<��ë�)��H�u��:�a�'yL��^6�	��{B���ɫ�l	����)Zm�!];�?��Ѵ���j6m)l��:P�n��M�`v	t��08������o�u,Dnx9rN"��kv��Z�a��/�K���\�wߞrb�	p�D���͡n����L���4x|,�?��Fy*1�4���ކ�<�O'�Xs�{�i�_�h	2ҿԫX=�u��Ĥl�/�,-ص����?�<t��ɹ!}lH�C�_��Z�9���[��L���ǋ�=NɅ�#"�2�V����6�蠟��=l��W��z�gO����D"�?�BӬ�Pi[��G"�Gx��ON3�Dq;���í�vÄ��1�W��%r��^+����`y����=�o��������[5�Ֆ�PWp��J]{���i?Dp�2��LʻwO�0�����(��h!}���A�Ks���~NQ��tYR翪T��I��Q�z�ɒ�5	��m���}�:�B�(�1X��h�n�!��<���t�:��$lc����?/�.ɵmq�ژi����^0�%�򊐫w�}+�8�8��݂�ZKN��S��i"(>'���11��Z�jFv��C:F�αɎf��5h��m%nv����r��6Y�Rh��A�xX-^�4��@�v��*R��Sϰ��[K�wx�6V��>�C=<��tٴ	�7���go��1O�ؠ�jIj�[��қԝ��� ͞,�3�3_1���z棆泊�݈�o���b�Z�p�Ί���|PĘ�w]c���*���0�`��'�$Kn4@����� ><e������\^ϯrZm�wUq�pH�)Q��=X�Vɕ��0~�yO�$<Xї��;����Y\hH���<�Y�xuP$�/q*�r7��b��ςk.s�;U*s�&3
�]6[ t�����T���v?�n���*�� ��/f�.G�q�����r)����^bb��E� ��� \~u�h"����)������� ��'>8\���Ky}}�n�Ѕ�Un��{����]v�w�qc8�U���ls�%0�[?Q���ϼ����U�k[;cPn�*k�{L;��t��*N������+�@�u�4��Wk��mo��޳T�}s|8��X)�!���S���S�98��f��u]5��#��p�D C��/�C�=X�x4���Eݯ\o��R�	�c���6��{�6�Q���Z��`��Q�߇�Q����_�hJ�==�ǧw�Ib���|��y~ѽp�:l�kWC� F�TK8�Y�$D�SV��XGeg�J=r��ޖN�K��Ѕ-Ns��v��ƴ$�I+��9�)%&%y"v�$8q[��ٓ,��>4RX�I�ٵ��g3̫W)�7�gcS(�xG�d���-<�������3l�&�d��A���nt��C�\ݱ�dZA�1kzeOO��d��.�$}��Zܐ�"e�e�d�mkγ�LC6�\����q�!�Rb,�œz�*�!NwB���E�0
a?cc���H��0�!��҈F��p9G>D�){��N��-4��A4rJ�jQ������F�!V��%'S�f�0�����W�A��(I�ꡋk9��bL��S狀q��$]v�H'��a�!&s<z�?�Q�b��j�N�����Hk�������q���MUClN�x����`ى����;M��8��{�u^���~/���L�Z�f�iH�C��'�!����dУ8�i���A�|��x<�$
��BaL���t��K\ļSV�IW���(��А
=����U�Adr%�D?n3����&��&�8�B��և^Y�0�0x�R��M~
4rT�h�?���U<��݋TC��1X��G/����-|r�iT��%+�U�A�I�aBY!W��A�����Ɍ���$�!o_���Q7R�/��׵q��P��N�����R7��L-aM���ᘻ�:~�b^ø�G�����6��+Ly��y��<�A�.'{�}��,�j�{�!'O�;z���1��6���a��n\/��`��7�������;y�˾>��A�Yts8�-�I܇�5��I0|vvbdm""�(�бT1�e��9=�v�q3�_2X�d5(AԬ|]�>�(���_�e���
�����>��-G�.`�bF"mo�^��3bqb >}����?1h�V�����<~�=�0�������}(�?|�A{y~1
�R�a��)���BL��ӹ�	I����mnɐbR�*�O��w[nI`��KlDCBٻE��p���U嫄�� $���E�0�O�w���������^���˳�%�3�ٸ~Ś��c>}��U�c4#�58T��iEq����|^��F��?㤪N�!%6�B�}s��8��z��6����Q�s�`�o,6-H�vx�H���b<}�G�}R����m�,v0h�U ��24){p�+;֝rS��@��	.�W��bv�dQ�L�G��G��_�e�Z~۟0,�������d���^����*c��O?���姿�$k�����|����vu� ���[e�æ#�Ӈ���ֽ����k�Y�f��}b�;�{x�N��k��k{���������lZ:��8�:�s�v��~����b��#->G>g-B���} �z�	l���?���~�������ʏ?*xm2�lO���O?�(#���r��<�{ŀ��|T,�h,ojݙ�!h͊2�v�Ԟ�}�#eA��&���� $7r��s�Q3��}��ޞ�����o�ʷ�����lsߔ޾	���'K��O�>��O̛(����i��wb�_6����b��C�oz���p���y^��l�{)��SO��z�0j�lph�@��+��5��??�:U�b�sz8������w!�����G�أ�֞�A��"��{��`�8`73^HhH��oV?Y�S����Ō�Ѱ�l,e-,#=��*!�a{R�&�ڮ��s�1ߎ=����G��3��Z\���ע����c�����������|��ɮ?}��B8O���dH�PgF\��;��!�l :o<<?�"x0���@D���"�I������U��{���2R�_�G���2�He��4.����c��V�I"����#c$UtR�2N.6���]=�OHÞ[y��,�m��������ᓉ-t�LT6���jwxf��]��X��^)FoUѲ:>祥�:
D��.*X2�G���!8g�X�3��aS_�
�`��A��$Ԥa��ћ�:̂'�x�%ޝan�v��V5R�/�R���H={r�
7Rº��M�4�^��7@5�kZX��9�`qÃ'hF�l�2�Ԓc̩
M�����`쿻�F���AhH�`��s�#S���4�LFn�mrLp��-�Gy��p�/q/>�C�@։ϛ���e*��"[�ZsBb�H(�����U���c���
�~4x^����u��gK\\�>� u�������r�R4��!�F�"Z��c��%AŽDF�x���*s�j2�N�t����ԦUpឍ����=T*��UǠ�a���M�Ի�3���Ih�Ϟ���!���?5���:�<U�.�S����<������������+p���\r��:Tz0C:	cݗ�S���.�-e2�|
>ʤ�]�)�u�[bߑ=D|��R�9�r<�e=��NQ�G�b'j��3�a��$`O,P	���w"�y|��8h��Ռ؋Q���r�=V�(���\��)��*�ϖ0*�F]"�J�_��t��p����]�ȵ�3��y`(�&^Z�nHcQ��x�����E�Xly�]�BJrjRc�愣��-�_�rDMa,�,fx�:d5��n���7j�����9�[Gwn��G޼�f���ݷ���T�������<��E�ȋ997�b~�T��5����8@��m�9���!�i�Q>��aH/J]�=v!�9N�e�ZU|Em�;&y��J�E�๪NK��Mvג�;J$L���%�]��{�?1�A���ΒC�p�|���똹�T�U���u�_^�5�b� �(�
���!E-q2���g�h�S�yO�*L!8^b	8md�ODl]Y^K�a�/���`6��'�F2-k��O:|�p�C=��&�&�N^����F0�݀b|x��]��_������>��J�b��RbV�*���!�iqc��?��m���(���qS�_������ �������|�E��Fr+�/q�th�#e#��5&���:�����7)�I<(=��(i�<��+Q�Jg��lГk�g�Yb#�Ԩd�ݥ!]Yqe�ˆq���נF���H�,f��+ƪkkp�e3C~�7�c!I�@o_�}-�y���kt��=�Ed�5����񮁙ʠV3�e�>��'P�0��9hԛ����z8=zv&�/��Y~'���8����_#I�'�	�O�R�CS���s�J�=��dG��l��Q���N%H
��/)a�
���'���̗�(_�K��b$N��n�?�e��c�Q@�$�d�*߮��?�MM�d���XӶ�)\e9+{��*�=ı�hW�H,vꍗɿO.��XV�dց�	�&	>p���z�������P7��G��Ȯ�m�n�R���)Q� �J�_öJ����9����n497��3�{xx�J�^�Qw��9�lw��I��}����9n��W.�u��dΩq��6c0�S#�E�݌��ǝ����b�r2)�O��m5�{�l�l���b��>:�c��+�����*�����E�&*m3���=�,������/��
a��/e5���E�A4����[U��ƍ|Z|Da����a��sX�pp:<��iV\y�<���c�3�,ɻ�������_��:��\�DL���~~�#m�O���67��w<�7i��G��۽�ڂ��fx�U.�Nh؅�篂���b!�bL�=�t2;9�.dbD�au�!q� �U>�L^�nY��I�S��D����I����F�F���c7i���MZO��J�������sx"�E>�ܷ!�T�),���i�!T�b]LX�Nr�~�^���BX��_�xtWgxʦ%�D|�m�`��Hn�]q�n*���լ�x���#�K&��A�Xj��f��<@�\Z����u���d��v���TIB���&LpЈWvVO���>g���S}����7�MiDy�I�q�z��-2/8�����I�FAK������j��8������G��j61���4z�I"7!ѻP�y��,��97����e������^4���If�x��ι	�#�P~�&:D����H��<�֭�d�����7�z���d�5.�$#�i-4��]�x��i��Ž*�d��=��@��F�P�[�|�O�|���q�M09�M�{�a,6!L��Ⱥc���7�-o�L�r�y���r(��x�-YiZ�������ӧ�f�aV�|�r��h@�4M��`¾Bl�1��y�-��U�V	�$�k�C�d�?~�Pϯj���F�Ϙ��ō䇌�E>G<=;X�y���0�k�9ε���!MۡX�Or���,�=$�F���o4��Ҏ�&_�	���v��y8�a�
����'r&mb-m����pzsMMf݈J�
<=�=b�#K�1ڿ���"����4����� ��7��6���2O]�L+*�"J[�(Q�?F,ǣ��T����T\��/�3We8M�mƞ��B)E��<8�z�NL.�$^�{�k"�>h�j2�F�  ��IDAT(�aQ���#�!������H��rL�p��\F�L1|���T��U�q�-N�%Q������1����Rb�F�q�s�&�z��04�ѱ���y�Y؃O�
�0mf��\I��]�=�v�l��Žϩ�"?�;L�_�;���/��ɸ�g�J�!��T�G�G�S�FL>�F��W�tU�ep5��0���q�ظ-㎃I����q ��^@),�����Y���Q�\��BGA�m`I�����l`1��u���V�UÛb�P�ƑBgH��� �g��5���9�R��2��ݶÔ49`��A��t:(F�q8��܍�վOp���Y����n�%��͍>d���Ðխ��rb&�nr��ƙ&�	5��>A�-���{gd�0�e���d\Y٨����OX����I�~�a��-�DƋ��\N���k]����S���P��L"؊�!=4�j�7v��Ho4;��5�#M��w��?N6�"���la[VDl���C	�b(��ms-KO`,���*�?}*����S�O�0�!����I��O�5��6�]u{��n���y��}���ӫ&v�0��l��92A�;�:<��s��u�
��d.�� o�J���\O�E�\FjP�7uUM��#�<*�G#�8h�A��ɥ�X�"47��}�0����I>�+¸�_?�������`����p7��vik�Ս-������������7$����s�+~����XIfj�Kc�;���<t{�D�Èk��sN\�<���5T;�q�/��}�9�p��|G%��
���$en�1�	mK�HBN|�R���d~����Zx�x/H�R׾�7�*Q"��
%����Za�j�bo B¾�'
c-9�w����4y�#Bv�l��B�ª��~�m_K_���OO��8��� [�KC��
�������|Pxg��xs���4Ҁ�K���5�Ӭ���W�w���b��?#B�\�����?�s�ր���������2���f���M���d��.�ѝ�/w�=ޕ��M�l��%{.Y�W3�f������p����q�-�Q�adH#Vc���j/z�P�/�X3��4�G���ٱPO�䲬�ү4�/6<�Փ��Pl�]�c�da?I(�y�>��,?��6��_�(��L~�hFH�����LmL�_�s:��Yq�bz�c1>�@�b�������_ZoD�v,y�qW�8j��g��zY|8��ϳ6;��%x�0x�V���V�&W%�@Ė��;i>�(�{���t;� �����7�}����zR�m�T��~���y_��0�r ��Df[��h$�f�����X��
皑��d����vu�'�>TQ}��rgA+�(b�'>�
n��$��'ג��>&W��`aJ���@&�)�N��'����E�Tk���j��چ�Q)5Q���H]{���֖������c��ݐ���G��U�^��?ݳ��j%�����g駏�7S�@�������q��7*���mS����3�s
�O÷?��Η��R<%udu�e���)4*����^����g�����>_d�iS!�K��܈��?}�h/�{�4⯬�ޯS��}��#uQ+�ݪ^�E����]�����wØ~e�������I5�;)	��U�	�S�CP9�7�-�G��D�R�Q`�f�!顶n�f�b�ɀ�]���deV�>sd��-���FeN�F�{�Rا'�`�P�bt9� |qD��IAX�����xW���?�u��g��RR$�=Fy+[��d�GoU=��~��za8�+|2.2�M����<�sk҉X<�ZH��}� \�1nl�E4��w�Ϗ�[&V��kP����!�=��n����K^����'O/I��Bt�@i)�^,2����[��@�B�y�����$���#���Ӎ�!�	'���7������O팧:�g��j�#^�>��8�f��!<M�Dm:��ƶV*w��WJ<2��9����t{,T�"��D��!n�9�u�'8�������a�F�����E|�8�Խ�b<�f5�v xv��(�*�*�*u���fI�Cx���R<H�����i�V�yS��n��c"���嶣	
J(�u�C7r&aD?��Qx����(��i޽)�|�����U��%���&�Q9�jH7����.a�x���%�O�u��\�Z���i��)Ҋe���~�\/J�y|2q���֮ςJ�r���G�N�������ua����t|V��,���eJ"��L�R��T��X�,�(�L��I\��M֩e����[<	����V�͞�А��(�9��E�M�d���a�Ae�>��^��l�G8�,�F%ԇ�zh�~�)������͇�����{������=��Y8�?�?��*��ɒ5*ް�������s��b�%iY�Z��C��x���Ԑ6�cB�N�3k�'%��q*������"��SH0aS���ּ�3�_��<[�':N�&�p�_>�*���P�=sêR�R��+�QN�Q�s��K����a�7j�0��$�?j��%8&��{��^��V*��&C�,Y� ՛��س�4����Ud�?��IgdPђ����>X�IK�:�嵑��qL�s턈�s<�\�*'�a�5��=I�u�p�
�7�ֿ7�5����d8�0 w����I�����ɒ�����<�ށ�U��I��ε���0Rή�tͥ�X�29�j����E���+������s重A'XCGK:$2$�����k�p��Um��������`D�s����ũN�vv@�b8Ǿ�CT��̠�4'���,�ɉ�Z����#����d�}^��E�N��T���먅�~3E!�Q�t� �nH�R�*1�~�R�>��1�$(�p��f̬�*ݤ3�����R�
!����\��"��'_H�WE�y�[Nf�����?��_>�2NM�֭t�qzO^�#����&f�dQe��/?�"#�P�Z��c�a����@�PZP��0�2��U�_�TeId=� �ֵ�ٓ	�"� ��5��ʁ�������8f��F�h]��.]�L0#ſ��/��P��Ƥfu�����ϟ�U�����Ce8Ǩ�^p�g�7j�z��˷��7���@�	�A�Z��M������f-7h@��m�oI��\J�e=�`f�X�v��y�p�G/l�l�(��J��S2�z}��g�ޱ���F���!�E��M����܇���������!�R��s-��CR��%앟����ix�rt��(��֍�p�)�߱��5��m��$�9u��8�۳!�)s����1�[#�{��i�]y�u���I	)���m 1�F�Pu��gkU�]�췔e��^�)���'�X�:/U1�(�PK$;`p������^�U<2�"|���er�dz�T��=�	���'x�P���G�}�����`�jD�������OfKz<�l,"�"t��Z2��h
_(���O�)k�W!�_�n��]��a��c@̳*�� �⬙j<O�	��c��ƨaH_L�t �3�-B����\b���#f��XT�9�ƽEϮh照����=��L��X��d�[5��m�St��N��Ʃ����c��Eqf�-y�ԕ@� �]�%�E�\����h�&��]�L���9O�g>
c�E�uMH��Gx����mo-yÕ̍�Rp���32���6m>W��dFݒ&�����$k��k���B�u���Oz��ʆ9�B�p���yZ�uw�O*h��B�u=�����{��rk,
iN��u�Y�P���o�Ye��@�|44Q�vR��8�I�t���/j9�Si�ߍ�Y�ߑz9�C|\�ׯ_$)�m7N�߽>��Y>�W��:���e��dNVBY0�i0�K���J�Qx��H��h�VJ�kٱu�.�0|��gfE�_A�bC�u4��Gz�%��Be9"Ssz�m��)�	~�"
M�qp���k�BX���US���
�l	h{e���i�Ģ�w0^��[�ډf�إ��_S��Zo+��I���fFP�mR�����wL�9�@��&t7هK��л��R6��J���;�>�á
F�e���&#��{��G��6k�-�ĎD��TY��_�*׃�KR�����6NO�G�\2�ץj�
%��p/���U�C,�?0����O��@��T[��kp��5?M�Q�c���d��dڶ�B�M[Q<i��Rj�������Ré��$����Ɠp�{�È���{�\�|��Ѐ���e_�ʣѾp_���aKT��b�Q��X�Ij�.��{Ql��PI�.Z�c/26�s�T��Z{��]t�Naf�1/�%�0'ӱ!�i����z�(x�ŧ��PxCd��� =��J[�o[ŏ�Nso�c4IB<��h��h`���m�n �S��X-)��}v�9����q>�~Jv���f�B��m ��*�}7�-�q-��5�V2�T0I2F�)v��o=Pi6stn0�l��m0O��Du<TpdQ�e1-U���`��:E<���m�����.BWk�)զ��#��f�iS�#:'���ܨ�Nt~Uj�� �ѓ�����ɸ��`��C�2��L<�0KI:`���aSO�7�J����=_:�U�
R��g�?4�>���`�}q΀c���U��&��U�y�Gg�2�����AoFg��j��a�5�p���(+r]X���e2����QzLE�.I����"�Uct��	HlOjܧ����U��h$
N���ő��D�5�A��{�hK���篠 A�D՝@������ڷdSE����8B���<*%�F!W���qEpS4�!���/hOtfu��кB�r����5 �
`<V�T[�i�c]͘�G�%��>|f0z�� 	��)?�f�Kz�R�j�S��r�A~63"��P	0�(˵�t��$�TŐ��)�����Zy=E�Kg�|kt�b��U b�#�G���<t��₯j�oBkB/<�P*�=�I���{r,���;��R�E�*FL [��a�7srD(����x�4�3J`�O&��ywN�q<#�!�ed�������jT���U���.I�޻*��tk�A��R�̺��X*:��}Cٽ��j��q���S����yk�9����e[aj�@y�|@�4}Kf�J�|�m"�#��2�A%Ho��R��;zULP�~���^Y��S��B's�Z<7�GR�Q�X��+����jNx���{+N����~M�e��ɿ5֐7o�M�ʆ�:[$�(3T���wjZz�Y+����g҃ƍ}��`�rX����U*�t�	�ޖ�{3H���ZJ�����>D�k٠�d���P���b<b
���QHjm�5�o^�!�;��ټi �!Q��x�E'Ka��>���(���1q^sӡ�<�x��ڇh���z����zc�1�f���+�3Z�O���OW�Ru�K(nZ��J߫	&����+��&�\��Q�kkߞ��H���7���n�}�lָN����q��s�,�,3�Ÿ\p�߽S�(6�l�)�m���������o��vF�a�z>��Vv״�mz'�7���GO�I�#��������8�[�K�u����\��U���M	��j5Ȟm��Mۙ��#�`�(+X8�4�d��G7mӪ*�<0X���>��@�&n��^����}Υ����*@S`of4�����zS�[5�����G�K�Q]���iꌌ|F�L�=�7�o��Y���U�"�roվ[J��ci�=Ɖ-vrW��D�����"�
b�jݵ��X9ׂ�i=���M�ܢ��`Lp��lO��O�Ol��uc$J�c7R�o���n^���]�������6ڰ��T�t��*Uj��Sz�,�&��B��՘8 �#��y����
�g�X�}�l�LN���yeӦ� �]�[��݌�x��M)�˦z<F�1����
�"~�ԗ��Z���}UHk*��p��vN��Z�H����γ�d)�N��C�����+����:�x���@���*��Fw��pc����\�1��#94�6��Q��D)i3G����P�d�#b��э���D筳sPA��a��,��q�6L�P1�Q=X�e��N���EI̚��^ǌSJ��Xo�L�ζIyBx�-%��5B�،Ψ<�D]���@P����'zyLv�CaHs�?�!�Ù�Wcr�= �3�?G�����j��MW�V�kS<l���U�Ӥ�ެb1_�*��<�IOi'n���b�,���Z��(`��ex���e6��bD��u㝏&�	�
�@S���A��4B�0��SN[b,����	��zF�Y{/1Q��׆�����������<�R�D���K�b�o��}1L��h	@���oE(\�l�Ų5�V�34!b�آdq.O�i��SR�Mw��,x�!�q�s<���ä�NNp�/3�O'>�ҳ��U1�V�EJ)2�e$��j8�r�Ǟ^�@��5�Ѵv1sp�G�׺����}7���ܪ���4�u����	1�>V�4�s��e8��ʹ�!�u*�D�1U��6��6�m|�GHơɎ��G�%aX͍9I�j2�E�w��NQL�, �5��9�l�z���k�@���u=ߗ�^K���2d���ςh�h	92"<�������z�k�y�#�g�Q����)UL���C��UK1|YjH�"m�Ӌ����CI����T��{���l$�JZC�?~��hI�A��68�N�+C�@=|��k�ڊ�7SVk�+vZѺ�`����g�m�`bI����FCB�H�8��	X�4S~zg��RvH/ъ���� q�����${ T'[K���갉��I\��z��RG������>{K��)��frKy�A��{���!�^U�m�Tn4����R��R~h�y.��S�ECv�uæq��d��z�kִ�����0zľ�WJ�;6F���H^N~0�Ţ�&,)�2^Z�eݺ��$�b��1��53��q5��)�^�:�����}W�'��l-�4����Yᔢ��2���T�,�%}����ZUܙ������giqc�5�;U�� Ts[M��(���y��0�%5aH�n��©n�ڣ�@FT��YP�eޤ\��_��币��a��1���ō�K���;,:q��7܄����1� Qɉ����G5��U����1�d\����Vh�x<�0N��4�E�F=W���a�dJ?P���О�B�@gC�������gk�Cs,|Rz����]�Q��~�1���I�1;Ob��Y�sSR®ʄW)��,�?P9���%Ww�F��q���4k�� �l�d�B�o��������Y5͆�m�����&���U̬3�a"���t@���08�c�,�s�u���J���_�K%�-�5�\3F����Z`t]�*�'��V� (.���e�F��>*vX6�9	�+�:e�KY,܈�����p�0kv���h�+�)�=KXԾQ0���f�͜0�M���by�6�li��F�R����sc�/�c��]�$M)��g�&6�͞�FOim�U�r?;���$�<�o<'[��p�XJ�����p1�w�M:�Wt�B������^��R��dH���5������΁R$uC}�>>�h�PJ�������5�.{����8qPUoJ᪇o�cB�
��ɠ6�1�%BzϲZ�!�j������Z�,Īz��E����%�X��%�xX��V�^�U���i�k!Kߣi嬲p$�@�Gj	>�ҪSn��41BaiN�J;����W(J�|��[�R䟹:L��qn��Q��_{����B1|���kr�D���FT&M�U��>���	�J;��������8�Exs/{V�Ұ����~���	�WmϬT̃Q�L�js�����=���%�!��#%ĉ�`��d��Nޏ�)�|a��Uh Ӡ�}�?!]?��s�Y�h:�a��X�á<=<ɀ_��ȶ���b1��4Ŗ��·��}�<>8A����=���§��
�b����2�'��g��w&��*��s�@��.�Ҵ�8���P��Q~oSVo=�ߞL��h�� 	a����$+����e_@Z.���*�#�}fM^��m��r�+Ġ�f�0���,M���`:��W�C{ETe������!?<j�$8�����j�R-m�jg�T��Rs���C��9��[1��X]#i�:�����ۊqF3������mD���״��z�x���ׂ��,a���d-�g��j"@����"齚T䐔�6��|h�Q��FO/Č��R��y)��l��҃9͠��4�#�1`r^o�*���Y��{��.�;�j���j����Щ���L%����jnp	�)�v��1�P�K��y�.ë�]M�C��$��Ӥ᥮��Y>Q��ܖ7_���7)
������(k{�+B�0���I�����f:Z�#'"��M����9�(�i���n� B���J�ߍ���Z�o���M�6dP^���GA�a�h�c�q2E(-��bSa^��yz,�s��x�C�FO�ه��*T{T1�&ɯ�GzWKNmV�µ}P��є�1�l�9O�a�ч�M������o�ä���Q%�mhDGr�"\�V�G�z	A��Z>��Q]A9�a�Z$Yv��}5���xTc	[��V��������I�����D�P�1�����dSxV�zc|���Qc���ۚ{F`�5i�2���m4^H��w��C�l�����,��`���SU�c�tX��L����K��-�3a�j�+ 5�#�MOĐZ)�"�����hkEZ�X?��4�H�2J>��jҪ� ��d�*= ���^n�|�4�E����
8`�וЊ�g��o���E��U
y�pް���������óR�o�9�ժ������	����X�m�^eFu"�3\�+�MQ���`�T�f��q�t��G+�<״�)���3d�L$�ʖ+��So��nH�=/�Q~�Y~f�T:7�«�Q]̨�PĦ*>j�Լ���{� �Z�G���!-~�����(�s�� ��J�I�ʤ���]';(����� 	.SWp��Swj��ah��}���˾��^Η�x<h��~ߨbD}JB��E��Z���
������,�s��I��}\�l��/�'�zY����B��*Ǉ�X��-75.bH�>��4"wJ%~m扎fL�P?�Ʈ�;�T�]�O��@��
I��6nY�\��.1�ܓ���N���X��Z������õ�߬�vh��Z��71��eσ���p��D����R����[x,I�M�OK�!i���rLi�����F��MǶ��!�1Yl]g�(�K�]���]QL��4�i�=��v���ֵ���8J:��`9֨x��Zh ��W���n���C��}�њ���E�2ȑ����B��5��m럛{��mt� .�qp�V�\�EJ�0�1��8P��0Ŕ2�hb�x=��*�Do�*��#��ʦ�.��Dn�8�j*A�탏��`*G�&z�.��ƞ0��x��S�q�k6������z����_z��'�Nţ?$�g�eMH}1Ly2>�������Y��R3@jd��sk��P���`)���H)� �E��^K2�&�i��a���-�\�	����W-�[�ӝGZj2zz}���A�j����!<Yō)��u���[�7Z�lpΫ�d	�#�!�Ca�������xh�M��h[���*�`��,�m+��T�Jb�����W+J�Aov5Lu��|Uᝫ�d�;�Fd�8��E��{�G`�U��mm�a��hQ,0�0M��U��]J��ɭ>��	5���դ_D���ZG�A#����m�A�|˝�Vh��
i�bP�(�.������$;�^j��5B����l�X��3�#�ƖR_��/PQZ��{�fq_�|��RE�'7.��5���ڎ`QS!�:��eČ�J�M�vM�g�y"�����Ed��d�U�M�]` K�Hk�1zM��CL`��G�A$��P�V%Q��?�� F3{W�����C�������og(��@=�����o�trB6(Kt.ʰ���q���Fq�Az�|�I%�����A	�7+d�X==�׵�Kf]��V;�j4��ã��o)aFn&�T-B3z~��)�����L�D�7�B��uH������e�Y�f�S�Ha��ǋ;��`���t(�"�e�aX�{��.�O�˥W�N�$�NQ@T����'S�>����ċ�n��k1Q1�=��^��˫�$�{,��aAHE��M=�q0�~�8UNL�@@B�KD�U�j5Hn�+Z��|�Y�i`��)lm�Z��76���k�/�I�릘���-�,	����]�{�P��Q;#��Ⱦ�;��}D�uxrb-3̓QI�u�
�n��/���m�����U+	����-�C�r�ʪ�8w$��ʖ��CͶB��֛~�̙/��˙�ua�U,M6��!���=N֔��������E*�{(���j:�x=���C�`6�&X��}��Cpk���4,������2�̧����d�Z��j���>;�F<�z��:��3NcC��� c�1��n9�Re��-B5&oj���W�!��٫*��Y����rP�������(J�/��^���T�Ζ.l��UPG	�WH�]�`�P
�kMX���W�����A��i�dh$ýG;FT�Pr���_e�һw�c̱���J�,5��d5 ��)�m	5�/��f����d�1y�7i��R�}��t��<jK�:���v�＠����������g��Hݰ�P��m��#UO�RO��(��_~�E�`I&x;#3���>X��b��7��~E�#��iXoj�2�~BC�D�"N)���EPG3.'+1���ż@�_�񽸆��U�J=�f˛�r�?|�(τ����G��â��F%U�e,\z�� 5f��v�4�1�%���jI#�P�s.B�P|J,zR��p3"��j
��O�<u�7O���xh[�t1�l�j"Em���W珸�����(p(it�W��K��+ŏ� 7m�
����%ONf�5�5���Ƃ�Z��ؼ����*�h��֎E�W�O�1�5���˯��"����� ��Jj�B�N�n@3k�g[�ë4b�H�C�j��r�����T�lT��\j�KP�&0q��_u�Ϯ���.�M��_�����עB�B=]�CU���l-�ci��I�����PoC��x"�z�5��T�Z�i�C�{n&�A�<"n�5�xH}��4���e7��e��zz��C�a�ELFq����uY�ۉ�Y�?�	�	]Mv��b'�Bƙ�Mj�4�;����?���m�n7��A�1�⡱�k����?2.q���zޫ�?��5)b�����s�O��ū����k�4�j�DO�h;�� �m&j7o⼱�p(ݸ`��b�-��H�YKo@���iZgH���U֣����e�L���-�m�V���K�1�w�v�41��ű#�a��o��!�s�9R�X���⼳��f�<3�Rμ�����u+���b�u_Gg��wV��yI�+`���u-֮=x�wb$��A�ĳ��f����
[�H�Dg�lڪ��՝�:0N��+X�P/&Ծ���uއ�!��������=�k�	S��|b��H�d���F�� m5�|Q��t�MC�,��T��������y����PA��B��׉�'ʖ���$$&��K5�JR~!ћgT�঺k:(�P�U��kׯ���1�*��qCZԸ�l�{�ꘁ�ߛ�����i�	���`\ԓi�Z�DTJQ�9���we�ٰ9��XIi�n�������7&�b�x�n�量Wċ�%RZJ�ϞT�O6#<�!U�S��5Jq�]^�6N��Q7T��<5����H�\I_,>i�P�.��R�R�V�xEZz
���v��X��?X��� b]<r`8�D��U�RA�u&�R�H��4�����״�i��'x�b��rh��]�z���7�a�w�\2�t"�fr���ږ��"y���Q;[9�t�R���'0TD|��x��t;S��l�0Po�@��Kf�pR�����W۲]NY5��A}��@l�^m)�J�X�]�n1C����v�Ӗ�I"^�J�Z��0��:)ߛi6%�qd#��y�P��\�0�8�U3�����س��0/�ْ�S�Q�FLi�Zc�v����W�4N��'�Ji�UZX_�5hYQ�0l�r��R�B�h�Ӕǹ!�Ny��oL��+�(��<!7�C��/�	G(����o�T/��3
�k�j�f���ސQ����3���?����sd�D2*�Rt"Z����`P�.�E(b5a����.�DSA:ʾ:kc+]m߽+�?|c*F�4m�>�N3�L:�fHI园clW���Vg�LIht*L�߫���sZ�]w��BJy ��'�f=�7<H��3Ƶ4pQ��`�T�����Ū��!0W���ئJRl�����já�!�����K��6�w��/m�͋��m�L��n��J�� @TJ��Ҷi���e4�W��*@�,x�Ha&W�Υ{��u���;h5�%N�24�B������OdD=2���������V�x6Q��Neo�l'�����0����4�[(��,F�!��;	�᭛�|v/O0Kc#CI����Ѩe܌ղ��������Ca�h3e��24VS��N�[�U�a�����?Z��}���˦-���=�9�z�Q:�����
[鑆!%��@#��)���L�ө�H=�X7,�Dx���b�n��+�e��~�_5�%dt� �=��ì0�(�'�w��"iz��\�b��y����=ca:E��p(��I����Q����}��_���?�mn�G�lи���Y1y�H3˅�3�o=R�rwƱ�Y̷���j��[k�j�M�(~8h;_����)Q�n��ꕃ��.����7��oK��q�i+Qן'�Plc�h+GA�U+C�ڿ�^LjP?�O�]�ͫPzEm5`��.�$���/]�2���Φ)<ق͘��1��H\X`L'�c=��3�C�zrK;t�B{b6=Ofz��C��%K�p3p�`A������emH)�C�D�( 	�����"�y�����I��[iu2�;�E��|Eb4�u�M?fZ�H)I^���wQ?���F�;1��2��<T�d���G�`&������*�r�ar*��������L�_=�4���KU2W��H��Ƃ�K�c3,Q�$0��Z�%��Y�)H<Ѧ�.��j1E�ϫy�����Y���.�'�۪� D��S*�j�'�H�`�OD �:\7�)�(2�W%��-�a�o��S���;g2M�{����eN����!�P�H�D=��GԳ�V�0���4�70�U���`#~�Ŭ���48n��w�%�&�&�$f����j��l��Q3�}%�bGʨnbop�DK�p��A	���;����xM4��|�����J�]ʇ��G�Y� �01�5�[�ɐ�xR��h:�u��X�K:8R�,�/[5����g���]��������F�����z|\����C��b�q�RHzу�����d�Ӑ���d�zJ�U�����|0��M6���-���MQ*�V����ĈN���j��Ѝ��HkQQ�}�q<���10w�/���S"|n% ��j�u��� T��O9 *��͕�T�I��(�Ŋ ���G7XjH�I��X6܊
aa��!�3K�^(��^��XiL��i��>���ʵ0L�t��w�T�a�R���	�h���n";)�^�{TS7�m�ʹ��,e��O���mi��Z#�����aU�~����b�OM��O�{5&z����1LL����LQ^y��T=H�����H�4f[����%��f �Ι7���\B�S,����hl�SP���q�Έ�� ��Ma��=�Ź��?�&[l00X�~�c!�Em1�+X��'o%p�U��-VP0����9��@D��R�o�-]�ܯ�������Ÿx���o_=���+�$�k�*,��ãy��x�b�Ce(c]/��+B��M�J����J�l���:�)ITU��b��d���YՐ���y�h�E����8m"ƣ�CE���u]��8���K��[g�L֌�&\�I#��j�1~�6��t'��m�a��p>ԛ=�sT���#\�x�r�*��������ٰh=��/_�����"M��B6�ꑑBOG�WXV�]�u�|U1��A�(�u�
��z�/4q�}<���*3�GG�|K)�B��Z;�V3�az���dh�mf�2�?0���#�i���@�i�Z�&�Cy��zɖy���^�����#I�"r8J����c�Ci :q���Mc2��������n`��eRY��}�e;&zT��-����v���o틭�e�a˂ـk�w6I/��W�u�QO�p������ӏ��p_�[K/W�̮W�~�=�x���E��I����B�&b��X���J�sex�fՏ�b���D�';�4��}8����`�~�7�Ҁ4٢��,�2�JTiZ>���P1T)�02t�p�e5��(��K�Ř7fH�}Q#�r[4s�6�øfN�qk\��b��XPN��tVo����سH��B1�! �|,�ǫ�#��������gŅ:	�U�'�����������>ȸ����A�k�b�X/�~����͏z��umy-���݌V�㠐���Z�o�*N���x�}�o�Zܠ�/��"�-S��%�w��V��Lո�z��(40M�$�`��;~z)o�����gZx�t���ܪ�ʗf��U�4L���
3>h#|���5�nlc�D���XX���'��|2��<����#�I��<3����JC��yf�6%�ofH��z�cKb����p��h54$�y�sY�[�k�n�6�c��4�t�����?��O���?H�
�X	����U��?��,�=_J��84��9�)��'ث�tٍ�Y�M�Z=�H�RjFxoH�_��ؐ�o�-��e�s����$R��7�W��Z�x����Д|�&Ja��xJ��Q<m�B��M���#0��M���i��W�*FN�4�Uc:�uVN/Hv�i��s$)�������ہ�CL��,�"��jQ���{�����}D)H��*��?�]��~�8��Y�&M����&~Fet|ch���{ߑ3��������vs�OKy?��;��]8�6Z�7���"QC�kReP�D,�&2��"��][Z����3��]oC{���u`H���~�v�{0�՟�_��7������K)ZY�u7��O�5��;��<5,B�r���<˖ԙj5ڍ�
�4Ƥz8~��l�z��ܚ��J,Qf�Đf�up��w��LcK�F�������:3_����M��\��c,���ϖ�G�$�&i!�A ��x�e�="�<T��E�����CT���ry8���I�v4���ߜW�Yr�LpW�U��U*����YaƚvQBGc�����-�I{����.�G�жf	Γxc,)h�X�J�MM�Rr���I˜��L��b�Đ��ek�\��a؂{ �����'�#��
��g���}(�?~�q���_d��o׫g�5IP�NF�:C�[��v�Ƅvb��~�U�ᒯ">����|�$��YD�:����s"X�Z���Š �a�4�?)T3֭��!hs�=����h]"z��zt��Y&�%2�3Yk�at[�����m��LhoL;�Z��l�w����xs;�>v�ZW	�섣�Q�H؈0E�
�bj��&�x2	ɸ�Vb�^��S�!��ʷ����+�$r?�S/A[n��b�A��&
{P�$�b�� ����7��8��"!��@<Si����x�2�3H+6�EJ7a@�U9Fwt���vՒz�=��'��J1%���k�<�CK<�jٿK*�d�J2�碛�4�&�{tC��0uS2�0^��h"CiH*\qxÀ	���)�r�5L=̲xf^�2�|Ґ�#n�#�<�e,�a�<cO*Y���ma.�J<�B���)�g�PH(��tM�K��֦��"\&�ޤ'&a�C�����Yg�~�۹��aӹ&^�u�L�T=lD{�)��(颂4샦̍�Seu��}?P�
�1}=�,{o�e��9'ՄEߤH�Jc����8�8�Eh��}��ù	�h�j�7�	'��7�����"�B5 ߪ��h����EB�}�D1�d.WK<�K��{V���s�v���h�<��"d��� n�V�(�I�ϥ���3�LR3jƕޝ'�������]~Ag;e�Ԓʁ�贿~��_m1|o������B5��}�o<G�X���UU�����_��p�G�Q��τR��x��|�w�r�'{O�<�(�T�d���_��Z�IgR#r�y�&-�� ���u�M���0H��oQ��D;������8,R|s
�N���Ԡ�
�����FՋ:���M ��a��Ć���K!�f^���Y�2��Y��t�b�`l�����b����R��ݑ$G��� 򪬃����?0�����/;�&����k]TD�<2��o�De&��������;R�.d�\����z��������])�'��E���k�]{I��[Ș�=A���a��o��lr�ܔ��J#f�U���9\�����h~}�O����.#��J���W��
��aѮ��^����
�.�އ�����Yi�S�yJ�H�D�5;�3��	����v*�fbs���,=�FY�����h`Y�'�L �v���X�I�R ���43��*���^f�K�5���SF�4י8{w ���l~����vL��
��k�h	��c5��rMR�Zn���7�9��pL_TfK٭���Р�����n�Ĳ����n]*],�0dI�ȼj#������Z����-�����	+��--�K��4�\|�i`�i O[������eC�h�A�Cp�9�e��@ry�i.WΤ_,��'�&#�I�Jgr��Yκ�C4*�-�\|#�ȝ�O��l-?W�{�B����?X-=F�2ܕ�C�� ��?��z�ʻw?m�����)���0�!�̃�"�<���<�pZ'�h��^�����k����z �@?����a��t�Wдޣ� )�m�CLzx�����v�����N��ѵ���+~�C��u�@Js�SIO�E��0���C���L�ӯՇ�>����?�H3#m��A���lf���	D�y��A7�,�N�;3��%L�޹؛�a7�F��Q�,��i��l����=6�4��t�w8���nU�����֯��
�7�*��-1�h�!�Z�]D�vF���=���c�Oκ.wV_�����s>�'u/������eGsjd7�D?}�F �G)�}_�e����<���}aw����o�����?�}���mz����t*�MU1�>�枲Y���7o#@������Fm(Ϩ:��1}�z��t&�r��N:7S��v�4�p��L���sr�un�X��NP۟�p}�_ca���D���s� �O尖��c̓#�����$��X��9<���u�-�"0`M�_.�_���;��H##�5��A�zӴܿ���df����wp��kՐH'�Ӽ��t���8^sO��nt8�eL��͛&p��9�6����0��R���%��VQ��,ý�X�V_`����Á�o��a��w�޸�6�}���?����wi�.#�۱4�T���:pߒrR���.$~�©��¼�;Gj��1����8�MK.����ƦkY��+K�l�i�%��Ve�f<���BXJ�_�,q�M$�mf����}�O�-�z�X�\�b�h�,`?.�nĢ�먛]�oA�������7e��tX��zՄ��|����LK�7�&�߂h��Mf����;�zh�=�Ad���
%J�q�>�fR�M�ދ�1694�:]����+��'�Ӑ9T
{+�,7����Q� v�k�de���=-^/���.��jRIOn{;>�"|�/����ً?|�#�,+$�+Ma�KT�� ������#X���m�`x�Df%.݊U�����1ف�.���6�������6�ɱ�8h�����3����J��=.��Yi91���\�l��������k��c9��^�D��+�c4���B'��=�q�+[��͝��?�;�ӟ���3R;t��������S��D���yU�t��+���O��JA��6T��vA/8�ۦ�ʌ �bEAT��H3gP��v'��\ѣ$��kn|�NK��5�M
J�-H�l,*e��UW�a'6؎C�l�n���Ȱ��	(I��U3�([��	���>��p��G�1ɑ��8��X�bbD�m˦�o����ّ�|�t�������*�l����?�/;�J#��GI�	J�#�\�;�J�^<l� 69����n�#�0�M+��j._.��l0J�LmY��^�J����<�A���4Z5��8֣6 �^���qb��~�\gsE�t�7�@H���Η��(q����|\�qbEC(��c*�A�����{��U���>'�b�9�ơ�uM��xj�uXĢ����π��
 �A�O�[X�ကi�~/88��2�n��7ǉQ�4�G�(��y0T���.����R%��,R��K���g���?X;��]+���s��av�d�yR������e?/����Ha�$�@�׃P?�ܛ�N�Y�c
"6�r����<yl?p�_tۍ�@�-X|:�l��D�ؘv,^!��m4��x"�)26֘;ŵ�yD��4�fQxfe��&�n{G2o��F!���ow���$<��&1.����R�[���K��_�'V�Y�5��^
��,�b̌L���V���A_g��2��H��ImsR�=8�:��q![���-�?C�S�ݭ�]F���|?��dmv�ﷆG�,�\8J�AZ� �Z�E�Lo,B-�1�����Q�2k�8��cs˻��E���������+�O����e��P�������W��O�JR���ӻ�}�>��c�S;׼��Xm��ٳK��W�伕~�n��5̮���H��-�`^2��p�[�g�a�'��i 3��8�\v2W�~��Hϲ�:��$�����o����˟�L�'����x��yIB0i?%O�t\)%���p�����Yj�H��wYe�u�Ԯ.�>S��ߟN�]�Aw]Z���ԍ�&�*45�֤}�>Q�e�b���
S�j-���^�vS�(/ڌSIHV�;���V�J50nM<��Ԁ���)~�Y�����b���"�y���M�=
�)��CF^%,�ospa��P���YY�,��9��u�Ԭ9<�4NP=)�CH���dH��5��cA�8�������B���ɓ���u�>h��咢�s(��p̂����Q�����C��dh4O;6��QϮ$lJ>�d_�9�W���m�a��O�,�Q/��,���C�����؅*� �榉�ƗKޗ�	��Xc|����ᢱ������|�K�x'�1l�y��I-�c�Y�D���v���M�GZg���X򍱑��TF�VJ���1�fV�,+1�og���y�9h�NT~4���F]���öR^��|9{��I�l�La��ŀ����`��Qj@M�ۀMs���gd�m�צ7��^��- 6t�����.��1tWr(��ţS�,tQIn�4�mи���eyǒ,�FY�R�*�g�rO�nHq����4�<����C��Y�E��%�� ӣ��jd��o�d��H������vc��и�s�!x�7���3a3>|�(K,�ƵZ�DUrf��������qH��Y�ڨ`��5� ��a���� �@����UT����ǿ#8˶	22�:�H�r����BM��l�с�\3���h�g�#`����Vt�����&n�-	�f��S��-3]E"^`}�����������P<1��i�
jU�Ċ�]j3�<v'lv���z����V��w�w�����X���B'I�;���Mf$��, ����XG����{7$F�b�@� �v
����yz.;m��lLU_�!7��>h���[k���K��O\8�C%us~�U�/;����!��42�X`[G�[��\� ���ʚ� �va&����uޑ���#�h�n_��h�d���]9��j�9�e�8�l���A����z���y��3�M�O!�|H:�ihd����an�x���
�\CS�d�J#���Aԥ�Bgs Tm�z�wwz�]�_�𻠰_g�T�/�w��Z}�wQN_4;���p5�����\gɡ9yt��#<:��$�t`�[�̾D�������T�3��볭�����S"��zX\7�/#q}�n���xnc��G�]9ዯ1GfJB`���%u|�~�=a�j��{�VS�:�{�ZhZQ�����y����z��޿���WC�T�v�o?������Q ���Q��ZjF�uҡ�F�7eC���n<�/z���u���/�9�O9�{�E� ��<NQ����1$������q�7/��Qb�ӑ�� ��^�͓�Hrwu(^ˋ������Y� x���:��w4�62��p�&]7n�k�� <:�u*��v��L��|?��W)T2#�f�vE��B,�����H�������sl|�ldg
R��H��E��$v&��u��wx#}-[56� �;�����Q�4�84��
)9�����޲[Cn�N�\�'�JX��&�����c�u�.)V�!PVeշĽ�!�D�%��������Z�#X`�Ә��j��ُ�Hec9/��3#�5]�����=����q�W�mG-��:�z��f<�Y��O��h�:�T�]D	����`\������s|H�kf�*���iS���Ã�b���\�� G���k�k���'���v��q Uv��
�u�m���p��id������X4��$��bI��dwo�^��}Hn`(l4v���э�m^�x���4^��F)z�k��O�c �'��~��X)��<w���1��[I�4�g��MPe���*\�D`�F���ޤv�7}�mY�+�%s���s9Ks	퉤��ՙ�7d/UZN���ɴ���.���~��.�Yu��,g+��-c�������(��|怽��{�6I�x��'K	{Y�͑��w��$�x�&qI�Dru�sҽGA����Q^O4|�qͣ>��y�f#k80c��A�ް�����;MX�HW�A	��{��	��ʽ8*K�fƃ�2p]p���ߓpC|Y��C� ��~�ܿ!)O�dB��i���۽��1ꮦ�l5ǸՁ�k^�8�����u�
n�`�c~:9K#h����>�
x(���$�����ת���71]�뗌�8���Ĭj����:Q[�j�Դ�1*}�{qu -��]֠/Y��r�((ݢ;�r��mGpR���ݛN���7^�Y�O��Ҭ�xΓU
���M��d��1��:�榅fy�W�F����!0yJ�
�i\����3�ΜG�=ǴeL̘�#}�ad)s6\<���G��+�d3��%�����A�����qy�@jQ#�s���\��Ȅ���QM\c]<k*& 
�ă����c�k��&e�*�W�L��u>�����q��t�%6e`��F��.=����)�!y��)�2P���+�4Kus=K���� y�e�r~i�P�y�C޶�_댡^J��� ��-Mmnb#�p��8�!��Z���쮲hFׁ���� �G�H;~��Ǹ'��8�6��yu4��Q~�����"]�b�V��dU����r��@��^n"�Gm[�@���������o�jV�D{��]eJ�[�1�{h$c��c�K��ݹu]����������=�X�-5�\jc��GQ��%qFf���]��s�Pο�J���Mcr���V���	*�,2�ZC%# �T[�9�9Q*� �?D�B���扇��;�&@Ykd���X�5p]�M�1D�جS�[�`��(�,\f�Ɨ�|?��H*-�bT����%1���K����|��5ARp�y7�r��A����<i���d�uh�����w-ŗ���(�i˵���p�e>#� M��>[QW�����y{<�(a,k��>|L���� ��-�!�%�c�8z��7ԦE���}Yc�ꑎB�R�%r���x�j�Yc{Q���T���Y�-�Ӝ)��,��p���@�*�Q޵�=6Ia�R����D
����Ʉ2ҁv�P�q]�L(ͣ�)$��k�6ÿ��k���(���}	ap�ĵ�z�Z���)��4ơZ��g��,�V<.<���1+��g�"�-�Yֵ22<���.d'���zt6���7%�:'����c�u�mv�9��F��)^��2k^��k�"�]��U�]I�~��4�rJ/�DZ�&�~¼��N0э(T���w�(_\�A�����CH`j��p�k�3G�?�s\Lb�7=��8�pL�����]�yɃ���r�:�����:y�qZf�z�ӴW�!�Z:����ǇtU��ꖙ��������������+�<�Y�����^)s<���gP1e����Sor������j�Y���þ�yc��M�B4H��%̢����17cwf��Fs�V�2�;e8��"�r
B�|
�%+��X� �iv������XP���APP�9"�{��^���$fI\5���T9�p������^��%��pf�x��UR��$�׫�7�2QȊ��N�dӯ*�*˦b�����jg��A>����Ϊ����1H�SA�\{C�?>�c�^�o�A{7���l���x��q�@��ْ.���JS�7d����J��1���]&4u���,��C<?�҉�y�"=+����Ę斲KI����FW�������Vje���7;��2��i��Il*qH�-ʱ$��s�-5_�躯��/nN|�^ԧl����L�z��?�9Wd c�f.�����m�r775�Z���4p�[�Q~]���Q2���
,�&ۦ�LR�0�&Ӄ�8lط���� ���,�v�����A��K���Y�ڵ�����Y��J���Nv}f��J�x�~/���U�����f�w H�h��oqRO��Sr��v�^�8�j��s '�@�5I;{|�/0X x��m)Rh�!�o���V��p�5]��ƹ9�HǒJY\>>(����@��b���g����X�]�N�'����zph�XGa���9��Z	��G���)iejܪ�h���q<�lyX<�r��ˎ�w�������vXկ�:afw�R �}�F��ZLJl�?f����)��~z�����Ac��+��1
l�[/�-�:��ܲd�S_���_��C���MY/&CV��<e�!i��F�M�^v{K�9lřV�&�@Ja!ꡇ��䑣��?����0��6�G��-;��{���A�� �%]�{���Y�kLIy��WƟ�	��9X�=�ˬn9�Y��ṏ��p�!�Ixnϝ�@��S����T�gC#ș�(�Y�~u}�QJ�Gl��e���ln���I���q�`�\�cN4��P��U����`��ZCe�k2M�]�G�>i�|h��i����T�Y�3��ʸ!	��YG X�D��,Wj&@�����3#�
�b@rcmNH(�z��0R��N�jVM�6U�G/E|�|�x���J���1�ov���i�v0#�kNӍމ�~`�����=F ���訆r��}�Tj�>#���CǾ�~ٽN��Q�]F��?�\�e $w]���d�D[v��{��T,֯_w�As��	[���{:�Ed{>`1�zy�llf�m��ʛ�JZ�J����M �N��:fyu��Bg��7�Z഻S��#�H�Df���c���3��c�}
΢�q>���':��S�Q�����ѣ�C�;�R{�F#`���j�q�Aσ	�y��`��.+�����<�8����<=>3�GС�7X8F~f3�f�3����Aoc�<;�Z��Y��W��#g~������?�5W���r�pů߾8��#a <�_�(	h��H�JS+�fY>�=u���'����8̿�:�7A��,�B�ǫ�I����UFQNc2���]���7�F�dҎH?��ⲗ����{�����0�%���	� 6J��Uc�����V[��x�rI�i�|��ȭ�S�f���FV�j�c�z�\�����i2�'КA�.�5�tjxC��_�%~
5��=!�Aՙot&������t��7c�y�{yΎ/�`V֓��GNK�Ů��-G�4��0nX]���Ħ�x=��O�IKd���{�y��UT�)L�nA9�f��J���%ɸ��qV⛙�,��.5E�|�1��.60K�.�X���s����-��j�9��dHe�dv�tO,M��	��D�������%���������uh�{P�����G�w̆�x���\�K�ן����w�ބ֚�60�`�(�Aխt��k��W��=�3��$��i�՟�����,k0�I�V�͝̊�X�}�2�Q,�UA����\�Fj>����k�� >��7�b��I�Y[��4��׊��}<D��T�%� �pu���D?�T>}�\>~�P�����?��X�v��g0M�Ti�Q����;��׈A��Y����Ȳ�,�ԞʾZ��F���ɘv�i3��lD����0�f��4&JϏK\˻8�����R6^�dk���qk_'�yh�!��B)�w�����O����1p�HEc|Ee��D���y�ωmƂ$
R�� 8��.���l��[T�$-�����o�\Č�:`�XT�.nGy�[�zJ���۫r#��2X��ܟ_U1c�31z��ˎ������]�&�zDݰ��b�m�O.M�Fa��"����i��J�O�4<��rh"�"�	��0�wJ�y��|��	'||a�e�e�_1����{�d�>5t�z~�[\���XcM�����ndi�Pw�fh�M��v���F6� �%��׉�Q��A�C(C1�V_m��qp��p��,A-6��]����cTfݧF��5�i��K�=_>2D���'����UڧO�@�Gdc�w/5��a@�o�0=��R�����f�>8����k��0��ب���Rn,%�l�����{	�Z;�h�]ǔuM�J���>=@��Z��UJ�U���%Fp+G�7�$���!�Sgb9����f��;V��yޫMW�R:��(p2�LM)bXq��;zؐ1�B�9:�=UR���@zJ�!,����sy��t�Cc	�F�Jn���#�/���u��D�_s]Mբ��H������s��n����. ���H����e�^����Zɡ���*�u�!q�i��aᆘ;��޿��"V�x}�៴8����p��)��á}�h���eӇ�tz�~�`{���nZ8�pꃃ9/c�?��m��3\k����y������V��"o��Y���FUQ7>ab�S��glp7����d��)=]�56�i
Co߆%2��j�2�~� �g1E3h�w����LJ���*�0ǭrz>n��`�%����7���O�j�rKp��!��H��x��g�F�(X$E�c5o��r�d ��4��lٴ4n{���dbs<m�|U�=X����#4�)��c͡j�>���=4�z%ؿ�*G�R��������UD�/5(�%?��*�^��N�}cc���R�x��徴�t�k��l=�D�F%َ�'���A�}�.�U�N��bn����X�A]�{ʂ3ep`�� �͚x��?���n���Wh���3�q���T�~�ٻC�窇�zCX-|���pTUM��g]��d㭨�1W��p�i4W��t�7���<6����X���F��.dĞe�q��Y6A�QY4��(�X��ۉ���by�e�kC붧 q�Y~�H��u�vҦõ#�J�/M��q�)%���Ą:˫vVݴ�v�Zl��墮}��1q�h����$�uR�R��%��9�<��ڊ���E&}b�4E��2�V�:����d���0#��p�Feૂe����������ݞ�k�ɺY#��y:����$�F�U�?�ت
ɒ�=_v�>��q�(�� J��1Fk)���y3g��>��O��e�{��_x���^~?DА�3��k�A�(zI ,!�F���7�K|ă���m��L�3m��-��`�����g���dԙ�l��/�%p뚳|*�O�]f�IL;7y���&�鐴`U�`0�Ùl���������oV .:X�fǛ:��ۢ��F���,��B�����T��#� jH�.��$��ق`�h��)k�͜�F֪U>���$�ɦ����+ ����Ui�&��Ȧ�ϊ��Ƴ����[�w��s���ɲ�J��8��fɎSl�mVQ���&�ϴH�"�ŝ`_3g�{j�K���gЙ�0�s�S���R� G�nޕ�%�t��{��0G0zt)�7w�|�hg!FYt��Ӭ�LL�m�5kfY��L�s�>��[���(���R�3H�g�E�D��F�P��ɭ%�,�'1��s�J��w�
���O�YS����ÕRiJV�Mf-E��%���1��pp��������q��ܬ�~��dN�?v�@�Ct���������Z�\�}��((�2�ը�I��H�l|�b�j������Q�k���_S��� 1���׳�cW+�m;�b���aǪKm6��U7p��0iS}� 5�,׻&�u��74X����bS�f��M�(o�0��t�I���â�:�$��,�+o��_�ZL"\OAs��l�a�������Hc�ȅkML+LׇX�+������8�<�uQ���Q�"������֕���#�͐r
C��'�}��a�s�O)�>��D�A�Z4&��q9ˏb�LX��w��Y��C2|o𜸖��q��#;�,\ʽ�T�^�^�% 8���m<yj�>�s³����ޡ���.��[՘�Ds�r\���,7(ӡZZ-Fi/��.�&����y9�fW��hA����ʺm�<��~�Nw�P�����լF�4Y�����:[�1�`�Yo��P�H�s�F#h�Oi���R�{Q�����y��@�
�V*�3diW?�
q���r��*��_�,�ۿ~�Nj4MJ��d_!�e��#�(:��T;�Z�s�f�LwR�m3`_�(��u`�p���m�`���%������G�Ny,owYW_�k%�CV�I����)G"�ɰѸ]�#�BN��^Cj� ߁g��xe�M�Wt��e�'>�\�jFd�M͚��Kl~�=<A��1��M
�~#^.��[Wy�e�s�Yo���U�m4��u�5�E<��CT/�	lbb�$��K�GŠTF���/�ds��ڗ��"h�a51�$�IB&�=X�zJ��+�A�bjk�%y��N�(Ј�%��?�yS��@��{9_�E��f��q��J��U2U��� ;�A���x0��`�\�X�h�ь�d�Uto'U��]y���k��J����FT-�w���ws����:�S6)�bu��p[��g.r��҂ʅ�@��(<d����ώ]`M͟i�Y9��������t�#��o��d���ɨ��~�n_�h;f�!)4/2�m�6�Ng�@>%��A`�5<o�_�g�7j��y�p���s���F��{�a�b���\��:�p��w�c�{��M�bǼ��/�yIE�4Uyfd �\�U?���i;�*h�Mˣ���)�� ��I*d�8x�q��3������u�D�Xk������-��(:��*	ƀDg4nFEc�\ٺ�9��� F����C?РSm��[��1�-����t�5���3�z�y�p�E�-^�*�/�h�|��'��h8�*�	" y�EKZ*���]E3|S3�"ik�{ �9*>X1�fJ�t��!�1ɕs�fVt=�EŜh+,�&�^b�sd^�b6�SB�{��M��ؗ��HYU�fl�M-���:�C�������F�
��"�� I|Ɔ�B�ldб�1\���1G(���<�R�8��2�F+I����8e#4d}Lb��ٗ�ۗn>UA�Ppq&��%n�u��\́�f�GV,���E5���l�X%�>����(���>df�d�8���T�@��1�s-Vl����:�� �4���ý�%�7q�ѽ�x�(%�����y4��4/"VS�.�s��S|��>�|wX1�cP��}���<�@�~�� 43�ib�:�x/��^ơ";�S���@�d&���j���R�ɠ��	���o�<ש�y_Ƽ\�GY�r����Aّ)��4�qݪ��L�.w��E�:8��{g>D���N�pKH���_dA�y��F��9s
�C�Ǹ���דБ�A�b�tHH���]��3u�����������3��$�6}��;i�PlYgx �/�﵎{i�Ӎ�q� �Rl�G��~(�7�\���؝ɼ��{23W�xZ���r��(�Q���1'uQfp���=�,2��-~7�%|���(��\*�=+>H�
�����&�L�cf��AA����p���nFJt��k�$�f�mݸ���~~��y�n*�a°�g0xE��RM�W��t��&3���ڇG�9�k�����yx����0�7񞱠LcX�xX�ɗt�ٟ���/����m`�q�U���02����m�O[����V���v��b���H' �n6��0Lï�� �᳚^��<�}��(19DNs�p�e*=�v�������i��7ǘ$�.1a�[�k�������f>�}V߅>�J����Z #�w��_ޝS��g&(��"�Z8���<�Hi�Φ��A��`F
!BAt8�$z
3����RLWUZ�6 MY�B��3���]м֥R4;�)�vY10�*��u���*�^Ѥд�l�+�ѻ+���m���y���4��2����iL�K��r���v�i�k�>�)q�n�:�2X8�4.jL��&0W��lASX��?_&0EME��k�v�n4����d/�zeײm�}���{��������I�.��Z�B���֛�"d6VnB��Q\;u��؝��=t�-��쭸w��#�1_v������zTu�yM�Tbd	L"�Y�o�5?�qoc�Ƴ����F&)k!cL�^/�X��zt�y�.�!�Ri͌1�D�?�h�8���;�I�pG��E�{�]O�����F�3_כ��CC���Lp�֚��.)G�l���$�o3����%����	��nG'���3S79$����ł�ϭ �~��cnrf�n�x�D������E�}W���#�t�)�k��"��@Q�lY����>�����,�N����A�Ǭ�Y�Ѱ�!�I�\�7VZW5�Az������ׁ��]U�k\�)xw	g).�F.�|A莋_
�6�J��jR;��t�)wd�u t��*��ܠM|�|_\h�8��R��|j���`v�'�dhJX+=+�!E�z||�)��U��i*�P2O$��ƀ���x�� �ΐ��n���4׸K'f�O�V��NQ< *lpkoq��t"�	]޿����������̸1�����N����e��r���i�5j&޻v6F�^�P���D �R�&*I�[$��h�ވ�I�視<�S��hL����3H�`�t�e����UH�p����ƚ��� ��)�JӾ=((�B��vɹ��|������x�ǫ�����9V��*/f< ���_��c��ڊ�y
��M'�2D4J/W�4jP�o�����ڰIzȊ��*�z�z	�ε�2�Ai�k�!m�A}��Z+�?>�zxH��Y(�k���M�a!b���DdYN�0cf���������PN�k�4VD��yW�e�J�jD����>�V�	��.P������Oq����MA`��=�	�O���]��
��A��aP�V��Yɧ n6��[�$�Ts櫭]�"%}��6�ie��G|*�l*�(!cOG��:�囡[�ch�ե4��$�߼(�g�E,��8W���uG.���O��g6�r�y��v�H����x�a�`�>�z{�+�k��3_2��ŋo+�MA��b9�9���H�;��C���9��^�6�S_gqx{-�%�.����|�M�t�P2��J*����Fv�T���3VT�L���I��T;��iP�>�f��=F�Y~�]�QԤ�x����/��WKYt��mnZnТ�� ��12���%���G�����J)E�Y�x�����Ш�5��՘��x
�=��/�8��|��&�h������kI�B���l��u��Ց�.sML*8;��,�:���w[Ȏe��C���3�!� �pU6���7���m2��e�w�KֻR_��i��I53��ն��8p���<>Q�	�|4`z����^����~���&�.����A������zj�z����	�k�B��<	�<e)�����.*N�V�`�΁x���p��9z��ˆ�o�t
����!2�]��P���4��l��6"��(+G6���:��*�#��6�}w�=j����+8�6��7�N�a�2ԕ,����@=�ڝm�����q\�{=Hco�._�M��U5x���m
�Z��}��_ML�,j��A��0{(��`	ʏèk��Sn"g���pl�%�h 3�^�@U�n�ޣw�ۯ�qݲ���!��z�O�|���O��9���[�JhMz~����N���X�'㐂hĊ#b�P�a�iAc��sJ����XaVٲ;�'(��'�Gqm������W�c�
�<*	�*�4�r-��WT:���[���ل]�7pӵk��:��5Pa�:Wʟo�n�<jCJ���Y��w���jS��'6g8��X��۝ܰY�l&/@�M�j�Դ1 �1N�Ǉ�(+��q��3� 1�����:k�\צ�#��m���iH�b�L.�TiZ�sC�F^�F�RWe(�7u=K6炏��+n���b�r�.�B].sd��c3E��y�}o'p46h�G3kZ�㩜��M�R���h���>(o���#�7�]��]�^���ِ����Z��m}:1[0Ab�����sRrz��[�c�e-���X]Ib~\7��٭��#�l�3��+�L����}�qM�P�7S��l0�PXc�����C�$�c�^F�:���$W3����?�!̔m�KŽ��!,�^��� �O?+㮬�'���T�7�uK�E�Nd�&��F�`��`��������Y&E��a���TK���>�tÎ=�
ٓh�`I�Hǿ���G�X��e�Nj1	L�r�F#b<���YK2a���R�ŗ��j����.ЖRR������s�`J���FI��8���5U@|�*��@z����K�.X���0a>т%:��n���v�SQt��z�)�'��eW'��&��8�@j:�Md��h�7�W�!�D�*&��[�<='A�J"��<)D0�ri����!�LM�?O�f9��ݟV->�"��V p�(l���nРM:�2�8��)�(�#'�E��0�XB�H`JP`�����Ǚ�y;Ȟ���{��4ω㽄�t8h�� �"O~sX]2[�ڭ,���ɍlR<�&�&~�3�Šr�k{&L�C�X��JCR�G��Q�5*�q�g�Y%M���(v�!�"+�5�\.iHeF�Oݴlh��ow�^��v�)�	���(�쪷ʘ�Y��E��y�
a��J��$l�@:�3�Œ�YD+ޘPC�l�y�\��,�ܲ�j����L�*X`����������Q0�5�秤.�`�A8 "ǻ���d��J&�Gsn��'wZ�wu��x4Vſ�D-w�ɫ����X�d��ڡ��?�㓴�_��.8�<Ŵ�z�l�9;���.%|��	�X�p�H��\&�:�g��vx��<Kg�#nd��c30�R�.v�t�L�H�K�R\�1{�F�`������"���0āt�ǒ���{GFa���Ecs?�����N�����n�i�����5�'&�ݏ������5�{䝟�Y����l̊)�d	mL�g�[��}ɮ��I��
	��ri��lks`&�?c�=�������{��"��R��}�#�}��U7�A࢘�9F ���4&����q��Ш�K�FG��$����'�6xmX�Y�`��� \�U��Ɯpg�kH{1� �@O��df���`��.#���G�����l���)�M8�A���A+�)I�D�&nʌ��pcSd��;�1c�
�̷�<�N��U[����g�Y��σ�.���ϻ_�Q#�*F��q�!P�M��n؋���|��-6�iM$y�wY@���r<mswu�ƿ���� ��t:s�rMgz��ѝ{p��Kw� k,�/��]�Ez�o�]�4Xr���
\&W�m�`E��c.��N�qΠ�fU�3�q���4맙�Tq�I&�u1,*���RV��Vxy3�`�rw`�E#s��-�hj��xM%��V> ����O0I�������x-��(2"�3un?������X�bg��Z���ԃ��a��Pח 冉��Z#K�rG6�<ΜS$�Mgw&�����l��!��]�Gݟ��=�j��K�G�/*	���k�}R�l���9+6W����ӻz��O<�0N>����6��)`����Rs��.ON4�/A��ǽF��b�WC�x�N�7a�mc!{VN������Y���.3��&�9�?R-��PV��£���=|�JNZ.jd�X���bsyQc�B�fIf���/6�l��ϳ�xT}�Hޞ�rk�hT�Ø�G�G~���M4�EZ}>N
ڕ�HI%3?l|x$R�9H�[����c��4$�(sNj� +w�6d�P؜B�%����]g��E��KG\��!�3ZK�jQ>�ݭn�^�D���P��@0�"���a�"lS�8� �_oȠ^��ڲ���V����y��FD��p�=�v�0�boD����^NA|����Ƽ^nY����tL���XV=��Mì�vm�x����+�W?\���`V�C�d��;��=�	���)���7z��N��Sz�kr�G�%~����i��m�� �uű?��bd�A�oB��p���0����~vӵNq߾y�U<|�E����+d��'�N�J8Goļz㧆��su��:��/���!�oЂ@���d��L�g0g�{(��] 5���Q윭�x�ϧ�*����`�&�(���$ʒy��@���7�F�|�ǿhG 4���<A�i�Yb�?$�����-2U�S��4:e�?��sy���(�@��ж�,��i�͋H�/�m����Yɷ�R4t����e"�%4�x,��1�r"G+h�Z��.L�#u�d�R.`�<鸵�I��(��<v��Q	�)r4D�k��%Cb���Uv�y��4�~�$	�~�-�K@�ۙ���;����ئ4���-���X��B�(9ֻV/�F�Q���<�#����,��FF���)�&4���l��a���We�U�h������h�$��c��_r�ʲV?Lv�۸�X��#G�	�����RH���Yh쿆��(~+y�X�*�(r,=$HG�S_I�/و:�s(�_��v���(��?�Q�	��7p��F؛����_��_˿������?h:�����.>n��--��3(fpDG^��0(T�A\�l�[';C�YsI)������V��@V��5�Y�_��'�J��d���JT��	*x�#��`��&���������X$�m�L�9�o��]��a��Es�(�tZ��*!���es�m�:�Q��#���@�-N�����K���_4�Q��9��X�ӀL2���׽eh� ��2�Sw���R��wc��\]��+̰9KΘٹi�{1�H��,�Z�	Z�mɥC�z8��.�]hg���AgM��I����r����n���B��A��ٞ(������߷��"��K��[\�V�ʺ�ɩ�jc���p�际�D峖�f 6α�r������)��;���f! �����kq8�?��G)ccb� 95GY��5a����)�:	��s|��Ici.��:_��wJ�q�cP��o8
��e���)�xO�o�����R" 9{w80~2aL$@p���r�"�W� f*���U�l�|��޿]~z��&��@�rp~�NG]6J	�`�c�����������?/�kY���ګWo4��T|���.��{M�u+j��n6]7�R���3%��jU^h�{N�v���n��aSi_;VĳL����#m�����`��O�y��}��I�4�5H[|��MVT򃯆P��'����x#TP�����-(�2r�3g��CEo"t��B�c|úLA�Y�[5�uYY���xy��m��
%��m����|w�/��$���E��:@��b�yv6�MVa��1H�Mǎ�U'~/�+�fj#*���)D���4U�jcc��\
��˷�����@�>�u��7[�1t�ew�#MhH3�V�v]�Z��-8n�[��Z	k�F� �	9c<6�m=����2���Q�}���D'}(W0zz�)2�=�:��w^2X�<�Na�i�����D)���bqo^me���NhԬ]P��D�h��M��XS[5 ���Z�{�j;�ߗ��_c�}�C�����/�}-9�G�<<r�*:�`���F#�����ğ�IPI`�:��{6�^?N$�*:Xa���-�_~�u�}��޽����z`C7�n=F�8�z�}��A�܍ʘ����V��%��X�Ț��o�������3�- C��ʰ����⹖�MǪk���q�����2o��\+ºTity��!?J"�7S��3ZsH��f�X6Z�6L��,[�)���I�����8�K�ɲ�$&1�� 6)�v½�V��ӌ���YoY�z#e��rߝ�yT	�aR��:�í����kt ��m�73���$z>����i+޼~^���	��ϐ<�4K�����Ix �M��|t��0a����S�H1qS�$�E�Q�k�������.n��%����ڂhh�g(���yY�sЀ���}�ҟ��o������m9�K��x>���t���M�n�����)��o�x�~�2���O���K߅FԒ&�x���n�g���)�����i�\q�@���@̏������o5̖1�~����C���6������(����so����*��p7����_~�����+9���h���K�I�Y�?Qm�޻�8Q�SE������� ��K�w7P�u�@z����9/�����K�1�h��@f��*=����䙃#��8
�u0�e���W6��]׮�xݗ�s��^��@�4W@oB.��˷���{�ödVW~f��G
"N��jTA��@:O��s�UI�w����Ϙ�R��E9f5Y���^k�74�na�� ��Q.6M婉�c\o�v 	/�Aq��8#%=�-��W��^c�����[wZ�9�"���'f�[0����%��>��l$d����o�7���?M����@zN*���<�OIu�5<0]4����Ag@-2�-9mAb}�C�95�-k��sl�w�^��#!�V�@��?���!����S�}���Oa�Z�~p3<�>p��],��n�׺vKl��rbd�v(-���K|�N�3����[@yS~���(���z��t���v�##}�@ڔ7���m�����QB����wRf�6�����˿�e��������ӑ�>�sd�ӈ��E����c4N~���@e�n���ˉ͋5�i����ś���U�QU��իf��z�chLt�c+!��脪�
��/�v[�NCT%?m�_������#�iD��X �Ϙ~K_<���m��/��P�{:p���<�Ên3p�E=�C EF�eF�@ʾcW��D`	*�N�6*z~X������V���۶6����a�x� �@JX��?�N&u�Yaܶ����Sf�L`���ç�ш�d�a�:��"��~�i[�2n�����f��k�hI�����fP�����(4S.���/����I��^k￫8,���H۽)'�&J�Kz����
�]��6z�=G����l47&�RvdV�]�.O!)tgm���X��JL��s~y.��~���"�SL_T��w�۫�C.�Z����ھ�7����5�[�C�Agz���|�z�r3H����Q<�,ż�F�&�O��!�y�1�<ؤ����Jk���<�S"��̠���m�j�U�bNz-�Zl�]iM.,��wB�8d�(	�>����o�y�=�c�������i�D0LQ�c����:^�����m��0m��8K� Z͛�~��9>½X�IЉ�z�d��a�ulb��N�3�)�	^W:i������W)�N����iZ��֑+��\hd���(�(F�fqǊ5�?gf��γ�IC��NF�0C����X1-���|�"8d?$�=�������}`c�Kiuhp�1f�0{;�NW����=.j�R�.]�Ĉ���&����k�t�5��K�+E��h���N,��Mpu⋳���a���6��?呺�'��h��߲��aG����N��ݰS���Y�96�^�VG|H=U��W	gopT�3�\�J'����*Wp]��,M��Ը�3��3���Wuc	|��9�	W����󘔞1�5��A��g�������`?��l�R�j���k�ej՗գF�� �f��[w����݃�$��P����2g�u����ܵ�)�}ג��nWg5M��Ϡ�l�����B�`�ؤ�)U��f��LFDP\N�����p�o5n���ǪVy�������=m�]�I3�<����ء�R�M��t����W?~���r��P�u�K���p:_�a��f��]���[�"��M13M��9d��T�gL�0�gC��T����?g�flz5"�7
�	ԩ������U�,���>_���n<U�xG�"�z���jJ�FT[�hc�j��R�����Fd�K5����ņd
9�6TI�7-ſQ)�;"����?�'<7��9�{��B���Wq�$�	A�)R���J)��m�K�Q�������j�$��kUI�]͔Guɉ��_lQ� �#�>��L�"TA��bnN�
*iT�.����!�|I��&5����@���� �'�~_���Y�j��ēNH�̣d� F0>`�A=z�i��Jk42�8����ˋ#F�>xTӐc���YV9\�+����o��Y\=CIn�x �C����������h^<2���_�G1�<k%�Ǟ�L��!>�u����|��AR�>+�p��5��ף"���4�e��L��e�ւ[uc���|Lk �x�ׯ_���\�B�ɖ�TΩ��u7���\�M��8���M���������H���ש%+@�Y}x8��l|�p���z�d�����dFO��]\���)5b��Rtq�B��U��b�'�i�
�C����	�h@v��{o�gN0(rs6�=�9{�&3��1Z17�v'��.͈�0������^�s%�{�{V'��>�4s���i����$��r����V��^�]�K`�R[�U
s����<+p��qy��F�|�5�����Z�0E��A���x~��i��l90�:�I� 3��&<|��]3���C/$4����<_scǂ��}���3m:��f�_�>w0�AOI�3o
	%p�i�]��bYY����a�L󒙳-аI���=E����C��ô��e�q�����)��_^�1���M{N7����ks��M#Jl��2����qP�M���\!�<.�|<f�ya���CH��jf����}hB����a�A�����L=�G�꾶���TZ�B�1��"��A��n|F�9S�O@��a�ϵIr�黔sN�C������[a��6�p��Dubl�'�2��ӶN��D"����}!�-%ǌDU5Oym��A��J���X���*٩�3�i4�3�CS}ƚ�����^����t�u��f����ˬ��9��n\
1{\4��/4�F��M�����pS��5�0�Ʃ�3����j(U:gEĢLҋnU�A��1���{�pƆBV�VC`��"�����B'�++��Ў�C��?~������pfj��n�,7�M�<hXN�ѝ=D���51���׃Q%6��m�?>�Դiw���n(��u��g�����z8� ��FD�����^�;��,F;�T�� LàU�5�(��-��r8B��^�9\�il��|�v�@i��5��7^��P���2������9�~v������m�|��8��2X=�ʞ��P��euPxtr4à�[�޸t�Z�Z�qEײ6�o�.�q`b�c4W�T���½9��U��w�fmR?<�X���#_�F[�wm��i�ML����ГCj��dw�-9�P��19����YZZk΋���<��H��Y�;������6�E���m��b��Ҿ�d��ǚ�i�;6��6t��	\����$�e��3�N�4Q^�β���୪w�q%�Pq�.E�3�̼Ff��j��]��K4^�m�Çn[��.H����Q���Y��^wY�:���(������<�!���j�ǅ�/������k�^8�?sb0A� 'Й-�{��)�.�y�E�)u�n������8=���~vL�P@"�,����%,���I�A6x��iH����v�0���E�,~F ݂l���1 Yed�G��)Ue���<�{�`�v4!o���n��!��i�Z��s��:ˣ9x:��Y��X����6 ��J�ƃ�uRd�}'��ܙqxZ���8�T����w$����L���Ȝ!�	�z)bdظ��3TJ�K}�U�	P���mò�Nd���ύ��l��zl�-@������a-G#�H��� ֔�Mc��ʘI/3c>��63�Y�	�n麄
�edc����-���;)��'���>#����=BZ���k�J�c��,���H/��:�#s�r�vl#�@�N:͈�4β�C��5q:R*_42`��vZ�{�B�f,H��8���N�A��ҵGJ�^��0�8IA AY^Y�������E�����lP>�����^,�&��ʝ��wHi��Y����s�!��t��%���O����`��#K�x��l?)"�����ebm8��V��[nv���9>�R�vI������Ꮟ @k�U�n>�Je3B�%c��X)`���e
�f �M���Õ�(lukX�ȶ;n��H[��4����� ��`���3R[c~����Te͚��fR4˔4/�������?`�H���V���>F��ږ����l�q����
�:Q����dBCW�>36V�W�;oA���n%��>끙v�N�2���GŬYM���s��3Ҩ<�hӢ��)� �v�HW� ������O��8i6�ܽ/��f(mj(]�w�}�b��^{��0������n)��PQү����[��<'���z�w���Hu㑐;%��P��$bG���'bVi�- �[���#���_U�]�"���>�{0��%iHwHm�Nr�:Q�23��k?����`���~<9�hɪ����(�	�tS#{?�%���1�0C?�����6)b]�#x$�mg�7N���La���"#
�E�E����[d!qM�����a)`3s�����z�X�`3hfX+��j��13��5�La���zq6j+���1���H��u��t��\O�-'_[#a��oǷq/�:���n�9ع6�%��>{��V��M=Ⓗ�|Ƅ��3V���o�k��~�ؐ����`h��~݉��XҴ�"����B���¦B��u�������x�Z�y�����tHKS#��f,��o�u[;�m�[t�5%�!���߾��I���A�]�i)�X�M����>������6~�U�j��ƙѺ3Fm�t*��� ��q�:�@#���4a8i�9O���.=�i�[�����*CsqCf��%�h4<�a4.x�J7]���&�ϟ5��V�:öV�R;jګ����s�gv�a��z�`	��A*���T3%�^t�'a`si�%���&d�[t�ϗ,�<������&ɤ�=Ǧ����5yKk�ɦ)��Ĭ��dS��,6�R�'�dP"���}`�8����������o�;"���� ��=�"{��ŃfEy}9�y�Z��2����X+iF��#��6{��Y1.��[���l�r�2k䦹�O�+tW���焙օx���i?�r��f"D��I����51�i�����9�oL�.��뗀U��� ���/ |�Q%�T�,�h�tg#�ޜd&&e�|�Ʈc�*�=����ܘkS$Ęӫ��O��v��Q��'Lt�%����IHk��A��}����D��;�S���Hk�]sû�eg��L20���5Uv�p��H��{��$�-6P@I�]x[;+|�2I���'^�\w��
����dt(r(ˤ+���X��7дF�B�ɀq-��9�v��� �52(�<�T��컃��#�6�Y�?�c���=u���"�`��zM5���0�v@ P|�v�ػ3�_��Ee�2d�N?�����U�g�8P�\�H�7�jm|��e����S�����wؔ��]m+igN�Aj�>�Qgv�*������_������P����aݸ=����,��ۿ.�v�&G���f5�YW�V�M;��e��9E/�����-pu4z����%�(�i��~����XO�Lf��:��6��wb��1K�v������C鏃\�����޽����L�*����b|�O�?������NSXz�b=A�R�dʵ�Q��Rlc�������9��9�\��&��Hh���۴jY+=�Ը
���qB'M=�=�k���x:�L|��c���Fxg��:wAtG�7������ԯ��)���^�:z(!��Q�͘c�S]��@{w���3��f~P'���\ߑׯ����hl7�S=I?Dz���.nT�1���31H���!O�jW7Gi�%,����#�{�˼��� ZZ��W�P�_q�8Xf|�y��3�?Gv�q�ɤ�12�1R+%�Ѵ�kHM2#}�F`��WP��x#b;84J����Ÿ�0�Q�������DF�������}�Ph�qPE��]��8��C�l�,��[�I�����/�Z^�Z��FV�U޷�J���Y�� �ݷp����Ru���4���v���-��{7Cl����C�+�t�)�xNg�lz�*'=�`�g�?}I���0㰬��K6KuK��1�l�n�W�,�0Y-r�{�~�f�>o�Ћk������B�L��2��7=�HϚE�Lt�d�9|`��P��+b�]2mj�f�C�cN��#	�N}���\*~)�1�<z�V�<�F0M�V�sF�a/w��{e��˺�F��t��SҠ�E��%����5B���&��$��+K�QR��*�����=`8�H���&�%�"�������u���n7'0��B��vh�������WX�9���ȑ'_s̱o6���/P��v+6X�;,Z� �g��孊��y�=7�����Qp�i�귺['���9�I��m�ֳ���;���!' ��A0���F��_!� Z�[K��S�~���/a�ۅ�}���~���,����ʓ�Ԫ�-*>�As�a ��������ޜku7`�����gr�����Z����qݘs�a@}�n5MM6f9�cm�σ���l�����*�#����ܰ�D	������P����S�LUς)�L���^�5���ʊ7��[e��He�m�ihHҧ��>��}}N��k�15w�~�d�7��p\���Qjj�%��{��P�t��Q�P=�ȱ9V'���M����4�C�9͛&V���"�I<���z������u�����k��8��#�ҊL��v��C��l�G��x�sZ�B����@���x�%�OG��W:��u9�z��BU삇���u���@fX_�9�酓�\����.�6�<U2n�y�"C�شȀPb�$'<���]ޘ"� 8��ec���������ߙ��Nq�id]��\5���͡��ղl��q���^b3��$��Y��Rw��EC�S��7(�b=�z��uMI51���;�ͧ�W�0b�V��g�,�z����0���,A����C���<�dV��\(�>|�������u%�vpŖ(�L��ӈn�&�F?L�����~/�l�~%�i��Аk�x�#)a�r�rȃkq��b�{�'��k3������C��j'L�6o1Ew�M4w2L�	��� ���hnĕ	�R�!R��B��f�a����D��^��qT!�(n���(�/\�5��1)@���.�5	��1�/�:]BYg�Ȩn��@��l�!R���ՐG��L��ݥ�H�d����z��=�. X-�*Ӝ1���x/�t��d��͈SZ����Y���|δ�3p��8��#.�\J�*eUK%���-��qd�()�a}��̚�L:�E?�H���I^��a�7�'}O)��d���iR�Tf�z��͈�BN�c�;�F���?���
���1	���2�%sμE���>G��,%���f�L�ˋj`{^�)��{<���xDW��-2�e�xxq�e������Ǻ��i��Lь�C<̍�cY��և��M�k�����b�8��w�ky�X+��hd�F�s:�}=�J��ԅ�?;��P�1k�-���~���{����V%��_���#pd��7y�j^Z�6����D��qih^�J-YyCދ��g� \/l�NI�µX`{ JyzE<�x*�TJ;ՙG��kC��+���ԜS!ƒڊ@�Ϙ��1<������C���1�7d�hV�*�ką�MԸ�k��%/��ן��j���>#-y!҉f���x�"��k��� �NBq�J�
�QF̤���ZeR�d��"iX��j�̡X�?�B� m#W�^��&p]�X�wV�6Nl�8��C_g)-��-K���Afㆰ/{~�A�����0� 7/�)c�-�ʮ,62)4�jg}��}v�1��WHro����,�׸w������<׸+�����鐝�#����i�;݊�ʱ$��/�Gl�qS*�Ld���r�N�6�b�?��n���B�3�%�˯����r���}���D4��@�'M�r����VU�F�D0:�˚��I#�#(Tä��Kn����f|tM�;�[��[��x���+]����?�����~� �7G!7Ɏ�iБ�P[*������WI��'A��sϫ�v60��=,�u���>�S�+a�j
*����a�vŬK��:�I�e����,�[�CW�O"��8y��Y��@�g��^�4����5���Д�
��!���Z�'&�ݬ�:�8^����ܿ�]����A������{*"�*��$����ˉ%�G����+��!��lz��녃x&�A���/��z	x!M�j.��6���JN�18r7�� �.��$����ٸ\cu�Y�Űr&}t_ů������(��:M���Hhd{�# �t���-� ����-�5�#^���9��2���7N~hpHoH����==kP��>���pP!2!����8��Q̮�4��;�C���X�z�3��`�����[�fѡ��cV�Tp�a��\�1�T,��Q"�Q������M�n��������m��;�d[ra�N�������3.�������͟x�at� ��V�R�VR���*~z<�q2g@�!���~^ ��z{YF�:�mz���Kpzeds�w4���>�1,��>,v�Zv|�]0�7Ŀ�j�&�����'7�ڦZd�zB����0锜w��2[�]�n4�4>�g�;��N�Pu҅7}�wRυMao�ƀX������c/ը^U=���_������&)�D�C9:���ֽg����Ɔ؁g��#4�-�uB{5v��+���!G�DY"��1�F�i��P���r�۾�Ħ4�]6Y�;������N�Ğ��*$����3J�5��Sx��~��(��c�^gN����l���[�ء5����������υ��^�;����⠒J���5
�UB�d������{uӬ��nm��/��hM��d�l�ֵ[�C�a�AqV��I΄�����yǔx��U����;�zF��ό9H�j�����z�>���������F3g35�Tr`���C��^_ϊ`���&��I�kCI���Y����-��ki*�ɞ��]��>g�M��6�c�`��V:�.yHuR[F�ܶ)3�x��{�>`�W�_?�$�+p�]����#NkPJ�V{L̶f��~���l��z_��
6 �A���\Ԏ����J��g��h��t�_��.7�8>N�r\##�A��4S�H"�Z�E�ĿXwfn
W�#5��(�K���Q�t�����ڛ��63S����l�,p��BVw�5Y�y�?ϻAn��A�\d�X;��-���*j �#�8���h}{||�S�QY[�_V�g�2|u�W����3ز#\��0
j8�i��{3i�6i"8o���8�Х��\��F5:�Į�����2�tz����1k��͢�V��xt�\Z�4�HOT�q�Fj��{@EK�W��i�V��=m_�8�no�|l.h�9�V�������pA#>���(c�L\Ψ��&�U�}��C+�N{_UU�=�����8F��Z`xI1�0�p+A,��;�I�2]�P�6��7	�9pV/XO�e��d/& ����բ�]�қ�!���zP�����0jG���mL*Ⱥ���dm�/ ��fV����8��F�l�t�k��G�XxZ|�^�����J�nr�)8}��k���Y�X5���-�{H��t����3� ���N��|�I6G���;8���b-A�Z��$52��x)Q-I\e~cc�daFmG��Q��R�*1����F���}t�=�oV&u+����LR@T�ڬƣU~ �Kڲ�0WA��]�e<N�D)��
u�:���I���|"n�Z�4�����=E��2�b6�\^  �[%�}%�;X�I��e�+�sx#��9d�o�8�PUq$L="��_>�l;H9���D��ob\�LOE~��%Tt�t�b;�а��	�'�����$������~Şϻ���O���`b<��VZC����hj$*�r�X=P�c���/����K�r��ʿ}�a�8�0�n�<�@��;�9콹9�m\��l�&8c��HVM�e:W�h�5Č�P۝�M���{�����"�wi�C@-:q�%kt���Nt#�N,wB���|��:�D>�������'�=�$K�$1$"2�XW5�r��;|  ��?�Nng���Y�d�����{d�άr6���2���nn���Z:��ٔo�d$��-�R�kz~5/CD����c�B�����T���Y�s��Wwp�@��8�	�A
�hRr)1V�V�����&�>��|,t��4%�^R����
��VM��� ��[F9��=�A�3�#�ͭE�}6Ʋ�8J���V{bun*FOp�q��TG^WȊ�mQ�a,Ȯ�1�d�\a���ZT�2[!��Ї�����9߾5�M*���1���cR8`�|�*|����*���b��3��s7�c����J~=϶�a��uU6_�!5��V9Gqu#�R��u5ӥ�+D@f���)	�)CW���2�"��IK��b���߷��]$��hҦlq�I�(5|i�Ä�+���J����QL�!a���/�CUd�
3�z�0�����0�
��B~��M����CH'w{Q�z����������7�.�%~����?�̽��+X/Q��ǵ�,39��Ob�<C��Xl�����陑
�g��)ͅ?��.%���fQF^w2�z���._N�o�����!����Ϸ��26��E��2�.��^ #�>�7��{��h׿��m�>�%<;��$B�4�l�puAn;��Q2������3ǂ�G��
,*:��XD8���C�j^հ���2d<�%���u ���U�����5�@��#Ow/���U)�� �q�>�v�N1,���Dխ]26 ��j�V�>� ��vmq��$J���}�;���<ff`�'���`{�,�i�5�
uV����U�v�<aD��ߞE�@�on��)b��F|��ny���y�}���k����/�R�Iה�TI.���s��S��w1�n3!��\4�F�c</��0W���GR����5�!���+�5%�����3��A���A�mf^��3�u�C���'1S&A��,k��:P2���F���7q�e@yV8��.u�K��]f�E���S1�)���OmF���5�67+�,l��c�`���2K��)R�gm6)����t�R���1��zqH}�{�%`l�Ab��DK��>ŔgQ&R\E�T����u�"�4K;*�?{u�X+�f"���˵p�2�Ah�����R4�4����(>n���!�� myb_��(%��W�v��uv�Đ��j״+°����$�C�X�U�M���ʹ��ar�*M
v����E����oʗ_}U����f"!�����Kcf������t�2�X��3�g�A��].6ǪER�|�{�[i>~.T��t�e�ud���ͷ�w1�Ry��TBõ?+�DpO�w�j��=�Z���Xr�!	��,�oe�T��7�1נ頱�e�i�~AS�kf���4Y[��셰z����ɘ��ʲWң��4�6�3�<�wr��}��_I՟VѸ'v;�:�CI�ڽ�b١�Y�>3R�\`�
$�]'O�Pm�\/1�6���\"(��P�T`����h>0X�t}�cr�D|I[yf�S.�i`?�n�!�N�۬�ﲴ*���O�1��Q����k�R���g����]��t�W�LN�� 6U��HTDv�k#��_�����
E�U�+��%����1�Hky�j���3��mR�w�Tα���}쎕
���42G�#����i{��1�c�XV�w]�Fd�z�����)hR�ؘ\�ѹ�Pp�6��@dC��?�<H�_~��p�.�'�`�lh���.���6f�����rCo������ ��,�r�]���'��^�q-���(���:{/1>8�j'��KEN�<��^�/.��Fp�ȫ��E �I@�p����&�"��b�
�4S���e����i�{��WG��iF���?��RD�/�b����3@�ˮ����zftrk;����EU\���ILZ�(�)n�5.ɟ(�?��`���t	��Q��j6�@#��Pu)��W��bJ�*�ոp�x{�nB5�c��[���6�3J��8�����esg�AtI~f�g��R�g�����$�E��}ۋ��2<)������Nn��_Ӕ�e�:5^Gi�h��C>"�ɱC0���!(|��Z�
�*�J���]Փ>`� l�zaQiة�!c�s�#����eá��)�㺤GLN��U ��r٥��h�Y��c�
T��_ �~�eS��'�ܝN�����Y��s�c-V��}]'}�1�e�K2��Px���ShA��鮀@�&&���cb��H����F+o��@�Z�>���^���^��w����(�4O?�r �Y=|�Pt���Iy���`:�@,��� 0Zx?A���HS� B�<�X�do��T��@Rr��t��l�@��1��P��Ϻ��)����>��a����>���2�����賙U�\�}���^��m���?�M��	�ҮN�[��n%V��J�馕�7�J3.����ԤL����Q�����F	6���	��W9^����a�9N$����T~ `A"|>)1E��@��X��$�!;��4?$	��]d9�%}�}=��^�@VR���1I���1�Z�Q����<��#���|C!8�����p ��)���y��dJ����D�a�'��SG>�"�$ ��Z�P�r�Za��'IJ\�_}�uy���?6���(Rr��nxP�T���Dd�] )�HG}G��:!��k���4��W� 3�E&q�C�Al��i�vb�̂0��$���#uW�'U
�����^�d�Oܲ�N���8T�b|��wܿ��ǐW��K:���գ��)�+3�]�W�N� J��B� Ho��5�#��X�H�T��pS��ٳ�K'�`e"������]%ܻZsu[㝼��KWW7���j����G�Χ������SoI̒|�zc���'Ƙ�z��}<R5>�m�3�?7��wv�Jxٳ$%͈"�3F3d���0S..���6(����H�FJLż��i�]�vĄ�}��j��OC�G�6���W�6��U��=`��c�-���$-�^�S(�������I��z��Sb����7&EۊظVu4��J$,�(�d��	���Z��5�Ȯ������6���R�~��uh޼y]����}�P�g⣲�� �!e.�]qI_��8�ҟ���%戓�JUW�釡��la1���"��\��)鯂Z�{B^.($���ߙ�EtV�n^i�ٸ�iX��i�s�1{�ݻ�K�=��f[��a��݉��2��4WQ�vc�|:'t�����F��Yȗ�$�A�g��lpkۙۃ
�O:ݖ��/>dYZ���c%�fs�Iy̞�O0E�р����db5J�����Uoƒ}�j�S]3Nv����$��I��{\��mZP+o�{�IU�gNC`E�y~/y���HP�e����`�1nܜ���t���w����~���3���b������ǜ
��)'��t:j�}]�ᦅU�,�k�~���n���  Y�$��UM� W�pgp��e��"1L6��@?3�DJ�Bl���la`��8QW�k�-�r\��.�.rd�]:�Ϛ~��1gy���_|Y���?�?��O�Tr3(U��%0��\q��&Z�p�օ����C�h����a�I�dp"�۵��U�����V��5�n)�գ��3�k������Tum��8~}�7�T*<��g�fF����dS�f߮��F;�p�Qѫd��t��l�D���Pzᒻݒ� y���fե{p�
�n�X���J�2ةՍ٪�asMR�Xq].&洷�	��6�R�X��t:�����4��t��}ڀ�C��,Hc#͟�H皑*史8?춱�}r���',6B$��,'�lD�v7uЇ�mt��|
���Sf�P��v���e������b��/>�r��w��%�����sp�t�r�n��_6���!p���5	/r��0�V���[���}8>^ܤ��L����M/���#1>w��Ƶ6�9'�<gl(����(�\���M������f��t>p�����++��É���v���G���e�/�b �o���M�ԴZE��JNnН�Ì��d^J��g���;7F����d!���J��`�� s��K�y��Խ�58hڪ�Dq�555
�tg�p�%�L!��(�1T�� �� ���9��%v潦�d5��>�2 ق��x���y��=	�
]�zt��I�S&�~5�P_���{�6T���k�7&����CO���3�,Ϯ�^��PQ�8ϱ��(�d��CN#d�h.��)���(a�s�����ݭ��a��ګt�}R�g!�$���:w��RiF�q��NJA�ٶ���:��+&%��͖:�kl�7b�����T�o��5;YS�ҍ7dor�,�� x� �]<�����z�d7W�L4�ʪ��vP����C��t��
ݶ\5���R�����w
�AX� ;+��>����X�*�Q�d1[L�"������`yˡ�(�>Kc �E`�>���Gy����F(�o��_~�e���Ct��d2�r����Z89Ǚ��Z��'��˂��o���&�M)]�Ъm�:щ֚qF��B��YdUx>������Kz���=��(�l��)�#V�ڭ�b�I���"��`��LG�Ԁ� Z�Eާ�tUF�1]s%�,�{�U����c�b�@7�?���}7\f��R���*/�#�]
�X̥���ZE�<�X(�b�\�Sƥ%0}�����;U���!�;fN'�v&��|�����ϧ_c�'_��T��ʵ} vI��Xfv������.��D���/p!�� ���x7��5���oI�o�wڬ⡜P���B �%I�[m(!��4Y`�����Ƨ:N���A�6HD���:�Yf��i,�Hb�S7�q݃l��61�;�Dn�#�J�ɫ0O�r(��l@
���	c�^L�,����:��ˑYd�n���w�Cd��}������hP���"�qTBȈN}~�s�9���X��P��n8ĵ��k�����p7w���%;�Y��ӎ*��Щ�� ��/��u���(�LA�F6�ݐ�7JI��#��������U2GSe<^σ+�Ę
(�-�[��y����v���Yڡ6L����x� ��`腁Q��M)9^�Q6��~UE�#�E��R3��Ś�#�� T�b|����>�]f�����R�xiYK&O�x6*�w/�6j^6�ڿ�w�i -Z\n$�x��?���c7�"�i����p�&�H_���fѤ��ؕ�-g).�[a����˙<�H}�ścS�
���Ac^2jL�zB���*lL
�:�p��3P3o���>p���o�^{�Sӕ�q4�J�X`5X�
��(�p��L�&;
6Qg~V#/ؔ���.�R�&��i_���iX���]|�8|� !��Bbd�. '�j_n���7[����X���������F�e�����V����+|�;V�Zx�w�������~r��Y��rM����t���I�]í�˛����߽�o)(g���pEљȼ�U�=p���Jc�e1)@�Ɂ.�kd龜q}�y�/l�̟�ا��Y�I@�,��q�s:(8[�dW[jv.�=���sb���?�X;sD�6���0��Z�o/��I��B�Xjѡ�l�V̲�j6�/���a������:-U��x���~WZ!�� ��K��fZ���������_|i�`�^"2QFw_�q����.��i/����t'��`-��`�c���g��Ѓ��E]=�j��z��KN M�����cu�c��S�T�l�>U�}"����#���x��!H��,K2^
Q*�8�#�M���1cJK�15�������#���y�0���bk�<���dU62I��uh#�%�:���>�����TW��88�8��|��|�����o�)���-+e��.��b�t'=Җf���ϣ�Og�47<R,F�LuS������ˬ�,'`���';K�Q��B''��Fq�l�-� W��������]�(��^!���X��KU�ծ8+�#�&M�9!p&�{vZ9wn���!nP%�ǞX�=�c�h`w(5a�#lU&�$-��0W���8y�J�t�$W�Άw�)�z��:��ý\'���W�UP�ɫU�}c��9�yD���覥��P������i@힆�� �Ͽh5���."�%��O�2zi���.���w�4x֤Ƒ��6��60d�l <$Ԧ5q!kS. �g`>��m"�M��lw��5?��շz��9u�N[���6{,��:Q4��+=e8�h�J;����E�q'�D��1��q�>(H��ӡ����2;M"��Y�8zӒ��DVv�7ؚ���X�ꏸZ@P�Jtj������W�/�,_��H���#��lo��X(�}8e��'9Z��M�e�����Xh]�V\b��5���5�+=��@y}E��gG\3>���N�Tv�#�-�����N)�7.�"��de�w,K�JO�o�����/���['�����V��A���-4⢍�f�52��0	�\�������L}�OZP�n���V46� �1�eQ�}Ⱦ��ȠI؅:Ʀ���u<o����d�p�oVezd#
�Q�k��>a-6*���+�{�Z��e@-������I6{�D� � ً������]k�fr�SŌ�3>�� �5&���o\��=�Qr�{��Y�.�L�o9_%ݖ=l�:n>��P"G�D�nܨ��	������H�8f��kh�~�)V!x;��+�vj(�B.>�3*��!Q�J��}�4�F.d�M����o�ʼ��t�Bz�����������ge�T/�H�����eL&}��oが�����&r��h���J>b�R�Q�I��#X�%��	ZWBL5k1¥~� �g|ཪ�ws�&ɵ��xU^��yL9�M��3a��ͷ�ˀ5��6��<8h�bnqN�lȞa��e�o߽�.�?���H�;4	�:i�Ƹ\����]�A`]=�.������(�h�.�`�Ǟ�>0�R���k5ՌqY2�ζپ��E?1N����-Gpc�e��Y
�s�>�zxo�ў,�m���8�{v�����9���:^�$�^�Y�
�m��$��K����0%�7J>8�G�f���_�72��aB�0>Q����)��Z��ΰ	ئ��*�q�Ş%pB�*6EH�o�qh��@?*0/�'~H����>���b�	1���r�H���r27~_�/b�D�����C�q��K�l@} �`��k'�6�OĵL/�~����Y��f1Q�C���B�j��{̝��Ed��~�m�/�KR��p�׃�w��x܆�2�un�J�?H�"�In��r%%�:g3d	�NQ�u�.����GM0am2#�TȜ�D:��^U �'���9,�HƉ�ב��),d���Ͻ������~��
�T��������;	9����C�Uc�&��;������b�V�������3o���DՓ	�jRЀ-�0���{h
l��W�Y������/��]K�����ۺ��J���^=4��Ÿ�I�ԈFs�]�j���3K���灔�88�q�r�2E�L�v�a�ՓT�̳��!}��6�dŬD�&k��䚷�Ժ*F0Q�/�p6MS-�"��{<��av�n�!&DzbNv+�f�y��:��/;����Jw��Eb�KJ���d�8�0��|�m������w���i��^k�+!p�:lg�Ц�T:-FJ5L�'�rlF�8^���'y��)��s�gqo ����#��S�3)Ll�yD��c`�h�{� � �&�\g}vO����ʔi݅UG`�UZ��뗋��� VQo��cε��1P�n��g�s' 	�'�L z�f�9x�&l�,�}��e����{�D=�_��iw��"�7lJ�H�=f�6��'�$��W�#�"�A�C{�*�Ҍ+�+��4ߙ�ui=��W�?kO�f��@ox�� &`5Nu]�-zUN����6걓��;�Z��^i'���e^�f��P�eD�'�Ԙ���[	���l�G��#�eǌ�s��dɸ� Ύ"6p�l���Ml�lH�FT/��|�X\�sl\|������Ѱ	_�+5%f)�ω��w�(B7Qe&�*��9��43�����J�Hjj�n7ʚ���q�Vå3��97%(���jZ�Օ(��H'�5��(,�kS"!Ԛ���,Ia;1�ƴ��i8RT�XU�����1'��W_Ei��3	)gٮN8�����n��`��(�þ��j��f�F����饨Jxɜ1��]�1��6���D����d)���������>�� 'R\'��P�Qk�?���=�� l��O?m��?"�����/��x��V�7џ����s���}W�pks�������5̜<3HUq�>3��Kb�e''�Eb ܃{x�B���W�yj(f��x5�Di���ke���������>�	�Á���0Ǌwנ�O�~��TN|~��jgtL]��eT��@����@ʧ�ԏr��ޤ}}ĩ{:�EFc&|�����b玞I���<�v��1�����1��n��+�n�<z-4O/����x�'��K��\ѿi��zՌn+�� �N~�Zdhp���e(�E#:o����i���򔿍������J�� �$�[nrQg�1���T.f�Cv�9#-�(�P�&�����>pb�2��G���������W_�"�-RDQ�#y�75VZ�u7�vR�w���n�aټ+� X>S��T;vd=���>Cq���	�f�rs*nYYF�/����Q�w�u��s��ױ��P�X'���w�`�������DE@���\8�`M��,�df��<����f�x�b\�u������ ��/Q�@�p�����z ϢҘ罻��{mHJB|Ʊ"�Z���Y"	�$�N);�hLo�-�)v�X�j��^����5�aX)\�8]xyP\6��D����7�&(��'�3��9y�TJN�SZ��+gZ"���El;dO�R��V�.:�A[��;C�DXȸcp.]���s�h 5d�s�X�.Iڴ��wv��M��l��qJh� cb1XX�������IE@8��.3X�ۄ�5T�e�p���}ƙ�}Z<ur{�^��U�x�?�}�0�s��X�HX�gN�`@��C���u4���6��/o)k=�	 ?޾{��CfC��+ )Ȟ�+�+o6C(�n,�[e�l�)�-�b��Y�4bcv�F-�_�Y��5G�����	3c��f�� ��?��K�e;P���6�d��pܴ���>`5O�=�cvW�actUF������$�2���k��/�IЍ�R�=k��	U��b�>�Q�OVIS�ꈷ����z0e囈d��<{�����1u#�����Y�������{͇���<������D�����_W5.#�����k�i0��cvi����Gc�C�5���:�x�UŅ`G�����9/:;�Ke ��MЏ\��TK�dL���8nx�����5ʗ���ZO����~t�ƀT�����_��x�5kX9N2�a����<��)�րot��'RJ��£�������@\�P��dH�^A�Axɉ<h�A�c*��i�@�Zt6I�;�E���\�cˮt玴)2�י�>���*�s��]
��9`8�U(��!G(}�����Ҡ(�̝�\�u��*d]�@αF��?��c������-+���^�4.M�<���g��?�e(|�Ӊ	Fe4l���:��}��[\PZ�����N[��M�&��9�Ιz6�p�pm"�H���F�����{��m�ջ̦s5� `9���e��೸���/ۨpW8m	B�ìTR�*������68����k�S�Q	5���k������L���h�!�\CZI���2,# ��Œ>ݱ����9��f�Y�:N~x��׻�2'����!�+p�@�!ށ�j�� �}�O�g�I��>�Ն�N"J�[����z��{۞��jt�/�UyM��G��~�"���1��N�����X;�����h]p�ʘ�g�U4SR�<CH���N҅���,���3i��%�R`1 �$���M"�Ɛ�K>|��>i8����ߘ�;�'����*%[�* �҇x�9�}�#]����z��2�3É�P� ��؈$�)U'�+pA��i=M�G\���;�2�N�a��Y`���O����e���E�F��|s1��.���7����B�e㎸+��1�����i{0\l�3��������hx͕,�@�u]�������/_�d��&���:����9I�ґY������a��Y!#8Q`d�ޓ��@��I�r�ќsF��R�k����EpmΨHk0��uU��"�6�4�I	�#t:#�*724tn߽���77Cv���1��	0ɔEF
Z̐�Q��5K�;�"#����iv��(���"#�e�$��I ���q�C��6+2�/>�"v=������b!E�&�[]�	�}�b��/����|�͗A{y��m8:bA}��Eཻ���z˓JM�L�9�`"#b�O[�q�,1���)u��������\�S��v�M̩���r��H���Ў��Rͥ��gB ��N&w�!��;�q7�B�(�qH�w�c�v$��c�,�5���o�)�|�m<§�l-�s���������G�@��^�%YjC~�+�d'�UpH�8 Y�<��8X(�� �pO��\�����%^��l~���o񖀓����D��=�e��Y[��MS���>�d�Q5���|NfμL�;�&��-��~�_AISƏ�#H�1Xq��E�ac�������%�|�x�c2)�:�7�Pz�\=<��ڍ����dŌ15�>qѧ��E��ׁ��������M�L�s���R��%7}M�;��A����j�n�^a��'F�"G�]�>QLt�W�e)�Ow��%��;��q3� �6sBE�X[e'<4���U⺌�>�i�6�Ȕ��9��3�P��(2(��hT@�~;X�&5�A�oS��H4t�S�R6*���&r%�^($BE*ro��/��j���;	�~'A�6�dL%�;�Lc���.��v9�)����DWׄhd.�ǝ���Cy�&���܅���A����8�8���,	����W]3oؠ�a�3l=�%d����Ę�-6��|ƴ��3N�	qݐ \؝��y�=�"C�����%n��QǺfv���Q�/k̳���3Ձ�#F���e׃ʊ� �dc�Ɇ^*���c��.1�[yM�0�]�]S�;tSwH���h���^B�pC�J%68	���ۀl�l8�:�ٍD"��b��r���խP�����x�/y��'��40���Uj][�S��h+*�z;�c�]��q2�$C�(7*��i�e��yJoo�$��]f�Vw
���f8O�{�/�&V}�%$ �)	'	�P�v>oA.2?����@L?K�<Kx�����6*�aO^���c�m�=%��(��6�����@�Rѡ'9�U�a<�gM>�0�U��a�I�Mς%���>,���D�w�G��DؙkԴ�|�����$ �g=Ŷ���1f���yC���4ixU���C����۳�����l-��
ݛ��t!hp�P;����_�ں"�B�K^��*#p�����*���P2�����>��/# ����cв7] ��d���{_X��@�Ή��O��N}�IJYUSw栆Dw|Y���W�К$�~��\8F��'ڤ,ܙt8
\��e5��$����z�����;&A�*q�8�� �Em��qφ����X=�;&#��y���E ��X���M�&vmm���7�i �i���)y�R�(li=��uɓ�4� �����MR�	n�jY�^O�^=��,��LA�R�"�g�E���wB2R�0��y�ir��5OF��wZ8(7V�����2O�YI�����):�;np�����Mx������$%��Qn����L�:GYW����ӹ�ٝ,W,\���Q_m�84�P���C�	�,���M�RK�%2R9����m�RǸ�mpFQ���h� ��-�e(*}��7D*ቩ�� 9���*��{���q�{Rs�q�������V8aW!,�$���⻾y�yr(��#p��᧟&�`�;0����a ��{`&���Q�S@���$z�j�[�2t�bϨu������:%�m=ȆI=�'	��|�a�5v$��kg<�d�q����\<G`�A��ljH�Ӻ��Hs���I����D{���5�k���P�'��C��Ω]O#B�{����]��[h�hئ����'a���8}�I��i�H�t�bS`Nк�^�(�M˱
O!f��C���a�T]��`�/	���<�T�oŋ#@�x�d�����>Ep�N��:�u�cy�����Y�|��R�*Kf�.��W���!��e`���w��p���� ��#2��^�[�g��,�ҀjΚZٍ��0��Ԟ��x�EG{-�Y��6���*w!�KK���f�����e�e��#����ct�Ew�ꡌ��a��PX���������If�1�/��ux\�k��	6���i��L�SU�"�(�r��-Cf�ʇ"�!�h������Hh��K󮛳B;K��a|��%'Q��\Y�CJ���&5����ʖ���;�p�y,��r���s�a:h8��N���E�ǆs��I�3n��p���.�gi�I-cW�N�Fp�M5Z�w�q�:��б��Z*?����^�{�{m�,���|�6#5��%�>��ul�"�v�N__�OE[e�����/�*�e,�������US�CŧS��6�ZK�T���/�!D�8��6�s��Nc��������e�!zB5��6ے%l,��T���q��,Y{��yW�M���+�4��rf,S�N�@������-)B�Px'=
��Z�9B���,ߘ�x+��[j�&�^��O�d]��ԯ�D��È��,'�h��Ӂ�C�z��p���xĕ���@���8�u��a�,=�,�ӽ�K��޼��u@�u����	����+	���-�Z���s�t�Տ�6��fS�e@���ﶬyˊ�����T\O��������q��޲$f��;( ��Y�JW��gk�����f~?|��t�5/5�hK%���p+= 5L�LLѠ6
���CY4�y7�?|��ho�X��^u���g��;[���2W���y|��O��oj�	��3E�� ��܃���[]�-V;g�p��;@ਦ�Ms�r2�.5��6��-U�OVY/C��@�]�Z�S FMXx��~'>]i����>��fe�&K���%��OC�nM���
�{�w' ���{��+��Xl.
/\���h�*U��@36GX��s^�1$��9�˴�����TeG�4�:�G�����ɻ-(�����n�}�GȂl�� �e�r{�.!p�}����0��Ha���`,:��ļ6>���%�v�&��&��b-�l(�Ӄ��I�+i��>)Ox�W[���5(J����D�Qd�Z{��(�����3l�����m\/t�����?~_ d��^�d$�W��!�6[v�kA�c���u�~4��n�n"����˯?She�8԰��q��A2��M�Q�|3��'�ظe�V�p�0ƺHD=��Γ��NZ��\�Ǩ����2��;��ǟq�$��pv�tS�j���jcٖ-\���b����t�<�:O��� �﷝�:&���U������慻9�Yk/"���A��G�O�������4�,��#�N<e�z��{�"�6�@ו�_�����T��T(
��i�?𪕸��,/�S���^.(\|4d,sM��yɌ�N�}�$�(Ё��n��o�S�L�?;�I�QG��'5nŋD�����\����P���R
��v;�����Y��s�T���n�x�F1b	�bd�_n~��WQ�Y����Y``�<�z����%*��Q��>�p�0xZx���>�|�����I���������c4��e���"�˟�����x6����θh��k���/�Ͽ�T~�������=�>����qm`��|�l10��5O�|زU�L�T�}e����W�A����57*���?������~�É%`��!�3|P۠B>W������3���٨&��"ړ���%����)�g쿸0R� ����4"F%��x��`�A��Iך���j8�,T����YL�NE�f�h�TI
��8D�ݥ��m�uEw�laPҖc~n7֘���Gkr�0��j��郒��L�ڮ��M]��?�G�@�}��wf�Q������3���2��i<P�>ޘ]=U֪uh/�*X�V�Sg"12�FJLt0��󒁗�W,�/�@�<ʼظ�/kH�m
A���%QB�U<w�h�%,9٥��C�Jg4��&=�P�������;��3�.OϮ��x����2Kټ'���T�  H�x��&���$�?�U o�C&l5�I�|���_|�Edh_m���_}8(7������dG��V0]�9uЧz6�`���m��~��ϣY����+������.\xǀ(pq8aF�6�pJ��!�,�SY���Ѕ����i�j)f�w{?*�A8(�4��xOyu6ga�3E\�q�UǬ��UQ�)�|�QT����B��v�i]�OaQ��R�b�N{�V����7V��U����
�k!�����~1`�=��AՕ�G�'�S�ޢI{Q���ā���d��>��şMݮ��_�������7Q7LK�l8�Y&6ǩ��P�]]GV����!H׀�8�|]8*׎�q����-�~&���S���ʊW��(;䃤�(.AN��{�r�g��b9��:�3!�<2�k�Eh����h.���,�� ȗ��D*��޽6�����c4���a,�����(�d�Q�5��KW��km�š��C̸:��4A4�~(3�C��^_�y� ��@I����/� ��쀋Ҏ�U|���B���wo# _p9�\2o�nd�����L���Q����c����s�1�9��;�3�-뒐�+&<�[T�<xԛ�O?q
h/�¶)�Ȥ�����b[����<T�A�B�?I�ד��MN7#1�x��CCV~�+�ݸ�ɹ�c���Zd�ۚ� �����5�jM`�E@T���/�����^�Yx��O����x~�,��&?Gmh�����hj7����n+uMG�V�	b�9��n�u����EY�45;�K}��@�����M�TǨ̫v����a(�+������
M��J���EAe�9a�p�TY�{\���R�cн���.�{�ۨ�s�|��0����.7��9l��Y]�fP.�]�0��/)���(�_o�:29,�yR']�w���w~�H-�F��)�x���5�Iu���c�r.�Ł����T+�S��=�-���Ki�7�̷=�Cku:��RK[d��(m������~��6���;�Qi��{�d�b�Q=��`���+3\��Е�{��qN��.uk!�{�	u��Z�����&��?�#&���b�~/��>�`���`0|H!�j7�"�o���C�k�u��!>/u.>}�Ďɝ�5�y���UtC_�F��#��ʹ���=}�G`��KT8&�m�jew07��z��{c�gJ�)y�u�� ��:�u�ΰ�:�Fw1X�'�<�l�3Eq��m��[� ��̬���wn�U=�5	�����FW�{'����k�h��Z�XT^�\���|n�y��e�g�kQL�ci����W���Xl�l5 y:��N���Fٱ�Y�W��;m�(�G�B��j'5g����˖������񚇄�]�J��l�������t���;9F =KWx����Z����6�|��mf���jb.{꽎�R��\o@G؎��U�@��Ӊ׿�-ց��;�c�2���6����x�g4�Pz#��?H�
����7�N�� \�nx�<f��s��cZS[�5f��k�'��X�P5�o�|���Y~}6Rq�� ��UҊ��lJ=���Ac���D኶k�!��ϳ�B��ؓg�#>�\�_B����k��L��T
c��O�ǵv�~߃�,NjRE�V8*���y��X^�����tN5��=�a���s����[/��U�c��`��m���Y���Tux�`��9�-J�|A�<(|XdO����8�iK���ԤEsQ�[y#�9��a�2��<�|p!#!aRp�7��R�ĝ�D�Ņ^���+ڌ����q��
D\�ܓ�H�HKL7��5R�Y�I�+_������p<^��J�ԡ��>m�� l�>t��C�^��Ț����;��
�?|���^�ad�UE��a�lt~u�a���g ���+���}��1 Pt���hL`�J�������&���@�/E��]�_���.dgo�3T��R���o"���ߕ���"J�z��}�R�SI�|C06�9G6H �/��!NP�)p�n���60WRs��hئ��5��;�������ot��ܻ����x�XCƌC�����:�����c|F�,���ͯ�i��t$K:�4=���?%�ӏ�	��f� 8J�gh���I'v��1�\�<�CPc���2���N�,���A�3���.�UnoN&�,h'�Yg��1=��x�`~52h�>q���"'���H���l��kD�X�x��b�cK֎L���u	1��`lNt56>�J���3��ZS��"�x�J�(/�Ag�lPۛ&��}�d��L�h�$����<	���i�,����g��G��~��������+N�л�0���+u�_�B�-�B�g�*cB#�0tK��i�M�@:*��: E������7Z��(����}���u���_#;5���lo����a@��A౏G�mSoµ��D'�X0J�%�|ڮ2�fF���z^��Hf�ȉ� ���3����������/.o>��|����g���At��
�>���_N�q�+6g`F�f�_~�EP��%A��.˫�S�NGX�q@a��7|���%�<�;�M���όJ���s����������L������o���E8 �Ò�*�"��ᅍ���$���������NN�?jk��YS{����R@��Y���4Df��z-�U2/J��X�%5��\u��@i�`���ԣ��6:ٸX+�"K2��i�B�E�X9���'�+;%mTCLիK�G�b`�xNz�h e����"ӵ��5�)Us�R$��jX�{$V�y�TbRy�r���2��XϢ���?B,�y2��[t��.#�"�'�3��x��ą����H��ڍ�g�YtӦh����씧|�rkm"�C`Y�f��;u�Bc)�y��O �]l���W׹@c�
�$�ӹf���D�o�	L��/>����F����~-�����= 5��n^<+_��P�"�2Q���=(#��� $��'�&�N�@Yʋ-��)��C�<�2�_~��@5��^����z_���������ٟL�tݮf�*��U���@
�R|�g�X�O��b��`��_�M7�弹'�zv|�Z�u�i��0f����SY�q]�˘͗�g�ЀV�g����������C@78،�#���A��޿-ϟ��%���!n���y��*�q`�'�eF]JzGE�N��(���hL���(T�����!"�h&�j ����8�ٸ�d}35�:�.������S�\q���ׂ"̤e���n6W����'m�7x��G�N��\�:�T6����[�ݶ�9�r}������Ԡk��uf��$W�}���c����N�
��o�_K뛾�-�O�:�EM�0X]����=��Q]<C7;�Ew�=K�ȴ�-z0�
��Y"���2þ�;��R�|�7���X������l��1kQ-����#C�	k��1���@!�a,xȠ���h57��FH�=j!�U�v�{ G���!c���^�޽Du���>f#mɶC<>��uy��M��}g�w3�Nx]��QG�xR����������PA�ߥ��NUK
0�����f�j}t�Xr�l�WB�+-���H��_��۵{ ��������8�^o-�^�V`:U��q�Q
i�;�O��4�!yʆ��O��x�]mB��w���	��s�k)V�
���9S�Aa8��C'LN(D��]�(�k7�K���Ȗ�H�8<�$9��(w��W��=mP=�Õ�f�����0�"XV�=���/��79��F6Fb��ͤ��I�D�����٤�S弝�ǱY��xc'���Vwo���a1*�eI4��_xF-�ƚ�g���V��#&�C�7ǋ�7T�����,�5Me<�(=�G���)r��t~��m��F&u#�b"��eiG^�sΆ�|ox�n�/n��e�[���#��*;�� �lX�[>"���g�2	w㽀���P�xI{�"���ڂbf�\�ic��1�&&�� ����A��XN���[~����>�\�
�v1�nk�}�C�˵�����h�][X�l���P��-A\O|�>���  ��IDATߋ��-�y�]��>���N�'�<�B_��W|��.�m��4�Al��LX�9�:ÿ��5�*sbT3Ͽ� �R�ڄ�^<��[��8uO�)Rw�$E06�㡤h&�����@�����YTU�k�|iN]�u���p_޽[��G�h���A��p�_>�`����%w�f����ɍ�&6�`�����:}Dd�l��e8��.6�i}��>�t�E�f4��J�e��xt8��@�ˎ��H�����ҝp�F�Ө�2-��A�o>�S}����[�Mv'.^����x5�h��bx�ȯ��>K!d6T%�Ha��8U*-<��)sg�)�,:`���Nk�eVVJ�ƃ7Ns҆)^��h/!��[���ܬh aQ��oʷ�|]޼&&
f��b �Ա�C~�Y�zw�|�w��)�|�M����M�[�_~��Ƃ!U��Z��B;�E3�6������F��})����`�vh"}��F�0 �]��e����ʇ��۠9��Fw����m��1�R(S��Y3R����)� ���$��u�x��: �딕\��PSSHdM/*f�5��k���	�ߕ���o	�t'xOɢs��t���Z� MF�u�h�U���Urx;N;��g�;�p>`���N��:^Rk�2���5��о���0\f���D~}=	���Q�)��aZ�e��cK��W������PV/���Ҧ�˚����i�]�KQ>�c�y���	J�WܳO���AJr�"����e��7X]?Ǆ�u"����}��7p��A�f(�,kb=X��7��o#a�<Q��^l7����\ѱvC��SN�-h(]�|��@Ou�g�BQi��5*HA:I���A�����*����8�iZ�S�P�F/�8T�3"p���T6I(ci<�!DD�~j�Ll(@A�߮/�]!��RV�e�?�����y�9�9�z�Ck�ٛ�R���Px���#1X�|8G�q���̑[LR_����v��Ӓ����}r.�c��lJ�e�W�X�$�&�t ���Y(KZ'E����澦fm;*슫Mh fG!��[��� =�d=����N09��r�q؅�8��X�HL��h����}=Mi49�ZW��.�MY.i"�m���i���OA�|r6��1��б.����Ac���=�D;bVY����r��8�@�"��q�>��8���+�@as�R��&���0)t|�k�2��;r�����q�E|�O���32�}�A#��������c��ǂ�� �	Y	��>���o�9&_���f��c#�X��Χ�" ���/�y������U���e�k0�F.��p�h,Ɒ��rR�H�!T��Y`��]�|�YP�����l� J�{͸��R{��f����5d�L~���*úy�(���`�� �#�ZCЍ��C�bd��R9�旆�������O�6Ξ�����y�}��2��!I��O������x�2������<y� �^��u�����?��1=O�.�*�����Y3��Cl�Tx�!�Ɗ�9DY[|v�]{J�ղ��6���K��2��F�X����1���ML0+>��L���:�Y�߽�eN)WǄ0g4l�۵&3�C˅UV�$n��9����Q#�ss@�N�OJ��:8�z�@�|�H���Iٸ��U����eqt	U�=[�l�A¶֍�ccV_�J�<1��1���@�C�����@�#���G�16gC�]�$`��i,lp��&���G'G�W����u-9�Ex�j�q�w��<�C@ WA�:_����K���J_�Z��B��^n��D�(X���
��t���v�Јrv��|Խ�H�h�BX���ͩ�	�g�l�@j�:.HN�E6�VM̀"���M���8,�>I���v�o����J}�x��3B�C�4��e�1����eqt�����Ѧz��~�Kg]��.��Dl�M�]܇���l:�ݟ=�A���r�?0=]'CP� ����I��w�+�m2)��Z���n���.��j8����2St���^\�ģc�����bp�N�S�$��K4d�<��t�{�ntʸ�5��S��j�rֈ9�p�݅~/���LFPɀ��e��
�O�1����ϋf�Em �����c�Oz/�-����ׇ��5/�.G-�r/B�$A�hh^āA�Z�iј(�AP0v
�y�5C��M��`����М YY�	������+Fʷ��jQ3S��=��v�L(�T6�������jϮ>Ns��av▢�t���)����`x�8dH�����==RX"3RfX(;�����������%���:l�b&�>����k��@D���Y���޲��^������ �Qu7�@�(#���=�*��@+���T~����e�(ȏ?�P~�(d󠌕kq����&6��|S�뛬0�8$r����;'��2����������ʅָ��$�oQ��,����n���o���S�S�����o�~��Ͽ�A0)�d�z��p����K���3��u]iK�q�u*�l)�#���$���%��J�kf����`��A��؃�cMF4,`��vأ��W���Z� -V~���[�Ł��HQ�a�hxd�S$${	�Ԅ��z�fDLEIi]��1�&N�����\޷���~�������j:�?�
�d�Υ�"t�B�d���-ܬ��b�7:�σ7HG�3튥�΍�i��i%Ǆ|s쒣:��$���ߧ&��"�-婿xT��1�zz�7J'��}�]�`9_~�6JU��0����~|��82��~��%�n�RY%2l��neI|�^�1pD�H�W���f�JzJ,���i�X�@��h��C63kS6Fq�"<qG�����QLKR�X�a�}{��ɻ�V��}6�Ɖ��2���Q���~-�%��Y�`�*�/�����w	��G�=���_��~�{;��QnS+76�̨��˲�&r$ѓ���� &����={����k�������?_�|���px�},_5A_�s���� *�����AL9WG֞�x�2�՚��`�(�+��O=�5�F�=�tK1���~-O9�ᠱV;@S�隁���J�� Kq��Z�x�u�t���nt.�@8m{��m����Թ��f�����t�6�>)�/��"|{Z\�Z�΋dy¡|��K�U�|��E+�v���#�����Re�hG��jW2+���n���X�婘"����v�Y��d�}ts��U�),r��a��6)F��0��[d?w�F"0h3}�㣰�ƍ�߁b��e-��wDC��N�Eo� �at����x�G���۳�1��<�A��n0EI�%����ܨJ�a�������TR
�;=�1������������[p�[\�\Q����qO��Q�2&dǯ_3�����+���#N��	L���.՘fѰƱ
�x�x�������3��g���ա��_�w���)��u�Ѥ5	ܚS~r��E�|_<nI:����j�'=gU������kv�Ro���&U.s�4��6_���|��=�I;�o*�1r�wÒ�E���/N|�����=�"J�=ଝk�ی�x��JZ��+�%�q�?@?tf��_Ү��H�������z��7�-'|����&A��~��N��x��t���>F�0�@m�@^@�H�ߧ�.�N�)��I��T�-pȓ_u�y17v�����.��(��+}���TP�-н�)F��Ѳ����D�bF��#�[�	-O`�hp�u.����H���xu�_W%�p�f	uu]1�=�H=������ڡ	�##=����Gs6C����\�Rz��!�lD���{��������Cu��g�A�@����������������Ͱ�U�����
��?
�-5��T�APBs@��cڇJU�?�c�z��W�7'�Na����}.@-0��a����Wo5w������BG_�Lf�/E+��;$�u:��
pO�rc�L~^9i��b�����d�w�[j7�2�"�`Fz/і��8���V�E�$����Ie�
�"Fnփ�9�*�؟8h���FV,O2[]7�x��}φ�f�A�v:�1f�U��g����'��l����?��&�*���I�����K�ɥo�0mԯI��&@Y��[�:�,�`㵽�հ��lY�(=V7F�R0�T�:X��K�9UD��X���<��/1Z�w��׻��(WW���� ��l���uJ�&�p*&����o��SJ���gP�y���M�%�h#�c4i����]d�6U,,���F�̾L%�&�̓I��������G ԰ٵ-h��V����@e�_���ypF�Ɂ�vG�1+9����(,��,��V�ml��Y�ڠ�f5'촐8���8����M_,5s�e��ξ'��8��t�2{�Il�G(�o��/�]�U���<D ��>�2�e����v���"4Q��Oe�J#򞹤J*�(��+�����������(<�x��3����.��!�(UY��eb�� 1k�ӏ�Q�$��X�3��b�Yf׼5\T%�-W�����ൟ���S��|���3e,տ�������L]Z�7�?^ ��T�9GlJ�^3ၕ=�������iv�y
�<���,�7i��<f�	������8����?�Yw=�,����?���'���A3��Vc.��Ƥ�N���,��$�S۴���ߕ�U!3 2�㣂ω�2�� G�o�5�73h��|Q:�.���޲�����g��C:��[9u��t(��7���!�l�e]Lu�%u{�Qh�zѽ����DK�W!%xw�<2�'\�y�*&��䲛dwf�>��;mY�a���,�j4]�Ze�C�1���MH��JA��g|�uU�ULg����T#Z��`%������l}!.x*�����U8�v�O�W�c�5�2���A���{�Q�p������UZ3��˔3�[��Lg9��x7��!��|�/j�ӕ�!8= ������N�׭i��s��	��]�&��贸�|B���%��IH�>Q����o�5�_�y���,��Q'>������Od.�E��{�L�]���3]�w�кa��XS��؏9��q�ܐ�I� �ȴ)�a�Tܗc���t.�w�����Pxz��u�'Q��<r� ~��3�"@"P#-G��u������y�Q!�b:׮�>�h2���0˳3K��*`�N~��3"�.z����*ȡ�A0iZ��eb�t_r��t�}v��/ބWՋ�����תV8��'�13M6�J�!lH>d�b�S�@z{'�)����vV�*�6�8������e�.|t�52i�A�'|&@R!xk�2rخ�!���b���7S5�&��8OY�[l;�G���&'�o�ZXE7��	{̒匀���!���K����]�Vλzp�q[m��B<ڬ����{v�\�vP [��gC��&�ux�bĦ>:���F����<�]��~s@+�4��b��f�-�I�k�nS�V����zp-ހ���%n@4$`�L!�ҏb$s-�!�J�A�/fE����|��ӹ����8�y�U����+� ?��j�KMe�W_}2���_ߖߐe|���UF
u�)4,��)Q�2E/r߼�T�{	i�NA4�-{z��e
<D�>�ʌ� ;�ef)֓�o;ZHk�d���!����©��fFhT8���GRW"�R����*Kr�o��!a�\U��pƋ�xY�c���N�K��X"�7yn��g��������}r#-��=�#�<��~��DZ�|+��0n<gFJ��}�}��(���>�8���p�o�鞥tU�EcEp�Z�u*�P{M�H�a!��vD�f�
��A��R!�0��F�$	��s]��a�����"�u	
��c��2΃���i��.I��P3R_/�C"��2���k��u5#M�o]R�q�,���q�T����k�/���=��]TF7�������P<���Z%��fPf�Y)'�]�b�uF��.w��?��å�񔾙�������vgr�@�Es��kk�Ic��[�|S.%���A]ʁ�͚�b����A%�&�.Ơ�ס6�V�������BlZ]��5S��\Ӄ�&q�����t��2�<�m)����Ta�uM�{hJ�I�4����w[��ߣR��w��ML��V�C���l��
� �'|��.�)g�p�>o�Dٍy�C����Ϙ���]��N����D?׃DU|p�%h]S��9�J����m�Z!;�����0u���C��&�t����^L�MբU��Y1{�m�Fs)3�&1�����MMj09� �A�WRЭ���������������E�	3tM�6���&K��֪M�S�6 ^`�Pk�ZkH3F|:����NB�=�X����r�%�L���tJ�F�I��.:��^~�}O����ғ���<>1t��X���g��V����э���ލ�!3/� ��_��KhzFp���� E�l��
.�F)�M�!Sk��`�N�.�@o��ٞ��N�#��������|9ZW�^�!�좊 K�W�x�_����7+��ch��S�@PQ�W[r����Tn�o�ci�W��JI+�暁��������������fv���m\�B�����<���
MC\̛�y��ġx�ֳ��2R�j���G�H���Uф�؀ԙFVgv��Z�f�a'����@/˚��e�ChLM]K�I�a�ks�CY���{����*�޲Wu�c-���8#D����r�贜�d�}~����I�3JR�� VS-u��=j��wc�H���R� ��Y�3,ӝ�c��~���MO77�?ٵwF�6�yZj���f���dB������#>���tb���)f����H���^�u(h�$14�6A>��Ѯ�C��P 1=bn4	gQI�����L���,�u��)@�Q>'Ή�� �E������l݂(g��S*�t�pW�iM�q��'�N�>�)��y�� ;mj{��U��t��z{
y�I�0� �o��m�F,39�tl<��
L0Q��v${����V�8Ȱ	���?��`�i������E{�������[f�h�Dvs])��G�ܜU��b��Kn�_�ɦDS�l�M�˷i�Rg�:���G� %�@�������97iCs�n���V�{gIʍ�y��6��w��3e��������ֺ�a�a���l3���`�6�A�4�e[0��q[���=xP8s���1ى5E��Ks7�}��C�oi�����kVc��t���C���'0��
�����1����E�DJ�˙S�,F���hz�؟���*�c�*�����k�굃f��R?�ʬ�i?�G��!kC�r�[唝�x-�K��X�X����Mau~�vp�ݕ��d�F��*�)�L<�+�=7���dx�#SZՀh�+�1L|�b�p����
Ii��j\y���kg��O��%��i!�\ ����r{�!��Pjڂ�*��9cbE�r�*�D�$�?�! ���q���۸V]��\n��L�����!�o�A#�0���^�0p�C���Wu����]���e|���x�".���gE���`P��Y��Vxj�tͿ�}��V?�{b��ա��7|��*j�<�6�
!����A
{n��y�����0q���J��u����3��s�k�\Q�`L0�"^�)Z�������sm����Xէ1�4TR�.��Zi���L?���i����PoN���(Z{�� S.�H�9g{�����i�����D��H ������xg橖Ķ��u	G��\����g9�ҝ�,Xl�~�rŠ���ͭa��=H�}���w�Y��~4��l��ն��L��T������V�)��h(��-��>�o+�`���i~�L�#��-ʀ���4�1���}nw_���wAm��A��:p����n��]���A_��:p�z��O����F�J�R�M[@C���g/��B�{n����v_
I�iӬ�c��n�)��h�t]�+߷�0�Ȑ'Nt�Χ�����	f�n�z��yx��@@/�Q�Nj�q�l��	j��^9c�������1GF3�j�	+X�����a���'n����^������aIf������g�6h�����9D�K�G6�յw5�I����,Q`�� <Ѐ�;�"ڷHR�g��^f��Uz�X��$ᮚ���i6��4�E�ާG>)�JF�Z���3U!f��a�}H�(H{�o]~�L�פ���z�8b��g�2���Y|u�9|�����M��/�?K�#�f���.K�LC(8������n�2VdG��F3I��R��s=_��d��l+�pp�zHy�c���cmW v�6���Ǹ쭭��o~tȯ8���� 2��B�����W*�8����꓂i��M�����һ���y'���(����fP(�Ϲ�.��5�5)�`�+]i� ��(d��S����lG(�X��@R���!��`-p)�a@�u
LT^�2O|��-D>|�n@�����jaq�kL���M�q�؛�m�Y#"�B-^����*�A���3h��-ᛑO���҄%���I�z8���vQl�ئG�92�
��ì��6������B�Qe(�_�;�V�yټ���pz���c�k��mk��&�Y�O�$���N�b�|DT��1�Ҝpܨ�������0|Ռ��J-(������p(�P	"36�s��et/A�#ձ|���0�>R�σ����97�²�Tq��L�����|���BJ.��f_�npK����g�^L�Ш1p��1��}Lė����Xٸ�c#/�U?�|/�f���:�P�<�!=�&2��xy:(v��o��t!��	�H�49��2��Ha��`j�2�9C���1�:�l��W��l�:�4'�D�������ܘ�����}H3���׌vO��b�G
�m�7&�0�QH�7��k�{iZNp���v>||�������(�L
�#t	���>���l����䁖̎�T��M��������\�a�1W|2i]gañDs��׽h��@�L������<�+�sV�7��x�!~�.cm<6��,�g�_��/����w�r�ػ�N�{ǽ�[Cym����z>m09�V����9~�_X�(��B����Wp��U$�/��� -���L,�=��Y����dB��d7A>�0��Axd]�������)��"��Cܽ_rʄ��w��:���#n4��a�g�!�{�A�3�h�Z���ʴ��{и梲�*{��n��D����{����ՃG�6>Eh�.S.J��c��5]A�&�z{�BW�(�~�_�iXO:��6�	��
�0[wӍ��Ͽ�"����B����M9e��k��繍�a����hfK�	g���>��r+���O� ��ǿ�sBx����S�Lk���n*x?(m����j>���d���U0��)x���Z7x��={�k��J\��V�xh_3�&��v�%������΁����x[�Յ��gۺ{�g�hL{��`u.���2Y+4����K�6���gńɏu/'5RM����լ� ZᲊI?���T�#�S���v�Zb�ɯ����zj��TK��8��Lc�8����9�*GO-E"�z/Z�GC�;��iY��"L�v4P{�iE	�./\�z_,ú�f�I�u�q-<7\'ZtE����28�.C�"f;���£2<�r\s����״R\���������#��h��Zet`I9�%6�����M�𓺉��Y.�4��4j�������%1B���� �G �b�8$�NI���޲��q�B���̝Lf��)N��C����z�n�UNj����(?��}������T*���FMhb<�M�譆J���|>����bB<
C4�t�Ӵ�:a.�~����V�@$\�,Ns����m��9��,�Ln��� �aai��6;Y�������j�u��	�tf/�k�,CMgM=�S�Q�=��"iXm\����:�U�w�R�M�t�Ƅ&�����2�ܶbz�S8$2RߌR��ی�6j�A3�p�xý"P�����.EL�
�G��V�h`���-�H�iF�WzX�Y� �6��^`u�����Z�)��2���A�62��_5Ia��4��^o���R�EYKSI���*c����M�=�0��< ��N�ҟ�.��&`�:MiA C�̍H�W��j堹y����D�얷�5�8�V-�潺���:��a������ut3�����c����c��pR�!����AU@,ϼ�!��6+N(��*U��_����>�ry��}f�2)]�=!�Mﮕ���Y|�`7�Y��9����Km�������:�7WwQS��X��vи�a��{$(�!��� Ty�c��&��_����/Q���HM�*����i���X�d�ܗW�(Cn�!�8�g�����}�,�]�z����2��I���nbܴ4i�o��z�8J�g�G�b����N��vX��4���b��O��C��]b!��FF�����]r$ɑ��{\���
�*���r8�v�����2�yCv7�PH��׺���Y$��9˙藝( 3w35UQQ,�����'~�<O*��S��M�t����͂w���e�m6�f%�O7>D��C�n"X���]���A�n�"3����Ŕ�a���`zʃ��Ʀsu�f�e6vai�ꀳ�̠ź(�3E���
�~
��q;Am�N�,�Հ��L<:�;+��%]ދ��Nl
n���0�,��A\\i��Y&[�SE��Y�b�{Bɿc�#� ~�� ~��r���VT�䍦�y�kŜ�W��j��}�6)M��>&�b��SVU��J�D�\���3k� +w�#�6��k>H����o�0m2/u��QY�-Y"�X���s� `�_�52�A=_�\S��U�c�]]Kg�5ȭY���k;��og�WB?�Ȭzƾt_d�W���&�V*J=S;�4̉
c�����?���v���{�;�Z��(�����Y���T�oN[�,�y��f*O�B�P�Q������C^`(]�OY>pE�`���"��f഍�e�O�"^+�{��H����u�}��hDl4����m�4�_�>U�v��j
Ȑ��	#����;�QH�8�ח)qY��@���.�1
����s
{N��B����r˚��O���/?�İ���Ҳ#�Q�_.T���/=���sP]�}���I�R�t1�d�FgA�V�/w�3PF�r3�Р4��cv���or��,
{�}&� �3u�oDo���Vl%s�f�����,�C��Uԉ��=~��М�*�\�&����f++E#t7d`��$Q;<��͑HL����5*��'~�g�=�'|�/�,K1SХ�ȴ��s�@�ڬv�s̸fk!>^~�x��<SjJ�a�ԝ�	���$�1��R�E����w9v�Pw�X��>;�(H��3�>�N/�R9����|����+�����P��"���!�~���O*�2�E�F��Y�k,�}t�Dit7K dR������m����������0dَ/�8o�������L�N��YE�����	k`40�Y@�! �|/���b�l��'L���s��1��b8`�O$��0GkX��S�o���.�k��ʪS.�C�%V�Y����I�D�� ��̟�����qA���Nѥ�쿼إR�5���$�F�g�T��u�e��T3�P:݈W��۷�۷�Rl��͏�|.4Q� ����$�e-��sc�ڤ�5��斮�s��YT?T�J�=}�Y�1+M4�N��**X�K�#��rۓ�3�|��*���`��yގ��;�O1k��]��!T]^�g�C�\]�(�׉�vo����}�N��:+N��R�tͰvW2�n��=�X�]���@%�Hkc�f�yRu�y�L4:��;�u*��~�'�Z|S���0<��ɦF�U8���jH�{��&q`x�2՟�pqȖ�0�-�o����Ϳp�/뒥I��5�T�̣J���q��@a����W6�~��G,_R��a�#(�W�s�Q���n|�7�ƅ;%�0T� ;?�y��rsL��Ԍ��Κ�����c�ۂ%����_�o⯃W�����5���Ҵ,F�1��`zX�54���֭*�p��������mU���`�8L�y�-��z��!���d���c� %�[��G���@~Q��|n��L��P���ݧ�xm�|�� {Kv�`\�M0p�h�In�U� 5L�=�q6	�t�2t�Н��m�4���15�x���2�U�3��8G&���wXJ]��w�y*�u����̤Bj�s�w+���Z��\·���`��FC�"9ʰc2�����uu|ׁ��P'��0�z�������{��9���<�*�%�g���É�����h.�$�@�i[�b�? EɄ`�E�@�����LQ�+}ɊO�QV�uqs/դ�ۮ�*�*9=K�R��r�$���*~�L�����������	&�d�%7E8b2���z�εs�1�9J�q��{J�q�;�u�$ h૯^�Nde(��x�S�FՇh@���� ��J0��ǁ�<ӲbV%�0�m�m�����kq�]UWJ{�NՃp�"����Q��#��y�0*���B�'뚕��Hp]�������m8��C|u���c�����^Q�����nQ��z�4�@�m3��Sgy�
�;��D9�a�ґz�DV�&���5&q_�;��-;�Tq�R���b��e�.���Jdanژ��L����ו���}����B��������*�KŴ�k�&c��q	��+U4�Ү�U��e�`�y����6���&����6S�oÅ[p�\f�͡��J
��a��hfou�1.�S3�.\P-��5�L�F�Qj�^��app�4P�q�e�#X(�f%L�x���a��L�P�V�u'p]k�~���i�0��[|]lB�~��w�сq����+ΰ�X)�pS������m��S{�
�����d��SO���E��O��9m��Y�������llt��Gܘ�-c�l$�1��<f�!:܋c꾣=��>߅�SnԶ	Q�+aY�Xb�ŕ�>G%�r����
JP?|�gգf��َ�I�u��v��[0�9�sz��p��(VUs�&pe@OB���,at���v)�d��ş[EGwMA8��ȴtؾ̃p���-Ȇ�-����)�°�M�C|g�`HZad�K���d�Jr�m�U ��h_�@6��Ftݷ�E����8�:##��	�̮�nD��U1L��ؕ$hr	��
i����'=�px������C��:�-ʄ�����3N�=�l����Aj�i��ZXHk��C���RͯL��&�s��Z^	S���0�o���J�o߽Uix���s�6,�i&x_]}��>3R��)�Zx���*#�Fj6�i���:4m{ܷ߼�'�?��?��a����'��'~��oۦ��ӧ '�$��=�ŀ�fVt5�i�`�2�e���w��wߕ������g�Pa����Z��c{e!|�?[���EKY�0_���%!0&�L���e���4�+<�|�8Z�"6���5�WF���)�ߐ�撟K���a���/����q���P��}Í}G;�;��]�>��6t��h-�@������|���1�k�i���챌ƩrY���}�����sY�w1��EsP�i)�?ex�A ��vH ��sb��H#˴r?^��̽hyd�\�rB����8�����9Y��ڜHE�=k)Ⱥ����r_�>�_M =�w*��^^��mP����U�?3ԦW�9�Oo��D1���R��_��?��*�*��W�hf�����|�8E�f<��S��%*��S �{	n�4 �������F m�����~@߼�E���U����"H�b$?2�͍��NT���6�\E�l�yьS���}TS���q���9�6o��9�8�0�1�S�p$��0�υ�:�8�lI��;b�k6"����}X"k0�V�����f��{&�a/�k\}����9-*w���
9��$\��Z	�s���2Mi����˟C��/巏����K�n?���G�����F�g��4��{ҾUT��\�`���~�¸��
�Y,XYe�Y������R;��X��C~�&

 �@��@�osp�mRfI�]M��Z�\�UW&�k��TkҬ���^9��l��4��_�=��gi�Ms(#D��d#0����Y�-�ݯi�`rc�����1CĮV��=�������2{�f���Y<���%6X	\�	��a��Z���.��w��w�����ђ�
�<KL���Ҝ|���u�V������XJdbKr��3}u�4^d~�	� �+k��G%CNu�Bxn�)�#H�<�d3Ɂ��#�J���8g��x��/5oN9��6'y��$�e���va�w�9�]s��<$���Ķ���H��P��>�	¤�r�����B���m.&ܗ��M<��|���M����Q	�P�z:�Z������� �Q�=6����MnX]���Qy/L�\Jd�yH�5Ƌ��E3c1���6���p�>�A��b`/p�>)��A�+?��.���\<�7�2ј�{�?Z�8A��p����e�{z���Q�2x���,TYf���)�)�e�
9�D��4<@���`��	�f�H�WZ��j���J�1�����A���Q4���j�ղ�^ex����d)�_Χ[�ߗ��ɬXG��U�1�}�@�`�}}�&��S�|�gO�ipg�-@���@�N�������Z�a��n��>V��x�<[�,(
}��5�s��/WV~��1;;�ݠAYL��(�)�1�hc}�N�m��,c�ͥ���I�d�k��bmH�}�A��ӻ*9�Ċ�Nu�_�2�\=(ܙB2{)ҟ�{b�6ⳌX�3�'����w�6ǭ��?���CI~�j\X��iPcm��x���5@P{����iul?Tzת9n0�m��?���y�]엟%N�)�7��(�RW�&���|��4�&���a���e�� x3��~��Z8.2h�]��]�aߗ���4���F�~	��1�o6B�	���<�1�UJT|9���s�.4V[�ԣ�]TE6��A�n?�,��:�0c�؃l��(����.�;/�AaӏݣDZµ��}�u "|3� �B9lB�=�����H�Q��V�����u��s�U����u(�A�jzw}���������jdm��2˒A��h�Ԍ��{���-rRG�E]ES8���:����a�(e)�N��P<�CԀYD�y\%&��/Vy�ȈQ>,d82�[�%�1�fN9;�@z8�W'����3j��l}�y.�Jji��4���u[�R�77G�kjA���k.���&*w�Dtl����&�w��x�,�����#P��P���H�Rq�Qdof��<1��uf��6�yd�B��m���b�	ҰV�(��˿������|��Q8�OY���`ĳ�w�BAp���D��9IRmb@||T3����]p��bM���4y��I��a ����)�a��ӓ �K4Q��/��n� =Ji��1���o�^���{|ޢ�D��tp�j��ʹ�E=���\�j:o����jU2��.�;5&�]�xo�'�U^�j�-M���F0�
Xe�N���u��nV����jE��$��H�_��.�#⿯����U��73R<O�����:�F��'�`	>}��rIc��]���B�������٥�5�>sT-d`�
l����y�{j��.aUw1&J<��F��Y�d�}\��,!8�M Sm���k��g~����x}�JB\�;�qL_�����Z����2%�'	b�	�&�*M�\��rtq�in*�%\�X���J�Q�\aB_�5�ΕɲY+,7����ǘdy|�ͿN�Z(YZ��Izۯ��/��*��/�J�;1<�>�a;��������m���샎�GeM^mMO�!�y�
6y�lҎ��Zƃ�b[���p ��ݻ�Y?�&��l8�;۫!���5�A����_�� DV��tf��|W��]��ޮ��/c��"�d_��͒{{MU`%'���ǡV��4s"g�]ҏ���ág���2���R��՞�[EU���kl���m�3M��|i~�k��RI�J	�xOIHD�Z7x��$���~}tW~V��7�8�^�^����&�6���a!�>�t*����i#��S��b��O4�7KS�� eQW�!S���������_���Ngv�倫�[#�`�h��o��J��S�$l�_�p���n0�c�0�S.QYV�� b�n(3�([Ks��1���86�m-���%���LY��ڔ��΃��D�eXɠ[�-��=�g& & �h#���NZ.�1Qt���ŽBP���L�������O���筤W#�xv�A�T���f���(zJz��S4w�@ uy�������b~'���S���n=p�A����*2��ۗ$���p��ÇP�*ѐ���N��H�@:���D}e����/�<�*�U�n��֜l5tG]�]'�>�T��EE ��C�Oc��ޑy.���$~��@��Z��@_�ރۛ�7K��6��X*q��	��x����g؍�y��49�Lׁ�ҴL��1PW����9Ú�C��^��
��t���8S�xq�5�e��B�k���kDF�i�{�O<Vb��ɵ{�R�H��K��ݐ�G�(��;̉��Ϯ�'p��X�w�Vz�馌iS�.3R�[<��m�
��gn&�~A����>tQ)N����@>G�9)2�������J{lLa|�E��zJ�C6[dC0I�%Iٚ]�Ӂ�V���<;�ȄrI(��k�*.YV�w<G��ؠ,�3#�F�������?�ݲ���.��4���-(���	-�'f��Z���@��O�JWz�V$����\�F6,��)�.��n'��DPΩ{������'�������}���t�H(4f�܋��i2���@!��*2WR�愸���a��jR:������xb�lF/���T��r��S�5FUoȍE/����.�!?dS�t5����eL�n�}�����������Yk-�?�p
ރ�JV����/�w�ޅt�%t[�!�T���Ͳ\�	���(����/��x��@<�0Q��:�^C,�P�c�-FZ�JPg�Y�!3X�+?v�W�/ty��	=��N!�[�u��͇]t������"5!N@]�]]� ���cF��w�������e]�kԲv��g =�n1қ[b��%��\F�'F 5V�C����9bxP	C��̓��%n��5`|#�=!{
1pY���Kg�5��]����W��n�ajT]�ՙt�������X���Ǟ��B��[&UL�E��,w����?3�y�f��ھ�u�㩻�i���n�}����9�<�Yb ��8p��2(~�	zM��Z
�Ja���
���:��\�g�X~���b��_}���^�Za@�\���7~G�����9��б�Mk��z��*q��ԇ��Jި)���Ͻ׉mOUp���\b������S�-TF�['�RMB����̨�\;�����R��?�q�ӆ��2/�0`�s3Q�����d3��PKƷ�;q�M4�Wz�]�S��d�5t�򺏓G�Y�׾U�7�~��I:���%)No͕+�00WˠSS	���s����áR���w�@�a�s�{�9��L��xt����#���tִU�y�Q4���K���$��R5��8� �SO�Y�SB��ϸ��:B��*�/����2W�-;��jW�,���l\K9�>0��xX�/��*�Hl�����<=^¡u_.5(v���m:�M:���AX��HC���o>�&���0Bl���O%6'���!D �P|�Fm�L��9����>��W�_�y���E���.ɷ��=ƙ�
h�"HB�?�^����M�k��$�� ԇ-�Z��Kt�`2�9�6q(�}�<�x�N���m�a������E����1H�?���T�|W&Kp6�>esNr�C��FJ٢&�����1�l�Dy}a��\p�����>�v�6̂�_��l�?��W�P3S�t��-�Pi������H���*.fRy���i۶_k�i]�Id��>|�'o���|߇c���.���]}�N�o�4;�$�K�\���d)Ԍ��	���5h���1�Z��8�iU��K,��m���,>�5s-F�Z�a�ټx!�%9k�q�]�=9�0��,X;�$��EF��/1��;�����-K`T(	{�AW��)f��k���� !?��^Kf>Ź��S�T҃��)@%j<�$9w��,�b4"�s��lΡ�������w���0��?�(���=+�q���Fe�1w��W[���¸��ޱ����*�:q��G:ǄW�Ȃ9c�˯œm�,�gN�!�d8ĸ��M~:�����v���'ѷ[PG@���
�{f�m �J�!���)��\�8�8D<�[{�k�˩�= p�z�6����@�πr^J��b?_����Ͳ�.�(N�H����y^��IH�c�N���K������%�a��=��	ASN< �>gbe������Á���ki� CPL�����gZ��u���gy�#]�����ȃ�g����eW�AjF�{�h�W7��C*�*�&�K6�y�E[R'ؙ�1�|�t�7��s��'���F����%ʺ��|�^������6>F/�m���{�������#mT��)F�uʌT*T���矸�+޾�}�n���Y08N	vBW����X��V͌��y���`N�))��-�9��߅t������� ��Q�q�`�̔���A/�y=q�p�_o䙆u���!�A
�9��*��#�)k}�w�3 �H͜�)��Y���w��kS��1?�d��8[[���8��Dy��W�_DP�WE0F�����Ge�����/&�N�����&O��������`��+
��:�f�Z8ݨ���b��D���d���S���^�$���4S_�yw��������,�b��)�Y�x~J>�W�a��	��'�I�H\p���)L��Q��9�x�~)V���� �-۟$t� �tb������Z��`��XӿJ���'���Qz!�*8mV�S*NOy������I�T�A���a�b����Ooys넻�}�l�"7��%���[##n�Ag�&�㔂d�g�=����H�7A�3w��ж8��NK�mG�
��%���ڞ_�"ޏj��ı'�5���nn3@Æb]�A��P��خB*���S?����k�Y��C���Þ�8��yW�/5#+a�{�����u*;�UP�J%��>����?�#34�~�����&�?�;��9�h�⿱�����IQ��DQm�Ϝ����۷Qb�x��i�}6x��y�ÎU��~N&�����x�߽{�l��\4�°�Cs���'Zd�3��ɦp�<�Εn���
�2=ixq `��ݮ'��J+x:H�����l&��qU�e�Y��@������hX%�������r�=���,LL\w��l�Y��n���Y�h]���X�vϐ��]��넱��[���σl�+<R�,��b�����'�ˋ�S-cfj.c�-!�'E��OUO'����>;i��N8'��A����HE%Ѣ��s�3���;�v���ob�ׄ+�g��B��'�;e��&ӳ�c��v,�n����=3ҋ|���|XGKX���Jɛp{����^7������C�t^�zC)_t7�U�;$&���gO��i�5�)�$O����#��,3l�GG��`������(�Ⱦ��8(��Ǉ;� �Y����]��"����/�=܏{�b�Ǹ磈��~��������-֬��oY�#CE 7����P=�(�5���.e��bM�bX\c��$���C̦+ F������ .!kc���5Ք�>���ܥ���u���A�����!�c�<º�r���gT�Դ=Z;c��k��]4��;Y�L�H���!��Ӱ��Cb�OOUO����~ga��A?��qSȰ�n�ȫ�+�H���c��j��6����M����vב�Y���fSl)��+G�h6��d�%��&���꺨�y�Jv)%ʩ.|i�7@ٸwv�������� {|��
�9M���;[�bX�m�{�u4�v�	��D�g�wp�MG�_���k|��?��?�	<�\;d��L�,�xf�C��iqSOAZn2Rw~�gzN�MQ��AT"f����n��X-0�x8��l��f��h�Ǜ<�k�?�u=�۱����_P�z,�Gr�m��.Kt��u
�\�2���`J�Z���]���ZwP2n�.88~��G�z�l=+�o�޲�o���=�3d�*E������?F(�fd��k�A��3����U��?��O���%5ǁ�E��z�e�G2�ސ�"��'�<]�L0#��L�%��Ԃ.�\3R�.��--ŵP��\��:�}�@���cc�h0���>ǐ����P��-��㣦��]϶�ց�dÅM��;n�K�.'��:��wŕ�S,%�t�m��U�q*���E0~jL��s[�����������oF�����H� Z�e���9�~A�j:�J}�RԦ����xB�"�SӐm�FbN���58eh+�ݒ7�?�M�<��Ǭ~���^R��(�J8R����g���#m����62 ��92x6G��TƂD��ݜv�����7��y�&�����~6/@Cn�`q�~%�K�Ҽnk��*�i'��@�Q:,�� Z
7�n; �}�K*�)�51�L��#���g5
Un.*�)���t���q��n���?x"e�qQu�q|���:��`4���|U���P�#�}�M,6*Hњ��!&��y/�F�m�O$:��\�:�7���8����ϗ'fy�`��������Exء����c�&����4�LO�\4��߅��3E���6j�c��6Dڧ��8JZ�wY��K\23�H2,{�5�Xdw�ߗ��������DNK���]�o7����������.&��p���R!:��+Ҷ�h�t���:���!���
���䥝�kjۻh1�/2�6�u�[�c�䳙Zp�T���>�Uc�ւ�Ԉy�%�<4�}v�G��RC��h\~��>2��cz�.x��Ң����R�Bɰ"�����c{ &��\R��e���Y&�V�����X��\� �2��ڜ�d���������Y�����_KS'{f�/ev��@�_HN�$��eu3N�1�nw�a���.lc�q�񿔌+O�5u�Р��w���_��9BX��y��gW���Zb).�/;`�><q>����������7�8d�@½�Ͱ����o޲�|p��\��JM�c4"���-��@������A�+Q��X�Ct{�l�\_H���<Q��ٵ��!E{%��9��5�Ws4�P��=�����0N��l%�w� ��b���V�/圛}Y+��,O���4ɇ���	G$)L$�J����3nՅ��\�� ���1q�qʽZ�1j %�wx��X�Ɗ��&�@&̋b�V�r����m ��d)��P�U(��tK��u ��~�]2\��iҸ��������	��i�_�-�k�{�0w���@�2b��齻�%�p4Z���!�Cl�9&5��1g�����RK4y�UӴ�g^���.�-��p���kf@����s#�A'
Eh���m,k
���tj��*o#�����O�>0K�H$6:�&ў �:mL�d��K�m�S���z
���k�`Gn�������;3�Ȇ.Y?{%t}�h��bi	�텙�2сYX��i��r��F�����Y^1��k��w��A��L�������4�/�����
m>�4��Y�;�����m=>U���&�����̵`��=f�_���l"��E5���R�������o����r۱���dY̡��� >� �� ��wwK��?�q �ґ������'��Y])Y�e�bZ�9����A��:���,S[f�z�XlȢ!��zU���z ��)x0���j���{ux0�K�=�RO$�C��vekTF�0O�>n�{"�{��.�_�?�8�hZ3R_/<���646�p�3�ps1��Tlb�����D��4�Y\_m=x*��ҴC�!�7���T���,Qm������<� ����|�L���c�`K%��O�����P7G97�"C	��~����?���/Rf������1�����=���?�q"̘�/^�����_�;�5Gb��0�U�x�Y���X�Os����:N�S4�� ��`w.e���J�!�0�`_(�EFP��J�� K�)޲�`�A��.W�E�5�?7��yAWU�n�5� p�!+7fV������ՐqUÌ��Fx������(P<]���U��`���H7�ͮLHB� �����/Yv�ٲcg�]c�fXf	�^qܻ[6��UG`W���j�Ah��I���^1��ɧiv�X���S�3\-٪��F���Y��Lr��\����C^/Q�
��g�^4�A.5���U�����`�k��Ʃ��W��j,�7U˕t�4�0ph�w�l��re,�v���>W�������]��R$����HG�bA��X"�X w�ҥ��q�� *�@�f��wƁ�T���I����0'��[yG��z�@�3�ee#��:�7��<���>>�JP���ŮK��NڟbZ��vM����[��k�ܮ�;�jb]`�A}��"���6��湌��p�KN�`����w�H�>0��j��1,��#���FԐ�/]bU��BUΣ����~_e�8	�=R<B�ͷ�M��1&*amb�8�&�7c�i��T�����HqN��[9xn�83�\{?;Xj�W/�O�>l��m��5�N�3�]�Q��r$U�1��O�������9L�.���\���J����\��D�j�!e�'M�ʹ�"���kjةkbI�E��)��9�6Y�Z���k! ����N��*>����]Q�i�I�����I��J�(t�.�{��Hi�a����n�������Z����k�Ef�,V�U�&��ϐ2�h�Q5�Z�e�v� +XI���/XG��<�;��Nx������C�� -$��B����'
�;<I�'�ҽ"Fy�g�� 
�lvU4-����ޅ�L�����:_�$�&�k<!Ȗ5G
�ѺyDrs�����[H[Qi2&"�8p=�Z\1!��K��������%^<�b*
�q3���ʄܙ�
@C�pBuH����&iDM�A�D��I��>~T�&�9��V��Ÿ�SQR�B�ㆠ6A�h�����a�� \s�r�MC�mБ��0`
x훯ި���60�C� ��?Q��#e��g2L4�Zb$Yx�'�&���et7����#��jm�Z�G�O�'�N1z#�l0"ၘ�K����O���KZgҶ���goz��l�s�g��s-��5���$�75�w�>� M.���� �am ����NA<-�Ԩ�Z��zb���.E[�������Wx�|ք��
Ho����[v1�q��gbq�ͱA4�x6����Z�4�Zn8��(�MĽ,MW�^'砣lr`#���s�x�����d��j.�x���:�D�b~:������e�@�Ȏ�[��̆��.��7 X�r�7��Q
H(���Ԍ��@
���Nie=�Hi��W3�+��xщ]�:���Y�aWr�3#-�tX��kjQ
��'�aps�s&��[��>^h�@\K�["p��BF��O<^�Щ��mc���4n�>gR��yQ�!&\�����GF���ÿQd�f�����o�|�ꛯx ��NC
2��X3�Q!T��<��*��}IȬ��<*Hh,��a�Z�k�(�Y������G6������2���w�����U�{%8}��q臄�j��N6՞��$��25Mr�AW��LנT��ǫ:�u �D5�����J_�FH_z��H�>[}�}�&ED��R�?�W#�k��Ԗg�̤68�����g���د�H�PEa{u��>Lhr@�6��c]��щ�,6�Z��I�8le���54���|B� z���9T��A~R�u��^�(�ڟ�aQދ%YW"�U���x<���e6w[��+?�224[���n+���x޲���Y��Gt�?*���u�'��q����ڂ���}��Y�y�x�%b��>�9�	xs���p�Qa����l|,�-X|���m���N��Z*��香�l��y����׻��vd铦�X�`�gV���q�Yr|֧U�K�iɔ`��tʵb�̤��~u��Rkfd��(��N���i��_�T�?o�q�NA	Z��#�ȶ��s��a���@,��_ʿ��^�y\�-c���^�ం��=�C>n7��%��!,u��ތ�*��Wt¬)���uS��Z#!����9q�I�����:e��pMq��u��[�"�B�0�P4�;P�!���!ǟ#�;Ӝ�w��X<���Ont������.��%2Y\O�������TT	�l�y?;�/�~<vy-9p��k��p���9�]}���2�8K�A��&�H|��K׽�u +�Ⱦ$6c@Z�ɒ����5,�w#�S47��n6q��H�6N�%AzƖe=n�g�$����h��dC�~x��m�R���!N���
�w[ ݽ߂aP�>�߅���)O���)����N��T���qVQ@@�������[����ɱ��R|]`��H&���ö ���X��N��@=
l.YU]9r�Z��-�Dp�t'��8)㇀���P��-uՔ���/&��a�;pS��&�d�|�C�vp� ��᧟���K�j�ڞP˸����3_	�t%Љ�5�o	���a�fo�z������	���D0�t��q,�?=�~�5iEaC
����_�l����^�|�d>}*�sj��YSm��m��2N|�*đs����e�U��C��q]BT��}B<H��k�L���2�9yv����g����qv>�<������z�!yp�����1A�Oqv��~_��T�':�GOAI���@���X�
`/(�C܈Xꨯ94t����D�2ϳҒ�+���6��	lȿt��(U��`o��>�x���R���|>޶�s���q�⍭w8�p�/,��M��H_�E� x@���k��X���-|���cQ�̞i��ʹ�`NEm�D���R��;D���莛ma@_˧�ч��,)�)��j0������Rw+A�Ң���j����(N�������������w����#x��?�5���m���I?m��@�2O5<+�u��C�XJtL5^jq�\;fp>؞�i�í#���Dռ�$�(�T8ѵ���ϳ����&׶���	��W�x�2���,����4#M7���Tl^��Rv�ʙ-��]\[T(�@z)�����0���H1�
�j���!�MŒ�#;vT�u�H�x�+�e� ��5�L��v?\g$��ll�|��DxP��2� l����C֟����2�SfMID���Su7�p�M//���"���ce��EC�ң,e c<���7������E��]c�S��p8x�	�YO�]�$�9�:Zw��tO�ߠ������J����E��9s�e��I��|L[�uI.�50�n҉6ש�>h� *Kx�H[��Bn���:6X�
57~f��[�!���	7��K���%�޿���C��1�b؇��:�L��E2��(B�3�H�er&[���TT�?`Jf*���G/ �k.��Os�ۦ�~G�Ydu)܏����ۭD<޲��������_��� �F��$ħ���I0���&�>@��9�DֺӔӶ���'fF�(�2�ǘ�Z��|<�����Ĝ�x� d�qؾ�ɒ�Ko\�����G@����>o��->Rĺ� Zm�H;�ñ&X��9�!F��ȂD��/<��[��  ��� +͇�3�]���0F�"������ן�����՛a������EԵ]^��cW>�W�ŋ�+y�77/#�^�<L�h%��2.�΂L*�х���@d��5a��x���X9=���ӂB��2���-@Mg���%)�!& z�|�f�nL���P�,�>��wC	ח�_$8�#�}xM~�3�f�@!�ZE:�%� ]V/�<�O�z�UXm���sZH��v�lܐ Y�1XSs�>�fB`� � M����"�n��M�h��t�b�5�c]3�ﭚ	?�	���_�s"(Y�v�:9e��dv�"|s�Xoד�>���@�ɩ)Z�xm0��(��Ϟb¢���=) "{?���D��b��r�t�N�gf9�4�1=�lE���E�݊�;m�i
+� NC�n?�D�?�4�p/����t^F~NO�A�L��������`zn��(+�~��M����&&��x�ߧC'�9����隳d�.O�,	]�"@ޜ���&�w�}���l�� ��=�$ӷd�C�uRݿgsO��S>�br�I�ٴ���+���N0�c�Y7�| �2s�z���%J�h<�5��bt�5V,x$�/�c��3CU�t_3�uۙ��B��9��f���5:��t�aT���KmƐ�+]�ur��W���{9̊t��nS�H��r��Օ+=�K�#�p�������?�����?���h��
d?��83=i��#8�{77����5���B=���f�r��r�֘XZ��AX�^-MѬ)���2i�(բH!�TXSu.��Z�!:�5SO�FN��Cp���d2�W��]J�����æ��EM����$'HdH���>PY�$�gP���\������(�U8��E#O��
R��6�E�q:\"��R�B��0��-4Q�cO* MXg�e��qrR��s�g�f���\�jaоo�:ݔr�M�.��d�FE��9�q	,� N��/؁G#�7_�w�9~4���Θ<�M29<q:��q��	�h���/^�{��%�ws_get%�N�~���b�HM�5TWf�h83¸�&�j���=�7�p��J@7����*y^�0�*	�5\�q��Ͷ��C��]6|,�"�ʧ���'E��i'��@z��q�_�C	�⪒̼�ꛬi;����Q�N�\�����K1�fS[���	�]�X] ������V��7�\��Z��+���e5�)�>"#�M8�i{
���h�3��3 -q���"
N�@���I�����>�A��3�)�E<�x2+�ʥd�'��Ճe��e�o�dse5�vΛ�� C�5}f}S���9�}�X�+62Jdr
{��"��1�ى�=>e =�8FE@�]6-��W���Q���i��sHd%J���9�@�#�8v1\BukM؃ԣ�hZ��?�x?��k��k����T��!�G}8��I'�- ����gd�>`�׾d�.�-�����3=��"�ӖcV��SP�����ٲ�O��X ����2E�}U����4��N][X��-s��c$遶������XQ�-s&.��b�I���lѦ<-��>wj:EO @�FCy����'e�_]�NF��ɴ�#���F�ā�
�=��5�T��03<$��~a�#c�Z�J�On6>f (�9�G����}f��iFZ�F۵X�e-V��	gz�3��:`���7m�'�\���J�X���ol�Wߡ9kjfMk ��yb��X�4'H���7=�[���?M�ȧ[ٰ*0�a�l!���L�qWҦ��ʉ��}�SbKƎ}�׸�iԗyȊa
:~���}�}V@��s�җ�}�D5s=ĽH#�Q[�0SZ�:R��l���t�w��1�K��������44��:�4��a%��u�{"fU�����-mL�$���9� �4!���sd�͖e�c��Hć=��'�)TD�f �
Vj�S��"!��k6dS��	Kb�����p��l���'�4�x8&%)��W\3@��3|��s�y���M4m�����K�y<���J�L����*.
����y�7�!���5�`b�}�s'f���4���L��ji�'u%'i3��rZ뺣�%F3Ą�i&��U�k��.�6氱�9�<�h6�X�� ���Z'O[@]�!Q7jMha�q�Z�hAz)�saFSG�9-�U�JfP�n|��s��;���)k�V�� ��Z28U {������Z�'S��M`n9��"s��K)���'��L
Ze�K�1��_rI�s\�g�JO0�F�t�C,�����E�;�6m_�x��W��ݓ�� u��r�I&	��0XC�c�k��j߰Y�I��:�dR�m��~#���T-5V��V�S�&>��2Ppr1�e+���v,�jg�bjq�Ptإ�-K���'�%j��Y���?����� ��H5�S�-����9j����縇��;������K�ks]#��f�٤E
ρ� �W��s�&v�'��vR��=�(1�'�)�X���DK}A_��z��K�8�������i�2˝�c�儀��1&��ɇ�U��'Mu�A�r[˜6�Sd��9KM4N�@A�8�����]��}R���5mhhx�mG�D��fJNZD3�MM��I`���a����Ű,~X�g����p����Q)��E��VҲL)�/p��R���g�e��rZ��i��%7��Z�!���Θ<Q?E�Z�,1��N�92��}����49��%1䔶�2F*o3�w�_J��Z��(S�z�&bm����&�Fo��c^3z<�F�8�P�b��� O(`�
�~B'���ǧ�3r��z�xmu�OU��)50L�=e��<�4�������M�l�=��g���f#-�;'�nd��$�������L�,���V8��"��Qe�تy��&��:ց�8ܽ·UU�9�W����6=��{=�*����ʤ�M�P�g �����ߤ� ���� g���Z��NF�������e~�j����`��Y�;NS�Kć �ٸPy�E�#��>���.������x:�G��%�cuB���O�3g�T��5��x�$i�ɒ�*~岕���.$���}�U�d9��.��v��5�σLbV*�sd��F�=��(���F�G<�pI3n���i��P@��i5���|�<����s�
��B�ťi6�r�����~�s��]x�nn�<dOG�:݇o7�=���%3IP�\>�%"vAW�E>�8��G�y��>�Y�D>��0�����8��ۥ��dmM�> �Q�����lin�ԇ(	N�=�í5�&Ɛ��3�լL���q�d����n�fn�����r�����1U�TB�K���P�ܼ�Qҡ��k�	����Jg�������,[�{����3_<�%��}W����f�_mE��_�塹��	TU�������@��q��ε�9J}���p�ׁ_�PGO��YYEw�*�E0�{�f��V�qP�+J�ژ�n�A�U�#:��5��O����eY8��Lh��A_�YY�{I���U�ɧ6����k3d����\����R�\Y���eA`���9��$v7�6->��Vڛ]'u����p�<�L��O�gX�Δ���3_���ǢY��ǧz >��r����P6�.#;�n:��p�G�X�}Y0�ٰ�� �;�9�!����M�{��	�5�^����{��KP�4ذfl�X	G9=��wIu�W(�ә��}��k��k��ϒQ�ĵDv���׵�0���Bɫ\ݸZ�r����6���:SK�Wَ�������Ď�W����.���$|�wS}8@���`zTl�������}���k_+�z�\$_�=A�?��J]h���Hɝ�8�K<l�Y�F$O�<�|13Y�,��Zl �;�<M/cH�B[�0�gw����ύ� YLy8�&1f6�2�����zfxnN�AwB������=��/}<?�4QIk�y��M}�jU����� ����k)�LY���5��C�=f�bgR��V��+�clof��6۵ZF�?��E�1B.����N|�)�<fH�梎��)#�H�����pfe���穝	���	��	�17�����G*3i�*���߇�m����A<�����EXvۀ��X�����f���@�uOQ�h,W';Ձ�	vəxJ��i�^jZkc-D�Ԩ�}�i��J���%�ֶ�v���i��3MO���~�ld9��a�s_��P=>t��Y�|��.��%���CQ��U���¤�����)�G[$�	GEvR�=��+���uio|��J3]�]�]�6t�`N�y��M���
�?74ok��{ ��tY���B'z������� ��1!%r�>ħ=���A�t�C �#��U>f�2<�KdȘ���,J@�,��l?�ot����k�l��*���r��%����NϸWV���!q����(���y��טl�^�v�Ye������>ph�,�)2�%8�]Y-*3����Ů�������Ԅ�ի0�������&Gm��b� Ȫ3�6zS��oYM��j�C������_��0\I����N�Dؤ6���]�.JUi������n��BhИlK4��[�I���V4��C� \b�4��?Ԅ _j-_R����A�>���@[�5��:�l9˞�P�j�WMX�}�1+V/V�#�d�X��Ka��s־��ݖ�3T�'�M0�v�M۶B����#�q���xW7��¶�+e�)��*�0� ���֫���2y���������]͂����D냇_�J2A-���,�m�[-�K��3�j���d���ǃpB�X��j��t>D�%�V:��趒/�������hq$\ �����7E����}~^ә̭�#>CR�b�RR��9S
,cZi]����R��|�ʎ������v�<Dy7g�J�M/�P�Cո�jI�efoq�'�������k�K���4�����
㸡�MD<=���p}���^
)GS9�$�0��-s��v?(��y�3޻���u��u�:�QE��>��މ��_}�-� bx�c�^U�����}��~��0���z���]r}Ծ�*%6tfYό�N!���Ῥ�G<A_ժM��9��Rg�]�@[R{�#�M���o���Ȁ[G��uļ�|����_	�>b�k�v����]���/����,I�U����!���.!/ɻ��J_r1�B��D��\��˚KW�IS*͸%-����&,�D�s�'n���'���������	Y|�SY�3d����0^��rNK�1���U/�r���!��ԃ�ŲZORAx�Ćp4d[��b��e:ܠ�̾�5M�}@�Ϗ9��Nr�@��D�K[���r��������m�/�8�u�����B���Xw�|\GAYR��g暍�׷������	}���"&���u�bYj���7��u{����E)N�aTB��ԻKd�,�k�6)K���t������ͳ��W��>���b�`B�����E�64w�������h����:I���96w1s�1_k�2�ѝb]��3�c?�g]	qo��$*�)�k������9� �áB��T'��]�d���o��m�z���5�����ia<�&��{R��\��]i�9K�dG�Tu�&��}���ܲ�OL��O�!�(;�]�V���s�3�w���RZh�A�xblj���	�X\H�����u�=-�DFl��$2 �1/S�/�w�U��>��J,a;�5}m���� �2�HoU�S��^�fzs
��'m�ؔ>L<�:E����-k8���_�	!�Zm��i��RS�T���P�����\ތTqz�r{/�1�RLZCńT�yy�Li0y��`��^�d�̴;Q����������.���(��99���uB��]�]��a���=BKȸ�%��̆��W�⽒n��Ur�����j�%0쒓b��y�f~�/޼����r�:��V�A!>�0�u[��|�,J2��K(�h�l�
XKf��{�qR��>z
�5�m�p���K�i��nxpd�Ԭ׬4��l9��j�jicbf���h��=�O��&H;Sb"��f��N0]-�q̍��5fܿ(��]Z����xӱ9�Z�d�!�ۜ̉�6$������w�T�P*��vpq��H��>��.����f�ѕ�	��U�.H�u�b�&���Q�n�&S�t��jM=Jd$K4����v�y��)p*<;�������k4{�m�)�'l�I��-~J���+�4��ih#�C�٫;�r������};G9�gp���¤`�k^)�O���tX��<�mY��8(\�\?���LR��B�ʴ�c<W��x�0De������ݾX��)�us�9,G��@�;�@@�ä�5��^�w��F]"�-���*V鵚ڿ����<8��߯߼���*�h��9�u�V}�p͊��`���VL5�]�dB���b�7]��$�,
�AKt��&dP����*FЧm/��ST��.Ka�w��/�/1u���w_���`�ą�w�N�����f��Q�57��ڻ)���)�o>a�G��Q�k�%B	_�Ǉ��ࢻ<��t�!�10���I�'�I�yM2:~�X�(ݠ�'9��2�~1S��F��A ���t͝C��l�����Ѷ,��t��#8B��WF�$���%�gջ(e�	B��MBt4�(��w	�ēG���,�!7+���z���Gv�/�bz��H�ЁF� ����G�mf��OA/k~�קXg�43v���Eb���ٗ��<��pn<_��$�9�ֵ��.���{�f�QƂn*�R�j8���i�N�����o4֦ ��kc �O�W�l��֒��	��Ӏr��9�~�����S��& W��ǚ�A��3�e��T��8x��Vy����D4}hǚ��@���cp���7Z�8R��Y6��=9��!��-��#�mf�\���IQz���Y����Ӈ����kR_�><ijI��g6�@�W����'�T�<��U�>X�2���2����;��}0�_�����ge���>�o�V/p�T�������ЂK�+_���`L&c�&����A�1�'_kOf��'Uo�J+�����;�����2�nw�Oܩ\�"H����O�����B@Ĥ�
��NZ�}t��Hh(F*�'ٶ|���@T%�箛�x�����\tW�H�1�,��u����K��9�r����6qKr;}oDn_�=q�@:Q�ڢӮ@q��g������C�ϐ�l���
l�Ֆ��֙h,� ^9G	}I|�4��,3s 9�j"�z�e5����C�[�W{�n�z�J&H<\|_�z0�����}��R	m�&0`���:�:L�Fa#����w�ԋ3��"��ր?�����}�f�4�SӮ�{��.�}Z��4�M����n�UV�V�u���cy��W?����׆x&,&�'��uA�ơ�c�ׇ�ϴ1������͢��.;���:���HCFjf6Q��>]$�[S9��B��t:���ۖ2���;20�|����R3���6��K�����܎�w��c�\�i6L�>��,T-� 㮕�"�x���Fx�]����,r��p32#��)|���s�U�EӪ����(	�-g��[3��Ȱ���=�(QUr
�R����&�Z�y����I�~7�<�i�����!02�}�s�
Pu�?%�|(G����Ll��L�ko0�D�re��CN�N�)��\��l�́5��b��Oh��E�i-��3�s�$ �N��Ժ�3�0O�쾁��'�1��fܰ�>?03X�~�9��s���(D�������-��G������Xtk�p�ɠ�l0�e����e3�Qq���20�� �%��Q��>�7Y췿s���!�/������c`�*�=?lҞ��T�I�o�-&�C�W�x��|��x�w��]��2��%KQ�WⷂW(es�}n������i��Ff'L�u��t,ns.�����k�.F_dܑ�g΍���)���Ӌ<e�B�*�88�<K�JY�c3`�~�ޟ ���;���#�����Ŀ;#��<F ES�6JS�[��-VmXk���Ă����ײeLS�m�LY�g���w ,V���,\LTV�Q��5BQg�}�� �?D�&lD��N���+�=�u�7^����ˤ�-�}���<�	G��R+���T�C��=� ܚ,U)*�*<��Ly���@��\�����1�����?���8S�O]��댴\em0��+V�ox�����t
��p������GqfZ:S�v!��4�K �s��i�( L��F7�'h:h��&<>�o�T�IK�D>�cz��OvN[�D��٠��̹��V럯&<�宱H�^�B_ת���:���d���T��-J��.!U���N0��9�%N�jג�C�䆎�&����yl��v[٭���ƽ�A�@ʏ�WJ�AP�;#�H��
��yq?�ud��W�>�6yÿS��$=K�	k�8�m<�W�X��s����Qi������Gv��������~���J
��0I��c��=Ž��WQ�H����Ȏ/ղ[�MDh�κH�s�nrŽ�{���@�� fw���;py�l����x}�Nrqh��q�h@N��z�Y����4V;�.n�}1�����y����FZ*m�)��t��#��_e���%�ƨ�N�]��]�%~~��-EV��G�#
�İ���Q�r��@AO�R� �㘤�d��"���z%���{�4�jp-Z,��Rg�e0n��#�����u3����yi������ts��،R,��Y��)u0�ވmAk8d���PM�T���ׁoh�7@)�~��o��7؁w~T�2�K�)i��-�����pC���5B���Ҵ��4������D�a�m	�%���n�>�=]5Mo���t;�ldU�F^��f"մ�ˠ�i#�S�� i�B��op�s��@���k���:�΄I�5�^�<bTW�Ō4��lt��&@�F �~�,���9�=@a�n��V��:��\��a���"����n��pi2�v�F�2��`ָ����1�qi4I�:0��*����7���9���<�ԟ�z��-i����& �������t(�򄌴�����}�<o�`���>3X+�+:���XN��h��.K�3�Pc����N�gn��}���u�L����\ũ4I���p(�P�SV��m�������k��s!�\�-�����P��k�.�B��C���V��:�Vf3%E���(s��:��v�od^�f\C�9�8.���@���<��Tb׀��'��!�Qn�`�,�S x<��r�ğ�j�xz�nK,��.G�{�����T�9�ES��r�)"��/�,��v�,<�C3J{�t���-o�>L����]o)I�M�+6>� ���%'���DԳ�jϮ���K��x�kJ���P�*K�-ģ��/V|;�X�)�#��+������{�J�'7�I�r�jn��]�٩�w�#���X���BIq�"��x �#�^�����
n�ӈu�cֱo2����H}j�bq�V�ť��0s�%)*Õ�PλG��9�,�x��;S�l'/#q�a�u�����@?�C9Y%��oޖo߾-o�~� +n��P�8p�vIO��$�Xl�ۯo����Ş��є�
� F�p<2[Sm
Qm(|N�{����l���O)��e�mS9���9��*	d�nHP�iY3�J��X��bRDYԁټ��	N���ɭ����i����NMm��w,�v��1'4������-���uEM������@�4�b|Qv��rj){^; *|��1��!�z������ꬪ� V7��J���F(�[��gw�O�-�\2�f>��������g�aa���C��gTS)�}��q2�s�n�FN�a�r�*��K<t�39����f<|L������XGD��d߶7  ����/�P�\��zpr��h7�����e��s��=�F�ɏ���V�*Rrd���k>)�&�U*�?>e ��D-�t!s��16K�Z�SK>J��;^�1"e?���%?��N���N68pY��ݻo���,��O�T~����ÿ�������J�ol���N����onI�Ɨ&�\���e������/���"����=\����~u�X�4�1%�6��6į�ICn̪XU7#J_S�hC�]w�ɺ�]td�xnO,�Bvξ�����J����.�<�Y^����>-B�����r~�����)�F��6z'��/X��U
������P��-�kM�߾O&����H��cB{y�/�v��0Y��(��gp?�'��Eը^Ǜ�-�_u��̒U�0�`r��z����ό+��9,+����e�y*�n�KN�m�܈�,ｏ�i��M��PQ[����~����В�Jc(]�awE�/�IC(~���*�'��+AWgT�_��[���<u���
s�����ׄ�6�Fz�G�_��h��e]�N�֛%3�ظِ�������Tl3R4(� ;e?Rt_������<����C�ם5�8�s�S%���~[������������|^�g��2[舾�dHw _mпE �F���o�߼�*�u=d�q�������}P6�Y��x~|N�>���s�*idfE'�a�Ms��E�xEF�4n�N�Q�8�4{�:�ZNN�_1K����� ��~�M��1�ȆFi�Յ �M"~���dvK8l��k@��5�A���jDh�]��w���� ���^m���o�����-�����;#MH)�8�y�.Qj�G���K@s`�%�\��>��3��=>�G���]SN`L!_�ʟ�ڈ�k���le<��җA0O�j�%a#>�]5��t`4;�/?o\_AB��c6�Z��"膫����gz^���/b�Dއ��o�����#�U8 ���ä�8�~���i�W�mZe6a؇��}}�b���L m:�k��2�v���qCJ�!��k*��&	{�bVVM�8�\�Z���A�G�hڟ�� �`w̎Z�E�>�ca��
��%�E|P�Qs��w�8s�9j��D����m�b�D��>��A�q����.�T�;� !���Yb�8�u~�������7�Xa�P ѱd�r����y���%�?��3��j�'L�����^C����5��n���P�����&z:?e���:��4�f�C�3�`� ���cg:�m��!f���<�������@'��2>S6�ǤU���T����I's'�j���<�u��`[h�b9�T7�jp�!a�黨�bͧ��$\v�*Q�:o�F	���2DzM��.
v� �kӹ�p=��l۰M�P�������j���b<s�f|�u�*	�����C`��j���k����������8�����~4��MgƟ�G�wqy��W����_yTt�tF=玕�;���-?r��ty��*������/:���"4�������F�I�w�h:��
Ej4�mʳF.&Y0��`�Opf��φ�ۆ��͛��W_QG3�{*��(�ǒ����j*�Ρ��,�8%���b��;'y_j�4���>}ܾ~�w��>I�>�ָ�=<����`J�	n�IӇ�KW�ǫ?�̂��\X��1��@ ���,��sL�AK�)����^���z�Ce ��½����Ӣ�%�(��
;�����;N��r�8�*ԍ���"���ƷѓS��)ֶ���q�.(3�l�D�dC�+��#�}D���^�뚴��1g���G�a{Ox��|T&s �+�p5{����t��Y�����Am�u��q&�N��P�:&>K<��������J���C���Fh4u�Ŕ�m�s\��T|�6�pM�t�{w��r��=��X�����z��T�3�v8�S��8���K��)���G���~�RJ��O��v^��k��3�R2;B����%��5� ��z�p�5����x-��#^=	�Ѩ���;�t���3W���M���1�~7r|ᐉ"����{��c����V�o�2�ZS^�x��7��%?z1ne��-�}�J<���]������PO1]�@��>j�QrW1c^��蕉`ڑ'MܱD0�8�����o�F����C����`�BN,j���������>$��N�Cn�{�q;�)A~[Θ�a/�P���=Ҋ�2f0e,*:k��뜳�����/^�~Lѽ�Fu��}���;C���%S0�h���Qih��(����U��m����u� �������)������.�L�t��Kx�1	�[����^������sׅ:��b�mZS3U��Y�b_�Ȗ�V�8-��]<��<�#E�;S�E^&@l(m�6)K�Q��(��	O㙊X�w�|7�X��6]��d��X�]Wv�Ӯf�_��ͪ�����@fGMJ�S��Q�T�J� �����p���r�񲛨��a��E߭������)ѹ�-��"h h��ق)��� ��sH�1��bs���V�2�TRpk�aC��cŔV���Q��/DC����v�댷�%�����YRŏ�O͸��ۤJ!�����!�_Ra:��].�t~���<����%��nAb��rV�_c�-���.�����z�uz��lN�S�t����sj��}Nj��U�Ÿ�h�L�9�A��"HM����fx�)��	��Q��v��1#%�T(�%�\���E�|`p�窻��KdT�[첔�]��P��"�Z��#�i��E��{Uk�f���	�i�5���]:;�c?�ڴ\��x<Z����\X?v
�t��Ӎ�!��5�^�������*��?N\�)�`�Ch�l��a��?��G#��eWϛ�<�8z��)Q����gv�%ˣ5�o$����v�����KM���ؑ�)���7p�J�UGM�!�YQ,�g�g�'|G�R)��b[���Yz<'h#h\��nu|���p��G @�v�mޭ��$7��N���ٌAg{�wT)�  �8�|�F�d��ap�rd?�Oل!�Li���4qU��v\�C6ָ�l(!X"[j �����i(O/�x�BE�큀�n9qm�_V=[�O��
z���~ `��
�����0 �^��0K����0���4���􉃑�����<��Aa���wI���A�`��C(�K��ݴ����uêr���� d��S��Ug&%,�x=2;_�9�����k�e�?+���`7�B�~gP��?�QJQ��>�j���G����I!��s`��Mx��JE���?&�;����4�8��G�`�4�>Y��
[G�4�C�v���5�ڃ���P@�zT�k ->��/jҜ�%	��P������L�����
Q�\-�m�a�J��&'�Z�Z������bQ��"��5�}t
��#����b�XPq�.y��9��x^��O/^�S#J��MⷃrOLid@��)o���Ǔ��^�1SEKN�Gooz;������_���g�fIC��|0��)O]�֪���ߡ�:Ӫ���'6N�o[vv����	��Au����ߥm��l7N舕�*d9e`���H�M���l��sy��W� �p�|����G�5���±Yiǎ�L�� C�nf��kbY��E<�ʴkH��&?������^ۑ$I��9	�Y���|�=���s�av�{���d]TD�,�Y3}�E�hdeA���TEEE�I<`"����{W�)[	�p��fe\��1>Hj:	�ȡq�7���6�&��xs[5.��ʾ0�l��6��4�*�w��I��B0��0�#e�� �EQ4�D���>���~ q�AЄ�O+���^C%�����3+�R;8��$���+W���>��(j*Ji�S�F�H[���$��i�d���&#5��&��OOt�����J�I87��f}���.Ū�t���U�O����
���	��VX��j������~�瑪���T���%.:������綉����[����g��G�s�)26H(iFpCѵ�N��c���?%O����f�a��Y�.�/��Ϣ��=�A�M�^�y����y��u��!]J�GZ�Θ�hF!�{�ρ���w�i�m2\ |����]g�is����������oݳ��#�.���(�I׊�# ���`�s���	M����Q����:�Jպ1"�<�����L���x]&S��:�kř���.;��^���j�*�p�܍�P#<6��9�L)���$�4�Yt�4�:)J�g=#Af�;ds��߬�N�P+��o߄���h�n{�!�3\362�H$�u͌o�s���Ѕ���*�Z�������~��>�m�0�(�?���9�Z=w����i�E�V־f�K�`�ʣ|3���m\D��r0mJ�8a�鶄).O��'Mκ.k�P������� i5b�8/sf
�(AAA�.�'[����_�?GG�%۾z�����Jט���NǰP޲�(b2�Z��Z��%	���>�e�mWv�3�A��^�LnE]Rak�s�Į�X��3�v����S �ۥxC��cg�$�9>�P_p�B0C�A�4��)C�]?D��f6RN�=�FdT M|߇�K��LX&��:��+��I鹣u�*�e-o׺�Kut��&ˡ��gb=5Sv/�'z�T�w��W�s��{��V4�>�*(Kǐ���0��=g �
X؝�H��r��:�ߗM�֡�%*�\���_�z�����D��������~��]�;���w���C�T��~�)��ł����d�H���7�XQ��k��C:
W�x0�2��4���?�5_C��,���bX������˷m��w��#���0��_��`��}嬕��������"�I���"�X/��J��74n��[+�3�[[�a�M��'1�}tH�-�y�(*��)/A�(QR۹��+hz/�'�a ����t�n,|<U`<��M>���dJR吶�)N��$7v=e��Fz�ṑ�r��$4R�)�"���Y�9����YZ��/������~��i��c� � (�@K����3�Ev��e�����������E�$ϵ�:sn�z���d�'ݎ̓�m纫��ns�N�*;�-�.i�?e����@A�v��E��WT�Ᏻx�����Q��=��~��(2����^#W�=�9\Ʒ��A7��2U���^�w�Ux��^��	bD�=X
����
P�2��;&�29����x~���4<U���Y"*�!3�6a��h��}�r*��]�? q>aUYL֋ l����Φ��
�5��ן6����d������	L��1f�"�˺��ҷ%��E�����:ɗ��2]��s�s?��WYs�4�HwU4�6�w��"^�i4�>&H�8����L-R���#���Iʟ�S�xGe�#�43��&f�Z~N� �T�?�]���9��3@X��j�ݼ���R�R�x�˅A�WCd������uL��v �q8?�z�l���iE��?�O:i[�	��0�~Ն�^+g�q�y�|��rQ�#K�,�7i��03cp�>w�K�T�gD�s��`�i�iu7�����0��Z!�Avǥ�ݘJ;�N���n�t��M[�g8�$'dr��쁅�'4�l�;����\o�}4tx��om6�Q�:��fo~�JGS��ÊJ�3�a���p��>�L4|����6�WV�z㸓��tZ)�Rj�i�hаy��O���ǽ|x�X���*�Is�N�
�������������ĭo�o�ݟ��5�&0�F.d��g��e�ܓQ%ox[���M�	�ߚ���+V�!�%"M�|�)�fS~��0����1�b�$U�c�,W���S>DAJz��#���|�n4��㩋 �<@��S+VX�c]כNe�g�y����g���H�>d�v��&lU��zr!��z:wWU!���4=�90�)}���EҬ��/w���w��ZI*������5�c݀���ԯ<�f���UU�J	?����1�a�ǥf���u���۔�F��^т���5\�yn6��冩\����~�L��.2?sC�l*yOz�u��,c�lDU��!>SCi��T��I#\K6g�e�Z��}D ��	�
�t�E���w}�_Mi
f���l��7$v�jx���E�;56���1m:9I����V�}���\y`�~��ݖ������/��,r�nu%c�I��4�̹�J�n�H�\�_dnFw��RT��}���Q��Yu'��\�Gz��v3�!΀��j2�����?G7?�z�<l��wt</(!.q����Yt��~>�~�/Ȍ%�wo��F��>|z���pO
��}�e��ɛ�>R��!���t[t�_8�	퀟~��|�����>mY�p�2.Cfj��I�� ��ipwO �&3;�$����v�AYB�ߟ5.�L��a<`��d�k^�	|�,�JP�
�zj�Ѫ�9/� X���N
jr���:�mo���ܓ@~a�Χ�>�4AS�>+wVG�|'\��3*�K��w��.2{\S�N��� v���V���|����t4S���� ���$[�������kx�륑b�B����f��t>�A��+�V4:�9Z*Wqr֥]
)ĝ�2�AJ�ˊR��2m���27�ێ�r�$ׯB��m��n'2�ei�˲ˇ���u��f����F�*�jb�C�� ୕6����7]�x�Ncl���	�ޕ��**�Oe���P2����Q�
�r�U3|�P`Q����u:(����C�g�I�����R�Yv�(���@�_�i8Xp�M�Aĭ5+F4��I:���U�;���������Rf���80e���ݩ�3	��Ӽ�����A���xN4�v���������~�Y*� )F<�Ɇ�/~σ��E)֌�KWՒ�p��Ț ��5@��>�:���
&�t��c��qϑ��?ż?�w���*C�Y��� �{�PL)�q;;+b�E'��8:�۽���������\��OSn�N��"bd��C�F��z,���u�h�5bZ�����>��xx%�7U��b�Y=�e1�p��H�棓���U�h6�e+�j���;������gM,U���R}�����ƭR���2�Z!|�_�W]{㤼�~!Χ ���3RO��,]�����P}�o>�_gQJ\ގ��"�̥�n}�,�+�2H��0 ���#;��]Ⱦ��r�y�;��I�S~���q����l��ö��ȱܝ������_��������-t���S̶�D�x���e�����D����a�<.����>q�9><LA�U^!���e��>q#AAW?�8���_9��,#����&n�I"& �k s��v�k^�v�$�t����fU�c]O�Fp��u/û/_�D��t�l���Q�y�8{R|�Y�nZ;x��*[��sMB6��%�w��jz�U
8�?~�����;YĦ���'������`~��4��Y��+5�����LoB�� W�*Np�IJ��߄�Q��s�f'��A5��C���6��q����&�Ki�3W�Ff�s�����z�����,÷(�~��9�yW`�Y*����	H����xb��VUk��u���$:-N�,{is��g��� �C`��u��������v^}}��t���i�����^*��g^9���`0J��b��@�@�Zm�ٽ�����qm���%��v�R��L��X#���=������
Iw[f�>(J��7��r�y����t-��?�ٿ�������q+}q�8������ز����s�r�5 ��4O��b�<�/���%��%_̾Cc@��h����������c%�&Nhl���c���;lȤ�������>��
D�I����v���x�X�O�yhFV&\oi0��dY���[�U�`�d��"2w�!Sqc����=)���2�ޝ�o?�Wٺ��
ci_�XLA��o�&�:/�m�qؘ���~�g��2�@za?�FnW٪��h���^���楸d�h��R�_$��wc���X��������$�N<lb_��V1:�f��r]p��c��d8ßL;�n�jw��B�>�M�D�X*�?�����,`9^ja$꯺7�-Zj~ږ������@�'���-�f]nL�B���SdDA��eDH�5���I3؝>�*���'�_�!Q��j�BD>�J'-��M`�M�A�ԲNc(�G���顜� 5<�z�����
#��54�@Ei�I������?�������@����	S���9߿��F>��2NRL*ɞ6�lD��T��yfs
_�8x�_>�2ﰯ�t�F9渗��A
�,��%��EI��?���*��Kf���s�N�B,����߱�F�����Q��s�C���1Q��L���h@�(׮Q��g]��ڇiov�]y�U������}&[���	U�����Wr���m�n�����1 R7���+�v�eiܔ�1�3]Ū`��c�-��0{_ҋ<1,�yN��h:��t>�b�����2y���Ƹ�{��A}����h
�{u�8�i�:�}��
=�<�g���[�{[k�LB��k��j�ۃ}l2��V��j۪ +�7�^�����zţ?ID�=}���Z���n՚��&���'{�_(;��ဠ9�oِ�����p�Y�j@](���5ښ��=7��N�K�"w��83��ih5��=Cl`��&x�S�T,� ����΅�¦aa"�B�r��?����Q~���#�3&��?���N��ӝJ�O�s;�#��I����{MNu����>]ʗ�)`�о\Y`�(^��1��턗�.z��;~��~�B���
�K`��}����|�Yq�C
��!�q�B����5>72L01�R/ ����p8�s��_,Gyj�WC��`����5r����V�G�7iM�^� �wp(9��Sn]� v\G�925'9��J���fs��[��3����y|���Ý�	T���fw֪(J"����]H�R�T�����8�v�� �����3��?<�G 
r� �`�������;�#���GN�u�c�?N]v���T�m�/��Y�$��l6c����k�k�����2��v�$1%ߎ��Q_���TiT.��o���eb��5�Mp�DM��$e�
//�lV%�d�x�������q<��K:<x��
���:V�کXz��6f��<��aBaJ0[��d��((ːaOe�扌�ܫ��uCS������"��b�x�e�wЄ�]:�t8
�!4�\����(c�|�\�-�]�_]�U�����!)���=�E�/75,�vz��%1�� /&0�-[9C�s	�'�x��|�#FN�7$��|�j#�K37zm�^����1l0l�;���n���u���ρ�Rq���lҠ�k���;e���7w�|tŢ&�e'B���V���,<� ���*�C����矻,�I._�`m�r�!N��j�a5��K���;��E9�\S�|� 5Q��Lz�ES}�/�;\^�Z��hG��g��9�MoI�I�޽
����O��R�j�[��1�#��J�-^ږ��U$� �����?SK{Kx�KJ_�S��,}�8��1N�A��y��O�I��1[�O>9kK��;��5 ��&� L�󲞢���w����UD6��u�,�����D�C�����q#��B��~x`Ge	0V3J��g)�ܔ���&��`�nz\����}ϭ|O����.�9�+]1�X��@��^D�
B=���-"3�˺ُ���AW2��x(���ii�����E���8�/k\я��iv�K��r��e*)O�0wq]@$�ߛ��k!�޲J��R{�9gq<�Կ��c�lb3_<��^e���EpQ�}��;��tȍ=�I����6�����h���I!���Y��@DJ1n��D�$^�*L�1��X�]��v��#l�)�1��u�:R�֤�x��|D�(�k�)��5}��0���:�� .q|�O���j��*f���߮�op�6�d�����u�ɝ3g>9J����Õ��@�6�g��ȟ;i��1Ƿ���(�<c��%�A�k̆Ƹ-���'���X����5�=��~��tK ޼Z�5\N�"��-*�w͘�sv�q�7ŵ!�����اǓQ� @�uX�Z;�x�uK��+��$� �'����lӞ�T�y�2���sX�O�u0gP�����a����I�'}k#�X����:�n��d�ꮿmd�Y�h:��r���i��ف�@Y�/)�LݓC�"S��w����O���V/M6�d��;���~ps��JN������8�Y�@7ub{F0��E4nD�i2-��ݐ����H~4)v�hss�͉%������CX|�PBa�.�R�{T滫Mb�x.9��r�B:)yJ�Q�+B���kb��U��>�-X�����lTe�m��v��{�=�_Mi_;e�K@�xe��Dn7�pӀ��.��D+��{��r��t?��=��au� ���n���!?P��H�U�B�ˎ��E�Y����ɑ���4/���9At���U�Hi��t&���Gzm�����o����b��CRu띑��D�ׁ5�vl�[k	��x~,~tϱ!�]��U���d��9M�X!P��^e`ڏGy�Y`m �ڰ���N�wC�8��)��Z[׍Y��8L�h!����&��۽�T���v����1�	���N�A�4Y5$�g�*,kN��������<	ϔfC����A��̒]�9,���c�O����4�Fʠ�!�k�2�{�T��~4�i�*3��+kf��i�Y�Y���B�������N�9�1Xdy}�q"���SjkT��9�6�r��f�QU�xq�����L߳jܺ�e���_�������[?�d���ԔnU)_��i��%���h�����EtG8Č���z:��ۈ7V�d+�4&`����rf�5�i�;I����7~h\w�,:��q���U�x��otI���c۱sF1���xXn0�8eE���G���^�$���3�Jf�MY͵[C�=��&v?�C/`�9���¾{���l�E���f�$L��h|uူ�g�(:�p��9��թ9��w��c}ob��4���s����q'Z�-�������1\7�T���k�Y���)3�~H��,ӋԾ��S��(�1�N�R~����s��'.e��$"���I�ρ�B(���#���hN�w:%�M���U�g;ꖵ����c����g�~)�߯�z�QF��������3�mЇ-]��Fų�X��%��	ۍ�l���zm�R1�g3�!$U��˾Jا4��ϑ���b�S�)�f��*����Ds�8i}����WN�V�Vк�ʚ2e�Vc,N����}|Rs<rigNy�ԓO!n�P ��?�:��h�&5���j �ɿ_�=jr�1���Ԣ��s�L�%g�$�9);�n�0X�I��᱄��y�;�A#�&薜 �b�UË�*C<�J�'��s���m��I����-��~���~JQ���	��Z)����Մ#����{(�ј���:�["�YS���M Q5��\�fk�u����K��,~���7�3h����d����s�^��_q3sȩ>D�˜TVH����gp��� um0�R��3��+� .�q7����ϋ���զ�&L<�Z��X�p,��0/�c�ሻ���>k9O�ܪ��yni_A=\Ki�Q�+���5�q���g�g�;��#0�pR��W��l[,���\Ҏ{M YYo���z��g_�0�5��Q��e�����#.�g����f}�ƥ�5.]�$�*ߣP���c��J�ͰWL�8mY�5&��ǐ��S�N��9�"�hC=����[�7���#0��Jn�m��yf@�˝F[���E�S���Ox��	;�|�yzƻ<������"P����e�^� `�I%[	n��0!ٹ� �Q�S%�%�������Zf�����R�"])��[ m�l�=���~��(��ձ��c��*��C�kpIn�{��^��Y��>df������9��b�3�Uv�Ywj��^����OQ{<vE�&�*�\u���RXyִ��,�s<(#��(dy_<Y�,��8#�B`��}� C\�
P�H<�		e�P�z��j��)�tzIA+�ה��
~��&����A�CP?�D�Xx5m��������ϙ,�Z�W�Z"����Ƕ[UK������0���� �Iy#�Kro�cNR_�e(W��9��]���q�As�P@u���µ%R�sTzU%k[~/�hsS�{`�#ۂb�U΢�d=����
�K|������w˜�;�sd����"����Y�f�`^��/�=��E:����2.�NU���p���%��ך�#3�Qx�;Ü���'oķŭ�d]��Lu1��Dդ\�2�v��8x2�i�-�m� ����IK�ɵ�4w���R��gUV�V5�`�u�Њ�p�G�����l�X�����k.�^3���x����s��Kg�r���`�M@�N�+��+ENju٣��)]�d)2�yN�Ӳ�G0逨\�'R�0�4#Q(f��s��Y��Sy�0[3�*�I��e����/5#��"��η	U�!v��?}+�&����m��s�~��xRlRg�~��`ĲT7|�#��8Ҫӛ����SF�|Y_5Ub���!����<E������X��yMQ�g���-���"������K���Lx_)���$�x������tn6����p�Ӳ���&��	|��jY�o5t��vF�g0#�Nk�t�Y����hF�`^{�02�P��᪦����Zf���1\ K
d�1����U�,[d���}�J�`�|G�]�6.x����bD�����qp-�9{	g�Ti�!2eWf�_v���J#���3h`v;�`�=���7�k��]�Ed��2�*^����~���R�2G����+9+;F�I�Y���.V�wr��q�e�i����#����j�Qv��H�����g��NE$T��§^ι�>��a�É�T�Ⱥ�|��f1�zOy�8�7+�zo�؛��U`4����D���ƞ���n�,��l�՗I�P�!�9�q�WJ-���kD���<�T�����Sr�4i����t&�!���� ��9�����c����Z��׿� �J�5�ٌG�PJ����)t��ۣp�o�l��M��_C�Σt�@z�pσJի��3�T���L�`�x��4�����"���T&J*�1�Y!��+������jS�2U?�w����Ỹ;q���տ�����R����sL���KY^�h�\E��|6��r�*���`z��Ń!��@�&z�l�,��}�-n���6�}TD:d��FP.�Yr��,�S1Z��G�Z��l����:Q��	��,��a/w�52I���+��.�a�� �����:}
k��-����y��0��`�3>&D��^��u�Ux�l�<x}`��F�k�S������π�l�.����<�e��Ȏ�<�k�2OH�����n?׬6GD+U�[!���\�k��}��8����m������y�b~�rS�s����`�]x��9^j�`�jv�,�ܼ�� v3i�l�_`CU�b�C�=���+���?���g�����B�m��MCΰ��o��Z�����H��熒�D
�x�oZ������zs��zyvw1+�6�YaY����lr^���7e�^��?��s��OP���?~/��;�@/ �4���UF:P�g��%Fp��|�}��o����������Y��j2 �B��������VV��N'7	H����yϗ�e��i�>�L��2�o��:D�b6X�e>Z*Ek�S�3:�b`��2����E�2�]��[e��Xr�[��PX�����Sv1A$�mdj��_2pO�9�$�F�i�H��m,�=�k� =`հ$b��5�L8c���H��#������/����1?w	M�_� �ۥ_t��y��w���:#5��b����Ig�HE�Ǫ������ϩM�8��Χd��\,�唋�V
���3�Lk��U��Dpnn\Xa�x)Z������)�i��<��� bG�=p$��4_���%-��x�]./1{��K<������TTHoE7�#d��A�u���6,dʰ�L��6�_�=�}��1g�B�˚�
���ݹ@�p�t�C��8H�U�l�Χ����i˸?��,!ܶ����_~�F�R.�w]�bZ���u�EN���>��������My�?n%p�%����9�`~�B� �	Y������C�-Hu�,���!���ch����;��C��޴��TY���Ҽ��������A7H�
�YҒd�@��f��.�1���2�^�~�6�ٴjEj&��-Q�+;[��XK�0y5�Maz���{R&��u�'�G%;l���KX`�#���T���G$��)��2���u���)��]�;��ܴ�. .(o��B+m�A��lJ��p\x�]/C��+�#�0^���I5����/<7��Fm�����-s;�V��=�*P��%�e�� b�\�_ҵ�����&n8Ɖ!�.������l9��@*�(��zg������@
�P4�5�6��@ ��P�0��)�it+w�@�����@�,��ᰋ���D�}z��|���x��c�����P
N�݀	bAl7~ �|�Hs� �Tt����Rg�c�@�Yٛ�2g�J���L	bDHQ޸���m�T�<w��9�<G0mC�]��q����u�>K\L�HF�v+^<S@��s�y�OUd�?|�v�0ᩤ�?������~;T�	�s�V�C����1�&ͱ���C���H�.1�ET!|�@�����vZ��ԭ骡�[�﬍���cC��qX�w�D�hL�#�O	T�'��I�Kxl:X���˵	�Pe]�po�F�k�p ͉�yJ�'])I�+������xO���)�E��I�N��Y�7W�h
_��}���i�����v��#���%m�9�A�r�d���ҹ6��y�"�ax�mٰM�b(�/,��f��?���0�kd���z��7W1h��k3 ��vpd�ù��7�0����Z_g���.��T=�։�f�w`q!~ S��!���ٮWEsJ�%��\�q���i�`�/6A7�QR|���ȓ���Jz�ة?D����Q���:
��?A:��q_���Hˢ@z��Yi4��]���=�xB{�3K$���ve{?�بo�Ǜf��u��=���Kd��J�|+{�E��#2>*4f#�T.P���_b�g�"��{�-�sN���������ݛ���o?�_~�%����e�J��P,O�w?lY�����e����\�,tQ����=3�`G�i�NT����ɡ��Ʀ8��hL�M���
Ń!��P�
:�JM���|��lh��e��p�ʢ�cj>*��tU��NR������I�W�Ʃ�d�!9��f��A���r������:������MG\�@�U��.�*7
|�\f���?G �����~�C5A�_� .s��1�Y��gZU̪����tFe�L�u�r��1W
��1,���K���N������
����2/�V�k�֜����fiW�&�_RN"r+���a��1�׾�!�E��Z��^��3�}9t{��Z``k M�9ۢ��O�8V��U2E$�/���B�׌�)1��0#f{�R�aVJ��52�lܲ�~.(�q���Nwߨ)7Qd#���ۅT��}n(��E	�R�����A���AGEَ)�>����v���b�=�0q�0��� ��rB�+y¸.���ٰ�#�)�ˋ��z.��3s��Ɇ�Y`*D&SzQ�(��Lf�i��wrKg�œIb�>2���R��@����IsE��Z��@�a��ö�ͅo��|����K�`#X*�t� sO1ߴ�f��p�C�U�u2W:O��S�����t��X�a6�6�+
�%���T9ᮻ�T� ��z��\^����������I�li�.m��t%7o�ʼ�ғ�n�Ĭ�i��ÈC�R2��L��y~1�YH���9�:�}��ݫ����Xitb����F mh"q=�������G�O�*�щ�'�a�r�Ɩ:���B*�G:c�\SkjN�,!���x�#��	wՄIX�vUs�+]^`��Q�~�=�Xt��XA�u)��ꋄhDG�� ���m�~ز�-#3�ֶ��M4Gc����\īj	���M���[C� �
���We�3g����N^Q�p�������|Z@d76���S]�6.z�K
;�ň#���~W<�v����I4�7�����϶rt�끳X7A���jd���SS+�m��I���1�PWXgi��Nxݕ�ƺ�94�w+6�V!hS���8k�+@`�UM�����'���*z2�)6�����u�N&����Fgw4q�i��!��|����LV3ȯ�&�Q�<��٢�p��ݨ�A�h�}"˽�� I��\Y&�]V�QJ���>zO�XhV�5������5�vm|�[��E}�E�6����B$�G�[�4��b��j'��8*�N��Ȧ�7?K����+x�m8w�cZc�B�H̕�����6A�X�)�����<
]>��	Z�[ E0�.���!�,�ycdn{?w�&w�_���� ��1�����{��	��;Z#pw���#���$>�z�\�(E�l!��e��vˊ���+
,kB�B"��]4x�����J�8��LꤞԵ��SBϪ]1?�P��I4tǭO���1��K8l��$}Nz�(^���E^�]�_�*́���[
N;��jvZ�����l��/��θ� N1ɷ��j�ʪ��fk��R�JMO�PW�ig��)cx:3�`D�F�d�%��W�=����Ƭ���w�|XG"�4_�o+�5��1L�8���J���8C��OXo�zp4�	�WN�圿iJR	{�g`A4)�w�A�1/��z5�sDc���
k6�U�n�j���&�5���������˟|ys�jX�@3����M��]'��I�6D	��ڵw�� P�m�ՙ�/���9D@��������DYLV�ܮ�0���AW7�73R
#�lt�h��ib-!)�$i=d��fM~��-�~��j��l�>���.&x���(�	�#>P����ޅ�ɞ�Y�@|X|y��ml�"C�6	^):S�mُ���y��3�}jL���A�2$_��C �+<p8a�6 x1l�����+��2�8�Tn�t���ͅ,���*��r�
�;���#-]KM���Oڮ?I�م����,���\�� 9�o���0�f�v��k�J�,�Kt�cd��?��~��?�Ϳ�����2���m�Z���@�4JcV@\c��G9=�W�_q����v�qo\e�y��t3���_~�6�ω�����x*qQ�{�‥"�Kz���A��;�WU0\�)���e�zE�G�A �)�gS�BY�ĞZwU�|�/�VFʘK�`̕�t���.[eD�$ �
�������K��BG'��,s&=��m�Zb�v��CʾA�l�EJ�1�h��K>��W��=?��̿q� �/W�c��w�52�T��>Pc�� t�S�+o\Y�geūI͐^J:� z��\���2L���#�(?&އ��-+-�1A���E�C� =JY@N���z%T�>��zK{���H�*�M�`V�j̢�s���7o�^� �.�n�e.Ehv
���(�����s����2~��46#Z�.Ӌf�`[��y(�Fv'��֠5I�)���b�jt��e|�Q�Z�۔����r1��)��`?�*X��:k�n��y���7��ؽeC!hc�Ú��G಺�ؽP�p�Y1X�&���>C�Mq��*uR�=���U��׳��rjhqe*�m˜ڧK{��3�d�5�5����i���W���IG?��Z��	���`��y� ϟ��lS�^s�XLෝϧb)��S���QX+��2s�\��i���l�9��R�Y��T�&40�G�B?n��xZ�r��l��wq�z��,�R��h������j��C@|�]r��d�ұ�|��$e��.��cjf�>�V�LO*���p��x�Yc��̎Q����O[F�Kd|o� \�1��i�|�{�U��4���NЕ  0��)P��&g��@yﲊ���NG��AΘ��!v-��)��,XDgb��x��t���¬L�fUvJ��p���;؍'P���U���zI�	��!`��5�����v���xp��=�E�!hz���}J��}x|E�U�c�j;�%)�	m�}�$�ۭY�ǜ/
�s�?~.2������+(a��P0c[v�7l��&@�=�(ziӆ��X���?���U#�[��EW|N��������6|��𙥾*�K>�SMi���(܀���}�~��������,|:�cf0|m�\c\����[������1��X�A�X��腦X�^n����D
��pнfnxt;�[��[O���zI��X�jF�S����MbOuV��$�=�c�����<����H��D�A)�	��i�OR!��l&������
�������l?�p�:#�,p{�B1���sՠ�uh�0��*���:��cl%�����^�Hyd�ߘ�57w84ws6D�Vc&(��6#u�R��,O�u]m�}�8X��նoH)�@�������ޕJk"}M��'���D��"E��]^���n��>�oX�7|��u#KPe�(���=M �&�vs��~%��r���*9�Y*`F�{�Ā���wx.��e��<���[z�U3� 1���{��FL��t��x�T�p�}�`�ç�U���k�K(����)e��VP�2Ҹ�-F�OZ����en��'v���� �R�ڣ�5/��,�T�(;�2w�L��g������ ZJ��D�g�Kӫ�6���]I^!3��|	��Ҙ���$x�6��8u�{.#0� ̅�z�]��ϫ$�z
���-�#r��Y��펢��j+��d�c>�'�l2I���nh2ɾA�x�=qo~хSW��'��%�Ʒ*�)M�&����8��"��#���M�kۘ���(�e�:�du�j<6���Q��;���+u�M��x���4�ډ�1g�}k�W	�G��i�9�tc��^��k�V��?S�}�ܜ��v�,=�f͢���A�����и�)D�9'L��(ɯ6���Ӑ6-~�kI��k�t+696�srO�P5�������y���}72������>_�Z����:���o2T<�4�j4����W��(����F���N���t�w������&>\ȬM	�{�ڮ�&5� ;i҂3�T��ԅ6�R���R�r6�SBh8}~�T%� ���&::��g�z��(�I�>�Ɉ���I���.�AC�^P#=d��fC	����2�9f����1�Ȝ�F�}�~�~+��`��0]>�� ���0"}��`2����niқt�_Euri�6��g�&NI⦏=絙� P����g��g��+�r�c�VI�{�����${����(�W���C3�)�;�7c`��'�R�}b�Weie]�˼�`p�fT?��l��t洔U��
8g8
&��z�ϟ3{���5��@���;]KŒ����S5{?P$bax����~���N���������ON�{���{+��>�7Δ#k�R������MFm�V�V�شDd���e����V۠�J��y[�4[�M"o�B�����3F~M�8]��������ec7�7ʬc����@�M�g��4ik��3�7>���2q�љ2@�,�9�PV+�W��+�6?o6Ƀ6�?� �#�����$lt��;w��r�D����kE���<R�=����i�BzpL�&ş�ՙ|���^�ԥ�E>Ձ 6V(m���/P�~����S!��}��{�]�8�	%�[G\Ϡ�|�Xln��}qx����0�s���kmcH��9������F8�>,>/"��^N��)�.���[���=�\~�����������r͌�M�
b�v�C��(���s�@��I��rƾh���P�M�Q���ߞ�*}'�0�Z��uκ\�H�b,��o��rfz��@Z�+��M�����^�,����� �Iez�x�c\�Y����I{Sr�C�{6Ogz7��p6j?0c�9N�} �c�#�,�!^�ą����4?�W�6��F�|��5lW��>��O�m�&�����Z�(L ��(�:;)�{� d���ɻ��_3Rlk~" b
�⹫�^Z�ūʒݼ�����h�t�I�=��[I� ���?�?��#�L��x7�{/�4���[q<ǻw�#3���c�72N�f���;��E �&��N�����H��(���f&Vf6���� �&�_�a@� ����X�x�UR�k����1M�O�w��E{���AY��X��H�tFc\�L�
`�|�/l�D6�����#��e�{�J� $����ֻ�V������5����#�c����Լ`�����ß'��}1F�k��x��9$�.����ɰ-v�1I��#���l	��_<>ݪ�R���5��2�D���S7� e�O���1�cik<��`zS��ͼ�Y��V��i9��y�Q}�����u����A����!�:����TJ����;X�`�`���T%*�G������2Rܨ�@qڮ+2p�h����ė��i�9(jDm���$	��z &��ɬ�N�Bo��t�Su������5קYybrt��U�c�:�i|T�+*˧�'(�o�<mCa��e���M)��4��K��D�,<�kʷiA]m���MA������<jgB��˹|��$�EߝP^
C���yxf����>o�������~8vnω�?-��B�g��Bpz����-?jы���_g�Y�w�}n$d�>��Ŋ���w���҆��o���p"��p�M6�e4�J����ް��p&����0�.�� �!6+��(�l[�,�5Fj��~�.���B;�(j�$i<�Yp�!��U<s�:Ġ��Ȑ�|��@{���(�=f��e�d����ʎ�8h(U	3�h���2�)�B|�AS�c~�M�H{`XSɸ!��ԫ�)D��,v����q?�*{��>�M��'�ph@�|�U���V6��d���C1�k��s]^��7]�t�����K�iy�����A`ۂfH}�l�AsIV�{��-�zۤ+�~[��d,^oy�������%��7�sP�E3�l�v�I��*)R�C��\lz�����&�<C�2F�w̎߼��?[jYh�jp�ԙ!:Ѝ�͠[�lΙm�/�{�N��DЬ����)4�"d���O���R�A�I�7u	��Gᰩ*#z��N`K[f6�.45X�0a�����x�����%2z�&L1�����놛�v_�|9��}���u�A	v�G�3����W~�V�$�3�44�[�]�� ���u�Mm�A!6���5>'�~�u�2��^�b=Q���;&��EJ�n !��(�q��c��`��t?�z|1X�n�U��t�<�4N⸛q�	u��-�2e��J��c �Ѹa��tE��㬾3�Vr~�O�f�X]7ϱ�^�YF[�p���c�\j ��"&dz�&����.|ä��L�?�J��@�u��sOYd��V�/�����&���"k��iT��ƫƓcnU�#�\�6�}T��7X+�7��n5=��䦄�y;�M�݋0�����$�j�ƓLݘ���'{)�1�B<�����=��O_e�s4Xp�� 7=�ٲtuD���w[���w�>�������#�g� ��ec�(_pS��=AdDc�1'�$fM?��d�Yo" 2���(j��lK�y�5��Ev''�hF���^D�:���8��.I��?=��T��Y��(pL�0�B�]� μ�W�����'/3��v0���Қ�sQ���,~��2R��&��9���(��4��[E�����?g0x����Q�0r�	��#�x�(��َ�9>R�b�^�y�M�������+krp��Yރ �/}m���}`�P��3�v�W1��gg�n&��~"������5fK��A{�\��q�}��	#��/����pd�q�b�s�����ӑ-����+��(m͗!V�%�:�XL�D�oe����w0]o�O%#��S���%�F�_[��v�}��S��h:���Uz8		6���҂�]��(nDJsb��ǔ��@<�Z�ܺЏ@��'����]�����6����-��)+]���;�?F�>t�*� ��nv'���5������Q�13��9W����#{��f)X��)P�M�R'n���Z�%�O��wH�K<g��gȡ�B�#8(�c"K����8f�Oa=��q�{\�=K�c=(4�JW�%J�#U��RWao�*4|͹x�O$���^-���g�FYflN[֖B5��4S�%���������j���ԤX��x���R�d!�P2�C;��� ��u3�{Ҹ�����C��%�E�ks��Y�g���D[T�sW)���D�b#��L��t��j�y+�R��?G\��V��?{k���qX/�8���ZI[b��?7���0�M��=�.K��{�l�Q^0N�-q5�DIe�j�� Y��J�^s��D���S#N�AΘ8��d<�}����փ,%&iO�?�����=K<!T��q� ��)��>:܀�ep�2k����������D`�u<_�jw$�u`�猦�0#���}F`3�{��b+cQ�T�D��ƪ�m;D�4���@.��9*K
{<�i9+��m|6b��j��u�)�U�U��D��,1�)N��i��y:�s��if�m�e�	�wr�)�0��ɑ�R���Ig[WPI���[+<ί��(1;rG��t�<�ʤ1�w=��>f��g�"�{]q�A�@�lg�#ѽL%bf�i1+���O}бVA�},��U�ö�x���"��]h����E�4JF�G�8���Q�&�D�rM�c4L1H���
m5�Ӻ�=`�e_
E.�Ӥ��P'O�\���76����M)[�í8�/6�l�3u�r]�Xmi�}�zj�6�+�,g�8�������5�p֚�n��Vw��CҢZ��^��|oƷ�����5d�A�lt������
����hm��W�(N��7ǜ@��)������C|��x�V��<|I��U��ڭ�y8؟���h]�D��â*����Fm�^K�XS/I:M�DǛs�g��Ĩh�3)� �x�p�:����P~`�68��p�ʪMx�cm�w޽{G�Y��˒���׫�)C���
������T�Z�":�J�t��=џ`p�ش�@K�>�G�{y�/�&��M�"�j��l�����2k�]�ʒ~(Ց��Cf~}��a"\v�븫��y�e2�V^�5i��`�ǿ?=���l�E�u��\�����V��� �aٙӄ�.>/ /04޿�7Ɵ�NZ�Cb�d+�%&�rm���}��-��L�����x'�F�`BuK�sHpc�*I����$̜X|��.�J����	�\�Wͦ�+�R�,cl&��9�T�{�]4��YVtn ��h,.��f �w��PZV/�d}���A��5�N ��ǔ���VѶڒ0*�`򶅳�@G�3�o�f�L�"L�DAiBz0��L0U��%��x�xmtÂw��H�e�4E��92\���#^�\)&	6�9��s���v��6����;��%q֮���}�um�Q�Ly�V^ e
4\�OŘ�x�_��	�� 1p�L�2�|1������g�M�M ��X�� \��/OdMi�]�����U�"��ԎY}s�ǽÅ�ld��������;L�8� ��f��Z1m�;ƚg��L�YR�U��������x���F��YP��Bf��	���y��������`I]��z�fX��STd�ځ"�!�A��=�q?2��z��9��àY���+�J�E��ۯ�T��+��� )�=G�A�K�Qp�ȸ%�"|���k�\n����S����zE����L��͊J�qiB��|ب���<�������/7�vX��d>��������w����fn`�����։὘�KU%|]eÁ���"�C ozmP9�x<�x��q��~�L�T�َQ��I�f��}����SLو�~�Rlv�=��猪C�Z�L�a��l���� ��� �k*���P�S�"���u�������%�c/.&����>�>*Z��ucJ��BWt��!���:��[��b�6�����q��]/�!)���2{�	��~����,l,�+�QEM��`����V��\�szoF��k�5M�MB���# Ws�f��C8�	B�r�xf@EjL�#)��a��������U�ͨ��`��p�p�0��'��R4n_(�XJ��1���L�� \��I����IpCi�* 1��^$\�mV�n.*���賒��u�Ʌ��+�>T"���}�D�#��۰^K��0��SZ7a4���շ���?�*,��fM��s���	a���b	���F~���>��N��]i���]���T;粖<��^�Bn!6jb�����-����tb)l	�(w��G�*m�ÉO���8����{l�]�_�ŤqB<_t��C%oG U�0���c��{������6�'ܼ\�1yt>i��}-��ذmS���Q���i�V�|U���S�)���&��jD:S25+��+E���!�V:�J��R��m�4�����F3)�OTosʌe"�5��'��4�vV�
�=L;e�+���}<al���~�C�	���"p�3-5��>h?$|��۟NɅ�ʭ���x��eפ�]������t+P ݿ�%ۃ�iנ��AA�JU�m0��J�p �p+�VȹO�P�{��[��H \c���}�;M�տ��d�?e�m*����G�V#�)�o���#c\��}�r���Ԅ�z��<06�<e2j�mN܋��wS~��@c9f���FV�$�v�ϣ�)O���\�O��1�}�H��`LC ����v[��.F�{��-!��[���d.	E��!���K<�.�C�ɰ���h)�^Ʊ��鿡?e`Rv��=��x��q���{�ciu8fi��XZE_+/���Iݜ�����2DI}U���.e��G  �N�����,*1�k���BZ�HN�&�` ���w>N����pH�典�ul�&s%����1_<0<�M��L̎�����Oze)#�ӟ��#���؈�c��a���>���t+X�����%���bkl���ݒT����;pƞiF���}��V�y���x���up}����+�~�������^���uS�n�k��Kl��س�J��������^�������N�Q����zpz"�;Sd��X�N`���������h��hS�XZ��6+]o���l��'����v���X<sݐn��R�O&���ߤ�Ku�n�3 ���k>������	��%��i��z���S}lbA�yL�G��q���ze�?1��*�����b�\���Z��7���H�u�ϦHj�~K6E��̛j-�]Ԥ��>cJ�����w����oݨ%Oxz3I�|�*d!��n�{/���~��FoW�W6<	�j�!��]�Փ��_n4Fv�W�ǇIL%�����b!�J;�D����L��ǽ�w�U���FsBTQ�`���˥w�P�Cs�y��\}ש�P��RN.�S�D�F}��	�8�4�bv��y(�	��'�	5�9�eC�O8-�$���wM�hYd��=d(ёǥ}ߛO��)��o_ߢ4k�\��U�kڃ]x>��i{>~4N�8&��S_��#�8��T�Ab�)����SG.�S��1վd7�⯵���`$���a񺝞ٵ�c����k"��3�[}=_�]���c�rO�YsP0���(N�>��3+���)���ՉY![�L|��{�c�Z ;�0K��o|lR9��T�k�μ:׽�H͍�P�!�q��|R���=�؝4�p��El����x>���C�büX��㺄p7�IL��sC�6�12#W 9�L_o���z���w���cB>��&�����F���[�6��"��z����O}�Z�b��2֋��yp7zo̮��z_�ه�P�L.�vX--J��E��@�a����3���m�s�*���5ýw��d�ě�A%��*.ܿ�=�
���jư��ʣhm��KMZ`&Zo���@g��.��}�=37��U�>sғI�)�����Yw�������^�3�֩��5���f��U�������im�'��=	�*9�B?���E�9�pM�]��_���bFAw��.@y�����ǆ���v����-4�H8�F��(�]$��xlԧ��T>���I��X��4�X��{*O"n_�^��sl2��¾�6����Z���MS,ED����ݨ`��B1�O"���QSC�KC��`�w��I-ߖf�kk�&��@5��Ȟ���X
�/�&�8r���l�x�t΃��1�7_A���s;��1S퇍�C��ȵ��F��B1q[MҸ�3����=-Ό�!I��D%�zP�}��Mڱ��w/GL����F�+'	gB�SrINE36Nو:����d��'m�&X~�?<�]z�_�lk������P� &�kA
R�?
��=�4��	���j����h����8��_Ͷ'�4�k���I��8�R����S�L�tU������kM3~�4(��d��v$������7��T�6�.�=&'P���{��E�H�@�Ы<��~�,g��A�29-.�=͑	�cX��z��]�4:0~���~+��Q���	SG�����^i|��7rU������9S�N�0S̔�45���;���.<qcQ�'r��΍�K��԰��zV�������*��Z�u�e��Mðy6w$Y�?7I'�n�A�������E�x��}p;�l�ϋ�x��Ld���� �{F� ��O�ʯ��z����G��`�� lr�{Џ�	7��K�ӎ��02������$]/t��{�֏]Ј��M�.���D3� �D�@�.�W�ŀƔ��*���{���5���Уows͜i1���ݮ�)JY~���6�)��/̸1��@2!�W;ER�hD�lՐS�ɡ�&L�j���Q*D��C�y��,�кj,���G�!XK����51m�(�(j?e��� ����W�}m���JqbJ�S٥d�R��/^�甓:a{���s��n�#d!nE�ĩ�]��B�
\/LT�cɮ������>���Y��{�H�pZ���h��f���=nA��1�v�_b�b������GPy�n����PUq���Vd�x�!tX��L/=4=���rJ~溊:ӑ�o^WY�z?Un7��z�An�K��>G����Ex;�Н�E	8�&��s��~cנ/lЃ	��k��;���=6�:xO��~/�ZX��8���m��SfTlz����$[��]�2tj���j��v(�w�^8������6�#�&��t�Q�����>.%�,"NZ��!�Ϩzt�^���\Z��K&nf�B�0ɔ㥄�(ޣ���$���"L����P��8��<t(��J0,�ܶ?��;��A�3��59�.ߣ1�����Y�$B��.qO�ڥK���Y�7�E�3V��/�N[S�ȁإy���&��Z~ ��f�{3�c��� M�pw�n���ȸ:�J���|�~q��^�װ'�PkQG7��;y���t"��q.Ҹ�p�02��  ��IDAT���~ FFX�v�Tו�N���;e3�SG�Z���cz$�B��!H�g����c�
6Ps���!D�\\��!�҇�o�,&I�ɻ�tE.*/[К̄!����	(�k��&��ǃ����H3��;݇��.�a��y,�?������"VMH�����MIT���CmԤMĶ�Tx���m����௎
��s�K
���cN���}��=���� ��C��cα3�Y��N$^Y��\c�{��`Q��9��5fs���!JT�d7|y�߂!� T���?	V"�f5�����7����"���˥����B�9��y���$�N�w{Q��4�R}x���A+*��q�s��{��1�<���R���^����9Ox��P�L>r4� Q����.��[+;3n�κ�3G�C�F�"yE�}��U�WEV	m�.�u�E�H}��:�6Ğ�^���ʭ������I�h:��H-�onr<,l3��̖%U�������ę3构q l��,��j��h%��M7_`=�W������	�Q@f����{FFzO��I�2Ә��2Q�:���s��#����h=����O:j��I���Z�z��m�����>K3S:�>8��e��G�#�
!�z7�[�o�k������P�rז�[R ��}��I��|���U�Yd�[���w������ ���6$����ӏ��[Ъ�������ߛ*"�"sX�EYG:On�E�郦�P"V�0x��5���~���}��W������C�0tQ�XY���g�������S�%���;����iԗXK����=���oNuTREfR@ΰ�����A�8��^B�L����R8��	���5����a~Z��>�8��Y�(.RI"G{[�{R�&{X�BV�=��4ޖ�E�y�];fasO��&��x�>o�<�2�ه����2�{�{�V�%�H'eA{�%��}��8�q}���=�|@��}�עnh��T/WfU�z��d]k��R���3�I�ϏN�1u���N`���I�/�$�v}�N������D�>�s�+ �&�~T�PܽA�=.��k�٘S4��jDP���.�%P��k��Ut�,q��I�ӹ��@�Q�:��	3��v'JLbq:ÇI@���xe��e����q��C�s�-o+�ʤ�[���.�N������Tӿ��������Z������n"~�*(�w�O7D�� ��{��*�%No"���=ߕ�=6�$^�E�����t��ڮc�{�m= s�񅪨nd2A��~�&]%{��l"�V����%����sm��n%]���}9���=TA���7�j���٢�O��-R���_�4p�y��d�t���0XH�S��.<3�⾆�����ہ_�e�y۠{�}Ϸ��{t�E�����}�����GZ���Q��0X���o ��A�7C{�J�]E"?�Bj��S�W{�JИVMU��Ҁ���Y`��)U�]��;Z�h,!��Nz�̢Q�# X��ٹ'u���\c/<U�;�j�A3�^b<�c��ox!�:p����C��exo,��d><��&s��q�T��<	�%c`�bF gss��Z)�زD�ObN���"�R�����������Yq?�����Ӏ޼݂�{*�G�f�M���,nB��u8�bY|/��1^g^���B�`�*F'��-����e�O�p䵛d�r���$��#��F\G)���-N4���T�9��F��t�s��u�N�ֶ�4����y,���U]��٤�8�EzH	�3�_������3��R�I�*%��"k�~�����g��n��X�����OټTCj/�6���$7rsŔ���P����uyн�i����6o�_��W_U�$�u�ɛ/�BϜȥ�x9�4�"gP�E���9�(&^�}�t�W iZ��ɴ�]�ى�dUn�=��d̘JD#(=W�%m2�Ȑ�ϋ�86�8�P�)�e�ۜ:�T~�2�ԝO4?l��v��3 �������V�q �&-eI�ҳ�����ۛ��En��PG1��F մ�ˇ-�~��r�5�(�� Ư�&e�Ĥ�!��xMd�?��c\���-�|8f�&D-�C�r�zpg����ChGqQ���Y4(�Ϗ��A��Pħϟ4Eӑ�V�214�{e-�i�Sgp�B]Kt_~��i8,�`�/�=/��ܐ�i����UE6�ʲ�'>��k�6BpY��"G�7Ҹ�J�oS��ڰ^3a�	I5���iQ.���M|�*����9q3^��7�ii�`,\�^|��s�}�7T&�z�,�j��6�v�bĚ��n�o��Ϥ�V�
���3ES�*�%gS��_ߦ?��n�Hk��^�a�8*�A<��jx���>����z�����7N�����c�1|w��g�?W�,��]3�iI�kv��s&�_�9��~؉- ��xϡ���T;/��Ӑ�� �$�ǝbd��V���<�	O�!���<R6S��GP�Pj�M^�bAc|ũ�]%�!�^�On�I~���G��)���1K F��a��A��R���:6EEH���o?�����X�K����U<�l����{�&p�J�IG� :������!��K�j�Aɕ�9ѡ+-C=T���{m����e|���@�F��2�r�\��Gubj4��M)b8-tg�C�/�e~(��]rH[��6#]$'�*#�M�gV�I���s�X*�������+�^JWkm�����=�4WP�L4�Yq|�~m���1��4�U����C�7���&!�����+�L\kp)h������H�|�_%�Miπ�㆒�ã�\�p�`����Ė��
G�J��/x�4���ο�[����2�w�⟕��4�i^�q[h�eq�X���x��58~^��T=	e�tOh�@�C�ng��Η>()y����3O0�Ud���:������e˴h�6��Q8g�Kn.�}�Ic![���p��I��t:�[Ui̱��Eb���[�;���6��� �`^��^�I� �_:v�*��r�'����M����
�p8_��V��wR�Bf��X���h6����Uv��<�,�jP۳j�I��SW]�E2u���Uk^�c�>X�x�ƽ�6�w�d/�z(��f�;�*�3�z����t���n�P������̀��4V&N2H�"q�t�-D$�^����V�y Q�/�jp̢3�}�8ܤ�`�Ι(t'"�b�A5�=Uyм.k6jo�A�[m��0�+p%��=�:��Ԡ�5�a�뫔���W�M��^��&�T�kv���BI���d�K� ��˳�O�)o���)MB��W�';��AYj�u]��.��@-���ށt]S���A�3=Ɔ@���~��c�l�@|~�8QF8dp�_�Ƃ��,�Nq���1� ��\�������9z��39Eǒg��lA�[��M�Ͽ���q�\���XRpj���N���eI<u@�#kj�PA�o诵$�:9�ީiP���tj/�"瓲l����Fr�].]]P[F��4�Ϛ����u��^�f��$/rugP�'^'XԔ���8lp$�B1�}6��3���v
�_70�&��<�r,v.g^MTc�8rdp�5��qe�,7�_X����b���@�l�(�����S+SG.nm��s�F��D|v�K�)�n/4����g��S
�X]�M�j���f����n��hN�9�Vշe�dfT㭗O�cI����J����H[�������Qݔ�]��6��+>�N�}��n��k�d�^�#�;�c��[��cS��$��f�{X,{Uhշz�o��T���H|�����_"=�-F����^�T�3R�,Ъ�>@�	�� �AJ@�� �\В%���� ���݋��� M	���ৗ��g�W���xݾ	�4�õl9y<)^B	=����H�3X�i���@�]\+o��)N�I\/��u`������膚i���j��޽��#���'��d��.Ӿ��KþډSP��Ģ��U�t��-Ɨ�����L��ɲ�F���T���mv %s���� �.P�LU�=y�]C�p�T/4��P�1!�� ���4����w��^�-�_2<f�J�p���&}�e�T��z ,��:��z�m�Z�a��/F����F���x����1�s���k���Ag���gcL1ǉZ�ދ�l^sv�o2�.$���8�5����7=�����Ϛ���Ж�U��H@w �~<.�B��V��͂䉸�\p�:~�.fQyj��O�X���t���o�z� 4�� ���ł&�@����Ʃ�U�-�1g���G�����1��t��F״�'8J>7i>�Qx|$Q�J�K��9�l�PK�0�&Jh��߹�n���Xx.˝Ӵ�&���gE B%
Y[���'2�7o��T�DiR 7U3��J<�����*�uo�'�3��qXj���)2��uv�=�rqW�b��i�X�\	%7����a�����)�˕�YA5<b�?��E>�����0b<�S�ڎ��j�QKYV;Q���(kn��X���9H�.���"�Y��kЯ�A�^2uA�C�W��
��!�f@$U	���$�x��vKY�ػkr8����鑭�<������=�o�T�J�&����u¹6��\�R��f��?��&ʋ�S��^+�pA0Zf��5������R�%��x�+4����2`䥃��&�_�6���<Ź�i�0�_wM9��7 ����b�rOy�����/�)���ܘ�5���sR��Φ��Ά�AԜ��P1,opv!r1����R��0km��(/K#d����=D	�&��&>_l��������xN+�L�|�Y�r����m5�[t`	� ������O?���xt�q�;;�I��~�F܏?�T~��/�V6�>R��|f�EY6�>������t�z��z����u��]�Oݽ�R~�2E����Z ���K�l�Qٰ�I�y�����a`��`�Rv�����:�Y#�9��_5�i>�${*�K���ƽ}�was���s�У�YMމ}�5��lYtߨ=��F��lχ×�V<�Q�=�Z�=�)�@C%L�IQ4?ڇT)�w~{ 2�f��{n.����WM~|q�켴)�_}��͎��jm����\�Γ�TVU���R{�I����2=�7���h2'E�R���eZ'�[6�v���3�K�Y��˩ ��^Ԅ��F��@��P]
����m����`����@ ş#� �n���E�n�3�<�s����vBʥ�ׯ��UZݺT�j����%������=]��>�5dSg���Ɵ��v"����O��H$~���K���#����В�8�E#EUu��@S,�����I�wI��zD�H����<"{��n���K��pannC��Q3�c�/�M��y���쭾E�j���X��書�����FLCJJ\���.�P����l؎F� Cܫ���y�ۉF�s���p9�[���dw��bMN��]��c��T�)(Z���)Y������0�{W�ik�Wһ�"��b׫*��"J�)Ӷ<U֜��d��Q�:�����'��;R{8�%g�s(�&�s{^$�s�^ԁ��:���*_8�{�:�n2sk�!���:���43*d���{-�b&�']���X�Mvz�m�h�.x�4����H'5~�Pە�0��5����}����{�,p�~�1���\/�OU�Sx[��U��#��g�#ɓq�g!p���dMuEq̅����x��q;����q�G�tU��Pz�CR<����m1"2rj��:+�ł\�j�ԩQ����ny���Ƒ�!��:kR��BMI��IVG_��^^�z3��Q��|���1.�_�����.���x�T�Rn�&-����M�B��Ïq��Ui*'b��\�������Q!�K���E�qрE��*Jk���%��c��v�Y��0w�E4y�b&�bU��¸�[�+�긝���E>��2��ܜ��
���2�����:�bFض�NGr�q���M�[$HRD���C�ȣ���q*^1
n�>�ױ),0��~Q����z.�E �L�[g߄Ae3öWz�}N菮��Ҭ iN�a)��ئ:(��AT�J��ƞSF}.%����I��1yY�l��K�(����y���V���g)-�K����>�
'u�w��C<�&�xB%���q�.�M��rC�ի��ȬHx,DC��8=&���M�M���(���2�h�,g�;�⨅��]yI���{�W?蘙F��#2Hsb
�nc�RἚX����|�b�$�D�����������C�E�.�V���#���=C��2h�OԽ�� ��!<s:��wG>�ė#mq~3��%}B5!_�D�tg����7۽��r�4�Q|SD*g��
��3�M��q����ؤ�^"¹P5��L@#�q��y4xv� u]F.����d�.n^���b�1ԩ�{��UB;a��	�U�?���@�G��!�z.<b�~;�i�-�6�L���+���b�{��g:~�#!��	��
w5W+1=�Z�Fg���	!W�K؎�I�����~)�_�zB��t7�3����]�n��Y��>:�X06�/8�Wڇ����TV5���V���&�����Z��'����5�x�F>����K�K��UEt���m �`,r������lH���t٘���G����m��eAj�Q�>S�|�1t���j8���j����t�)qG�I�~ئ^F8���8���15q�(q[U��^|���OS|Ϗ?|�.��xhhP���F�Ψt �O��=�>	F	BD��)���T�Ksh�r�8qt��6���ȧ���6׍�;Rl���8Dҏ�r��` ��A��3�F��ad`H9ǇT��.jJ��>J㔢�t*q�V[�S���a
skH��?��:݄3!A��:��קa�1f�Ӏ���f�gCٜ�72�o�{�{C��n1�b��u��QH�H��b���KNw���x�=6�ջ��h��X�5��64���p8��P��b,%�ʵu˥	�|�yb_��7�QҔ�L��i/>F�"���K��D�2�p�/]U�/I5���U,��l�دړZD���ìt�E����Z�ٻ���#_Z�O����͈ʘ�`�Cm��E�7JD�q ����EG�iΛ-�2��� y�R��[q�Fc�@�uR=%����؜��������7ٻ%m�|���4��#Jp7/��}
(ț��/��P��zu�!����~�����ϱ8!�3���nd��ėc69�=���b�$ҪgU�W�k����!��yC,���)^�ϴ�'�Ց#*��戔��F�l�؆��!���ځ�3^�+�v��xm�˯,�mQ�Ku���xG#r��ԟmOJ�ǡ*iݤq)�E+:�hKn#Ү]W\o�g��dHQ�CD
����.x�0�fv�Z���y*\C#��4'��x���H����	��ރ��#��P�Z�lA����掛 nl4��ب��,�g!w.�=j��|r��כ#����9|t˹��\��+(
(��'s��}�deT<}8"4�%��'7[X5.��E�=f���ڷ]Dj������ x��
�����TzHМt���x��:��]�u�ޘ�-ʓ�t=[��1�Ϯ�1��DǦ*�0��s�QX�چZ�m��Tg7)�4�N�T�+1ψ�o�ݽ�XY�?
���9���p�zѻ\,&,��(��9;1��x���<��B���.��:�$,\$�2Y����hWV�� �1�{&<I�3"�R�A���bӓL��l���wq!��`q*"�HS%~��yI�n�������O�o4����%뒚��G��v��Oc�0���\0XU� ���x�Ւb����#N����@������EG��Tih6n$0U�5�k)����i��#���O[\�ް_��h<�
&�䭶R|	�Z�0�\o׌�L�_f��I#T�	�wӂ�T�"�x�u��m��T�:�v�1P�=a��Ep�Z����V2i�V	�{��q�ZcZ���!]�g�@1i[EY�H�"w}��7�5أb�G��iN�+������D��?y��kg�犏YN�i��T�� �;%�peRم0H�� �"�
���aR��[����c/؈��fK]:	���N���!��~��>����\a4H��M�>���ؔ��,o���w�q)�w0��f�ӆ���Ť�Q�%�b��dt�*n����ES�[� p�,����7�J�{�60,��3=&m.R/�d�Y��e�qY<�kz����F��sMo�0�j����~ۮ�#goVw��0S�}\G\P�8η��� ��"���8�T��w����v�^�������ޒƧ�na@���x�Y����{����=v�yFu�ӡỐ�9c�u���Ң0j��P_6Q�Q��]b~M���4�tC�� �}�1M<p=�=Vj�^��2�ل��4����ޘjG1�v��m�Sk���u�T2��\�������J?0����!�/�ע�T}V���3�~|\%�z5智+4���,T\X�������W�"����JjD>����|0��O�֜�b��ԕhHQ {�N����Jx������0�2���CL�m�4n��9�������$!e��Pm��5@��;�<Wj�S�Vt�6q��QRͲ�wgQ�]�lZ�5��� =+d��<���M���Gn Ec<����Z��#����Y�A�F�rM��Y��jG�k��G�jޫ�k��v��G/Lz��xn��\`�kQ 0C�%Sv���M�U�|����c�9�����F�tϖ^;�0��{Q�lHq�WuW��1��}��Ga�l�ը���B�B�x�b'�(�f�D�U���1��@���c��=����p����+q�9qP^�UtAgY���䗛!����d�^���tO'�;V ��� f�k-�i'`A�P�Z�Y�ON�׈"Ӷ�dc�L�%��=տ�3*�1λ��|�'��ִ̍���R}b�^�]���M-�(��$�m#^/�n���t�r��C`J0Z,L�W&\�)�%��JW�G�A���D���T�P=z�&��!�������W���@�h7��X�
���v/9��������p��|n\�P
#K\w>"R�7谰E3������=�7mBwO-�ȃ�t>���Fy�S!� Z{&C���L�|�齎��i䐨/����"$U�Y����3�����xT�a�?&�� ����-�����^S/��5�@
�5�j�0dt�h�gJ�W�_���j���.w��3K�*����K�+�{�F��8b�V�"7�圆�:
����G����	5Z|u�����g�ܢZ�'�O��]��"�ahF� [�=f搆����#�'Z�o�#-Md�*��G��p��Ӎ
R\?A��iD[9I�$�"��[����eڿ<1��x�c�9�֛��2�BG�nѢ2	��&s1�r�����̋{".�~ࠍ Z�B�̂G%�ՠ�\m5�!g�����g{����4PQ���^&�	��n��{3�k=(�J�ǄoĸDUu�L�R�����#����#a/B7{���^�*�V���-k7�� t)���j�R@��O(�˛�*uI(��hV-MՕQ����2^޹/�;~Wj:�G4l��nv.�������_o�c��X/)1�h�8��`�#��;���3�i+�T��bl��?)����㘱����J�&S��yK�]9v���*�&N*����e�N�A���z��K�}�~�ߜ� #���k�߉��h}��z���m�cP�=����uk�rܲ���>+�5�Q�N'M,�`c�A=�7�훫�̖�5�f�ĝ��V�b��r9Ĺ��FѷT%)��D��[⥶��cj_�8�hY�%�np%��{QO��EE�=����QXt��Ţ>��Ӑ�ct������Ά���T��T�$Rc�{.�B�FA��q��t��
�
q�ٶE<Z~KQ�hL��HF*䉞�k�L��J#�eH�����LV��f��CO�4C��Q��.����M���Q�#GS�
Et��"1�{r����Z��x�"H���,Cڕ���p]
+���Ǜ�����O�6{�4ε�d����N�[R�zeF��T����EE��O4��!�4�����6b!^J5�{5C��#�d��3�̼�������ib&��&�$���_8읱��kD��H����:�6֟&��ʐ�]���=����vkBa�׵Tc�jM˷1i�U�hU����|��b/��Ŏ�-��k��@e*[��u�C]�D�lU='���}Y|Ԗ�?�F�����ڜw�Q�?q��L�vU!�ѠN�4�%�~ȋ��/eh�������v�P�(%��Q�"���h,E�Z�����rtH;����Z|�=���t.>����S!A��.fD�+�*�ָt
�"ƬH�;�Cr*	w�}o���Y���n��
��b�����x��Um͓R�t%�
��%�Ʀ����A����� ��RQ�:[�q�%�r��"+s��q�7�.֪��Z+5B���s�G���Ql��i�^xN"�S~U!�����k�����K�4F4i�gj��;-R}�T�Ņ��։E ffu��;�R�C�_��MF�c5��+�3S�
 �b��� ��%=���\�VS�`�DC����Y�!��Pä!t�9Y��0pVW�����?iY)!�}�����.��J�U-fQ4��۔U�n��v������o��I�����1P��>YOcZ�b��i<��[K��`){�v��/F�g�M	�O^�SGeWi��tGQ�aH���Q몍��P�=��A�k�ۭ�����+e�.+|KIɱ�iQ>׊�0Re8&ٷ���̇�@L���Mek�Z�`�t��&��-�<G��zӺuiR`S�zu��;�J�5Rfij�wu-Ɍ�`����VQ�J�6�5F�����tV��I�Ѻ�Οm)C*i�Pt�����6�!�'�?;��y��ȹ�V�E�OO��<�`�b�"ϕ�ٹ��zLc�%��Nc�[���	~���(�RA�#P���р��0
��A�]��#�^%�la���_O� �o!l�; 6uc�Q���Ɛ�<9AƲ4s���6-��.�(�,�Z\S��RP�>)��
��w���b���?��il����Y��b��hѲ2�4�ջ�S�j��6��\�Pz�=~y	��E�L��=ON�G`��?�@`92�~�tK�����`�n�B�Y�M*=đ�]5�7��t��?�g�rArc�� j�ӚOv����4a(
@o<�3�MK�xȔφ�Y^���|!P��P���f��+���Y����*�⚖���\Y�ݶ��aX%*A<0"I:�5&W#�!�����Nfe윘����HqUl�� �PU����e�d:���#K���h�=��_�vP�ԟ"J<����4Gh��󪢌��E]����A���Ǡ�qr�C����*�qO =�C	����zd 1d�w�a���`M�ym��g��4�د�<�M�K5#�}�in�QI~�I����YMɑ~�|����u�"�	�2fc��*�Lxh�D��*���{�bl?|]=6:��q�}h�#��\�[ո�^7ʘXM�=�Q�huʩ�f�E*�P�KG�?*��ڊ�t�aa��!������Z@��ϐ�i?I��`��|�8�X��\��nP?S��ȸF���W �A��h�y]�9���;�9*�9��.����5���s��^ڝ���g�%��"+���D axb]�:�u%�9�ms�<Ε����KyAҪ\�m�1���)b�[�*\����H��Q��3���kZ�_�L@*���%���*ve]��n�(9y8{�������6�] �n婳�������LS��w��A>FpfH\�(�>���M�1��~�8t���]g�_Y�[��WR��s�#r傒��.t#F��7_l�zqi|O(�mN�bڿgt�jn�ⶸ���0�j~����aL��(`V䏾}e�1\kr��}�(�ef5F��>�K��c�\~j�M{ �XF�ɚT� w�:��U�э�8��~g��{�J��ߏ�8ztd�n�&0y���S؛�ӏ���аYXؠ�A��
P���5��W�gbj���^�*�ö0̡�
��pocCG�ŞC����G����q�/T��zV�b��"�&�T����횿��ƦȢGH~ 7c-n�Ԯ�;1� b��ո!�����P��0Nq���]4I�U����:!�.q�e ԂGd4�W�a��݌�]sJI�5F���&,m�[�����*�Ltw��^(��u����>6]>��O����jjp�J%/v�����*b��BG�fEة�����̏�BT�D��F�,��c��{�"��BX��Rt��1��'���}�'����g�)�jUJF��L��I��6�X���zl�;��?ӽ�� Χg��d&mй�3�-��R���`v��$Ak������,R�^'��撲a�ZI�J7�P,6��wT�
7(�71rz����ܲ��[Kt�`;6�suT��/[�AZKQ
���$��s�7L1X_��u�����C�%r���׬���V
��>�*��c�Ɗ���j@�۟xCq��r�W�kaHQ,�1�Tp�� /O�5�O��x؎���٧K��N2��؀7��]WG��(��Tx�~�r3Bcy���b�ޓ�uM1��:O(�S����9n�rn9�$v��`}��s@�"۝	��]���m���)Y���Q�u"��&(;=�ӯ��R�?���Ջ�>�G������>~��H���5y��ً���5��C�7�o���t���9�����U`��-�~�ɶ۹=�"��r�B]�9ڬxq̈́�u��K��*����9�b`y�8/�/���ð6ƍ���b@⺿/��1�wռu�X��N�u�������'XȄ�.��
�L�(�R+�U�����G�����1��C�Ȕ�N_ �l�H��V�d�s��ZF�#gjT���_1���X��\y�����`6�ǵ��&>��L���b�z�q���%�0��H�lI���3T��|��z�x/e�թAD�Q���K�F���C�[v|CbB�Ȝ8_ø������zT���J���젇�rU��I�"���Շ��,��y�yDF���x�BC:o�eݜ��?!�s�8����0�QRܭ�X3H�����8�I��ݜ�V��T(R��00>�Rۄ�4Y�&�օ�:%e��-����.�B�"�E���g��x�+�Ό�c
��"7�Q틞=c��7G>����ǆ�
cs/E�I�h=^��ub�Զ��DGˊz_U�6Í{���\?z�Ȋ���z�X��Ѩ��|�7���E�'�]F� ���E�0$��������ߌ�*"�W�p�<�:�ѫ.R��,÷��V�d�a���s9~�1�������A#�R��I���!�~��T�MWٛ��ɬv�����Q�n_�^�����+nk5�� ���X.� 3���n� ��Y�2��M�ƇjH��[�x���D�5��'U by�޾(���>z�;F���:�[�r�:"��xzu�ġ*��s��0�l
h0�a�x��ɐ�ۿ�!�.�)RJ�l�!�Ȳ��cbD�l�\�H��Érf�3��,7B q-Ðn絎���g��?+_|�y�h
j�j/���
�������B�Y�]F���34J�'�%ƪf��*U�K�ԭ�)�*�t���:����/�3S�eɓ���*á�uL'آG�͞�񬍓��E�0�[`=�f�a������Fd#���b:H�����A��=�7fƗ���X�ZL�q�H8�/���=7�|O��U814N��Q\�!0��Q�Z�,?��$n\��������,>�1�x�*U�IDj��$�YY�1f�7��k�ݶ��gV� �ŗ�>E����8�O>�����G�E��o��v3���z���j��X��Kc��U4�#r�W��Y;�ʇ�����䨑�TcagEI��Z����V�!7=�ڛ`O�ș��ۈ|����-����.+QY�xވ�^��{�Oh�fZ�M6�8NŤ��0�FąBJ�h�B֢J�{�=�@��@��Zn(O�Ņ4��4Lg�⭳GSD'����M���[���+)�S���#���Z�H�u��WQ�����R}ިU�k��9�wM���b���F�hT�%��{c���������]J�A��Y�1��H1
Og<Τ��b�����6���;hin�m8��#�����y:"m?�}b�*r`سǌԶYv����3p��g\�C�Fj�ZE����&3T"����L��CK�3�4���&�s|I�K{�W�m;�c=B�@�N�(�_Fu��*�kA�l8N�wNѝk�m�s��y�y��~sԐA	;�Z�k#GÛ�H�&����M���������W�����џ�w���wk)���[=�񖩥/�m��!�͈Uf4�����!"N�kR�'�o!���EvD����=͎J��X,��Rq<��j���$2�hIS��0V%��e�.$��Hr��G�ؔ��e͛��Ѱ1,W�*�*��v ZI��s�"�3B
�]y�s�d�9�9�8C	��B_�~U`�G�i�cl�(�D��G`Dq��Aϧ�xWGq���.�,�x�T��X��ɧ�s�8�qG�v�P{ū���ciLh�v]D�ky����f�^�1$q��7�4��;�}T��\#ϧ���1C�x�Z���oN��#Z �hQ�vj��R���!�T:'���W���6�\�H��j\Qz��5�+�R�jV�G0K��O��1��9)��|ּ*�m�yqm���s��l���d�=��b������k�sٰsME!������S2�v���i?���DFu-��7skL�)|kҎ���sW��4�	:�����s�S����;	+��	��:t�K92���Srn���z��nN��^΅�<f�ex�����l{�c�%�v	QL�z���aC�E�E���I����F��-�F��k��쮣)'��������{f^c<����xs�F�w����9f�GFpc_+���E�����(Nݟ8n9",��14��<u�]dl�UY����	!t��ɛ{���,��an`�>�fzmdd�u�J��}n����ê�h�8Ҙ�e9��a�$\v�X;5"�۔�R��
_C�!��0�#����߶�0+bZ3[1��c��tMD�\�S@^�Ͽ�"DU(}	�Q:w8�I�-�����Sߦt�� )��V�Pf�o�%�@%�nQ���Y,��,�T)9;0���1*0��=����E1�5�#)i�tp}�e�QJ:��ݹ%4����t?zAՊ�>2u�Z#�**�)�Ǎ��&�1��'�ψ��A����7^���0}:�811�4%%�ZZ�Zշ�(��K�@Q~:3x���l}T�`��]�e��I��o
%c�#�f����~v��F�Cu6���t���f�ɑ�R�z�A`�6���6-�C���<wG�����~c*����r�Sbp�<Iͽ�F}��j���b.� �A���FʅG@���̭�5$yȪ�}q�Jӭ��M�(V0C�ǖ�]y_8O�z�SgQ��<��iM���~
C���h�Pd��$t3翳��XqlY�N��o��H��f@Sە�&�$�'_�lL[��N���X��U~��b��ߥf���L03�={��J���z�3���,�ͩ	1g�jL�X�^���������oǊ�k���F�%K�l��uf�O��ZϽ�xj��|aR��n�޽�}����e��D�W��,�0!E�6��&���l��Y,��u����p�(��FR!RZ�MF�����!��19�v�'��宖��9h�"#V,��~��NA5j΢L��{�g�u��7C�,�Y̢d��L��9���i͋��Ϟ���)���{�5מ��u�@���-�Aao]k{cF�p����l��_h�Q�¹����y ��C��وn:�L�)72�mhmB�����"�#�PF��5.uMb�\�<!�q/?��siL\�aX�/�q�~�i���(���������$ֶj��2����H�RG�G����#�#�ߌ3^y]��u�P������y��ߨ���#�*F���Q�%u�s-�{�}�Ԭ�"zҔ6b�_t>6O��^��%�k�"�����e���"/���V�r��)Ys� v�~a�Z/���-�]��6�iD]�O���u3/�]t:��=��~�)���J4��.��b1)�`��>%զ����\,1�$:�п�{:�������q-e���Jy�E�ݤ˅��^��{�1�Y��"=HvܰBʛ�^J��מY��+\WU�!�|�ѳ�4��يF^�?�A�X�&$�[U�9?�Ƶ�,�l�V-���R/+�ہ�|+&��.������ǿX_��0�f�pNW:ɘw����������䀻��!��s�n7g?�Ϗ�D��O?��gB�g�kQ��*��.|��>q:eO���!fh!b=�Ё�x�6�*rͭ���5�4��ocr@F�����crfE*�D�6��d��9�2�*�y��MD����c*��.�$�#��]~S#Ns�B��\ǻ���R�*�6~�Aָ�OL�hG�~����F�n�&n8���m�# پ��]ҨN3'�F�R(x�=�ܐ�2�-��Ze�h�fXP#�'��jPCZ#Ҷ�^1=��݅JC����r��P��?چJ�3"�C��t]�X4m��-qQ�1�S'�h��[�4�qqM��s�Q���H�ZU�����e���f�\��-�1�FT��H��l��� �*��?�k�H�v�Uo�ⰻ497X�rϐ�1���e���w)�|I��5��#f	���<k�֢~��#!c[�ٌ�?������#x�����~�*��6�Yت�/��~��7��}�)��M/_���,��������!u	*���k��ǟ�w�}W�����Q�X�0z�#蠞�n���4҆��߶�����_�X��p�@���V�h�t�S�v�sD�f��Ԉ�U��yg�h*drˈ�w	��2�D%��& 2ѹ�k�\I�����CHT?��d-iHT��P`���)���/�e��N��Y��5"e p�ʔ��H�nn-���qF�Ci�O�xV�t�گ�OQۦֈ��W����}������E"�&0�#�R�f�2A�YR��I�Ե���!�G	l��ז�����,U������]��x6���^dbbMA~��co�����-N��e������<�!fZ�ac�Zz�ƫ�=�ړ���;e�x����^~�S��Tٰ���W��%@���	�"F>3btj�����" gʔ�S)�4�q�@Ȇq��_8]Rs���?g���Xޤ��8:��H[]��u��L���L���>R_�aP��q�����w׻r�g?��ry�BS�s�;��9�-d40>��%"ݟ�I�)�JX�X�Q�ߢB�*8(1�繖.W�g�q��������lǉ����I�p��̸�V�u��	p�?#��3�*�l\��9�V�;�����y��T1�4r����*�ߨ���:�aDb���~X�UU��ΐ֌����L[d�����J���e���T���	+1B?"Zl?k�I-�i�l-�AQ�(C3�Ȣj<p$��Lk׵n*�ox�7�HYawʍ!lå���Q�R���Ðj�X�H�7�M^��KP+��s��� �]S%��W"
?�b�'�22�!���X	�R�q%8����I�x�°t`�Zf��R��=�Ǯz��pԽ��,�° E���fHM�	��3���3\+`�A{ꚬ�:Ud
G��/?����O�.�ѝ�h���)`�p�f:6�{E�B�#�hup8D����b���l��L�
cX?�p�A=px�b]!���Sh ��1��_�`ǋpQ��/!��9��c����f�.ځ�����,91���Yu^�`�<���fAA˪���,;B%���?A��+�a%�u�U�9⡝���:vP'�L��Ei���u2�֙0��ua[tpp5[���J8�#��ΠVL�v&��&����D�{`����faV)�]���'1ӎ�)+n<;fYX(Jiz�V2Q�ww���%�<k���0�b��!�ڈ40���!�Ξ=St��~��W�\Шd��y2jTD�p`���R�xđ}�_�׈T��RQ�H{���Fb�ӆ��ōj��y�E��������ѯ1<o<�;ص-�O�<���m�.�K*7yl��$�cS�(���8��-���T0R�~��t�����(j�F��8�2���E3�Uq���}��q5��Xܺ���w��}Q����-��2R;��ݴ���K; ��/?Ә"��:x���kn4ڛaH1�.�^�FJ�0�5
����.i,]d,2�Kp���82�q�j�m�p���pU|�ڜ�U���1����JF�Z?����#8��A�:�T��R�LݳBX|���������o�}U�8��]��.?�+O&��R���K���_����OF��Z�6m��{ѯ�-�j�I`>��!��lW�:Ŕ���*=�O���9�&8��0�B�?��R+�A��"N+�������=��	r,�X��F�R4���J�nr�Z7���n#x�%��6!=e�0�㚴&W���Λ���!+�,M�5��IJ���{<ߧ%`[<).�ϛ1�1x�B���Q�ڼ����Vr����0���)>�BP`F����Fט�L6GKn�L�)�:\�v�i�Ny]�lH-��@i="�(�m�.�	��%��R[$��Au�*�h���Q����J9���6G��u~|G�6���O��l�
��`_��`��W���p�l!6.��9/�)���� 9��A�|iD_�Aǡja�X5�G�����J�5�f��o��ВU�k�ƀ@m�è�]j�1���\�2%G^���0�Uk�����:�f�{L�<1ޙ��ʍ5��|�裭�si���B��-�4��je��-�U��U���z���hχ�����\܋7\]�1�d[��7�*����N,%S|SX\�J�vf�׵')cDM�g�M�ֻ��A_hU_DsQt�墬Us�4��N�ƯN��vE}���N�۹j�wѽtU�8^Հ��_�1�|���~�Ba�1�~�(�U䧼'չ`S�h����9���J�O[Z��8��T�bʉ∧���ZII+%#�Z,�(�c�V 3��u����?㘀��s�Nu�"�I��VӒ����IBK�~��mctw�~o����GQ؁����SFMД�S
� ¾��H��)��8����"K�ɕ��x�?�~��e�)�/�c3�y���'9,Ns�t@�ևJٲ����m���H�$�w<F1k��zn��ґ���,�7�E�Mg�]�e�"jդ�M8�v��<�X�6w��=�F�{q�"�&�49��KNeVl�u�U)UX]ɷ���c�|�f���3une=�iȌ�/�wY;�y��\*N��9���E��B�J�ż�~�<R*pj���9Qqo���YԚ(���<�K ��j��n�Mq�0�仆^L���;��N�Y�+Z����5Ҳ����n�,����٭
[,��8/�qτ! ���E��`R�ƭ�ś�e_df`�4F~0.x�S��f���l�M1=s�Z�N�g8�F�̎�V\��oRg��Pr|�m���嫯��w�r��謺'QY�bK�2���#5v���ǟ�:"B;D;������+�l���o׸Ơ)Eg��Qb�2�^�W�܎�6<�5�o�H������{'>s�b�y�WICj9K��vP�5�?ѣT��ȬG�	�r	︍�t�^unžOYj�� κ�z6�,;�m��,��\�UEw��9�C��;x�?1����C#{p��W>b*��!�!ጦ�վg�k/w�[�Šy��R�ة�D��I�?�"R��x���K��S	�4�98�*���Įޕ�w�aH��T�F�5ʀ{�C�L���L���R͎�I�$4c�meշ�I7@��\J��PĪ�"RG"BD��2e�u=���s�I�H��.��5PG�\q�Q 
8�w~�Rߤ�o<���*���6"��\P�/[�X�
W������(y����YE,��co�kq3:5+��Z���F��5-hK�����P��G+�v,���~�Q�lL���j%�Ћ#RЩ~�"�I]җ/C���?��vD�Q&�|���h5���f��G�3�:��L���,�7����l�uAΙQ�&_8�j!x�>������2�ttPD���3����f��mW��D�9h�_��})����1�n�n6�������mՠ������V�������4ŷ�"~P�㍴+z4���E
��f��wHc��M�~@�4�ۅ�[,E������+�Y��b��[�1�6�JI���*��3�;���������T�D��>D���t!�)��@�S��#T�J�8�kj$�˸�fH��0PQL"��*g��K|W���c�h��-��0r�<�z�v���D��Q��S��Oʖ<�#<p�F�>3Ԕ©<0�S�P�KR{��Y�����f�5����%����(C�� ���\��j���{��Zώ�c���nxꨮ ���|�(�s8\��h�s�~)��[$
c
�j#���sf"2i�,��L*��Q����D
�zU�f1�t8�SJ��]�&Vg��jƌ���cJ(���Ԙ�O��e`q�L�"��`�:/�ǵ��4s�j��⼮Yl��Hv��4V�wz9sVm}/�fI[� wm��Z�j<�:���/��XR?��;.�=tv���;�R�As3Y]E��ZS+hlܭ�@�ń�I�D��#E����m�7
,��UD�ہ^7�c�,�w%SsM�r���%��ԧ��jU��C��4ҁNE��"����-�rH��7�9�"i,BN0��>S�"E���1]�=�ʏ�����I��C���w���6��H����T�z�����!�D��;ҟv��b�K����^<�7�����Kuv2Cٷ+cX����c��l����=����A��}�E���Q��/�^����������B�C*D�hU7�V0����A�
l���'F��b$ƒ�7yDf�x)��5��j\\��RKw�~-�������o���~�`cn>�m2��Q�M�[?me�����r.�=v���"�
��gh�Z���]n����Ұ8ڡe��3�[mh�l�	wM$�ϩ��G� �ZB��7F�uO˭q'S�<�����x^�����.L
鮕Lk���+� 3R|��p˛�g����h2���nz`p1WF_É�U�M��N��C���>f+��؍��M�<��@-`]�����6bGT�"	6��;��b�<��Q(�L�Xo~܊�_.�0�G�I��p�TuĵŦ��OU_O�ާ��sxn+��{ދ�^'�aH�����E�C�f� C)l��oK�6�R*v���&~ٌ���=Ry��CΟ"�|3f�)>��\�^�C�	F�J��V�R���>�~B+���__�����g��_~���l�i���kyP�N�����Z8�s��i�tq����Q��y�����'�.}�2~�1�H�7b�$"s��-;����$�J��~�z���]ُ~�9e#A��q>r��.�k�A^�X��{���<׌�]V��;#�G�y�b�>��{���q�/�;(gj`且�H��aulC�3�'�ߪ�Юf�c�Ac���GF�^�<�򇏮��!m�T̓F�߁�����ɔj�Y��8��V�(�Hznn�E�M��Ж�T�:~׭�����GsgЪ��M~S��g�u������R�"�]X�q�7t��u푯�|8�!!��ל�c��c�'�܁*���b���6)� �,�h#���M�o� ����"�E	�W8��������cEC���ﭰ�o�2WxL	haB�����p�u)�L~��8��@����a/�BY6vB�~��w�~[���W�O?)�~�Iy���a�ax�	��޽[�ea���|�}F���<Ρ�tٮ�� �}\��Q����~��1k�ш�e�k��g�30p�0�)3��bOrD\wz�yJSR�JWS[ޫ}T��u]��M��xL����gqe�9f����F���#�#EVM����(��+�j@0)2���$����2���Ň[#���Dv6��1B�("]��8�/� ��w�A��6Þ���49��|X�%�_��,5����3)˅4��M'�50��EV��"=�Y8�Cj�q��/_��"����Q�!�O=^��f��WE�D��b�g� z�w#�ñA.���X�$����@��i��(Ea��G��ǏH�x`�ww�D�m�RLU~RRlHG`�6<���͸|��7[���f�87<�l��S���rj��ӺVt�C�`H�7SfDh���KtH+z��5�:[��~�ڛ���)���+G憌(��et[W�����z]�w���w�bT�q�P��)�B�n�}'um��9*{&���v��~��wq�Xk��ʛ��d3���pA��������:�)�?k�Fu�ն�5��f��s�����<�$V��,Jj*�
Q�ҽV/�G��Y}6�[��1]<%1�N�!5vV]�!�P�C:�	�۱Z.)��7S,������2�E{��E���Zc�=<�5v�R���� m�q�b%���Э�w]Y�aµ|�0���/cs�Z�
�����n���XtMG_=_\� ���B@e���ZT��ٖjw�B�
����ia o"�������`�KV�=���P� ��[� �!��[c�*j����h���nf ZB�%|~��X�a�tn��g��uI����mH��v�h
��+�(��?ޫ�g�Xa���BV1���F������-��.!�c�m�AYC��*h%e�i�]��>�y�O��6�5���G�ڃ�^p;��G ��h�I�r*x��͈�M���$Ļ��)���{�D4��﴾���F�����~�Eekc����g5�QlSAqgH-�oԁ�ŸٴP�I�a��rf��_��h�05��
���N�u����.j"�)�4�v܃2*g�C_U�n�*p=}��W	�6��k�B�b^��J8��d�P�b��|�\q�t�]kEL[8@V�F�MTZ?w�dH��Qh���jL��K���Un��H]�"�A�1<2>�#. .N��
O\�EUwa$g��2-{T�'g;�E1���56<��04�C�.Q�6I�Q�%��$�E�璚���;E��=;�@��H��=�3E��j�D�|���)SO��;U��E�����Y���l�r���k5����j٬V�_C��믿N��)f�+"�!ϱ�������f�	�)
.��@b��!N�6���3�Ӄ��^Ʃ����q��6"5(�F}�NF��eu���T?�Yѯ�������)Y8�c\?�8kEP2Z�{���HD��}_�Y�yH��Aw�we�h��((�Q��'c���(��p�y�ax�n�����Ѱz��m
#�᎒����U�8**5��Ա�(���A��"��� ϐ��.p]���G�I��x.X��cX�d�0��^GWᯑ���S���30˥�u��J#�iH�$���hC;V#�bOO�S�`�c ��i4ԡx���Յ35)���,n!��W�����}8GUn��E`�
�\���J4�Z��=�|�ߣ�Y�������HU���Ű�Z�-��nu����HK�W�H�7=��a�(�E;�5�|�;F��V��Fv�?/1DMv��%(���?#�}��Щ|�I?� "�
#�s3�������(.�}�
��� pX�#,ցf|Ϥ.�Y�����ҍ��y����6�ǽB;�� �������I r�p����^m�����]F�2�V ��燓�!P�������oU\�(�ir������+�;�)�ݳg���)��fd:�Y���-�]i�&2�g���H�׼?�����'���ܰo��])�}����.�5�y��ٜܺn����v�������kd���;��h���}Z�b6�Z��0*mO���ȥ婢�7�"b�q=̅��I�޽��Z8��g9�x�p6Y��4 �?g�%�i���� GDq`t�s�Ũ�N$TĹ�������0=nț:~�'=�15x�����pA;Q�"�3N���K�<d�psUU􍶘��:���~�N���/���*��Y5�;�bRt�(>�$[䅈�_~+��y�m�g!:��?}Q>�����g��1���]֥D}Rj�i��`oOd8���T��������1�ch/�j���g�ך�~Uƭ�-��Xa�pJ�?�T�9��+D���r��I�0��0���sQ�p�/23���i\$�H�f�[^��	t�g���I�ݵ�Aj�����*���#G��NC��fԦO3C�� F��\(#�@�_����Ogk�2D=��	~��z�7(Ԩs�&ѳ�Z��FN�۱6�Êך/O�{��њj�5rP��]����хQ�.u�@[|�b}M�ۂU[ds�Ŧ����Laj#R����\��'�l�1Ń#%.ۉ�'='7q�۸كZ��%���
�I��c~�ma=f�y��hm߿1=\|`��B$�6�!)S�w�g�釒��{]�3�]�����S���ļ�ۂ�9r��@ŊyJ�uRw�H�U��2��ϊ�%�(�)`L�h���;��k�#�kQ�䩙�[��z��Aq��_�-� <E"�fSM\ģ��p.�-�f+�G$�_D1J{��{�yu�̄�J�8����1��ᜧ[�*X��WC
����}h�C	��}���O~��g�p��)�
0Fo?��PdY���}��8W\�y��^���W�b�A����Ґ&才��ms��������q���u,�-��:���F�BJm�.�?}Z�X
�,K�d�K,eB���>#�Z�b�GQM��i��କ5����P��ݎ%�Rg$'��}�z��U�S�̼w��a�#ڲv��0~a��m���}S�Z��Q���h-�����(�M�u�,
)��=ᵀCa޽���WQ)�ᩔ���mh~k�BZ�Eަ��*g8U9�:���ߞ� Y��o��z�����cl��*gB͹`�b �c�I�2�e���W]CCO����^lIu�����b	xaL�|�ȅ�tv3��������y'�8<�fvJ���a�@��~|>8�0.��>ތ�ˏ^��mE���3qa���,Z�h��[����	r�s�MF&�o焨�$<�x]�_���9����C��W��?DA���p�V���y���KS0�9��rt�}� �gk6�ZgcX�7~g��ؓ��k>�5��)�]�Y���8V	M~x8V=�
��Ұ��͛ ����mw��N��ɤ1)�:��*��0ɦZ�]ک�4'6��9�V9*/[~���������~�X	�>�NrIj�M$|��,�,�1jŐ���Y$lb�=�������:F!6�sQ�t�s�C�*Z� 
7dL+Lqu�:ra�(婎�����(���K��M��Ɉ`�s�.��-��B��IF��鄽�{�ݝ��k�%'g����(61JY����Nf��=��bn>'DIP��1�5*ˈp��ӗ��-�E
jL�aloM��[C
m�P�~�q-o��]Ch1Ez�h����E~����+��4��=�
op�f�P���{�p+rAvS7�\t/A&0n���8����7ߊ�L��~G�y��9��6�|]�؎����p0�_o�	�'84���(,m��NG��<;�j���nǪLt��
�YFq���4�=~j$٬@Z��Oc�7�ǞSe��F���Ŵ�[�Mf�XZ�v֠���<���u�T�5Z��
��p����4Y�Zo�u4�����<q�	�Q���oXF,rd�����Q��nY3nl���!���rj��۝Rt.�~�,�ʂ��V�S���q�47�-A���;ElY��lH1�BF�M)�,2p�MQ&�����_�UR�s2%ޤBQYӐ�cd�~?�B�>QfayQ�ע�nW1��tÈ.�:�+n�2�=�R(��16�5oy-)��+�eE݄�,	*w%ǳx\oܗy�E
�+�NH�q��n����2�6#�oa(����,b�M�Gډ����_��Fq�Π�[$����-`�����9@.�CP]�������F
�����\)����z%�0�?G���m�����o��pR{c�p�,؍ZC5j�I��v{�t`������8o�m��'����"A�)��J� �DjL��x���,kٍ�� �O-CQ�Swvڝ���A�;H�?� v>������
�����0���l|�گ�h{��#[�+V�r��mr��i1�>�5��4��]��1V%q�?2��E���h�Nw$U�NC�	��C�3��8zUF�4cφ���şm[��4KZ��ݲW����93�ѹ4e(�^4QӋ'���d��R䈮�0�3�i��#�,i5�N�Fb?�\E[�<�5�>wW�������$(�k洖�֚��Mx���QR��3u�fα!�s�63"B,�����sbఒ�|�RGp46^p5�Y�*��B
�]�Aw��Et��)����>	�g%/�%]U+*h8Z�w�p�p�	-��Àa�w�H���ϿG���P� �t����w-S�(�)p:�;i>W8ZEWpވ>��~����V�����$� �kP��.ڤ�a.�{�(�F�z�T�u������m��L��~�yD���֠�Y�׮����>8bme'Yp��DO�KN�u�ü�Q���)���l��{R:�1a&�/j;��3�d��vk��$�ڳE�����},jIe��r�����Ol�fs��*V���T��G�	Y���)k/s��#�t�+5��҈f/�M��]�9��"Z�=�O&��5����%c]:�%�e �Ɇ�!�:�a�z<4���E�?�MC:�M>hV���FZ~��bʅ��-��u�%k�e�"�6j�ƈ��Ն�3��W�:U�يo��`ҔX|� �uX����	NsUgg�A�cA��(�=��K�ԙ6��R�k��*T�_}DJ����M�޲��d
\�U��Gr��!:B�;�Y ���y�r��]���{��q���RC���F�H�9��oX@�Z��'|�駟�?��O����ߢ�t�Us:	bՇ4<���0��M��ѭ�k:*C����/��	��}ܯ����q&LP/�����:�<z�˺/X\[�
�O����B=����Zh���d�m�� m��)���UЌu�����p��9M%+܆�ܮ�����Ų�xM�Z_<�&ܼ��l�@��^Ly.�X�=��ir��u��|;� ۜ�zl���`�۸�c�����<��?�K���v�!m�����Βa'А|���W��x���&<܂����.������{����F����Z������Ѩ7�uM���^��~�U���80��B�w]m�6C�����ٳ�R���Jg��Q�gMk(H�̌Z�ʫ�#�͢�+v����w��	�����L���:b/��V��*���:��m��0�䍲�m��A�ĺ�9��Ȣ�҈��3i�D��A��zyK�!:�%�򀽻t��X�)�=��E���_����d�RBT�9��Y��J�����vD�塚c�7��;�5�
�<�� xZgw:��b�W>5��X���u�,^kc�[�=Ũ�f��t�*W%N�/0�9�Y9�B T�$���;��=�u������e���5%�B�`,yE����ȸl4�����:���!�tۂH.�m�^;�����z�If�m�NMqs�:��\U��}�#���R��s|q���������4ྯ��o�Eԡw���w�F�W��h!�A�ޒ'5v�4*�E�u���=��7�s������֙L��Q�NY��8�����C���{��n��D�FZ2v���X���NllG]X4G]2�"�[ve�!QSz��#�80���ֿ��aЂ<�Q���A��W��Ғj�.Ϥ��~"r�{�V֗"��s��|T$���+<8�jt�����)���J���F����8�G�̓]�k�(��>ݢ�?o�(i�}��^��wa����0~�M�]�� �c���"���!����t�m��Y?�:�8\�����~P�����k�߯���b�u�wY�΂ ~8<�#��Τ|o��x�B3�5a
���k�~����%s�f���6M�Wërxq�(޴3\c��j����a� �ܨ�w�/�)ǚ�cp�F�i�U_u��o\�;�t���t^�'F�N��c�L�KkPK�s[2BuJY�����額A.�\��y,@���>�{7��RqJ�\v'G����}��fE�璋��e\��w;.�"�o��I�#l��I�G�1�$���x��O~P�.�M$b��:M��Β���&\ґ9��+#��Ė�%�Q,���%�@�dBZ��Hk��?d���+UJ���/������Q�gn��3��J��iR���/u,�"�x���+��뺃(��6��®S]qn���ۺ�X&�)=��o��-��X5.k�R��$U�A4�;�k^R��m����hG�$�m&���δ�K\WXd����6^�Q�t�#�;Q{l$KW�_����ډF7��c�����/Ű���-�����JZ�
ծ�X���jT�0�g�]M��{�U�>��3��2Z�>,q����C�
�.��d�L��������z�����t�Ր�A$�q�`5��@�<�T?���h5!��!����2�6���J{yA/l� 8͸��\���Vꗁ��Kꔍ��+�FaQ��.�Q�uO3����x
L��Ȗ�\k��U �Ŧ6)��Qo��q{_햺��ޅ��۵�E��G9��~]�R9E?8�����1VZ���@_�D�+�_V�S���T_�y
��@�P���\+�+|\>���0\�Hm@�T��*B�u(��z4���a�W��*����,@K�ߨ�Nv�Q̈�>��s������崻IgV���Q��������va�q��bJà��hi�|��wuV"�_S�
߇H:&�n�8F���(�QU�2�9��fu��a�%��'r��u�m��|.��8L�pc���%N��;�"b�^������!�ac��3�!���g����!u����9rV�3{#��yN��=$;�T.�	�������Ycs���i�;�4�M��vȸ@`���.5��xK�;	h��nS�|�ۅ���Q���%

�4�У?���Qh�5�!�hy���]��H��E1���R�7	O+��)$��<:�����ңN�t���!��`���"B�N�:mOA��0>.�#�ш�ψ������.���?S	݆O��g�}��@�1�:���"��)�!sc�3`\���?�?m�.�� �s�.)MŤ�2h4���ӭ27�V�Ҭs�ݶL��Zz��v%��sD�������
B0�X?�/�T��X;�/0eD����K!%�EL���g�!F:>���17�4	�X�4�m�FF�
�0ϐO;[K��g%����7;砗0~L�����@��3�\��Qo�ڣ>Z���F�������p8�u.ָ>}��X���լ��!��p}�ɾ��CR3tP\�1+9��މ��ة'&���I�k��F��9S�]��U�j z��T��E�9�֌���e4ZJ�6��!����S��r־� ]q)]S�Q�)�_��C`���hVM7��Kc�ܜ�ٺ0�o���~z�������X6���n���n�G%�l(�s�9����)o�jS�C�,�6
aH�������^����w��/�����c��1x�Q~wL�i2���hFx��an/�v0 ��ҿ��/Q�7��s6�7��נ�E���X����mV�,��J9��c�����E�1tn3DW5e���>x�72��H�h��t��i
��gwv���tO}�03=���)~���èk��<Bpb�p��,D���ʑ��Y?"ړWj8���.����E�tI��4��$�<��ru6��P��p����z�b��,b��o�uDCzK�8 ���D�0�_|�����V��gʐ��Y)�1�5l�#8ړ��(K͝��}���Zkt]+�Q3xm������F�������m��ɢ�	�K�T��M�s*�,�R�I�"+U��SϿ.�+��T��:�t
h垵iGe�ʒ��nw�����j�2���]6(�$��k�s�[�5��cG4�݃�t��nt��G��*�3��l��4
ÕS��V�5�s�l�Jc�}t����`��gI���R��5k��tJ���GN�|��]��Gt/�.�s\���8�b��3#�y��mW$�Nɏ�`]w����I�hs�~V�I�>�I��v٭�l��9���]��،(�\K�:���H{U���G߭�r��Q��F�*�I��R�ȹ���q���2�*���Q�t�k~�<F���%�D�;LB$׆v�OoѦlu�U��M�R?L��P��{\��`�����|/�����x�Á��̵�`������ZS�r�ܖ�N���5����K�����\ܡf65��ĪQ�*s�Ͷ�A����=U�{W�z���2�/�]D#v�H`��;t*���86����(�4"�4���ÐD|O���n�]j�L�5�����97?6��U3Ut��)kױ�Pp��ʵ��hI�x��	g���X%�.�N,�����Cj��0��������y��_��fI g�e�TD����e�M�$���9��>Ȉ:�+k��(��MU��Xx�͘[�(Q������?��d&���01��\����ET��k��񘥦��ӳ���h	�H���B;mН����ls��%��^�����k�[:&;W�!�;������b0ju��Xv�'�H��B�!�/�9�4Z�Y�C��]�c�&I\����>�!rV7*�<XTAJ[�E�(P�	L�A��z\<V��^�r��%�B���"�J����F������}$�z�/����x}�ٔ��<�'f�W��N,Θw<q~6�}l^c}�����.�� �jA�'}D�x��VcY|���
�n���ے�tA���0�N�p<���5h�R�xh�ȡ�Lה�s
R�~��0=X�Y�e��v5�_Oݞ�#"SA�1�3?�zJ��#�"�5hvT���T�
�VP|��˟���)�G����?]I���ގ�=9����7#��' ;ߦYƠTgx��(�{�9��
̈��z66�L�ɱ���!ź�J=)�Eݹ��T���,�hk
�;.ˠ숑:>�tj����3��h�����be�WN��H�5��U�9Z�I$�W�M��-D��s}��t5+@&@�F���p۱��}���퉨�ڶ�c����͕\ٵ�$��J����`Q��)��j�'�������y/Z�*#�NbG<W��q��	��l���:���}�e~bH�DX<u��d�[T�>܊Hk�i���̋i���Z���U���	-*��p�"u�y�i{[��'OAcPuӂN��k�J昆����;FFE.刦��07��T�,����{1o�otzϓYw��J<����J�T��˟7X-iAk*����B��,yE���O5��0~'�,J�FcĒW���L.��Q ��B|J��lpd�`)Rj��55�Y��yi*"6d�n(g!�q誂�e�~��(䬔�����rS��k���/��(4���x�~��>5��ˣ�vh)�H�J���Zi)�_��q�Rg;-�0N���A����Zm��1)���k%��q=K�� :O��Yb�oGqa���cmj����y?�7� x�h^��V���t���|&������~�I�v 1]�8�^�*/�]�o�J#M�c�w�������iIE(z��6Ga�S���J��b�(PSMk�|/�Ջ�d,������ǻ.M�3H��s��o}K�H�����~7Ym�ۅ�5m��Q��꠮{E^-�LX��I5t�O}Wv*�2���+�ۧ�C�F��1$�ȁ�pd&�tgʈ�c�1-��NQ����/C�������[�9h(J���/��R�ԩ-���ߡ ��H�_b2'����g����[���uI��}��t
���B�8�����R���v~�y*�c-�hBa3NbuT+�@�NLqCs�l�W�GN%^m��F�W�i�}j��u���i�G7WZ\��Qc��(j}�>>�(�ПP�F�R������U�@���T��p5&\�{.p��~��7G�<֡�x.W�$"�Y�:�1v[����^Ȅ�O-��\[c� �]��s��DDG��U����wh��I�3�Wu�2ݗ`<r1?��;{o3��)�{l�#���w_c=1�J���� ���Na���R��E���蜹v�=&Q�0�Uu��i�q�v8��N�ya�m�g��a��	���d���ت�o:�n���)�?��,�ZT�	w[%ѽԈ
\�"Bx�HQ�q9�8q��a�葑��=�ד�h|����e3WnC#ԝ���Wl�ܾ��K�{B���U��;ӈ_/��hBw���!��ڦ�}x�M�Z���?ǽ�����r�!��*m��yW��k-4F�*�t=#�ܫ]�g��F���/����o�OY`r���͚ɸg�pL0�6�������W�\�`H�V�8�5�M��c纇:���A���Ru�K�'�n�s�{~<O	�$�#����b�0�j<:ʖ[fgf~�8o�e�ƃ�:�ҨK����d�,��eۦۯwV�T����ڐV��ũiQ?��R]<B<fy��������!m�`��_���I����d���$C�����x���HQl�c�8�C�Ԉ��R�|ʈ�T"�.��o���,�h|00�Rv'eٽ{�E�p��4 bV�Ų��A��[��7�V�a%�=���>�C��$�"Z]aV���X>�;�,��97,���r��F|7�5���1��t(��r՛��/2���_�ߏ��ׯ?ۢQV�?�{��-�P���������:��[\꣨��/�3;{Ta�J_E0����Xv/��t�<2{�(V0Cv�dD*#6P� kz������#M^oM
��F�G���x���T�b�S��>!'!����ӑ���Fx�;v�5C�]Ȋ�k(����*ϔ�������%�r�(�6h��*�`g�����2�+��{����ω�{���E<�x]o��_a_��O�y�>��l���^؄�z��R5�35_��PZ	ZM9ǵ���X!�]j.��	|�.��.��P����_D�t�b4��Ԑ�A��!n�u)�Z�A��WsJ�
'2��E.���"��fQՑ�1��9ӳ�b�����y{]Ǌ�e�ےF�8Y{1S��@ ܑN��w]v�DBE!V�ORf*�K�϶��(���H���{n&8%��0ڦ�v��a@`</Ѳ9��"F������4-<}j��p�2��C���[u�C����a�=�x�j�:x�0h:���a���/�����Y���5H�PA5
D九CU�Z�Da	�Q���,)���\��Uųz��N��8vDs8�A?c�H>6v�3W29�i�U���f�L("��"��oa�~F�>�Q��ШRtܭ�S�rJ�!�J:��d���,�u��X�IYՐ�xy!C-�]*��X/�0�p���LH�65�֘�C��M�[2^�	�c��q�ޚ4�m��#��T�="B��O�̟�V�>qU�;��n�,45Xl�*�"]à�����v�Q�\����ESDI�i9M��u Į�j^����?$�}�F��	x9��\TI=t������h��-�<Cp��NB��9�d�ZS�X�w��1d��k�91Ǽ��W���d8��D`lB��x,?x3J:$�5Ƽ��.��t�������bRxg,��#�h�(
E�����QFJ*1�|�V<��9�6��˚�����I[���,)"��c�mH-���榉�}O�:#O��Y���3'<p���ypG�����E��D[lz�qF�iD�px8��3�<�a���9��\�EE��)�O.�\�q��UǱ1	s�1�H������OֆM�J��8����G�A3�I57��&��z4f6��T�6HW�A$��L8{�W��g_����Q��	�RL��~l���ר��JV�N8���ħl*������*,
T���T�rڽL�k��!E�-����!�U<I+��3U�c�=��⁛���"��iG��`�ys7�+pו�ô�Ò����@=�(�b���2�K����T����&Fz,��"b���{��Ҧ��XFW�|�ICz͡y����zS���k[Ȝtz ��D J�z��<RD�5�3�s�t^a�bX�VC���v]����#�<q�0��P�b�[��Ɛ5K�ف�g&��s��'eNYxd���\Ӗ�����������q��-������ÐZ��$��7"Rd;6�7�Z�kK�DT��=�/\�Y�r�юV�f�WE��]�Zz��e�<4$�?F4���4[��ɐ���+�x�~���\c���͠���Q�|\�s�-��pB�CR�'�r���4�Jb�}�tp�@CBQ�Ђ��q<ƽ��5���^��׼v�,m�<"�JSG��Cl8����Gۛ��q$IW �%�<=���?l�ݙn�$�@U�infQ$u�ՃEudFx�����{i��$���sׯ�@�.��COX�Ar��$���_��
��_e�]��ᒅ�n���Yz<4�7qQ���)+	9+�Y/K�TK������7���w7�\��fٞ����Ξ�Ln�1i���b��U��n7ǖu�"�)>#wA&;���-�,_I�6��ⶄU���*f�5A����D�L��=˙��$�����=Đ/�|����4T���ĜA;X�#~~��`�U��盤���c6{ч�TkrKOSU�7_�YpFಡ�?ݱ#�꺇�{fa,%#C���'TP������St���F�B݆ڟ��c�^����U�z�;`�y�*�>�;jOV)���<}!t_[I7��m�:S��r)ל�1Eύ;�ќ4�_���=E�G�O�nz��!���)�{j=�$M�=׫3��z���>��Z�~W�Q��� �ܾ�:7��hwz��^b�ۍ�7�����_�w�k_�t05�:�MF7PO�f��LE"�
�5Q�8V���e�����+��H�E���� [A��<����t�m������Ae?�h@U@�?S�98����N���7�|ZA��K�����cF��Z��p9�[�v���ߐ^�
�t"��zY�Jڧ�$�5�2��1��z��?���R�Q��R�.6̓#��^�
���]�+�/m���;���i�{�Ԗ�kv���k�i-����R�(��Z��,L5��"ؿD�j>/��sՑ�tU�>�A\r����:U(��Kzv٨ժDE�1���}���Z�7���I�K�Nl�jc��^����E9v�]~2ஂ�d_o���W�����ӧAw�(J�8�p��!�Xw'�N:�P��}�n�\Is�Ţ2{:�brp�CԦ�)�Mܳ�Z�c;n���$ǁ/� vƜ�p�I1�VtH���5�&w�	��7����kM�w�I�m�Ѓ���'Q�Vaa�Y������8�YN!��1nJ4�����!J��*�j��+SMR��3A�:�9pyy����K\h˩#��a�ün��G�V�]g�����rw��*��i-R-�n�7�=�X�*�I��i~�7	��Ԟ�#���$M��l����r�F&���.���G l��9��;y��0��2��2j�<�!��%D?���YS]�mv/�=1]�Q�F���h�!8B���鲳`W(�4�B�������S`��^6/d����ŚƵ�e�>O���M*��%�Z�pbhM^��+����sM'98|Y�ĺ�hs4��'��&�=LQ9��^������E�������*ؤ� �� �� �ɥ�z�����1�W��� �v�#f���@���ҐO���^Ģ��V'O+�V��t�m�=���,�tCg��m��!�'�]����h�}���o�Fr��}r��s�|\���L�n8͓�#dCX�������������o�dF����x�;ix`�I���ʎ�������ÿ��K\���F�����-�S��SE:�<{u��B�K�Y��u������I����f-��yR}6v�OќB)�(�uI6�f ?�L�jy�k@�O�!�k�n��-�t�*@{���
��l��a(^=�{h�(G��3#��G��C��3!Cw!�&q@=9-4d�G��$�`H�;���gZ�|f���b�[���f'v����"e*MJ�^//�)@mKd���'�d�]Ng�`f���P{8�rP�
�2�Yn���� ��|B�QS]�T{m'DD�����堄�d��Z��.K�k��	d��fCC������������a�����7��;��%�
�t@E�set� Ȫ��s��|b��'Ɗ�$��������2u��'
�7�)gk�l?&��,r߾��J��&���2��Ϳ�����+����[���-cq	vp�Ml<i��>�R�"�u���wఠ��������3�ƠjQɃ��2��֘ePbp�bb�������g�Pcv}\�f\��F�W݅v�N3PK��S9�j����@Yj��X�Y��7KG�&s� ����#�"me��`bv�57�-�Ɲ�#���yF/�ezA��B��ћ�d78���V9҃^�Ճ�r4���rZ�3C9iZ-Wc��16*J?�ǍƤ�*8õ���(��N�"(���:=��I8 ���/���N.����@�sS�[�o�'b��Ab,�x�ֿ�&#��2�}�z�������C.�6��O|~�����I��#�V�t�}{NћC�z�������Z���0�):��Ԥ���]��\��舲�!�����p�Pu5)����XݽrV�}�:�h�*fCZA�4m.M$[��.�j�xʟ��3Jv_`��κ��<����[��.�BC<&Q��=���:�!�;Jz�zn�0���6:�o��y�vdM�xP&�I�\B�$��؄Ѕl8h����ufP9$��R�9�i��;i�����C|G�(3Y�m-�6��GM� ���L4Up��uks��YF�"�����$J#�~�̏�)�Y(� �\¿I5�)6�Sl�
C�Y@\�p�<������Qaʟ᪬sTv�����A)��Z��)���,8������h�5���BU��7>�ǒX3�*h1�P�8m�u�jz�v�fp�(	F�����O��},���5��{~��h���D'S���uh�P�S��r5�g�E#�d ��{�w�_��!SĎ
��"��	�������
�]��k�X�ȫxn)u:��N����i+JN����sw 'm��Ϧ��]��k��N\\)׆�iV���7+Q�ǣ�ߐ����W��:��Az�vus�k��"�?<�wCI�쩠�r�F�R1G=SL@�;�I��\HY>���-�6�GTL��ׅ	j��\h�D&��T��猍���X/>w%�.�$�H8�ZE�y��K�@�����{��8�{�Μ�>�x�d�^��~�46&Kύf譵YR%����?�Z�&�#���c���E����C�øn޿o��G� ����0I��$([%�8���P�����p>~��(�0����%�7?EC�Sy��w"������_����*�5����~����im�J ߼?>��qGU$���<�Lz�C<�C�0W%#0�	Av�	�Q�9�m{�r��;x_����ϟc�j�	A�f���G9�:I|�����X�
$R�j�1�n���>�}�uP�8т�ҟ>=��xo8�pXұ��`Ҡ�5�0^/�Go���F�^瘘�0a�=�}��碵�S�0��[l4��ju>Mk���l;#�$�MY��ɫ�^�x�ke����w)/��
�8^eñ�z�H:�c�W������Q�i/*M:��@ܳ(-k���I�\b2���K�[��qҌ�׈���Kx�<�^U�����Wf�F�DE��k-���v�1�`M�'c����5؊�u�ȼ �ahW�K�3E͓P����\��#�k=�ѯ��Җ�N99Уt�Jt�\].N�a/��1샑M!���	����Qvɸ.�PT] @�u��X#�{�z*�Ѐ���h����Fc�Âd�x��P�w]8�rg�?b�J�O�M�u���:�����?
Yt����90�y���}P��}��9�i"�5�W�
rm1 �,��@��w����M"�>Ή�r"���������Qd��y��O������9އ\"�o���I��?�(2a������KH?š��A���f�M�����}ܶ1���A��䃄Vnӵ���W��*�i���0���
H�T�����G�`W��+K��k-�/'*�ʦ�#ַ,�R��6f��|������m̮��4x��ã���@�A��b���o�5�}��B����EA���ZCЃ��,���7�v���"B6��g��V��ܗ�0�lQ:z��"�<�΁x�S��t".�.8���� ��6r�,�l�]��s�QS"H�r�� 1�¹�{~�A�v{��e�nI��\@�����MA�Q�]#��ks YB)Q^�xsd�����9>J���q��(��u���T.�1��^�����R����#�b����M��Ƿ���G'��Z(���&���G�VO�J�2h8����>���,?��kc@���[�W�e�	Ki7/���P^V���>V<��L�C�e�0����X~��;�ϟ^i�c����8��m���Ĳs��Ʊ��:����.�~�6�H�>{v�cp"���<$������q\���qd�x\d�q�1�z.ဨ�x���ஜ/MϢ�_G��&Lr�dlg)v����z����3�k���҆��)q�_�?�l���DT���7�+u��&5��.
��6*g�ݾ�#�f����<�Ήz��d�5�i%w�����N��Pl�Aafr����t��M�$(^G��}��F9-��R��jx͛�uIk)
���6i{��)+
�"p�s(���s"��i4�LD�z�Öt"���¨�T��ކ|�U�O1�ݕ8<^� q[.�T�G ��U��׽U��Ɔ��4�X����N�)�2Q�������t���,�oH_?F0����3�&���h3|�h������E�1�V�����Lm���A�]���^"�}]��E �H�P"C �k�Z>��%��g��X�� ��� ZĽ��w�����a����JTS�I�Gq/������1_��ܷ�AΚj�3i�3�8�=JR;��J8M�b�E�Z�k0O��8��tן��9�n�u61�zyu�\��s+��f�����q8a�]�& ��/���@�ʱ�7�dwL�hY;���9W u�� s�I�^��gB*�@ϻ�~e��6YR��J��[42��;N���m8����Y�^4	7�\���frt��D]e�]d]���;/2��"�F1%t�EH�Љ�M��s��{��뚳���`(�_�I�A�ڳK@����|�G�6�ͳ�ЀO���͗�ٳ��N+��*>��W���5����c�|w|�3�!��CK����-$�@�ڢL��A�!X��#3zz<EF4��g���4�YjH�P�6�f�(9�m�p0$pH]`>}
�A����gpoH�zzzZ���Ncઠ�m�ff��4�T��'�7����/�	�ϟ�˻�~����4�2���5������xo;`�ȑ�a��������~(03BFZ�C�����=�@LӞ�ȅ/ܛ�;�Jg]oǚ����t���XC�g���M/Yu(s�D��FjV��X�rTz���l��N�])��X� ��}ߘ�ڀT�'.u_b�����Y�E�1�!�g���Ω����zY���4�N��N�ά׍w��j!fKm�֌��%v������5�Ly����{!2@a�������<����F�]�8���C���qȔH2*���D�.#���.��i���ZF�.�
ϰb�F�L��=�i���D�P���'u�%���E��ڙ3�cgg.bdQ��cr�(,��-���+�	�^��W�ϛT��Ӎ�#�\\�l��fA�9{�Y-�����A�E�?�|Ytd�ȓ� �m��lݪ�!�R��'e��I�O�t�y����Yu�	���&XP{?2Øk7���z�oR'�2c�'���*����h�@D΢vE`����/X�`8s�Pƶ]���s=�������sw�<��9b����[��቗P*�4Fv�l���1֋3y�q�I�
�1&����Ou��� Iȝ�߱6@g{~f�fyʃ���M�̓�b����AL��Ǟ��^z��E�-���vS���+v 㾭�ڴٴ.k�4u�`k��d��Kh7��EV���qm�(�lu�� �L���|��!�N�V�Q�� ��[�@b(�֨֊����7����dvϠe�p�<�;�&�O3������N: N}ʾ�l �K	�r��N8 M�2�cw�����SC�h�$�CM���S��u�v��[���6������{��[�6���f*11�o]�[���
��ѭ�MG��YJ���Q�l�����q�:`��B��48�륈�9�%�?��Oy�c<1�"eL9�t<��f�82�z�`�yB���)�Z�g��Ee����^�
	!-L�I��l����ŭ�E��D�9�f�]�)����׌���L	x9\X�w�38:f���ؤ��I�}/%OYŁrҰAY��O�
��a '
�#x��VѴ��D��!5�?�R�nFl���f��(�W�V]�m3���M!��F��Y}����y�������Z�>�߇��'/ٱ$�TдH�J&9�V�|���G�{���?�[����ԋvc�h[�Y�	ߜ�s΋�bw��47(�����B�˼
nZ��!#m�Ѹ�lt;�c�.Q��L �:�(qv�C�9,��:��Z�0���,��!PY�|���>��q�'g��5�K^h/�b&�e�p�#hE��j £�\�ө��i�.阞Y�2R`y��u�(wH�-
�2R�U-�=~��1I:�T�I4�S<�cp\��x!���ۏ�!�@���~����u\W��m�m�ue���@J��W��{�P1ե	�5���ag���Y�f����˨ό���C���,�d�葝O·�~{e�$�[�7o�i����\]��P���އ%�����mHL;�A�+!���z�`�)��ک罸�@sוR���kC�o�F#;bʟw��U��E�Ӏ5@�^�p}N�Ep(���$V��vB��cÖ�C�����?��A�>��Q�GG���s�w�E�RS�=Pݧ(p~��U�Ө~%-*�g	~t2��������HsZ�� ���)�2+,�1�G���EK�?'U�����]JB&ʏ'l©�"��z��/�v#+�N�(^�R��S;��5H�A.��x����&jZ[r5�f��,Ѕ.��+I��,b� �Mg����B�Sf�=�j�<@Mu�F��4��C
���M4��ؕ�F�3��妃U��ڠ.�m���XJ����pd�H��e�u��H4������5�;XV>3�Q��E�A����kN�W+p�Lԝjg�س��}5c�k�m톅�����@�e�Y�$�֫��^���#56��N�%R��o�@�����;��ٱ���-�b����<j?@����y튣-p�|؅�^�5�SOy"�k���~�K���Z1��l6�@���b\�ӆʠ���7(�gG���g#�i��oc��u�"Et�y $�T6���YV6�"��}��i�D`e�{ٚM*Ŧ��d{S*E�� ն�iVԬbu`��C2e�)�/�S<;��^�Ag�r]���P����@�g ��"��ɩ���Q<�v��)+�D�-��PI�C'�G	��Y{��G���:�2��|zJ򼗨qPܓ���u -f`qz���fxC��K]�J��U���d���ꉁ���Gُ��<���%�r������򗫺��T���$y�t��j��dO�)��vZ���!qH��Uƹ�W�e�IRZ�0��<�	�a�����W�w@Q�۞�d�h��Zn������(�V>q`k�ٍg��9�}���At�x����*���/��Y4������u����Z
��x�rs�Y���͘J:}�VGPA�~�<1��βXG���yNT�@����+��=y�\7�n�
:[��Ak�3��Rf�x(p�eS����Le�S��4t�%q�:�ϸ4�閥�3� ����)�*ŵ��̦��3S���Ag�L�&�����sy>�'8��z�E�b�e��H/1�s8&��2�&g�P��|�@�=?Jo��1��A��x/�J��ׯ�����D�}��9p��Z���)s6�\Γ�>�ߡ�8��r��2����`�x����p=qDl�ęnM&��D�EA���_����ս�oyy�,����Pl�TI�#�)�u�v<��QA<̗gk�.�[���&��L��6�$~�A-�N�E}�T���*�܅M����IX�*F�C��-� ��b��� ���Ӎ��Kǆs&'}�rG�|?��O1���-(��L�?����0���:Q2����tk����w:�}/ޤR(T�vnD�xx�}�H��ٳܳz_{��vF:@����c�M��]���(�}8@:����ܺYT���M��K��"��Yw�/w�tSFjm�^��m��@fO�������x�d!����M0�)2��כ&ep�%/����c��ڙ�Rc�1Y����2�~�����E��w��V�"40�?����X/(��;�ie�a���n|t]fQ�?��~��j������g��T�JT1v�{��拌��Z^8ʫ,ބ�<Ħ1��K����E ��XN�H��Ǣ&!}w�����)����?�/:D.z���� ���ݓub�q��JQw���:X�ڥ�gJ�i��j��JJ1{&�:�O���A��R{��Ą@��k�5�?���m�-��F��"��z�MNc��_Gį��� ��Գ�1gt֔��iW;�E4�Q�ZX�I�-��&뛆�S ڠ(� ��) �E��>7���k�qRZKf���dBD��v�TWf �tƯ���?���1OS�Lv$i|>Kpa������:�gv�դ�@��_��)��U�#����#F�48�\�]��?��l~��H"�^)׆�2���U��1ˍ�zzb@l癱�0�
n���~F����X!��w>H�ً={���{#��b��.&+��h>a�}�v)�SWXx,�.B�A���+���w�0H& 6�����:��P¿}���{+�����uVy���[����8i�b?ZfQA.��:�/�=�/��N9�΁���l:d-�iv����kH|�b�����=�P�g���c���@8�4�[c��]/�t�T��{�԰�ޜod	���"��Tc��=a�[�w�L��ke���� `�58��E�G�����{��ߍ��;$���{7�콦ٝ>�f���&�7�l<�	��}���Cn���\�q�^��o�(`��]���F@�SY� �˸�����b�:0����x�v-��73
�9�<ˣ��%>��A�`AK{e˶���l��%�X�F#p]լ��9�1�[��Y��*�8�j|�Q�hp ��cZX�1,>h�A�f(uC���%Ki�.�+�������� M ��qm0s��?�ԟI4;�^���_�J���b�G�X��9�����}C���������=�c��|&���q�,����I~���di�2kF>iGRײ�B45	~_�`�`��cTdNڢ�dt��f�³|��D�(��/̽n�K�\]
����M�[7Gs���t�t��Vj�/u:r�(��Ȱ���H�{��4�>�f���b��V���%����X�+Q-��I8i�i
��B�����%����X��K�m�>�d3��)�S֪m	6LMׯ�2#�� �U��e��JXx��G��x���
)�|J�Z,wO�M�9��M��6f�4U&��i�A�<vC�Wף��YQ�����Bdիl�䅮�;Q�wkx�[�x�tVĶ�4(��iu�  !��o�������'�4��tV�Gf1X���p�7<��+�;����1��?���as���߄;���V������Z�1=q>~Y��jV���	��93(�}�>Є�
V�8$ı��� (�i�w��k���ӎ�{��)���y��90@`[�ەk��������fN�5)����*�#^/��cr�)����SB6uϲ�������p��"�[��UMKq2��0�4�Q�H�Cp����T�2�#<ΐ�T��CvQ��MUK7��y�X���d�o����/]���>�BAu�%��%�48���ڹ�KzH�/��[�����;��=�[S��}(� e�4��O�ւ	�����5��:�U�)i5�TU�M�pY�7���t�[<����H��S;�M�����}�p�j]���'v1Mb�S���i7�Ry�6��P9�p��"�{��l�
����Q�`�*}~~as�~[�w�8�!nR��s�ĩb�\�ul6H{��_�o�mN�0!:;��q����.D�q���Ø~`���ld��\e4dN��ŦH@C����3�|�D�0�>���Mc�^31n(̝�2���U��V��1(�|z�u"����o7lOE�|oN*M�Zi�b8fO�t�,3�:�V�#yP� ���b�w{���oѕjC�ƌ/g�I�� ^�2�4=�4��	��mKHq���
������^̓�w�y�i��T�Z�����S������_��^�m�:��u��	�ߒ�]37(ğ3�jbx0:�~=!���)J�SLEt9�L�^�i7���o���B���<�a�{�h$��Jadv������ )�>Ȑm9ι���5�N,-��Pv{͸	��	�W�=b荻����x�uEP��`�������X��Մ�?<=
Ҙ3�<�#�,n/����8=��o� �v�q���9�u���hx �GV��v6���J@J6K��-%�kB��9P����i��;��A�J& z_+�u�"�?�߹�<^k���y&�T�7�d�+�v��T�Ǝ��k{��!x3��^�Ǯ8�����s�M~��b
�>�0�K^<�Aέ�g�=o)GB��Ps�|S%E�ʸ��3f��M�/ga�� �aί�F
��8��ޜ�G�i��?�9�{.�X�t�����F�"�ޕ���&�6�Ѷ�7��[�֓����ds�䲰9T2���^¢d�M�2d�����o�����>	�\7I�ֳ�u
9��\Oݦ�o7)3
`'��}vm�Ɨ��V�H�ͅ����nI��x��3�c���k��4'�z6�u ݄)35���ծ�%u)Wa�fT���!���~�v~<�n�U���9����\�߾��Wo*��ש�IXup��L�)����qN�<C9��8W��X��w���9�g�������pQ��nuܷ�@�D���R�z)[M�E8��)�~� ��[��?����� �
�l�1�@�j�M�A��]���̫�#p�~xT�q���mP���U��QJSn�ڕ�^W���;�y�G@��$�}��л�^m��t#�!� [N\��-��)0r%���=ǟO		���R��u�i�U��P#���9��������x|�#m�h�rs�48gt
u��PX�C^,�ͳ��������a'�L$�Q�|�]��L`le���-q�%����d��'d��j��V�F�Ӱ��qk��'H���JQOzK��e��ϧ30wC���A��D�����Y� �i'�5M�����.��\�_��$�6����D;��d��!K�E�����gI�]�^��I��a�������l�8h���x�Ȫ������-y'�k~/�24����X\^��?���O+��>_kC�nV
c6��u�O�q����A�F��J����Y����.G�V�=u�4��|1�
���fp���)���G�u����2{��㯒�NL���ł9��cO�*5ĵ�|��ʰ9�B�o���pH"�l�cvO*��¸���'���Wٞ#p�6�Ȟp��\W��)!�1���C��ڑ��EAT��lp�&�C��v��o�2��mjN͍:Ԡ� /�3G���T�����������a�SK^P���I�.`�
��B��\T2+����LRC�`0�Z�=\�����9N��T��Y��jC<����H�H�ͻ�!�j�l������B�r��tv�;��Ҷe�V��G���T�L���z̊��ޑ	�>P�>�	�\5F��N�̳�~ȞVM\��_/��[���X)��*�7�+�ݕ�˪XνuD������|�߻zp������M��_��څ�W:���Z�`��h0AC �5�����J��vCf���T����8��hm�|_���T�e<���`@FMqh��w�K[��-/%�E:!�RR���:½�=O���?V?C����^[Bk�<��^��1���k���.z9{&�/����u��'��E�ON5AR����C���)O��M�ʕv�1*&"�)x�)�S���IrA��6v���<e��`C��Ħ��ER����s��GM&���"�������fT��R�GׁԓV>4��٢2�U���j@���q���	Xg �U�zu>q��^)U�^�qx�\)��������M�Xg�x���J �Q��]����%V�+Ǜ?��1/	����5�Q(�G6H��i�̌��Db<O�{�Hm��뷪���vS٧��v�@35x�}�V*�t��(?W'���qi�5/T�����+-aH)���a�M6	�{�F���s�NU�o�4`0�kɷ���m�lD2�0މ0�8�,�=k#hE�{ӠΞ��6�����HF��މ�'�t7���pz�d���Ғ��j�1�I
�����v�#����	�������\3Ҍ�y�kǯ�f�f�ܰU����c���B�l�A&N���~�D�CNk�B�`G<jZ
4�.�A=)���h�\q/�Q����(AcE*�]��tgW�c@^�sm0���Jڔ�I�y����G��
��u���USP%��a� �i���J �Ҧԍ�l�p�\M5�7������T�������>׀	�Z��:�)����� o:��>�lF��u��GPb}�"�x�')�b�uW�~�����%a�P��B>D���b7-���.�<�^BԼ���3����%�T��##�J�*���3�|fL�a���A��:.�g������h@���9+����eAZx.POJ`pHU�j���k����M\��㘦�̲.BI>d���}:S����O����d �0A�a]-C��Z��F�����F���O��/m����i�u�a�W��,�\D^H��Dƹ�m�;)�HE�I��i'��<i֜���TP O�Jpv��cg��ݙ�����rn�����kL	3�7v���<�BMĀd���(%he;(&&Z����ߋ�����"�����`s�.2�ۜ�Vˇ~�e���������'MѾ��K��	_��q�T��p�2��iL�P>�RL2��:�����r9�st&�����bdM�����9d�.):����Y����`�!���'w��9��<_4���q՛h�I3��).O�h[��g~��w�	��-e���{���וz��!��k�M8p�^/}�mVڮC߫d�d�(�>zQ׼�|�C��:�ͭ\�Y��<�����uO���S)�7�ЍF�gK��xc�{����s�<����&�&�%l�+� �'wi�O���[�?����W�)�ea�|��9qb#<pAѨ	L6�.��d�[���QB�_,��K�F������Tm�>���X��V*G��m#&��}�_�s�{sF�Ƿ����g���~w�z�&��ޤ9��W�97�)-��O���e2;09�.`�9H�����<j2{4TRJ'�@��^���� ���������wm(��P��@����]2{�}��l;��ْ�p���~�(��!��Nn���� �S��/�l�L8I;7�Y�I�4��O���kD�+zз{6�½ ���5��t��Ra��HKi	'�Ze|�N��Jm��C^j��{�f rd�щ�-Я�q��ٙ~f�Seܰ�h ��!Ý���C��U��A��0/��P�B�:#��=�ŝ�z4������� w���$7�J�u	�@�0��k��Km_�9	��
���;,�n�56����;t���GS#��$죄�x�;� ��5�ۮ�&�ŧ���7k)*@(C��	�HM���ZD��*�X=AUr\�!�go�H�!��W�D���Ec�k9�?��S�6>��s� ���M�|�x(W�KJ���|jp�oU��S�=΋h`�1��������9��+��zaS.������������n�L� �0������*d�󭔦�C+�*=�����M���l4ua�\9�X,g����0ډ�����h>-�~������$�]���<W�H�6���Ī�J�wgہ!����C&�GM�AWT�����\���j�#�}���ة+������:��Ӽ'Q8p_o����[�s�w��N�rruR����|.�8���_�Q���j��o���=/蠓��h�����h�#��{���[�$u��NYbn�#(ޮ�$����0�S.<�#uOM{�t�k�1���2@�d�Ň���X��2S)%
��]����&+5�a��6��,�IB�{e���eOy�q�uH�j�� �q���(����K]\�Y'���yT*�CG����NM�.��7Mm�eQE�םe����A�5��;��>]��=u�k������6����<[e*ᭁ���M��d ��ds�\�q��J\;��Yk5醟le��A&8b� �ö�$�:����+�*a�h���o���2ŗ���~{#�'��Z��v/�N����E-Av���������W�^R[�������u�� RZ{ߔ|�;�z��8�9xQ����	�y��J00�5|�)<�H�rCsJV���V�r���sXPO䚢J=MY�x&�����+����o��m���1���8fM��u�9ȘTo�cU��p�t�~Z��R9�Wv�ŗ+���>|��y`^$4dG1.��r�Ml8�Ү��:���%q*y�|�������o3�Mݓ�6�pc���%�3��ږ:yG�{��lD50�8�Ao��M�좻�`�pZ�Yf���,��9:�ƣZ/(3�Tz�R�8�2��6��Z�|?��f���4���{��{M��� {�	'�L�0��.�T�-vMk��*N������b`َ��nnW� �C�e2�C�����[
߻z�&ݯ(�����4�v17PE�y�Qz� ���p�T�y���= �	�Q��#��w\��"̤F����~gC	2��N-�^���d�v`�Ӄԟ��z�u�V(~����x�������@ho&���Õb���*��6�(�&��c�݅,��aO�7��_<�	���͵�n��vRP�xv7�F�$&H��q��b?�;�dsȪQ�q�/��T	<�عIrNߛk��u�C��W��I��6%��G32c��5�ˇC�qA�G^�恾�A�)&N�v��M��D�B��o��+�,j2!xDV"�l^�,�	�����c����%=��r��NW��uW��fGW7�DʍԛmK�z̸oc�w\o7��ۏjȬ���P`r����:�d�^���� �၁����-;�7�w��Ip23�WZJ�Z�d �@�Z	�83�mIu0h�td�6�ǀ���X�-�l�L\g��@�I��n�����*�b��`��Kj;`;�s��V���nj?|H)-�'��
fPߛcB�R!���	Wv�\�ig� {��d�b���ס��ņ�5�e��&i��]��X̹�FK�G���.�X�.�Ya���MU��*�x���4J��'��Rl�FG���q�8�2�v#�&�� �
��#��{��%D� �̋v s#��1St�Gv��� �-N��t'.Z���{���Z���Y�0�3��v�V�K�%�$�ȗ�E�&���)K�Ȟ��R��.�IN�&�GF�X6 -���*x�q�#��4���9�\���8=u��C�b�YsN��e��n��Z�|�>"[���H*�ҁ��`�����rd!o��fɛ��]��ΰn�9�,Jͬ��kP;�΂�~�m`��56�q���(��U"�eD�ٲf�lZ���!�
��f��������8�v�@��6�U�bL�F�p*��؍�2�i�0�������z`�7%I[⪮ڒ(��]���6m��)���ăx�q}fNW�gӚI�s�bV���[4��� &��|<Q��ja4�+j�Ep]��.�;��zC'�	��/�Ocs�w-�\���tk�v(\$_ܢ��l��[���ݞ%U���lB��Д"{��p(�C��6g�'����R�Kل3�$�ki����ԩ��*(ߺ�J
r���>��˞��`��|�:r��j�˵�N񾆻��ϒ]y�}�yv���0)݃\eP���(*�W�t�4^LӞ���6wWL���ߔE����ݑ=_�{�s���@pg��2��*XUC6���2��1[7�JWED2�뛀m������RU�9��2������D����yL���S��0��nB�$�"vVw|}a�ى���8�aF�q������c^O��H`X�w{)v��{��U�j٫ÃY8��|��;7T[m�]a��׺l��^��`���,���FU���w7��d���M�j[�D�C/w��jjc~&���H·���4eU�K =l�a
�9K�*uv�TS\H]d�}��$�%��A�������PX����|�G���ARFi�믿1��ܕ-
_��G6�B�/��;<�z��&�n�W͋ǍBgz���5G�˅x�Ό�I��f���l��, �K]�D�4��%k�Iޮp:c�}Gs86\?���Y.��>9�g�� Q������A��T�Oy}Z �AqU� �˛�2,�+�6���|Px��z���a�=zH��oӁo;q7�z���nE&>�=��!��6}����	@�;���{k�"4��H���;o\7�Z�c�ӉV y�"�T)��PN��'G��xJi��y�0êe*�{嶎�4wݻ��d 1u�ϓL����fx$�Ьqg����y�:�2�0�xx߳I�tb�1��N�0q��M�U=�{o�-�������Ҿ���l����.d~5?��=%����ӧ���|�M����`GfLM��xS/<f�N����,c5 m��w/�>O�|�P)'	-�RÓ�A?S��=�?���T=y[�^�6�H:K��������@��C�O���g��ncf��"ٓ_�剬wM�u�Y�.)�@����p��=�F01<����"��g�w����m"�&F�<�T�yV�����q�`�����)=��F��e�����4eҍV�=�
O��'��Toj0yw��P3Dp�R�̒���ؠ��8V�	|ѹc�|:�0��XDzqݬM ��Y4}��;�қ�������A3�W�����Ca.�߿�5��#����`������k�9��cI�*$t�j��-k��*�M~��u0ދ'(1����Tŵ������>�_R��+�3A_4�8F5Z��[]��Q�r�8^��:%%�_:�c7��s�̀pK�i^A�9O�S�N0�:n��A���`���8�w�^��w����4�04�y��z��;�7��������C,��, R;��O<�����8~I�7��=�0H`��C�R���i$FH,�Y2n$�AэS�~Cvf��Ւ��&|qxu�DWk�v�H��u�B�X�D�����"��t����R�}��XX"�>Dx�yܪ�gسt�(Rk೓  TևtC,Y ��Kb���	��=O�9���С������x��fu���s�w������ij�7��CND�Z�sl��_#�Q��ȕ�͆.�6���J_E�q��p��V�e?�p�����������@��d9�i8�d���������v��GB!_���y�^�F'�����.�J��t�-�&��H�z0��n��%c����u6NH�D��f|xIz�=w�2�\�8;NFJ���O�A�y�#�Fs��&`�l��e�טj�ƻ��\ڗ?y0]_Se��P<.���2fi~.;��/������eJ�E���4>q��y�Lm��ׄn�P�ڻ2x�T���F�9�k��e3L��6��Y�V�n�k)�4��|�hSX�a`v��'��fv��^�ZQ�P�r� /VKj9j�@��
xa�Cc�~}b_��B�5lC�{�}�M'��l�q'ecK��<�4D`}L��I�Ђ<!�8�%{`�lѳҊu�,p9��G/��m�����T[�2T:�6���݆(���A�BҼS4�	��G%1��ާ�ot���K%,w�IO:]3��ĩ,'��~�k��)� ��Y�[[ ��dG�����1��]@�G6���+��Bc�r�sLY�t0v,��!��l�Ԣl��{ ��6�.�ec�VD��z�O�"�6���e�Q�v����u]��8m���FE��Ѯ���b���7��%6��?���f�VO�U�`ΐ��&K���U�{�������^<�͋���ub�Z�����*��ZvoV��tYFw�אS���"�����j.i��;R|_�y����f�H�3����{ʛ~ϗ@��5}���At5��{P܍\�(���m��jɟ��U�j�?�纃<~d0���40߶����#a�x�%'�ꤔ�i<�ͩ�MSa�kLY��@ځ�׮EY�z��Z�Bb�]�0�,���b�\�(m�w�D.��T���r-V��m�0����MP�%��dbn�Y5Fi=�U<��_:�4
9)��N���lP!�tox :��F\���ǭfל�@�(9���J�{�Pk"klpXw�݄�>AHW9��ő&P�mW'^�Y���2��E ��އ�g�A�a����~��'��u�b��n����������d�5 ͳ�V�u9Ŗ
M��`Piq�i�m����� ��cy���n�yѐExa{�Ėƞ�"=��o2���>��~���{�<y#P�A]�oL�c��6ܼ�,,��r�l����D�:sDF5*&H�&/4b����
�����QS[W�{y<�������.�������
�.�P��½AF
#86�^�Y�����"q���tw��^����ڢ޴�r�@s�՜�:�[�=�J���,)��v[�����Sq�~�m�^Wm�q�!Hڌ�У&��>�<�G���X�t4W��Op����
{��)�y���JR�~ۛ)_48�.��r�\����>r����~���F�����.�����[I��y�lJ�5�~n�ƺ�>�ҽdF�,=���S�Y�k�O�Ij�5\	���_��RS�/Z@_��6x~'�$�z�q�]j)hG�P qf��eZ1׈�]�v�7��g��z��91�d`�����Y_���ḩ?i4nf��n
`�tJBv1���x]u7���%�	۫�Z��%R�.���Ϝ�gad�},���`�Nb�z(cߧ�%��$M,����#�nKR���wZ�������sٴ$Y9	�%��t�c[�um6����o�=�M��n�����`b��J�o�g��Y��7Q�[ı.f���Fl7�5�`C������x�u�]Z�!��}���n��Pu�xK�=�W�L	٘+�^��>��z���F���׍�%��ɍ�v�t.'9�..��z}.KQ�ݒ��,���0�8��O���mm��u,���u4�m��]Y)t(>?��=��YY6���{���{ߙe��Nr�+��a��N��o��c����a ����B7Л�a���jRJh�0*��6z!�s�����@�]�Ɍs`Q}7�w�.(�r�PO�o.�7�Ln�鲲1��5��1[�AR۷�5��Y�����I��FJP{�o��d4����8n%��i*��i8�M��d�x�}���g[,�a�E?ц��?~:�
7vUU�"W�k�ƺع�`��K�A��#ػ,��m�V�#���U���x�X�֔k����K4^;�6�ei��0�Lq��4Ռ�np��������`�����鋽ݭK��?�2�n��*����FS���MN�t��J)Y�sj?)�;8����.A���:�l�((b?0��E�7e��.�{Ů�+�)�#K��^Z3�:�o��&D��Z� �����1�wf��9��� ]c����M��E1��j�o��~�0R��?��΢"$�ZxdV�vG���	��T,8q���� � �R֪1�2_�ų�8j89�js�>ﹸ��\�c)�ŁB�%�2܀h�j3L��$Rl蝍"p�(#H�۶	*`w<4Ew_���ٝ��pm�[�y�r�-5Ե����I�A��"��IM$���.��m_�13�a����=�W�>΢�E����Ȥbn���x�l��a����X�#(tZ�&��⮮ ��"o5���Y�~�ᴵ�otf�\7�V��{��XC��8X���q�c�|������'x�F��9��4	��m����^�9��"�yO\%�r�ޘ����%f�5�"���>�1[�1�$���^P�֜x�qτ�Tq��:������&�ld$`d���SR4�^!�8�J��5�������,-��y�-��Ɖ���\�C��F~�LQ��C6�����T�8����X�We���OK{\dd����b5�[n;"���Ơ,���Sg��V�{�w<�D�Fwt�t�ŵ q�.�
r�H�{��j��&;w�������1���Y�\Yf��=���x�Z��;��߽1���`�L��q����In��q����j����������84(f���������u(�@Τ�E)�f�kT1P��^HG����|��m�}�tࠡ�*އM�B�ے�5,3epۅ���|�Vy�=Ƥ�A<:/�����)�qOZ͞�g���4�!=ծϟ�0C�9> pX�� ��]���/Z���e��w�T�g u�#���ΌY׾C]ۤ��׏C[���{f�Ūe%L3p<����ة)d�a��U�� ��~�jZf�T�_'D[�E�),��)��@s#.+�I��"�:��)�Jʖ����Oү�z��O�O�#j�a��=�`B�i�T��C��8���]�l��r2�������EP�MxF7�]3��2���P�b�p� �o�W��z��]E���Ke̙3�����P��4�����I�(�Q��n��a�ު�5���0�7⠊�e�G	u>O��G$�^��Y
�*�6�Yn���iw�k�E6K��cP��Vv�C	�0���¶��\;f��Ԡ��+�_���C#�1fS)Mkڸ��ۘ�ff���b��HT�l����ˋ3
��UwЍ&�nN4k$ޫ��)\L��JΔ����t��-�X����_�_��L�*�FC�+:)w������Ө�m������$� �hk�u�&h0_�N;1�ܟ�S�&���8s����Q��l�*�£e8 c���/��䜽G��������*�@�������N��?���ฌ��5�jb�:K�6�B$d�)�y[�Ӛl�`� ��.5�*3���z���|*{�\�1%P �Kj����Y4y�@�b~5�۲��zU���|��S��z1U�x�l�;���Y��3~�kT�����?�L�]J4�8�0��c��S6���}�ƴ�K!M�\Śp�$&��+8�q<��)��XR,�ɂ�x<�#�����Z�KS�VL��wU~��b�球��'��vg��(TR������U����{U3�ǒ<� �ע� �j�źC���-�q/O���J�K�Q��%	��x���҇���L]�w�TMD^C���Cl"���zkϞ�_-�m��EW�\���SO1�9�{�S5���)1H�/��s���H;�/�hT��Q-��4H�xWf�8��;C��<��uM�r���*��{�k�5ww��}X�"���_7����bF
�����L�A�B~��L�4ѣ>�HԹ�%6=���g,� =���&��a���EQm,U��������������o�9y��7�*��H����!`GU۱tw��04p�l�1��XG5C�X������4{d��3S���W&�#�"軙�\��I�A��:c*�����:��~�H!����{ٞ���$,9�>��><$��
�
mYӟ$�+�3ҾvT=�y�6�i`��w��g���Z����Q���u���r:8��%:�vj��j���0�:�~#��a|�0�?�89��
�{f9l�ؚ�6�<F�u3�:�L:LjQ\.lB���SVd���Q��\&���40K-�6\��������8�1l<�_��
>�8��G�\�;��	Vx��s���A����T���)�E�&��D�Cq�=&���4��5_��Dl.�LW�c�Wӷ�u����Oi`4��'�ZS�ƶ
̙Z�)�.�J�vL�8E��uSe�	1���R�˒~;7)�{��٥q�{��eP��2'q&���� �\�!�B�?;f6��^�]�0D��{�%�rH��bsS�c��f��v��F�xʳ��x,�EM�Mx˷�n�I
��p�8�4a�o�%�+�VPM��~��U������s\Y�C�זj2�3ՋzUfm8�}byZ�%u���XY��(P{{l�o�ynW+�|so��ڱ�pI��nb�	��D��u^8=,��~)��?`pN���^]�꜑�0�J�.��w��4$�M��ʌ���l
m}�T��A�%��8wދ��\�=����s�HLʣ)e]��|*�z����/]l^�W��w|P^1KHN�̲S<S���5�D&+���}E&�U8H��.Nfϡ���^<:��/Һ :�R�}��s�4&Cv��8ɞ5�����FJ���&><>�WC�s��B0����bP��g����|֩�$���-` 7̐eq<q�fu(���b6ҩ�>�۷���K�/ov
R���į�̑Fg>L���h\�.H#q��,8�T~<�P�D�1�w��B��^?�N��G)�����!��՘%��~3�!���Q��t��,�ƪnn�Q����lf���[s<дQ����4]}��@��{���Swl�4�]�hSh8\R�������/����5�Oݡ<�k�2K�.�H������:u�����qF�n.1��j7Z{�T���k�(��Ln�3��:����h(šmp;����]L����D�'�e��\�ʬ�2m�V,ٵ�5�3_�v4��/Pq��<>�vG�N�{8	.�T��3EE��M�����I��Uf���R+8���O��|]�57Rq9"ƅ����M��ᕒMw���f�M�5�N�^��_d�k<'���e�AC�Hʇ�L�V&lƀrBm��������o��x?�I���(�_4��(���Ǹy��L�N�9Vo�����~�&�îN�k�N&~��}`q��{t����|>��D	C,`�:��;�3%��-b �p.tۙ��y[xx"P�>~���͝]��p��,��"�lU\�muG����RI]zc�^��;o�N�oɡ���X�,����`G��jJ8|� ����9��`wOAў�&��M*����"վ�1Q����(׃�8W[��	y� ���4p���u5[����m<�,�����ǚ��<Q�;Jz$A:����^��3QO�U!�[|&���?�{
���X�3J�d �U@����U��/^�E��F%�I�m�t+6x����<�bO��S-�s �:������.���y�\�F݋@���Wݤ8�F�����^"��=ǉ5�V���`11�61[>�	����4�v���莯�L�YdW��s��@�`l����IZFD���O?�F��!��Qc>/��-��d�|/Cn�4�Y��~�����ު�%����ܹk��\��qAꘗk�wy�����g���&���҈�p�]�l&=�u~��ww��Xxϟ_��ʒL��G0���4o^	��4a�1\��c/Z�R���@�I�m����2�ڏc�p�l$z�����*�<��zS�c��Z�ۥ��*c��x�6+�VA�������]$Ɉ@�je��?�������a�#��`s�Hc4T�b�`P�vK��h��p����b0��A�cŲ�<�C�g ��tw�*�E'Vk5Y脥\`��N�H{�S$?�����P�G#�����u�Mw��#㉅v�/r���x}>��)�$/;Ħ}
a��nJ��41�ߋ�5�:;��\��6!/���k擟��]v����$^7�K�k`Gp�^K�����ī#�w�|��z�f�<��4��Q� ����t�h��K������뱝�mv-����O�[����J\֦j�qe�W4��=*Ni|����M4?�L\t� �F@�S7EM+��]�=1-"?+�>p( ��V)�h`��|d"��-��t��p�������/�^nV����R�<�r���3�I���cv����3T�f�f�jj��7��/9�K	5�ㄱ��i�~cd�t9?�5:��=S�� ���ˍ����=�b��"���3��$���)�l/:�)KM�w��6�*��hś�W�E������q�����̊�a��GPK1\K��j������+���@�%���}��ŮP��*l�,SG��_o�rT��xFO&�e�k>M1�������$#���x� ��irK�i��:%ǉ��(P��"�E%,�=�ׯ"�~���du�w��<ܝ����b}�^�=�$���SU���yQ��w�¡�����Yt^k��@ng�O�n�K����b���/�������)V�F�h�L�wqm>?��L�A{�e�����:4��P_v�/a���f�����b����?|�X~����M�>~�ݻ��������ԍ��I��0+T����fyX3̞�U
�T���3���� �羞�0Y֪��9��ɐe�fծ!�	�6�|���6��ж��u*N6�cIK��hhk9�8��ם��Ǌm,�m�R1�AnM3��A�C�K�D��&���?8c͇��]M=⒬�����@	�`�z�����j��n�k��]V"���f�.7N�����t�(گ���[�H�.fu�\n�}�&�������}w�~3���W`�_�H��\7�Y�y�����7�6���pKqx@�V �}�"�	"v�)Ze���?�x��=.�X;�Y��f�r��b4/�����U��:�[u�Blq]YNL����{PHƪN�tO �}��G����^T,ݰ������{+����C`ԁ�{P���_5�>e��f|�;�Ί��)u��Ty�����ٷ5��@zd�0WQjdT�����H;������������im�~����M�.YC�����u� H��<-t��#,��{�UN�!��ou�o�N��h���i�b���>Ӂ0��>��-Hd�X���!4�σCy��Yk�r����#�Z!��ּ�4�S�&�c�{�;@���е������T�gK��JtTbx���ɒ*�e�����!�%��鳚���,v�;���𹑑6��w���j@�Y�j��*��V��d���d�۹��EЯ׎����%��7ގU�\,_�)xG�4T�A�>nH`:��J3h�Ϙe��\�I�_n)p�S���Ţzg��N����͘�x`մ�EC���q!g�����h����A��c|d.�kӠ��*�̚f��)-�ۙ4�ٓ#����st!�e�O��0� j"�KņS��7����E�Π����7e�j;�כ�0�#F���&b�!���:�p8+����O�M��B+��[�+{M��L�Q%�u6���7a}��53�,\ra�2yS!w��w�d��b���n�Q�_��u��3�롯���A+�Ը��=��6�L�z��H�7���-L\��~��OA�rύΩ2c̃��\���-t~��[�?/�����o�u&�	���[l�t�〴ݲ>ST/C�D��rvܰM�D��K��)~���ߧީ!��ڬ�_�Y��?�?�ROC;�������\�a�M�\���_���ߊr�.�Gi��-F�8U�;՛���E�8&K�Y�)T�i�{�4Yƾ���Y3髀j�B`�s��j����bsX����#��\���΢�+�'?�^�s�DVWH�Y�׷W��:Z Aw���������:�Nm��44S�-� A��ry.z�@��;�����AX� �|<G�*m+�/I���Olq�o�5��G�H�$[�tvsD��_^r�r���+��@AZ�����#X<P(�Q��i'�)�����kN��{v��(s!\.�6��(�ͱE&�������ǉ���ʦ�y�4L���G5�o+"j\��CC�V;���5|��������{}�+i��l��I�ޒ-�k ̡e�~/x�%`�G*�������p��u)ֲkBM�/���Z9��!��:ߥ����YK�R�������S�'��`�E(�pl~uƸ菛���H�!�C�t�}W��V,6�	3��C ���}�(�n�ΕH���S�ʓ�;ǒ�sFQ�_�W�Y��Sd��B��'2�����Y�Ƞ_xn�8�K�4섿RG��3�5_�y�1�����T)����ܫ0�-��Q`�L�]�{4�.���{� $0�@���>x���-:�8Hx �
�]ⵝ�����j��cp��{�F���:!(,1Yrk2�i/�~<B:�&�?��Lenǒי݉�Q��+�:>��Ǻ<S�
%-9��<��Fut��Ŋ�K�+)Kl���GY��\NҫJ��'�Z�����6:��ߢ{�2v�s�b��L��B��3��W6�S�����T�z��B��%1��]���oB�B��h ��U��YuH-�_��A,?�uͪ����#��`m�:%XǨ�e�?�k�av	Z�q�n�Y�-N��um���{g�O]�GbD�AH�:c��L-e���%���FP�A��`Zt����N �X-|"n�yDc*R�wC�$���q�r���t��i��R��*6���cMч>?e�N�Ys�z�jW�MS;�^�!.g5�c�ח� 4	cG���M�1��wlڟ�����\��	����Q�?����5n0��#���^���������x�Re�|�y�y�r��1��L�^7/l�km֔�YX~m
���kԶi
��pP��&�*J�-�[�[�a��(S�*V\�k�Ӧb �
�>Ȃ�#CD��z�{�R�e��t4�ǲT�Xf6+gޓ���F�2��&�w�ѿ�\M�'T?�Wa>k��P��8כ�� "2ʸ��!���[y\�L��5�����.�� �X����/�� @��<q>}��;��y����jθ�5,��Z�������'/)g��U:�U���WF ��51@���z��$���{O7}	�v���KQ��}ի�M���'���_v��&.��6"�;2����K�z�jHO�N7'\h2n{�\x]N��TZ4�ƒ�6����6�`�gF�f�ϱx�i�#�^@����w�蘃���������#�{��mQ�4�>k>_0 ���L'�h��
���V,��	���D��F_����/�����?�Y~����`�=��?�9���v��>=��S��'��15������q.��m� ���g~����#3#����SN{%�c��5c�|�8�V��ٷ'6�T������c�`�?�)��*m�����r�疘K̇{|�{�s�R��p=p�����5��~�k���1��!��1��u���G's�z�*�8��N~��yM����X�ޣ���x_�sֆ�PvN%�q\;`�ͬ;˫H|-d���(����",�A�m���X�s��0����s~x�U�b�0l���jm\V]԰�^m\ԍ��o=���Wu)�=�E��)�kIa�
Z�M�":]ca�1:K��w��+�Y��]bq�@�8�:�<�izƆ0�Z�I�� :�I�E��|��<�aO�; ($�������w��(������~*���=���'6,��	�����X0�$��.V����m+vR�B$���)�'��}� ��SN�,3�g�od$��Ս�,�v�Ɠr�׭�T��w�E�~QG]%����8��%�0|&���uu*�J�溘)��˫J�؈�:M�T1׮#��VEur�v�|^�*a�%�㯏�5���]mg���zg�7�0Q�&_�=X���9�C: bMvv��P_2�zϱ�G7�+8�
 �f�m�cf��6�0�`�瑱��q�r�%k�����,�G�9���	���d�:*���4�Y�R^����@m�'�}��H_4�*��h��-rͪY��٬<�[���G�ϛK�7�פ����ڶ{op�ٵ��������E���KM<�P��p��7x�:�jw���8�E�-*]��H��9�l��cࡲpF@���I�S�_�I�ۿ�[|v4���U�7�A����l������_��n��7�|�Iq\����*5ԣ�~����������8'�u���fH��>��1ex�)��x���ه̢Ln��R�R��^>�����葝]��.�*M�n"��P�E������\^OY��A"+����|���h~%S���f��M8+�[�y�y�~�,iLݴ��%;����!�4E`	]TK���!<=N���������R�U��9|T6K�b�!59�m�
Ǭ�|Q)��e- ��^K:y*�wי�!����n��Gwj���((�r�Y��Gr���4Y%J&���%|?T����k��k�VA4��ac-1��WϲR���X5��A�3��Wm�1�Z�2����m��X.r��D���{�*,;ݸ��z\o≙I���ԓ���	��H�u�B"S�s-j@�ۺ$%���Y��ɹ,W�@I+�^��eO���-�~�:W�L��?&@~,�!��OG�_O�I�S��eׂ�$�˯���z�R8�۬Idſ��ׇ���)/R�)��u���E�bdsX��6�lU܇^gH�	�����P�A��� �&`�cs�@C�<�'�e��[�e�������>:�H�g��;�V2�i�հ7�����(�c|��msbvQv��+mQn�1U�r��R�u�=��iu-~2�E��>�����*�	x�ڕSfq�����:p�جQQT���,!kU����+=_s��0���^��L�x��.�A	j݄�>����ۮƝ��zQ��|~���u��)�>�D�K�D|Vi�>\����6X��wod���"#�Z��S����7pxM �|�7^�_UFT;����n�]�f�V7&O�V=]1(`�������M��h[Qt��񧼁 ��OkRglMRDU�RR
<�_ڑ#���q��'�<t
8�@�s	������w�>=�����G���"�������|�m�w2=z�o�MB �t�*S�G�ʇ�<��c���ߒ��@Z�G��\޽{_>��$�G��i<EP\%��MP�(�3`�.0p-�Hp�L��awq��~���-��s< k
!���%���d�wg  ��IDAT_Ш�k�i�C.R]�.��;�lz��h���Buy~V|����$�Fx]��n�k�O?�����=:�/���3\ҳ�=��Y�\�!�[��ά�P�(��KK=~(Q����߹���z"=�1���0���ܪ�3G:HW���cu�p_��K@�[�Y��&��>���e���>��E�'��vi��({�69��I�ڌ�]XzR'������W��(�  ̚�i�vDddՀ��j��bLw������ps:����Y��� ��f�2�+k��JX�)��1\�3��,�*?�2��Z�f�TÿSPe{�1��l-Q5��jZ���ؗ�h��X#m�W���r9\����0Ͼ� j�wY�ه��:����0��[+��>)aF�R�mB��5�����������4�ꥩu�B�*U��A��E��5�u���纋s��Lӕ!,�ACz�ѷQ�qS���;^#i�a�r�=i8�U��Oz��^��m^�i3���X~��O<����Z9�E(:�h�u�y[��s��AOCva�7�s����<4�`8aDϸV��@}?�S����VZ߮��d^�,GT�l���p |�w!t�X.�F�N[�S�!�Nk\cqw���z����r`l�Ez�<�qhO�~*��	���׏���}�~R<8y�cb�P�ق�Z���8�������B�J��'\es|x�[�aq�t�O�����i`�-Q��4��;"B����ҁ��o9�5��j5j}�_$�D/3�c��㐑�_O��3�x0_�	5��'z�{J/V}ZG�UF��Hv):�0/�P��5��%
M.����
k�v���ѻM�|�v�c�pbWic���ڈ<�RJ[�����k��T�Jb��s#��~5|��TW|��M��V���^�C˚a��l���l,�r\�a !����Q�=��hk��U�8D9�)�X	Pm|]��w���1D/���^
������=1Ϸo��t��mhѪ�Hp��P-ߞ�c>��:�����"�.��w�6�?]�A;�Y��<G@҇Ioj`V��c���Z������eh����B��N�ϛ�ɀ�n^��ݳm��J�ghO�B�쐾8L��Z(s@C��)}|������z���=Z��3�(�%X]CK�D�7�J��q��c����WZ�{3͵����[�8�-��l(ׂw��Wm�L���1�R#C�D�>z"]m����bRtQ�����$��m�
>"�a'�sG�.i_���޴Ϋ�s�!�]s,эb-�T6�qA��N�sF[�5j05R	�d�d����ݜ�Z�/�&�%����B��*B�X��`!�~��ۇ�Q?������V�|K����0���k>МŲ��,���O�&Bf�Ui <S�<3A�]`o}��d!��N@R���秒���l��0wiۂ���]ވ�"����NŜQ����@��Bch�V~��c�05�?��c��!��u�>�� ��Kr�3���"Qu(u��k�������"N���,�{�|����e�Ӌ�gHTUR8�/�Abm8�'?��>�������F���� RQ�F�eh�띥����-�q�����1�H Y���мL�Ơ�*=ku�x���R\A�{9��ɋ�flL�U�S�J�D�Ё��""gЪ��=��9�E'o��}
# ��һ<�XsH���P:Jr�D�W�ċ��&S��0�bոw�k�o���� e��5��|�1ͬN��	%+�1j؏�j�.�^�B���je����2����߂M#��K�}�u��X�<�-@�^\�U��<s��:���G`���u���ΐ��o�]��9	�-V��U�W�`۰�4�,5NƩ��>K!�@�z3 ���kp!�Pp�.��ʎ^��ɖ�����^℣!1[�T��8t90�9�$s�p����}L�;^#���=�z��X��E��pX����T�Z��=��gR���HZ��zp�:P��%�3d>��8~�ˌ���駔;��O+g�s[��q��Z&�c_�yh"Q��`/ң�$��$�7o�D;�}(��~Bj�mi;���)g�un5vG����i���lr�Q��JUw�-�K������T�ϓG����a]�tVc�9�aHo�9���Rn2$݂F=�������z�\S	�]�~%#���l�51m7�62]�5L��Y�o�#"��䪟V�6�<ٖH�{t��v�k=���9.	�<0Bs��0Ta��Nh�����H�9��<C��#X��cZ���ђ<�4��Sf)Z�4CY-p�Y�tu��3�Ԧ�72�R��J��cyh"Xl0��lt
!]���;"�K���a��Pa�G
�pa�O�S
�ڐ�#%x����ft�G���P�ϫ��t��8����d��Io�Y�J[�15+��6����Ɇ�;�#���D�
Fߏ��_ߔ7o�2a�k���4�ǌK�1���%؍ ����m��u[�2�&ч�o �_��h�������},o߼�C6��_hH�وZ�׉�%��9J���==���p�ҵv4�E8��KB<(w]�g�7r4��X)j�H�X�S�L,ѻjI߅��^Y�`R��.E�/瞆\s������c�j�lޯ�����lc���в�Y�Sb�ɛ�^(�[��|��L#��(���e�/p�.���ե��G���ɋ�6b%�Ĳ�����Y�����^,��AY��d^G����0�kӮyA�������i�K�d�q��\ȇ�acʠB4�bPV��rs:UHL_B��2G5ԅߤS���N�X�㶧��>E�׳3ͧk��⠰Z}��k{MUa�q�|��ey��=�(`���N%�%C�2_�w�Sx�"�[)~�ČX�
+�!�œ�g��-<TP��0l� سRk�-v��P�]�N�����w$�[�B�5�Z#�Φ��Q�Ϻw�QBwme��~L~�zA�R�MxV+6QKF�Tq�\a24���Kf��L���\Yk�li������v�MIl���G���碽Ū*�l�]�2K�W�J����&i-�O�Y[o_� P������2��~��Wrc�>�hZ��f�@��u=G��!:q��2�K*�m��V��8e�9z�9Z��}.#�{*���n���՞Xr�S�ut΢����)�I�D��%W��d�&1�J�xw�8��i9tŦ�ʘڀ������#�Va��c��`+e�@�~a��XG�9#�z����_�b�Ν3�V��������8+i���5�-��	(����Wϑf�Z�8
��&�o���^���k��I���9���	�����<D4?1�r�b�GXD��jD�4K�ɺ�,��G8)���}� �Ђ(K[�1�7 ����>�p��=��҉B/'~��ç ��)����(�}��q���Ko%ޡ���a0���A��yd�(��\EW,Z3���2lK�Z������ e(��_l��B7�eSC?q��]���(t^�w��&ץv�mK�f��s���z��2�䎒��(����224�e�K6����x�+�B�e���wFJ��j��y�l
�3��*N�/��c�����_��^�#�C���~`/��p�z:?Fbv��}n����Y%����1���^���RNY�4�W�ZHs�G�~-��ڂ�����w�k�zg��2v�c�,<�-�<���u�P+:G	aU3W�UI��9n0���C���[m��-��Id�1���F�L�,V#-I�͕&�F����ҔJf�?�-���S�y���'d�6�MY����J��)/��1q��<��"�ڦ9����2��õ�:d����)�t��/E���.�%��j� �~Qo�%��0C�*ŉ��g�O4��Q��6�{�٨����b-Xm�>1�5� L}�ف/$pQ%E��i���u!�:�1����{��C�!z_ݤ'���?(*�tű��A�	��H��OJP���3vAV��p>��ċ��LSRo�uY������g\[󐌔L"��B[w��{�@?	ۭ�p^B ���ST=�`��"�ɸN1vMx�59���H�������c��A����q�>f�11�$�*���w'��ݗ�f���	���k�n�Ҙ.���&���1�+�������V׶��������͘�O�XXy3(	�N�U�xj2�F/�Tu�2ɄL��+uc%�a��Y���BV�KϠ��������^<	u.��O�՘�JC��� އ��H��O�$��һYU6���ƶe�|\zf��J���h2꩘<����̔��W؏��z�U�بv���۵�����_)��.�pUתr���W�~�p�*�[��Mܖ�z�,Xm�iB��nf�)`�ǺR5L!�(O�!�|,�~[�ʱX]n��D��P�%��mMFAS�_�\�ɳns�H����� ��:/E�B�5��]�$7$���X��~�]a���K'�(V��q�A
���)J)MΗ�V�K��61�6��S���5�3�4T�
Y�^Eg�r��l�2WHep �8o�K<��a�pЁ�W�V
&�Ǯ��~��ג�y����ʈ���<��_gHWc�/M�a1f�k�}Ye>|�P�qs�ͅe�
"���m����)Ú9�jN����pg�%���dh�W5o�"�X��0Rߍš�z_�*.��<�VR��+���m�z<��!�fL�	�gS�}��������%z��ɝ�4PVvghop>�t1D/r4�rz�,�;Ѹ"q��%GQ��cSx��3��k�9�җ:LNJ`�o��>&<��1�wl8�e����݇��um��㰁��K(��=����]�]���Ŀ�mRoe�=Œ��2�1�u1����ܖ�} >-�O����B��2�X��	�G����f4���6��6������u:uU�:�3�w?��������ݽ�O�At�ct��Eb�@x|�]i%��t�:���h���&~�;sn-�]?F��4�5ۺ��U@�@��h��>�wR��ۮk���h 9F�1E����!�
ߏ������S�tLΨ���^P��<m7��	�LU{ DŘ�ܜV�4���H?��E#��;l�nh=G}��!���z�5Sr�������o<)wͬnu^~���o�-����l<$%�ݹ�5���K����tzg.�.�� q��Ȉ��3'�NLюRHc�'�������Ǣr�fեx
=�aȓ��0)S�Ds������C.����4���V�tzJ���ȭP���!^Jk��Q����횝�Ŝ�۪9��LE�#��=��f9�}��x��d�qm5���{yՀP�]0�7���f��4�ZIj�'�X����������0�}]oݪ���9�c�}΢"oF�qC@ᕺ�����1m�H�V_޼���ٌ!k`0n��
{�R�O���J"�'��a2֭\T�|z�QX#�n��*��O�mU��rr�
��j�:���8��t,�џY<Ğ����X����r�2憮���8���@LP1!*�ҺZ���!mK���X#������1mCb..A�������s����B�l����1�p",����ɫ_w�4�����H�x����ρޝ) ���ՙ�IτiO<����u��K,�p�b�t�ߎ�CPO��f��S�2�2��Gڐ^.ǀ'f^g�
���.Vx����2,!Q�h���Ю�f�(2��G?| ������c�4����V��w"��:�yyBw3=���]������:��q,q��Zg�G�''�PFr�9���2W^0��݌�{��kߪ<�	��sz,b���2rAU�A2��e�����X�sr�}����gS7>w�H�<Re��������`�Ix���421���n0"Ps�o|�Bmp�=m��Q�MJ=b�݇�����1�w�w�R�P��
J�j��Y~��Hh��+x�������( �/��yI�W��԰6�H�?�5��[�<���������mmC��8�ܒƆT��!���>l��{���'a���Q�Lkn[�l�I��������z�w��29cL��t��S��n�����1m�Yu��5�n���zV���k�DM�YKm�����`eǝ�L���qc��n�M���w�0sU�,G�ml���8_js/���9jȷ�eس�jj�[��P��+=OʥV���~�S�G]ʰ��7�C.��=��B�?0��k��V3P^7�����x�����4a������q���g�uP�(0�y�����Z]���U����t�\�V����(�Q�f�K 'by��l��܄��rׂR$�b耇c\�i96�)�8Q$P�}���p�ǥ���w{�ڠ�^�`��5'��,��C�3���b3đ��zꃱ}z�oxBo�W�e�o�s��7�����5�~�%9���C3�����ƻ�5j�wN��U�I�os#��5re����G�%g��O���Z]iʝ�JͶqLW!�Lvt�A�b��Q�a� ��c�8��L�b{.��[�T"b���OYI�����t��_.j���'&���]��k��6)U����po�!�hq��XO/�P�9@�����[�8פG�h��hLˇG������q�5z،��HI���NGʔ���R��h~V�E\�S&��{���{;�@�[��J%tk,N�M�,/��u)kz�N�8Ӌ��|�j8�s������](�|R��50ג�K������Nԡ���Z�^�*��)��2�=;������;���r�����B ���	"��R'���������=۸���y�,�&���iYU����L�؋�Γ�}����!>U,��<�)��Ω%
�*{��X��^�U���:�܂���F�ڙ�i[�"�+�٩��&�����:0K@a��'Lk�)>7�y�����9eb$��?���)�O�"�d���լ�9��Z�A5���0,����;p�JQ�76���,f c�0�������� k9� ��3{��úm�����%���%���{���57#��0��OO!<�D%�H�����1����.<.��Z�!=~g/X$���h����ח]w���w����!�f����\�-���bv�C�C ݡ��]a��9fcRcz�s���bdY�^^����Z��!�+������bq=*�84Do�����"K��J��2_?_�\ǁ���=�'óF��B��J��V_�꿎u�IM��W��5�IɡO��NF���ܮY^i	��#Iz��k�]�.�s'A3����5Ԉ�Q<̉�w�k��tH�b�ϣ�����Kp�������:P��1�]�N_�;���P�P��w� �AX�io��ZD���V�^�(��!l����	�6�Za��bH�|�OY_�� 08۟�jh0�ZI�5eB+�,��z��ga�
�t�&5�]2�b�5�/i�$66E������Yi1\�g��-��'�!|�:���j�γ����
�X��dc6	��Ճn=QWx�K�.6��aq�񘇉�������	ä�x�Ww]+�Sj}t�P�Gc�U1��iѝ�sP}���L��U0��r^��rD��G���j�n(�!#��8M���y�P	�B�M�y��ɨy����^��"�GI�"�� 5��`Ms����r7���R=�n��~!�?uC@#ԒX����z��4e�Z�B�]JK-��ژ����s�r�+j@5]Iυ'J����u8��L�
U��J8j��q@8%��n�Ʉet�<t]� �߶n>�W
N�����z���Ҿw����D�����t�rm��f���^�ǟП��y��!͖a�<W0;ܩDMD�K���%[�Nzx������/(pq�%��U}�m��F���8Gݲt	�w��1���$�D����(��Ĥ��"$r�W&������(�[���Y:�?�uL�����ˮ�o3ε��U��"~'Nɖͻ�}�ډ�ΦV!�Oz�U��Ɋ���B&W|�3f����:0���cؗ9��;�A{�9���	8z񥊱��UG�N-6���Fu��|/_�q�_�	A���1'W��C����ǽO���'ەz�.�'+@-тZ��DǭJeϹD�ob��~��T�@��'�C���'m�Q|�4�+�Bs�{�D��*��9�����ݻ�����D�g3�`T�*ϗ��]*��7uo�*��U�}��cG�f0t�&������e����9����,��.]�FѤ�R�]��5�i�O�걷��jC�?[wt��1�1�����d�»�Ø
��!���7*�0��'�;,���ݧY�/��2{��uG���P
��H����8��zm�ſ�"I���\L�$
׼do{]>4Fw9M�q�Z=G8=dr��,��ܰc���X��k���t<{2�Ui�͸squn�ّ���#i�h 3ҿ�nT����$��MWңv��U@G��`1��/(\�S]P���G�>8�T�%#��$BT�������&�	O���{K�9����EMťU�G�땺PW��^M�iH�=��w���}d7�	���B���k�R&C�z�`��S��� y��n��ZC�������t��z��>aER���?ʎH�ͪCa��#0xV|����u^�׆ԥ�6��)`�<۞(��{@y�(KK�#n|�]�+��(i64U�k�o��@��a�D����K-��t��׮4F�όi�	�k�=��BF�dh�厣Hףկ���Ah��_��D,��֚�9��0�_lO�o`p��r0E���t�E����6qw0Mj�p������d�&���o�F�@mA����Yױ����0�%��*�0\a��O���#��.@n�(o�>�b��x��J�_�,s��w�E��O���(kJ�����T�(H������^U@x/[
s��������a���$�3��"���%E���Q�z���BQ�!���8��P�Q?�~�.y�^쵕wŏ+��U7�+�w5��;缃!�rBc�UnΆt�����ϥ&I��lBK�}���x�s��a��3���yx��2>MkpX��!2�P�"��/<@�Ѣ::�ؓpl^F���W���J��Өu��R$aH_��"qm���K�z����)���.�Ϯ��9�lR�e��=�-qb�b!zXDao-WӶ_�����'jjȯ:�Zٔ�=��$�^^��6%��x�zb�7�<���6�<��$���0A���qی���8�. �Jf�5hCV�M�����@���*��	RO�7�k�ͽk)3ƛ������:�̓c�kRk��U]|�s��ѳC+���g��DSN75�H�BS�c��D[;l�k�5��YO���0v����R{���7�Cra$�������W+�׎y{��9�[�2�L�Ҷ�le�w���/�B�Ob����Cm�k�l��*�����_���^I�5:Td"�rn<�� ��4���t�9����x:���˗/��>�����.�S��#�]�t	��EF}J-Q~|׳��"�ƹ��Yg�a0N�gL`>| n�!"�����UF�o?q'5ҘJmU>GnE^5�6L��]��[wQ��h7�$ݚ�Ve����ǅh�M�&�mV	��L��I�r�jﲕsTҕ<$��uؒK��ޓ}t^ך��J��n������{#���x�:����k�ȑTu�*��O/".g-��Z�j�{Jqe����B@�O�qAnT��Ss]����I��J1b�@��ϥ]�MqfZJ��9�9���83�	���|I��������ʧ��vw�����y��H�ϧ�\�]�iHc,��]��q��=#%�'�(n�=P�)z�K��OC!��WM��~a.$�H\;�H�/�� P�P�{���w �B�/<|���a�n���g�q�P�������x�?�}��J]�}*-�(�h��)�xBj!})�����ﶟx@�}� ��J��i�5�Iu�s&��?N�؎�/�W_}ɍGm�O��[�Ic��ׯ^����|��W���k?�'����e�eR�ٽ)��Cm���u�����.��To�
�"��}ˬ9*!�dX�)o���W��h#��*�u�ϑ���u�)�
ׅRS9���6��=�܂��Ҥ���5�6+�;D�3|�8�I4I]W��ikT'z���*����=Ww�p1�"�h��N|��a\4����reL��Ue��1Ғ�hkH�&�8�R5�s=��wt	2�1��q�}[x_}�u�*44�]M��\�����	��a����m���ꟺu�5��}p��r�նa���C��-�=7!�N�����Q���W0�w��ײ�a'��3$u��}���<�Ż$�l|+�]e�]�s�J�xw"[c���-j�c����]�ɪ�H栖���7L�`��~m�%�hxP���R$������?��C�����c��-==�5�ȗ/��Y���_��	�����m�|�'�bl��#[P�t(�`���`����7R��q c�E�~�X�~���������ͷ�n�T�i:�p��хa�G*����J?vP��4髰�f����p�g�`�Aa�h�Ib��ZZ�����s���������*����[��Z�����X#�t)�|�� ��ƅ�~sA 0t�h��Q����Ɯ�!��z(gY����8��:�NnEa9�*�x�EC3h�p��%��hXG촓�헵�R������#m���H[�SM�T��{wz�UQ`1�*
�`vO;e��mqCe�� � `r9eE�I�fX>���x|�a��w���x
��'�0hC���=�B1��){0�t��D!/����}/��mzk���lP��z���0����ؼ�W�!�a��AV_|>\e�aX�㐋J��$"���P4�ڟ�_�
��T
۴�&C1gn����Eu[ASwA���W�%;��q�Yg�U�f�Wqp�0�	,�F=��p�].�|��a�JDI�A�e'գ'
Z��1�	hi��st���z�"��q���2��P]�z���/ʷ�~S�zyY�R8��!g; k��^��"�b�c\;�lF��J6� �^�ܡʧ'�GIk/Q=��a��%�X~�1�ΐ<.�p�D�o?F�]p��e>�������f0��8fՒ�E\�[����m�ђ�K�:�5�Gf;�jw|?}���u�ϕl^$��NU��5����{���o����gF�?��!5-��T��>}\k���'D]�>)9�l�IG��-<p(����`���؀���*�<+�f�&�s�$���"�%�{R�N�FJ�m$�/7�Em�2�<�ȅ�V�ۂ�f��R�}���nO��x��ó*z7�b�R�����&=;z�x�p��������O>D���`?ܑ�l��4(������|LӋ���-n�
�p��%ۊ`�[?�i�����kq�OO�Hor�s,/mB��۞�|�Uy�
$�G�d<�	�A����z����67����KW��'�~~������'�#�u��e��'�b���;#Q�B(*�Ǖ�f�N=�����:-����c>��~��.��rŘ��>qP�6C4X�T�ڌ>��iN��⋢���������#�051H�J/wc��F�R���)o�'5F���>e�ɂ�(C5G����n�����[���
L��ҳ���]U��r��m���3v���i2����j��1:
Ko��\��V�k�1fw۠?��k议�?39թ�s���0��_�!OfǢO^��f���=	+Y\_;��B���ә�"�G������I�V(qCC8�S���5����6��L�w(�c�L��=qx	u�L��C�x=�������y��-%���O`x�����C�F������X�\�0���$O6��leN"���L��Q�Sxg8�C0�;9!u	��j90�`C�s��5�]%��m1��!D~��{��ڋ��.��g4��5�	�Ib^�����_���mPU&f���n�b"������������s��"e�5[ ��a��`����.��g�ox��ާ�u1#Fg�7�4U��H��>S��D��,���5ƾ����oޕ��OYb���7���1_���R_���б��3�'��w���-��_��8�L@)�d��ԏ��ʓd���EG�Btao��񖒆k���98<n��0�����#����b�W��z�:4�<4���������0�CCO�xf�""`�L�~N���ձ�r[�;�F�RѠ�����,bM|�����<R���?�[&|����3܃�6�JH'�UN� ��0_��摾(?��3�?��s`Kj*G�8��Sd�JcDC`7jr�km~��a�����E��n����%��6���L��[G ���/�Bd(��<Y$#�PN����=�`�x���J~D�v�cC��Ʃ/�
?��MP�W���N	�ɚ�2�$��3�����c���������n߉q���#��?��C��+(�+wm=�U�q�g��v���[����曯�����{;l���T�6f�8��"��z�ۘ���w�����ۡ�[��`���o���-�Ex���w����c�jlH����]]���5|+A�w6����&��X��`H�G
CzwI�1������5�g��Q!�-��������ٯ��e�|�T��<�`������ �?��Ss���a����T5X%������P���j�^�8<r?z\��]C�N�xb�=~z"�	�] ��tD?3��՞j���􎸌A��>��I��8�]�$��I3?�� OQKBb�lo)��R��*�Mll^�+�6��+m-�X��TX��K�k<���Ҿ!5ϲ>�u"��X�lU�.�CK�8W�{�h���M��;���������O����Y�iW�I�QXNp������������[.ns���a�J,d�7���81<�!`b��йD�B��RxxJ [�%\33���cL���SP�;����=�܅��L/Ix~��İ����n!���=���RO+`�7I�Q��MO�x�3a� �j���T�_m�A�T�N!}&Y�B&�#�x����������eL!�|�������W�y;�9�=�m�$�o�v�)�2�s�D<<�c񓚧��J��m^8�>�dl^��*����l%8�4:����Ŀ�#����q�$�3mX��3���k�,��?(��蕱�r�V��ϫ��I*eE��F��I��%.
��:%����Ն�ɶF�U`څ.q
��c8-s�0�����G���!Q�ͣ+jS\"��=�>�a��}͸��ۯ����liS��_X��W�xCB�;X?�����CgfhCz
Bl	�ƈ}s�!~�7�E"U��l[Acל�|؅Qjq�.��tڻ�1�nCߧ0�]�J)3DH_�R1� ���&{)E���*p=dT�$���"�vOh��O���'��(N���&b��fdDeP`x��Hw��Ϸ���u�'��t�=��q�����?H(e�K�<��~��M�0������g�7Y.�y��p{;0���`P�w�L&�#���f�%\l�%a����~*����f�ߒ��7���J���ű�(�I.�뱹�Y��"R�sJ��f3�KV�� ]��������)�m�١w�ד�}6�;�B���!r��pTDL���!Ն��^x�(��ݷ�rnp����?	�`>�lp3��5- 3�ASO,������N4�ǧh�3$s	�~���yO�$.%�2�O�<3����(����qfS+\�Gy��Q�{�����X��y홧=D;pU/^2��Dqe�V5�s���}'����[v����:����ꚗm*C�Gԧ�w���Q���/�?O�s�j�^֔wC��P�ޱ�o	��
X�ǃ���Co��BZR�Kʈ����ݲ���+2-H텅=���^R+S,+W"ܳ!�6��@���8���/��ɐ�l���Ķ��&���0X����Ɗ�[^��D)x�Ґ�F�a�fD]���Fx������1Ï���矣��nbsQM��w�&���維�ٷ��[mҳ��慝�O�)�c�~C�=�.�l�8�0����e�;�Q�7
oM<�[Q*�/jA���j�����S7���:�&��"Arz��`�����<�o"���p"�]m�a�����]%[ԓ]�(zW�3q�/7C��������s���'��lb��t��1�p�w���Ɯ�E�Ѷ�t����t�жȁZ����=�2Bez��n��	��K8$�N?��N�� I�zH�Ť�SP�B#A��6jj* �?+j`��,�,T�ȑ"��<P\��H�uW�b��|�.%�ҹ�=��ӧ9����xCȇW�b����M�\��#���s#*�o=�L35o��Mڪ����P�«p%S����v�&s
�ݴ*W$���F�5�����LцbYݭ4����U���E��y�Hr�C�ñ�:d��gy
j�2h�v۾���9��C(�/)ʂE�:�{�yz��D��4�k�*�w�� *H�jt����Q�y�������JZn�Њ�����8��WW)c+��I���cS����ƌL9���N	���W5�T�!���~N^������R���U��eZ����	��E0�h'�V/�������1Ϣq����7�D�uM]\+��Ç]�B؁��g4�싵����x�9���ڄ��L�������'�Q�ծjO;&QJ)�g��5��e���\�}{�4E]QYEX�Ɓ�����������(J���58,�]���l�:F!�iU�RJ\�Tқ2�-a�z������ΠC�r�+�sm����"kae�` �B��|iJ����n�p�M�}-�S��Q��l�5��pMFNk`�L!���=s�]I%�]Ы�.p����ث�Q�I��c$~W׽�Њy�0�}����7Uo�s.J�kE�ffp4�.z�8��d��wݛ>#�0��A���Ccdq�1Ĳ�!�R��K�^��*����f`��_�R����+b`��CӘ�{�=WrO�!��k���ay�L��,�Q)��������XC	�Cc�X�����_���G����`(��bN��<��g�u��¸�;zL��M�;6�8�wi@��f���Y_t̶��,����!6�ˏ�u�]��aX�	Ǟ{|RKo[0��pI'�N���[>�e�Ȥ׭_�3��pm���{]*������1Λ!c����l��M�>�6,tԻz+.��=���+�^y��zi9�u�}���Gg�)<��ôL���,���"ؚ���K���ܘ�����[�NY�p�/SXp]A߻��:rJ�?R�@�$n3��!d���A����X�Ŋ�0\��h'�ܜ�bϸf����sY�΢�x�D"4�j�_��{k#�V����ӦRS3
Ta��]P�`�0>���n����9����7'�*���G)2�!Kq�������H�� ��u���Ƣ������ߕ��C��_���B�ɐ���Q2ȇ|.|������������x�ΙG��9����5���D��W'LM��plHa��>����f������=	���!u��������w齐�vW%ۖX����%�Yb�P�Sԋ�PF�)hi��0BC��\_���vL$a�2��pv�"��u����=�ۛbؿ����m��`�@y?yo*�>�%"�Y���v#�]����
�i��6v�z���4ϭuj"L���Vf�`��J�ĥ��=�v�}�8g��j62�S��叠��oՈ�����?��e�9g�-a��	�����V&�'�v�Ľ8|J�t����D3���x���ǣ���a�%,�)q,��y3$�~���ڕM��� *�{I��)�����IKe�����N�i��0b��}O��v����,�g��..��a��2����1�x��/�>���mM�2�������z����1$��������葂�
����Sļ���bx� ��X�3��?mzR1�xP���)p�����j�"��t*|<K���<�&��ȚF�&��6cx]lo\��$���
�witi_!���HK�Zd&�]��6�i����9Go$W�����鲂�R�(�{�.n{�Q��zy����a.B�,�kۉ#����7^�^*]XQ��dr	��1��
�?#�y�qpT�׸��;�o8HSO8���v�I����k�(�:�����J��D���6�����g��`S��B>*1���K�d,mD9�}Md$�� �x��Z*N�������y	�>����(O����\��D��ءfq�1�JWZ�i�k���B%���$?D�^���,a�Ƕ�Ϟ��.�崮)��l3C�X�.�3~U�/Y���^���nv�R2�=�%��B��k�&���z�6��H���DԻ��-�uFs�l�׭$�j�Q�OCu��t�f56i��>��u`��d����k�ؠ�5>>�>���>V�6���[z�dE!A
���:ĤIqR���`�j���q�y��1�-Aj��%��V%�ΧS:UKbI'�/�y}oQ��j��b�BPs�C�d�h��P�&��W[�j%�`����_�f�s>K�كdn8�*#6��O���(��h�G{�X�.-U[�c0'�
2{�
>$�dSqw��b�|η��oG�Հ�����m>��o�Zsl֮v���$Y�<�]3	��:P� k�����3pa����˸���Ioyf}-�Y}ډx�E�er������\b��x���6Bć����X`Y����5��Z@�%�_���C�{H��dR+�,R_8�)6������<�Xý�!/"\OlVx0x��@�z��%��,��m��#�Q�!\��E�G���AI3OTf�����,��ō5@,��o0ڡ1�2�cx�k�^>03��F�s���R.��>��P,�톘]���Y]*�*e�FI'�� ����~�	�60O�;�|=��}$Pv����Œ�u��6B��Ma������p�z(Zs�X=���L��v0~���9�,<��Z��ԥ#����9<Y]C�
YW?Tn5Ǧ[��H�ܒ�!`*s3d$���5�ԙ��@v�`���fdk]�ӕ��y���}�mDM��=�zTt؍�/1�Hp�<u"Cf�,E�WlQ?3�����a۞�����6"���I}Hb�ru�t�i�1L�\�&�7���|��^}�6b��������N\��t 9�I3��v��9�d���#v�'�M3��I�>�{��5|NW��Ӗ}���z�!��I!����J��5��?���p���d��]�����!�)-Q�e��b� a������7����k
i� ⾔9�D�(�Nﶟ�e�XJ�t��� x/���oh���ص�/c���Ӏv��	C,k�4r7���{6���c�B���������)EHv�Α�]Y��q��f��07��m
d@�نC��.��X�׫4^����`��L��է�Lq���	�l���o���?����,g�3��1�E���wsť��]�1����cO9B�#~��~������� ��ʩ��%��o#�~܅�VeY�ç��+�a]"�dxNFTv}$���������w�`Y7��^�`^&�ߪi�}��~����G�?vnߨ�U��76��1Ro2sX��Fy���␥+]/�B�L���h�)4cS�}:�uF���ym��$����P�]�Fn}�2!�&���L���R�y�0��L���c�FscuR�b��IP���J����gE��q��;��%�Dɩv�� �������|����xU<pS����j�9Ƶ��I�)�/|P����F��&ۊɈ�ϡ6!��ÛS�(f2@]&%Z����9��:����<vg����c��.��I�wƗ�)�����I�"K�cJ��w�>9����[� v�|P˔+�K��0�_�\�7�|C���1�:;N�.��[@�0W��C:?I��E���J���.X	C����]�&]{war��'6<G䱬��>;�|9g$�Xi�s0`N��R5��՚|V�N��K�;�B����[����ϵ��b#���=Ғאa}pK��#���=�e6
��ye�&�r�|��	/8���=�.���'yFE��YmL��%�R��q�{���{�+D���4�/��P+IL�Q���:i$V�`�eeR��$���=�4�ۢaF��Kb���j��Z����l��q�ws��J�<lR�s�I揽���,��5���$<��Ÿ~���̼J9��w^%�G���3^��#�ܢ$��9I��5�q�P0���xd���jD��ܮ��F��2.4� �5�4�݇��^�!:#A�g�h%��:E��[%a��a"��RJW�<�CKB�0�qX8W�l�Y�����]&O�������S;vY)DJ0�/���	Z�Z��	Q�S1�a,�p;�nFiZaǰ��� ��o`y���� ��b�u�ys�WQY�)����
��qﲶ"��ۧ��m�"�K2|ҋ�h7�O&���J�duD5cY�xxo�Sx���ж��g	��2��hKK���w��]�x���$�*y����(C�ΚcV��Iƨ<��F���@�V�.���J�+����~�"g�B#��DI�1�������Ğ0/�y�sH!|LRxv2��I9y��X(��z��\���?Gi$ƚ��,�������G��?��+iX�ٞ�q�h�gx:��K�߷\�
�V`8\��@u���0�~F��%v���(��ږ;�@�탄�ק5C���+�9Q�q�8��+�}�֐�8Vr}���m.��?�rI�v���5<�6�y�lOT3}� ��Ƈ�m���A���^�!�:�r��2�Q����3R��F:�4�'�'��Ȑ>�z�u�Q�N��Z	d��%��Ү��SY(=�&����9�l8Cl��Vg�X[�I���>ց���ݫl%�a�̒���X��^|���zZ����N�,c؁r�����#+�6�Jnm���kK���}nN���о�@;��p���sT��iO�ւ=yNn�R���x�҄^��>_��(��� ���gumo�6�!5�1�@q�N�d�C�85J��Tr��~Hc
� �G�>�ZҐR�g0���p��s��")"�_R��=�³���a\������4��t2Ieq�t���ު���_}�q�1�UE�1�����=�'��Ht8�>E).���'T`�8@���J�z;�!������,1�0��@.p��-K�WLf	�y|����t~9�Z~��M��]�����c���[��B\D�K��6�n	`��/�܅�Yĸn���0�<saA3Ú'v=�G��u
����]��*����SV�����֩�{���p��˸���?��ch�v%�	��TU�X�k���Y�=�ġb���X��Ú�Q��sHoO��L���2N:��j%��}&�����I�]|�y��'���?{4��C���&w��s��鰎�sc�(� �`u�>J����U�ҥ������F�F|I'
�P�9D�)��_�,��޾5�.�d�uR�YW�z�X��k�%�������M܈(�,ۺ2�G��>��2¬�a]�G��2��&;fV�8|��\A�q8Qj�ݻ��~(���/��'����@U�%�������n�u�)Y����>�C	���oB�D8��eM�#n[f���1ď(=�^����7�-4O����JOV8��V����%�v�d���O�����K��E�7;u^8Ň��S�y�.��O�S$ N<h~�<�����xQo#uT���$��R�x�p}�:[�
���N�.�!�S,VY]{�����Y�#ˋ'	q�;ȁ���D��qX��柆���y�C�]xhd�@�_�*���c�҉��&I��)���Y9n��?~M�[KV��A�s��{�'������zϗ��լY�e��P�%��ژ%ıd�!���uŽ��9
/��TB%�u��v����8���=������g���df�G�y
{<'�BZ�վ{�aux��\�[t��9BQs�$v�1đ�ĉ��%��,j�:���QU}�^�U8�R3�����<�a^`�c`�a�y��g�hv,��RXt�g�7oB�|=�2-F�0��GS�7�v��/����Z�O�+f2Bq�)�Cp��M��a�=�B(�/��j�ܴ�׺P�Z���������	E�j����c�ш��o�oyM���&�l^�/0 ��,=���W�����c@u��`!��"��͟���)Y0��`;$=�Ɓ�5
��i[C�%b��6f0�0D?��Oz�7��T����kU��~d(���k�&OT�S�6� � ե�c�ŶWXauCz�gI���׉93-l<�2����3�x�k�p
�ou׻<zU��uȮ�̶/�Z��0�1�X3��¿�r�R�O]�(%�Q�G�ޟ��b���$~���0T�tP�A��wGm;���w���SG.��ƹd�j+y�\Zz�v�?��?�a^�Ol�=��5��
黰D�eRykDI����M��.�H�>j�w� �z��a3�E���=Hb�0Vؤ΄2D?�i��%h�22���x�s����$x��d({||�x���]~7�3Y�I#����������t<,f\76�K.�ĵ���*���3	^��e���������R�5�`��Q��~~�p�}o ���8�0����C&=�{e͟�>�B��X�#���a.%�b�#�YǇm�u0l�ǵ� ���e�M�ۻ@a�w̃����-�As'�������'	Ct�,:�v�w������/��F��O���w��Z�!�Ѣ!���k0��!uj�Z�R�vM��z�pw{a��I�b+�����~;���P������'e��i��V�F�6�=�|��7X�R�'�qs#ąn�.�6�8�q�1��MA��E-Ä\k�O�T�7k|�Kէ��NF�KC���j;{N�Nc�!;��c�UEߪ셅1����,��,�Mc���?2��G���2<���#-W�K<ؑs�Oe���(�*)�+�	� ��'g4��E��J�5/L#���c�{���E�"s3Ǧ��']E5Q%3�}�,->��lT�Q�Ix�O�'nc�Τ�5����f(�o���#S�'F�*��JX���$)�
���^���X�6�����
��}I0[��9��=�v
���Z��2F�Q�6ju����P��-�N�oW����{�-�A�c �O�t�S��=$p��t%�$܂���?L�F��݆�4mJxaJP��v˰�I�0DNRY��M�{�:��6Ը�K� ���ǀ�`DѠQ��.��U9aI�飸���@^��HԍplB�#G�LCr�k� 4�@9j{=e+�@�b�+M�oE�X�4��T�+��ō���*Th��}��Q��2}�X+�*:�)�mDI��P�%�_�F;ӱ���}�K��P�7{�J[UK9����`��y	' ��������������3um�����Cõ����e�L��{�K%k��%^m%�q.c,
��{�%iH���4��s�]�P~~j����l�R �FV=��  �����;�2�v�w^�1�	��租~REKp34}�g�!��)��c��!0����i���=�C����U[���x��\5�@�Z>G����ڿIc֙�Q��Cȓ��K̽�9�m��D7�!�(��g6[�B��$�l��WBD����e2��_T�b����>hX�f�អ����#�q�xF"3n�{����Z`�7��<�]庁�] /�~�R�����?D�s����D�H�d)97�<�@��v�.��*���ό�p8���OC�l碄g��F�����B�YPK�y�Y������k��Q&��lBMz��!��8]�mX�|�����d��CeCIOѢ�L�"��,
믩sm��V%�l�!ʥx��On�'-ђ�5�l��0��V�ħ
�E��Z�[4�.�?�ssFN��6���t���հ7�8�į��}Z0V�J-p����>���gM���$�O曣`AY2`�
a+�\CK�Ǡ�z���Ln�0�
�?e���/qx\�,��s���-�)<§�6�;&�Jf��!�Ӑv�Aݲ�?�ޏl���S�>FI)QR��>�z���������t}���}|b)���
W�t�WB��:�0,s�w�5�6�3�.I�_���J^��y��n���$0�,�UA�O^�"����7�}���N!��"�i9�p�irI�|EO��0��d���a�GK-"3G����� ���v:�M	9G�O_�B�#�o/s҇�pq��4W"��zL��Ԯ1s&�������&3�Dy��G%5D�+��*����Z!5���(&��ó�I��Z���;�0'�fO¸�q��A��w?�[U<��pV�T�#��'�L�j��¯�
Lcz(�ɉ�� �:���$Dr��Ё��3V�sa�����%��T������@/�fy��c��ܰ5�x���r
5�'��St�<� �t^t�||b���<���X������䰆 ����1Z�I\wɝAu#JH�܌��44"Ӭ��!�����w��γ{�wN���!��=�w	��a�tHKu�8�NO���9���E�e� d����cp;�[7�&.ġ'�AU��7�A~�"�yZҘ�!�ü:zN��C�8�]���X���;$�v��8с�?�݇S��kܟ�	�7�I���P�f�����(��((0>�a�k�k�]�����1qыү(S�F��{hNUz��C��X7����qb�1��9�^K��[5������3����#�-�m�X�s}^+
��qm�mT}�Hd֎u=\x�R�Suc�
�q1VV�k"�V"��g��ז�?��9ѩ0���d����7,.Nf�T��
����h,��^I�>H{��^�٫'٪8y�g����Y�
I'�l�:�u��<�x�pY�3�Q�?k� ��6'��7F\�L�Y^({�r�v�>nV�t�3#���
��VŦ	�*��ƅ��*YfW�0q��{d�
4u���F���TK	sE������tʺh%��c,%��t����fh>���}5�����üϾ��-�rp�}�n!4�z��LkV.ל�%
G��u��za�<:c�8�%��5�������9���r<"A��l։�b����s+J[M	�t�+iT��m2�\y�}-:!�3�,K4��C�i,$d���eaO�1�	��!�Z�U�"����x?�	�g�q��1��.f���]����H3@��k�p����L�I�J�W2�gz��t�
�퍖���&�Jz��^����O.�BHm�{h�#U(`umf��t����.��,1^4SS��!��c>[2�����H�X�Ș��Ϋ��W���=��*�ӻxۭJ�<����D`a��=S�ݵ2��6Y�m��a��J��ҷ����R�Qj��ł��VVhD�A�+Iկ1��e��.�l�I2���K���x}�v�{��k^Y�m>\�#�C)��<	F�F���Bn�1c�,�N���E+�I�$�W��Uo�#f��$��w�'~D���I�:��^��E�H"��E-?���{�z�H;�mN��z��[�Dey�fP����t��1i<��x��k/�9��G /�e���n��,p�==Ȼ�o��k�j����cDe��jRY��Կ��_�p��
	1�\R<�<�W98���i��ڝ�n��̕\.�	���M��;镆�6�Ø)�tLQhu���ɦ���1�W�����[������4�!CƓ�	�����,j�a�A]zs�4��@[��E�B�����F@<m�l^hP��xd?�W�j�ҫt��}�j޵p�|j'}�0�A�Ϙ�y�0_��������=�uۃ�x�6�'��sx����ī��`����4���� tPȃR�i��YJ-�5m�_;qE��$���ڠ�^'��{X�7kt@�I��S���8�2�E�CO#�J�ٙfv�l�1���0�sxS]gOt��mm�3{��DSf���>�u�GY㲖L\�hԎ< Q��ǒڦ>��BU�a���cw ���qx<��C&�����F>"�%�����0�����>4��0�i���������h�=6�]�t&Q�(%�p4�z�w\�r�g�������H�u"��OAӺ/��}��<����`�T���`B����G���In4�F-ib�����S@H�
r$j�ЙB��1��6�^+�e��a���ц�1�W?���1�DYf�׶�=�к.�P��L$�c_d��;t2��<�����v�-����q������x΁u�"a`�K<t]�{���]����*��G74^P�[5-�d�*L�ז�;Wq1�圸�At�~U�	���BBor���m:���'��K�dH�Q�xv},�9k��Q�v���+�X���UX��6`_��H����7w�=灰DM�#�W�j�!��ջ��?
^�3�c�z�oc�����j��3æ��u����c�]�K�{S��,��ac�J^�0V�
�hbUVR7��X/N
9����Q�h�w��aw�CF�g��ֺs�-��O��iI��Y�͹g�Ɋ���t�@�-}�+���j�� �A����lX����5R�s����]&��HVK��i<�{z����!��#i������ 7�x�cj��� ���2!0SU�P��3,_hXݳ��*:���Z;?0�"Xa
�B�g�nYq��mei�P4���Aa2 �M��pE�*V���>C�0�d�슉C��u���1&�ba�j��=��tE�a�� �{.V3�Tl��L�nk%d|#��Ơ�^%��r�L�Hx"Ad愠��2���q�=�4��E�0V�n�׸"1#]��e��`o�5mp&j��m@i֜�cH�Z�yQƾ�Nڹ;CP�lԆ���t��o8+���֐�)�D���'*V�(�Duޅ#R�+��:s�>6:�}��Jvy���<�[c{L�6K�{w"���`��z�}zo��?�ۭ��5t&� �]���^R�RG�����3���N�.�>����*Ʉx�!!�>Q� �"��|���Ԭ��ظx��4�G��&z�~gL���'�%5{op�UM�N��uZ�6q>���9���`��W��]���u�R���<������rKj{���B)�(���Զ$�7�g�&���.�_O&�?X^S���9#Q�}���Zoץ����QJz�]��2�5Y`~.=>�	$Ew�D�����cH?W�cSH����r�yS�U�C��d�Gh|c�<QWr!�B�+
8�X�
���)����ީ�t�]�;������2^�����W�^r�]� �ld����R>�m��n��v��������Km-�sqCps��YK�Hm^��1�وWY����:��~8}��?,�p�vS9d1K#����e��q�^����BK�6����DG�&<��MAK|1BjT�Z��k�.Y�VnK;z�8��;���*���r>?~ʜ�x��=�NQ�r��Z�)n�)�L���Y:`��y���`�3�h���s�uu�W@�ځ+K���2�lL��v��:So\��5�t�ך5�i[y�Gzݣ�m��ӹ?��`9���F�E?��8��3���z01Ԥ�Jh[��ۆ�N��A��I咧���%0$	���ԗ�{	�����~CR.�r�U��jYZ4�pc�l�8-a���l�ݺ$�d�6��$�ӑ�l/O��	�W�;�\/_��^Ay���%,��
!Ђ1�f�|WW�&{���K$È��c�*Ԧ| ��i�*c{�bo(<&Z�����v��n�`�LCY*=jH:��U�>O�I�3�p �������k��Y��mwA�P�m���;\��CrNbC�֐�}3�QaS���5 %W��h���@�����$v�Cqa�UU\�gnťH��=��z�"������41�,��	��@6マ�t!�к��À��}B�7��|(g�TӇ�Pey����bB�^�~�_?#�-�l���s�����<�!����U	!����
I�W����2r�w#W�V��z]�
��_���~ICtg�����7�E(L��wo��l�hlk���O%��$����C�}r��_LEA�U��C�D���\b�ج��d�o������~��O� �!#���V�I�X��k��C��"�\*���?�Vx3+��Okx�%�4��9�� �PP����f���Ik[d��}~^�d֎F��]&~���A���R8���t���f��q�<x��Yyq'��T�^�k�����=��8�a O5�M����q[g7�����]_�2Cޅ�R�{��x]��m:
h�|'y��.��e��|�����C��P�1v|��%�f��^�SߥPP��&��b�쬄���v[���*��#�:�7g�4)26C�nkf������{ᰬM	ys�`ɠ#�:���v�J�Qc?��\�m�v�f���d*�Ms��7�����z�������_;$��P�l K]�f T�M{V9�)�D�}�d4hG��w��~����̶���Px����Ր�Cu`�����ET!1��Nl�n���#.x_8 �O��m~�fL��l�S��?�")y�k.(q��������5=������m���qϐ�`?��%k�UB�*
U�&����$��D<_��4eB}_Ss�Ԇ'єzZ��8�D;hh�kdPZv��nܚ���(��M��$��ɭ��8����!	'CZf�Z�4%\���=Q����p4eK��� JOOe�~7$������u�[YE��{�<nƒun�3� x6+��C��@���9��9&�n�!`H���iL(/m�tڜx�����s����Oi��v36Z��bW���޾|��Wعs�30*�
���ژ�� %���A�"=i$[��-��YF(|`�>>\��,��׫�}����}��c�t�����\�X?=sVۖ�w�B��"؍V�
|��!��S���1��N��d����ڤ�����vaC����jn�Qx�_s�kF�3;��?�2�5��Ꭵ�#�w��Șdy�~F���q�33p��L�Ȣ	.��&oF~'.;v>'N�v��4U,L�6DdG7�ӓ�'w�C`�ڗ�RЧ��䅒-kV�H�t����	����¢϶a6�2�5Hֵ���cc�Xx,w�X��C�����l�q�<7o�yP�.i4�`��rF���y���kQ����M����(�mM��(WE���/K�Q�G*Y��f�|c� 4�۾�6<����C�6��q�7��-8h�߾����Ǉ{�ԕ}v[^�|V�������QZ���G�����0��ț��'��ֆ�V���ё��*5�����/�S���Ǐh�������O۵QUڲ#�͈�#�Ð���<R55���Q���,�r���L�h�]��<��=�$��n׾���N���{�<ExCx���i�!�CLC�dֺy�=U������$I�b�̌.]��y���,�C�G�I؎�S����W�%U�P�]I-Vm���[Ѯ��>������Ë"�wI�0r��7McM����?0��V�������V�z�7\�_�4�WV��]��O�
h�2AG1�ݒ����%��H��ϖ�Rkla��/�
=X>�޾s�V��x�x�떍�bJu�,;}�:�%��Lc)�����$�E���LZ��XI����jf��'vt!]_������3a?�p���c=� .v �ɫ��B�W"��s���]�����:��8�Y��$J��YR���$������w�p��!�1Re�W6��w&/w�o�B��8?�_�ܞ���_ыe�9��`gHV��w��Q��ܨQ��P�T�gw���YTm�b�^j����	KE�.BZ���3,URt.�%7����[9�g���@��ah}�񐸭�z�����:R��k-� k�(�=q�����L����~:J�H	cS"��1��1C�����Ո6��]��\������Ⴞ2I�H��!�x�VE�����#���m���ui�j�s���g���x�`���Da`�����t�K�l����ߘ_U58���	�xZ��)]d���47�1g�d`;mߠ=M�ū|;�ָJ�k�ey���ܯ��`��KL��jt���t*��Z��"�Դ��<~�V�08x#G�?��f۠��a�������~��W�s��j1[{Y�N]a�@��M��:��Vf�a�u*�|̆m-��MRrQx��9�P��vy� ��Ð���w+<�5�,����y�.tZ����)��<��� �m�σ��%?|(�͈�e�u_�e����>1�_l�ź���u�a�
l����K��fK
�������B����ݭ:hx��>��P��a�ޖ}�)�w
��]�V�NC��0ڨ�W���~Z�zD��.��<EDW\�;�7D���!y����d�j.	��Q,`�1�B��m��F�՘&�����ϠV��ަ�>��{���=�b��0p|a�1	��y�V���ۡ8ӋUe�%D���������?K��v��/��jd���Gʯ���7�+�����C���\����wR4�Y�*0`W��Bw#e}u�����x�I�I��FU�ifЇ��/���c�0���|�&v�<���"c#|��������<�c3���2�m��:A�2��m.��+.�'��*���y�MN�B޳�MtX|b��������D���+gI�A�����VϥU�u�P����D���I�q�D�VY_N:��gx�bF�K���NzK���fr��Y����!�pϐ��a۸_~�U����JzT�8*�|�����^����>]���=����<��N!���,_m��:�xBQ��9:��$.�#ؐ�`�H�h���z�����q%�lxN�� x���ޤǆ�o���=�S�e;����,}4�� �������?�R�V��Z%�[o���n?6%.��:�)�HoRe��h%��k�B��*C*�^�=%����g)T��w`�@��ի�������.#پ7�`��]���~f[�Q_��V����Q�?1��Ɔ�CZ7���:�� �[��5�ChNeJ�B�H-]e>�Z���1�B�m���u� �q�Z���	��ZE(��>��,Թ��Y5�k@2�0nh6�������n`Ha�ݠ�3��P���o�����v��!�َ��<�1�'I#��`����>H�Jmƥ����(�%��p��υ��C�2�9��`��6ـ*"� �j,�n⾸��J����.�zI��ң-�Llv��/�������2��#���*���5������s����_��C���������
����q�L��_��(S��,�:�����=ҋ�}�/^��������?ŵ�܊���ٳ8�#2��ݻ$޳|v�^Ԙ���[���a��1e",(D��*�ּz��?co��q$FfV�t7I��fg����}����I"�7�:��473�(��TT	h�P������9>{���~��r@�Tΰ�'��]��웈�:^�7���B�����;P߰��3�!am���K���f�l������{�߃�̲ҧ��ǈ��s�+ƞ1�#
V�{���Y�a6�{GG��,}�% �(P��,��q8�߳��7z��^�w�ڻ�[]�)��(���s����E����۝��]bb�]V'E���\�6��#T�i��Is"1w������+R��H�+���a��Q�O�H����O?�(�����}_;�fF����L�Er5��]�/�F9���g�_�V�4��g��=9ApaGE\׷�����%�����d�`ɋ+��6�K#%�=�ɕ��%�uH�f,l�s1��l�;W�md[؋C�m̑Y��Z��4�_�� �?����K�2�!�|������0�2��gR�>F+�V�������D��zۈx?x�NJa��i��b$�������p��?|����횎L��'���=� ���5)~�e3�WC�Y������5�+�5X	�Ԏ�U���׮���U�9G�l@ a(�Ȏ-�٪�Q]a�c�0��Ӷ���#7��^�`�QQ�5��	���j�b>�(�"0勞lh���V�p$�K�} �X��!s�]iݎ9���ꝲ�ik+��N�����/��4�i2'-�u�摶ofC갳��2����YVd�#�pu]�ϔ�h����>�g������B2�ť_�P���$���4��6�:�`�1!*����@4GL�8�R$K��NȾ�0`�K��X#�:.�G($A0<�sdP?�
>�X����
p7E�t:����D�c�c
_���:P�����I,by�)}7L7�׬F�v�8N'yħT���}Q����t7�AQ�t��ԣ�I��J�ge��MNm��P	���
�? y�M��s��>G8��CM?	���əY��К,����߻�xL)��M�y�h�)��! D�^��.ƚj�L6�JyT��!�^#�ެ;��=b�~1ָW<L�k5f�ی�]py/gbӅ����]�Y��(�1����%�(�0�C���W/q��o�8�4��+[���#�_�@���NIOt�s*����Ÿ�ÁѨ�MCr�t����:E�S8n7����4���~e�~I{�e����W�}{��J[�wԟ���y1xm�"%��e�q&�0`��j3�]sq>9jQWL9�ލ:�X@��)��V!���>2����2aR�#}���������O����y+�X���i[�0���q���+,J��Y���ҕ5Ðv!x{��S|>��+gb1��2xćX008�a�z0v�ې�c�E#��H�����';�fѱ�!��G�I7��o�zN��2DU���,o������R�Q��Y_�"�))U�v��'�������x�?��>Z��!\fa�'�M��#x�3�=��9���$��G�Y�������F港�R�$��Hw:l:U��H��=RWŽ���jZ������H.UڰK~����!�ǔr>֨��юǽ!������sQ�U�߈lP�W_��BΘ+F#�J���-�|?��z������sxPdUY&j�N]�C�{~PKq��w1v\K��1BĴ`F�E-�Tw/s(o�ƴ�m��u��qH�M�>q���:�L!E	�ǆN�o��l�j� ��.���]$. �gYL}PP����� x �D���tL�m��u�X�z���-ۥ'C���vǘ$`F�@�4!Ģ��!Dq��/q�D�Yv�Y^9*�]�l��q���y@�R�^�8��;����`���e��c�n}$+^^N�5�$/�v�~@�i/l�ka��p
	�$E��p���B�	�.��y_��*�p(j9ž�0�vo/�UyQ�x����M<ewem�*��Rw]V��a{`gؐ����1������e��nG����;uJ�w�	�b:�R�%���Fu����1i=6�*XG{E��kz����I���N�#�z
�C��&� s&+_�$��I.�+��b�`��I�Y4/�=-��7�h�AR~&�7��7J#�h���VBA�dS���4�NV��� u��޲��:�E�YM�$Hzg ����ImR��ldY����2*���"��dΪLԽd�1O�bü@'4Z#����7�,�7������:��&�K�}y��6�����Nde���D��܉q�(�9
��>/B�Yc;�-a�c���(�����[B��B�Hn��3k�q�/��-kme͖�l����]y�V�b���[�����g����d�/�����J���ڮg�a�>��E٥��P�R�[�O0,�|�@(ĭ��0�����Qq�&E*0ե��Z�c�J&����ފ�6��//'2ҋ���]���ʨ
G3�r��}�\�xUr�M�e�9Z�.�g��T���e`H�糄V��;#&8fXLn5��CVEb�M�7�j�J�"ӘY~$5��u��,(M�����0��o��o���£��`������-J<�mªr����x8$�g e]n����K�Wj����-xbJ�,}�ྑH���P�Β��=�N̒�.�g��Y��2_㞿4����'=;�kIX /���J�	Q�4�i�]�h����|Wa`I���S�"���>\��w�����@���M9�	u�˧U�����80K��D���hNG�H�w�����q���1�["L2���$V�q
�{z�*+1iD���~E.ݗ�����X,%w���I0�O�6��%��/��B.$UT���-%�`D����$P��f������%�~�XK��g?tpf���Fq���;���/c<.���.�R���#4�!f�M�6��������0>V=�5��c�wC�	�kQ���8�[m��ۑ���t2�
q��ؕ�_S"��wd�EP��4�pquT��<�s�]!����!�W��z�71�RZC ���*��k�j��(���|���t�)i=��x3��d����5GF�1�6��%8��~���p�z� >I�kʪ�h^:8���P�6���a��P��T�Ev&2��������n�ID��ꃼT�5�6�6��rIWu����Hm��kT'%���������׶�L�nMյ_��f�a�B���n�����X`/�7{����&'��G��%�媖�+%�T,g�Ӎ����n�k���֒H��H�t���CQQ3n�2�p�I��"Ga�,<�)��1<R&S��O���a����&p���/ݮ���FZ�}�	�؛�F%/�m♗�-���Ң2@4�Ʌ�7d@�jQ�6l;$%s���Hx��0���T��^��U"�ӵZ��� ��vip��y��
O�<�亳?�f��\�X��]�Gb���E!�0�b{��׷���"���4�b'g�We��]��:���6?�oh2���X�Y�{!c!Zq���4�M扞�������՗L6/sM*g(�ђz0�8���"�j���Zp�^)��(���Y��zN����	��I�[���*; 0�טA�S}~��לc��|�{�gOr5����k�R�GҚ���ԕ��5'���Y��=7�Q�T����rRVSt���v �wE`v%��9��,[mt�̠���F���AE��@�QTT%�(OnH!�S��,kz��ĭ&yaK-a����"h����U�E�L�����^C�|�����wa�������Xy+��"C�T�a��)k��9���}�� b�����)��q�{5ɢ3���ܜI�bxgv[	:��I���;	�����o~�5ᳱ��P¼�$N�Ćղ�7�~AȞ#�Ì?���|�F)����`I�{�|O�T���ͥ�.9
8���ciY�,u/��k��5��n����-��r����0�8��#�Xr�j�:��b�5Ǝs�&����9y�~RM�,�H�c�8��ry�{y#�fq�|[~�`�Ũˌ9����_#R����/�H�sV�,��6pǵb= �2�۽���� ��;сx*n����� cK臒��G%\�,4�k&�m�ر��7���T%[~�mb������lP�+�|�� ����J�㼈��b�h��]�OC��BL�
-n\�FZV�%Ɛe�ͩC<�a�CCaHA㘩�c"s�:?>H�O��P�.V)km���۝|WM@8䞍�5�j����odn��𧠺 �YCteR�]�Э�C�S"��#{�!u8�E���]����aXq�.5�[��4�]z��/w���s���1�$��րDv4<�;�2#���°�-���܌ij9�('}Ì��-��[����S�� C\1�-5P�lM����2�Ɖ� ��p���N<�z[,����Klb$�X�t
.��l�����`������:��u�K��rz��a���t� ����S���b���];p0CN'e��Kzڟ�B&�0�DV�&1��w�#0�H8a�`�p����)�ۏM)%M���g�*�=�����*�ދU��}�[��馤V�6�F�E�W� �7�m�#JC��!�6�<�i/�%�)��a��{�5�B&br�Ւ.-�����kc}�n��)�,��*�G�S���-���dp�3�P���Ъ�<��P���{3Y����"&�r=�a;�Cf0$a�M�cM�*�-�xH�4y�ܐɩ�^�{A��4l��a'�)l�����_���>�0��Ҟ!�}����<Ix���J���3Ԯt�G��s�jQ��u�T'ϐ�u�s���W��{���hM��5��7u�WI&�'{�q����;)4�-������0\�\
Q�� =�ș]#S_ˁ/�4�C�v<��,��M������p�G��\�kNTfg�N��(��(wz	x�����:L੝�"���E��8�	��#���?
��A�ͺ?�#���}�� �@� �5��4�>��A[{<�#)�h�6"*E�0�x����?EH�z������n��-��fd�u�����dl��Uv�+Φ��Y�{���Р���E��P���Эq�� ~���f�V����-ڮ���e��$���:�\��H��g}�a������I�1wT���(��|3#�V�(9����z+mm��=@bUL��17�[~��7n``	�U��.km�S���T\��&��T�=��޹K%�j9���~����JS�z���!�Uh{S�� ��\ƝD����I�Հ�4b+3��=�IS�E	?��h�b��o|NNo�Ezv7 ]F
��!��x��G�H��Ø�yIl�=vjoq˨� h=wT�a���Ab����~���M`^X@q�}�w�|*+�T��MlN��`��s*lB�37$��`S��&z kA^����G	����˜�x�T��iQS�H����JH&/�+EE�?Zh��;߈��v��,���o�w��>�O���)�?| ��|I�����w�s�<O5I���X��I$'sW�;6;�u����e��9�a ��=j�`�XD�kE�]���W9>-NZ�+��4i&� 2fX�ޅ�k5���Az��v��t�QhM�|<��;���}�^3�gq�!����Ƴ2��b�f�ݣ)W�� ���̧̒��paޔ��R�jl�������$=�Z���ͤ�MJX)�'�����'6(K/Q"������*����f  �WB�����З`8���9�ZO�?�han` �E�!Ø|���lw�m����~g:����˛����`1����QɵP%Z��1����#ta�g��*�{���b
D�&������C���P���<`�B�k
ܠ��Y���#w }����k�S2��A#���X5?�c����a(B���O���ew���"o�����#�����(�9��hk�o�&�+w;��Hu0��c/���k M>7*���������������Cw2�NSڮ�w
�i�Ae{�H+���UѮW7qH	���vm��I��&�ZZ����#v�kV�"�w ���|�yOyj��ΗKPW��#�1�W�ʐ
#5UTz�꯭N�V��B�4Z"s�DJ~x��z��Xn�aR��@%Pv(1�](�@n����O65SM��*6�T'���rN�r��
x�-ԉb��,N���\�
�9���\P��ק/Q�!�h!�D{wW�+6ڶ���������N�N�z��E�:V�X�vM��B�-<�K�
P�`n��S7��L�'��m�Yj�Ȩ$ͨ��I��0�0
n<X��C�����(�T:�/�z&��훸w$��w�OOa`�6����!�Q8�,1z>�~Kա܀:���G�c��j{S0H,Y�����Ps� J?~�nC������}�h\�蹗;2�K�dG5��,}�_m�ʐ�i��n�C�Q>z�>� 0<(��ケ�������������fB4�ߔ������h��D��]��*E\��ą���+pB�0+�ُ�V�yRe�޶��M/\�}����A5iͣ��8[o��&��=�Ѵ��x��k���~c���b�t_}C�:;�����j��	���$�"æ�̰z~��X��`�v4.���J�:���y�;v�a�i�/V�
�`��Hè��,b+�9��\5���v�P&:DZ���S\UxG�㟢~z����&���{z��=�lc�F�=�=�D4 `���?n!��X��9ل�yM�PI�6�SD䇁B(�(L�^Z/c6KH�X#d���Q�V�t4������䦦oJz�˚!�H�1��o��TB;��a��À8h�����g�(��M1�`:���L�������S�͔��#�dF��DYl�mgk���L�oL�{�#������r<�4'�"�1�m�ktx,�9��I���4 �b�6�LH]�#�ヮc;�q}(�E���	����X^�ϗ������������ט7JlBbW�#��.Tۆ�%t�v1���X>�s?Pkk�c���	�r���w_��i=��m��������ޒ^gM0�J�S;��ǵ���Ȗ���LAkMK�\������%b	^�H(����?�J�ۼ�������������!H�Wf�k	����H��]�t+q
����V)�O8�m�^���XlP䁌¢(!ݮT'��Zx�%qXj ད�L�v=����������˗����5�*����EaA��L�y�SOq��
7_�I�q(���E����lX��Sx��C���%�����:HB��L}���캤*M���6��۸-oi������_���?��Oq��!0�sA�	O�ġB�<�����_�k���a=Z:o����D��Uh]U��7:	��px`����ت{��l3z�6�{��p�ᷳ�0���Ѳ��Qz�>,���ӟ���kzbu�_��桥�W*ck1���3ߛ�a��p��QūX��y�|Yc��#��������)
�7�J���-��{���N��D3?�I;\~p<�w؇����^�P����I-��/���RigQ�AO8ztO�����ř�������=43�Oc]���>�����&#�ũlٻImj^F�Y�ɀ�u�� wmYS�:�E�$77Jwu��L����d��V���c$�2H�b��_�*][�>ܝT�z:��F��^��pJ��7���F�R�SfI)6QrX�JEull�*&�ӧ�[��a3����&�A}mhH�ğ*�j�X�����,LL=�b��d��@b�=
�õ^B-�`�O������5��j�=΃��df<�67Gxx�kcEۍe��1��PI���|�xT]�zg�8��z ~���aH!�����a���H��	��2;��ڸy݄�X�ġDCJX��3��{Jhڞ?�C�=PU!����;te6�+� �x^����9�Ž��4�he�׿�5�Ƹ_J��Q5�D-��Du��H���ʻfS3��44�9�ۯhF1"�h����y��Or^���bMR�Io��ivg�Y�s62�)DιO��ƹ�|/˗�w�7�.R��U}L�A�?��XF��PT©��^�z�a��f����F�	���۲�Δ�%�m6��E�ȩ�!<��Q��E��ܲi��ȉ$r�/1H�=�3�Ђ9���t��v�m��[PP�%8`�����mH��{��B�k�߮o%�vH�Td5�0ٞظ�$P��D��|mH��P��@�ݻ?���������O����#�*�4��	�)D�jJ�-��7�R,�����?'���~/C�-C�҇q��|x�1���X
�b��1��?΃�*ċa$�{<��J�9�B��n�dx���[��s-a�xl�58łb�#�X���D�&�3�p��u�=��_�e$�c��G,E-Gܶ�t9x�_`D�>�p����ݔ*�!+x�A��i$$f*���9`,����Fi��(�(�Q-�%�	����B����N�!�"Nl�G��u��Z�F������k�G������-.JF@�ݏ��ZK�=�*�\��:|S��e̤%bM�0��H�U���6���R|� ����k>,���<���e��T��g�8w���e�jn�:��<�ր6����u��_U�����K���d����E�j���z�'��ߌ����s��:y`)�ܳ#ט��J�g���N.�rw¤�
�CҔp��q�ԋ8���{��Dۀ^��B�t�Z������;���-���v{�k� Y�-ŵ������q�jX�@#J���/� ��pK���rg	y�kx2T!��-u�_�x���>�t9���.]��`��fYj����IB��O��;�z)���o��@���YcxyC �]352��{���u:%7�H�!��Ir|m�Y�����7�4v#���|�A�C`˘'7p����7SSg�K��O�t/R�Bb��������� �P�kj�D��b�/��\�v���*L�y��+���6���}��UHY��y� ��\A-�,���悮)�n�LJ/58*�a�Z)��
A�ߵ�����Y�ƈ���M�6I�(��IJYBo�����|=w�pg'S���Yi�O����K�Xq�8���˼ġ6P�>�{bb� ��^�	���`�L�v��w�қ�o����R��S��~��!��cp��l+�\4֏Qq���m����h���zZX ecӘ�����I�	8��0��5W��hA�m�',�%��������������I�0N�P����k�wެ�5��!�e��UA�T�ҎMo �"=�1�j� ��N��$���HÆ3<7�
���W�d|��n�X�4;a�����$����&��)#�^o�#�F&�޳G
�8���e��b��B
���d3¨ņg�=|�MmN��J�c��������o^=��y�W����q8Q�e�{�a����-�5�w�tf�ۏ?�J�҉�8;�0&؆H4�:	�����WX�k	�����db�%�Л��C�n�L\�@d���S���|��Z���j��^0ڣ�I@g�����a��:/q4.�d]�j]�����>���|����12vK�h����,�|��+y���^S�h���'e����0wo	�u�B�[�n�fu1}�U7�S�%�v����m�0�A�]�����h&�y�ġ�I��~����m8���́41a��#i��Kdv8T|z�Mj�ς�����D������q'���`l�3�oC��]�3Q��v]�̆TViq
x��=�20��Ы���H� ��п���5����5	� ��w�ƁЊ�`Ȣ��2�a,7C�v�^��r#�ʐ>=똡646?<D�N�3t (���yV)�˹�;�(�k�i~��=�<�O�_��J��)q�g}���cs���P�)��A0ScرM���Y�\����I�7^c�n�(�D/
���M��{R�\�����)"iɲ�s�4=�Z�%�L
�ĺ
���E�t;�
i��n��S�sF�@W#�d0"�5�\K:;p0p-L�����ihP7M��S���8�x�����>���B�p�9�`�
IW�	&�9�=�$^Ӄ.�����B���Y�I��4Ȯ���b_'�k�ii�����f�������i\_�H�_|_�u��{�]q=y�$�
��F�̜�^v�v���X�Z�pE�qB�rb�P2�
�e�+�P�xy![�&����~�s�h$."[�*���f��y���?��B�m��bivYed�$~'���X�?B�0�d	 �{��L�n3�X��((!e��>��B�
/���9�uӓ;8�J<�V�k�g^ۅ���3<�)�N�dƈ�*��ł�̡��O'�Iz�k�N �e���"�þT���}�����O�В���"����AqM�M��m�}��B���h��a�	���� �6a���vzHZ^s�P)��S�`��7��!��퉯0�g��A&���cC���q �v�������d��^�6��Ř1^L,.J����懶�3�x���Y����{�μ��A�{�Aq~��6�r���L�iNN�e�J'MgteU����%?'�1��e0�-�(�Z[�{��p�%��������]W�+�V~D�L��wu���˴�iD��O�T��o�T;����Ѳ_s�-��dj��n���M�f�6keG�N�D��o7������1�Oj���.�+VQ���![� <F�F�j� Y�Y�L�/}$
�������&�h1��]���s�Q��b�IH�⾭D �j��o�ah�nބ�3�F��wؾ?l_/{������<�q���C,�;póp�$9[8{J���y�:�%hf���
�|A�Fk ��{��fab����/5"�X�x�n�\�U�&d��;j�Ѻ��ց��Y�k�HP|a�-��篟Ch�k`׷䃚k���snLd�*q,Y�vQo0"x/�0�0b�����
�M���X�o�$����0S��\H�m^����/f�5�N;�.G�l�hٌ��`���c9������z�[���h�Z*#g;L
 68���pjӉέ:u6�$�7�M�2Y��QUێ�6>U�S{NC�ίA�ݏ�-��Hܪh;���C%�Os�p����]�Y>L!;��g]g�җ;h`W^ҊE�η;���p�u�������J�
{)�k���Cd��L��(�c���k���Ϻdb��nj[{��^��Y�N�aa|��>2�l-��N����u�+��z��Q_�x-�欮��E��ɨ({�*�ݥ��HG%Ix`\s�Gk�b�{�=��s!Ro�ޤ�R?8�&Qc�o\tOq(�f[��I23ܟ��^�>�{�U���,t��\S�R[|�;�+�j����p��3o~���&0f^�����#�9z��U�$�Bu3(^��:�t�S�a�@��{�S����zM;��dX�YG+�Q���)\��s	#��˩��0h��C�8=�RC�+�U�Qq8�������	#�P�|odn�j�5)1�`���Xv��)<����xS�ҔE 0潔�Kw��������\��믌$/ّ��H@'�IG��E��K}\OW=R�ש��/�JjĖ5�O�*�d	E'ɛb������$�	����o=Rf���ҹ��N�T�G��JE�Fsf8�!����3ae�Gʒ�蕔��U"�0h3�S��h�-7�U�!N��W����}-����p(#���%�A�m�GƆgi��m3>��(�̉�B/?{ܐ�\,D\�w���a,������/�q�SrSN�H�c���(qoT�	\p�̥�';aֵٞ)b���+������)�ŚI�B�Mp;��,�[���82��*���F�f��p�pHQ�BUubџ?}�>D4�%��3�dx9�!u�H��}u��ݮ���k�g��-�7;$�T�����8*4�ݐ��=$��=���R�u �h6D��B���ꖬ��m�݈Ra���8̖�	�wT�r����GB5h�ѓ[�'��5�#a�c����b��M�JO�G�_��vۚ�*g����o$�MO7=��i_,#�ݢ�*8��<��M8K�>Q�А�2�� A�5c�l7��&2���J�V��I8�OG�k�.�[j�Z2U���j�>�v
q��kM���I5�1�ᥭ)v���8h����D�Ԕo,W!��/���1+E��׀G�+zq,�����Q}�v�����|�U��uc�$Ai���L2�� o�C�򮾯��B����[y�EgU҈�h~�����OM��$�^a:���k{n4��9��z/�v��M�:dw�|Vg�}�:Z�ؤ6�+��:��v��-��=��5��M��ϙ\��5�y����c���Ϝ��V���T�n'&2ݓ��2�t���}�bzH��>!�eC<V��^�ưԱ׆$��Uf\W���ι�Y1�a^q�BWQyz�[V-���L( b`Ik�F�	x��vE��y�=8�D\�X?1���2OR��ʒW��Ki�@[ϒ�]�vơ�9�I�����e[xS�\{�=�2Jͯ�J��[���msO�����y��>��>*���MM�!>>����j�x��(�8�K�,�2����J���>P�xk]�7�u C�l�(���֪��x 9�k�D���(�f'�|���L��*^&��2����q䱭Jp��pC�ә�X8��7fNy\�XݔĳQ�gu���^a�9�{�Ck�^��f��<Kc�<I���6�r'mWc9���Zۤ8�]db�������&|��!�R����M�k߉�ʓ����74F�DI!N��ajV�d;+X��GC��{�S?n���
Y��X8C�&qZZ��K����`t�_&;G%a�I^$�㹧G:�Tq_Ŀ����=������cHF:R��׾���)�Ö���q�)�o�A*Mq�l{��Z,zF
$I���*i����S$����JϾ�c�����;�a�#�{�3�C&5���א@t�eb�,��Co���R��E{is`�j���e�~M��>2S_��|���Y�]��un	 u��)1�7%�m�N�O����*�lF( 	8
ps{q ���Tg���1x�I�a�@6������B<��;�|p�ZE4fƿ��.J\��S��T<%~~K��4�X$
wbiw����S�Nɫ��ha@㹰/Tv��hn��N/Wz�{�z?�<x6#p~���w$������d6۫��2�뚑D�Yxa��ڧ`�R�r�uS[�P�U&���ˬE'�U���]u�p�wl�֢3��90��tr1色�pMDuؙ:0�K$p�&vC�x|6�<0�s?#S �IH�d��z!6�$x3�ö&$�0p��q$�:`���?�����Zד�5Ԡ=���M�Bl1.��yf���(��a���7[}������w�V�����r��ն�O���]4Fڐb�̓��o��à�����%���I.�������<����{�kb�s�����<��l�i���e�1x�G��a�LcZ]e��"���o�]��:�^T2F,��EaYf�4�>��H�w]#3���o��..��M��� [�̵���p8�� G,ȵ����P�p�Mg��<DSYz��__^;.=�/&����R�zOxYK}J�x�^4��o+�B�k����J|�2�c�"brgm~O%uWXE��[w� Bv��H��5��n)`�y�D[������"���3Y���оq!4ELO!�x����<|{�_{�f��늉�U*-T�#ݪX*`m��A���o�AP�����ǲ-t�gG��%�9�kt�Sݰ�Q�ipA����Ε����X�{B2��j�5��*���{�6���,,���G���4��'��c�ӗ�o�ڎeP� ���C�;ڬ�������a�v%�GT�	�ar�h=�i�{m�''�*!w�oA<&��<�.=wG���C8�~ʱ[h
	�7�1�w6�J���g��kN&[�R��f�~�j˷�}[3���N�Q{|�v ߑYb�z�>� ��Za��4PL&����7�yδM�,�!��N�IwcNT*N���Ɩܰ��Tc���<��&�{_+�G�#D�W�v1�5���Z���/�S1��f�z��x�˚�=���
Q;�w�J���L���k4�QQ
�@�}�o��d ��������	(�*�]��e���ȯ����Z�*a�Z�v��8�ם	��� ��	;��,���uE�39��	�c7��ҊxO�h"��t��*K�q'��q�>�{��E�2����mvr:꺪ɍ0⥲h`�.���pXGL���V����#M�k�N,^���6h�&���l�֢k�5:��k ���;& �Ŕ�x�J���]�kz��!��&v.����t#<�;�ͷ		X���y�9������g��t��F��NX��]-u^��ҙLZ����iQv�&
�$��a͞m1��|�P��'��=~��Z�ۄ�=���u��AV^\ԻfV��k�c��/Sn:׊����c�+<�RuM�yQ�t����ڠ�=���m��4�����X������-$����q(��L,��g����=�R{4r��Pc��wj�G���/��1Q�3��&%|`��*_���Yd��:��N�a�'���b�D��J
Rr�U*�U������y��EF�V�WY�-�e��ΐ.����lb<�B��F��q����6���]8:}2�[��5���k��^M����W�tM�G]g�>aL�>��zLq��5��O'���%qX���D��{|���
����/����v6^������5�19���K,2ƾT��Д�����*5ئ���
A#`�'HQ�_է4֥��{�]����!����?�h����q��=^�א򄭓��k�I�v@õo���%|_�!N�x≁G)�+��{e[ {�5\�ă�R�?�$B�;�u��]��z���������=����T�X}�����̺����>F� fe{�u��#�������f{^L�p,�[�P	�h6&���x�J��{��N��h-�J�5?��^�Պ�!,��'$d�ZvyPZ9��Ƀ͵p�]8��,w�1���I��O���`��yP��q=6�L%�"qٻE���x�'���>��M8�ݍ)54/:���:p��Pv]��6�yPX��n#v]5�;�e���Ν�p����x�u��;k���FĆ�E*�*ʞc_��hbWrAGv
�(�Y+/�Y����ԡ�Ȧ�LX,[��{��"Wt�8�c����p�H�C� X��,������_�����p#D;e� ��f|VN�z�y�A�������i�M,]�^O��7��1n����͝��R����Hj]~,"R=�5k#L�4D5|�wxj�A1��:#ۉ��s'#$]�>x�!R�Vq���d#j��bC�W/i�<��_�t3����_����qa���;y�ʊ��5g1:�x��^^g>E���o�hӌ<G-i]׻��r�K�V��k��=���J�]��]z`�3�L��^�1O	Dy���Ax�`���:%��"��݌�ݦTkzMY��8+u��
싸q.���oӔ�37�q�n���	:WdD	�l���/Un����F������C}|PD<�d"*�*K��hM#y�P3bՕ��(!��Z(��X;�v�e3s<�Q�]
W-���`�/Z�M�u��Y�C��\��M�)s��3�� Q�cѯǍ
V/w����X�7�R���v���4Ѻ��u�����N����o{�2J�$p��eć��bB������Z8&�>����<��R��^����LU8]���,��J��k�C�:yэh�L�]��٢���k��G��BlF�m,��zR��ކ����V�>F%M�x�p�\SݑW�	Wy.�{D%˲�w�����x��=�c��:ݱ �L��UZ���V��o��8 ��/��gQ�,j;rI�� pq[�"�}��d���s�qm�]$���[&@��UOϭ(��:Fu�z�]��w]BH6r��X�p4�A%�s����1�mcFf�	��å5z�W����G�}�@D��������0�K%���>���ޡ�p#:���pPұ֡����n<���c�0P�)�%��xs"�s�C ���LNE{i1jܘ�纬�3��'	�D��f)ECb/7���)�ɪ������������6�ڊv�x����Ա�O�s@��!}y��Q�à^N稚�tr�juF+v�G�i���s9�3t����|����=�-OV/�rvQ�D�4�R���z�
M�+
�Nǣ4<��I���U�\�9��n)>�9hY�&��N�x%���Y�
�ǂ�6*�~(V�!��eS���ZRd��8�.�ܐ��wi�,'�eץ��^jIa��l�{�־�z���$�}fuǬ�2~�V��i���RNnQ��%3�֑���>*�X��].�	�8�X.<:m��|�ڣ�'@�����㲨���YO�.bWV{��v�{ݼ�]1����Sx�oh�u]���lFW��sB"/�&|N=�(�܌�K��C>�a�)�6V���2�+���*i[J�ب1�S�4�� ��A�Epz�9���W��䱚Wno�k��ʗlJ؜x;���.�B��'R���Xv�/����L<��'���1�MCZ�xLK n�*#�B:�ol'����z�D���y�����l�qr�PY4%���
/.]t=1VNK��P^5ܫ»���ny�j_��M�o���
��bO��s�Cz�Wm��ٍ��������Q�kUon%��O�n}�䅈D��`�{��H=�b�됯�Ē���6�C�0���X�~O��d���s��a&5��fzPc�R�+Ԓ�RK*ãɹZ� n-�I���^�}�QLk�Q�a���c��c�k��U�@F���H��5��Ns�#����H
m�'v�u�ڲW	+^�T�^���ȯKdC7d8kc֮
��C�.>d����oE���f���'�;cr<C`�Y&���*<H�7v<� �T���V��4��a�`D���tR�$Ɗ}JW-�ݲ�W�d1�I2�U��|�=�Dv�x��m_�!_��;ϴsh���דM�]3�tK`��N0�4/�	���!��#N�4h�K�/lA��=hĂB�����������RccaVK
��C���d,���b�l�[���g���	K��i7�̸��FE����QmS(g������A���97P�2*jTu��)c��H��H|>^��M)��DL�H���u&��uU;�[⢫�yW�������u��a���r�.*���?��U	_1�z���eY���cq�������O5��ʳݩH-kf��e-�W�z��������,��J�pZ�*^�$^x���]'N�`ϰ^�o�����יִW���x\�����3E�U�A9���������(a��wQTIUb(��{�um����hC,O��������&f���w�%�<Z��/ۊ�|l}2�՝~}�V}��
F��/@OJ*�>�IM.��=v�E5d�����O��\�ᑋ�����4�u�Q2*��a�גX�iN/�]$�G�b����eᬀ��|?�ȼy2Q�%Nil��
M$- w��SY��rR��m�� �sd�a@v��V�����{�YӮb�� I�s%�nTqBu�z\��6��w%�vm6�&jfU�C�%B�m�a���5ծ����llx�7�[F� ��-�?���X�X1�Us�^O�`��\-ڲ�ڶ�e���.N
���ľO��Mw��U�Ȣ�-T�w��o2�J�p�rl��N�:���;d޲��v{J��^�䯖��v��E�\L2�9(^�z�)4f�[G���S���:]!b�\w9��{��.��?g�1x�Kh�^�Ě"�mL,��s��#�X�{���E�#{j�&L���8�4�P0>ꮤ\��6f�q���Z��lp1pYM8W�0�ˠh�&����%婵���w�����i�;/�%Cu��|%���wq�_g���r�"�db(�ǩ�剕�!Y9�)��>H�ԩL�T<�H�왘Xw�p�kS�V=&f)��5���&yb؀�2���C����{�?��I�*K��9�Lu+��5��R���I�&���<�R=��*��Eet��4�0wY\eZ�̅�ǽ�}GZQ�d��1S�g��V�xA������a������9��)�:�L�)�s2g�J�(��^��<����4�Ri�cޗ�f�E�h��:7�z��-*�̵۩rN�n���W��R<��X���1�Ӎ�!D�1�HbfDf8��~'Ϟ�e'����]���N�PP�g>=})?��S@](|	�-���-pO1��-_6㈯62lB��y�QU�����U>��J��HyVcj�t�@eN��	N(��-���1%�����R!�bj׼��z	f��Z���z�mZG���U8��j,�C����z���[��l~W���3����5���"�޸��*<RO�9��r�2IE9���|�<�úg�-gp�Re�lH����:��u�Q.�����$�	�#}s�E�M/�y��fQj�p�5���{fZ���@wI�Q���cV�"��=1���/�ѳZKT���&�H������:�Hx\�����{�n	�A/�ӎ5����v;|�1�HAW��ޔ�R����`Α�|��x��G�;��d�����2D^��u�z�j�=D~e��" x���%�����k�N�a����(��|�kQk%W�6����$�̛�7b1��K�E�:������,>�,��ƾ��~(���b6bP��厞��"ܥ�\2�/���:#Y�.��⸖���qL˭mK_-fRiHb'�G��z�)�e�nkYwe�3=�&����֚��gz69s�`$3�!q�HD��^d�'�f3̣�������&#On�@p��{�f�XE�,�kk3���`eҦ��;��}��p��1�>�o�`-2�פ_i��&kWT�,���;g�&�tà
����
��WKV
!�����cTN��/O�<^�)��������!D�Yy�x�S�c�ba��M+ӣ�S
3�M� �5'��ʫBpư����>���'�9e���{��[�=y�5�1(1�z��]�~X�O�"!�j��6�����u��f[(p�CD��F ��u���V{��H���P��p��|G�1��	=��S4Un��?"R��<�獱��;&|�����բ�QXk��{eK8��(ʜjR覆o�g����I:�WF�r�c_
;&����N>{��7tÃ�9kW?v]��5��k���AM������k~�x�Y�лo<'������͓�Mr3=���3�h��0*+,*P�%���D�T�f�(=���l}�d��SE����V
O�7����!��^C���OT'���y��}����S�L$<Z'l���{QYtZ��6����7a���N�������P}�6���]v�]�,�"�|C^��{�X�_gO�jD��ט�ǽ�/+�w�^��#��yR+�t������PM��� �e����t��a�Gv�k���u���N=��!0Jnr�!�Ƙ��̗m,��s��0�ͪ'\@�J��������)Y�!��J�b�0^ļ���L�i��RĂ���Um�FE��<�kI�a?���!a Fe�����y��w{V�BIOKvC�UC�C�8�ҹ6~�~�!���J�anΈ��&lF�© �أ��k��ߔw�.���E�~MZC��O����6?m����ln3&¯����6i(B:O�DTU�u��j��Zj��N7�4(��oY�k�4�z,KU#ϧ�݄�.ٌ�d]�dc�,�!�p���ܼ�o~W!�^�>wG��|���� wN,5"֋�s�a�V����.K.�ҁk"���Fqz�f�K[6�w�D����+U��4��}V��[3�Ъa���K(�������k��=�p�S�l�a�uJ�플�e[c��{��ʟ����F���^�u5m��c1f,�}�.����RT��#1����<�t,���K.pX��rhN�y�/݋�
�W]�!/�VO�EG�h�R��B��p'ެ�*�&Ml��'�]��`7�$���O��6�N���x��H���,�P�cq%��65Th ��V�֧H���Ed��䆯v��4�����7�bm�4���������1m=S���#�����yu՘ti\pC��g�,X�e��du(�r�>��j��H:B����C5���m��9�W7]���е�ӛ��2jS��r�u��F�EQ�p�!r�T�c����J�N��
sU�hW,��&0�8u�O#1Mt(��c��� s�@w��'�pN9y�Y��!x�8�nW�-����	��΋��a�J 8�/��}�����9U���8iA�4ٻ�G$��v"��k\�}W�Fd���ø�jZ�q�2
�X8���C|�b��J��,�i;���B�Qx��Û�����b�5Z�`�,W�.�!/�n�x���y�0�h�8M)���j��lc�Wj���P���q5s�K��-ڍ�k^K��'v��N�b]b�E����,k�*��h�* ���:�F��TL�����>�
����K�o�W��4�t��H����j(CW��S��J,uPwԙ��W��K��׏zf����ߵ��?ڛ<lCj:AhQ�)��ȯܫ6-�g�?p�CD8���A�.''��J��E�����~f�R��6᷺�kaC8��pmWU�����W�˩�OMF��.!m��C�Q�˪�IFuJ8�%}���Ȱ���y��B���M#�0�ُg����B��rn��}��x+)^P������Ҙ,/h��L���A����A��a�E��n�:�1h�2��V��uM���x��Am-�ā����� �2�J1���TFɲL�u\.0�E%����{�b́d"���k
�Rq\�22�7&�F����6�)�����d 7���Yz��ż阌�A�P�e\E\��k'"�o�j��
tb���M�C1
:Y��YT��	$mG�jH��^@C���)Ա���a��U��*��cF���]Ib-G�n)		�g��Кmd�p)�����ְ�W-_��_�[���-i�-{��%�k���=��1��⃢�qx���&=��n�� ����n���E��y���f�نT���ر�g�C�Gڋ�%�8-ѕRl�uYű���y��)k�@�b��N�v~k��f�=)6`0>���:��瀿PCp�Ka3���>�(=%��3��f�Ӆ����5̵�q�ILS���h�Ø�@�1���>�_�����X`��4�_�Iq�>�
����U��e�x��8�f]k��V��:��-5��e;�m[W�o��}����5��k�I'п��Z�y��01���rUy�"���%%oy0'.W��V�(��[ɚ�5���F��$&z����g���N-�6e�g���$f�N�揓v�9m�
tW��P�ڌ�5��/�{v"O|v[�(��~���Ȅ�@��Q�Z=�Ю5$�����3V8���i�n�>�o�����cӷ	�jn��GZ�@����v�Hca	����=r�����Y%��aEx�
�%�$l���cO��r0&���=�@�o�`dFu���'��d���%��j�96��k?�4���z:��V��O����:��Px-a$�&��l�f4nC��ޥ6[�*&Z��أ�%����)E8�B�CK����ZT-b��\�����،�.@�CׄR^G�Ҫ�M��]$,��l���L�y�h`�����Wa���4Yf�-���&M�5�H�H����T���X�sɫ�ѡ{c��}���=�{i�rkuŭbp-�,�/��PT%���A�ҳ3�)(i*, Z�D��/����WW�i8[����*-ks :�s/�I�2��pT�Jv,��uU��W�������)D ��wa*ٙ�ὶF�WM^~�&3_߼G�gB{ߴ'�$6����7�S��F(�bRE������<�I�GX�� b*/�-TH�`IO����µ��|����|�og�VNJ�"�_�밢�Z�y2����qo����d�{�oV�M�'{�^��]�	O~����jVK^މ>,�$�0<p�|����!N�c������Zk���	��ϊ�v�c��`��Rhܝ�ˑ�YM�Y���H�Q���(�ۉ�*���ZLt՚��_Q̔8sSFo�Q�����j���IJR��
S�Xq���c�(��rwh�=�L�s&9ZCw��W�۲�`�:ו��u��ap�0�>�Ӊ����6'���4Y���)$�6��F��r��[�ŞpzÅ�Z���ƿ��$[(��9VyUf��	2�5��Ŀݣɏ�4὆�%cVn5����z�I�E��q�ZX���HKNX�������O/ϕv�p׋� ���]X굗D\�xG�+mHټ���K@o�Bod{�L`=J��I�V,�R��A����N.���^�x�2s�Ϊ���7cr�|XуXR����~�������B�k���uS�k���$�D3�,�ѳ���DX�_>��:d�߽}������n���g�)=?�z�@f����$���cj�6��!]��'ʚ}F���W���g��:��:l�5��Đ��j%[T_��0����_��&F�A�k�������n��p_&�#|��R[�_����Eq����(H|X����F��1}*{��M�	#7O-L��A<�5��*�}�����\���=>4����߯w���I����I�A��u���[�)YZ�]�m۞ؐ&�D�C���/�m/ڞ��c��?}�֤���ʐ֬�-zK٩�E��^���2��h���ɛ.V	�����$��ca� p��zz��W}��d�J��;6�E4$���=���(�K<ɓ�*�`��A�v���7i��ITx�#-@l`���W� �څ�e �]0ۓ.sS�RSU���]ӫ�CN��4W���,�|O��*OМ�v�2�.�����s��
��oa��1a��&<�ɧ��+^g�Rk7�޷>ܳ}F��^��J"��{j vE�G]�m�5��:�p�H�!�Y�t`�2���ϱ!(�<�QÚN��|��Q��Yһ�BQ.ZH
�b(h�JJk���"g��]I���3¢��tĭ������azc�k��#�ӣ���E�����ޢ�`�I_v%-j)�2�Z��۩�K8W4ص�i��u��Yts�c���_-�	�i��_vk��WƳ4xWJ�@��Q]j��J�PV��T�?���±�rg�M��tx%ʞ�(�67�{�g�A��>��,J�_�����L��~��&��<~�m|���D'��J��9�cj9_%���%�>&e��Z�W�'�-ԛ ��ϗ:ָW�~w��N�K��kT���W!h<��١ .�;�Y�b���O�ɳ)��v�alġ��lQ�)H��1yj�.�$U ���B*��B���b�쨹_�o&�H��MY�� z&����4 P��A�>n9�ɬ�xɇ��b�Q_���%��ji7�A��Aǵ8#��h�]$��R�/
��@:ņ�t����'*������O�c%��]�?q+%a��#��,����کo�r�F�ڙp�i�=�t�@=rb
���ӧd~�3#O��(�|TH���O�FC�C��������R�����ب�k"{�R���kRv{=�ad�P���5�MN5���mwG����ҙ8�buF.i}5�6���^e��W���F�I���W �2�^��{w���P?�֯	�����y3�Q�=��DX��G���ߔ~�!�"]�.�[P�6�O�2�Y�����>����� �UZ�;Ȑ�HSV�B���A�y9�*3���1�>�]�n4�U��Exd-�;K�[K���Hӱ&�����2f�lƲ�Å�UjBJx!{����AӁ���8s	�Un��nA/�	�c�WV��6��]W�|R2:({X����v��Z0C0�Qʌ�vi[�&JO�@�� �#�i�1�Wg�����*�q��:���;[�&�>���#"ϫ��?*�(&�&q8L�6o�rԡ�KU,c�&ޯ��P�B%�U��Huߵ�m�u�Dy2���&��J'Ls(.[���*87�}�Fg�Vޔ��.�V��Z���eؖ�t*�Y�5k�R��;g�>��߱�u瓱�Qz���qI5��H}�Ixd�|��WjR2�[[�2LiN%v�>C�e��劒!��`�]�+�����YU>��|&Y�5���+U��M����a�k�o� �#�͌j�a�������nI.�q@��t,��'N}f�Oi
'G&�#���m#��_�ەr7G({\#�����>W�Rm�.���_���̿�՚#�U���A�5��&��;s�GpTw ��~��.��%s�a�<��Sb*l��Q��[{h���G�w4up�?�ˌ{�������> N����c���Tq������L(�`�}����k��1��Yk��~޻���vdL��zN�ߝ��`<{�]T��Y`��c�����}FC��!9��3�;/���0���]��X��O�iD
\��P4��н��ߗ��`f�f���~�TC졖�RF���Ң�&-.��!bN.�C'��d�mB��
wJuA��9�,������X�;E$^b��f�
Nv7���z�]gע����N@����ow��x#�����$V��T�/��u��ș[�WKW)�X���G�B\�a���YJH��lP-'F��]l�����_����x�2�����}\��vVoX�zK�x��
��kv��0�W��ɧ��:B'̾�=��	Zp�"���D��=�j�m�t]f��S~MV��y��ૌ+>J��T�p!��C�v�]x�"�TY���(|�Gʱ��P+X��.�I�$vk�[f�W~6���1^�É��5qVg�]\	��H��\v��K��b�L]�A�O<q�X�6���pw4��d�W�L]��d�4E�%�ׯ�ၗu�3�{k(�p׵F)�h��|��<<I��\�^��{��o�x�L:�#��R/��nc�'1�eN�cO�X46���e-�!���J-��0?�#����!�[���=��J
X�)�+@Y��X�g}�<^Y�W�_���s��i�=��P8�v�� T�Tn/p'tR�II��a�l�)1�(=,P��� ��Z�!��D����7��L&��o?��'|���}uH�A��rr��T��Ξ3�!�����eb/2�s
yX~m��1�u���`�OYpb����$���=��T�W�*t������^�`�r1�W�pMzT���1�Ga���yʄ����'Z[THlWL7����5�Z���=Fٮ�9չV�ti�)L�r.Ge�5KlT�����h_k��^�"�(7��б9�����u/�2���3���L�H���ʊ�X�"�I��N�α�Ux������h�c�u?ġ\J��u��2����hc~���>���Qګ.m��:>��_'�Vҧ�������rQ@�!���^�4��]�@Hp����j){�֡�g��cm��bm2*���������Y}�H���y�ʂi3��}3pMY� J°W�N���;�Ђ�;�@:�q��7e�[��5��6+���k9���vV�F`�+z�WT�yLT�Q��`9����le
^ʚ׽�g��ݡ�dW��Iz����El�(�KO��J���lf��Q����ccٴ�)�bp�,��+g��,�J������b^�\*��ZoaJ<�uO�C�n�hWҳ��/湫(���+�r�5���h`�VN�sOOĒ�^߮���-��/���<�a�0�Az~*������;b��;@M�lFN���\�SVRU#�1�����q�غ�U��zZ����H*�R�vv�QT�I���hWvE����ʳȠv��w�B�gu�8W�0�/�ad�6����׀Ȩ�&�����%�v�u��`ɚz����L�~8
LN]v�u5ު�C����7��t�����:�g[��U�����r�����~����z����WU8��q�XǕ�A�G%�����r�$�Eq�MV���ր����r20x.�+�e�"�(���.��n|f��n������6�P�Eg{O��3� ���qW���-�V�R�x�N�B�j�j�t(MJ[�
a^�;�F�uX�!h@7ʆ9�����"�b��� k.&:D�|��һ�r�y��Z1�"��a}l\%�\Aey2�w��-ϐ0�1�NQ���խ�ſ[���3�Ɲ�ɝ4AyȄ"��k�e��ϯQZ��\�`b�@����jed�]��k*�ʬ��ޙ�[x��wmw��2K�����4-�$���u��	����*#{�UȈ��jL��~ތכ�S'm�(M�����.�/[�������"E}f�}�y��U��5����oa��ر����7���x'��)�s��V��2�w)�R1P%?=/������#���G��s���;�Z�Sw�z��#�]������ꂉ�\�r�a9�>�k����ˀ�69heB���u��}�.I:g�@}��Noyn����%�̤���]I����T�-,����΅���@��̃�ix�xN�<; Ng$�JI�0f���DBeύ��֒F��	zi}aȖ�Q���>.����Iw���ғ�����XފJ����!��Ɵ��T+*��SV ��g'�M�Ë�ܪ�Uz��]Զ8��%������`h0��y�l��y���G��a�o��S�~a�`jԪ1톒n4�7F��K�͎���ǌ]_��<w��c�S$��zd��h�)A:��;�{���W������*c��rۀ�u���ǜ��������8�=�JeH�O�;Ц�\��
]���h�`��9�a�M�����n`��0���V�i�5��4�4������P�<���V$���&�w�v�2��u{�[����(�"��������҉\7���MhR�W*��XC��v�r(&|w�bp�W
[y�TI5��Sߥq�ڃ�B�-��k��.E�9��Q��64؈c��w։ff��ϝT�FR�8M��5��P�;��A^(�.czc�`ovS�X�Z�$qm�U����MWI�����|�!�� o�vf��T����|!�c^خ�6��C<�=K@)/�a����Vb���l�L���smS����U��k���a��`�H:�X�W�Z��+�w�q�g���;+���T�ٱwה�D�*-ؐ���hZW�{�r�e��өn��;U�R�x����7���|��!�EP��ۜ��4Gq}_�X�]g�� <���,�X�M���/�^��:�O*�މU�z���O����3.�1�u���1�꣒U�U�K���ժ���b�4�.��Na�t�!u� ��s���Z}����=����$?�W��"����Lы���DI6���GTl����/p�_�n-�}�T�I9dg�Y�u�!*���ֱ��$�H�M	���6�-��>fe�Y�r�GJC
lu��{_�NMۘ�FI�P/Ah�K�z+�/�{ZtJ�#*C�^�q���I�H�!y讓�XzP>��p\��Y��0lw������EU����ݗ0��z�g����{L��ue9�׶��>p\��_��ܳ�;wI^�Y��Qҝ0s�!<�E�NF���:�7F�	����WľP4Ќ��J��6肊�"�6PWm�}^��~� �p��3����)!*�NVmYx�o7C�����|��L?��S���ۛ��n�����	����9��g?'n#���`���A�{R�G%�;o�W0�_������z��<��x��5�Ӱs[��lh���2�Є��1�d���(�t8�|���4j�^�ڵ�h�\m��������Wu~cP)���0ŧ/U��Τ���N�8d����x]/5qBos*G)��|���f޾y����R{���?$>\�g���V��}�ކW�\�<�
�'���p��r�ȐJ$�
��0/�O1�0j�-N������~���a3d��fj-PrP��}����N!�Zq> Qb�ڗ���Q���岴�Ɲ7�s^�P�to��iv7��D�!������j׀U�1��sh�&EK\����xL\2*�8bp�#�h+�o���W���Պ}��U��Ry�v@-����x�1[-פW�8�0�n?NFE�'޾�uτ�SR������GBzO�_y/�E��%���c�哆1�I�4��?���ۯi��9���7T��t�z��I�i�ik��͵F�N4��<E�Y��vuOmM2f	+��7��WiFV*�Ҵ�v���n'�Vo`��᳼�Evy	ٚ�lOq%*v4U��Pib ��Q�]�B�5�Nt,hj@r�Gk���9��x���u��5!��D�1^>��iJ	-���u�lI�N�x�yI��K|�b���(������0S;g�"9�z描��ݷ�E���qd��D����^e���/5�p�P)bnҤ}��J���UICL]QW1���g�e�Ϟ�AX?�:�3kG�bm���~	��0�1�`N\K�зrX�	��t_I�!���m�Z�qa���A����gy�c(vUϓI-�=YSC���"n�\���y��9$��B���r�VC������r�����DR����o�h��K-�#a�`�H�w�-k��Ŷװ�0�Ad�U�F�5���_�Sݐ��7���I�I5r�Mo�}I�!����o�H��r�.i$6��wF%�B���� !d�W��J�XP�F�P�����x������C�����Bk��x_>��P>~�(���~����`�<���w��o�-�����trN�y'��YO���!T���*i���fm~���9*N&�V����ph=�K�e~�¾������]D�0�x�W�c.�m��������O������5��>~�@C0I� Lč���+��o����p�DT'>|?��q�I:F�U�0ø*������S������l3)pGa��ˇ�C�Ł���p���Z�!�A�A�������"o�^Q�-�2�~�n��T�O
����ݽ���j��|Q�5���I�I�G;�ų[�pZ]&�H�׆�Ѫ�!8��u�'S��r6�5�kCK��r�0�6l��X�&�/�H���`����������������oY&������{e ��oZ�_7�~��(%=�4����U�����Jj8$���gu_fZ���{N�Y�Qڀs9��5�qwҭ�?io�帑,n�Y�v��˻s���?�ͼso�%�T[.\@��[D0�����lfe� ��p777/�je��e���UOo`5�Y�,��Ř���y�(5��a�nb&�;7'KL�w����n�~��݈ޣJ�!�I�bJ�_�zI�F냒�ݵEg��5зw/������<FC0�x�d�e���׮⼏��6�&�_���T*��?E�80=��yO"��0ϼ�q�wS��{��MNn8��>`m��Չ�� X���Y����1O		�������<y	87�;trU�0��z�]U���\,�l,蜐��g���C���;�֕7�.�����ʅ򼷷�^^���v�f��%IL� �t���J�V��@
]��� &V�E�K��4DS�V�~��q^���>�CFo��x��e`�;��S.K���]��(,Թݵ�
�D�ƶ��ҕ�WlE�ڎ~��V��Ԧ��XH����wK���x��ϓ����ؙ�DλG$0l$�]7����
��fc��j��I�gJ&���#>��]�1��R�`�vY�x�#�������W���^z!�|��ۤ�o^+	�{��E�EY�DOlOa��$���#k����y-hKq�(�\<ZzzOG��^B����onI#�cѵ�eT�]Ȱ\G�bO1��"|��O��2��H1|?I9
�ߑw+�&�����X��z��=e�o��l�(-p�g�wi.=�$�'�B�&i�n
�޸���c��\�1C~�Q�I/QN��w3��O�Tg)�"�a�7$C��A��<���cn��B����&�^/N'�%��L"��:�� J`�--ўa�Ǡ�B�z^����B�s�D�k��m��Ebv����r��1��|a.���8E�-Q?Ye��ps�.P̬�Q�n���Ι��B���{�ŶF��xJ�>/)�-�i� �l#���9Y�ϫ��kv�nW?��Klԕ�ƞ�)�|��C�#Z%S�1�ֱ��|���s��;�;:1P�u-:�?��}���b�.1��r(�&{��}���X�����]���%��������J�Q�&��>|�A�7�n�_�|�L"�U�^��7<�.�X&h�_M�=Cg�?�{)��׺�9x���M���	��ŋ[rH��@z��PD�Xũ�f���������F�'eT� ����`nj� �-=T(*9��y	}?||�>��{��&^ב�ZGS6\��F�U�GM}^&�)z'9�c�;m����a,p�`|qm���J��qz<_,���y��m�S�p���b�l�wN^K�������uЮ�`�R�Dv��+VD��@CH���������SRiK,�:��=�:	f��a
����QYk9"Sx�؜aH�Q����=U-��pJ���Q��!'��{R\e:fC���S���~�]�%�a��p�D�� 1Ίs�����^�d�+���9i
T��E��	<i�x�T���Y�^�-�']m����5:ӐV;��M�l�]�`Xw�܉�-��� ��x�[��!2�S�G*x@��-�gL����#V���SH���ǔ�iڎ}�1�d��ݨ���M����/���M�>e@!j��#���o<Gx����+B��8��n,Jߞh,��?��=�����~/�*���}QB��h@��c�G
e"\���=>V��rC/�~lw�v����,�	^��~�Ţ	!>�s\������o����n۱D �c���M���w&�p�?���'lD!����-�|E)�]�U��*�2�9�<�����#�ae�}�H��	:"�����bQb��@d@�Ї԰n�>|L���W���74·	�s�U��zcvȶ�F�����1Ģ�{����miC�4���A�ݹ#k�tR~T8�~LA����(X04UwЊ]�v=�܎c>�~�N�M�%\��=6�}�[��;&os��/+�e��9�i%B�&g�M۲�7<�� �>ĺ�g�w�r�X��-�'l�7���f F�w�;�99�k��.*�9�:?�y��0?C%���<կ?��SJ%{{���n�x�2��T;�ɑ��"�w��)ė����8���U(� �]*e�s:��Z��C�"����(	�{�����BNx�x��������D�u?�����;>0";�T�םq���ijڂ��+ZZd$zi���?�g����W���d��cū�嚰)�v����.�GD��O?-����IK����!e�7���m﹡2`N+�l7˫��+�*���>2{b���1�_�1%�S�G�X�⏏bJ�C'�-���cA>>�>1����ȧT�A�[��
�7���נp1�E�\�����{�J�jYV�ʉ�����2�Wq��n����pe��8i�xzZg���_�{;;ic�k�5�B� fCk�O��$];Q��	{�L�G�q�%�����wW'	}4A�D5_"�\��3a'���1��,-��l�y���E;3�*��D��l�y|�q�V��B�)'��J��-�X�\v0���o���6[�s?�~s��J��.�֢��~4��B��T73�S(�7*C�wm�1أ*0� �W�ccq1|_����_��z����aL `wL�8�8�F�=m�A��&g, ��Y[s����d�g��q�bl'�1f|-D~OC�ب�tՂb#3�D/
�Ft�Sb1�}v��1)�^��x�{�͖s`Rky#�f�&y�H�L��Ѝ2�0\�7�2��x¦���^�:r}���%�X�G��~Z·��i�F��"�!�EE���hl:8>5����M�Yo>+q2�ksFXk�� �����y�]�xo�?y3�|M/C����Y�;�1�w*�#x��B5s��7��u�y/��:X!B
�˙a�6� ��5D���{�C���ыж!�=��xraE�(i2�p�po�4MIf+Y-�.�"��T�"��!�u�"RD��xy���:[_+��F����e,��/�Ϥ*��_�;��Z{c�uf�Ύ��w���`Rt��~uU��^+Nv��`�_��l2o/��Ljxv`(wg��2E�,_#��f�ey�K�i<rM��7��_:p@y�eAX����;��y섛�����L*OOr~�r��mf{��J�um�3�aHʈg	G�݋.�� 煨�bD?S6����cj̫�"䑞X��ǻw�;�K8�٬s)��$/��KдC��F�&�� �o<Gb-=/<؋�<�kLṹ.z����y	M��y�.x���=���4�i2��k���8����n).S�԰�F�X&�f��5a<��☙x��mDfYZ2��cz)�R�+�[ݓ� xa�xi�J�z��2xrH6��WQ��S�LNFS�
�B��gr-c���2��U��GZ�\���#��NRTV�.eCz}M)'�T������	�����T��si�.H�,kВ*�l��nV�_��7��������=��h��8�?<�B��Dty_x��n,gv�s]�o��1�&'�����GQ�Ty˓��pܘ���7�2K�b#K�)佨C���B_�ÌZ����X0"�u!ϋ�7d.�0��Ы�~�P�q���<��z��sm7��Ԙ�t�=4=�K�7N�F���*�ι�f�,b׵�E�e���$2*�_��7����EL!�헋�UE�E�^yLMQ�r�Vx_�>Ĝ)�ӻ̲�'�w���r��L���dZ�9��A�r�<n�ϕc� ���.��!�����E��?��k=Mj��j�*R���M�w�^�g����ѹ�1�xN+4O9��b�Xm�}Ӛ&��F��_Z�#	馀hi�4�L��|��1^u0��|s�6m�i�N�R02l:�U^W�t����S`�K�����쉖��i���K;�Ͳ�;�������{M&��w��.��09�AF8��M"N�����!]#�O�OM�XG+%s|�P�#ͦU��E��SЖ��!isI'��u��P�"�'P;㚝�%����i]����*_.�A��""�4n�5E�������=j�#��Q�Ѭd
զI��U^�|�.X/� ƄP�z��H��
!*iR�J�c*�p$�e�ƺx6Zt+��]c��n��Z&���a�?�����_���{����{z��5y�H����d�Ԋ�c���<-�� ���a����
s7ߟ1�Ѵڨd(�.�Kѩ���;����iP��GF>�Qr�z���<����������$���-��)�,R	ׂ��t�!A�k�9wI8��KqJ�~�\�܈Q�	M����/A).wI�z�[�SV͊�t�x�!&ݏ�X;�<I��.��g�ꂻ�� �S�.�a
WX�z�;�Yq�}³�8IJR�"5�$��F�{�Q��E(��}�/l��m$����5MW����gc����B�-���1��a����v�^�D���� C�
$%乖֨nP�kL�nY8���ь�s�lK1L���F�x��` �%�p�4P����}��t�<)ک��[A�gM�$���N6�5gj1��!킃��&=!��4�Ԣ,u�g�h��0�'N*2
F�$!��0<,=]�yw����FS�1P��uC4M��@X�����I�Y	���:K�����7DR
�������_�i����p8�-���B��$�1]2N4R��Y������?��H����].�w�Ȭ2އ�p� ���>�cj��9�3$����� ��p�����&ϑڸy�0O��r+碞�� E$�Y1��̶��R!�He�EoL�18��\ٷ�Á{ Y繶nn-�<��@c��X�Ѐ7��\Z��^��Q5$ش�1�m�3�uQ��t���K�F���Bt�ק�V:����P�:2������]����6��o0�/=��p�@%%a���nc�3xͤ;���	/�\J$<���=��Q�͡1�F��e֏"Ja�h,�p�2;��q�����ͳoS�Aۅ�!�ζ"�z)C�0��`����D����I}��1Z��Z�6�͍s���4aD�!�A1�Hq��m��D!p�Cx�����E�ۻ܏�c���ӕ-�8@�z|�s0�i*���ď<�˘�4Y�h�n��JeAEB	�o���x�2����i�x�;����Hu]��t�^<ʮ#i$B0A�}
�(�t�c��'])�F�*C]|GT��﮷�t'+�S�S�Im����;�����F����*��+��S�%�D�/�Br�O}Mycè�[[�S���  ��IDATPYe��h��(;1L>����� j Mlw�ˢ�c�
8?P��i�P��>VGU�U��1T��WٺK6��IY|9l�i�b�k#aZ�;��R���Ą1�<R�'9��LĆ����
����S5��l�$�s���C�ɆT�+)����R��\e!�����`pQ�O��U���z��J�[B�.>�Lm>�%Qg���h�E��7r�����6T�����{�8��Q*R}�<do��.��&U+�QB�H�4�������+s�rc��n����+��C���Ix��1�mh�<!h�/�7�Os;g��CC�-w���i�����Cђ���@"������s8./�H"�l�e�A�ܯ��8L� vL~�7Lz_KA,WG�a�yN6�l �5"��JMܤ.����g��ңmb���عbsC#���r�y5���)a�pV�a�jf��9�?)�L�@���K��Q���*�)'�\����<4NY&/�h";�ceg&�R, Ǌ-r�_p�\UUY<�<В���񼦚��\]y���Q@��t��UrA�RdQ�7è�NX�#���\~n(���~��=��Տ>=3�_!����_3�ƭ8.��*�,��5��h�4,7�B%���e�:��ء��1ӂ�KS��j�I�T%̬~�0�c�cp^ �Ls���[0h�2����F<D�RS7��N���2�n�^�e �Cy��2Kn�����e��FoM��y�<E,����\�&V_���$��>H��l0ɽ��Y"M��%�x&���!��2�����h�����C!����j�2E-{���)A�Wu ��y{sԝ�Bd5�&h=8vo�d�%�a�T%d�ם8/A�K���Cήt�uRr�)�*�����̕]pIY�f��eq�)Z��#h>��4bZ��
��C�����Q��%������cN�D�h�OA�p�P"7*Ҕup�	y���f0�_�����yj����aqx0W�~*Q�γ��s0c�Ic�� �E`�e���ju(^�`-�]�/ �#3dR.]m�ҏ͑H��[��ײ�_V.=���{@��D�3rM��4Iy�4	�^�=�s!b�h�	��!�X��vp	f��c޻���r)����:��>F��Ꮼ��*��ց��.o
���X��OcU3�(/d�b�뙮i���l�H�mB�t�F�'���Q��l��>�0��ȕ�-��J�c��X�zS$�0�0p����:)[�!#	zh�f��,C����TBAD�aB^P!�c��j���BCm�%�6�V�9�t�]�O�t�u��G:���:xR�����KR�Bų�u)���|�U����������S�iˌ��j"q%�PT��[{�1��pO�㮚j�҅��^e���H����"�@�
a�ŧ���6!w��4#a�D�Ou��,�s|�b�s�����]y�}@l�g&�wxٗ(�H3ƁT�h�q	��y����D�C��Y1(��lt}���x1&P}�z�!uCL'�0?��i�y��Ќx�)R�e�g���{4M����C{�S�*>A��	�H�x
��|�OX���/�Z�o�ʕ@�020�o,��KN&�Γ��N�v����YgC_�@0�����L���sL4z�{�L���w�sD����e�m�<�<>A��Y&"����B���Jэ�^"5=�>iLa��H�� j� CD̩����kc*P'��|���d=fa6�^?���1��	���af	�"J�`Ԕ�$��~�w�oB�c�н_�S<E��0�i�^,�BS��2yPG߭���|�N���x�00>���E�בOc#�d���&�Z'��k�͉�)6�>BV��8���x�S=���
%���7��|�??���it�����=�(�;&h�I��X�#˹4��ײ8�c�^�����)��󹌻���	eVMEx����d�x��[֭�t��]$�����׃ǣjXE�%ʙ�F�+Ӿx8�W~S�Oבy=z�oz����3��69;��A;]��^X/Z�n���@�'�j�M٧�ꬌg���̬i̝�R�\�D�Վ��x\�i'G�F���\V�����	Yw��7����5�����8�q����Lc�p'K_c��+��[NkVbWF=;�c����&&#��6�Mn�V���r4k�`ln��{���>��2�i����֑H�a�4���[m��R|f���(�����> �3H���G1�i,1�������K��^A�qoY�~����L����N�����)B7�{w�|A9DWRs	��ep���7�T�L��箊���56�ɂȎ���"9�8o(�xV?(���:�6��q���r8P�����Lرtr��,|�A��������R����e]
W�̈+,5���{{mug�����&Z��R���qiOm2�LF���&�Md�\L�w�����zw;{���K�38�)ڀX���w{����pw
{�a�c|.�z��^�Q�8Z��([��Ӹ��i�d6�F?�������8�ӕ!�������m�x��%+����U;ߵ��m��3E�e:-7'��I�\�C��"�]��4������_�_��b��u�0���ls�=o�A"��8�2!`��OU��>?��+{�\ΜH����B`g=4���2�P�R��Ezё���x��s�XtQ�G�q`��JT� ����a�~��0,��I��"�B��,)�O�/�%��U�2zq�0��p�3Ce{��̩u��y��p+�����ł�y"C
/_�u�lH�4��(�u)�G��U}���[.2(����y�P�8��>)ǿ--6�����0G$��ݍhW�Qv��L��d�`8Pi+��j�"�#̇��cA�����~3�w�$CNY;u����9����p�b�Tk�-<NC#��ǵ����
�w�tn&�%C_E�ϩ`��s^J97��.��8.�+�dEG��$�2K`��M��C߅�9�s�J���9�a�ٕ���SXy�_rb�3������<R�dʡG��P�QKa�KX^���b�V�̸�B�C��R��Gw���u��U�����	c2�uj�jX>�x�w5���I/�!�7�YO��`���׭<'R(�������CVW��T����CJ��PEb<6|?�x�@c�a���dC����V��^Z���.�7��L�d��Z��g!H�5���nh�`��3<��������{XD�w72�n�B�c�� �t��3tP�R%���>��ݝ���x�!�b0���E�H��d�ժ2�߈OyD/���孳�l����ȱY�J$3<.�#=lR�[��<�)�����U�N�,���65E�[�1�!*�MTx�0�R�zAhO;M�zMS���Mꜙ�Z���A���E��9a%��"0��0*�e�+�OB4*�<��������i� �Q��ې�aV���٨;
�\x���4�ٌ'�/��{�W3)j��\��s4�d��9o�H8f ��n�4��Ɛ���E6��RTd�z`�ƵJ��f�pF��0R1:��o.*S���ւ�4����rU�˽\꧳v� H^�e~��p���K��]��UY�%9��#�<�c���a���̽���*`����g�_����Q��91g�1�\��5�$�^�]��?ޥ�>.���2���q�-�4��<��A�Lx�sN���u�9D� vn�;��̃�B-;ڠ�F�#��\RM>#,<#�{�5�?�MC�ȋb�eW�`Q���㑑E����4l)Zu#I!&�Q����q�g§x�G%�\���bPV���1Z��>��I��UpsN�\Y�
8��g,^UI�W���ߩ����&�A��`b�U�J���>8Ņ�g��ھ�c��QZ�iZӠ*���0��̥�Q��sc���c�.���=�!��[.ǝ��yV���`��R��U���y��<g��{�F���}�h�n\M�*���q��_�����WZ����<�v�yҫu��-�Q`1Ñ��դ�S��P` $�fS��
����:�)���a��hC�:&�0��.,�o���Z!��0�0�W�މ���U.G�Am"���>zѻ?�To�?���%������5������bpc
"�)����*���O�6�f4%D`���oC?3�R���Ӂ	�!J-ɑ$��z�&��$���>�M���v��bi���%�י�ۜÐZ|��G'-K�ɋPR\^wauƞ�ߐ�{x����_����)�u%#�s����Py��a9�{W	nq�iT9�Ӽ�}��chx�Q�s{��8�J��� y�G�NP�'c$xԗ�<�Z������K?�]�E�����D�AY�s��X|�B����K��_⾫
̎�+��ؤ]԰�뷦Ja�\(����*�#^z�J�Z�.L�̛�%����N���Wخ��X�^�(���X�,��I��.����*��i������ў< _��]�K��	����,��%g3�����C���}��c�bOq�=� Q�=�߇p�<x"�'؆We����b�1e���v	�_�o�v��+�e�n�r�epD�j��ۢ����!O�,�?JC���.��X����+/�\���X�������>!�a5˿��	,�3���J����gE���IՎ����XC\ML^�]l,cL�K�6ɭ$�q�}��bs����h.JD���OJ�IG��J����P����4.#t���S����P�s�MGx�e��D&l.��c3>h����YO۔;4�i�(��oZ�)�ٳ����q\�B�4�Q�����Bvo�]v�9!��%�ߚ�,�,8��;���m$^�����U����1oǱ4�:�ο��(�E�-���t�5�Xz����`����$[]e��Y�c�{l�.Ӫ��4]j���Q����O�؎0� �`�VT+���t�(rF����M�����.�uhoRrex��+{�2��6R���Q�kL!a�ɜI�jBx�m�&C#�&N^�����97A�QT]t�mצ)��Vb�x[��r��ᖎ�:ވm���I����ي�<��V��x�������
�R�!��?�	���{�yb��q]sg%�A�H�*���/o�^)p�U���h̭� Ɓ�<ga�j�r�Ha�mw*Br�A�����#�7uE�L�_�+4�E�t-ˇes���-��"ه��k���n��,��D>qL>}����ӠO+�}V�
)>-�s>�����te4�mw�+x�z&��!���x~�j�Om�S诺�\��}�TIVV�r�Q��Dx/d
u�50��<u���FW�F��� sa
݁N��S�5ݪ�kz#��鄖�:�`]'�JQ�H����B;�\����0M=y���4?�4��>�{��I�MS��S���9������ƛ��s���I�%S(�H�]���.(N���y�P���8N:����ν�q"������jǻ�&pdH-���q�����W�>Ϲ��jF�����z��tYwc�^위1����%:`n���:g�6udh~���RA��S���{��-E$��q���5������C���O;���&}����}o{���s^��h�*hx��r�~�9W"ΏS6��U%�S���u�僙>�P��$Oq�po�\l�+�6�ʀ?�?����1�pG�+E8��-e �r��k�_��K���.�/��Nm�QE,n���J�޳0��z/b��%��M��T8k��������z%O�x��X���ɵ����-\�.=�pJF�Px3��S�Rj�ioiHk�w1~W��I��ǣa��lW�,*�v���*ڥ�N��M��Ѵ��wb��#��1�wu�9vWu�(���o�i������Ƴ��<�aL���đ��&��� �k�ŋ}�o��ֳ�d��ܲ��-C�c��`�L�c,tL,�ﮌ`�C��ϱs��M�@�&�q�x���� 퉕%��`Տƥ���\S�N�R�*�m�~���s$B�M���t�s�����-.<�U�t�Nkn�� ����6�+E��&�W�bN���1��s`K�g<�D+Q��	^5�!��E�K�@�xȘ3�迅�ۋ͛�)qxJ�H�C]��@�(]'wh�v�N����H��P�?e�-��Qrj�7y��zOǌ�q�-�#�s�,���S����<��m���C�����=���2�0��N��I����r{�Ґ�'e឵�Ѷ�ڷl)CXp���Zy��C���(
�C?BUfk�sa^J���6���+�ި�&���$���7��4�]��C�omʌ�&�_ӳH��(�((�d�d��9�%�RN`{|�6�ŘV1ͯ'�j�EO쑆�i�������)�5�!�4W�����G	�L�,<Ҩ�c��0f�4Z8I�=�"w�L�r�>�D�H����JS��L�m!TYGIh H���92��tc�T8ڊ�k�T'E�w~
����xۍ&�.M�͑�-B��-��>5A�A��]FѲ����LVcf)cg&E+k{ɉ#����a��-A9�v��GnX¬.U�Wi/�_�s�#�~Y����D�8�fv��<n��\�dkJI
쮄u��Q�O);m�V[�wӯ�N�C�Q��DT�����"�e> B���XL����k��VM�$,�y���?��ۉ�9���Բ�]p>*)�X�c�ZP����;U��8A34��jf���h��Sf���<�F2��D�L�f���$3�Ҏ�� �2�`�^�S�E�zHQ���!���zu%�E��E
c������c���a���R�v9Mynφ�lc����+����.0���ޣ^O�!�Ě�,n��]�w��"�!`C ��6Ё[� �N��Cd�Ι����H��@_��^B�b ���XJ��'.�I��{�}�*�p���qno��ciQ��YVO�;X 0�02�(cܚ(�LA�bM��vx��!�ҩ�N�+�ğ�wJQ�\�
�F��p�ƃ����ƈ�u�i*��<ct��""�8!�va]{y�YuW�>M�FXS07'?��!�W��w�D�OA���:,�x�	>g��0sq'ݙ2�ax����H&�ޭ+*�*�FB.N:q�jC��}s!���J���Q,�?ERF��"�����x��z 06��U"��9r	1gm4ovQX�}���ǜ"��=�K�S���Ӛ\�m���_��rTR�)�
�1w�����>�{qݻ�8s�#Ā�Ԃ'r,��S��ں��(A��C�W3��x.$#IĎBA����UEh��
��k���l�G��Gې�߬�5��1[��6�.��]��.�]��-#Z���"��А�dH1p��C�%=?T�DX��hCQ��M�ݴ�0Ȅd��W��E�3�à�$(���;���w̾��3�y�g/Q]t��]������2˸������e78�]܍+���������V�g鉎F`6ؙ�R��O�����
���a2*��f�9:��t����j%��+}W�����l�Jxh}Ty��	�˘��)��-�h�G�C�����)��Հ�_&='$-og�G��	R�tZ$A��1ۘ5�ԇ`��$7���Աm�eU��S��1k���.�N!�܍y��%�;��c(��Qv9�F�l������^ZES�!{��(ヾHF�I��El�۶�p�3lP������lG�S��W*��<����%���L9���=J�����؟�'��#�Y;��r>.+55j@⊘k���	}�6�Բ�G.4J�5!�9u���U��X��}�~.8�1H��1���7��j��Q&����f�������b(�ĂG�`��q	��A���$ٷ���T�<��z�y���D�>t�:5F�A��Zp�.���7�~�ԛ	�Z�����ڻ68�dkN
�y.+��&ZY��-������&T���m\W<���RL�6x}���Y}#f���K�wT��7���snr�!ƞO��-,�n+��������s]����fڎu]	I��]L噊�q>�+��w���&�O�9� {)�Der�*n9�\y��'�eG���#�A����Vx}�ы����H���ܠo���͐G?i��gvy�MO��Hs��/C�����*��Sb󒶩� ĭC"�d�K������͌�	7���b+�/�;���b�_T��`pAm�駟����Ɉ����[k��1]6��@7��_�.Ag4WYc;��V���YI�ψ� s&�A��=������6��f�U� Rrɕ�Im"������k�����cri�@���c/�	�I�[۵Z����ҩ���v��`��v"���1�H�\i(5�B��Zє_��H�p`2�c�%y�Mϛ��x'��(t�j�kgWr��]�ͺoU7ѠEuap�՜�ؐ�ĢE�:��N5�E��sS�4qLMS����uZعWV�G3��6�Km��Ԅz|5��89y��Eg��,�.3\J\����>f�i<\���
";3�R�'�����1O���M�I]��d�8�56w�F�DjVD;�&YR�j՜J�����]�����c�x��G�#�@��jm[�0��5-V,���aC�d�\��	g��ɛ����E����Κ�N������]E�_5�ϭ蜾�h���/<�"Ag]AS�ܒ��i;����񯺎5y���n����q� ��C���.x�ێ�Aл�������d��ذ'�D�55�/ш��=��ۈk ��������Ń�ڵ-�xƸ�q�F�q�Š�)p?	�����H���D�U�d����7V�a%���X��~��#�߯Cp��J�����3A�����a������k!(a.e҄6�����U���ݠ#>��4
�a���x�nn\����|�}��e�Z՜r"m�7<0Y���>���a��2-J���]=Y�@�@�t�r�l\������Tĵ�%1Ŧ�W�K��=���n�E=�sn�33kL�����C_3U���f��s$��l�8�!^2�ĸ�a[�E�5k؞�&w� m�1�]n�"�2��Yb>�ʯA����!�\ѩ���]Ń"�i�N��N���x�Ϟ�v�G��+��kƔT��x` �����Aw���lXQ�ʒON�[���җ,F�&2C���τ�,	g"Ivg�t}���>�� ���vI��dx~��I)e}�r~�
�N5�h���<���R-�k���FX]�*{�����/�B��xٓG/��0E�ᄽ-�7�bFQ�[a�ؐ�������!w_mKF�<H"��7@�ݶ��Q2����������	����ڥ�%Qg$�.ޣ����\��������� ̩qױ+��^���><`c���~P���xF8d������1zw�o�&�Q�1)x�NܳKE%qe-�92���W9�"w"f�K�$��M�'^c����p��v$��Xc<f�k���6�H�vc(�[ fb��.Z9CC0{r?�g�k]k�+�j��N����L�gf	=�i%��0��.�9a�-�c��~�1[���o�C�6"�E	$$Z����ÑaC�n��z�l��T��\IԹIW٭��]�^@c�O&��x˲˔�̟𨰁��[���6yq�D[ʘKJ��c�X-I���a�-~5�OQ�}���8Gd//�>�(]\�!���h$�})�zr�^�>�FuCW���"�Ι�秫R֡8t���<)��H����5�	��/�Ƣ�PJI�3����Yb3'#DV=��J���Dω	��<���#`���x�!�3n�ίg��iL�x?�`�E%��	�q<�E.w�+�c�s��3�0�L:�e�~#�~^�!gx
������H_Ef�FS��&��V��`��jYG�F+� y���S'{���K�����1n�}1�p��T8���(q-�f��]{%���F��K$�앚cZ�%23V� jP9�n�##��Umflw�ƙ��N�`�'��g�V?Ex���髏9ciM����:g�bfE��26�%������f������5��Emrn�>X�N��6�5�W�켟�����Rp����}��榺����B�zƃ�	��VDo�K�[���n��Kf�+~���W�����X����c�x���y����1�6D9m�N�8��g���&O�K�g��&���}`���NA��=c��������H@A�xp���C]�>�C;����8WX��fM���B��w��n�*��� ��oB�%�=�u������X.+� H�f��Pk�!���~/���b���!O�9��	:a嚣}�U�6�@��C����2JB���<wBQ]��y��w[�:I�p����lQ��F��KKn�v$=)���ׂq�8��$G{�Ӝ�T�-ojF���������&��6t�+�S$�Y�����(��Xx��K��jK�?������9xN�G�*��q*��BR���&���5�����H�}Q�PL���ڐ������n�V��S_0'�R1������l	&S�d�Px��`�Quò!����U�h	��Dٻ')���ل7�C������^����Ի��g$fOS�"�>�hbh։�9�D�¹K��;�j��F3g�YN���]^�2������uv�����d���)�9�ǁ^cD%A�P�K�%5Xӵ���YGey|�D�#�p����m���H��a�=^�sj��T���̖"ژ;y�h�����:0�&��C�ҜY�*Rj��S�>o�K�������۪��gET�����X#�Z��V��U�_M�������\9B�H�1h^M�rv��&*�v����+���>�k�u$}�/����ӥ��l��S������� ��[q]`�Aߪ˽sR�+��rKDX^��}n\+K��i��~)ü��Y�IB0�!��:qh����-Cߝ;"��g�	�=ɶ�H��5Ì}����N��V���9��0�]���n�j#����$]�X���\D�E��<�x.?���+�6��A0�7��OgC'aܾ�*@���x�7o�r� *��,mă�XM�JR-X�Dr,��Pܙ��Sag�0��e�V9�M� O���iO��dvAln+D$L8�S�n���7�~�Gc{�Cqs��8�1����H|hvƽ�8�C�ŷ������H�f�3�h������~FU+���׼Y�sl��O�{�H�Z��<�ې���p�E�xP.a�*;T���j�f�-|����p\SzJ��#�t��Bg ��k��8��J�[%��}��-Q���6�.wP�XQ�7���bH���1��M��%�"톈j��~M�p\]��4���L���hx<�`wr4���*�>�/���}֯%}w��ژ����@��y��l2%*B�|�eeꨋ��2E�O�|�u���9�}����&y���$m�%"��+P�re��̞&B]ݤ&9	bH��%�W���I�,	��U"�U޸d�j���M#TQ\ͷ��b&����v&)g��Ʀn��<��s(��`�3��Ha
�!k���)��U�5a��ish��,T���nB�x^󜮼Br������(=T)��0pq	�T��>ۖ���R<���7��O��*2��H �wVfB'(;T�jRM��XƗI<Ѷ�`a��)������;ww7���S�=��8�J's��:pe��HV�P����KV�z���J �kC�(�!�4孉r'���F��v�2�&0w�+\�s�)UWT����!$����N���M��^_D���K�r�g��!h��z��)�zI�����]����[�o���㻹a�A6n�.��H��{��1��������"��U5�<8q�{���1�Z�#4܊������w+$n�]!�w�C��V�!(t-ܻ�+\��)b�2,��y�İ^�� �EQVG���6㐙>��U�L�`4I�C	�mӔ>rw�B�LPŐ�,�ۖ�hO��"ߓ�/f��}`����y����yr�>�36������Ԇm���G�?�o�"��¯��Ǽ��C��vT�VA�W�>C\m+%|���h�7C�%�`�=��FmP|�y,d�CZ5]u�]�C���%��V�06�HN�{����͖������z��WB�(:�ΰs��T�����!�]�ެg{8ກ�tY{�1��x���~��ni0ב�f���O'��Ԙ�[W�6�%
��ę�h�<����%��5��E��-a/�`r�7'�,�}E�J)(]�\��D�e{�T"�(�T�jDdng���Md�o�K��ό�@\�sV�n0��ۚXz{	'�����5�4l�37�:B���^)�Yk�/�����I)y�hu���̮����jr�I��B��d1#�$t�t��q�;Q�d��|u�x��P*�/�C�L�mԕsw%���%,1xOؠW�pN�Ñ�ܱ��kNr�;��7�R��S/�Cl0/�^�k��[u#M�N1V�r��1�"fS#��0�?l���Tb�fo��Ʉ�%`����7V��:C5��Mz,�m�]W�S�#D���}{�?=E�M��I�+�7��]�v�9!�ǜ�8��a, +��f�jbc���P���4O����q�)7S`ԋ�r����b��2uY�p�&�t�M̑d��~�aĿ�!]��]tW8`�X�R
�������0�>��h�4 �Nv����<n�=����mx���KT�T��m�zl�\���W�M������Y���q�;EC�/f���x<0G\>�Vα�9���Q��$e�.ӛ����l��f�-C��ک������9l� 3X#�T%�W��z-fu�2���������4�6 ��P��I���������8��8�>v��>ǍxZ<�6��P�aHD|������յS�$(���å��R8��	����E����R�a��zHw'a��A͸<�@��͆�Aoj,�)L:�ډ�P�	���#�����o7�Øܓ����fW��7�M�,X.�l�\�Ŧ}w�93	9�P�Hno@���)&.�G�)p�.2���w�T�j];b�nZ&��2�諒��]�ʫ����-�0�l�r��.����t���@���K������5؟�չO���H2"<��|�jJ��i�$�x��;qbI]XsS-$���훷�j@��
CJ���c��mN��������Q�-����j�����Ԥ�%��Nz�f$����_��-�S�7b':sk�H��#5��v�Ϙ�b�L��zM�_nC�"�#C^!H�x�!0فg�Z)j�"�ms����yNn�Ҷ
�aH��g�q����̌��!3��� U�deE��_�u_㡳�|��/���!\З�K����l�r'`$����^<!l!%�G��
��/�!/6y�&�G�ʈ�NIv�o�h�9L�6�+��i6�H�r�u���B#�	�j঺��ۻZ�N�������Z�QgsK���E�4�:�xOH �,(ã��%����ڶ���6�x���88y˄��v�LB{�Wl��8���ڸ�Ɏ�\@Q\���%��:o�C%�p�ʺ#tfk��Õ�;��pC5Z�����D��;���6,�j���?�tSDT�m�>"�p���v�/2�(?V��h{�CUrd/��c$T���n�4����v�>Z���Ŏ�Z[���li�1�E�0@�C��0�b�,�b�Đw�r;7��(ڿ�������A�2t3Ny�?�K�]@s�>8�a�nK�*ZS��)g͕�*��5Dk���z�Q��d]�	p��*��1:����ʭ���8���=7��u������J�#��ԔJ��c��iﺴk��dNaf
���!���<D�0��=�7���;���V�Wig��2U��9H�[�r�+�RC]��_sQ�0n�%�r)d�����k�ׁcm�˅�W�h�����n��b��?�����)�=S~����m�/!w����K/o�to����T��K�
�.��|F��������}�.�+1+��M�To#���J,(��]"���ϼwmNr�59�B�ɭ��jD(0����e,�jV0�����+;v�c�YBN1eڊ��P�W��\�"TBC��������@�Æ�^�yI�0z*�����͎E�{��àc>L���ެKrs�̉��3��1��RlL��Օ=M{�b�
���2�R�K�V���!�D�%A��p8�y��T�����K�z�\#���n/�T��g�ț�߷U.��rn_�Sj.Y}�y�*�^�MW�9Z>t�����~��lSR��PW��0\O�Su���{�1dC�e�|iy;=- �0.�Z;Ĵ� ��u��r
N|�S6���esά {�;N�m6��@�>�d6�颤U^�1*,��lc��<�*�QdZ]RGjɬn�۝zr�Ӑ���\#��Ř��x���U�,���e-ry��L?]�Ncľ5˸���lu'g������zu��`���z��҈�_��62�T���2޷�/���������8E�\S��s_&S�Q��gx�cb�������!<�B��|����g%�#Gt��\ "�$~$�����|3��%�&��я<ɿ��s�I��,�#�!uG�1".i���]�w{��	�s����z���n2}�1�.��)Fw]�������K�ٍ2���M�,�!E1Fx���͜rI�;ǣ^�`���p[�2�`U�wj�8_R;?x0��XG�S��Wt+p�ϼW�d2�������霍mz��lG�lb1��=�~��U����}@���Mh�9'������Be��#��;ע&A➛���
�%$�p�L/��V��'�����x+n���Ԏ��SZiW��s�Xvu5QFX�q~�
�{�X���P`�W�7��v	�N��m4�p�/��9���x=Rzp1�ct��VJ��e�����ĕ�*a��<�����y���W	7���4�QE��6��N˸��.s|e0T5��nk����=���P��9G��[>�nJ-�Z�9���ޔ�8�t� L����y���ٚ�:�
/W���%��h1��@��1���T��I���^�z��k��[OL2��`_��=�3ÀJ�f��%��
����=��n�n�#Y���XK�K9��+��x�/��
�5�I@�mЋ��rDF�!�c�K�� :���ec�e1GO��:ڲz��Y9��+UkS��p����YU��"�UG��ҝ���::j�'��[M���4rs�%1����Ѹ��<_������3�$�zcn�����e�t�v�N�c�����}�u�M̹��g�Đ[���%lq�{�j�p\J3�h�ǰl���!3�c?������q@����m���Iҍ�!��L���U�,��m��D�������e2=�9�X�h� ���A���F�7���ݤW���:����@��y� h!�;��Z�F�u�dL�,�x���wm<�ɖ_��+�t��*�/�1ƔKy�X����}�w�M����O���۸�{�ܓ4��+�!U��zA�nu5����+�fl1b�Ô>}�ϡW�`k�@.��	��"qq?�-�������?���I�����=���ś<��#�H�lE7О`�h<}�~��46����zا�4
3��0I���7o���}������xhK�Ԏsǁ�����a|���F����������e��::W���B��K�Q�]�y���x�b��uj�6�n���u�ڂgN�D}໊Xq���=+������+m��,~�hP\��p�y��
�sl�EeQ�e½�;#��s	ӝHz�;G�n�Ve�W�J� f�fD�y�W�ȉ�d�z�J����[�|X������m}�o
p�)J��a�0)��9{/������m��n�]|�g�0��'�jҕ��V��ZR}�8�9��4��&��dVWO$������{�����;,��͊���c��h�a������&�k�L��vd"M�2�!ii4�(" ft�����;�L��k�h	!�
�Yh}f�,Y;c��
��3o���6�Qw��y��MX�Ȩ#�D:σ�t�E�^�x
�������9��O˩)�����Bgv�2�,����znsd)|���!+�K0f1>���!��ǟ�O��-���i�s����ç�p<-��,�ܔv�l�6��|��m����Ć��z�����o��r�S԰ҊpEd�œE<%�%�߿��OB`4�T::��z�VT�����K	p�� :T
̐D���I��t<��v�s�T\E�s��"�8V�I;�1i�>J�G:�=H�_�C)�&W�1a�P:8ݝ�/���E��7�0��\���S����]8���l9�E6�஻���q��Y?�kW�Y><L?EWhgeI]80^i�P8�-���)X �#ue����G:��u��u�L$Q�4��g�"הJ�8\�}�oA���9bR�B�*�T����}����v(&ҧ�md�&e�������<��wT�?g�-���i,����~ym�s��u��D��=����j�/����bDOT臤�n1�/_�`����B�?��K-��H��mt���ky	Lh�VzJ�
^���O�u�C���%d=�I"̫U�(��T� u'=�a�+��ό ^����+&A�m�X.�&y�����%�~w/�J�|nX��͔���l,�N�<\���}����2�(���u���P�m�J��p��(�Uŏ�~Z6�?ӧ������x!	�~>�I��C�0�0�^�y�~���?���`����������/���+F��w�|�FБ�&�	|��o�r�)?3鈱��G
���	M�9����	�w�r�j܏�Ζ9���~0��A�h,�f0��{%l�k�ޤ�v͹��i�"�9-�U:�Q��TրP⩋�Et>P[�
�{��Ex��i�ᢡ����\�l�Io�o��@ö�ŋX*L���336[��"��*�Ԩ�0QA��$�S^���$��.k��XX&�~A����k��~�;��o>��X�,��ɕm?���~E��ؓB9�e�<@X�x�ъC8�6cdH������V�Cb��g�ڹ�|2QFMё�	O�G�[���=�6����D��~ܬp��@|��Q���|�	ju����냐�LJ���K7�;�����f;y��g�q���0[8G�\Q�V�޾���U�7RJu�@�X�?+05����g�c83tSc�đ ��ɠ)�#���7�1CV���XN1����WA�W�!�r�"��	���7��X��	����Z��_����_����Y�.��6�1f˛����%0L/pm*�6^5����.F��׸`�Y#������74h�3G.�z��Ⰶ�+���P%�po(2-ĵ	�#��݄�ng�:(���ؚ�B�t���pQ��{�� ���I���o�NT�#n6��e.����3Mp����IT�I�a�s^+9ǒ܏J�����t��F4��Pj?{�%2�}��k��=
��Ե��V[y���hq6P�,���*5��y��1@$FT�'�[��jڐ��fK��^^�ƀ9�J�hC����\�<�a��}�����r�G�g�>D���g��i���2�{������d�����|�(�ؕ�N�(X�R��ǳ{�br�0�O^�T�*:��R���7�z�ԕD�h8�R�K�jwV�U��Z.�:���A�P�[4h�y�]I�9JW��e� &�=Q��cU�H�i�b�/�X._���^�,�����o��.}��w4b�Nܫ����￥�������8f��fk���������՝t�2J�W���*�]E�w�;`Pً,�7�s�{�����׋ф�y"?:�:O1�$�2j�j�'*B׼m�_s���qB5�ؤ�2+�9��6ox�7J:͜�Y��,��Ê�������Ms�(������in�ۼ�Ԙ/��/�|1��!�S��{S��`�h^.�|��[s�E�%��ls�^���=�P�����aH��u��4�~���!,��H��i/���M�+�ΉOy�~]������1��`���vhkB�1�#�i�1�	ə�)0��*W�ecó �/߁���k������)H1Р �A>P��z��XT�q�����d�Ɓ��\��-f]״[�ߴ%�Q��8���� ��7K��-ѓ�b��n���!x�nG�Rי�E��p*���x�G���w` ��ɤnJ0.��Kg��Hs��l��jX���au9�o��7G� �X-F��6(D	�?��<�g���_	�������^�����O	���[15L��:�31fC��jh'�d�)T�@�#�̞ߨ�c�j �6�D�_����s	����@��M�{+�{�#�d���+�fe��]���˜���]��Zs}���<�9��������n��=+!:DiÍ~�2Ow�d^c�g����y��HM��X8p���}�^�i��0�)��.'p�y�G�ϳ~�ިy'�/��־�H�U�)��N�Ōa����
Ƭr�c�ջ�PF��-��V�C�`C!t�6w�Ӡ$E�c�l2N��Jd�=�8�n{���&��D�m�i"�ާ��^;�%$[Srm��C�:�<��?�w��C*dE���h<Wa����n/V���G�o0�K�Z�ω�ϡ���Q�)1�<5�,��s�H�.���j;�ˢG8E���ZQ ;��@B<I�j50Y�ٔ���QPTc��ǜ�x?��4���ᔩtSH2�4y��!æ�ӏ?��o���8o@X�����@O�UA�h�E�c5�����-���jEDG��D��q��[<�r#bBF��(1�x���_hȥ�����9��b]E;�L��f�LC�j���?�9���ܯe��q�����A{E��"��W�ywںUۿ��m������=�Й���%��Ys��a��:ڑ�h�3��A1���ʓ4�2��/�����L	}Ơ�cP~N�nU���A���ĩz�x�]��J�ꎜ>��&�S��2�0{��C�H|t���� >c<EU6MrC0�ש�p5/�~o��؊��^D���w�ty 2w��ar>�i�,*�Zww|l(�L�s��a1�x��t�B&��I���d�>5e���;���l'��D�����e��MT�zEX7<g,Vp���Ar��V#�hEb5�6�0l*�4Q�|X��6l<��rb�C3�>,Mxw�=h'��~5rj�4=�(��#�2]Ox�?��st�L�F���Q���>���kF
������M������e<1_F�U��h]�1hEl���镼Ub:v��w�r������x̠�=U�Z�$�Tb���+�������NZ�AA�w�1ccAD"1Ϊ����0��_Rƞ!�)���|F�����{�'���D�Z��$��	K�'Ut�OWx��H`_��T�х�<�bD��m*R�*��q����)�o|�&���|��>����hyvaH]Q!���!Mj߻5|[�9n�T��  �v�]h�Ӝ��"4ڸ�{�	�{8 ߐ�ƚ^{s�-I�������0��k!��E{�d�G	�T�=�|��ux�=��x�B$z9����/���\�&w�?O��>����!�Cq�U@�V0eO����\�<�.g7��U!ԘG��
�`:DM8&�&o�wR�xY�jHW���K]�\�q�5��7�]�܆"3(X6�%��8�i c�l��v��׺׸V<r"2��8d��g�}�2�y�6}����}g��0L�_d����{�ws�������y�d�}��)�����Qe7D�K�V-Ԁ��DT&F#���o�����G�޽��>%ť���Ue߫Wo��m⸂�J��1�Y���æa�
y��@�*�C��nal���u`�q�9�L�N�*��O���&�
L��H��
�:����$�Wc�.P��7_x�^+�1,�)1�⸺i.t6:)YP|L�Y,-�k�(/g����v�7!�ڀe�6���R�����-B]��<K�g:gж�@��3i��N���6↍<R-��H'y��)��q�D��a�&(�kVBϳUh�rN{'}XL\5��ۧ}��1�v��=!D�
���?|\<�O�V�`(|�Lh�}x`7NH�a3px��pߝ)g�ex�:ҡ���9���Iʤ8.��H'4*d�.^S��������X���O�,��"%8nr^���0gN���U���S9.h-�ˈq�kK{%ЦHxΐJR��G�뒾����J!
�kÆ���q:[U��3�ىs������sot�ϟ�`��J��e�6o�8��U_{z���s����I��p$v�����ת���H ^hϬ�(K�7�4��+p���cF��M�Q��F��@�[޽^�9�*!��r��j����_獎%���i��a!�GCW5�I��y"��UC�*W��T��M9R!{`񜛱4 ��Yzh�����9U3Xd�
L���HSع�wϟ)º��c�u����R����Ӌ��R����X�m��\r&�]$�����h�4��U
ÊQ�*à���}N
�抩��-=�M�W�QGޯ�
+\q��ߗ���Ű������V��S��٪_g>���x<e>��J]�e��)q�Pk�����ד	!y�
��Á�		���;��� �#<h^Έ+thtp��ܣɚ�� �Km����~�*	�a�~�fy��,��RʃJF�,�՘��^+����p� ϡu���	��D�����ԃ��|����n��5�{ 0�*E�d�T�-��+V.�����t�/��̐~���<�:T���0���LnaX<\�\��D"���=�3x��k��H�k-$*��14q�3�s����͡�:��X���ղQmyk�j���p� 6�M��4���{��HD�ϔ$j�,k!dv��~�1ob��9c�8wќ��?e�Z#5;>��R�W�+�!a�d#��(�cR��vJ��kH�p���$�ֶ��7hO�L�YS.r,C�^@=냃{�{��gā\���Y���\�R䀹�md��zC�*Φw�3�R��p�$�a����r��T[��#����P���}�Zv�4�U�}�}�ʐ�x��"�F�E5C�D�w�MMk�������|�>Y�<�.!_hal���QыtZ��� `����C�h�h-N} e�����Ta�k0ygO��?/c�*��/"4��Q�"�c�)ƃ����^=zRr��^sI��f�1�!�r��s��T�P�e�C�%�Mt�-e�H�`LXu�d�}�~Hj�	�Q�f@A�r���4�#BoF$��� �똏�By,s�&6{lr���?}�!}|���ɱ�mw] �x���V�/��hvK�&s>�X�$`䍧��R�L9�Q"G9H�/ב�d�<燊��t��[�Ug
X���׻*@{��T�h<�q����X��B�չ�*�d���'GƵ!��Sd,����\g��3٘6
)Mՙ��h�dI��}���$���Y55᧔����r%�$�$�N��$,�H�X�͜�}�6)�[¢�/�M�v
!;�=ڻ�F����lı����D(#HC:�#qq�'JoT��F4�YLSeH�\Dzn�x��@o��v�2��٨�$%%k`̇h�P�3���;��O�5��F�ڧ?P��tgZ����L.��Q�=T��n'�Mn^.�EY΁qN�W��?0��&	pjQ��Ǖ�]L
�l��cx_$��9��5�����͹	�=Rx��,��T� _��c�ґ~�1g�?}��͎b�Q�&d���3�8.�����R�o�~C�:0B#5i�u<-ǖG�t���%.h��F�$lfxR�g^�M5��6���n]^�:��lE`�xЈ�8����e�=ۮ�����l$OM�������	hm�q]���)����>�?F0P�
-j/O{�ִ��4=TQ�;)sqL���S�m_پ��h�ƪIW;�W����w¼&�_ь�9�p殄5���B�R�a޵���2�Xp��|c�Τ��Т����hʓ�������v�����@X�(��g�v/u�u��n�';�dd�Q�V��h�"��c�F���*�qTP��m�"E
|�Z��g���'��mt>�՜ͯ���)ZN����t��8&�]"�p,L�t��;BR�����}�޲jG�4�V��iʊ,ƠD^����Us�PN^Pm!{�Ә��%5.ᥱ\���3u5;�J�O��B����	Z��q<ED#e�5�2B���u�#7l��D��l��������2�q�ߜ"Id��ןKu)s7E��e�織x���+p��]]!���Ű����'}�h���a�M%�=��S�/�Y��Ҕ���M&W3V҉�3{�M)jP��AFxtr�>�au�@�f`��K�Ũ�_�7_��&�\�����dIm�+u����Y�_�������x�o�ض9A2��%)�&u <CG4��nEޗ���P���3S6��E�z��`,�������EB���ˇz,���t7[a����9 �dq�ݻ?*���� �,}E݁]rU�b�p_@O��MD=���ˤ���l񻻹ͤ{֛cG�B�96�c4�c��[*�x"�ӂzfQ�)��%�I�����K���V���4��wO2`�qbROك�!Z�J�:ȺCl�Ǝ����R�tΟoA�j��S6kCT;b�(tn������Im�72���[Sr�R�M���bq��v�GJЍ�C��3�4�I7A@?e);��VK�X�8^�!�qkW٘�>E�!�Oz: }�O�(qNY��h��n����a
(`H�=OQ����
����J����"<�ip�����RT�5$��"����el xnO�h�UaiS^<���D�%�m�f��܍�i��$�X��b�����y!�dJ��uŒ4��ޕ��˧�i�̘r~�z��h��4�2a��i=�bb���%vqV��0�O�!A�;��?/5y""��E�rQ�SV��y��(�iG��X�d�������\�rmOO��}�A��J��F����=�-�ت^(�q	C�9}:]h����Z���b��Z\Ӭ�ވ�K��u�Y�]���SS�(�[�?{}6�
�ֹ=2��1<3d��:c����Ĭ�J�����U߿�ԭ��=!'u!P햛�SH�ɻR?��X۫��.͙�P��!]�Zg�3�I�;���aՓo�:x���TȞ(������Y߻�B�i�"C�ce�4�4�c`�dy,� �p�$�`Y��>xYC��b⓰�%W��[����c�춱R���^�q�Ȝ%B#U�UD�����5���#,������ �?���9���r�-�QѨ�n�vyn�*���<�s�����^�:��ht�I�3�ڔ%�q�u�L�͍Z�Q����5@����<���fj�0��b�w}eC����X�Da�<�ݪ���-$D�9��5�z��lmC�JU:��&o���3MA��8S'"Q�w�t�`���a���ĉ~�E;zz�G�󪖖��&x'X��ʹܵ�l�֑pi#��%�`X�7�w�{Qկ7�z�=�"�#x�kqt	���<.A7��ا�k�A�Q��m��:%���7?�qs�1�T����<M`��d$��,3�c&%n���0oTQY}K�c��ğdHy��/��ʨ}uT���<Nt/}���!��K(�b9P��U���C�Z���AlH|b񁆆369�s��o޾Y����#�-<I��eLnwڠ]Y'q��3�PfIY�p�P����Hś��Rجq��c��� �#�6hv�1��U�m\I���Κ^�pu�Ӝ�>,����X�3�{�!�/TΆC��zf�M4E4<DGi��@&���W)_��3e��<�>I;��u��T�l�Ӟ�7D|'�uL��[�QK`喛�|\��钡&z�mg����*su�������C}󟔈�p�J��{k�D�Z�up�t2x�R�ìE�$�K2W�]BJxiY85�C�n'��Oו72�4�:�BY�^��i�-�5�� ?^�?��?s�#Y��S��9���ܭT4����]O��d��ޓeOjL��Л�(���ٛvG�$Ib�G 򨫻w摻��������73�]]����pw�\f����Yb6�	 w35UQQ�b��F� JVȔ�j[��*�Rj7v��[<��=��x;s��'~9YP������f�Bֆ��B�8Nfq�ee-\ے-���BkiE:�JD4�p��P
��̵m�%'�tД<��ZZu]JM�!� ��X>W��U��ͫ�*w���*�#+_|�܃V1]��\$�#ۗR�)t5D��le�,�=a���l=z �T��|�p_���F�Cm����]��$%�T;i2ֆ7fZm�}IVB5Xo�rl�ڔG�N�l��!���~���ӣ`=����g�p�p������s`ct�O՜r��2�u��η��c���se�����*���k�)��GBײO�jg��a�.w�v��s�-�Yꆦ�ͱ-�4<��lޜL.᯶2` �`�;�����cv�N�W%$+�Wl��Ģ��kB���ܪ}��T��AEguSI�$
*��ԩڻ$g�ͩ�T3����ИHXf9��!q�+�M0r�^^*�<^I�R�(�Pn2ۍ#|o���$	�	^�!e��0�P��f�; ��b�� N�x�w�q�U�Jj?S�/o�'�*8�Pw��m�Xa����$����$����i�M-"��pM^_�\����gW��|��8�.kÄ�!�}n�����T��^ȭv)]�g�acj�:WCa��:s��C8�!^��?~���}zW��L�T9J� ���y�6�Mn�b�]�ԖvZ�]/	
�<a�//��f�2�3��x0��a�@KNj����x���R�ʠ���7ۖ@IL�� ���߮y�q5���}�(;� _��dZ��.�֤p���_V���k��a����4���R-���e�����`�B�P�9%h5/R������t'`�()�u�ϕD��b�z͂*; ����
��أ���*�w�C�$���"Bt���gss�I�����>7%�A�F׿�Hqf�]���կVw��Q�L]�$+�63�[ن�hTu]���C� t�F� r/��z�y/��:2Ql�w^�g7���.�7HF�*���f�6���Bޘ5��Ha���kWtM���J�
N9Z�J���C�h�Z���K\-�Ji� �2�~�L&Ͱ�f����m���a5#�ԬF]�c՝=O��zY#�'O�2#�k�R�VA4���*�lq ��5;	��X�{�bU�o}������q<�� |����ӱ��R�h�R(x�������"�˻�qO?|��ғ�ܿs�� *3,&c��osBc�L�iC��)��Wր�3����A�aZ(R��E��u��j��9�tew�c}=<�<�t?����]
�.�7V@�H��˄e��v�=�n��Q�	��Rs����_C}���䲰W,��ڼq6g}��\&� e�Ud3�����jF/̀H��l�٩�k8&��J���s�]P����d �2>
F���ke���-�$68�U�ЦؤZ9��������9��,k���.*�����kp��<q(�l"�dTqmSb���Y�\��AY���̓`�����&�{.���-�ͪg�|����ԎF��\A/A4�^>'U�X�f���-�]�י}�����x�FZv���մ�(�5�{��+Gi�R51�qʹ9��9���� �
�����P����yM �]�c�������o�e���5ʲ�&W-�����$cػ��JL��Z�j�6��>�QT�)U�M!,\��p�2����_�ıyD���϶�#���	ߊ/ueO�W ]��Tȥo�誠GA \��7����vo�5�����Um	\�NemJ� ���_�=���|��-k	�b�����]�<W���&誹��?3s9����H�N9�mW���.c�C�楖�����F(����'ˌs�jQ�RD�r����C�k��Vg>��+�/�+��*>�uo�oiC?�϶�+�v��R)TyT������A��@�\���.��YVO�(3�N(��T�����J�=��@T�+���dY͈R��Vz��1t�1[���F����KyM��q=��V��W�T��v�Q5�K;�]%d��P����a�Mf�W� �<$�rYls�;�2���p�^G�>�N��o�fk���<]*EI��R'�8����E��P1Y�(ax�(�xY�ocC��#�wU�svCs���j���T]1�F��eׇ��;tt����(Mu�rn���s�'؉��*�&�������I�`�L?�3�
��1+M����w*��E���$D�Q��lú�4�K� �H�Qq�^�.~��2/�ґ#���ə�����X�[M�:7��n� Y6i�vn�	�efr�윳�Y�x&a�K��t���8$��PZ"C{�6>���}��]��D�yb�z#�	#Nnh_���������q*�ɲ �B�7z�	E����K���2�*��F3�
#AL_� 81k9�K�v[+���?7�N&�����a����Lt{���F�yWޫ��# FK@^�\���@:֡�L��N9$L��A�M�@��?e��`���ؑ<앵�����6\U��b�=lK��>\(i��n��)GF�'�OQ�R�Ҫk��Zs�_^5�|y�Ը�a0e�\�}.�w���A����/�#��ݽ����u�M8&��=�@j:��XY8��/�.��컈�OT��Ņ��W�����g+:����P���š��̓�V4P�Ĵ��:5���o'����U�;X�H��ݻn�O��5��| X�4M�`6�G��
`h���¢V�:m�L͞`u� !=
J�����e��N�m��=�7���eM�\*l��d2V�v������b��f&����q�jfL�<�Y%�����֧� Wfj����|;�õ���J�����?���j�{Rr�Y>��ù�0F ڊ^�,e�wQn�W8D�;75<>��_�x��vM)%$`e����Lg���|��#�k�=(�\�B�l\M��q�	W����ў��K�y�u�o��v�VX!YQ���:��ܦZ�����d��D��#�����iZ�}�Ɵ�ftv���-q��ȡ���o�[�c�YU��g�u��3~:I�>f�i��������$x�Y+�]�kD���_K��뮊J6_ת�a�K��2�J������+^�JN��xjKPJ5����oƃ)�q�)f�}���V�����?f�-��+C�@+��!�e3p�7�M{3��R*��њ�^�i��*�^1�t�͒yk��<1AOB7�)3wT�Ѱ�N]P�{�mr�e�Hq�^R�������O���X�ݓ4��l�4ͳʙ���`>�Ue6KE-X�"k{��H��W
�h�f2k`�AY2�C�����׻�ֻ+�:�T�D��z907���V��~o�~~wh#v\Ȫ�'7c�:�H,���ȱ]��TBm��@}:ߠH�x�un��Ɋ��6YSi荄�$��xr����܍�X��\"����3�G�ܥ�|7>gLUi��x�v�Б����ŪW������p~?o3,%0Ԛ,��gM�<ص@6�[ �C� �7��1`~�~G�Jg�	X�\��N���Vԙ�Ǒ�Zګ
��"�:�!�62��6�����T �����YdQr!W�s�	����E�S���;������z-���+����{��J��w�S��ѕݪ���[%JJ�5�n-����g���k��]J�)����ͬosm�EzHM7����$VGm_�-�$�T��n/<P�\��XXE(��������/n�C�c{�w]�B��HU�o/f���ظ�q�cF*��h�*lyl8�%��lN"�����D�����Pr�sY�/����%��󽙋��v��R���9�tU�`r�i�ќ�<! K}xp��o�^:��������S���0`L̼R�3��,�Y���L06�d[MԱQ�f[�s��c5|����g�l�o&�
s���a1gWΚ{��	�i���hK���_ه~�JJ��L���R�����L�ԭ�To�9\�R�(��c�����8̳:������S+��Zt�0�H�!���� k���u��=��֨k�N��L30�`$'?����2�� ������d�-[�~	�ے���)�?&��Z���+1q��haݯ叁4L�}7����$����\C�r��ΐ���ܵ�3R�ͺ�O?��&���g�E����ހt�[��V��m����i���_�k�������s 똡6��a|�SMĿ��^|RNv�81V�����QF�G�z̾�Vݩg�l�73�K�W���X�X3,���TO��ṫ;���Ӵ0���V@v��6�p��59����)��0�q�QB5j��zeԢ`u%)�y��:��k� NKd��3�t+�/|wN��=j�����$w�'� z X��7zr�<x��l����bLB ����8?h1A6�����٢�S����r����lH&�g���|h�0�v��w�4?���wC�K//Y�F+&X�փw�����kz��hG��

���Xu���{g�ſ��/u�L���&AY�0���Ǌwʉv@_W��ACu_��I�O���Ҳ�L�-p�����>3}D[v�9n�Gj<'�p\���(C}1�d�]۹0����+��TD��������e�Pl���fJ"bL���r�h��0;���;a��IfcO�Ƣ�xz؞����:���.�Ɏ��������l�g�c_��x�?�]�|�Wc���I��ga\)';7�NG���y�PuEx [���yq�{��gk�t��F���ݼ��I�:��I�k�����#�_d���qJ2,:ȿ}��~f�:�I����Ar7gq1{F���|4��#�\�{��S���
����矊\p�3��.��*Y�<�Xg�7��v�#i��WY��<	�r�n,YC(�A4��\3�Ҳ�uP���Edh0	\׫���#�b���I9�]o��,��X3�Q�*p>]+_l�+��w�]ۃ�oa�'9Pt�x]��VoZj%��s>���d%��믲��DҏЎ2��s"6��I$�V|t5a�M�T�=�Qn�2�g�ð��R�}/ݽX��*V��P�y���蝶c�2 �޵nT��m�;���Q���f���&\1��K�"a2u�6��ѳT'Y��R��=��!G�����K|+?N�?;��<��z)����K�5�2d8�J�))H�9+c���E4}�����I ��S׫�x��=���)b���������|�O���Aԡ�_H�8U�l/�4��x���0�0�e���P�����1���ʵ��?���U�,�7�$��g��9�P6xwV�ɱ[fw�$ie��
s������+�-2��M��t��Ρ��]Wn�2냃e�=�-m�vXK#V��R��ɲp�o����*��uW�0����(��L�e��S��?�<����`�E��Q�K�D��^Nl�j�4��4ʰ����%�~k����m��e�oqS/L��������{��*zQ�7�6V��\���J��g�'<>D}�����MW��k���g�Zj�v|nj�FMj1�p5o{���g�Y?�}��fb���}�B�J`�N�X��f�����Ev��� 뉿֎��lIܬ���J^.�uss��*F���řc����减Xf {�9�ۍ�������Aj��Z��9����;��~�!^"��gbKT:�SwRp�a	���q
#{��_\dRx?�_���,3�NA����Dǆ5�/����u������H���|��Y0�,�O���&���<��F��))��9�!=�A�=���]����R0��� �u������\�A0�����v͓��î5ڢ7������Z�.�K������=�~Cx���t���J���F;ԃ~�8]׆󆸞\$��wX���x��d�� D1��`��XPM��3��Z��v8���#1��(.Su��iWG|�Q��ҩRC�h�I��-�IW��/�\��ޥL��XGG���
�?�W{v:�K��O��x-�G�V��o����^.�l�����u��\'&Z�[m�L6ܧ*��S�c��]�Jl�M�9�V�hwU���ٰ�i�������7t�4���lj��{���&CU�^dYuLKK�~w��_*Ƒ�����٥L�'��M�v6��D
k�"<y(�kq�t�����������D�;O}
+P)]����� t����ba�Bs��,����U`�0��3�/��s04���=�_7#�X�"��ڼ�-}��a��M�w`��L/�_~�I>�)<O�g~����!�}&�T2w��=�F!��f�X�
��?m��x';�x�Q�����"��(��8�4�|l	ޞ��R�K�1(���<��t��D\t��޵ݷB��k��Jq��\�����}��;�RQ��Ww��k�8�<�&����o�X/go�V�
�^7'�OG��3Cm
���_�p�Fu?�e�&�$$�D#�C�4���&8j��a?��[-�� �v�t�����'3��@���l6(+e96���I����x&��>,�XqX�+��VV���e����i�y']Zu!d���p��Z�S�>�Q
�"�<��X�g���3�:k���ɻ��.���b�g��6�3��Q�t��]0�]@hI �E�p-���r�����MiV�I�9i�U�h1�zD���"���GM.�&O�3�dw���b����ww4�� ܳ�����V�u"|�����I� �f5��2#=q��\��=�>5�\FƇ�p�� �37Ȳ]���M���������x�����v�#�e�ˤL�}y�20F8�	��u��^�bΠD�ٲ�&bA���%6^�e���\e�]�鯩������<��T�җ�_�
bFur�%�����~���"uU�#��X��Vĭ�ays�hVۂ��t�d�|0���_��.w����E�w��'% �N*�:q�_�AO-��T��F���;�	��A�uUsK�ߍ��/l���x�p�ӟ����_~����վV���]�3�k%��L�m{���H�{~B.6�ý@S���SN_��@q�Mq0UU�����T��ˤ�=tn�6u^�6�'ׄp�Em�w�wб�:j[j��-:ޗ��zmk\t��*���|E.��3�c��w�i���v@��x�gnV:��ӽbP�p/6@�B��R��X���<�]~��9�������ֹ��Uy��X(Ͽl����3�6e���*���SƄ�b��t�o���w�/�e)1�j��(�ДO�*FMe�9�с��Yc�(`�=
�6�-(R��F��;��"���|�A�@�,Rg�O�i�uz7UɿX���F_����w��3ʭ)�Cm�-������_^>WFƃ���6�tlX�u>i"8sC��:���8������ٛ-�4w��ݪY	�\�����|��L��ޙ�W��~�87��_-�+�#o���<�/yz!����i���[�)]8�� ���]�T|�W[����WHY�졁���
&:���X�0j��Py�Z {�(����:H6`u���c4:#��w�I$d�x_"x�����T�o��s%�DqZ8{�a}w�}�-LX��\i�f�z#�w��H_gus�b�j�A�Y�����O!Ϸ?1mmA�M0ݳvj�5���s2��a�HuM��W>�&��k�@zs �[�[�E�ND��>K�����e��`���q�y�\Ɲ\��{h�O��W���x��~f`̜-�#����e�{�,qv��ij.=3�Ʃ����������Z<X:z����`˲���y������L0Fu�ZH��52w����L��?Y�X�Ќ��1��l�������5�/�tI�M'����L�B��qo��l���VN8�x <h��� �u��w�-��������n���PB���JHp����x����T�8H�:�zr�=������
��34b�V�	j�3��Liny])-�,����^���] �}���c���p��z�~C�ה��[Q���ָ�n���5�����R��` ����o�<�~!�����pSn��:|4��H-�K�j��u�**pE?o�)�y��Z�O[M�{�����	��9\T���0�:C��>N%c�I�/}�����oƠ�7�/��kEa����ochp�?ӮQ�G���.������Ͷ�#���ke��E],��b��f�'���l�4�>q�ܧF���Ha-�Sr���X;�6�f�L�q�O�N�/����pN�s�q$��_=Ut:);�=���l$m�c-Ii�(���C���-�<�{=Uy��0���Miz2ܑ�Zf�9�I(-;>��Ł!^o��"n��oNR)?�/����4VjH�Պ"c�׫n���4�����8��6���ٱpclt��__� �~ ��AWQ�&36N/�*���t���i+�>y��8y�'L�ݕ�md1e�>�2�GZy�cP&w%��؄^�ρ�F
|�q0>�Ú�R�8����N���U��Ҩ���F G�������ߥ�o��K�u�k)�'3��c�9��* ֆ�Q	of�a�0�h����ꤘ�+�k��}(P��4ݍ�P_���5Ga����gW#�[6�;������|�nf�,x��\2��$����Di��#�v���l�m��zk��"n6@����\ꌬ������H�yW`��~})�W������7��H!����b��"�XS\u�W�ǥ�'��y=�cz2ٸ�k��c����S]e8�����<3�-+����r��mdc�������:x$5�1<|@�ꤘ�X�S�ĵ�?2�S�}s���s:K->8Ny�c�
糲����uց�Nx�pҜ�W:d~�@Chb�dUS|�n�չ�ar9��k��݄��n�ʯ���N�),Ȕ 6��?~-�x��՘*4�n�K���3����d���	19�6��ަ����.����J���u�1{�������A%|�?��2PT_�}fV&��VL���[8LSQ"�ܮ�to",+���#�;�Wa�i�������{��8��G�w��U����+���Ӥ
�	{��%�F��x������.��D�
�냃���?G2�*k�1�����-@�z�WJ��Jw?�#��{�4*�n�fQ}����`�&�V�s�ҵ2�%����Q3��S㦮X���ț��/w5�"���L�����e���1ݲ=FY=:����Q��A;���%��Z��͖���G��_�dͣT��T�c��� ��;��Kw��~-ͧ��x��4��XF]ѡ|�J0�������Bc���V;ͫ1�⒝��E_��oZ�|}�=�sIԜG�C��vB�¿�J#�}w���K;\�Ԉ�O��y�ZU|h�O]u����ܙ�����N��|��߷����ݫ�<�\o4>;HDd߈B���;z�_O�2^�7��d����Vc���^1�I,�{m0N�����(�˟�K�l�R�0�AFH�{W����YhAY����M�HO��p��Z,����:|���%���IR�^g��:`���`{d{��u(����o� '��"qe��KU��%��Kl�����|y5Q~�"C�A�P�,2��L��~f����!�E�XW
��E��=JIw���6L�����_��mSfށ��K=�Sv0��[٨o�X�����#�v�Ics���ˋ�1�U��uWG�h��9��/Δ�~�:��b��n�
�r�3,�3�ȏ�Z�c�q)b|�&�v8=����MC���@������r=��.l
�E@�BK#�'��`R;�I�(K�XX�m��)�4��ɨ4�H�^t���r���y,QM�(J	��
\���,�� �^����3�x_�__�o)��,��Q������z�	M
d���ū���N���]�!?��N��������Q�"���'��u��*AG��
��!fO�dn�'��	��*�n��&�C@ȔP*���扜��V��A��w!����$"A�(��  �N�6�]W�@ F�(�.R�l��:�;���^����D��U�4�W��'r���ך����8���\M������6�����t-�J���b���:���[O"���+���^�����A���Hk׾��oS�҉~0�Q���|:qZA���N&K^�Cx�%����'OiL$��F0��d�Bn�,���/�9m�)��e���)K�i��/n��<,���J���O�}s�>J�H�N�#p�}�d�&�GjBn�8��z�)K'�e�Ց�V������?_oM̫��ص=���`Q��O[&���r�{m��x�~֚NZq��ػ<�kT��%~zd�q�.��912��()������=�TO��K��a����x�QNϮ*������տ�q:2�����6[��V	��E�MR*`�l���M���b.�γ�F��u2m�0
���k��OKl�A�F�R�����������~%M68��
-<��C��ÊǬ�Ш]ڡ�ks�A��N^���q��Jە͠��-%���n���ވG�VI��D�Z�� %xO���T�$vȲ���믿�#�4��d	1�Ɂ��Ң����(����:��i;pN�:�]�7�1.o�B��B�׾v�}�݇�Q���_��i\��6 ����6��`����H,�M2Ǉ�g�����#�2��"�uo/� �}��4a�:�l�PԠ`!�*K�}�n��1Έ � 穉PZVs
���p�5���4�U�8�z��'@޸{A���s��f>\%p}����K^���0'}le�|�����(��G�>����+�1��u�|�)G���6�bU-�
�p��O|I��n��)�e =���yRQ�d۰�ZWY	����Hu����韬.?�R�5���Rim����N� S���D#�U��P�ƥ�e�8_~�u_\!����� �H�d�@���3q�����
�����u>���l;
V�e/�@�ʵC����S���@
~�G�����|WqteM�~7b)�q\�/��2����U�����K���P�8���������p�X�n��
1I��3�=�A+k='c!�����5b��̿�"�Tl~-�4���Q&�t;�[�,���{j��v���@���ߕ?�d!�v����}.�2�k��2�.5�q�J��]#[�� ��i>�A���i!�_a��)הJ�b��l�7Մ��o)���R�|n�Tb��,@��.j����3#]��'e���jZ��z���}��md��u�a�T�����J��b���lG-�BF6�,�c�]$E	��-E�����q���c�:*g�8�S"K:X��s�o1D�@���#2Rtg nTDw�Y���><�] �|r!~j��P������w�:���B��������A��i9����33=9��q6׬�SC����@z^�u�/���-P?�Cű��.�V}WF�Ȯ<�%��A����@�������r2�k��t�c��De%���y���X���x�
N�w`�}u�������o�Q����?����O8�̀�PC�F�>�uw��2������=j��G��w&�ͧ���x�N$Q�ik?L.籞��;�bڔ�ܖX�ⅰR:J��-�׹��x�7�j�59�M6�i�oDQ�&��d�yC{�v�s�#`�-S7�qe�:�p"�W��D���s%R��_�j��E���p�����e
g��x�-
�/a�~�;������`qE������Q0���̒
�����.R��K)��k@��,r���9L��~b�s��I����P�����R�����K��2ƶ�3�p�8�g���L;S:t��$ʿ���xq��V�|��3-�cvS �Q����"��������ȉ��Ã��ޱ�����Me������{^���h�b�}�x�o����!܌�_�9apj>0��B�j�oޤx�7W4�w���L�
w7%�(Ac�܋��*˹��m�QX���
:>�t�ޟ�Q�[q��P%��=��g��5P���%��V/�^ko�,_��v�.y��7VL���<���IMd�m���&�k�C!�we_��m1S�k�'���g�z��^i���OU�����i�QL��&���Z���pG���>z�R�� 1?O^��P~�
��gdU���X�|~e��p6�'bB�IP��2)�?��h"��8%�k	i�(����<Iu�]��DAɉ��V{B�}f�S&���S�
�,z4�r �2�d��r��|׆�ٴ�r��_����BJ̕핛�ݳ������ ��A80����X"ne���^�޲�=��dD�~�ޔ:�Ƙ&��_ܡŃ��4RӤ����7b��Ͽ�S����ؒHɩAH�jy�)[މ�/x}|����ߘ�r��_������sB��y�N��M(6��D��ɴ��ަm�"�3����`��3���kq���}�=#@��δP�͖�����ֱd鮄o��� ޛF��>����r5�q�_P	�wMR�K���`~��'s�����1R~�A8d)�k���ؠ��u7��Y��t�	��66�'�
��ʰ�o��r�`K�h���v������y�����Qal��^*�jZV4$��S�լ����nݗ�|����]�P���~��{u�+\�u�-��3�t�	r�D6�����nv2^��_��P��`ꁛ�x�M�I��R�T�Jp�vS�6��!#��^0s_.hi�!���D��M+[@�G� �|��cU��U
6N:�̎M�_��(�CS�8���b�̏[`}��7P��,z}}��ݗ/�L/�T
��zy�a�,��R�	Jb��-(;-�QlZ(#Ǯ/7�s9���5�g�};L҅����?�@�L��`@$.V*��H���=�T����ȿ���/��_8�y:K�`5W�����:̈́��h�\��b��ץ�+-<N��zJ����9|PpvY��rsE��;�gB'�����'pY�u1�:C�-�ܾH_�`x�sr����@%1W��Ls�\�3�A����յ��\jU�@�C�9M( ]^��~�$�u�vW�������c���Z�����uTyL��Ca��ą8qh�{�����N�鋟]�B�8z��9'9g�K�͵/+�η�e�6bv���	��ث�Q�M�Q���,�ר{�q�6��z1�����'=2'N_u�Q�gw���C:{�] 7��2�[}��=���%ݩ��w'����@#A
J�������eL ��m�OO� =���Y�T�z/���[��e��i"wm�ApUiL�>��R<��q�l�a�<��M��n8em���;����q�����#�-E�R��~�r|�|��������3t��G�+�o_�0�'v�E��@3چH�Ye篼�T�v٧Z#x"�g�������Ϭ�d7����+�~v���8<�9��
5���8j���N���J�pf��i��?�	��\[/�t�')Y��M\�O�a3w�eأm�T��&��n�@C��yTwL.F� �V���j����k��T�ȫڶp���͇���$���=+�.t5B0۵��w~Q�΀K\F#�)��!䫛U��?�U�sk$��P���Ĳ�A�lo}�Ӯf�����7���;��v��R)%L}�E\�œ7���2��@U���NX��(*��PkuUL	��m� 8�h�La߱&��qZ�z��^��n�!��N��C����n�Zn���=�����U#����Lժ��U��4\��v�t��ה��q� ��2�
xVp����Fc�=f��P�zS�.�l��g��e�қM:��"���R�l4>kD&R�����C��2l�S���5��GvWTb�w:�^��]�7
����nK�˳����e�:I)>!k�2uЈ�>���`a�����M��0�P��6-ٵAz����_�cv��mt:v�M�Z<}���65�46��,���F67���_ .|kSX�_%��nx����,���dū�B��	\i�;n
QϤ~وK�)4'40�R�K)	���_�M�𑯅��Dq�j��R����tʚIG;�y0�}�u�O�+�@3�}w��~e���)ֽ���~�����w����Z��\�y�0�����N��9l��%�
(��Փ%X
)Ur��g�޼�uN㙔!N�� �hv�$���8�b"�������*�s��`lm��b��`���q�l�pT�A0~���ȆR�}^~⟾\�T�Q���4�@��&e�������D��Y���\7�u^�͗�A����+�HP��EY�n7<����En;K��efh�eQ�nf��l?3�xsH���K�*�3��+�6Ov����]Y�,�ss�~{/h�����l����d���s��<���-P v@Ɯ������ �kf&n ͞]D�/�a������'X!9�Ek��-^K(gG�Ƌy1�ܽ� �@6�)�z!.\��6�c]k�t���*�H�u��R��,�V���`���G�t��c��-Y��撁��+#&{.�x���d��\�Xv/Ǘ�w�2:��|:�+���Zi:�#[��(��[��k0c���v}6�([I_�s��i}��/&�"�=�|��dl��yї�-,�&S��e�T���Ԥ1���m U�X�B+�F�����x�����Y���"��a$f�N7��J��E�)�e�I���H�I������4Ը:oA0Z�P���3/]��K���~'���@�LP ���
�	��H�m�NlW<[?W�P���m�����,-#�٨��`b�{e"{�M��=��)�˫4���!*�B�}��2�q�nvrӽv���*�CT̏��)#e�	��C6m�,a��&�L��u��(lr�ؐp�3�"���f<�x�ceW71�|�{�b��?�t*�k�X(n�:�"�?8 R�u�����<�����/�Zۍ@��^���y���ێ�!�xTAk���µ�����MwN��sH�iPV}�=�a���ܰہU��*`�J�F�}Wa����M�rF�ᓢDJ�SL��N��o�x��p�e9� `���c�1�l�������R�7��@���w���{�\^b�������F%1�:؍�y�I!�ry���N&�&��1rP-��fX�@����@d��tR��3��p?0kC<�f�&3J�D��X�}�]�-덇�x8q�b�"�I
HT"_��C� ?��z�<�_��Y���q�#�}^��	�}}7�6�՛����昺�ť���@��3���Y�����zD\��m�H;������5��<
��z��>֬c��&Sp��B�ƙ�����ͫ�нR:���ᰄY��5�m��0���ck3T8�n~�����{R�ah�AM��-���C!}x��
�(K���{�RjC���X�!����^���zt���GCU<���A�@��X�Gi7sV+I\%౽� �5��kyD2my���G��Wke�,9��Z������vϣ��|�˰[��f�
Gޯ�7ӓn��b����}�H��]��� ��I�H������܀���_�|�aA�p�D�q�Mz���&\n̓��B���eX|S���V�z�t7�f�I�5Màϧ�t�b��M���C��/��CU!�wȒ֚����vR������W/�����@��-��H���:ƫ&r2_o�7�q>�R���b³T�|�#��֎di�����R�{��U�R�p����d��tb�����y}\M���c�&��󼡰Q}jU�k���xr��l����3����^�D�8�S�0/�Ц�`��e�n�b��~��rQa�����P!�o� ���bX�0����!FnG�>�D��z��ǒ�0Qfy�ŷ�������O.WS�p0�ƚ��6B�%}�g�a����t�PTOH�[�ڸI�ƥFq�����̓!f��`���񺧳�2�*�>���j��|�t��ܬ}������e�u���3��SK�#Ҩk̥���E�7ͦl��+�Ԕ�� �͕�8�}��:mq��#�����⩳�F�y������SE�=��[�̦�����@ ��1�/��D�����Ӷ��9�S�u�Au�|2��i�X���$�1�M����&�K�~�woN��c�������o�/u��(<M�K��q<Y+���r	.~vz�*d\ۮ.g:�#D`�@s�4S	*���T^K�]+��%
����V���/�ŝ�⍮�Z�8v����C��s�I""a�K^�>X���_������\�T&��I��V>��Xz� Yq�Sޥ�,�S68�>&X���N�#'w�ϕ2U��3���� s1G�f�u����j�p�հ�����}�&u`/�^�_NVC�P:�Bx�����h��1L ��]C�e�oゖH� �x�3� l��V�I||�>�z�[*��nh�A�AVN���ҴhT6��8��*x���+��a�r6�vL���h�i���7��n�#1�>}�?F������T;W�3����O��KM����Aʕ�)\g6:q�C�^�B^k�d���lj�'Ns��E��AJ�d��9v6[,;�$>�R""�;M�Lu��dů�<O\K�zAc!�DF�E�M>�Ub�����I���WMA���LgX�o
��LG7qn�C��e6d�e/��W�N.����U������
�g�߳�:x�N+M�|�k_9�����5�l>�|���[���SS/�2a�g]�X����ϞL<t��f��?�1�C��C�"�Q[jCZ�<"4k�W�[5|��Q!�~�T���*��4�����p:���:�">�w�޶m�
����U^0��u���z%������̭F��g�㞢TD�t��H�7�FP��hhTά��`V�����$>5Ϧ�I�ppj��4��z�Ϧ\�!��͕G��hyOk�;����0s�>���X��Mi�cD}�#l�_y�lj�sx���j+'o���D�(h�m��k�<&������p뢶��2��~V�y��F��9ܖ�?|t��f�*���bA"������[M��)�:9�,���;X=`v�n�˥��a$, <������⫛)�7��ȃi�ś{���*��Sv�XiS"߯U�*���]�q��Iq���r�s��J&�_��Va�A}�olNN�s�������;1_���L̙�>��_�����~E��x����9�C��o���%�Wg~b��MƱ���)#�iv�����첓(��K�bVs47V��^�q	���.Kq��>|���[�X�4Q`F��M��tXw����q���jE��2�s�p�J)Q�=���%6��-+��������'��]���?����%� ����y0�������o�+�G�2q��?X�4:	3�+�Gуo��KZ!�^���Y4�:L{&6k�cխv�I)��>n�oBg�Vw��m ��+ѹ��ͬ������FE�A�o2���Cqd/Q�>��H��*P%~�����O_�m	3�� n�>UA���� Xvvr�?�F?Y�Iֱ"ccS��t2ɷi�1�"FD�8�l�v)˩QfX�Zo�J����ѯ�����vs�H�����&��|��5l�?wIPO��8ؠO��x~d8_=�q��#��F���B���x���\���]�w�쀠�b�qf��O+�<!3����8
)Lt�7�0ZXe�<Hj�ԷH�3�����6���L�c�>d�y�>��I�r��\���AM��`��j)�c��0��bq���Im&�h��~������#����}���{LVlSsb�� ��\�m���5����<��R��`�- "�'q�U�K���$:D�c���p\��J�K'��_��_�P�ۿ�+?�vx�6SS�B�I�+���ĺ���~�u���d�2>��;�-NL��1/�_�?��:wc9�&������7wy���_�e�� "b�T�hn�l�q8b1>Äu(��2���}�?0�b�����d�asKmG|���T�� Y�tg~��ؗ��4Â��!
;ڱ�t.w�kc,��F	�$��Ju��uI�Z�,5�j�t� �F����W׻*U�k�;_�S��tu�5xD~N���L�`ۇoŋ���]*��RT��I�f�Y:�P��/[ �Z<��8�:k~ܘ2F�]��u���ɫ�v_�;P����R��ܽ��'s�_�἖p>{�KӇ|�>����'�׋�6��]}������7�"�F�5�22�qG`ӓ����.�4\u=�A��ڎ���@$e���++�4X�bSÆ�˟�ˠr}fy��uR�"?�􋼙�p�͖�3lCh�J�/�ٚ�f2�+��OR��_h�n� �oO߫����hG�'���fó�q�c��Ï?2���˿����X���ȥ%1����owilA=�G���/���֪k?Ն����I�Ib�h��O��߼��v�����H]���yc�n�Ӎ[ �->�.|��^�z��=�Z{:��3)��(+�����D|�(��+D����'�c��_-t2�j�� ~R�y+Ǯۆ ߭�@s���~	�mB`�){�xc
�ݜ�GԺg�$E�fJ*�\�$�E�D�(=�<�\�W
�`���9u�w[�����x/�W\"��Û\�*X]�.U����PR�hf�0(m�w�i��ͫ�X�����m����������J�NO!t�,|+[��)��9�����=����^�u�kt�NƱ���>Y\�	��&EUO*�P��S��l��
�A�C>�5�L��� ���\͓T�ū�j8�w�1��n8`A۟#Ix��o��2SBsi�T���>C/d��Ǟ��p�H[���Spq�}�]�>Ø��7[f� B���{���*\!c�]�Pf����5E�e��׻&�"L�)�+5	�j?�� ��O<Jbڸ����3b�:��U�`��ާ]�V��)Ş�W��j��=�KR7[Ì���%K���5�?u])m��}�޴�ޘ�0`�bܩ�'�v��"<K��RJ��Sj��^f��àE��)?��;	7�n�We'wz�?9k�ƣ��Ǒڥl�1���E�F�&:Y�2.�Ƞ<�;���3tw)n�����9�_�1k�/+G��|��;���:	LO���#�[�O����J�I��ڶ�m��8F��Z��YpUl�N2^�M����c�M�y�wlNj��F�y�-���d��13,��O��	GdBPw?nY%2�m3�c�`�ejU_�����~|B%���<�~bP����`���9�j�ƹvg����Ayג�a�[uv�ԥ��Y��3\5cN��`�o��]�!r�v��)_1�;M�]5�ò_���l��b����8�z3����b���&�M4�Dy+���-����Llbw^{�x����S���v�!������\�-Pa/�w`�H����\zޱ�/`t������t��ζ��${���n=<=�_��33n�@��~�~w���!�ö7�z�l���,η4�Xt�OAU3�c���D��O|�W�����P��d�]Wꁮq�H�BUV<v�4���Z�<9��H1-a4�y�O�N�R���9r|p�"�~>J�^_��t��;��q���R~����]y,��㲝�0�Cq�����v�x�l�Rfa����g���_[�Cj��Wj7�;\��Tʫ��N�X.nH�9�7Սn�`��Ձ��&3,x8�(������/�y8�KU��c͖��.�"R�,��m��(��X�=Q �/T��+�8����m�˭gPE�,���;~_�������>��{�9�b�B:Yٗ��������Gn�����O΢���L�`��P�rJ����
<����L��̩�x���ޏ���M��ܤ
z�G�ͅu���;O�
8sⵝi���+���
��>Ax[t=��H/����0���t�;�HlP����̴pH_�{�2�sM@�蠐͖��^U����=&�\��~��O�iYp0#���N�S�:�;�n��"�k��gLUa��� 
ϳ-"�=l���?�"�ʠu�zy���H�q�u <<�y}���7mkH
^{����80�QԵ��1n}�C��A�&�v{fО���b�}i@��N�{�~Hy.X���y��������w��&�� uv����|��C�8
������E_]*0����tw��ϓ�$�>Z���)�2d�7�}�s��U�/�����D��x���_I�|w�}H%�`F8Cs͡�J;vX��\���D�p��Nd/����޳n*�#��8	���L$����Ҋ%`���}aɉ��0��~"���,.�e><������
3 ���@���T��7�xxdjG@�0����6���>MņE��ּ#�� �O�	-'�;A�%�El�m�4gW$ڬ@ g�	�����o�+��+��sTy���8��J����<�x�Q%=z�������^�o�$�7Ԉ�atƟ �Q��2�1����$%��� �"ZU߂gۙ~F>��px���.�Pa
H��SρQ��%jO���N�F;��0^��6�pe��B����Kc��o`����5��`��GN�/���N!��.T��k#&��c�.��J���#�"�_�\3�t�������q�,`-�8��ũ�E7g2e�7" g����?����,�UvEv�]��&�g�4˄�	���-�����fѺ�$)?<ý�7'�W�V�Yj�⏦W0;?���|FgW���T|�G���6~S��ɺ_ ��.mZ��㺊�}I�Je�N���~)�2�ژV�����f��l�-͡�Z�g�)QL����r��B�Ɵ!p��P8"Y*��j[����Ar��Zù�Y	3yt�7Բ�g��&�lg7P�fݛəd2��o��<��������A��]/|�:��� ��p�QE���{�%`
��<HyhR
��(��wσ��Gv�3%��!�]�.)�f�
��!M�YW=�8�q�<մ�(���Jp���&�vnU�Mp^��ݺ��23F�ٸ����,�c�-���ƤٕY�{�X�;k�Koa�������@��6f��O	@]=���˷����)����`�2�eY�/��z�l��X�0��	i��F�hp���^��쁪v��Q��Ʊ\��hτᔇJ.�a�)S���)�g���g8@�\�uo���b �R�����ukJ�n�) l����_��M��T��T\f(��s��,�ۼsF��ܾ6l�wyn���K��I�J.6_4y�`*��2E���>n�BL/�,;H�;��b�e��?�䡇�S�뻲���04(��v��y ��<g�y��V�PP��+�Xwq啃j1͏�-C_I��<���櫍��h=`�\�K=�r�f=���&��GWrً��|ئ��CmY��y��>�~&�β���=����6$P��"�#h(��xp���>y�M�i�
��7ʛ3X3kHF�X�Zik�f������U��vBQ�y6ѦY��y<]���2�R�}�M��Y�i�:X�M�{o��o�f��(��xg,K�'c}c;Y���+Vɛ�@��Pyv�f��C������I�����7��rA|��0� ��@!�S��:�l�����1�6�L���7�,U�4��m���Ԫ�*�q�D��ݱ�F����q&�B\6e���pi�t�Cv�&��!�؝Ovf�d*(W�D!OBE�\�J-���H���ښ��ڔ`g�Ŷכa�W��.:]�f$��yV>?m���x?n��[�iF=J��#��뾽�'�m�����(;���Y%�z�;�>�Z�p֕�ԍZwI*�Y%�/�h�d��(���@WX��wQ��4�Nk�|��z��'ixĳ����u�\M}��i�i��}<5�3|����l��|'!�p�F4����Z��"B+qϲ�	���DK^&���PM�^fB���Ì�MH�g���H{��/�V{���Q�����Atט��h��u���[vJ3H��ĉ��S4��xS6�ѸL�d��D�S�̞��x��MK��;��R�&���x}i'hW�d��o�`�.����	T@������� 9�^T���b���q��kཡ���JÙ5��F��P����k!�CX�����ҩ�J>�<�nW7]n�����)�}�2İ:#��P����Wu.g��$�6��9��>,����0SU,��1�S����_�q��r�Ag(��O ��ֵ�C��e�|����`�1I����*=M�v�k�C����J����ƾZ�>ȁ�{7w���A����n�L�kȬ������揶+a��Vq]DZ"S�`D�c��y=�z�>E��l}V��:�?]ūU��k�%a"�I�e�恃�9WM��k���$ל9��J�P.ŰY�=M����ap�v � ��Ե��.h�Q���v�u�Vǁd�f5��h�d��xN��j��`�I�e���)��������ʰe���Q�&�@�((f�>�l��%�Hz�~}	�~�HX�x���e��\��]zrଈ�2J�^�c¤P����q���I���Rx�������"r�����ط��Nl��
 �jz��`�����Uz(\q��{�����T��Jf�]�����ܥg�@
��f㽸`����0�����;�"c�F:��[m�f�H���`O-��8H��Au�����3;�2�^+���4)[kFaFJ�ZJ@���������Z+v����y���z&/�����$/�Gf���z����q/�>�v�v�2WJa:�U� �p�+���8���,����ڸ3;�d�Ս���?:	�1�az��`�w*��>M5I�g	�����Ǐ<��Hb��s�O�c�1F����FBw�/�:����pk6��ܡ�Sj��>���-,�o�8�Ǌ��V*�sϦnלI6:��7e�#�&1�C�vIX�J]>gG T�7��i��D��7�2��Ycݸ}�Y���վ�
�s|oj0�FJUQ"�|���DGm09v>p�j5U�i��=Uӷ�˒l2y(q����د�'}f�!>�Ƙ�������tP�O��1�E!N\�]�Z��j�bC�;���Ql �e����en�����oϠ����չm��٨,�o�0M�k���}�Dϵ�~�5V��0�a�Ƨ;¶l�����~X��2xť�~2���7MMt-С��5�p���j��L�gZ��G�z��3�󶻻#��N���t������G=1��3�<���w�꣉wH��ٽD߂@�v�&�=.���{�h����Բo<�jF�%0q b�I�M_x��4�[�����Up_k��K���?�r��jW�����_�M���,{��P������oF�y��� �ՕO��=���Ѹ�;��o1Oƍ5n!;��?���tLCQH��:��(���29��Ep �����(��#5�����7�Yh�k��p%p�N���.+m���|̨X(�4�	ZK4%}��t����?��792k�>�å^3�N1�xQ���<�g:��!�d��B;�,��K@��7�+R��c짛;e����s-��a)�,��7��N�+㓭1֔��l�e�[�D&�2���y0�p?�f�%������ژ��,Q�᠁��Ws#�N|{;�U�w�)3�mY.�����Q\^��v�W���G)����V�PS5�OSWKmD�z�X(��tiUÕk�7\��3���J[B̮ջ��:��M���&l�t�]���9M�V����Yw�(a>��C���b;`��Y�m?�A�C�
�;���5�Ρ���>{��z7Z��Q�#�c��6�����=>-o����Þ���� �承���"Cw2Tz�܏e:M,7ɖ-&X3�A�i����S�\И��[�v�J��9x��d��)�Rk�c�c�swA/�ucF�Z�3k9Z?�f��0Zj��l�ɾB<��R�ڞ�q�@q#!�q�M���A�H����M#O��)3Vԩ��k\'o�Z��u���/m�a� F?=Jq��f�ʨ���m`y��*�_�s�\�4#�8%gDsqk������(�ǡ���R) EÊT�Z"�6�!A�gG���Z�3B`^J���+]*>�ϣ����b�c��M�"v�]��d�(��	q3eC{H���T��^��\$��Za����PY�HP�{mf��PX���h� ܗ��⦨�}v�V�c6����� �a�j��J	�[쑗�����Ҙ�^UU��J��.1R`E
�|�����C�q�%*t�b)�K�l�Y80�u�dS$+��+�	�Xc��QK�#_�hC�`���P�]��v���k2����Hs3�-��t���q@�4��f�y�H�lu�U=�[��
��(|�4lPث��Q7��%��0Հ*W��MY�.��v[����,2����4�5� 9���JJ���KiM���٣6�"ST�cv2�����`��4uᢽ^�8������?VL�U]�8jx������L��U����])q����q��۶Ŋ�~�[��p>��O[i�$�e����:�q�d���]l9���Z1-q>��������/�c� /i����˼f�ֶ��ut�)ϚW��g�h$m�W7I���16&Qr�cѪ�z(�ĕB��.1㛛/Θ��[�l���Y�&�G'��Mi����>/T���I7�wj��Ln����X���F^���qۗ��"�K]Cԛ��k��z5\���%>#�ĕ�@�?lz�De�tlJpL�HW7�?S��ӛDN�p��P)����kb��\qiʾ�qe�˛N�Z�����O���H�F�`�;J��_<m���ғ�[�,�#����J��	�\8R�K
-0^��mR��N�(��V��hl\Es��`�%�X��
��I��؈��h���J�Ֆ�������;�>Y(燥�oj)���m���F�(�f���7�@��H�� ���\!���FA*M��ĎA/���B<����:�.��K)Aa���p��TQ?HE}�[�ƌt;x�- ��������ޒok����1��>��tw@%>���Q��V�db�V�(�nܶqZ05i1���v��4��v�H��G|��ZaFxO�߂�ӻG�;�o��7�
��؟ �\=f�{X�%�*�_c�J��hm��r2��p ��2k�γ������B!��Z�b �Ǚ�$Ě)7y���:���x��(��;�NI�����e�'�`h��U��.�6��@�
Y�(A��ˊ��52�]��L2鸴�\��e�f�-����������O�<Y�@\�6F���D�٧�FEO��� H��v�3�Ȍ�D�㖑��IڱM	��!�*L)����8��4��LQB�V���ɢ�Ň���6��f�k����mŅG�M�yn��բ,��]}��$��a�_����~����N#������Wwt�T¾�������z��-�V��u<�*��/�~/����e��3��#R�9����~�:f~��� ����Hl�e�4,L �L�[����[�Z��o]FM�����`0_Լ�&��@��6���>�ֆe������6�V#E�7����H&�G�%ّ�@��������^���`U��s�s�ք������*�q��U;ƚ���(D�_^����+	�rc��'��r^*<�DTy88�@w��J �b���>�b�&����ul�2�ci�/#_#���ۋ���Y�ʬ7M:	W��D�Mu��|;ҾP/ .�����k5��o!V��s���W�)	c���?H+�� �{N��1c�O�`^
"{B�8KOQt�fO��ˏ?��e[9zF�HL�*�fj��"��jA�?~�/�����5_o"	��{7�H�򔱣��UV�&�+h( �\����ߡN�F�k��W�wS�z�4��vn��-t�����6�a7D��	)�'똲���2��J���H�E���h=>l9S��7�O<�y��TX��d}��5�M�.#�:4��1w�y|.�*!`uc�&I'Y�e�Yvv�+�+�'���//�<AJ(����>���	�D�����?���b=�d���������l�����J�@�5�Ġ�sp�����u��A�V,g1	�������]>R�ִ9�Sq��:�Y֚]���^��/^S�{`�A��������9R��u��O��������C}��G7������)�Qdb10	��L^9{@��2��e3>?��p�}�OSRd��{��K��:�ݦ��@�+����>Wa7�Z0-j,v-����4�����5�5�l�"R��7k}��DP�2�C�A�%.r8Q�s��l��J�����- �mlwϘ�M�u�Jp�rz6܊)�ѣh�(���v&�_ܘ���l�S�(J�8%�j��nڌ-e}��ف�&%��I�`�ؗ�Uk��P��3���I��P������� ,��[��]bhףJ��vX�X|X�q$͂�������G�Z=�"��Q����]J��-�L~��\}�WW�Φ��q��d��?W7�}ȺA��wV5�K��^T�@4I����Œ��j���d�{��E_�����M�P��F9�L'������Ⲽ9��@zoͬ��5#--S;�g��i�����E����	'���C���~}u� ��0`D��Vb�耱+�~�q_GTs
�_`alR:ǚ6�O������Bg�K��)a��!7��#�{��[��w\�_����W!4�j�-}�Zv�=�)ȷM$�Y1��A��^��{2ֲ;��Ƭ�O��k-�Ӏ�-P�L:�k��h��IXq�)p>��R��� 0R=�JF�ũ��u?��Z�C(/� �r�{��^C���� �5�K|t�W�&o�縴F�G�R��5����u�E��+E@0���^a:�<k%�<�8�L`0[v�r�>��/��
9J�K�&�M�d_�T4��7�]%pH�RR|�I�7f��J,��:Ү�I��
�;nWu��yv�|�%�1��/���W�Qg�eo��0D�Rez);1K�%X,c+K�$�eԳ~:<0�Q�	�˶9����<]��6��ٝ�4㣀OT"���T�R�h�ŌDM���q��@f�?�mD�a����+�L��b Ȍ��^��Xb�=z�cs]X�$����>�Z�*=��Y�n5Mn��+�O��Zc���[�
(���T)����ҾI�V�LO�z�3ۂܮ�,�{�Mi����p���O5~���)؜�Q��o�Ӑ����i�1�H9�r@�%JD&pjqn�l�J,s��#�͑ԣ7I�F�)�'O�W�Ndc����l���$�zq@L�xm|Ԕ]��)��X)�p)�r�9�Be�J��x a��J�n���τ��(�yv7V������'@5r�Q�~1w]��b�K��(�a׺�{�﵅�p�����l�4-#�,Vp���p�ƃ5�q�s���V~�;��s��~�3��zN-�(� �<6�8�Q�B�� �UӍ]'s�0X�g�(��h�ㆉ�����k}�gԋm��\;>~�ڕ�6
ތ-8e=������9/�|�רӘ4�������qY��������l�6�z���} ����-�Ë5��ɖ�iu�Ѹ���A1�gC8����vϣ����\b�����s�h��{U��UY�Bs�؜]����5�N�5�0����{=���X~�Q����~��v�`ޕ=ސ���s�Z���і"S.��,�A�S\��q��x�]E�EWn<�C���w�UZ$��1����o�Ի2-4_�3  �o��fg��=W���%i
aaH���'��L'	'�9XU�O&�Y���t�t�M&^�x���W黳����χ�w�s^Ԑ���7N|��cĳ��k��,�/���S�U�:�6�*Ӛk��䮙y0qRjP
*SG9�C�� ;h� �YA�5���i٦�T�\v����c-��,������B��`U"ken�j�
�L6U�P�H?������A%(_'��t;Rz|�䀺�w�ٺ�Gn�B��ų��y�����G�IoT��W5����,����u�i��6�i���=�������,�/�%ؔ�x�On�.�@38?=�~�7�`
�e]�v+5k_�;�T �Xʩ��t�hL��Li��~l:�vG\h�_NW!���=R0K��m�&�`)�:J�	�Y�$��ђ���}����T�^\������,���L>�nwp�(�t�������b��=��r�Zi�Jԑ°d�t�x6Q7'�Ͼ�ť˙�t!6.�{�Nz�O*a!<��n���2���~1�q�ϟ?��>Y�\*7y�^�i+\�?��~��°���zBX��)%A��jY�&�q��V!#�'�d>H��7!z�?�2�v訂^���h��d�ir�	^��r@�iN�	�RQ�Nѱ{�\�(�M�N�Y]�KQ+�z��K{�����Y�9�u�Cpe���z���^��n�]D˱F��2]i�����r{�H.~��8��,�����oAs�:3<�#&�`-~e���q��(�]j��a!��U?:+�%2�D�A9�Aj�&�����3��#�j�����@�� ����2j~>>�ii>�b��¹�
�Zzѭ��#ˏ�'>�1��^�{�EĽ�g:cm�u�Ī�n���m��-߬6�Y'�q�>*i��uܠ��t��7Ѯ��$��T�����.��{W����Y�D��qGv������NZ����F�eyA�U� �%�ɲ����0�ə^��0*�Wn�K����/m��ȑMU���gfw����a{����v���d>���7�jW��T*�y �@ ���#��1���3��<)`-�3U���_����V�������޿|A)*��us��c��QU35�G-<��^��1,U޶3�͹�����+�Ed�7�0�aHc؏.�=�l(�����JH ��qR���CM�4^�m�m��m����~�����?�I�)��F�ʽ���ȸ��3�[kk��v��̂�9��A��H`�R�l�gޏ"��]��y�ρ��LD-�����X[�j�ٍ���'_�!EJ�؍Iy�P޲����ʵg�wo�Z�l8����u���^��٘�:!��y��r�i���֟�<t�g�����V�KA'������6�2�G��K��<Q%Wm�}ޟ�x�ϻ�~�=w�$)7[���I�%Ze�}��Zd�C#��g��Q����C�!B������0���X=(h��Ҩ�V�"�Zuk��$®�)嘭�'��Ʌ�X��<Aq3���?��,u��)�Yg�vnj�v#�	!��x}��X4�Zyb���Bzy��^�S.<��BY1`�߿b#Fk�ی�ׯ�^��:�b}������{�����z&}��&}R��0�4(e#�5Ee�p@�����V�S�n��d�;�[��dي
c����ۯ�q����/���`"�����EB>ѓ?/k�*U���z���i
�ڙ|Y_)X<*T4H����`\.Y�4���S�,4wJ�g(y���SW���Qĸo1�0����}�^;54y��s��� @����&wO�4'�;���E�<c�*C�qq&V�е�������(���&��3#�����rm���d�`�j="9�vD>6�r�M/A]�Np��cܗڔxa����t��]n*� �+���["�Lt�X<?a�iB��C��Rق�d��MiW���?7��} v�
U����� ��q��d�j,([����C��K�PpU�@��W��B4�ͬ��f� ������}%�z�|co�%�-7w�3�����z�)|#���z%��{ŏ��n~�W>�*��Ȁ״9��[��%k�i���a<%�熀I�r����Kp�p"�y�:=*h��d�oKg�w9-̻g���ˎ��lz��s���l��fHW�\n��?�؍�o~���w#���?��)n���n�-O�:uyn,v���NؚtU!
>6����`p�ޗ����2�N���!:����(�=����,<�=+��yzF1�uw�}=��٘S�_�pftn7D�T�[Iv��v{�Oj�U�����ɤ�����0�1i�g��G	�W/,�!�|�M�lݛ����{�a؞q�qw�����m�#�vW������r��Wt�Z���¢�*��ȁ?��OQ��a�k(������Rr�����|��ND�3�����Ϫ������T�Y%�RHr�`��-��ƃ�����`Fˆ��%��	$��i96� �`|bA�g�fD W8�4�$���{d�'��΅�'b�k��b�U����[kX��,+��-6��������Ðz�Ӱ�siA�N�����e�� zf&��ؿ 3Z�`(
N�T��m�1mL��Bt_dY��6��ǁ}^�g�1q!��F��0o�Hq������/|v��2���+�ӈI�(��5P�j������yp��=C��qſ��Ĥ����G���7:t�%�`�9�x��.h�q��>�*�Р0'4b`� ��#*!�%y�77^7
4;�v��<X�h<��C1��gJ�|s��8s��r�>����G�ucJ`7F��AC���Ǻ\�h�>Q|�p�F���=i���m_��?w�P�E�h����W5:��0�4e�Y�v7F6�E��'����SM&�ϼ�0��^�ǅz��	;��-�Wȑ�'�I���Z.��� �wt眨`�����f������޽}j������mC_�>�}p-����N=县��;5�e���As���$����v�$�����UF�����*UZ�B5�7.y�+5@����,��,.E �I��ps�G�έ#7��.��mv���a�ipq������BݟWX���!fщ�N8P�Ѡ���c�i�>���>��������� ��o�����?���*�����G����'�왑,�ah}�m�Xh7����{dF�?C��@����:���D²��D��y�=�L6�g���V��ye��w����X�}��#L7o��4���+�����6�N�za�ݕb7sp6��Le�7>����)[}�[o�-�W*M��`��{��
�����<B0G����a�r>N���#��ןC&���e�3��-�,l_��ܸ�u�Jο^ d��Φ����b�׏�(���^������m�21�I�98-T0T��߰�:�$���7:~gH3�υ_hQJH�Ӭ�NU�X��%�m�ZӐ�f����&pdIW���-|��1#:y��7��t��[�(��B�ejx瞱y9nH������n�vb��6�������Y�+ۥ�@��9q���4�>����|�	|,�7�7�lV�Qy
��V�f|�_�O�|�M[_�d!+��I��ֿ2����+�k�)��i5
�%�i�H�B��p��<Sn��&��{cڴ>���}@�fgb��@��B�H���z+yR���cK	i�/�W���%ʐO��{��3�6^f������s���F���!��P��3�K�Y��8#�	1x��/��=Cq��&=����P��C�(B#�EW��
f6�vc�A�����9f�S��ʂ�l}�<��ȺXٵ����9����Ma�o��
ÃPO�u��!eg	�}"�Ƣ�;N�	!%h_�
8�<���̲a�+�|���Ys<l-���dZ{�8���m�M�Ġ�F�Ml��ATы��w��-������%�W���e�ģk�}z��C�M{�a8÷�J&P�#=�"ch���Ic1L0�x!��O}#����/ho��:�(&��H�)js	#J���/��ed!r<9^��"\�:k���>�6��D��]�O�-�g��q:m�R`}��gv1��� C�N�A�oj�n�Z�B ޥ���Y}$嬌o���ɕ� �c2w×���R�*�U^��/��nՐ��*#�<�N^���<:MI��8'���o�~{�[��������ް��ܓ���s:�c7`��C�	������+��|����sҘ�H։�kt1Z)f8�pb[/5~|����u����*���[`~�4��=� �y��mjWf�}�X����B��4Ҵa'|p���M�"�1���S���9)7�I|��F���^R�x���"����5�����W�Y��>��=���p�z@������u_�����i��,#5
f�=�����߽Ay���O�}t�u�ߛ���P4iM��<Fg
S�
�����e��oN�{y�*���h�H[Q�o%��[Ң��)0�!3���FR�V6��K�����-�����Ҭ�-�'VmL���ې!��yz��1]�	�}oh�<ٗ3w�����4��S�� ��ܫ5��pƆ�#3���0X8�������%m�	$d�آ���@�uԈ��3��к���T��N�f��ȞV�9��Y��ɍ�Qm`栭}`��A��q��!��3��=�Ep'���&P��>3�w��O�O�G��G��[��po!���p6nf�:Y���0���T�4d����޿{�m��c��û}�~�:���.�
Z�׺�:�u�9�k�q8Y�0[�&h���(�ܰ^�Y�P(a$v[^%7q̣��Ek!�����vO<I>�	E��ѷul��%j��9�������.D��6&���!Ltu�)2��Ǐ����}��}H�gWQ	Rgqʣ����>�ٲ���`����޿������޹�C���ݾ�9�\2Ac�i�x:E��Cx��7y���<���P̎/%gz3J���T��0Q�D'����%7;�wѵ`J�,�D��k��p�<�"��q7�9�aj�_Yx��$O�ps�s���a�RGy�g�%g���28�<���2�O����.�lz�o�B�"�T�缩F8�Gц�33j;d�����{��#ՂΩ�/L�� ����I�U	@�,�C-:�y�L��ϖ����y�D\zεt���۔<�#ܱ��ƭ�zg0P	;����^��p�F�vQ���:�ujFTl$8�"�k�pgE3n|m-M�o֟~��x]m���\�9�\}�0al̀{����%6ͧ&�^�T`c7�� j�[�����
��6Cݷ7$��&�8{c�{v�>�����j�ɓE#X%��^�qA�G?`m�^/�<q�90��mt�h4�N�ʪ�-N�X�9���t������NH��8�NT����c z�Q������Ă8�_�'����_=�����E��
*�4���5g�
(xݓ��T��^H�H	By���aP��h�Z�lG�Ոv����L�!�X=˩���t��5�l�h�����?�*�Dv����{�`xRo�-Ly����4p7��Ƶ�t�Q��ۂ�3:�jA����}�Ήu��s���I�=E��|�/�2hG�N�+�/Gf����
[]���@g��-�9{xk�=< �r����o]s��i�yb:`{ �m�Ĝ��\<�(�I���H��0������p�qlA1:o3�3�X+bDR0B�����I�w���0��Ȍ��Ó{aKp��;U��%���(����D�WEж7�HY`"������ZԿ&b#�>��)�-�2ڞ8gxui�y~`}�l1#T��^��^u����������0B�.7jFG|���G4���sim�}-�ky�=pR�i{�7��J�#��߯�؈��H��$��A8`�ܡ?�H��DoU	#D�b���[���@~��J ���e7�����g�Kpv^$�ɦʢ)V4�c������z���+��+y�n(Ƽ
:}�7����yF�v-��=B�����;�n���p�ݛ���π?4e��C#{ 8i1���:�i��c��#Q��M{=dq�@�[�&(N|�`a"w����96�NՑ��#[A?==��2#j���M�~�U�J*US�ΐ���x���T���\^pY	|Y	��xr�2���9��;��:GP[��� �-~{�'bkW����VϬ��L�������p��`%D־$�(Z3�s>�x��,�̵yТt�+��[c� r���Kx�H>9V�V*E��d���ب}c"�%J��|��y)X�r=Z2��?;����zW�[�]������ G�R�ݐ���{�0#z��0FҦ�x�)�*x�5�:���]�-q_a�g� #�d�p�hl�e!5��P��6%�i��4y��{���σ�#w(ͬ�Z���DuG�����<M��Qc{#�H2�SdWiw��a!�����l��ϤQ<PՈ��S��{��É!C�M_���0t��鑊� oQ�BKCz˲V0�2��L���	�V'?� F2G�8Hԗ��<�d�E��C43|� \0��Jm�:�[CM%#�dU τ7,����)��MyI�����j�Zq��mSgʱ��m��w�W5A��mK����:��ptA�Ul�k�]Fo���H:i92�'��(���>Oy��M�T�s���q�+��`�<x��@��IQ*;�<��!�!�v�i$���z�᧤�I�F[='�
���u(���9�������M���'g����̻g�-�o��x��"6�$�^[�L�	����g 6��+�������o�����^���eY�V�]"*�i�=�C���x_$�r��ॗ�h�ύH�#��K�b���3�b4<#�u.f�N�uh"i��D���mH�^�@�y����=d`=zΣ}	*�.厪�=��@'�2�ټk
�����]p�N�4Sx7G�8Wax��I�q���V�U��3X�\E%�l�-hpQ��6�
c���X~�s&#�Eb���	��N79	wD�F�u#�d���U/s�Ԩ
�W�5���Lj^\&�f���]�Kc���
�ӌ��n���T��;R&�n�Խ��x�H��!�N�1)F��R�#�Bh͵ḭ�%�P���8�[��#���4ȳR;(;�I���HN-
B�|������?0x�V&J�e/?�G��@�	��)@����h�������X����9X�yv���Jc�1�����i����2J��:�ʖ1ef~+)6�ؤG(/�v�����gc����/�i�4t�D2#}�R�<R�-�4Gخ��]�w^�i���M�SQ����7�g�yIj�jo�J����0�j�!u'�<�s�qH�C��\a�s����C�7��Ux.O������
*���7&b����3��l`wn߽��%�����Ql>-r�\A��~��S�}�(c�ߥ�g�d�S���u2a�-<����G����K�9��U	֜���-�*b	O�Y�$)���7�*d,P��DàmM訵R�y
�B��3��s�BR�mޤ�a�7�qg;�)	�Ф���(��	X4�-5��w���5Mم�x�HT�C��>�{3%)��>8�IQ�*�&�[A$1'�F�ĭޣ��7�Se����~`	��_��3C
���zr'�Ƴt���3�?���7/9c6������!+���2;��k�xW�R�h��]؝{A"�2숯-�<Ƣ��!	���$�FId�4ʲ1T��	�V�#��$��w�Jq���~D��ϖA��VO���S�>�<�2���4�@�|��]Ѧ��ww ��N3��R�1~Y��$ޤ-�f������C�I�L i��3����{xP�X)6p�fh�I#��܂���p��P�e���u%�[Tȵy �cԺ5�;�m���5��U])�k�=@	r�iD�xOS���$�3� ��S�4�C��hz�qǹ�o&��������P�^�?��(���qO�8�c���-�8T^	m�(b��?���b5^.jUn=C{�/����h�dr'���@t�x83*���: 4/���@+BF�8��	 լl�c$�!%�|��c-hR{O�Ak%9�'�39��!���}7�xː�4@�!���N��� �E8�(A�/�a��.��^ANsn�֎�Qy��[����;�p���B�����m��Y���J�<�%��ͳ�}�m����� �Q58սt�1�1Kg���8�����8�Q��2���)��$��r�vY����z�۩b��b�g)��yM*Q�����#�3c]tz�8l�^��)�����KƱZ���E4N�Vw�H2�a){%�+86��Ǎ������W�N�����B}�v�\�Z��DBx�~�IP�FM��Z���A��{�K������@� ���$�:NX����{C�&���9ZIU�^a�?�au��h/��cՂt`V
V{З
[*�$XMkU��A�z���}�� ճ�������?thB��@@Z�DNʁ����?��b7�J�"B��.$��x�4@���U,�!7����(9�qJ�%<��'u����I�ޗ�4�M�'{���n��ԾV,z��
�:JJ�jǁM����6�f��զ�yf�IoC$�tb&��l6[E�������&~'.����D&_�(�;��q7�,ȮdH�$�Ҙ
OU���^�u�0e�5��������5#I�dc�J����OO���׵�1!E��v0"Cs����n��#��4<�&C��:zE߷ɆCv��r#:�G�`�F¿6���~��`��Q����%R΄��d==��ޖ�)�=N����EY���>��|�>�?��!���v�lgL(a�M��J��x�+'`���քl�HeK�a2�A;02�+�H���Ƽ
`&���\.�L��q+���6Bq�C3�FR�t��j5�q��\�)����ݝ1�F5��*Y�Cq�&+�!��WC��B�c࢏�TV�#��z��^<
���Rq%�J́�i�<��E(Ӭ����rS����[�ҹ+�RcM*Y�O��<�<ĸ�@��6��'U�V�����k��������O<S��ږ�m�$B`H�Z��,����H�5d�����aY���;-�O�7�uO�^�����6��Q}��%
?4�0h��m�;��TK�̤o��%Ӣ3m:�{� ��C���Բ r��(��(@ˍ�G+�4�h��F V��=$���=ĎO���#T��a��3(A3�Cv-,�%J�[���%nM	N9@�ޑpF��i����n�� h�[�̼���GF��U-}����-��j&e�� �A�����0�����xH�8fì�T��ȸzB�8Q�AB�[��9S�t����T�觔?:E{���~��{�!��̆*a��"�- �,䏚73O�"g_^�d;,�X���v�Kȃ*>^�H>�JxGy>=�<S~K�=�6����Zp|s��<B/ �� �9�fԷԝ��������c�)��6FK��^�F5��A�2�%1��6��,T2��! ���b���&r�k8��vzc4���yX��TEKx��2yqv�� nA�=��k� ��(D�ׯ��?��B��@'�E���/1�G�֞�=#	�C��9F�D��	F�� (��l��L��Q4�SOf�'��|o�5���MWi8��rⳑ�Dɹ+��:YE�{��δ�׍�ajJ��nL2i�jj�{���5�1�����ݰ����Gvf�S�n(ڷ������{w=�$�Z�bH��Id�<��tC�N�(�|
C*��]Va��	*������}G�.�ą���F\��k���S��=1R��!A0�<����d�����P#Gr!w�ŧ�f�Sd�'ǝ6$�DAѤ"���l��Z4�ؤ��^�������X�v#�(#�F��U^u'�B����$��"c*O��j�8�:���C�� ���ѝ�ɮ����S%��^��%ճũg�a����~��D�I�sxB�<���sьi��k��`-��XDa�]�ЁG��&j��P� ƺ����V��v��|hNk�}evx�Ŕ*W�hS�herb�-*������h�&����բy2�ǘ�W=�����?�P�*�ݸ=c^"z[�⠇���ᗘ���W1�5$���Fz�7�G�a5xZ�Z��PJ�F�Ⱥ�p��df�B+��3lP�����恙껌�7�s�9�012�O@�>E+ZK�l���8��$�:�)^�� ��~��; jo��,A �B(��l{�t.����k�[f|��sy�6.�^�Dc
A���z��tW���k���d�:�^��v��|�Hn��	;G��c��l��5��WHә9�����E�$��Qk:��0FX/�L�򴭝�{k�/����GO�̱���� ('U���	��lTg!f���P��Ȧv^eա9��.n�!J
���,h �<��њ��DʖXC�ڿ����b��T���}��'����}��([�H���CKy�q�m�pf�Y�ʵ��	CzU'��B����R�f��
Iއ����h�� jeltR`������[��]s�X�A�;&��P��+U�A��W�BA?Ո�Af-H��Ha߄�:K���KO,�O��M@c;4M>�(�C3/.��Cg�	�5u�����������{����6y��p�Ka4��T��B��b�Y�į[�?.�s|�)��������k�x�(��感�ћBW���_���mI�1o�_u�_�$���͛�5[�Ki'2�!��7��p>��?�Ȏ4\K��Ʒ���-el#O$�7z�"�CUI�Y�X{��V�14�5�Fy,��EXG��2z���}�hG��=�k��� ��4�0x��ؕQG��W�20���6Щ��a�b��ځh���4���#y�à&}		Uj�C&6�v�l��(�PQ��	&h�"#(OZ���RS�B�>'����38��w�lBle��u����fQ8�2fs6�T��u��E�7�K`��9�U"?F�#�v�f�0�V��9K��f̈́��m%<�\jϮo����OȊda�?sQ�@����2���Y&�,��-�"U�s����ނ��Ʃ}ٝ��7�������v�L��?�P>���d��<M�`�~]=Awc����	��c-��� ,0M�NC�Tw�m�IS�f`��!6dx���� {��1��eKOk��B�qP�U6vi�~�}�PI�aǢoI��gE(>���kv�@�'�Z<Bu\G�|{!�֛B2�����3;(B�	�����zʋ��"�[`����A&�R��vm��V�s��7��Y���; *3�żj�����a�H�+�у�H/�B�Eo��|��*E�o�*[�'!+��ښ��Ւ0����*�.�fߟ}�3d�q��AL�8�q�!mgޫg�aD�`�5��s텈ak:x��l�;��8�m�z�u��~��~N#�Kl1w��I�<�v��ү0�ޙbY"
UN'�jFz�J��:�H#c�;��IB���m��E�U)8iU�ɕ����������]�u[�z�X�*̨�bx2麷&_�ᬩ�Xn�B��n�cxEZ�G�ֆ�X�Kt�;��&�B�ӳ��'m�ǽ ��\ST��ЈK�崧��HU�Dٺm�s��E1�	������hv*�IOlm�񬮁��+�sTC?�X��诬o��CZ��_�H�ܸP}�͓�N`[���1�FT�-���I��8������PÄ�AQ(�b�]ЉJ��Q�4�6$m�7|Ll�s¨c~|���!G��(��*�zk8��!�l����5x�4vu�n��L�Wf��1�Ps?�X]윆�|"�^�y�tj�n���9�{���HmM�Sb�2��\��}�l����'*S��ӲF��y���Lc�"y��Z��������0�7z�*���ƴE@t�:x��r�Tᗰ�Ȅ�@�:e�+��M#��j�<��h.8=+m.�O�)��N:n3͘`'Z/�����D���D� ��0�0$��I�$�F��da��ĳ�0��������|b#�=��R�����Z1]>6�� �+s��!զ(�- <*<� !�\ѫV�E��
��I�����uȠ ��KUіI7  ��IDATX�i���;l�y[l*y'�Pfpe$u�o�O0/f�Ϭ��}����M~z�c���e���,!���9ɩk�d d��"/�.$���qZeL�x:�I�5��~�t&֚k71D��A��	�')��u�t���Xɦk�b]HR9��E]�h��a
�^�=hs	OW����w��\D 4[L��֚����|��I&�o�y0�W���� q8S+֌�B~o-�U������=b3T�4,�`���zgZ�G��6e�E�PF�ɐ�W�c>y�w{wsj��+�Ѹ)ԑ'dX��m1�h�Cɾ;9ز�&��:��%�:��	��O� Rưr�6p�H`��-�s�t��g���,�qÚ:Ͷ]<��x��������M��&8A����&�`���!�P{���k۾=���%��Q�n��Ђճtze�٦��Au𾬋��񄐴�3����ɉ1�i"�'�D���G�1JhQ�|����;�q������1�u����$�qh���E$|�5R�*ML�T����HN��e?�.U4��B��yE1DJǵ���y�뚇?!�c�����S>/��+<5Js	?�']��^_�s��l`d4J�����u-rv����µ�9��lln��[���6*"���T���S�ǯ������s����5 ������䡆*��o@0�Ř��� ���֛����3V�.��%?S�\�����Ҳ��e�`�A&ë؅��Y��C�ϡ8h>PG��K��V>&ʓ���~�����C��ֲ�x��"co�R��� V�h\�2���C��Q(��?m�OJM�Wԛ�bÐ1� '��$2�s�;ٗ��J0d%�+�=ȳ��`OC�l6��-��F�&����I�B�s<S���ᴔ�����Fe��Y�����C�~��>��IG7v���zx�� @�p�9G3<;~ַ5����-_�7##i�#����Y��K��kp:O��v4��H�����o-�xKg��z�.��C�߾,�+�)�mM�
^,a�
7z]c��'�Ea�t�kX���@22�P�O��DDF�L}��m���������?����-O0�.�s�t�G���g����u�$1���<ٱ������P�F�s拶��b�{�ͤ/)��RTw�-�	}�a�����[���0ɶ1�O%�k�����Iy-��a�� �u���D�U�,��6S9j>��*�����fl�!�K���~������%F����sXn7z�p�2�)C�5�
w
%Hƻ|��2gC�0�g*�?;�ll�Z�����+ժTaT������E<���k8�Ґ.(��0q��8gba-��iH��J���%U�IF},ܭE�U,1����sx�)�T�F�")0�#�9����oL��?J
�%z=Ӡq��p��I*�t���c���q=*y��# �\� {4����2d.�m4��#Y��5�[�y��!lk�~����8yUC�Z�VB�W���ҷ0uc���`H��Bo��oƇ��6u������ZVǁ�#�����?h���@з�5z����68�H4y����.�ۭE@�p�<�HHi��_Z�<Ҟ*�p��"i��U6�ήI����5���}�/�a +��r�r>*1�	�]��� O�W��̓5����Ž�Oz3�/���U��u��0�`]/�gP���L�P���tM�PO>���-�pķW`ZBn��A ���M�a�杊� �]o�$k+��s�*7d���w\�-C\�p��1E�[a���֚������6��¿=d���e��~� ��
�ڈM%�+�,�0��$p��7��=���ū��B��O��Ao�煂�9D�;���s���-��_}L�0�}�γf�\k��;�u��qy8]��n�	���}RԾ;4�ԍ�9ᎎhf� c�m�N�2��u�>	˛G/�ņ^��K�7i�����H�	UG�2�m�*�v�S�y�7"�&��KV���n@�g�k��|�G�	3������ߧ}M]�����O?�N��^z�_�pb�<R���L̓�Õ�ɐ1�O�7�Bk����S��R�M^���q�k��=���D�_;�/��c����j܇�u�=�(��}T�����钺��~�hW*���g)ۍ�*�*`�|a��M�J+e�E� 5��~�]dH�4��8 )����YhZ�>4�p��	l�XJt�F�t�O��_�_�	}ޑImA#1��󔑓�r	�w�М���u�����S�2�gs�^y<\�؀2� RϨ�qxa4��r�C�q	CT��l�ǚڿW�=+�ҋ-OR�	�G����@=W������|]/t�j���(
�A�;��,�_)0����v���4�{~�\����Ό���~~��T��ӛG��"3�u.g��k�#������P��wnU{���5�k�;�f�D}fR����@x���;�i�XX��C���?��=������݉z�����),�m�ZfK�ݘB�BЏ�9����2_��1Ѥ9,`iz�����u��F�#�zuԳ�TB�xI�q��^���	�#T)�7-��v*w�:�N�$�駟=�8xu�]m��4�6֗�����׿��)W�"��F�:�������\e��)T�R�Ěf�>f��� XJm36�����"|� �V�#�4��>��w�F�*�\`��o�*��D� �
�v}��^�-.y ^3�Β�O��dz+m�GfX�gQ���p�*���uԈ�%44�Gz�`L�a����T�ދ����R�*��
#�O,���5덉R\H�����I�o��nkC����PZ�F�qh*�5�}}���ZJ$� �sp�ʻ.^����I����~{i�wO���Ș��12Cw{�	E�5�c��r�_+{-�5�j�������w��`1�2��7��Օ��F�0L��#�5և`����_����Ç��/n���/fK�pްQ�;�����������C���Z�$�x.�-7躙�����/y�Phnc�yl����y���}h�R��d@˟��^��K�a��X��	�^IC��yi.���ވ�9F�y
R���ׯ�a���z^��0C��<J3��e�C��OU�l�7��X�]x���M�3R�N�� ��^����܀���9��/7����]�,c�p��e%P��'����B�?)\-��K�]�~�Q��oYg=�1����eM����Rz�|+�LM�Qna@S��v�d�JIK����j򽷃�*c�Lxm�mG�/�'Qx���(�Ƃo=<�
�Zpd�[L_��A	n�XR�04�4J��>��'{6-�&e_"Yu��G��}�<{2����{=��(/UuYT>�C� A����*͸�8|��L��9;3��'j����;u&z��ռ�5�x7�c�x��}l��=��ĩ9L��~���K]�g�ӛ���a1!P�b��5�]DF��%��Ci��@�{�����P��U�҈�����GZ~,�u�����Z�zn����zߣ�xf��{��믿��Yϗ���/�/�y��_b�fVk ��99���~����Jr��a�����waM�L6������`'9U�D��l1�^#8a|��XsFï����w�֢0�Sh�<Ю�P�$�њ�g��]�����ſ�߆n�|J�ŦvbȍF���zl+�]/'�F�Z�������U����r�"�%~c8Z˔�Qm@�&%%}ٳ����>3��s-o��ꞡHT���\"lUqȫ>�HBs���0�K������j���z3�v���w����j$7S%��ئ�ac��q�c�i�&ܰE�N������D��,9N�ϕ�S~��-P[Ϗ�<�2�`N���P���k�-d�����kTP��I�G��u{����G++W����ٲ�\��a���k3�|U���0m~��Qdq�қ�н⺃(4��0�=�M�Rm�Lx�XU��H�SPVx��	~c�&�^����;;]^����^=%/]���F3lϰ����g7&V}d�����C�8v}����������w����F���mc�P=J���0>I�8$��pH֬�`d)����	�8�a��kT�}ߤXH��z�^�7�x�fc`��\l|�hH�G��&}�h���T�l��ӧO����ϝi|��э)B3`px�$ԛ�:����<+4DR���������?�I�+E�+װR�����K��MKt��p��e�g(��F��`7�-ɛ�\�?���G5��0���@l��q����~�:����?��%-Դ�s��kH��7��@M�"���K��"b�鑣*i	O��±T�M0G⠕;kk�<Q�u_��q�	�R������5���u�|�("�p�H��֋㵞Trk+X5�[������������e�SVӍ��yD�!�G���!SH6��GZ!p���;���.B
�?��Y�j��9���O��=�D-�f�4�=Rm���	��O���������o� �bt����]_v�?�6z�jG!��hS޿k>��D:5�`ߓ� �c�\5��Mrj�Ka�=��G���q��y��w3Z��ԖLPr�6�_��78Fy2�b!ݗ�����fs�H��j�6i1�Ka|;�G;&$������)�ky����W���PRN^�LOf���¸ps�!E���z9#��]�Bo����i&� ���G=��x
~&��%�ٟ��H�6t
�QR��\,�6B�'?�bnm�?=��6���(&����}���������d/K�(J8�QucQ�5-���нF�}�d��z���1} ����5hp6f�/��ze�9E�asCEC�?�W6>���԰��v��e{6;�?�Ǻ��ʵ)#)#�i�#�:�2R��?S�:���ϗ�.�v��1��2�U�rp��c@I����ռ{�#M���_={6I�z��î����mHi��*�7a������Ÿ�g��%�B��W
n���뿹�[`�^�9e�E_,܈�E�EUI������~>�r��(�˵$�m_D��ϕS5��i!�K�D� �lk� ��&c0�H@�QU�*�L�h f'�iM¨a���>���0��H�m#:������'=zMvm��|���>v�싿���/�^���+������x�dH�^�(��Ңe3��4�g����1��ȼ�� �	�k�2Tz��S�^jYݗ+=��d=����8E�s$���!<-
-�f0ͥ������땉�[%��~{+��^��u��(Eϯл���xE��`{�׷��y�O�����k���{sL��Vѧ&M�L�&��=������m|��Lv�i���:���N�5�~-Ga������� bm�Vig_�!�a	"x�ͯ���r0����`T��}�(/t[	�3����ڊ�ꆷ���^.t����M]��$��r9}utT}М��C�<�e�0�K�$|� yHCTGܖV�d���L����@��:�z0�D�����6ڀdr�Q�3H��B!��3���{�q�xo?.=�-��֘p���-T�ά�u��}j�݈Z+c��jr�H=����3� �Оg��&��D9RWό�~�ʡ3ͯ��Q�}Q�D��M�ߖ�{xs/�|�Y��+*p)l�^׆��g�0�;�t��%t��ل5�����a��D�V����F�VOgMRJ$��n�W��"�%� ���Q�\cy��.��J����n���˯�4H{5�@{4�J�g}�Y"���8���Q�7M��f�:g��-^��rhu�E�� ]��j�l^��Q{�ʧ���y.9.�dg���86F��U�﵃�����W�L�ފjx���7 *��{ ���Di�k@�J�����;b<с���3�����yH���P51y�N��>�!�	>�d�3��F�z7dcJ�-�HiFq�����;x���%�`�GzѼNYK��WL�M�1��&E�6l�~f���9Z?� K���oϬ<7Ǔ����*���<���fp�v��g������$~��O�{V�^<#M/��M��f�����/����'ь^e� �c���:�gay����:ƼO��_��/�+��g��&�!z#f��f�(�Vx�ߞ!�}y}�'o�����Ȣ���-�7��w����%�4�`(Rq�_�D�_y@���Zn�4���/~(��g�9h>nh�]���,���J1{$<q���Yy��0���K�A�ͮ[ʊפ��
����xeh������x�v�@L��<��m�Gm�)ǸO��k�A1J��phݘ1��[�.�A��):���3��%�?����^�B��������:_��߽�"l"��ipC���#[���`�M	�em^u�n��M告:h���rISw��#���=����Z�iu��]x>��k�d�غ����@�q��\��V���� �hQR^���]�,~?$�������"�ᚼ
UH��B�ֻz%���[HB��f*ʈ:#���#���U솰E��C�Ps%ff������B���l��R�kF�J�f�R���Je!�ί���;Q�⋝���y���gFv��+K�+��v���M��)��%.����no�}���EHףc*�k֍�#D�rTu�J
����^x���~��eU���y�9 �W�"�EGC�}�̯�53�J��>7W�A�	q��kO�0K� P�A��i�������Bs�x����y%�P��P5��mu���{֚ծg�{�)���D�a�E�E4j�\ғ��󢌗[V*0U���l��-��2��Ψ~���]�[��G/��H`�SW��?FB���bu8��������ҠNA�Z���=�\��sE_��\�����)f��=��RT��^S��ڔ�<�y�£�x+޶�N�d;�?���OM�<̓�K ���S��5���� a�虡��ױ��2����\�%��ၭ����b�F%N�pf)���"����i|��!��Ub)(�}p������1��{m�AM��[�������#-�G֢II���@O�젇	����tf�
�a�,��c$�������@!�g��a]f�	���8H�~
�����Z!5o�ڲk��K����%VJF��h�w^��*�9�%0�tK�J�9�nG*�	r9����%��@�q|�_L���(!��u,��,`��nٜ��O�(��>sf����(=���p�k������NB�i�o:�8�v��o��D�U}����⤩�8�R��sO��Pw��b�ѕ2��h����
��)k�O�\�2�[ܾo����ԝt�frJG���A~`O(�|�����qnC�w�a�a5F�V��hk�s�B(� Q̄��{)��j�lۖ���8M@�^�9��8�|�Bi�w[�
���.�Ր�[��T,����ܠ�ْ�^2�RwOc�Y�Z�ը��Sփ?��8�%�GC��gS)fXb���B�+�V㒅
��9��U��Ͼm�e��"��Yj�HS��{&�	%�	9[�/>9�f�،93��p�1�(K[39���[��4O�Dt�����6�ڸ�Xu��#�^vF�U� �i�g;M���V���+��9sb\ ]��4$�K�Ģz�o��k��Z1�=Ӕ�p��Z��A4��Ϝ^e����H�a���@^E͠��X�q�K'�,�2���QB(�����:�J�vC�ғ��������Ə���q Ӌ��k�R�H&x����y���iM�mv]��-��M�� ]*�Vd����u�j3���}�H�k��� LvZ?>2��jMQ
��Ή[�jt���Voy�(�&#�%�'��9�I��O�u_]~ϵ�ke�4��vǊ����K�	�FG�͟�Θ�v��W��&D��밐�
�k��eQd7OYJ�_�c<Q!輨ĒA�E� �$z�	�V}>{�C���~��Vf�{z���'�w��;<�G�*S��[��i��ѷ���S쯚?�s�%�j�z94�kG��� L[�8��;3s�R:�L�����/ѝ"<qFsF�b�NI1Wv�5��
(~�~�%M�&%��^K�����rE����^��m�v�1H�L��X'�H�4?����<ȉ��v����}�XB���6�clȊ��{��7��Ĥ����~>^���^s��p��!�¼�Fib�1�4�<�&�`&�����癉H����n	�>j��#X��t��:�Nćט�m�U:7���������<;�Nl�W�w=�d��Kcv����id��F,V�@�z)���HF��DWQzt34b`�+�E�����{Y�H��m�G2"l>�aa �����a��\I�fе���TIǳf��xk����I\���A�G�-�kK��]RnP�}�p\�>Q@&���5��������Q��:;:pu�I#a�U�M���ɨ�mm:���y��������
�1�)�7&r-
s�Cd�%A�Mp�][�����X�V\iv��ɱ/��g�z(��[4زMm!��CM���̪F����d�i CC�����nz.i8�ؚ���G�?K؎�{��G*�سm�_��X%�G՞�x�wϬ�>%~Dϲ*�(�o��񊗷��Og�������Y�8���3�	%��[�O��`����.K,kX��t�u�L�n\Nx����N�Ff
�bl]c�(<Jݣ_��\�Lu}m���� ����)ȡzy��J����N�ߝk� 	�d$����J�f�b��r<���|E����z�����)������D����Ycoz��
�i���՘�NY�G�q}
��E<�9���R!�g�i t�ߧ
܅�ԓ��R����DM�3�Z�u�q
���Y{�*���L����� 
��H�NG��o��йx||�Cv@�<��Z/��ER=�;���)�ڨ_>�}��������UDl��A�yx~H��G�L�����2߲�5� %_�m��n'��yT<L���Gc9�	���Pt��b����\��Sb��v� ^����W���S������"2��3e��N%X�.G� I쁈����c0=V��&X�y��Ku"���n����E(�]WK(%� N�}s�u�0L�k�y�<�J75]��tְ/���wWrŗ=z��F=�e�#���6�0���B�Հo[?&?��s��g|�{��ʒ�:_�o�9������ׇ����w~��g�\3n�%�>�/���q�8؄҃i�%�����)����X'eJ��[z�����`ֿ���u������F�p�������r��z�6��4�������gBQ�S�pc�}�m�}"d�P �w�g�tv�ѭ�����G7+ѵ��k9�'������"㋃�Sge=1�$+oA�pp����p��T4B��%:b�Sn`?y�,|șUD��d2K�pz�'�����dx����:��w*N�rё�~��V���������g�����}��'�PO�m��n�$ʾ[�n)������O���4�����:z`m�X�8p2t�xVz�Bu�Z�ў9�>�ث!���	+��Y�b�2˙���c���ʘf��L��`�3m��QB!p�4�����Cf��I>E_�{%���n	u#�ε *_�����Gf�o�>���1ƭiT�T�o��Ӊ��I���#t�L���?h�������G�r���� v��ri[��-��N���ƫr����!Ґ��ф�&UPϣv!�� �j�b����h�3��"��p��L��/��ɲ1Oh�-�"XF�*Ғ�r�y
�N�`hk��'�����Қ���B�����tcy�N���=y\��d�MC����*��0���%/!m�c	⟀u5%yZ�B1��� �2'&�.A(�M�kA0��B(+'���yv!�o��YG�µ{|̦hØ�=�+�����X�dA���-�M��e󨓼-��tHZz?�1���72���%��b�������px�Ej+B ��~�g�D��<Kz���g�n�q��{�����"1ha��̓Jx��G6�4��D0ڀ��|#�V{��s+I�i�}Vq�a����4E�DF�&|}��R� 8󠓟<��G-zC%8O����	����٘�uU�ގ��W�Ƒ��z�P�X
A"�P�d�{`�W�^��vO��y��{8^���y�n_,�`u��;�Eg��d6C��1eN�+�I�!��d˚Yx�0mJ�ʾ�^^�7�,4N�ĭB>���� ȕ7C��m#�b��L��4��Չ�M(��Q5S��(�[8YcTH�x*�'8�i�2#�p�+��D� ��D��� �Ao��Nb�L�W>M �[X�NI���iOz0�?Dj�8 nx���"�L�@R���(-�\�5�(0��{�&W�1Q9��Z;,؍ắ [?��D*�e��_��՚��'��uINȀ��m��ck��"9E����a��Q*����4J��FQ��z0P:���9��Q�]in<#�[��Fz�T1�3��d��=�Z��-9���T����@R�o�b�ʪa=�~���]
�����U�Ȳ<���n����
r�#�n�E�X�)��q(���v�R
3����?
��+}�6�۽I����gci��=�8�e�Cz��H�A�ˤ/I��u�`�p�v��@��0�cd�e*OpݶX�
��@FĿ�\�7s���	T�NWK��{�9�~o�Ǧ`�/�*��&e�;6��q<��	E���&)Wʑ�yZ�6�f����]��p��I�F�O��X��gT�",ϭwC�y��5=�X?v�=Jj�N���P��.
]�Ů�Қ4���צ�S7h=$e���y� ��H�� ���]ԧLؑ28�k+��V���\�5$`��Ud��h2�|eBi�k>n���l&L~W�\�?E����^��B;�ʻ"�DkpE[W��E�=�w���x�5 ���6F+ј��e���m��w��y���
��nأ��j�m�G�Y����a���x��Zmas����U�#+2Z�yMYs��}�ó��pT�Q�a�ڽ��H�A^���G1�ū��]�Ji���o}榋�~���g!�yzO�B��	?��'� ��<tk�e���H���np=���r�k�D�I��w��*.���=�,8�+Ac�&{�\������
����,�K#W��� �Ry�f�
 �޼?O}x�SRV�}϶�#+EfNl�@��>29D(�Q|�&�*�}��������$�
K�r%g&�G��{㵼O%��� �b(UQX��z_HL*�0��r0�v���8^;kK�yB#=J%�4g$3�}���^0�����w�W�PPcZ�������������t��VEj�5�Ͼ�o��&����U����R�"��z����Q��Ǻ�ٿZp�g��G?�F��[eõ	�/��G�oٳ�O��F{�U�\b�Xw_0��He_�����dx�ln�PQQ�O�62�epʦ4,eh'���
o�V_ؤJ�׾OlKb����BJ7�� C�F��J\ś�:�-�(*��(+F�ڽ7ڪ7:7NXTSRO�f��+~�>�B�H���$���Q##�k
�D(�{��f���I�Q�c!��c-�
z�2��s=���rO�AW	�Ŀ��g�CR��)ֈ�>g�����`Հ�Ƭ�+�H�d��W�47�dD
�5>ֈc��с�з�I=8T�%o����J���!�-i�[�����Z���=�sd�3V
RY��f�jFH��^^��:��5^46�W`Wn���#;p8'����{C:�ŕFT�?�u[|7�mWV/A�U�Mb�q�K�])�B���Y�P�YU�,���ޘ� P7|:�eZ;d�����]�T�B�W��
+ܟL� �F-��6�-'�o�rt��AAG2�f���5c�$�/��U���+j,���J�Na�Ě���<���k����m��7*���1*�&��J$d��/��#�{=���M^<�C�.�^�����s9)D?��m��jR�
�b�ci}r�#�t�\�S�0E������KF.�ےc��%�Gz���}�{��{=;P�A�JN0�1�{��[[��Ҏ'�T�T�Heü�˓E�B0J�ײv*OɳB��!"�nWBz��BgxJ��ʊ-	�g��!mMsro\��������N�!���z<�+6r����!�&R,=ڠ0-���K�J��?��IZ��k�2r��V°hLඖ$��56�}y�(7�D�V�0(٤���b6�A�\�F�[aP>�.��$�ɘ��|�%�6��
3uǶF9��W	��t����w�������Q�1��;
��;�,q��͝��L�lM�Sz�%�tZ�m�e�������Z[��Gn�|V{�U=�d�x���2������BG$�Svo|�1�Keg� ��T+��K�
�|�v��_��?��ڢ�iO��[����2�����L9Ӏ�~V26��S_�~V�h[5�!���H��16c�.f3@��r��&�+T�3�9�IkI� �qJ��Rѧ�0tS�y+ޟ����Pe��5���?�!6��	���	\ɛh>��8D�i�j�4���6&l6f5I��A��c\/)[�=[ve����vO���K�CL���-��ʲ6b��ۿ�T���^[����8\���6DS�����W9����0#��y���q���jk�|>���� ��O���L8%wQ�p�~'����t�9'��Y��dUG�	_[t���m/ܿ�N��n)8y��s��@�!���%+H�
��4��,<��T� �?	�c���=�w�KMؕ�մ�/7��ϕ�x�㛏U��]�1��\+n��VA��s%#����y�EJ�c*���yJX��$mD�U󥹚X5&ÿ4�<�C�VM�o(K��FaH3�;�������+O�,Fҹ�Z�~*��|1t���Z�׹E��D��$t-~�͘�3�>�{)����2�20��̀��[ԏ��X{[�m0��BZ��T?<
>[�W� %Ɛ͇R9�~�n8uu��u=�d�mOz�,};SD�=<��@������ocs�ʦ��q/�3UC��7̌�\��@����>���X���Z+/Q85���J��D�G�Y�Wx[�Ű�nJ�}|���<�շ~�{&�Z1�Ca4����ш�0҈�w���W�Z:���[w~埱<Q�x����c썭 ���p���������.�/�A$s�
�]�F��y���g֭�[�	%���Ys�T� j�����?�QXm-m��M�+�ȯ?	�7�������t�w�R��x��FeH�������xc��0���{�)����9yV�v�Z\>�ŐЁ<�Ɠ8-�a��)����{�%aW �X���hl�e�P+��|��9���=�D�?�c��·�D=�1u#�O����VH����p^�{��*��)�#{�Yb�eL-�{=����W#�G����Hc,�2��%Z��p&O&��:XQ:�yP�PHj[�!������h�^��gT;�AQ;��a��H��Z҃�i���Q��c�W1��h�RR�9��+?gb_��!�nI��\~�uam�5{��RyoJ���M=v���ɾF��	,��JD4j�[�YN��, D�T!o)=� ҅O�P/�M��h�Г����iz�%���^'.J����5��sEH~�N�or��X���Ky��=�,�*[�����J��<��縁8)���U�#�v�rduT��%���㖷�wo��H��X�v�Mkഩ���4b� �d.��שM}���8��/V������l�޲��/���/�ևxh�e�?V}v|��Q́�aS�[x��q�%�kO�䦸?�����(�?�_�"t�P6<�e�씚������Ȍ�` 4Q��Č���Z���G�P�ʁL<��'����"�����#
A���;��5������d��<@$]�:�ש#�5�U`]I���Ű�������4����o5��{[��.�?w�1/�~�܅�p(��K�#��S���AL�����Z�O�\�s��們fH��x UYHj�%F| Nh"kO��P����c�w-�s�n��v��m�E������y�s)Գ���M�S�ZJ�	:�,fW��8(�1È�g��]/�i{��%0�m:`*:��kD�*�)N��f�%�a�����B}]�B� ���V�hn�=L����Y�j��|P[@�b���9�c��T�i���z���^۰��m��l��fK��PQ�����dٖR�ڷ�mM��s�jM	g��g��w̏_�*�`>*C��C�ND�&v�[�62L�;{�q�1�z/���#���y��IN<Ķ��h�3"!��	�5��֩_�!�jwT9"�!�G�V!�*�T:��G�v0����oV���Y�R9&��$�'�>��E�fj����<p-*��g��[��+���9)��w:UD�͌��*�%ޮ��:ΧbH/Njwל�峲�]��ĄZ;jX��0���,�[��3L9`��.��k���<�8k)a�'��@�-F�qÑ�d��[�90��Dg7CH����Λw7fkR�&��*������zi'.����/O�~�=7��ǌ�8��uid��p���j2�-���]�fs�ݐ��J�x��Z���-��*���V�#�`y�7���V��=�%���R�l�ֽ�95�kNQQۀ��.fn��`�jV���59��%L�V6S�	�6�=E�ys��fz�����	�Zz�G"���XK��Ęסx�CJ�+hF��v��Ġ�[�f�3�ͻ�;���,A�Sb�M���BJ�^JI�;�q�#��l�)!�`��X��O��������5�.�	g<�%��`e������Nʃ3�'.����7��!���Ki��,��!6��@�GY;��r��-��'\�yp�$f*����6b,�[���]K;[�*�a��eɊ�~TfOC���OLS�_x�%�����I�W�<� 6y��s�ic�����mE�QW?x�a�$�+nz�c(� �3��/��$����s�x<(���z�7�ÍS��B7e^}-Y����a�y?PU���5�|��h�3�v��R�ul xˌ��4���l�e�QNzu��z�)�����j��V~�(uuouagw4\�T��ҹe�x��iD�labɹQ���}|h+3���v���s'�S����x\�n��������L�̑p��u
�O�ȼ�J��	%���	���CP1�.�?�EA[�bZ�מWa���u�By|@��j,����hd���ᾮ�>�*a<�K��l���9c��]ɧ����g_�6(ޘ�m��k�ɓ�6�?�p�p���)�=���Z�#mxy���+�SW�b��0|�Yn���gW���p��S���ٮ/5���6��a!�p.jnȃ|S��W�߳)՘@���u�TE�Q��ͤ�����bHÓ�ސ!Sh|���+���M��(�hdZ��]�ߪQs.����0�1؏d&���NkLR��Pޛ���Z���O�R`��S}L��hZi%R+2���D\ч�V#1����<M�˓6��&	"[�gF�g�pJ�˼��l��g��s�L}��cd}� 鱬�P+�A�f�C�-+�����!	5O�9[2�0�������j�+���ď�֖�ze6x�SQ^NJQ�'x�-V$�VЄ`_�Z�լ{?{cD�<od��T5-J�����E�+�1H������I[J3�6u,U�0@�r�HU�Y��3��b�Ʀ��C#
u	MF��K?l̑���f�%F�;���Wb<����Rh��k�7��$n���2����Xɫ��QRJNX��IC-.י��ƃA��Z=$������Y��LJ���Ǿ,\o���co��-1�]�9m,����-�v���H�J^���fFPՕ�¼��Io���o�JR�=u9,a�YN����w���n�Z����{�D�d�_uy"Ai圧��F�2�je�I�R�q\�r�����&l���1��u�Vi�s��0�O�a��Z6׼!���h�W�*��'�4���!����FU�oj���їB��ͅ���	A`��K~a�3R�P6Oy��UY�ۺm>���?Hhl��;�����x���d�Y�U'�xP��2*ԩڶ�1��w�A�%~YD [�ыW�h"[Y	��EkYi��}wy��*a}g�j�Z@O��f9+Jh�\8ĩ��{n��{#� ����T��:���C��,IY�������	L�U�
��L�Ł2NGY׮�[r�"��{�/��2���X)Ό|�a�A�\وǽ�!Z�܋9�r���qC��R��.�Z�ɃG��d����l������ܨ���-�}_�1�P�)K���
����!E)��n��U����p��[\�Q�� �[N��(Ƒ�e���cl��%���I����\���)Љ56V�N'�hT[�F�;sA��.jA�
�zʓ�,`���]=Pvu0�+�w��2p:H�	8��`ȗ�A/�`�y�jn�����KY�U�njl��x�z�
��n���Nb�W���/nEP�E����3h�vMo�^�D-�{8x�����!���t�OF��2ێF�!��#B�����в��݆�a�Vv�Uģ�Ud�{t޽F�.�s�ͤs�ۘ��"�ۺXC\F0K�F!�?��$��n�oES�Ác�<����j�TlT�K���C����DZE�-���g`%��[���7W���K[gf�#�Z5p��x&ws�����u��Mc �$�2A��M�����F�w���n�rS�DϒZ�����0�y���?�7a���O-�<�v1��_u=���������u5L��wLjddP�L�	�j���4���!�/��*~����/�E�Wk���񹃒;iH3��a�8���OZ���F������~�����X{�����z1��N���V�/����G��/o��)x�UW��yL���!\mb�"g����p@��d҅��Z��	>��n���\ә��u"Ｓ.Q���o�jW�T�!۳�S]ac��A�l}sJO����FBF1�~Y=��k�WC
�
k��Q��b��O�yl\�Am�ӗ��r���A���D	�(P�V^{-;�����5m�U�;�B� �u���ǅ��m�_Ƕ�k��'�����%=��H&PLX�	m��].K��Q�T�e�
�{Q�[&���U��s��,И�g^:[Ġl�1��cN���V����7�u�Uꖌ�P��@W"p�ҋ�F%:Q��T7p��Aj:��Hw�G|H�4
Ð��X�0���RZ��܌�z�3�y�Y��)>���#��CQ�훸�\��Lw 6�}��A�5���;��%B�I8�i�=u>�r�Ciɽܢ�G�tF��a�����m���|��ѐPJ��B�;�P)G�$������sG�����|N��?2RG�?�ߊGş��`+I�zў���VfW���A������6҉'m=�e�8"�r�)��a,i���~ҙ�x2�Sn��B�T����Z+�C�c6���n���4��������A�D޿p˲��0���Q�q��� ��=<����*���r��f�|?6����-�ؚ�Ҥ�e�����h2t�2*8 >8������X����P+k?�_���Ua�\�e�5zC��s�4��@����k�U�5�w��[+��tB�pL&��mwi@hM����|::��m�o:f�q��>pZ����ɛ-{6��h'�q+y����'����!������u%&�
��* �)�'Ӗ�`�E��n[��)$ת҂��~>��|�ѵ��>�.�AR2*|7�I��b-Ƴ\*2'�0
e!�^���j��o��;J�ޓpc�|O2��k�i�I���Ɔo�:�X�,�x�5f�HB!���6$f�&��0N�ʩ�b/u�9P���¬��L��`�������Wd��Z.�b u���	ȉ�)��vwM��H��A�,����ǁ�ʿ�!��9��y���<����C��1�L<�8w��`���0��6t�H!����ض���I�8�T�Y��C�	�-?:"�!���:0���+y�	rY���#~��a�!�{o�6�k�������:t�aԛ�7B�#y��0��*��� ի�=	+Ȱrb�O}1�&ߥ6Q�|��߭�79z��a�O{8�n%^�we�OzD)d�gik� �:8�[����7�{n�$�䡈z� I&# �8no�e��P�����}T5��[��PC4Пr-t%�������e� ��]��eN���������쿟O��!>ϝ�e���!��mˆl߽�{��xώu���5���������w���ǘ��A� ?[��2-p�ko8~8G�����ݱ$7��{Dfr�K��F��>����y���nI���B2��xa0�H�J�3!e����;0 ��}6���s#�g��If�A`JsSC2	D���o�W�8�?0G���������������#��:H�.����T�N�8)Y-��]i�y6����DL�ս����lύ�O=A�E�=�@��*��t	EzeD���VP��#��#���	�e��MKM0"s.�!� ���[V�={��	0�e-���T1�e�*�����k���T��$8F��Ze��ʫ�]��y�$3�]ɓ�I��M�X�K��K�3Ct,��;[%R$-���&Q�v����@��[ey�آ継�3�D����tx�ͼ���E1�Ϻ����o�i�oBg�"t%<��Z��M�`�3w#ބSdP���C�?��KR�.k����6�=�����(��O�<�r��^0���&�0�q���,�JB��6�Z�h�Z�^VK|f����*��X�q"Vb#�E��0�}��zX�2�.�5s(׏��$Bu�زY1�q��0�P�U�И���Y^E-K���󭊵/q>=o��c�oV�߸V���d�9D�3��,����P5�|��rtj�̾UJ*vuX�r!3%�b�}�L��l����T��A�E�����2�!~���eֵ��C���|��Ϧ{M�ϤK\���`�s՝S=�d����ƞ��y	٨5���Q_$�KI'��Q��f-�?h�0e�U����G[��U�{��<_��[�����?�g��4��]O�բ�ruE����ݖ���e)�6y�ZM���,)LR�����^AQ�N#U�f�XU2�W�4��;�IQ^*Ҟ�R�#��CR ��RΗ���Ÿ���<K̍��Zhn��be��4�!;-B*��|*}%"�&v�W�A�N��d�%>��\�q������O�^��V��������-
F�"dRF��d7Q��]L:�-�u�"���F�(�r�k�F��p"��T%�}�+���4����{�������S��;�w4��q4���US��,�eȹ	�R�rl�M�tk%.���Z*c�EȮ��<�3��5�hX*l=e�*Ӎ|9$��^ݎ9>X�LL%Z�.W�{(�@�a�ge�R�&u��!�XJukd����f>��.��
�O���&�����Gv�R�1fI�c���ׇ��%:�l�(�z���m�h�[wC��ZD�=������Dy܅��V�؞w쑜3D��@d����,�F��u1N�I���҆;؋�9?�V;eii�h�xo�eI�8d�J��"�2�L�+�����]�཭�-�:Z���sYE�Z3�{(8 ��0U�ԳL���|�ޒ;[�RWK/t�+ġ�n~�X_��*$T]�P����BU-�|��/#�ò'�P=��2�Q���j��#n��y�ʲ��K7��F*6*sc��%��B��v/���ܽ��<���_#�+Y�������WE��{�ZA5�h���C	X�]� �(�\���T⾠����6c�O�y+.��Ń��q���L/����i�X��%3�Sco��o�DV�W�����c��͑hWLV}I�=n��Ҹ��!�a�%����H�m���$7�n4�V����d��*�?�U���b��:��qR�֔�c��i��	��Z��ZG>� ](D�� ����8�U�p���	@���Kσ�wy�Ճ5�h�l3yY����y/�Z[��*����:�ׄjK���7P.z{4�Q��G2C���Zl����H��y��ǫa�]4�2|޴�J�nN��]bq�+
5��+�y~Hڪzy�e��g�)s��Z.�]¥�%b��z���m,[��7c�]J鬺ڸ�E���{8f�D�S�_O7}�b�lPT�c��ŎE��rO�ɺ ��D(g��Ʃ��B"�K�m��?Zt��A�ne���|ΡW#��F��D1\�����P|ٻ��R���M������J�ֿ��$�=��#/m��_+)U�E)d�Z���W�-��p�U.�� ]��>?�P������N@�7kx^6 `�2�ZPӸEL�ҍ2]6��4�3� �*��Eq��v_Ch(o�DpϾ5���9��銪�+�x��9	4U�eCo-�f���H+Р���%u*N�|.��	����9���ڕ5�֏��v.��~Y�Y|O� �3D��$�朝�[��&%t����T��בi*�HP����ޔ�]��"��oj�"����Kר��
�p�-V���O����Z�R͡���h�8g����iΡ�>F���b�Ҟ��2E_њ<�&�R�]�Wʮһ�$�e(��]S���h�D�9�j�Qkb��k���UO���x�2�آ���|u�7�$�J10t-k��MM�x��E���F��s��@��	���ƺ��wB��VV�qh���d=A�?o�g�*��Ik���dGPC/���!j�U�u���֘����"=�c�ɗkT�ӶU)�}��k���[�h�~��ʲm�^��Q�k�h��)%P8a����#7@���2^4�ə�k�Ak�\����2��ӵ����Jݚ���~RZ//�U��n}���aN%;gV_�]�a5WT~�2u��v �!�y�b��L%�
Z���-�J.�gm�s�E��U�dU4Cue�
F���狢k�|^���_����ĳt?�1�i�shM�zU�EE�g�}�b����М�D�e>�N4%��"�4"Ul H��Х���C~8c��$n�ҰҘ��H��4XBY�L�*��˸l��񔆽����k�$�w���I)fٖ�UԄ>Z�Ֆ������n����ַ�AP���z�!�����u&|�Z�,��MZ��OO�Ae*W���������v^�N�Xc� M�y�*�m=y��\�^�B^�gK�lE����������7�H�ˮ=�
�޴ٚZ&JF����U�Rs�U,99�Uiuz��HA\��,2{�]�D��7X��,��g)r�y^��q�^����؋�A+�N2y���u��+�OV��X2�4�b��_dP+J,�2�Gu�ɲ�-����רwݯք<��dJEl��(�f�=ǹK68�&Os�|��zn�<q�zN�2��H�e�� X^e��$��Mx��>OR���,[��e�*� NT+h��'򊂰C�%Kd��l䃪�hy�:��.~��m�
��׋�M��ed���FGuS����Vo��[n	�$%:�,Ua}j�_}�9+Q��5GA�)
��F)й��2�>��(6%��K�a�Yv$�3dU_ם���D3��Z���d���"��N���_޻X�ӥ��~���KgG3��6�<��F��R�Ȧ�Q�*��F��Nz&^�VW���_�hYkFH��0!��;���ͽo�M-e܌R�Lq�ԫs\N�{��\��^�x�)_�`v_W�KI�����^̓��ǋ�}��J�ni�"�W�����ō�U���Hx
�7�)����h�j�^3�}���1�����~z���k��ŭ�F%�f3?��YP}gG���﷔���_6ISj��%�%��EFe��u�=8�M;�T�<��w�ie� qn_ ������kb�m�1�]�ޣVjqȍ��yTM�My�B�1�K����V��~�z�R��t}C��P�j=U�J�(����ͽ\�W�/�!�4d*��#JW���e�
$�2�K����z��ac��fy92z�L���U#A�:��G��k-�q��?k���4�������ȉֵ����FS�������.-���I7d�cp��Ja�X^�������R�U��}�x�%�YZq��ma1�0��/I�I7��|~{�t�+���x�j+���AB~מ@xEq���sҷ���NOw0�z^1׎{ma��u�U^^��ҥ�ʽ�Q�#�Š���_W�yi�QK$��ߠ�Q���ҽ祐Li �2FGɥZjۄ������[��eL�Ja�w�9x�=�ߋ�2�/:Y^��W��}ͱ] &y��׫�K��7?_S@5�?,�yލH����{���q�˺
����y������cq�;�MۋUr��oJ|1UU��q�H+�7�n�	(>��=�$F=��ܻ4m�xM&2��6e�eN�(Ѯ\2�Q���+���@�Y�F�u�l�c��
��C�Pq���~gޚ�+گ�ՖP�*�K�$#ueP7ϵE��t��#z�N�r�pRn��j��-ׯ�|�i�N��iI�q�DC���,��(��j
Wu��gmk��OJ��t�K_��
|�o��17ܺ��O�?U��ԕ�ac�c����JW[��hʆ�ى-���{���gv;3��ɋ+��d�Ĩ���t)=��y#��/�����d��4�NyZ��w��������l�~�W�V�*6���c����xy��:�.��MG��c�"��������|�DC��� �nĽl�(8��K��H��i��
q���D��B������eLk�ZrNe47���S���V<�3iu��p�[�v؜�P�i�\y/)�9�Tf�-����1���[t�ɷ���鳾��<-B�C��cJ����H����J}�	a"b3Wc=pcn�����N�5��y�Ϸ�^<��]�U)\�b��� ��I��7���l4$�L��eZ|���lF+鲼x���ӓ�Y�E�ͤ�0'��qU�/c��ZkL�3]iI@Eh�"Һ��@H��kG���G��e��*U�w�u|�D����Mn\�Q��u����CvX����F��[�]�Z����7eu��|���{j�G��{p�0K���ϒ��Y�"�%%�7�Z�*䋹I�L��m�޺��$6��e!���9�=�>B�[R�$O2��������_
w���_!@G����8�NK��6덲īQ���V��3ͭ�Y�Xk����m����0gX"VDx-[S,á���V�=~��/�%�4�~����"�0����2��y��V�pe�hD����gS"ͺ��x���j߅7�{�> K���W���Ÿ��|&i��Zk����X�kh��r�
����BX[Sg��1�����6)t�t�U�ǧ���� a^R���Z,�n�����g�1�c_3 �J�8\�J�͞�o�S��YQM�1ֺ�z,q�ih5���D4�O�K��l���^�I��ۍ�ܳ�lpe�~u}^��)�K�s����)m���~�jk[�������"���ꦾ;	T��E��>��ؑ��wfۓ�YL�:��egh�^5�)^�R��F����)����*�M׫kP�`�ѫ�)�S��=�{%})y�T�l��#� &����g
���żS��޷��໗�~YJq��d`	���>��L*�2�o&��������R����Шȸ`e��o:��29�Ks��� ѥ�jv7�|ټѯ	op�b�]XiԆy�\7����&m�9�$x�}�rz�q�f~�����b�`;�x��),ukŵ"��F���h�ёP�!c��n����P*K!����fl���;ۚ�^)L)�n o��M�ι����4S����H����֍F0�t��w_�!ϋ̡2�y��-�:����N�d�#iY�9�^1$6ڸdb��M�W��՚��l���3Ou���}�|����Q�\�g��L��E��Jt��hc$r�ܮx�&�;�(s��0�����XW��\�a	���=�#TGh��jP�=����k�ҥ�oelrx��Ht�Hc�y���.����Wz�6�Y�mLV��8
ٜ�,($��f8S��"j��7������fzĝR�jw��Ԟ�-�Ԣ�j]���p�iY\+� �R�U�$��n����4�����Y"�l[ht��� W�۰GVݲzSRk������
a��Om�!R��?��Ӝ=?'�cK��J6�e�]�Z1�QRY]���H�������67�f{M^Vc�[���!������(�4��)Hc�
�Kk�ϩJ-(A����>iE�5F�\/��˒������g*_�^�Ȱ��EN%�,�����;� 2�w�S`��}y;s�-�6�7�΄N�����󳿑l�Gj1��r�ʒ��ut]�I�<�l��Պ$Z�퍡�bc��EHx���M�e��v�ï]t�����y+��:v��u�n�/g�pB������E�{a�g,i�=�7�Xk�s��I��A��u��ى��,��s���^%_R���spZ$4��X�� �d�X��Ms����ׅ��bT��k(���l�]{�l\7������$<�RW'�M!�%��[ěƀ�VB>C۸��>�R[<����4��\J��4"�"A�^8���X�^�)o_���`q��>�K��m��]`�|� ]nj��zl�zA�0�hf"e;y�� ��r�1�����ID��i]�u�U�5����s��Kl�V/4G�/�vM�����y�CC�SQu�+]�<F.x�@�o_���A٘��%�1�� L�w6�5D�z:wݒ�s���"e��e����NA^w�c=M[���2v���Tq��s����s
��]�f*��5�4{6�3�l�������x����"�d3��^Ќ[뗈�_ULR[��s&zL%�0��{ܠ�������Jt��;��OW��<�qɹ�^2��&������,��r����M��Ұ�{S_[Wzj�3������z{(^�Hw Q���b�X6/�����kkmn��8�K��X�Vf�r�b�� �M�7]��j���a����0������o��{����9ц�,{�.�@Ԗu�-6AC��
�U��qI�ƆAHt�.�<G�0[Z��+��5n�����{;s��	�!J�RP�xG�X����"�}���F�Y^Ύ�;Qْ
���rWEZ�iU����oY��'u��!B��N��Kkr:(�\��K҃i�B�W!�r^���pO�*�HS���bo�a��ѧ�H4/����+(՝sܫ�.J��yM_ob�.Qcx@c X뭻l������t5�m�'ä9y�ş�,�ٔ	P�*�S!�M8�����cL_�����<�<˖�t��M��r�IY�Ɖd>��M�kd^�B<�������**ݪ}ICA�U�.۟��Y��j��B(I��H@of�U���3{�m�̅��Ѽ����=3�*��r�t�òE�2/Ky�pGˀ� cRx��p<�'�P�c�H6�pnK�����oj�]��sf�s6����o[J�Lu�8�K�I^�+?|=���B֢�S���8�.0�"��kڛ*>�6�x�z�[]\a��µ�0)c�q��=��ܦ�fQ�b1H��8���!��K��$Y�򨞓<�h��s;kz*X��fhua���|����a����z hݍ:Q)�ch�x���"���'�'e-��1���1Y��*{R��#S�6�ە���\jL�ݥl�|����U�_�Zu��dMԲ�
�(�M����a�l=�C���%��z���{�LI�SG�=2SYR(Hۖai���._]�9ؕ��/��'@|�t-JQyZ�i�����H�9%̒P�����b��BƜLD�.��Z�Ǭp&�~xbWsrl�.��#z�}���q��mtť��"�+��1����E����m�\K�䐂��v�&�j�vyHbp��o�Cʑ	$m��"�j�(��P����.�6nC(=?K��+�*�dˠb�\`[/ ��5����aРuʡ/p+j(ni�ۓq�$P[�,�k�}	ۢ����$σ�m��v����x.����l�]��`����\xs���ʐ���� ��ǹ43e���%�&nm�����@H�[�F��>�j,l����%�Y���=ۙaG��s��lɧH�IN�vE�Xc����w����Λ���"��䝊F�~�0?�.V��_���w�nh���Ҋ"uڊa�Y
&����s���ΡdC�.B�� b�R��DϧS[l3,�v�����}����y�ʥ��ue٩]9C;�d<r����TZ�i��M��r0*�3n<�y��y���f�b����\X�x/l�q��ST��,R:�[�7@�n��;�R�z-�Y5-6H����!B�F���q��2��J,K��F!��p]��u!��"<�t��,�'?w�j�����	��ZE �)���E�=Y������MTN�	p�M!��\W��LzGQ�z�k+ `�"=��t�4���ihh��fw,!Q���b���)r�{Dz x*�[�hhy1����Ev�꞉'�\�s�k�ze��`R�G���{F��{Yd�=&�U�#V1� ���mR$�,�n�H���c�*"U�G"ѪL[KD�!���i�̨�\Qָ��ue�J{���T�n����%��n�xX�m���m��j{��P��0#?/�ҍ�}`!"p����K5W8c.H�R�g
��v�s���=���I�-=��O�B�RM~R_t��ќ+�u,��ļ\��Ukq4��ثMtu�:���H)"40
���I����L�3�A����!�C�yD�~���;G2K�?��ۏ��F�*��r9["�rvis|��g�-;3�� I475�'�����LK6�г]s,76i�Z{6���/�U!�  ��t�es�?u/

㾟��X� 4_�3;t"R�06J��b��@�mٔO+� �75�s����)T�!�s�1�x��5Kl��RH��f��R�p�І�5�ܓ��� H�����r4g�	f��8�X'"=�썮ȹ/C^	�^U�5�I&e͖�ߴ��ٺ�[2�U+����Q��=�v+t�V_�9Jњ��s@��TA��n@s{_2��=1kw>Q������n�M��^B�7\C���;C�qi")tL��{���+n���J�����θ�}���e�_W�&w��V�;��LYs�Lp�2Ae�9�ݍ�WI ȯ����]c��'�P�OɆ�\B6ۢ��F�����@�C"Cs�BZ�t�S�1�-�]�'���uDS��8FC�Uxm2�d꿇@�t�x�i��1�����74�i|:�:.Mͷ�^��o˘��|n���p�\&w�^�]5���'��s����L�#��v�=A�h�j����њ�5��K��(���3�L1n0��+c�s�P��Aw�_ho)���sE������V>�,���vI�r����K�:�SO����5���o%l��*�(U)�.���0�+NSV�^U���y>[SC�1J��~W!�s�B�F6�X|�����5š�}\��GB���:�� ����Ն����� �����D�}.	J���B���k�+��ɓ��rщ�%�&�m*̃9b��w���~�,d9��M�c|���G�z��x���存[�a�J���$w!͐C�2f�<�!��R�mn�I[c@o�&�M=��j�MM���!�#y����P�JU\��̙��3_.��%�-jޒk�(�0����Los䘎Cd�w��V�2�)��:���e���3Tp�5��=����etw�o �e�(�����������N[�]_�4P��*�\��	��	���HԳĢ������H)�✂j�V^:<;-����v��Xh�Ui�����}��l�3k"�mK��?��T�)�e�UA���c#t�h�T�/*y6͞S�� ���Ꝝ/�0MFky���759�ͅhLɅ�c���:n�xKE���{�AT�XmT�h������ln%����{����$eLJ��X&�ڹ��ؼ����]��^Y�.���إ���J�6�)r�5rG�z���~]�9��m=B��{�k'�z�s���Aw�f���,)Rq��{Y��R�dF���dR�A�v!xR覕��tĵw�����^Jh�_h��ο����p�fA^[ܺP���W���96��
�z����ѝ�𪫵�\�^��,W,T3B�(�N��%�P�Ew��{\x��,�W�IlK �8��|���:])�XǷ\��=n�j.����x��eN�Q G�w��@z=����=d�z��'󱇂�z4���T�R<)�.)��=�1�Ƕ��O�cp�c����;"u��a]۞���o�D���8T�$�8�kH�5�i��k�`�c��Y���%qj�FQ��}�����~���yW���άCTy���Y�L�#��z���	���m�"ou�$G�P����<l���y�'_(RCI���I����dx	�*�W�^/�bE<WV*�qY���S�{�JCq���=����)Ф�k�Du������Nܧ�H��f��^��8.�3�?f#�ڹ�|��|�	0��̩������1��߫F�n�g��F��Q9��D}�Is��fL�c��=�z�%ⷘ���
�!JR]�@����ҫ�F�qm����1b��D71]qO�V��l�j����Wg���d���#K�4�c�m�5&Z+���>,t!i�¬qBmK�x|��1����Y��%�ϫ�4��ɝ�z�5S�m����bgr^�)��N�*���^a]���佗�<�s�����D�%<�<�<�r>>��=Q�!��Uq��xA��y���}��W�z0֌<�3~5FJ��owww����~B;C���pյ�k�H�V�Hu�k�B/%�E]��D�r��K(�����Ӫ�P�6; ��u�4�G�Zn� �B7������z��ƌ_ή �Hp]+@C��3��qQ+�+�(C#�����(��l�Ce�{U6C&�,�]hZ�=9��9ϜS���l��'^�{��D�`��v%���W���}� SҐ�M_�ێX��C'4t�I�1�5x�K��t��e8K��23���*����}�?��U�q-�.+�(E>���tU1؃����&��׬��q]��=��5u��&�>[����ZY�o&]��3�g�qoX�݌a\Na��.T��F�绹��kd�y�Ǔ)Q\w�}��]T�܀�U�{���51���q/�rQhs�Ǩ����TcU��Eϔ����z���o߆"��/�Hщ������H�G(ͻ�T�0�T��נ�&MV���-��B�븄�!Re�*�
��$��ה͝U�}�m�Ly &y�T�(f�l&%;����j���x��*O���̮�[͂.>aBE�kیA��8��=I���n��a�!j���׬�(U��4L�Ŧ;Me�8Ű���܎����O1�.w�\��N��Ѕ)����[,Ȍ#v3^�w��(/�aɰ�-a2���>P�ސ��Hz�m�T�ol^�lw.JJ���)U_����o�Q���t�p�%�Ft7$��F�jO�c��5>�쨡�}���o�r9� �(ZKMdF��*lE���/���W����"��^1_x���%;���T6%Sj�@����P)A��H.OPn�&�lc�� ϧMx����� �S����y�1Q�1����eW�:��4�W1�+!ү��zU��HG������*�|�T��2��|�po����Ѭ��l�]��N
�:ȭ���n�H$HJ�)�pY�G©ʇD;YŲx����`� 9��F�;�Y� !T��0a�վ���/����s���Q	W�ǹJ���`|�1�6��
�O	�B9��kݳZ��ω+ڝcۘ5�"�;;:�v=�x��ۛt�"���K7�簄�-o���XkQI�n��ڦ���B |����K�&�nE������?P��B��0$�O�͓��������=@í}
�|~�qu��gO��I@����C������O.����)� Kz:�R�Z1"�\5��nW��V��דL�qo��^�tVR)� Ej4,$#��=�k	c�5��óL�?]~�+Ƈ�^��Fp(6Q�4F���Ӣ��``�n����Ye�dp��㊌��G��T����(N'�B���kD���2:�����Si5��Mr�l��7%h�GE�%�v�(krJG�.n)�(�j�04b���qL���x��PY:���j��'޷��m.D�V�E�`^��r�k��f\���$Q���y(�>���:�#���M����%��j�+������Lj$J����竲#@tg�)D���M���S|6��R]����@a[
�CYt�!��~?G�M
R���aۖP�����Ɛ�]Q4cx�r���Ux_��b���	��S!���?������(����qdX�Lxx������C�^�*�+��/h?�}�|�w|����c%��/��@a�}[�odX�2i�}�+�j-�P�����q(�B B�|�A}
G�pWZe�V�L���c� %���ֽf<+���3�5��s���@�J^�<ͱM����?�����+��9�]ʺ{�޺+`1��Uf|7i�т@u#��d�>����p��!�`8��Z�K�`S��9��1Ez���u����Y֧u@�J�������u�OP��V���sK!�>o�6�@����v8h1��~p~�Nm[��i��{G�TV$�Y��T��s��M	_D��6�o�D��<)�F�;�:�9�R�����Z�����:�X�xAyZՐ��&a�qѲ'O�&G<��MO����;��W=vd����,���0k���`��h� <�C��+D_��}�k��3(Fk��"g؋e�T�DA�H|4?��W�,E�p��a���fl�������O�!\o<;�H
�
�������d�C�2\w��$�}Ng_�K̞�KYO/=��v��-ۍ�%�o-�|�3�٠κ��&�U ]�H���T�^oV.�����w�T�Z{'���э��u�`H������(�!�)��JK��!�#
��U.XZ�}�D���lbpbL��ͧ��
��YdW/h3,�M�����m��,�fc�m����f�Bg�f�֑�hV<Ks��8�g "�*����2�ٝ�@!���}_?�/�g�ޞ=���Z��N��\_�K�i�3K��su��nf���I���*�(���>~����8�K'
�.��~K�yrJ(H�E\��ӎ��ŸK7R�GgF�O1�H��M��n�uE,�%���C.����>/`x�(ҡd��kk�5B�"�k,�a�ǻ0�;SJ�Xxl�������Xo�O�S?G�ʞ���p���9���aP��H��7�<��-F���
���9v�7�QB%��֩9�Ԃ�4#��IB��I{ck�ϐƧ��l�c��d���2����o�1Y2����<"Ż�ץ��Ɗ�b&�Vy� 7�;��mK��P��֤-��Q��ʳ#����l7S���~$�"8�EKcq�7o͊���/�Ç�� �! L���ú���u �ie����-f�>.N8.� �	eZ���72��8�ֳ5O��CQɝ�畕U�a*YF\삟g��,m�B�7���C�mm��P�_�8��*N�%>�]Y�u�M�>w���ڻ�6��8���Ap�3�������H<��Gs��Ї�7eb@�C���z2�~�����qëJ���m5ȎE�2�Lp�r�^z��/Śm����ؒ�'W�N�ꕃ8�������z>����yK7�d��̦˃!
$�0d��1���OxU5���dU.���`�����������N��a�k������c�/�fgc���b�8� %@��}��ݭ��$O�a��B��/	�L���0�x�W E���>⭶V�g��A�`�ݛ�!����G�� �9����h�����
��� e$�2]bB7�c��!d�E��\�K(RQ+4xh@������&��Ӌ-@e��^E�������;���������O?��aU�o�e���⋙�/W��>z&�q2�"����׊
�:��4�B��g+��ȑ*��PR������z|�R��(�`A�Į��U�U���x�/�VxV�Ʃ�%�"�٭�[����	��(Ct{�r	�3�(�#�Z�0`.1�_}�U(Q"���z���.����)�sO�����ɲ�9f��yȤژ�NX���=�JXA1z�nq��+�j�?;��U���ܖbZ1�Ȓ�*�]��ݻw�8ܵ�����==�s0��oq�+�����u��B�����۷�L�`�t@�1�R��)y�2���䝡�J��.(�O�?۽���9`}f��0oQa8��*�;�0�b���gH�����c��axA�W�Ŵ�aݽ����->��a� �Hq�Cҝ �"���m��5�>����_���҉q��1?��<$�ب�N[
��R�z��@ִ)��+Þ�0T�	<&�eL7�����Í�����}�bj��"iqCh!X�����}�ȸ��?��~���U����:�m��Y�T���?��zC�#�	����}�����r��ŬiA�������f��ȖYu�٠�!�N��`��ΐ����u��ݝŸX�ؑ�\I� p�0,���(�����X�oL�qNSP��N1��ި�()��1@�7���7��u������Psko޾1񹽿I��hڊU��@�٨M%���� �wͶ�н)>j-�J��>����גަ��uL�"F\�iUr�;��#���R��`,a�/��~�~0y�}��dTن��V%�*b&�pN(�Z�Fo�{��a]g��=RZ�9q����?������w�f�>����O��fw����\� b��,�
�3�B�\���<=��)f�;���B��sךԪ]d�eH�H������C"��B6�|tgi\�Ǉ��K�p�<����� E�gȀ��q˴�}�"w��T��_*�Ɠ#>=�-��%�+�آ��1& (D��~����cRޯH ��& �t,��@�*`���5�B�z3�+
������kQ_Y%�d�\z��ص.�㰉äU=D#c�?�*�A���4���.��!㞮�`��-�.XkYE��ňq2tW�M*�P�&fWVo^����U�~5��sB��\�)�Y�	�\-CӗP(X���/#��
(��=V�!�`c"�ǖjO>_��~Θ鲄��Y�Z==>��y
�����BNl�q�}�,t�h;�9!o?���B�����*@q@[�y�e&;�qQ(c���c��V@����_���8�5���e���ƓR���JJp�Q��Z��}(XR劜	>�d}ǳ?����w �{Ý/b�Q�F�� ��1'��ޮ����2T2�8�J���u2�S�Y���$Ӣ�;��c_"��&ܕ��_���+����"�[)R�0�䉩�\ɬ���b!�_~��·�;����_�$�3h��h�,Ѓ��:���^�����tr������O�����D�Τ|Q�N��Hҟ��)K�!��{��e���\���L�nDD��@]�p>XnX��*#:y�c((.�Y��`���U�]q+{�C#��+:��v?�����f��/��b����=��Y2k��^@xP���Y��"D��)b�ճxa���S�	M��Uqb3	V�A6��ע�=vW�B�{��������x�XJLW�6@COD�0^S0f{6�H�ҭ���dn��H�����^^:����$�Z��E^d��ԕ4$*{܋2�_���3��p �Sb��IԻ"�=e�����/�����㺗�\�lМ�%�)�Q9S�0����'e��(;U!,� �CZ7f ��*(}�-&+�x�i:o�Z2V��-M+Y&u���4,��Ev��FN�'-�V5��H�>;�>���oG%�P�ל�>�B9�_���0��Z\jU�O+�� �e���Dd�po�(L�ϨD:y���*P��x/��a�(����Ǘ��?!���!N"�[��f@_��]i���bx��ɔ���NP>.�'�.�D���l͓v����VK��X�h9BpS1F�ɡA0b�pOE��k9"4�s?8�i�1�\���}�[��5~⚘�_?��I�3㭗S�$j��ӟ�������2Er��UiT&�x�������:�ό/����qFk�$�EF�rV|�P�}^���7_[�U+J�a,q~��-~?M.sR��-VO�x��w����b������c�]�ڳA��2���ra��`��E~�uv}�A͈�;���[����x���ft��޽�sclqN��Q��'w�l���ΏO����0��bxG2>�(n�0ח_2��@%��ט7��Ֆ�%	*���R��֝3L������4�8���P��e���[-DԲ��t��
��㺴S��f�'��&GJUu����K�,.�ɂ����O�?�Ы�$�2�l�ᦉ/)�عP��s�H�͒3�-���N��U��i�ЛE$IX|��T>,i�!�0/,��.�=\��YH�>;�D4���r�ĉ$��K�O�z�}(1���d¤$����|q�'^#���{�gWlcS)#P'��-�@�X��o�ǧ���̅"Z��[^	k�v_Gk��p�$mjQS����������q�~?�_�r>�5���J�$s.���q��:���nYcs�QJg�b�����mF�1g��4R�GM�Ϙ��Fơ`�[��a��bA�2�<Df�	pL�L�&�wβ����=V�?D�&�R�Ԣ�nF�����P�%E�g���Z�����K��8�;c�-in�ښ�t�
�\!nz���� ���(�B�Cܧ�қjʍn�W?K!����o���o�ұ�p�����y6�X�z�ÇP8�Bt=n�}+;E�熙^�Z���9�l�19۹p�Ϫ��0����7���_�/�6�z涮��	4ג�X�rQ��W0��U�}�d�6�e��㧾��n��@���/���EĹT�1zW"�_�ɛ��� ����E�R�_�J�/&�ޘ�5OǷ��zk"�����)N%���U�S)|t'�����a\��B�??�4?N����a}�>�}"�� �D����,s}�.5b�G�ĵ,��x�]��-t4�w���++�U�CC@�?�����&Vٱ"3�'�!|VqE+-������(����!}�?x!���d��X>�<���@�h�U>���y��J$}����L���ɾ�q?�ThG�n�M�2ݬ�QZ6}&�E^����u�$އƩ�I7�d���N�¸4/!d��h����&b,l}������E�].5~V���&�6&�+�T֚��v+����s[|n�W�b��TRQ��57�¿q��R`�k��!�'���<0㈸��$�){��!�$f/��� ����AA�-���ظ�Ȟkﮈ)R�p/�qYk��=,c�5�G���%�0w������?��?V�D+[��,r��']F`[����;�t���&� a	e!�Y��q�[|4��Dɖ=8�_Q50R�~���=���Od5|��l_�n>�A�ӳ+u�ÆDuw��`0VV��9�8[�u�����z����c�{"�m{�Nɘl�Ȯe��1����@ō���F'2��Po�CR$)UY'�ϡP�%㼃�JHE�V�^�)J�UNL�|狖�U�^��!I�ǋqM���\���1"�#�?���a��g����M[޸�PHt�W�@�̙�Fw���Ժ����
�����(��¨W���J�J���l�R�{r	庶W����БYt���JU���z�v������(�m��Z��BTQ�X?OCS̧�#�f�{/%�b=�<`�pb���&��!+q<d ^�-e�H��4^�/��dUѝ�%�P1�������4
����;xv����qa(��S���p���Ѹ� ����/vN�O�A�B�H~�b���Ѕ���;RCF�w�F������PƔ��)�8�=�K4O.� ��RoW��X(�����n���7\w�Kܻ�ʍ�o�>b�1�k�BZ���]�4�;�A� n6?<��~��_}n���sɤ3��?�����;G�^=�F��crO� ˅n���GK��E}0�D/������|ë�X�1��s��x|^߿u����.�1K(D<��t�iwWy�Rj"�l�W����]����gCų�8��í#��� ����x�i�<_���*�*���_�2�����ӯT��|�Z����{[����I�W����z:U)r߸��6��o�=�y@�5BrB�f��� ֊�h�~d��Wq�8�z������K�����^��'i��� �L7ۚo�����A��h�H�sܜ2�p��#ӣH���/�;���5����u�.�E,<罻�8�n.H�ѳ����ӝ�K`(,���!�q�/�Z@%��|������X5�OO>��%�K�4ј�9�#֌�f�b6Z���p�T�\t��;�v��@�
��.��<�J����I���Qߠ#���b`���Z,�m�'Ɗ�E
c(�L�?�6�￰��0Ηܱ����5�ŀ�;�;��<�G�ޟ�Cx5�^b� s�q)�:}7R<�(F�ųܘK�9�����-d�l,[��0:�R��Ce�����O&�޷&˻�bޛ�	o
��=�հ%�3׷��)���UER��5�u�M���=��k�i�2Z�P����µ�aD1366Jo�k�g���P�t��\܇���R5k_u[(ّF#��Ͷ�^�������׌U[��+�7���XE�Y�Le(�8[����[۰Յ{{��
�	��n�ܯ��u��h�CZ~|F.&GM(�U��;/����b�X<AYq�kX�����?9O�C�)N��d��a,���3����,���ǟ��M�-�r����o8f�`q>a<�����L|p��vz(R�8�Tԗ)b����|�8����}祧�JX�tq��������w.�%�<>�4U�]� =�1�
k@f�[x�x_.w�0bE��yX��\��q�#|D~{($ݷ5M�g-�h��k��`���.�'w�ob�����#	�d1�=r�d��b��TǑ(h �Ǩg!�M$��2Wfh�N.�S�|��Iw6�"��qB<�Ь.e�ay3j�S]W��ɥE�X��m5_p�P�d@�t��#�W����.0���9n�W��BJdg�^��ւn՛�fX��ǿ�����3\����78�����]7^��h�=g�䩹��0�${�`KT�s퉨��l�6fBp��q�~�7���-�ƞ�B��g6�I4>�7������ x��g>쐈t5��.��z�J�� N���Q����$Q������ZRN�!z@��om�￶���ovO�|�M��߶/��2j���^X����F�R'%� <�0����-h��f����H´�n�8��{���)Qܳ�9]*U���CW��O?�+��=�iݭ�:,�/V"()k�] �A<�{w�(�ÝO*�B��b���r����Q����φ�n{�c�M&9.2l/<�[���yrw���S�N��u�q�莻S{�?9.�Oœ�G��'ƣ��\#ɉD����M�W������sd�3�Z�S�_��o��e�"����T�j��ܑ��F����8�4�zw��Fz�ɴq��':O�}�0�^֌y�(�)ۄT4�$ܹ��&Ej���J}�q}�R�����mA��� O'�K�AW�Gj�����|���"-٤���-S���+Z��Tk�a�ٶ n<l��N���#�-l�*�C��	 Z�F���P�Bj��)���8��7��3n��Eh�5lv�Q���M@��j��cq��Y	T�xR����.�:�Db����>3��v9��7`Q��,��r�������z0d&/沙�u��๕>���˷7�����Dm��deеg��ήO��4#/N�qҹ��aάф�8����l�c������'��2cG����2w0d�}#�|WE��?Ի�;*�Q�_�,2&��s�)�y�|�Pu��D�/xc��0�}G-N��&&� ;���"o�vc��G�X�'� �6�B"@@ٳ��nrS���W	Y�}�FB��B	�]�K�j�U���L O�������;���ͳ�6� q��*A�6��x啌Lm�r�<u<�RURsm����I�I+�擇�����H7�'����3��J`Z�%MN��1 ��{� "�n�*D$���I�V���������d�ѫ_p?IE��frHI�WuI��)w+ȘX
��3�����YՅ����n�:v@�����i
��w�sq�\4 P��L���u��ۼ���S�p�����1n�S�쁬��W%(�V�8N��aR�[裓�w{�b�'���t��T0�\Gۣʹ��-��j!���ͳ�֚�%��?������O?�x��\ͺ�xp]�U�=*qZ����%l1�[�>�ʠ�!���ҍ<d��<8'��x����U���a*Ҩ�h\����aI�dN.kU�2DH�⹕������-�g9�6�S���L�>��ZW��W��{�� ��17�ߋ���%/R�L�ђ�5���*o�yBV��Œ8�|=��γ����"��Wyj�ㅱ�a�=��S
��!C�,�?a���u�����5�4������g������&Nq���أ5����}Z�#Ăb36׊!��-w�dFRM�] }��C�$��M����U����4��v���^	�0h˒ƶ|��A�R�j�JU'Y��gO>d�]���4��N,�V�1#Q���Y�g|H��X��a�3���?������	b���|3w��ث�njj��K���4�ME�Ɔ��Ο�1�;e޽���cg�R�����K��뼖$Y�Ż��_��T#o(0>zl�}�]`����@lϬd����ў�|~::0IԠ��N�y��%9	�����z�=o,��t{��^����2�09��w��2]X~VJ����;{숌��'�5妑��T���:5�b{V_m7�����(�g�;*4UF�����M����8�}�`ct�a!R)]�c��a�����`�P�ry{���QT�E4��'B�0��Rk��cc-������?Y�<��zz��T�+�z(dﵲ%��=��4���������ɃЁH/9a�X����(9�w�&,p�q��0| pVYuv!JƮ�ޭ:(W�7�������ˋň{#!y���5G�S<+���gM��i�*	���ؓu�Iޞ,���C���{���Ǫ����5��gvɹ��l�i+l�H�w�kp�����j���m\��%{����)�⻉^"֊��D<m�(�%����ԃU-���&җ��ϐ�{�x���H�v�
�#)D\|0~�7���?�bW9*��_}eJ]����#x� ��$�->��-�&����(HGn ����m,������|cq�/�� i_Cd���k��3�qk�Y�Cdtq����#�"Z�!�er�L��yt���ݳo�A~um�&D������-5���gӴXǸg�2vIER�d�|2�Q#n�>�"U�}��?��"��8�O��",�)��m�Ⰻ����?c��+��"��������1;�yM��"��q`�KR[�'<RG��[AsYz��j~7�(��J���ܵaZ& v�s衆��Y��W9��ذ���a�����vAL�߾��<Z�f���m8�Ư��s�.�/^��^h�;?jk�1�x
����'�1p���;�֒]�G��8��1�jP58��j�������
���H��t��i��m|Zw��q�j�k�](s2�[� �J(������5�}R�D�!GQ��T���N[hfU�@�
����s�S���DCOA�"+� ȇ���s�}��,�����Vu���]��Ũ����K�I&d���}(`�-n��l�U�L���~�bƌٗT-�Ы���ØՂ
��QUD7��>E������<�\�"c�bO�2���F��Ѝ{b�O<�m�Ε������s\_� �E
IK�h������R�ݷ�{�~lbOZ��=���{���s�RhT%���.���K�|��E�������X��
�Nd�2���-�z|�"�B7�?o_�Ba�)�j�W(N�����Nŧ�E�+R�]�����_عH������+L�8 .�sxVeNVH� �9�hIIT@�5)s��Ʌ"���{�P�+�vp5���jy�ث>=>:!�%�f�NL�(�����ʀ4�[�����؆xOTH^ Q-��'G����w�/Z��H\$WS�����He��VE
��T�yTB}r%�geOT��=���"�g����zlA�m5���bq��g�?������HَRк���5�d���66�BIȷ���Ǫ���L�X��i*L��o���O9'R���]po���̿5����s&r������T��<\��L�O쎛��fU69�f�c��*�OM{!�+Jz�'��h�^��[M�.S(:��Crn��5h|Kq���t{씱��#�T�W�JC/�����Cª��	�-p&��~~t�p�&�'�"ǝ*:Xc�N��j�V/�G
�����s�b>XsƇX�C�K(;�C��h�����sW����t�Ϧ���	h"�^��ݞ���!/ >����`qP�����wW�(q�l~¹ =��	���߿��ד�]�e}�~�w�}�!�7�cB��	��Ǭ)���Q�σNN�����wZ�e��^K(�RA ��!]k=�������������g����P�k�7ǵU1d{�Y�"�C��A5�wN�BÂe/�m(F�(�ڄ� t��� &�D7��ʤ��˄�y�Pj� ]
�V6�`Ƶ����A��?����?�Lַ
6C��m�E�S(,�{8I��M(�~\��o�Ka�JV���"�``��7� �H�׃��5��ό�����4pڠS'�9��  �vN�ސl�n���]���{���hz���)
)6G���D�2յ�A�W��Fl�#�='��Y�F�\���KK�jY��iN�ڻ�����Ҵq	J�-��@{.��=�Xoqͳ[E}E�Z�E�]i�g�E`=�����B(�R`P+ƭ���'������V�)�e�C�j*��1�5�HX¹��˟-�޽p��._������S gܯzEVt"!�g �#���Z��q`I��ʬ;�cqw.d�Q/c��@Y��⮐��	��{��45ߖ[�0���U�M�}������+��"����&[�E�Ě�\)*{,φ[��T�Z =׏^�k��ֈ<���C2{m}��u֖�ֿ�6�U�]$�{$�$i�]d=�9OsY۪p�^'�@a�)���P w;e�S'I^�%��#7?�,��h2.h|..��ȴuL��^e�C�����V��<�ZH�q���潗�k�F��H��Ԥ�<�y��������G��('���}{��	�{����n �	�:��uڅ��{�/�ϵ��>糺m�2BC\����	�����X�FT%�H�ݵ���'*����G��1y������b ���^U%�J�.R[T"R�ڜ���n/�k���j�T��������w^4�[�MZ�sR|�����6�~5R���ف��ڳ�f�Zm��?�2�uѪ��dfR��9���Zat�\�}�_�80Q>w�?���v��L˵��T^��r\�==*g��'L�AZ��W14$��J�1��֤��9��-����O0.��!7�H!㪤���8"kE+N��y�jZ��,.��*��H +�=��=���`�6���i�LŊ&�ٶ����y��r�Ϟ2*�J�U�ܝ+Mzd�J����X��ݓ����+ � m�'��J��k%�Z�t�T�?	������'z��'��r1�$��J�$�'��|!^&�X��=�ҶRM_�t����)��g���r�-���}����@����|���
:D��	�QPO|y�n����Hd�JAYB(����*�Z
|K��9�dA���BS������51��{�c1���,��P����-��`
Jt'�%*/M����@d����N���}��ح��bc�ڹ�����qKCesnu��R'�o����سqLl?��S��BruC��a�8V�әat�TSe��8�_z	�nv]G�\�+dB�f��V=���0оS�N�]�Ձ��K���0�J����N�U<��#2�7^֊Ј�ܠ�_����xm7_�� M�4b����{��ِ��!��㆕)������NM޲GK\� '7^�$�2�]��?�Ǐ,�Ѧ�*)_Zҿ*\^�|�@_K4m~�(�Х��*m���	�T����bp{Q�Bc�Ȋ���g{���pa���C}�7N��y� �H>��0�
�b����q�����2ˌ����[�ekNoai�ު���@�����v�ɰ��S�n��w�r�1���
��i�� �Jj��e˺�{�l4����wn�+� �]�n�l�.�ώ=��nn��T��uj��]'�]^����=�.�� $����+�	]ԕ�K�ݾ-W.��}��L����4�
��}{���'n��h��s(Ѥ���n��#���}|fS�;�j�'C[�R(���9�-$�b��H���FƵz�~���j[����6���{K��2gm��x/4��%b��LGW��)����8i����)�S}ie�d���j��Y���1~�<��S��G�q*�)�)Dz:=�:�U���6�1�ρ~�ǣE�m�\�XS`��dU[�HCq��_D�5,���Yd�8!�ɗԾ�j�M��b�u�ܓ/(5�9̒C�A����n�*��"p��oCv����l���j�E� W3���6B�3�%���O�l�yu�0Hn�Y��(��N�i�a�R-����%�h_���" �s��.<`$52t���F-��� .�{��)'KRA��V#O�	�XUKM�HW�=�#v%E�k����{d��5 �9D�
D:����y�f�էS�'� ���7��?����K
�:&�L:�#�[&~��'����>DR���x����ܳ���D��|��/�\y*c)�F4,���$��tk�X߈9��8���mv&g�+ �h[O��<�W��S�C*�ը��]6��{���۷I�R�P��0�PҊ����D�*��M)y�:����pQ]Ĭ������"���i�F1[=����jK#{&o���>�i���{J������ ����4㣆|<�i�<)��߹������jYm��n/*%����QZ��{�+�s�
�����3�e|��d�IǸs�򥡺G��l ��g�EH�j�P�v�e����5~U�b�¥=F��g*��+Ɠ3��=G/�gS����w�{����~�IƗ�D�w�ΓY��I{8Y����
NYnm-����u�d(�'oF��BJ.��o��Y�8ȅ���	���:�iC��pҞR�'wpXA�/B��L��W��ʘ�$�ԗ%WKha��$r�u#��IݤQͮa��R�������
�eb�� *�98��s�=`\l���q��W���Y��Do���'���D��:.��(([_���QZ[A��{�
���Iq́ܩ\� 3�<�nb/��	@������ѥ,{���(g�*���Ԏq�{�-S����g��Sŀ.	z�h�-���<�3DD�s$�ΗdU��/e裄���z�t�_|�����ض��"Rf�TO�O����<�{v�����9��V&MJR������b;/sRu#��m |��@1�P����)��&�{����@�r5ɰph���ѧ+ў[1Hq�b�2��
����γ]�W�L��ۃ]R��� �������G�.F8� �ݶaq�|��l�|�#R�Z0\��׃#��Qaa�U+X��ַ�\� P�bU��6�I��ӈ���V����UH�11%�|Yj��?��A��R��b^���/M��]_q�Gߙ�6����h���q˗��A����z����������پ�
9\��3�a �"VW "�k>ll���}���#KZ!H� &l��>&�*�J�� �����a�����>�.hj�Y�:*K?�T�R���4vv��U�_X��F\�!��/�#�X�l�$Y5��ۺ4��Ge!3���f}��U'��������
��K6��ի������Uw��>�8N�M{d\E�]
�h�JxH�rO�n5��:�	�\?�͔���ל�
S �˩�ߙb) ���g�7�>d狄�yur��\�l[6[�$��BoR¤*x�s���j�x� �z3ܘ�1��^t��i�P���^s�nqځ;��(�����-[d�Η���|�>�*ە��-w�\5Q�<q7��9����	�y͋E(BP��w����	�w�|�R��������Yq0�MZ�y>���y���B�9�g5�8E�����qÝ��]p�Iyr�~
�h
e*9���xY;>6�:K�q��5h>x¤mb�эi69���n8i��IQU�	E�Eݎr�81�Ѯ���� �v�G��.�వ�xd�r�����)��<��%�!w��=�d���M��.��BN=�szfY�IN���ʧ\/���:��]��?6d�*p%@���D!R,�h��S�pO^�� ��]�"���g�x��P���8�Bʾ5�x]|�7�F�H�"�J�[���ܴ�Z�ظ���@X�5��-�RI�6�{�4�%�;\���7��Ƚ~�W당"�7��$� ��Zu1��]�U�C=h�o�o͞���TՊ��}����g����0+L�mev�i�<�W�xR�B����W��dwܒb=-��ޥ��w��u�0\����z|T��y��[Pdܛ��PZIR���D�\�0��ה�����#]�bE&�ٷ|&�<�@� M�L��S��ڸi*'e���Z�A�ùŕ���*�N]�Ll�f�V ��)1�Z���竚M�j��ŸY����'c��Ԏ9�u�K�UW(�%&��`;G��ϩP:?��wＤ����hZ4@b-n$$;��f����b��W��e9���O;�׌��o8���Go�|�&��D�T�J��^z�K��dm�����%m�=b����Y��A6��$xs�#��`�H�b	P��S�5�����!>�~�ۤ�''�ʲ��~.{o+&�d��8V��
\�����2�
�3ÙƤ�"7Q�Ce���(YP�߬J�޾��}X]Y	s�VntT��Nʕ7��^��ۣ�F�p+�]~2�/���������n��J���h���$q:R��?��3����D�"5>+*����(Q�yts��W�~~���~�k��G���㻦u��]r�+kB��Ç�gH�iPM��8uo���W�Mff��2f��f�0ؒ_�Tx�����}�si�YV�A������Θ,�l��ی;+���~�9�⦪2N������U��}-�1T�F[؟��8��̃ws��z�nĨ5�	���܂=���k�6n<���՗X�Qy�HO�ܽ�Q#�H��?����/ވ��)Zұ�F�TS?���_=~�־_!�q�mH�^L�77��~��%����95E���g��ҍI�WqX��L���ɮY��}�mr�e!]�}��=:���$w�[�~0tc� KoM-�_�h�Z�Zf�r"���ӟ�d�tn���u���EcB"��qS7z,j���÷�rq�S�*$?��C�n�>�0�g��C��/��x���c[�����s"CR��{��-ka�	JV16.b�Sj�}�h��@�b���u��Vp�R]KD�$��%���A�B��������%c��ۏ?N�̈os{��T�y����=��^�l���e��0nvHn(� [;�D7�d������%�J7�j��%K�� 0T�{@�0C��=C�����o��u�0c����9��7ߌ�/��j��'O4���)�+�v�9��E�����,����� !~p�g̞�,��Ay��l��[���%x��/��;ǵ��N�``���������o�7[�?$b� �B�o19���o�F��ʔJ�w�朊����t��>gB��q��p�� �Ɓ3���GGi��`i��S_��~>��]�={v���Rz�������8�X�� �`�:�/J�g��h�>&R�� Bc�VёVNn'�d�M٠�C��+�"� kQ��<zB#��aW�O���1ceJP�[��R��'�vu�fŨ'Kk�!� e���#$ג�烳�L� e!a�՗�*���%����@Y��+��˿�����{n���s�'t��|�|�-�|O���B۲h+	.T���6��n>y;�v�jȣ�]7���v���e��+T$z3���,��[�(qn0x4���õ����]Bi�H9�������
�Ϧ�w���θaRV!�������Y���c>�Jp�N*�V�G�A�Xz���z�#�!����q}Əv�`�b����"�1<���<iǈ,M�-=�Z|�[��k��?��>�L����Dh��wr"��♗�ƙ�"KHɝ�����Q�'��a_��R���`�G��k^�J���[�V1)���"��sdH���)�@,�\���b��?H�$5İ$Ѫ|��p�����pr4�T��\!����b��:J��P$8��K@��zA��>�q>� ���s�KxȽ����b|��ch{����d�D>�5�W_~e�Ol	ۖ���8�6�����{R�*J��F���a�^N���������c,���:�JV��I���=����*��R�K���bIhW�q�Ap:�{���T��yWiq�m=��֛[��]��/I���u����)^��]�����8�*�Xi%Y8�A��x��;o;�|��L�g��_�k�q���EIRS����nY(P)׀8�
�T}�~�d2x��ų����	kGr���1ҪP������mE�l�QWqQO�]���"��L�v�-�yX�K�؏i/���pqe:9R�L��1A��)`�"*Ū���Q���UҶ �)Rc����6s�=t��cr����������^}�)�Z.8{�Ԓg>��U��@�����.>����&g��0j�bX���;���1�=Q�:$1S:�1���}�?'������`���*-$6�^�.��?X#�'�!9c���kـˎ�����JV'a쭦�_�U�O|��Q��V�"��T�K	-*�l�A%�{��k8��������b藡�7��[��ۦ�)f����Z�����8B[P�7^j��v��v�KŮ�Q��L=y�喸WŢ1��E�3�@�)c��Å���8���+Cow��<��>;<������GשOG�pA>(��x�R>C9�32��]鷰���U��h�*�w��K��Z�9b�b������F������Wh����te(�W�����i��;1y+�i��+�����[�O�J�ҥT�BE�*�&q�98�`E��ܨG��+s/0M����@��T��~ٗ2K��E��O5����K��n�E�ͬ�[` fY3HO��'�?�X��!�2�2��9>�7�5W)��C[��Sr��ңR�:�{]��Ѳ�H�=#�j|�U�Ɲ��؍���ֲ�B����;:�1�O�R�9<���͹Yq4��`Ht��Ð�n.��<���jՙ�-ʋE�Y��,��P�Ns���k��c8G(5�?�Gۢ��P���ߣѼ��m��O������*��e��[�#O���]�)e��E>nr���q���# Ej
?Ш���^�6O��u�v+�a�\�U�"	՗�~g9�a�V79%K(�*�<dH�{^��w|���h��P���������:|���W1��Q����@�R�ኈ͙�Lڟ�Af��-A���q��)X�9�~��R�r��*p�L��p���C;�;m��U JV�^�%�Q���%������MĻ�Yz5f>���z�/� ~�(���P���u�4")s�u�|{(a�  T�8�����a�ϛUa��>�+	Ξ]����}��nV��#V���5���?��ܬ��̕���'�\-�d3폎Ȳ�E���NO(fp�����[�����
�P��bØ!��P@�8��K�\����JF�KW&8��њ0�^��]�Γ��<��Uf*A�k�v���)Yy���s6�|}��Ɓ�6������5�A>>�����Z�b�����B�{��tt�0�
�p>�;˖q����j2��Z�d	��~�������	���	F �x!ݰA�vC����H��c����N���6_���{-I��X4R�h10P��������9���.䈞��n���{d@y��+��-��"#\����CVބd�ucC�y,��"���
�~	�T;8l�ʭP�@���n���7�wU���s������;Rr��*�j���q��G��T��ʽcHJ뭺^Ê�ѣG��PĠ�*�����4F����J�q����!�� p��m�*�Q���<6;��xԠ>:qj�ٍ�62�7���smVR��)C�X�1,��n(��<ݾ��n!�LG��P�w��<���s=b���0��/����ĺ��+5���̆{�f�uB�vu&}�x��59W��:��YP���4�) K�+}��e���vE�g�e^�,���?�-�w���y�ggZ.f ~"���\A(6�-�p���m���k���I+b�(Mڧ&��T�4 �5ıu�1l..���dbmHպ-N����9�̴>���u���9M��Z���Vq{q���|�8v�L���ƀ��pQ��K���z�:��}��0œ1��ºN��"�k�Y�d�9�S�4���UE��`�3%�'�`�J���:j� �C�C<���O#�U1V
���MI��hʨ�HiZ���������_y^U0�U�6��=��=�h�`�oN���p0��H��} ��hs��>hkEu*�0Ћ��ƵPt�4�9*���MJҖ�U����
t^ܢB��E C�ej�=S���?+�<�FR��#��p����A�6��Mq�ap�_�n���)ֆ{HJEX�y��Cj��&��6e`5�0���z+.��/o���=4:��@�^��,�.�
=�1M�|L���g��;��i��Z ΒP�Gp�Tjb%]s��w�K��1�o@1X3��z��jU�a�m~�n���-��BP˧}��К+���@8�k��� �t�8��{@�HƔ����A�zE6A	ni+c&'f�If����ڟ?�ؠ.�ݍ5ej���j�{��xO�Q��M��G����h�MA�x=�T[�J�������C��)('W��0\�#�QDki�J�O�ll��h}L@m� f�gN��a�B�5��cn����߃�l��@|u�
�c���_��mӖ�+xh��`E��i�^�ާw�Ao�>G�4^���9q����-�mU��J���~�ņ��FuV��qzcNTb,�L8����?cx^�Kt��}ZK��Na�tu��
KbY BP1����
A�:�T]5�"/�.NS!��Z�z�8�d�c�r"�Y-����k^�z'<��w�;�)`�0D�T�G}�N�.?��|≭�Q�3zԝh0�I��Y���ĵԓ T=�!�uX�#�G� �Ǣ�1*LB���ɣG�n&�F�E�/�G���S��Q����C�TY+� l������4��+���g���`3~�7���=�,�L���iU��0ҍ��_�����Ya���T�����U�u#o�d�v�jդY���� C]޹��j�v�a����Ӏ9���͡���-�9�`>��W� ^\m\�<��W`�vpgbauT����-�� ��[q\�Z���ɉ�x���������]D��˜��WB�o�k�ޑ�t�b�Q�<P�g]C^,�6�E]f�4�[��*����_
U�WWջ��H(FF��S9$ba�}I)6F&R�ד�5�|I*7�W'��8�m9I�m��}�a��CM��zN�->��h��&��*Zu��a���W����:4�)����]~�	��D��afW!"1s�%՝�$��}���^���k�ixG_mXl���5�oyF�P�4L��_~a�x0"��o=K�C0��̏i��Y��d�CFU:�xd1��k�qC���a�^$T����1d'$�~���{��Y\J�<R�%�b��Ҕ�?4��`��R0��fS������7�8I���$GRI�\�L�,D���vE;p{�/���:g��L���4oyb�{�ݨ�I<���ͨ	}��\���dl����k�\mH�UO�t7�=��js}\�.[��q4����F��OKl^9��ذ&g�R�Ѥ� �g?��$�1#��z��w��0����R\�*�#�^����w�s�#�8�^���8��tn��
�����6	�����ӏ?��C!��([F]:8�voס�}�
���9�W�m}`�t�,�D�h��TvU�Z_S�4Y{H�^㚳�2��Q%G��ϗTZ�]�pxi�P�f��Q����H
��pASC�&�J�����^G���������j�<K�ZعK�q����������8p�.�>���M$�ڴ���d�(Sb-�f�ܚ�^��~�)���/��Ž��Έ��1�*$ݖ�����K��U�����zU`���Uk'�*]�`����&BE"E}9��#I�>���=<OUٍA\��#b��=�bb(n�R��[�jP;�~�	5�a ���<.��t���0�{�)�2ڼ���u"�,/�6Z�3!�*���\0cZD�� �R�������{��*P���ȩ7�\	g8T ~+~�V�_+J4��&��8�Z�6���k��gvms�鲑��gN
T��46���6��˲`(zW��j���-�>��1(r:���v�S��D>2�$��&f�4~[�LC�8�E��K�ӤHuڅ%�X҃��P��9�<������g��x�%'\��WӦ��Rc�T�*̓$�����Ȗ�l�
�D�+�k��F�T�)���f����s����s�Q��e�5����j�K\CP>���~i<��,l�q�ya�7��b�8Z���"�ش�!�q���ru��X�乥A0�B_�I�P��w�ͨ
�TbGj:=���#e헟�t��я��S)�j�������k���	�"�wE��?��Z�%Z[O�Γd���;��yZi*:H]O9�^�!�;+���y�L@�aH.�qrq������gp�p��yx�0��)/� Js|�r$G��1#�ya�M�'�)��DID�������sL�,Muj/.��M�7mD4���:~ľ���M�3@���6���R`�˳�XSv�D�(�54��*�hZ*�r�&V�L���,(�sV�+*��j��:��"o���#%\1Gڟ�z��%��a�Kk$zsD%gk)b'�����χ��|<�H��,�&��'��Uc�T;=���6���`v�C;|�қS>{*�����t�}���>ֽ,J�(nں�,r�#̨�Ћ7�)#REWaPeL�FH�������û�$ȫ`��eC�7a���Ts�\�ү�������u�o<I��#�`̔ɣ!}i��ژ��C'e�Ee/�}�3�n��x�p5�)��#�!m9qxaX�@� �:��$�3�=Z&~)��1��9�at��0g�n�5�>{�!i�*R����{�*�]��V��������Xd�-����4d�ԊYҐ.7s����r��s��M������߼yW޽{���n�v;�1����U`����d�ؤc����o�]2s�c�PBЃQ�a��G���M��P�}���U�KU�sy��^�2��R8��9=9��&��ޏ�M���u����n�=�r�4�D�7=���!՞Qg�0S�O�{�1O�!"�B!iq�YP���������{
��2x8O`��ɑ��l��g��=�E!�z�M�~������fF��!T3�m���)�B-���<�1�T���)<g�S{Yc�Ve�n%ߐؘS:QMS�G�uӴE��w0��YSc s�D��OEP,��ż#�$��	��Q,��`��X|rk򆬚#
#�*2z����ݤ�8�wX� l���׍�bj�GD <k?&�'�	u�P��7��d�.H�D�Ti�*ir>�<x}I���ZiI��;L�{
�pѠ��x����j�e�&D�@݈�Є����n�Z�Jnn|��S�1a���4�F���"����fJI8��,��g���Sm����u�I�i�����b��k�Rv�H�)G�(�Dѷ�(�Hڮ�W6��#�-i�0f2�08�b��j���aL��G�j^�(֬4NS�Y�n��N��m��KqKm�ܓ�����V�fJ����",)]h�@���`��sS��,������O��3�an��2���>j�,�7 ە,?+�l��Mx��h���TH�ӣU��.���!�.�A�v;���hW��G��lB�P<7#�׏(H5F�Ɖ�^�����"���W_H��5�(����j�6�>���Ԋ��ʭϷ����z�� IPWU]��e#�ֹ���>��╊2�(}^��=o@#���R��A$d �`X�y�ɕ�x�C���u�zY�~��7���FZ�,�t���/^�V���ܥ/�����(��8�"��.n��j�kH���v�9�W�Ţ�MD�tt�Fi�&���F�?)�S��"��:��cv�]#����%��m��>,�S˶mR�`��	eS'@�4�us��ɩ�:�ɉ*#?xD��D%>?5wy��w�gP�0��a/`_��^H���ui��y�Kd��r�;YHӓ� hR���E]��~��B~�c����oֿ㐼i��2qm+�l��Ş	��*l�a�+e��.�E�r��\E/̐rF�(B2�����3���ߒi��[����>��GX��~F�)��䆰���#�4X��\���s>y�>�E-�u:�~ly�&�����n}���7ߚ`�w�}g�
*���zy`�֟1"�l�_|��Arc�[b+��'q��7��ESt���W.i�E��>�4C�ԍ��u2<��~��#Efs.��$C���YB�����ɉ��V(5	E*��Bup��i�������D�9��h)�FW�`�+��\C��Z�c���*c���R7(�%/�/R?S!���,&� �_;ۧ�ŦN$�{�8-Re���&���eIU l<��v�i�p��t��$ں�<y=��?C�4�a�����ԍًG'��й3��x(�z���(�SSW ︁��U�蠒3[<B3�p>[�I���ûw��T*8w�8�}���@C�s7t�����Լnj��=�W=m&Q*�����:��V	��H==�*_�rtu90Eh�8k}�vX��iܤe �8��6�F��^��������jE�}x��5&���*,t&������z�HQ��6QΖGF�/���juX_����ܐ��C'Ux��*�s��ѐR����(�J��j~����F	�!C��(|^�Ф4'm��N���.�5���)wj��g:��A����iDo�w
$����ِ�xc���{��Rہ]O�Ȳ����[���(W#sXP%.[���u-"���7����"�\2+e�*f �����9FD�3g��NMΊ)9��6�x��\�2</
�R6N�b���=�Ԑ���ċ�tV��I�rfxD5���V���j��o�:��Q���� I��_.�H)C���J�h�&��*���	�Tl�JQ�O��Ε�����Nޮ��3.E��z-R+/M%��t��ڸ��<�u����n���.-`�;� KX�$��6ý~��.�5�H#��H��֍��&��ޱ[��,�a�R׵�P�g�Y5/κ�i�)fŽs��U[1�|b�j�J�� q�6hC���60*�-T]]�wk:�Ť�9��k2D��J�p��X�̬�k(�]S�#>O�ugN�|�<]�<��K��d��·�PL��0�����mp�`!�U��I�	,E��eq�2>s^�=��H�'ߧF��u��5�;����5�Kma[�X������z��̩~�O[���4|���5E�Y���h=�ͷ����K�t�
�����9��c�*�9~�^�]�j�T���F
�oJB��.{�J'?`�c��E7���5.�k���k��uL�Zw�~��Ee��9�FVv~��ܥ�(�Yr�th�y�C���:�{}�2����kae���W�`�م�ŏCtß�}m�;�Fѭ+���*����X#�w1����n��yCJ�O�A�kt��(�0٦�['@'�E����6����M���2�Qt�(4�scQ�q=���#z[���G�fOC*��������B�,]�r&Z�t��8�I�h]���T=� ��Gfsj�AU���`FfG71_��(	n�0Mda��2o|v6�� C����>9�����7��5aM��u/�Lf>V��9��iۀpp�m�4�v��D0~�j�3k��it���Iy�U�	����U@�&���>3�ɚo����_\6���?5"ޤPXŐroz����w���]I��m��}Sy����/Ν���b��\a��t���v���;W�ñv,�;�C:9�>� $�4l�,I�K��ܨe!��qyXS��t�n��ϑ�*���q�$�9a��!�����F�+�	��v �I3���͠��w��w��?���������h��At&fD���6�f�#"0C�ۯģ�RJNc3�w`���Å!��?��	OXQ�h���^B��`R���vTP����g�	0p=ۂMD���2������Ed��<���ÐJ|EІ����߫7O("�g8XW�v�0��L�¯S�T|UF�]��beh4	0{QA*����o�P�Q���,�����tV���\�E*��O������
�짳���8�%G?�\�>`]-
Kd-���0C:Q��9��^��mH�N�YٙhH</�g��P<S��V���Z6���wCU9�g��	��:і""������e��l���tM5}�>�sC��i$(a�����x�K�V�cDL��ؠ��T�T�¹���#�>�����x*=�t'���IC������vw&�l�-��:��\�NG�GS�_S�k����u)E@=������&�L����f��Tv��}���%�T[A��bbQ<ĵ�����&� ~G�����ɝgm=:�KE{�C�.+�=�Kr��GQM��8��mOO��8�߯��5*�����{	n++���������z.\���Ɯ��T�.c���MZU�3��8G�5X1���ZMoo���I�G*�a�OKy?�F����k�8�U��z�qΚkh�j��w�%��)�`��JQ�c��ДAm)L5�Є
�Hgj�sxP��H�ƿk�2*-�kDj
(W���IŦ��|�C8���ۼ�J���:���؆/`�v,��Z�r�Ar���w5dK" ��D<j��z�"n<i=�F�W���8�]xU��H�T����+-sN�䠹�oa����hm�
ޅx�4&�{�OPT�_�v�7���9Q����SdL��&�֩�K�|�9�:T��r��Q�\%Hѓ�kFUK�K49����%�&��v�a�^I9_�-Q�O��[X��f��˚�L#�F�m�sV�y�m%�V:�4t#x���'&~^1��Q-H�97���r ���l�{�])J{F�<��۷A3�uύԕ�H�A8�gkrr!y����\޼}kFgS�7J�P'�y�c��ɀ�T��0�x����Љ+�)f}T�~Op^_�������ޠډ�u`v@��߯����˥s����s�r6֧ع���܈F�:&]>a����!��y��F��>u�I]ʍ��ϼr�ɟ��H#����5EH<�">�.Լ�`���.�f�D�z{ĉ�G&�� B��!��6܇�gG��I�P�����[��4OQt�������QJs�n�X�zG׍��߫�՚���U�������J8d��v)Mᐁ��k�a-V���>(=u5����d�c9�)ءt6���F����`-H�i(N;�2C�}����יS_��jOԺ	�����Ë�R{�ʬT��lƴ������'�����l�����=�SoE�38E�6%��2�$���`*d�����C�M��+�K�jB�u���i�lL]X-�=���Q�u0�oo?2���#MJSt��e��n�T�:��M��&E��i*D������Mx�R$̞�����>6�u(�����L�unң+�o�܄�HY蘣�&#R�p6K�Fb�H��yp�Sr_�ۍc��.�Rb��E�`�pY�H�a\�A���7B"��Hka
���0k��}���-�W��W��Qh<�v�"�:�ͬ(T����:��`I�n��m�x&"YTt�����������훷A��\]A����﬏�9�F��"�I�K�\Έ�*��ˇ��_ߛ�Tt��a����������.�\��;��=e��%���d9�ַ�{fN������eLy 	e4%G_�}��>�;ƸǠ�;�r=$����Bm��~�9Q �^{��믿�b><Q�����mo�>���z�J�sAD���u�W�g+�s���8M��z�xI	��#l��o�L��j)q6�x��jr?�uKo"�E$�k{�fE���zw�{S�P�d+�2���gt�қ�k��^}?��Lj�i&.����hty�_5V�,�����7m��%�ϩyi�n��;&Q��%������j�E���'��k�`�\E�C�>�JO�=�H�q�@����v1ي;'�	$�u{�C�բ�yd�qOoh�M��S/��hT�K����U�p=$3�`>���1�N�?ygx���&r���.�I�M�n]#��u�P�3��iZ�N-KC�(�"'<��<p���,�Y�����~�������60���5q@Ιm�HǓ7�
{ݠÒ�B�~�c�Rt�<��V����.����(=����ڥ�����{��h�y�u���Vө�>b$f[6�I������Xk�3��0x+wN5���v�5?*X	�l�z4�SM;��j���a���B����(~9~��'�4�����?%鏀�(Z	#���=Baz�0�nlJ�8���n�,%�tK� ��a|��h��ru�Z��aQ�Q��� ��� {)��76�ҵ-ʘSM(NC4v��dj��}��i==i�H�\FV����զr\Dvn��C����E@v>��B�D`@Es�5 j��q\��HӤ8%j�����/0�����՚�,���ѽ�R�_u�\�#F͡g,�"����^t��O���q�ށ�u��������+�"g=F0d8�QzM�j���S;m!�9�YB�W�o?TX�p\���o�����z�zF�2��A�����N�VU���[�9��T2����Sݟz��o�����|L����}�j��O� dJY@M���f`z����Y�Lg�p�D1.�wTJ����G��H��,�E%�
Ye)�y���K�W�����o5�o����ٟ������Q=#�s��rY�����<r�u���$���!�GO!��Մ���`%� C%`�D��u��E*��M��SʞɳQ�f�/�4��w��S4qPt�ON2�~���ߣ �۽��0}xC���,2�ϑ�xo��� ��E��&;[��Dn��tY�9�ay�*�&�02|�,�US<a���6Jt�Þ�j�틗�i�:Dw��`�\^�o7v��wQPI�.>�*��>�k�9��!���K���E��u�{YG�E{Ƣ_��lz���8F��C8]v9�X:�}L3�N�GFቧ-Q]�<s��2���*~j��E�h���)�&�j����Q���:���VD*��Kij�*���~?�:���ו��$5h�p[F�h-�ߡ�V���c9�5J7CC"���3�b��R7;��������N�ąz��g�i�!����Ϫ�Yy����|�@ߨf�^�&͋/I�(���� z�zIW.�W�#��&�9Q�����G���q�'7����D�D�Y��Z����n��Ɯj�T�^��q�[��hX�^S��}��b��MQ�H]�wRJ�H��z{[$����h.P�G%��ɚ��ڄ�ňj�NC��06"��l����ײO��"�R�4@A[�����i��5�X�_�*�ީUT�G����o�%ǖ�g1����{�L�<<O���,����<JE����)i55M)�,x��l��\��:��q��4��,�s�ZXfaH}�� k��v�x�XO�&�g�s�68ǳm��r��NٴQ<2S���DtM]w�:]��q��X�3�63{�u�?e����F��垭���\�-��B��M/�d9�Y�s�t)��]SqƖe+��')C5a�M4Z�'�Ƃ������M��%~���h��� ��%�9���C$���BUY4�)1��铞��[�x��MDjyӺ�Gc2��:���=G	K�
���^��W�-_7@㇞���n��uD�@��OܹRmNimf�~����!(F0�8t8p"�S=��n@���m��}V��6��\�"#M�4cǽ��w��K_$���!���,1G�.�Rd�Q}��'�N��x։R�}�����Q�Rؙ��|�)FO(��i�@߬#%u��3c�"k<�N_�uu�4�ù�����Z�d��8�f֬#/R�r(�^K,��P�gp��� wL��J�b��}�ڂ�i?�1���9�M6h<6��&�53���v�;�7SZdnuV8�T� �EMdQ�yƵ�k&�±�Q�����H:���٭���>�-w������)L������?y�%�4��c(���s��9"U�[{7HGp��%�g��Q8�a'�ǖнύ�h�cڃ�Gm}g|��A+8����Rlo(�?�R�nLU�Tj"7�lz�t�ٍ��!z�h�<;��bw>K�|P��6 ��E��Ř�ym	� ���nh�N׀dw�%D��^���wvXLKz�t
����Xt4�(�ag���g���]��Ro\����XO8Q��9G\��EN��&R=��a�x
N���SVz���..N�G]��7:g������5� �Q����\�W�V>���'iڀ����Y\��j��޳���l���oo�ѡ���S����-��4%pu�ۄכ�Fr�y��~4�ޭ �ܺ��<��B���ޓ4�t�e�4�ʻ
eH�Qк��H�U���[����jC��B������T�4܈�^�ʘ*������"����M�K��ً*0(�b��@�!"�k,�@q}&W��Aw��mnYq��u5�� ��Â��8���<}C8
��VEJ�F��ܘR]h������G?���&��'p{�kC�8՛�m���$��p0VF�3�!�5�@��`�aP�T��ϱ���)�����$�"@�` 8����iNִ)�7���B�HB�k=����-^,�s]�v�g��'���~{���d�ɌB�	�	Eӑ�6�{���Ģ���=�j�8o�f�F�Z� �K��Z"��]�W�QG��X�f8�1ǌ0ҿq��G!�E�J�ܫ;6�8i 2����V����u�ǜj{�QM�1Ѡ�i�:�9Px�Lk�ۇA�����dkT3Ar�_�X(�$%���9�0���~�H������_�2J�
f�����L�M�wM6�|�F�xf:�l�_�@U�k��	�t�n��������H�$�1W���2�R,�rI�_�eĚ�����-�6�����WKl���Sy0��i��o�ug��F��^�i��bG�<`-{Ӂ�qн�l��K�Z�VP� ��OA���o0F;E�s�'g��5 L�BQ�H���G)��"-a��'(���-��{���9��g�*�o���68L�Y��&�1q�o�yw# �,�㜪p>/C��-:���u����$ڽ���_8Ċ������p9�.�$�����d�
b�6�WG�ZO�#(	G�SG#���!����;p�e����ं��5�����#)y�s����L��7ERM �{i,���_�^�j���C{.�U����Ft~�����3Q�v	��ȤaI�ß��kŷZ�7�vG�{Q)?g2�W��ƶ���_�v����m�\��`��P�G�w�q�h��.�[X�� �%��HE�xE��e���b���M���B���x�����ݾ��
h�OlU�z�x��Q� G
AD�SF#��q�}��;;h�?,ת2�Mf��B�/�
/C�7�r��~K����]�'Fp5��I��<��r!����)�]	��ީ��SY9��
%������&x���wC�ʽz�Ma�#�������ڇ�>���ѡ
sϮ��l���Q\��V�vJv�L#��$�ڐ�@� 6���	��0����~��fwއ��g!lp�q�ǴS����n����lE�Keh�Cʂ���F�h�L�� �1�V���J��֣Ud]?��c�l+����k2ٯ6 �a~�������#��%���O��MR�y���O]ǈB/��F'�"���%��t~��.
�9|�Q!������f¤�����$�3�t.�ն� �5��JX��{w����UC��-����))>��cH[z_�Η͍6��J�KvO��%���{��X���hz`��z�;/�ᰙƦ3%x-��y(U�����L�l�w7'����ZL�ٮ#��:"a�/���Kͥ4�ML�$����d�/įս��O}p�˾hb)�s��ud���.��a�u�S��.�&�#�·��{��F˴<�^zZ�S����]"�bRYک���%�%������ A��׫N�� 7����ԝ����L�p��.��Qg@4%8g\+֛i�.����K�1���5@��3�I���N�u��}�3�~F0<��X?��i��I�1z,�2�4�G��j���#�GƮN�e�j�>��T�tY>��T�풜8�K��K�^�����|z�ҵ0~���W������H%j�8[	���n+UQf�8I�5%�s(A�֖_�}�%�L2哃��}���������߲���^j�M)�:Q(��I:l���i�TJF����w���Q���m2g#�i�Z7f��8F>�<a����ůA�ۜ�o�_��D���c�f��)Uw���(@�V��Oc��n���:EI���������3�?�#�>�=��Z<�t��D��?5��|~0��$��QG�7�ԴA?£��Y��>O�<ԑT�i�g��r�����QpSS��Q[H���d�y��T���K"PЇpe�"��:U<aer5u�뻈�Ek��:y��H$�<g\�g�������o��jޭ�LJ�4M# ��R��h3Ϟ����Q��u<�A�Q<�T�tC���P��0��,g���@��CFimt��B��vpp�]�z����`�l}e�ǋ�r��(��)�cxwp�TT���%�&��z����H���������b��� ���ާ'�8��UU��Q�]p�$d<�)�����o?��E�~إ�ZD��c(�_.�s���T��"�NDp�H��j�%q������j�7qΝ���]lQ�*J����>�='��`KPx�}���	?�����c-�n��	9�������.+<�v�4r9-����������?
J���Yޝ���Ϯ����G����`��u�!�c��⣵��3��vf����l���Ƥ	�V�Z���4E�\���պϛ����$=9)��	��\��Z�uO`��;����f���І��'���O<j#��'�I�s�	��Z��g]�Q����)�I%n\�L͑�M���F3�iDJT����B�mkH�Aj�л5��uU%�x/�s�66W�6OD�0��!�,��)�lE<YzϹP�0�����5�8c��D�y�i�J��ڄz�
���0Gf���[� kPo�+1"�.7�B�O�&#�E-��j�� �ZFΪ0�)���e3l�H��$�b-5,u*���%�Ȱ/&6$7�� �!�7R��=ͳ��6USy��9�1{|/���M��y?�9
���q^°��&(kj�|=eH� r��ۃ�Ꮟ��o��7v�9{�~}]Mvǿ^Vߒ�l�7��m+�~��_S�z�����<;C*To�u23��a���n�(Q������ʜ�N�s�s�F՛�n���Ҁ���3�Ty�>u��R-R�	��a�^���q��Z�c[)����nw��9�8����Kߴ0�x� Ȱ71�%�,<����܄7Q��a5���N)�N�\�hK�Ϳu�O����z��3o�|0�O��������!r�3�F��pF�+�H�]$��������Ǐtalp��Y>d�J#	�-�k�}���C�/#��;�Qp�%��9Ei�FS���v�k����T�h8��8��4���(���!�9}R�Ӊ�-�K�7�(0��O%�gb��R]��~��4�&��ۯ����T��ȏ�?QyB�sۦaf��o�n��J���9ʊ��6�3����&���6��0�Qh3�~�z���K�L��+���>% �~y˶����1"�q�ǽ���c�����y1�͛K��}^�^"@��"�t�qj/���J�P�MA��ee��O�w�����g��Ŀ�*�@U�gWO5��O���;ǒm�%#�q��w)>���s}T��{]E�Qׇ0�%���9�	�*3}uq��fT�-�Ґ�MV���ʏ�.��L��C���<�ɣ��*�"�7i�"9���p�
9s�g�7�8��WE�*�ܔJ��ٙ*�TϚ���q<K���g2��A�ѝ�爵�`+��Z�P%Ew���	C��\w��#&�xj(Ǡb�al'���.�zȂ��<`Xe��T���>tK�,��~�Iےv�M�-ɳ���Mq}LU���0�\�-�g'N]g(�:u��.�`�0� T����_����N��J\=P� ^�z�"��d3����#�/Q����OL[82� ;���Y�F�	a��T���	��;if&����-���3�Xp�����4�`���,�2<k.S������)�*�b�{FTPmxEK�U{u)L^�Z��%��=|D��W�qP|�'^6�z͆��e
�*���d���PK7)�T�kէ4���H�0���o.�ei��UZ�Y7!��|��3{���P�d�DR�_U�W�D�-�M����[lVK����>'"�2Z�s��B ��J�i�Zoٓ�}�6�qW�-�N��H^��Ud�T�9�;{��5M��b��9>�0`
ҩjI}��E�A��z6�!���]t[�
�C#qev[�I;��_�εcw�p��=U�l�\԰A|�$��O����:ͮ�����瀭x?���3�F�p?��K���u(�۬!����R>ru�^$��j�����8@v��j�d�TZ���h,���Wg|�̯���{~B���	'%,��麇��Y���R-�[F��������޴��h�?2>��
:��:��A��hF&��s{���A3�1��ʐZ��EҼpy���Fc��t�v�`�#e��C¤rJ�VQ]GJO:��T%�oɶ��{}T��J�(u��'9�M�J>��ݷ�Y:����?��MC�<FE����պ^J�<�s���q5��y��KF���:h@r�:RCNI=���j%��ؼ%��,�4��11�n�,H)�Q"��g�����H�U���i܄$	3
�Ѽl����É�ˁg��wx�h���S��&� !L5]�i\�ͱm�Z�_jE͙c�{g�,�Y��:���ј�����KM���¡T���M��ދ�"��:7���:�k�F�uWזĎ�TZ/����k�kшX=O����󽋀{��=�M�,��s��z���OG!���ɮyy�dޓw}�=�+j�գv:�t�/��ܝ%T��z0�?����z'�@)#�%��C�G0����2��R���P4�B��.��9�����9f5{J0N�M�Q&�^u+���;K�I�
P��d�H%j����m��I���Eё�$�n��#/�8���ީ ��N���I���0Ҹ���_��^~n��,��a4�����3z��]"r�F�9�˿����8x�{�6�w<A�!�w������>X{�ٮ��q�5D":J��l��� ��WF��' tmU�-/�aQ�ܸMj�hZ5T��b��  ��IDAT4��mk�ŮJ���k�7BP����A�Ǝ;ͪnFׂ;����6-����0a_-��j%���.iM(����*8�Q!��>�8�b%�L��"u���H}�-���'��q�q��]W��#�T0��y��ѯ�랍aO�;>�%�������k߅��1$
jd�Ց$�2��鰧�^�s�T��0TA]K�8�Q\b �T�(|�� ���Wm�%�����.��ܲ��i,%
0��b�{�s�;�P2pl��k��f���|�dۙp�z�M �.�a���H�N� �韪�}��<��~~X~z�8^�y��(E?vm�@������?�`���~��A��ң��7}�b�"m�n?O�-!��:�X~������ǋ|0\�O��[s�'���ӈW���[�p\u��Iő!R�\Rw2�pp������6�%�7��}ui�R���
rⵊƣ�B������n#��,8�bŏ��3���d�w0��W��&�2��,�iGW��T�C�]�߸�J}QɗcA��#�4hN�62�Z�}����|�s(�*�)5X�s��I���}����E��@j�RĆ�}��.��*<��&>����}H�'���1a���`oj*��*d�����|z���2�Ri=5I!m�c�B��A�x��!�-�Z�B�ߣ��|6�9:�8���0OG,�m��cr"qs`LΧ��A4.:��x����-߸	6��)�r�n��0�go���33��ݠ 7�s#�|��Jd /;�:�0� D-�����?	z���I�U&��H����!y�����p/�R2�)Q^ߛ�'���f;@`�%�-�5)sq��F]����hb�-�^�R��fs���*�/^ܹV����qP��♍�z�%m�Ѥiq:ǵy�k�iF��Jw�d�3��?�S��L�zq���w�H;I�[A`쯓G�Z����\�qC���'�~Xm�R��W�t�X>A�hu.�7�7b�hm�4jd�����~ľ �6T�q�^0��c5�2��T8R����x�1�*�\�ݰ=�!��:�T��EZ�~9�"E���S8[��a_����-N'=ͦl`_�64���E��R�;7������!�V�RD��o3p`�900��8�V��q.y︙[�7o�2s�A{�6�6�`ja�7zt�,�`�ĈdP�9�8��B
��`'�m ��I������Ui:���s��3U�<]�ݙ��~��T�JQ�ka�����T�b��"�3��}�2��Q����޺!�3#)�)��gg+Up��q��FV$y���?Dz�ͅ�U���sBYp;�=���P��w�W"Vqi�4V�j�K�fR:]rb1�!h욵��Qvkɭ+Q	��B3�[;��B�ukFO�S\E�u�pJe0�˸�Oe���Z��l=+B�tZM�Z�ި!J>v�}�d{��+*Z7�"eFԴFO4Tl]M�c�o7G���c�gm���~��:G���E�wqI%U��^�~�L���KL@�5G�)*T�S�~�o�N�kj1��umH���
ֺ*:b�q>���6��)"њ�V� ��* �'���1�G��D���S-�*\<�G��uYс�m�����{��=�1Uꖔ����y
�N�<�ͫ��L�	�:� �`�'�x��G���8T뾼~�:7��f.)h���'�!�X��O:E�`*���=��S���n]��j���<�ڳ2�,8!a3,�H)}�T�x����&�>���Rt��0�	{Rt���p�g:��(d`�
���4m`�l�uE-�#|}�Ā訚(:c�*|^�_����n����=c\�=�#���7{I���xK�GNn=X��{��z9�yt^wA1���E�iT�K�����NjVEZKY��S$T���CP����߸��XO����v��Q�tcϧ(N����P5���{5�(�Wǔ�6;����N�Κx���K5���J�?�1��cp[GQ$ڼ��j�:�LҽJ�_]��F�"�ʺZ��o�)���h�Y-���[����2� եs�]�a�nXM�O���=p���׸����w��h��!�ya��Gћ�0�φC&buM�a[<��'���)'�yL`0�H��X"@P�4<b���Z�\L�e�}�ͳ"#�v��S)g�$a�d-������օ�лX����F�C�>DǗw$Ie���ޮ���?�bUo#W߈v���3��f��/�Msblո
�'}�Aբ��m��M�t�6�-.������e'�E9�>�����y�G��֜(�T���)̢�"A�&���1�[r@``��W��!C
c�lAJaj�Etٵ��L��`_�-*���`H��jjt��0��U7Q��7;��/6��Sb�yA!i��x�j��}�2�]=�WVC�r܇�\�}�{������[�]��^����*e�I�4�Uw\��N�����L��ij_{�0�S՟-2��@��"�lϼi{¥ψ�>K=��ԜeM�EUl, �L��M���J!�X'ۨn���'�����o7�rRuو�YS��R����7�PЁQB��f��NO���&A��?���z����=R<���)6��\5�Ŧ\N�X�4{i̹8�G%}P��4uE$``���?�aF��_~*��߽y�3��'�w�u�"�Sj���k�L�:�����/_���ֺ�@�
�R_S��៓����7��4�D��,�A�U�,��%d�}ں��E)N�3�q76�*j�LN���c���"�Dr��NG�f���C��{i�T�p4�PE��[�}tlT�*:1��
ĘQr55�[�q�3�u�����O?�lq�hf�Y��$�W7'��W���&�p��i�v�w��a�D�/&:R9!�TZs�X45U�'�^�vA����3���8$����+�����c��+&R���r�:�O#�����4�ؐ��z���o��䇗��&��!�Ȃ���}T�=�fZ�~�QR_��m��'�.9o��<e�g�'���,�&�������ތ�Gg�x���H��ro�?��QY(^��4
/��Gd|�'&�x����ޗ\��Y,%�u�%:5���N���Uiۮ��Z��o�S���-u6�ߤ���S���r\�(.�~�P�`a�4F4�-�6�Y!mn�]�G��ꞌC�~�]�%�,H��yэ�QՖ�,k�O�9]�К�Ve�0�����}-~_���+��Ql�jR�5���s�!��ZWMw�τ����{f۶��ĳ^{�&C��*AթR�X�$�+T�([k�`*��7Z3F���?,>��+�3�5^L�Ԟ�;�V�:���M�^�&�7o��a?���Q73��K�Ö�����C��2D@p^D�m�|��Tڿ�G���-�E}�i�%���:�➀�@/��F3��Ci�����<e�E�-5 _Mx��zm
	��+��S'1�=Ǌ
Cw��.�4q��mQ�R<]Lu���J��)oj3mn��!2/�ƩH�xC�GڈF`�j}T��)�n,z�3m5��
���v<�?�(ڍ"��;Í���[��	�k�w���#*�Rv)'>�H���4�(��oQh{�^�)4C�L�5���POؔ@Fk�#�<,�'.ȑ's6��"{��cО�,9�f��G�YzK�ib������W�}Qp�
Ք��a�#�P����T�u���A�V���g��S�k�6c5�P��['��Q("��4�k�}�u�>��V���>�s(���e����x���:�5�3�`�nn���>��0�^Nݠ��˚U�Q����ӏ?�
�"[U��EN�����#ҚF�����
����	'��'͵�G��Uj��# ��պ
�����&�P����kX6����)��asӐJ˓�MS�0o|.6���\���@�x����t״���P�,���v�cQ���T7	6DfA�u��EQ�KL#��ŭ/_�LT\�|&�Zq`M�V�T�T���aM�ؚ@�z=Q�8q�z����o����򹴡�Ak�l�%��F!i;�X����c�oMcN���74��
#��]I�l�	]�5iђ���q5��My����
���w�}�^ue+�	8���ׯm/=X�gp�y��=�;���gJJ�Z��~�����(d�E���������\��3.N�K�vY��������ER��U"m����s��4�Sg�D���u���� �ޑØ�v8��O���u���΋�3[��E�M8H܇ś��u�<ؗ�;�޺�-v~qn���{]��"���Ծi�Ѵ�u4�{y|���7�sCZa>5�<xW�B��8{I��i�3�ɰ��f����PK gO�D]+2y����I8QV�Ii����}vW<8�/yi�6~O���=+�鯻gi_v����b(4b��0�-
��_�:RHI��1�m�~���������x�Y������)K"�)�I�P�F���$��߿{�j�N�Z���o�[��X����Pn��4Z��U�-��:�X2}Ed��)/˛�~-�Z�D�0F4���AiFw�0�LGiԳ�w���鶺|`D������3kX_ԕqJ\�"���dxd#���%[�������g9D�3��|��Df�U��_?Z4*�[׾ꖺ���i��${W��E6N�/�ۇ���uu��(W�NJ��(��mHVJ���1�nHA?���n��Җ,���X��	�8C�|h41:��|m��U�W�%ɹG�H�S̓����4-rp��2Z��cF�����Z���z�i:�2̈K�9D�>+�FL��̱NS��k.3��B
I|\�����H��񟷈�鍷F4j�����_J TSQ)�]�&T �� o�兄�T]�X��AF���Jŋ�w��b�`a#3���H�X �)�o�FIr�)
?���#�յ�Z_��r���(T��� �C6L}ˍ�J<M�Z��R�Q���
_6��B�a�G�+.���n5l��am��i��������Ѡu�;���y`�b�t!h��� ��a����f�����:�n2��6�O�%@W׮4^a)����}�t�ڟڣf���I\:�e�UsV.H��E��Z��������\�9i@J��1rX�GZ��ҬN+��ZJ�;����Y/e����~�)�	���Wb���cI:"#4:]�K0	po�yΩ@��@�4O>�j}]�7��BD�Oe7�l� �O�Y`dQ3]/�{�]��7�8F��w���	��7�U��W8+���X��>�ɵ)��8wW6K���3�[�+���1ϭ��#�X��'T��M*#��e󅅃�@4&A�q��6��ӣ����<&1��(��c-����r`/�j*� k�-Gm����:ڇ�)�'j����/3�5���h��>�m�ׯEc3$a�vΫᓌ�h�q`Y����kQqS6�)c �~����E8�!v.���R$�lֿQ���ه��/�ص�h�D�j������iR�6J�̚꾸�su�OJ�!����y��A��gZ��nQ�X�{\�SB�#>�����q�n�c��g7vX��9��߸����+!���E��{Ҁ�O��I������������M�H��jL�������SJ���F(:����17p\ѩ#6@`���>�n	Q���\{~�Y�ѵv�cipM`Ɯ�%�[�BX�����
��?���0�k�X�c��&~�d8�9� �9���!H�ɢ|��H_���I49�thA=C4,gn�l��A����{rt���=ˌ�J�?��I�O�6M��+P�y��+p�Fx�&�a���t�ibEX�j=kZ�M�J�R��Q�ޢx^��>�3�b���95{���B4�ǈ&`H5�M�;纏q���~�hk�2��� �I׉�@T�߿_�������5H�%T�����B|�p�tɣ�����`J6#
#��%/KИQ<��K,��a=>��#�Y���o�ѨMsN�-�B���n3�߅C:�$��Do=�ų�&��&���'�Rk�Q	G�2;Dg�Q�|�:�h���� y��p5�	g?���oY��L-��	W���áVXb{7��I���=�zX�g�֢S�;�棋oc=�5H���0^T?�b��X
W�����'�ґ;y��č�����5�(�l���58f�����3���Raλ�j�%	�a���XI�fc��X�x��,>��ihx�}LQ9F�;d�|}�*q�#�gE&�I?ɔ6��~~�\�m$A#�D�i#���Ȉ���ȨV)5��H�T���,�գ,��%��"κx�'v��"n~7�N�nð�FǄQo5U��B���Z쳶����M��(4^A��S7�	s8W��W��o���HE�	_S�u�����`�l�VVl8lr(��5�^�C�jd�ihV��&���л����
�m���	�"��m����8p-U43B���[���,��A��x�	��dWX$��ɱ"���j�l]�@�%�0��)[M���p���~��ƻ����֕���:;�T�J%�.";cq� Vc���}X��V�C5KDB)
Dd���<�u?Κ�K�N�f`���1�Y*NĘ���9������UT9�Q�}UѸ%�'�a�Ԧ�"����
��M�g���.�2�(~`�C�m��v�9+u7�-$�����X�%nov,�>����z|"�)��&Q��Ƀ_c�!G0k��~'I�5-�kI�0��0}|��|��󶍍y�,� `U6�r�wC,gP���h�����y�$2�DT�J�m�Ź����cP*�Z{f+����'��x� r�vFHU���C���C���9q�MZ�=���,�]ʛ�o"W��u�������[Q�Us�{Y3Z���`ׄ��uB� ��y�"�����841ѱ�X��Z��a�H���V8r����i�wY����`�k9��) ��5µJ���{�#��7��������?��\)������LC��j`��f ������%|����pv�:��s�UTC��בbӲMV�XW�Y�)������U�P�3|�;ز�MC������Xp�S �CSJ۰`��G�����`��͡�)�Q���,�Q(<W��+�X�M��(�8�*�(���xh'b������})��nY���!UT!��FԖ�j��7�\�w��pPb������ ���C�ޑA�����´KRs��K�@Tĉ����1U���Ｐג!�Za1�~��y1^�<�C ��ǟ~J�^�8Z��6n�@.��(`���V���߈{aN��>Z�]_��SCy>��}R��GB狫�_9n��!{��הs|K6Y�I��{��*���:�\HCSWvζO���a�MU�J[��#�K��	�I����g�}�����&۸��ԩ�fܟl�Y�����G��$�i �EPU���m�󶰏`�O�S�]���w��)������eb��d3�j�;PR�ޕ_��k�5QT59?	��|\]���J�C���p��cm7��W$��lJko�-R����8O|�lJN���
�Y��?�������b�ܖ�h2<vޝ�I'��yӶ��a���j��p�W:�Y�E�1sY�*b�XƠ�yI����+��c*��<"%olr�x���r1��K\Dm���$���Z
�����|r�nQy��!:��E��X�Kfٸ��<�ج�+��:�V��'a�) [��7_S���F7	I+UV5?�;!����Zı��W�Q�!����ȞK��]��_]3@"(l��i��	+"�X���,l׳� "R�3#.TWmmY�ױ�OXMh�5j~o��x�!���>��M�&�>l��T�����iמ1I��|�6k��t�z�m���lI�B�a|PZ>^�3ۻ�>c��|�"%�a����#�*0��b6 PI
Դl?�f�mVp0z{�`�~���2�)�8�k������iB�V#��c~m����*����e��]��qT���4���<4;gU\k��f%�%����0������ �3k�X������Hq���#0�g�FVc�Z#�3�$�*�#�3��Wr[ M�S���(�qJ�8������{g�>��MSo�%�z�o7�<o�I��︑-�G���-F�	�MmeHe�j�U[y�l!L�G��v0ݰ�.A*����@��mC�K���w����`��t�G�+j�61,�AK-wqȰ�~�����'\�x���(���l���'�*u�S���I�\K���I�Wꖠ��sr�wȤ§G��p:�]ﺱ�o)]�ma�Ǌ�G�8���#�Cw����{K���8�5���� I?����S�5E�Q`jRR��;��N�H���g��W�DHm�6�����M�����M�^�ɲ����z�2�d4K��r�(:N���x�7G(��v��*�
����Z#�_�{��*%|�sV�u�9�� ��!�����9i�������Qݡ�"�Q�b�6�{�6d�V�B1ZRC��ep�=�#v��z�P�z.�t��h|�����u �4.�h�(_|��s�W��?zH��l�����KV�'P��bS���m�ҷY�hsC"�%��sc�ti����y�YC�ćƈ�ŇT�����ͺDa����GU�gF����bL��1*����H��j��!��C�����~��M��1R
)�@39�9�,*׾-*��S��%�}:�uȯ.5�9����m�d�ם���`�|V0�ѣ�ǆY<rE�Ml�p~�4� �꣪��!
�x�!	�����7? �ً�2�Ͷ3��[������7�����
S�uFf�S�7V|B�\����m��ʐ`��,U `dwWh�=K@G[0�hu��^f� 8���6=R;3Dhx��'c@�	��]2Ua��� E�N�� ����@�)�<*��x=
G��ĩ�(��@Ӕ0l�o_��^ߔ�8��3��B,�	ң��t�Ā�_��.�TI]��U��AR0���isȈ��6��c�գ���?�|n���󈴭#�6�"d0բe�[�h�����Ы�&�/J�p��f���hc�����1��4��}i�0�q������A�(̬�7������TĪg<aS�ۈ^O���z�*6���;�Do\����6��=;1l&���,%�!��W����ɢv/*Q����7Y��\>n}��!��DFa��^�z��1B�b ��} �q5���6g�9w]\�郭���0�Z�����Rl���?'wxS�]��\������5\�9�u]oonܐR	�k���v@�_x!d�(��}�'�ˎ<�xu��L�d��
u�X'c?�i�0S��VE?1�RPPCF�݉�FOb�������~�߇s�����s�����{rA�!�)E޽gy�\IÊϧ�2���ZDH��4����vސ����4���c�qc��u�ڦ:8�8��~]q�uV�nP���aːj
)���#v�=��o�F�3�p�# ��.Y�% эIUOJeL�f���ː�EL��R�>jn?��4���X�?���ǻ�p7�.F@�P��&0�F��B�*T�ߚ���`���W����xs����Ӎ�,)��y"'`
7���-XBl�BɽGcχ�e�$emX<,]s8i��߿�Ap27���ԓK��*��˘
��H�['�g*e�D��T�6����]� �iJy�B�;�*tKF�˜\�R��w\��6:����$�v�ǭ4.�׽�Q��7�&��DKC$�ȟ}�W�1����	1꒩�g��ӝW=�fwh\
ۆ[7�ZΡ��k��V<Gq�ٚ��G��	���k3���D��Ϥ���y$�"%��/Bip;7�9v��;��H���㝮�wx��t�=6�����w(���=ԋ��%��
��9�٦uc��Z�� �Q-��N����>_�������N�3�EB.�%����M�"����߿cM?��f:X�P��"�J�5Q�H��&��jOTTx{C��6�bB��� �^8��=hc^�i=�O	��sԶ�WmD� �]�q��L}4uR�R�'Uc�)ܮ�z�y�����0(����`1�s}/D#�$�ñ��,����Ԫ�r����Abˈ�S�Č��X>F���9��A�� �[a�U�OF�gK���H�9�������Z%�R�f[�M�5q��Z��O�h�m��ڽ��0�6��Z�zا$�W���T�
;��u���
XE��%��auS���c��燑B6(�a��h�a `#��!껢���@:��d�N�q�������~oYC �A]q���E��k��/����OA�E슋�:��mlLe4��������&}\���=�>f�s��"o\�YjP�P�U��SbO8�M�h�����G̜ A"AK���iJ����Pz�>�D��M칥=���?��7��c�����9tCQ�=��%�dQD֛�)3��/,%���=<�q�&�%s�"�[�̔o2���N�$�,���t*Z�9��9:����i�y3�q�y��~x8�CG��D���b;�yg���]�M���i5�[]'����~�.t���$���^}����1as=.�1!g��Dڐ��_�`E?+��	q_�=�_F� ��Q~\�z�I����P���FE�٢ \��M���zM�홌��_�Ck��N��K7��/�����$��Έؼ��sv�ᵎׁ��'��y]�ជݸҥ�q\���4>��q)���&葺����*{�v�&w����k{8BY��s�2�bWw��^�W�BBA�2&s�r,No�y�D&�P0dF�O��,\Q��^�'\�u�{
�c��Xq��*�;Up`�F�Y�t���PJ�0_vN����{���b�\Wֳ�MPYա��'[���)��|Ύu��ba[F��s>103K�a�Xt�6���1��$օ;'%�#	�PN�ϣ)�\.'Sg���&�7�s�pBmH�0	�S!�6��Re����
7���/M5�.6+�	�A�
ԖhH�����7��f��>fL�av��t���u��u2�aUǛ�X�\:y�t*3����������~o<QPJ�ۈv�#|D��o�;U�|��'"R�Q�P�hkxb ��羿���~i�����9e)�4�8P��/���Y x�S�3�h�0̈JŨ`�Qֲ�9ED�e""}�^r�0JV�p�9B��S0�|����s&������[ߏ�&�|�@�$��8#
c������+�JfM	�$��r���TR���4n}4M�TT:��0w�(�%�6��pWP�P�������v������;��>�=}tMb�y��;��GJ��^~��֣iސ==�k�	���5FZŢ�ʧ��Վ��_�Bը��8�R)D��ܥ��E.�Ns���"EHIX��2GX�y=�Cu�
���j���UŴ�H�6;�u8��b�i����ʠ+2� ˻+
%D*:��a�/67�uy��D-F1A��J|աg���N���ɡ��9Mq�¹���cgѪ��^ฅ�E�j�
Jͧ��-�V�Xa/q1�RlB.�{��_��X���ͩ@��5jl��ã�
��������$غ�j�Cg��q��)�|��(��!.��#*���8��2���ǲ�Hk�>,����E��b:-�/w�Ւ]��,gjx4"i?�g:h<���p��9��1ޤ9A�?X'���8����|O�6��4"P�c�Hgfs���X�3�P�a�����
��?J�SQ��s������{��|<D}�j�}:�P��r�6�$���Zim1A�� �h�Y����LJ���0�n�}C�	ָ_m�ܓ;�ٙ$J�&k>�:$x2���󣖥��U-���S��Wx�[�z�wXUf!��)	n���"��/v�C�1���4__g24�.�|��1Bp)�Pp�EhyJ��n�b��-�c.����&�uq��v��)�g�A;� ��:M8��}y�F�H�8�䃍�Ib("�ӣ����>'iO�u�a㷾�,Es�D)���t�'OUL��Y�Pr�=�}ai�m���X����oo�FrcR2|�`� ��(b)��;a��w������B��k�磳���R��"���]'^v��X�0.�����\/�x��K?�1\7 ��iH��3f�]@<Ț��Q� P�W֔�)����gqȫ�ۀ��ڥ�YcY ��O�A7�~��,1f&o�I8���pu9F�׾U���0��X��C�:�R7�� �p�ܮ��=�ِ���1t83F~�o����Dۯ�x���ch3�WD�H7�B3��f��:np�n�b7]|��]���jS^��M�g;�=*'�8��oKH�Q�:\K�bэ=���.�QJ���ztC)i���F[is��h(�H�V�w���ȓ�2�SP4k-0����֣��V����W嫯��4Y�6"�GO�mF9�8����3R^lVu=1U��,h�b=F_�>.59_XdE�����0��.3��fX_�x�<��Χ�R����zK�pm��,�W��Ӝ������Nmj%0�z(9���:�n��]'RS�Y_��qE�9$���e����=�ɢ!��hWT�ii� e\��۞�M���6�/�u�T-��=���gá�EU��"ņ��+b#J��ڻ!xFT{VԵibuX�_M{�$J��� ���\o�m}�Ѡ�!����_F����ώs#x�f�?a�a|2,�x���$�c?c?iԈ�>U��پ�!�N�ә�����������_�`���ć#'w�S
����zݵ�hd�)"�:�櫔�(�"k�Yt8!��&)k��j@�T�Dzҽ��xX�[�Q��!�F� ��?d�Do�h�@c�s�U�m��ۊmD�GMo��ɿ��FF�{�ٹ�DJ�0�\}߆h+>�QFaY.�zY�hn���l��S�M8�&'�;W�O��
͖�q1�>��p$�J��UOŜ�MN��
�u5\�w5�����;�X �dMS/r���R�٣V���xtm\ҶMϾ0�5ޣ�-->�m��.�wo���D��3��/� C�
7�戀�3��*�~PL���x4��J�QVi�^����mF6����y��Ce�65?��y۾�rx��� 9nO��3��9�0�T[�^s-3�3�	-U��""��6�ϤHI*��Y�f��Á8��ό�~�]��s���
��<[}�䐁��\��)�;-�����3�)nT�1ҕ��|�p'cJq�'�,�Nq��v�̻fs�dHe��O����͙��	>Q��m"�Ń��!��eʠ�m�)�Ti�-�q����nM^QM(��A_d���4i&������ņ����7��l�����3Vh7�����sZL���)����֙��}�bS��|����uF�z%UJ0��Wz���s��B�NU�,��ܣ�HPBX��֩单Q��j�������-�Ьl�}�����읾�qƇ��Ba�:�/6��zk��6��@e�V&:D�R���y̡.��*ǀBLJm��3��S�px������x�5�+�7��=Wx�R#eT�&�7�wEeë�w��B7n^DoF�[,:"���I���*��Fs|kd�~�u�~g�[���J���,-��֛7�>9-[e)�v�3lTWz'Ƕ1(D{�Eܱ��2��Ǹ�u�B���z�>�ds~�Ս��ѓ�fz�m�C�����_��"�1��z����(*U^��uY�!���t}�j6�p)�M4��^����T���-!�e������^��9�sKx��\]�TMv}n/�^���;'�F�W�$���T�u#��BI��M�]�==�v�
5�VUHPt8.��:e��f\���+C%�#�I�]����w���!I�ΑE���%�O��_|����W��OjҐf�����4�H*X��s]E�#" D¯����/�o^ݼ0j�����X�E䅆�!�񔔩�Qb��xf�������S�y�&��:o�;�S#31UT�
?��`}�����{�Z䆩���LD��c(������}�z��ʴ,���ept��T�Y%�Rx�lK�ሓw׭�Nc͡W������d�W�x��X�� Ԣ����w ���*���Y+T�j�;��������S#[4FE�D�q-һ2�S<a�t>Ť� ���y�q���ZM�h$����2Z5cA������5;LR���@���(�j�v�z]��:�Q�d���"�MD�ܘV�PvI�u:�N=�T������S�a/^U��]��PO�Dd��mR�X"В��i2��yY2��>p����\Вv52E\7��)6��7�~kt���֮ׅJ�/��HZ�$�w�."Q��de��C���P�WO�|�-~�����=�I�#��L$P�ը��R=�����ܷ�w\1Ӳ
@�7���#P3�偬���* 32���?�Ǩ��i<v��F��b!ߒ�Z��c���M�*x�ar1�I���)��m�
���1�s��[�Hݳ��K�p�O�L�����*X��'m�tu0bbk4vT|_`�@�K� T���g��$�p8���}��=����㗨����wl=��?��<>]AA�C?��qo���qqc�Yj�1�h����eCt�]�0"�U燤=�j�f�h����l�`M�E£��D���nӜ-�mg��W����~>��!�#rP���R)�������r>�T'� �눴�����[T�yn�]'������3�8E�zw\V��ղ0��4_��Q~��H�C���#��#9h^�iA���c���8e"�L�Qiske�-�1����:z��$*�*���v�.�IbU�!?��3��f�ty(�{OE�aX�̂P�v��v�}��F���m��wv�W�U׀0�eUs��n��xx�i��|\��@d����i��u(�B>�7ǈ�GNj�y�ff2v��Eu�)�� �o�Q�!hd>�Ǖ�[������YZ�-�-T2(؋d>$�JA4�k,J�c�G$!�9&S�RAH�������	9�CrI���1�WP^�R#1����|���?N�ёCl{��-dU�����FFo_�����RH�p�W��8e�������hum��#G�����U�!�8:�X$�Y9� lsj�<Ys�q�)���Q!�g�ɇ�4��uH諗��>sϫߍH��Y��T���T�?s�����i��a�����UuwYU���}���5����#R?�lB�V��^��\���V���V����M ��T,���È�����Q��ǈ����%��%��U���8��jT�H�a#�r��u>=�$ڏ7�r���>/Af7u��hׁt�\Q��>Lɨ�D��,�w��晕ToxE����~иvT��)�?u �Z4�/Tп~�hc�����LL���}b�>@��C���/�\G �껁� iF9%�: ����<�h�]E����~�xh�*J�ǲ�4O6�"�e+�Z�ʦƲ$O4(E�L��d �/)h<��N��pL��YY�S���_��R�-��mXpf�fn�\q@���|���(�s�$�(Z]@a��D�C�����[����U~N��b�~nE�m�]5�XL-��h�4�B;S�ք�1���a���5:����1���S�5�k�(nWѓA���F��}1E�tY��������e���-M7���j��������Q�_����hP����E���G��z5��n뻽%IނN��gF�x��)G�z����
8hU�ӧω]R�L��sv\��]��F�>�C(.�@8��	�+RT��T������wR���9�	0J�g�������z�~���v�cRV@Q436�� �����>1����x<�q���?伣7aX�����SUܡ���q�A�v�V"�9M��4}w����v���	���z`��F&������,zJ�8 �0�������&mE]Y��9��VT#��j{��扊�]_c�f���"o�RCa�sk$y��{��H
Vb�^\a�2�H�7��:R\�H![�]�F�5bw�J5�c|��X�Ε_��֚�s���y���$V�,�g�;�Q5S�hlD�Iu��r��	�mw$.���;�o�:�c�0O.<-q��]�طǏ�jYDwzmH_㺿1}�1��ڭ���!�[�7.���]2.X�E<�8�Z��.��>�-<l���v���z9o��~���|��.@��h�P���xy���ltN2�?d�u<�o}���r
��Ym�QQ����
�)��m�Q['`��}���F=ޥ��Dt�*r�,;"'�����>)�����UU>#L|�6X<�>���x1�V#��.�3#��`{�i�M��p8v��9(�+���|](�%Lxw�DV����1�!j>`q��]�Mv<5��|n���~��{=�2Xm��{w��=4��	�EN�Q�x�q�	�NSCxY���&�����fi"�,�6\Z��-����]c�~������Bvhx���&�sp1���|���b�زn*��Q],�og�Dy��6O�75f�T��ɐ.M�!�xv;i��L��+9z��,C���P����r����*�����x�+�WH�ݪg�#
�|�ɿ�|{Dn!��;4z�.��9mc�M5�յ����G��O���{�_Do�bW��X���N��������X/ߟ����pJ�
��S�)<?62�X=�s�mre��Y8 S�=��t��8�����;bL�.[%�H�6�9/|63`��@������9x�0KG��*����Yl�%6�vд�b�܀14���if���a�	�	�)��������y�]qX��b��Z�_ "W��
qq�m�k�4
Ǽ���ߍ�_ݥ��Z)����ف�E�&tネÍȭipY5�G�� �K��R��n��0�2�oVt��>r�q���3V#r�	����Ρx���o�b?ڡn�a�6(�I�8g�kպ;skY3�] �G����Q���u�K�,ΕQ���3��?�0I_2�v����X�L�ʃX��н�u@�u�m��ZԐ~��n���g$M�W{l�ǆ>�b~�s��j'���1n9��3Z0��)6I㕶e�/���% }�F�&Fa�į��$�����FI����੩Pyҥf�Ħ��s8����)����#�r4�U�$B���!�.W8��W|���m�{-I����)�F2&lk��/�w�Jf�b\0�W�OnTr���Et���������o��a*;�)�f��r�d��d^��}]�����[}��/�jj��(�Z�jH��sJ׭o�(z�kv�c����p��LM���hU�O������
���^�;Ӝ4)�y��#Hj;G���eyz��@���Χs�l���t �λ�<�S�����Mp�{'��Jk�.��s�J	��'ơ梅�) 9c_F��
E9N���_YB_X�����X���������w�?v���@�����ҙ�9;��j'4&�Τ�NO�Vc�P��V�p�l��<����]V|m�L�rO>�.�����J���Ѧ��p��>�J���s:j&�S_K���R��6�~.��X�)R� ��~v^��O��yR�2.9��V*�B�����:�ބr<"j|���Q�n7&-�YEG�Ƙc���dѨ$�5K��P�v�v��90*
x@cVއ�=�ѝ:�.�B�h���J�`=̈T|H�z�z(߬�]d9�&%
�ٶ�)\Q*Ν΁�Ӝ����i�~��l7{�w����4�=���/��Ic�`�#R��߾{�Њ#�V?�i5-�uQ��QV�#16��}�N�^3�e:�`�[F��BdƎ�|!E���g!S\����l|�p�PC�(.����,��B�:�YQ�M{� [ř�ې΂�Ᾱ�V�
�f�_^Ā��n.&�W�I�U�V�e�^E�՘Vkx]�����!k��b�v�ՉQ1a*-�ߤ�J��>M���IX����Ӽ�p�!n�X���7�I
��n�G9�B<��;�Ǯx�Bp2U���3��Y|��3��}�Z��]����i��Yj;�;
��C��S*s��ta��XN�H�US3(EG*�;b�Cr[�@q�)��6�]S,1�oۦi��s;F����a��i`>��ؘ�/ˉ�ա��f��>U�n��Ͼ�-V�����i8���=y����u������Ģ�Ѻ��6J^a�U��c��/��f|��h//x��|�p7�@�S��J֊&y�2���PS�0��b2q�OO҉u���eM��3��k�*j"ts ��5�9IU���^3�"��v�d&Uz��w��a�y^�������s݉r��h�ZT���oݍ�,%6fh�.ၼ#��{��Al�E��'�Anc��l��φX
 �,�̤����u���^S�5�]���@�����P�y)k�[e�_ť8h���`}fOxwƎ�9r����IL	�;�}���P_I7Y�����c��q�e�ϯ�ε��r��G�G�Y��dX b×�����XZl�Q�ݝZ�u��8�0��H}���5&:IH!$����	�� ��������*��:�����>n�*)��w��4i�.��]'cU~�
���˄�\������0�"a��WD�l�M���he���0��-1>���H�4&n Qt��t���Fƛ��uӰ��s�����rО��(%.|�����85ː�A��J�S�lp���Ug��f���N�	N�&j���*;PwO�I�T�w�F��fw؍2)�� �����_��vт���Ye<�!x-V�y��۞=��l<���_�1n��Ykt4��p�X�l��.�����̍P�:#j'dPa�v] ��rM���֠* ujo��U��UqR�]Y��n&w�r�c�y����RT�Wva<<�������!
���������FI�ƭ�&Up���fFq'�&�^~��p;��}V;gr�UCU�}Fۤ�\8e��0����e*��U��3��c�۶�"Ӂn�2��(O8�û��É?�=�#|���>��5��a�(��sF�~����+�:h����x�g�Lp��ºĢ���>�s����U���O]�T�*��޸����(gE�OyOQ��U%&쟣& DƤ�J��%�f7�xp���Z���4[�F�V���&y�!e�e�u�A���#0ȱ5����c]c����}�`�m������sG��D��g6�Cm�6v.��L���&
�`���x���嶜�����4��kE�/��{:��a��56�J�0ǳ �۠�A�
�E�o����Л�7���^81�����1�����`@ciJ]�����NI�v(��I�w�=W�������ujoS�w0�5M���������6"n�j��k`��̘�_.$���zӑ�з�B�S�� 9��)]7�bwi`�bn��I�d��k^_�s���V�������9 �'id�Ԟ@{_��k�撞�S١Q��nْ���:up�Yq�X��g�&�OK�X��P�{�eԍ�h޴b?�U9��l�0�����갔�z��9t��}���P��lN�4zU�T�������F��8W���p�x�Ð��A���Fذւ���eո^b�3�_��4��V4U��;�G�2��`�q�*���N����Ya�����r����{ŷ�,�*Wt1����(��o���(�I�#1"2%E����i�X����q��>�s#~�s�fv�l��f��`>w�EČs؏�~���k�YhS���V.�1�L�jZC|�r����Mͺ�V��J8_����e�
��%0�����3�2���LgGG
"���89+-px+?1j|j��U�������{��v�+�1�_E�a[*�5G� J���/��� ����ۨ��e�=��
)�`���!D���aq;�7+����2O�Gd�X��F{��?,��/�{;ѓ�J|P�����d4r�M��oR�z��w��7���E����n�\gqCa>4i隅����ne�~V!���%��|7ϝG$���y��ޏ��]���zz��,��a{΅���T�r�, �P�z�Q���� ��ᔾ/�"s�Ύ,t�0uQ�k�2��J�oqT��+�����Ο>�b�<ާ�@����L͌��X�b-�3�0���23��Lu_��N8�ԵM�Y�ۋ�����8�DE���	�>�j��"*m�?�q��|��_�:����E4H����:�������G�#B��t�,oc`��l�����1�|x�!�B�P�Ez���u�Ϲ�X���.n�����rX�'�J��ʡ��5|w��k���loC��6Sl��I�"��0���q�nh�a�����RT����3�+���__S��cbf6n�z���p<v �v{�5���.��	��%ػ�z�0���>K�b3������u�Yo�4[k/L��`�Vq�X`p�[�m���%�Q���}��@A�pY�Fe�
N�}�i~|�f.i/|���9-n6�%�)`/D�ls��&�o��
o�ڠ����wa$?}�T>m{��ki��������'I����=�S��:�RQ8�~(��ܧX�)+��	t`]|�ϥ��w{r��_ԣ�Fo������p�
�1�Q�8���o�7a@�//n��]G������I�����) O��e��F�i=s�|Q�Z�)��X�kB�+���G��z�W�dKf��3��P�~:,7��X�䩟���C�����a���ka^>�&��K���iH6ֽR�v�3၊�;��L����8�dE�7�~�X9�]w� �h�`�!�����]�8C_g%�bΟ�.E��kr����#�QY�@��E�H�Y��� ;s�DQd��`�)>��`"R�}��)�g����!��2#.�X��a]I5{HC�C�,��/�(0�:�&��Ո̾n���f��`�R�r�p�`|>qO8���)�K�j��/�K�hg�xK�H�u9_Ȅzg&_�u���J@C\�^mЦ�����n����������6��E��l�z�ܕ��.?��c����?�g<��PB8SлD���ě/U�$x��̶/}�0�!GK��7�Vjb;40Q���Q|�r������� N���&?s���5&+|��sf�9%��ׁ����P~���X��X�����]�N�g41)�E�t���uߗ����"l�������KZ��i�U��X�&"����]���T�;WK�n�G�8ͬ��2�22%æ���GFQ	�8h��E}���؄�-�$�����H��>����T����)������I������^J;҃�7��� |��t�TBG��
<N=<%�Ņ���ValA'��O�:�)��uF!M�P�:�U�����03;�� 
�FH�A<��fQr�Ŗg�]չ��#E�È"����+|����
����((i#�����T2����H��Ut��ɐ<FR]%Kv���{�����wUǲ�#	J�cW��&`�\XC=I _�����x�F!΃뾗��e"����cjCD�E!)�흨%l6O�@���i��b����=����v;�(&ng�$�~��b��!q9+���3���q�]�3�M:�5���FnX�����id����#�^�B�z|րlЌ�}�q/�zM� �Ѯ2d��,��`޿kd+��P����?�w��������Q�����ĕ�0�Pj�QC:z���q"(�� i�;���=�>�L���x^�qXp����ύ*�-E^�8����+9I����i�<�I6��V�%��)��s������	�;n�8�C�̩�ʡ\j��x}Q��l+�Y�of��#�+_��㔅�.�r��x�n�+Hۭ�c}�l���?IpeR'���UA���O���Kd�f�3�(REA����0��M�`T,��͈o�֕p��ƂEP���/�l�y&���k�������Ȼ.g��{�Í渏L�/lB�����_��r�RD��hH�E�1��Ǔ�Mx��y֥��4���S�:0`=�9�f��wfY��Q�<"�h*��!�s9*0�4;��� ��5���/g���N�`C�.��Ҙb��o���Y�������^{�.��Q�Qj!3�D��h7�l��Z �8�p�����Ok���1�W/=נ|�w��m�i� �IU���lF�:Ԩ4�N�E{��S"n���@s������HE~ݾ��A�G܄[�������q��4�K���D/~'��P�׬�ë��E� �Kz��}j���SL�L}UG8��-��I�|�ᨊ���j���_�K��_D�A��C�����?Ʀ�
�f(��l�+e������Et�Ӊ�g�����	���4�ќ�q	0�<l��m���8|_>���?�%�����]n�ٸ2�k��q��	��RG���Ѿf�x�C��)B�"��ʉ�6���!V6�XV�wF�KK�r��^�ws*a��c�
���pDN)?��s���?G ���oL���nBo����Q|b\�ˉ�XOo�t 6D$-
��I��G��n8��	#�$:��Ӿ�����@)�Ѣ�Gq{�P�{�S���sCW������sF�4�k|��� ^���B؋�r!����?l�{NF�y��k0c��� fW�z^ӛ^����M�jO�"�uW�����SU�Tp��o�EjSXY#vG�z72��8ȰEeK9oF��t�����n��cv$��7�s=�`Hl��$��b��U���B�w]ġ����+� ���	�'.<{i��z�JŃ�Kx��ݠ��T�!ժ>$�G�Ѐ{>�7�i'c�|S⫋�V�"(
l�M���>���n����>X�1p�QuE� �x�yI�N���� �y�V+�@�R�3��EX/�.sM�c���'���#k|(b
�v��ḚJ�UZK�k<�]]V&
��w$�� �zS��a�7�+U�T��J���p��g�u�e-�V!)�׹F�cFSYz?��ݴrY�"݀�R�v��g��v.R�H�\Ea����W�c�ָ_*=�g�0r>�G�X��m�0E�cdE����Z�+:����\�$�W��?g�m�K4���ځ�k�5����7/�<Ґ�m��b�ki�����	�'��1�6-à���V�1��`�_n^�R �EL��xJl�7��)��$�����&�u �������E������>���8�� On^��D�oZ�_��9B��Ak�_�e����!���|6""��d���g|�{�	��@�>��D��%��xE�~x�Plڢ%T�]���*������=����}~�EW����D��.�˔stb/�3��e���GyB�a6���Q�̠�.{�Tv��k��Q�Y��%ӮM�h�&��]I�67��v(�C�;��Z�(����ݩ ����mYa~1l\�N���\��E��a/Z�]Ϋ2���ꭃws����0l�����\ؽh#b�`�5��[�Ȇ��#D��b�F���M�M�/� Fa�A8��ѻ�F��?�vlN� ��J��O��0�����w׆����#lGͥ7�0[�i����M�o�%���-��Q���/�9����,���FzG����&v�t��oԆԞ���F?y���M�:�(��z��6��öؓ�z;N\���u�C	#v������?�����א�c�TM<�1f���pU*��;�O�|�<�@���ys��IA�Ɛ�#u�j�f�G�o�L@��xH�.���;���S���Q������ɝ�x>~����XGT�q/HGQh�!6�4"7:�ϱo\�u���k�k����J�P#A��E����m� �-����]�}��{�5ۜ@��\K[���J��{�^c��sT�)*�n>d5��M�Bլ^��c^R�����)eͬ�s�Q9�#�y�£����RY�2�q�LTݫ�3��V��  �s�>��F'���;�1&�*ru��L�4;rP��J���H��"|�48J� �b[�k�	�Q�|g�m���Z�PȄ��1�,5K�!�SDe<�[��ԃ�*xk��Q�2-��牎No"*U;gz��]�Op ����A͠BQ��U%>��y���pJ���o��X��$x{�2��a9G�Dt��C�E�WАަ6�F_���_�%x���o��?���
%`S|��q�� !{����ZӞ��pЁk�(�j&�ć͐���Р���+)L�*
xN;
{6��dq?��_
ǳ|�h2|4����Ѕv����O?��d\�v�!B7r3t�!�������4��r���3�qG����;��k�f*2<1{��y����`i[4�b��V�
�G�{�(�t�޲EU�5�,��ro�T�j4�b!���	��4��`i#Rub!�2}��|N6��||���ޡh��Jt��b2��"o�蠣���T*�����!Ea�T�=W��`���h����j
�^D�O���x��<�>G��p潮��r{�:%��yZ���k����� �F����H-v䂓4G�m���s�*�������'g� �B�.i�&Z���2��r��渉H�/����ɘb3,ul2^�I���V!{%D�` ���9{�M�N�^�Ȅ)!�)�?\Uཐ�춛�� ���q��s#�؀��eꆈ�#�EtD���)�+�"��*��o@4�Q �1G1�aՑ���d�Q��Rm��C�z�9�_���(<�ȳC�����!�@�"`��#ٷ�$�ً�S;R.S`�������$�q'^�slDA_��f�>�3�X��3u��?��|�E�4�L���xVq����0 x��R�NfY�����4��|f��Z�՗)4;��<�@��1#�q�h�>=1"1���ﮰ�0�F�ј��,>�H78�����.��Ql�m�����u����J=�aa�8��.3\r�i��2����b��j֔�a��e�6l3�(�|..�������(�y�4A��U�g���;2�m��ʾ���i1mH_KEU0@6��^̳�5ђ�
!��Ε�˙)ґe�^)۸f��T\F��#E�2��/�����9cm�͕�����?dDk~�!�i�w�P��}�/Yr�R	���0$���t�%6r�QnlP�9��e7��F:m��_J#����F�Bz�50�l�a�I��:��*J�G��B�}}�#��n,�ǉ�_a䤤ONfm�ͷl� l��(����f�c�O|��JLǞ��C����mT亸��5�����
,���(8����aHmX���Y���s:죰a8��L�\�&�{#�[��P�ʽ3�p����<) �h�q��.�h���{����N8��(��(8���M졯�ti���kvR��QIV�*��ݠ�u]���D@t"�}g�"Y�!2l��q��2(Ws��B7�he��!��m�`k�Q�%�����Gп4z��S���dH�ڽ��d�����fa�.�Iy�]kD[>Z�S�I)�GCU�A2=����tV�������g�dc����?����?���9ӀPOza�!Da��D}���JoI��=��;j��;��^9$�\�Ke\9z�Cј=6���1���C�5�
:�V.��^���ǿ!\AR�s�.N�=����x���H=s�$�����-f�G��;9�!�KAad��ܫ[�>Ԫ�0��?��׍�F�T4"����ȢY�I=�v�ϭ�״�N��#�����ݶ�����_��_�l:9��6�|�ݐ��!�֡��\�E�ֳ�FBN�2��Y������
G!��q���JY�]�P�^�7=뀛�ݫ��4�2'*g�i���R�y����(C���BQ!���c�yD;9��B��eI��Vڟc�gD�H�5�.��>G62��������5��rD�ۭYl㵘�?+@��]I����E��%���Q|�}F�-��m�.Q�����OGCZ~׈:��W0s�7�-,�-x�5#d�[Z�����$�k���]{!S/~Kϸ��uN�������h���D�G��TՐ�'��,K�ZS�I��}���S��KL�ޯ�e���a��a����(\G+��tDl��h�z 8�bWT=�R�Z�����z���r�����Ǝ�h���#��&��H����F���[j��$CȗSزK�W�*���l�_�F���D�%��F��F��ؕFM(��cT�}�.���ؓ���U�'6���t�
��}K��\�H'Y�m���k*k����Z�m��m��{�|iy���ಋ4/�Yc/�.&LU�X����l�y^��&+y�17E,���ܘa=���m�#D�C�jB8��LxW���\x��Z��I�������<:�m�>���H�2\�D���	�M�Emb���:尵��| ��'\���D�g�j�s�ܞ�3MU�ؑ�EI��3"�����9��ѣ!Y���AV���Ї�.�_��n�^.�Z�(v)]F����u�sSv�X�
�<�T���u}|�Ȗ!��[͚:)��zEv T2j</u�O}ya���х����Rq<�+*���P)�&�Gl��{%�U�T�-7~IC�H��Ydp�����q��+oo1��#P9Nd�1I�X�RGQA+��l��=�9T)@.p`� Z�y�=]�q�u퓦gV��f��QxP��jpDI��������s���`n�nC0>����t�.�}�WDʤh�l�3��窮�=�K�$��5�35��L(�Tv(V�2s�M�kH-����ڶ�h����>�g�pʄ�I��p����𷆴���Ɨ4�5��)jm���B��A�-��<Nh���;�f�Ζ�xc��N"s���m�wN9��@9�גl�F�!���Z�׸DJ�
,�uF��-�.2���$�Y��r�iܛ�s]C_<�#��$v�b�,���A�1� F���,������'��G*�
�w1����6�BX���|DY;���0�W��/5
�^?Iy���RU����h<*4�f�9`��JI>7j��_.z�q�D������P�=�ѽ�&����Y�#[l��|�w_���l�"z� kd�s\q�h�=5��Ҹ�)E�fRn��PN�@JU���J:��C0ӼK��(����8�Թ��(>�1�����>k�}�.<�۶�r~���mG�Ps�6Ai8�_�J���]��`UU6>Ϯ��_۲��������`��WJ�g5��\��������!U8�5��:�ۘ�*��Ԅ�Jq:Q�R���8�U*���8�A��7dcg��N���R����mק.$C	�t����)5�6��Vc]$�b>�rC����B'��r�h��H�>_�15|6+��J�n��Wg�gv���(���(��a��I��/�K�-���F�F?���"�F�0��U��W=�S1/�x�#���(�L��?��ާ����}*�?<k�'���t6�v�+c�,�B6C��2%u	X7�����"#E��ų�j�	{֙^}��"Rv��<0<>_���G�x�(7t��	�0F�{@����c�.'I2Ml3�����ԩ��8*����ݩ�Mdq�C	~�1��T�uU!�t�v��xiJm���,�͛>�J?n��s�L�oM�q%��~�n*�.��S4���p��|o�+�sF�/8��r����6�`q�R�������,:�Q��,b����~-����G�i�f}E��w��\����پ~��u+�, �]�c.,�����Z�"՝��H�Ý�f��g�n l�N��7n�n�~a�z��:Z)nx>DSa������kf�=��U�)��L��*��_��ѡ��va��;���M*��uP�@L�Z�7�n��������wQ%�^Rx���9B�t1|.�V0��Y������׿�sj,���$�=m�� ��8�(��:)�UQ�.3e��22u�meV�Cd��95Gk���E�t-�rR1�J�@b=�^�d�CR�z997*B�����`>���l��S�oR�5����7%�l�r���.�a�1.T�Z�Jbfs���8�Y��ng���T�^>��{�}{�/�{��g�kF��zz����0	GG'��y�g�V��萙�T�E�Z�2QڥZ#q�l��\����:�w�ŽN�sOS3�Z�mj�%g�����t65mM�b�������B�4�j�����=i"���'��d��cl>0����w��6��bg�>ϊ(f����{����I�*��9��mDt�����}@\�o��ݪ��`��_�dɿ<���뇁.Ɣ�x1F��4X].H�o9>i#*�!T�=����᧟��<P�}CΆ��7Cz�ro$�Wv��O����9�_��"�p����q��kC�M���z�9��Fx&S���t��o�$�
���c!n�:jzh��x��SU�P̜�u�����1GQtzԆ��c,ʶU�igDM�H�먔5SZ߻���N�~/��MS��8�,��敓9�hHG�6�\��)�(ڒO����:���9pp0�v'5,X�"��%�]0]xm5�L�!�w
�H1چ���������c�׫Z	4M�cQօ�אeT�^�`�׆s-�АVc�0�z[C����n�q[K��ʘ�)�uX��F�Ge���a�":���%�bPҮ�H�Y��;�qur�(�����g?���StP��SW��?��gu1Q���D��nݽ\=��V��(�T�H�� �9ђ�ަ�='��ip�H�(�!X�5���-8�n�� ��"��P��aK�1X�N��%6:���	�T���Ǐ[4�׈� �1�ʎ.�acA�	'��wW�5b�<�"n�EE�����0� �}sb8����@��y�5W-5舴a:b��!���������R1�ڡ����8"vZ '��J���GE--�t^�#t3f���}UQ3D��"�5F�_�U�4A� 	�s�cCm$�`0��:,o�>�s��l?�ʀH��a�=L�Ħ
������#��:nu�bC��m��v�5�;�65l�4��J�A��Ym���PV�`�)�Fu׆ϵ�ֹp**�!�
���ZC��������kXiS]z]h��-�T�ƫ["��T}����h����r�0����WX�s��Q�@��W�Es
'*����� >����K>W�	�"�SO/SO�a(	�Yxj$ �nȞa㱌���4�m��G���*��W��kN���Ew���^��zK��T��ZɿC�6ܛ�h]��r���ܣ�k�ty�4��:�;��bR����3�)P�q���J�x�߅!�/2�K�/v�?�le�z]����wKK
��h��mD�Pe@DG�XE�����`��E}�1��P�=��DL�o���f
An��Hs��@��AM��rM\��ǿ����|�@'�m 6yT��d.Ἆ��uy~� K�kz����+#Y���Jڒ�f���)jKhB9�u8ڭ��ud��o�G�<��5���-�vm�Ԭv�qi��b��K�����H�1ص* 9�����L�\*��"�O���D��"n�!:�F�a���}�#�;�]o�h��qxa��~��7.�k���ߍ��X���T�5�H��q{ߧ� P�t>˾�\?EJ���"���@1Lµ���9O�e�脱FS����r���EW|5���=J�7��!"Q��������Jjւ9�A�A�S���I��F{a�n�����Í�w	(Qj�f� ��0�\��Ҳ(W�
32C��E���27>�`A	��H�zpA�R�p��h��ܸ�C�u�$�q�����Fq	�����i�rN9t�����o$�wT��!�xk�m\Lgb��.�z>����p���n��,�L	�\"cq�4
|GR������<vb�1�P|�$x�A�km���e������:J�'��Jj)Q�,�������P5�Kc�+絭�8�
�`��X�V��y8��3W��q�Պ�:c��ν�j�����9���>�8�B��>��m;$�W�Ҁ��W	��ϔ,�HZ��8>kx�S��%*~�]0:m�(*Ǔ�ɹ|��Cy����)�=ƁG�Z��!Ҁ��J4c�%
PV%ꕶ�bָ�Q���%���bHL�#)���b�����<�s����n�^hJ�9��}:�P1�N��oQD
��CP��U���h5u������L*7�t���/�h�kYׄ[!9������Sa���E����70���P�%��S�Wi2%c�1IT���>;�@<���9;�n'}�N���p�1����[�f�3Z��c����%����z�s��[�ä|�0hr�O8'}W������Yc߰p�|-��Il�H黔��5�5�����¡���Q�Z����Լsb�����a7R~�Q��q��3LC���\���{���]U�ƈVVɫ��s���aLCCuI�^�%p"U�cFN/�f�J����;�<��m,Q��ν�:�Wx���)i�R��-=f<����h�k�K����|�%~��	#,,�~������0�:EdgC�CjH��?��vc��8��"/�匋�5����oN���f-a����a
6>"/bV�F�C�a8���O��U��lH�6�JS�ś@$���>���0<�n5�i"Q�l�Z�=0�g��*�2t8G�����)#�w\G�>i`�(N��cԼ��1&��5��Dq�T�#����(��
�d��ǰ�"��J��xg8���0J��L~]Ŭ����Nb/-�A�
�����V�˵5�a#ص:�x����ا��B't�4CY�Cn>�����3۷�g�=CcE���|�5�j��lyJvm1#����s%���*5��Z���z�r��w��s��m3�kb�SlT�yKV�甇:j��r���1�:��.	���<]1�qPtQ�X��p���c�ǥ�����Q�rS�UӬ�B�9j�����EЉ��b/�1<�W`�2�{)�*�$��d�5����5}�WD����Ƙe�
����������mh�z���ύ����P�f��ʄ�\4�ё�e���e���'����և��C\�1ו��"�Hgȳ���z�~�6IO~��o�a��L���EMF$\4��ҍEy����Θ��5'e
+��p�H�w,ʌ��<�N��᠊��^G�}�u)������!�+��E��k�a���Y����G �0��(�e��3��<2�u��
g��aB~�g�M����q<Qt���0�T�z��g{�N��V�X6����3떵 d\����(OL��{ ���PE�wwb��湫�x���N�*Q� �5� F�7���H�B���U��32βc1Ѷ7َ��7Bg���Y �_Ү�$#���e4H�`�=[?��a^.M�_XEc�Y��;
3�%��}]�6/L���t�P����샧!%�yP�y�1���k�t��������KM+q�P����c#�2hM��Ҷ�E�H#t��cY���0�Xj�*]�~�t�4 _oղՊx�)�\�#e�(}Ƶ�X:Z�l�����4n��|nq�S \�s6l�Q?ߎ����a_2��?���TK�)�(��%c��Q�~��[��^Όt<�.��ƴ��$��=8����bةӈ�o���q�Sd]_�7߈n�3�Z�X�ZᎽx��q�����C-��߉V�}n�~��r�<�B�`�|ID�떽��w��
��m��� �'�y�~S�6�X*�����%��ض\Q|vR;t]����˒[o-n�����^����E.\�1��������Դ����BMU��!�NېN���Ey����a2'�*��m�����9B|v�H�p݄�e9_=c*�Ē�ŔJ��'Q8AJ��%+���YS�Å�1��ƈV�j[P�:X�rT����.�;�T�K=�X2�R�IڇH�Xǃģ Dm�K�T͘.�#��K���*}�d�"=t�j��~f�ib���9�������e���K�Y8���^l��������������&����w͹-W�=���r�b��9�Yd{ v��8�ʴ���	�]��y�ǐ$�)zF�`�9�UD������N�����$�M	ju�PLs?>��������&���Ü���n%�|�0Ͷ����Zq~�E����\�#��w�J�m��.M���(��6���o�?����Ra�Ɛf�.pV��n:T�4�um��i��Kf��i G���������ʐ.�������&~��aeQ�[�|E�����{+�e*o��5��`�Li��T؁.�vx�w��0Hla���Z���������)&-;Z�"�4��
��m���Ez���O����#�&��L�_��s�: u�W2�Y^����.G3�����؝8�,����9"s52=|צ�pv02�ҫ��%[wW�u}�<|P�qc�l&���3��Ԍ�0e�B.�M����tɴ���£^h�k����&#�a��9�~��lһB��5�p��F�D�0:���y�ׄ�%��OZ�܃`�㨝Ӵ��v9$�Φ�x�;Ȱ�ӫ7>Z�߿w��,��9z*�.��M]�FѪ��P��0^���4R�`���Q��G7�T��s�r�kg���:(z��BSƱ�=��@`P��5Y�g�����`\��Fwl�6"�ޣ�`���T+CJ�����lL�N���Nݼ�7m�^)wi�Z�Rww��]�b�8G2�b�K)�*��w٘�na�/�����K��8��8��a]���%��ُ�>n�|���=E���i\
b���
Sq��?��������8Ɵ4];4��j�*V����nΪ��Q�,�ʄ����կZ@�+hFόrMq4Ƕ<�`���H�$7ϼ>d�8��~z��I�`-ZQ��X��Aw�Fqzk��+׃�#��eD�x?�?�!�/�G��t��
�7�7�f�{�eUA�K����]�$/�1����EY�݆-�eJ�.���1P��.��������4����\ڗ;v�X#t��3ɸ�'l%��U;�:q"Ý�u�/<����>T�+�y9�$x�j�&����{�h�Y��{��U�梳��Y�o�0�k��V��Χ����x&-��i"��)�bФ�i<S��������+S�J��K[-+�d��^�� ��6�� ���3�gZ�T��+��I�0�vZ	�莉�k7τ0[���?�T��+��mX����?�1��ɀ������Aaq��W�'�B�JX�$��3u����"�/���S�ꮁ5-�*]J��}z��4e��&]k���؏Y����Kx.�o#z���u�:���`�S�o��T��V�S%���P)P�o��>3�o��5���\&RW<Kl�S̉���B��H�$F��!����ÏL}!��h���ې�����k�[���ܸ++-�&��JIL��x�1±-��@c
��V�8�)_D%�����mo�e
cHq�E���v���7Ulb�Q�#�UN��1�I�;C:p�F�F\�����=�R������������K�{��Z���s[�~�����=ᔝT0��2��h`r�,例V�!*�>C�Wl��/�k]9�Q�a�N���H���!߼b��u^��aԆ�j~_`IA+��%�OG$�̇��xP"r�b�aېbct����b���}u��*IO�q�/p��N�yD��]PS)�!�r�]1=�	����t�CM��M��"Z�,U4*݇l���'�R����?d�NX�u��ȓ�a�HPn�V#}:P��|���TԎC��w|foB���������H_w�v�((�WA��L*6��.h+m眿����T�	Ro>��C�����M�m����g�S:(8���.��1Ac^�'G�h@����}��"�v�������E���Kj�"��P�RC�(��OI�0��~�9& �!aV���d��ΧT�
]XQ��ap�{�>)2�|�8{��߿�.����%��Cf*q�t�~V<7���
��}���:s�Qʣ����}�
��َ���y��o(rȺ�hp�gv��Hw��
��O�`�)"M�yeP[���!�
���0�h�bb�!ں��E3
 e̶+/��EqhY�sF���Q�
3-<$�go܊�� � �/�i��ӵ�$�m���ϰj�b���,��97��c�͚*F&Rc��+m�i���vEE�~>G��Q�����߳�c�Ջ���ܞ�Z�9ύޟ�\���Y���g1rW��Ey�)������Q��C� ll����:{#���^�!�����������g~.j���$�b!�p�p�۟�4��s:9��X	\������P2�3�/-�q�J�g/��If�`6K<f���u{�{�DS8,��(Dy-�9ܩc3������l��A�d��)'@�Ό�y��0d��킂U�2b��~���Qd���-��Դ�g X���&G2�M��Z��׶fd�`	�Fm�OO��4�3�g:�V��>I���+���ؿ��ʘ����*C��q2�����(��k�6�N_��0�!Ҍ��o�Cl�/�=�vLEU@J+�0�fK䔅���/ײ!P[<@�8.����BU��Bd��h�"_����`H���S�)~���)6����,c���#a]L�{����%�d��Y84PE��ǈbD�6�V�
����A����N�YxF�ka	8��(�P�����5�k�t�9�o���82����J���
�G��J[]5�޴}����+-�#l����,�jc��~[������6�Wl�.�͘2��BY%h���X�T2<Lآ�q��J��Nb�i�x3Z�QsИ6��|#������W��+f��k�jQ��]HE��ߚE�EQ�|���x�������W��~G
U����1��N�*%�<sg��&gO���+A;b�KuK�T�5�/\��Qo���Ҽ�kkgۉ8�0�cL�~:?��TzU�����׌EK�䓐����k�Y�Y���U��:+ƩL[Y�f��~��-���&�
� ��x�yJ��+�1#o^�c�w"������/�ׯx�=�؊M�L�u��5q�)g/`<�[�?���k�q`^H��t�5��R��!��)�gX ���-��JSD�������.GS1Vcp�ךl�`'\�Y�G���'�͈��z���@�\FWq���w||��CJ���R�$�_W=+��|�����qa|���o��}㮹V%�ڜ:p4��o�^T)��*co=I�_Q@Ѩ�4<����ϟ/q�0~�&آtD�h���_���{�S� �=�7�nnoum���aH��Xs@p�X&����+!��Cb�a���:*r�\���pMk��Itl���nc���10�2�o�O���ˈF7��TI"�=_2��Z\�{�g�P[0�i&��cv'����/�p
[�������t�qdT�_b���̰�ƠS�=���f`��]`���Ѷ��i��:o�r�g�o[^���u]W�j$Q�W�au�``��o�;3��(<��0f���Dj��SG�z�����X�>7&�(6?Z6�{�ZҎ/����2���F���#����Q+�6>Q���L�`n��rC���v�QTI>��e��}�x腧y�Cd��
�'�o�Se���۷S���=z�G"g׏��)AHѼ?�F�b��0�P�K����u�A��<U�����*>�W����� �-e��s��l�5�c�7Ñ�"zrKY���(���4����8	�ܤczU_�B��6��aD��3�/_ޤ�h�tQX{g�؝bf��q�:�IB*�G��YY5Ez��O�Cꞇ2o�tzǮ#�5on�e����r�fe��;�q�nG�85Vp��{5
l��ܥ5�jᳲO��9��}	���q�>vҢX������G;�F�=�iHj吴��j����������U��hP*6����z���v\��fm��+R��v��g�]gw�,TO� �'[�YP >�����1	oT�e��Y{l�������XI������|<*��l>�);R2V�y�JGZ�K���3�Iv5r(N���j�
�ot�*)���ذPN��DD�p$��pz��������Yx���UX\�-H��	��r�Z�I���i]q�Qx{�bG��I�:#V�ki[l��DpU��t[:~������Sg���ٙfHf1`O��X�7p�9���1Q��5�������=��a?�r�^�|��}���V�z�kA8�;>踺[_�c�e�Z�FWw�He�=��]-�1B��y\�?��V?,���Ԩ(ΖN�C���������g38pga9��[�+N�.��>�ښ�N�C$`�P��	Y#
{/�#�fM�n-�����Z^�F}�L�:��l�R��Y(��U�4��D6����'4���4���oCꉄV:g��1Lc�ʐ:��C8�����p^���öpH_�jm��VT�����}���\�W���DO�,�͛}<\OD��q.���N��Q�{&"��^iڭ�57����|��)9���w���&�G~	��(a�ۜ�m�⢖7� ���>[U��r&����S$���/�Q��r��"t�)����÷��׿���m��c�P����!՘�o��IU��Un+��0z��W��ḏaGD��te��Ց���<���U�o�A��6�:� 9s�6�"���^�I�B��j��v*�KF��|�t��Ǐ��o%����,�d=ԨlM��=j���a�!iV���lY$'���q��3攺�A��U���3�����X��y��[e���[ɴ}. t�a��yP�7�g�)W8e����1佖�6͸�,t����C�_��m�gTy�|���=�`�Rk�cw�P�c[�%|�\9]g3m�i�vMD���lH�hc*K{���� �a�`�ݾ7���jn��vW5}�qhD/¿�0��.r�u��i��}QD�N/��m[�W�q8L��{��`Q-���f{����5"���ϑ�y�����P����hq$���.vo�pDц�| ��~���x��G\_T';�0A�M�*�}=�%y.�X^(�oF�0��_E���A�O��x���өR�V�^�.��m]a�at�~�	�l*�#g����<(�h�Z�H��@cxNV�U���u�G�A�e8.,�uP���%��yxV����Z��C;D���{�&�d�{�&��=�m���~'%�7��G��Zo��81f.���
��W��bW2���X���";6����ߢL��NB��7�����������3i3ћ����i�k�fs-�Z'�:�m�:Z��Z����K48j�B����N#x��uknq6���ڐ"�Ҍ�*���߷α:�ׯ|�]��F���kx�*5��nE�f:0���}�_ѕU˿��/�=�h�T񬓢�I"kfX���x)x~+��z��rPy�+���m��������2�q�cV��� �RD�@4���!|���aR:����´(��d���a��)���9�'��p��B��u1�����:iL��^���m��Mό.�lP�^�[
��4���V�R
����!��`�J-��B@:�7T�w��a����Q� �?F-�e���>|H��g�ɑ�SJc���,nr�f_����u�D�x�r���xv��˶�,�}��)X���5S"�� �wq�`�#��R�pQ������	����h�8>�g���|�=�B!�a��"/��tvq��YHњц�@µ�rڬ@d]�L�����)���gB�i�?��x(�*��Z��%Y\��fc�L���|��5��2W!�g�3�{���s��&Ӽ�P�z,�-�-�\`��=;�\��-;��g����&o���R�^�{�7���,����$��:̗��������t���E��\��4�ƐZ?󠢏�ۃ6�cx����Z�:��^�9�ɒc{)图�$���X�m&b6�Sd�(�5�/��- ���n#FZx��xy �:&�=�ENN�S8��tqAo���#��"�
je{υ��"���3�)IG�İ�kO�(�F4��u¸X��a;4]�$�Vi!+��<Q(�{詛@ne	'�n�)�dO���׬��|}:�dI�&�����IǊ� ��!b�2܃��I�YP�0�œD�Q��sG���xO�f���&����k�����dG��XDߊ���?���B������m�c�5���P�J=>�>���uMO��vԅ $���9`p7S���p��?������������	��)���e��(�m�ÞY8/���\ �h���C%��p&�\�fH���0j��$�n�c����U!(�����>K�"��4w�ǳ@JO��2���ߔ����n����������!��$d�P���Rw1b{�ϝR�Xh=���6*��ۛ>S!�$C�kϼ��
���i��|���Z8��d���N��O�x ��M�`��zj/\#R
�Vc���H�MC��t3ZOY�;>��_��9(}QU��ӛ����}�Q%"RPn���6j�W�� C��3�Ut6%@����%���ME�����L}nr5_4DcFw��(FFԩP�!�c�z:q��t̌w�6����혃��x/��~�X>n߱��"��1t���fd롥b�eb��F���6�*���áS]gdD��������%�����!�Nx�h�`�����ֻ�Ю��N��b�TD���]���y;�CD���}C gRz��PCFo��_�P�:T� 3�,��p ���g�PO��w<[���f<�ƠQa�H��p��9U���Y�OR��5�p�`��U{2^�"�_qJ�;�z���gOT)F��N�QD�8���=v���j�3�NȦ?���:�)�[����{���������j����ٶ0���p���!�� C���
1i�3�6G�$N)�ߥ(�(/<��0^���V���|�h8H5����,��ssӦ0����c<=�ʢ��N��/�`z.�3w��7Ґ>�τP�p�Y�7{����3��ɰ��{C�%��?��]��O��s.�=j@*�G��}��k����Qtj=�S0�Lw�(��q�MP���n����t�>c��`�ņCH�������͌��'�_��.@�� B&�M�{�R�IŦ0 7��z�����.OrJO�.ra�b$��$�����P'cZ��B.���>k
A���)�`��6�
���=�o$<h��$�{M��Ɨ`���b�zZ �jd]�G��g8x_��(�E�Q���R��#����e��nʳm��[�<��Gz�>���X�s�Q=��~_2����U�M
��+���H�F�=0 ���E�ޭ�Ě�4��%�َ�[�] �����~U����!�?����������ar�Z�H�xE_�g�ϵ��bŖ��ag�
��T�}�C���kx��������U�=�|�F*3�2^�,%�06Gͮ�!��K��Lq�,�=9��z؂O$�u����gUBe1�MnVu�uX�H�P@��E<'�/��a3�4D�p�f�7��gB���o �X=�R�������|ԍuk.7u`���#�9�"�nN)d8Jt#���|��))Y04���}�r��ī��X�(�B6�g�5���F������K�Q���6r0ñH������s��1�A�Ն/;^�O�&��8X煎紭/���11�m�� @D�1|n�����[��h�x|�s��
a�M�)�����SMad=��E����͈����hT�����a�ʎ8\.���b�I���)&�iL�����PѾ�ʺVA��{|s'�_��?�|X�@��!��[�/��+!�����a&-�
��Ws�[H��7���6��� ��!�hL���^wJ�����D� m���|�L�X�*X��6$��`QiE\��UԆ��X�*
V�؋3i��j�F=>�	�G����3##zkB�oxﮈ��H�_�c�*⻟�E*��Pf�o����{g�v�j�)���`'�:�.���ھO3)p�Q�L�4��Tz��gu��JM|Y�ԶQ�a�.�O�b�q/�쑽<GV25{`I
U]c���m���O�i��r'N2��c� Gnx_�ge �n;�̈�����눭�6ď�~��&�`r��B�i3��x�����)���HV��34�b���*��?�J����Y���?�n�n��Jg�[�W���E�ׂE���cvΠ�٦;�AsZ��0��gwR��t�̕�m��5#�H�\�(���bR��B��u���J�la�r�ºG}��W���|����«)�X4jw֑��|���!��;y�^�4�
O���:�p�^��7;��}KqW�iL��zᪧ����E°�]�`�zHgR��KVxp[u���,��%��.�zH{]��ȜE��e;1�VMTI��w��d�`a�6X�Z&��t��4�Yh�h��� �0�`��^�����oj��� k�rVЇڈq��E:x��>1��QM�F]���,Mfõn�Gv̽�r�d���`uw,�R��{�VZ�,�p�օ�3J,f�ڨ᜻�
�	8a3�!)�7��Ե\��5���L��=��+h˸�,)��$#�3�N!�����`���H�� ya!�m^��s�0/^�fʰ�jo�F.��/1U��mqyR�S|m���~�M4��]�د���8;�2�XG���eh(��k�W�Tȋ��A��>6�E)}Ua]��I�!-���.,#�N!.UϏ>#b{�*��w���Pa�ޫ���]w������$��W
�6c��ڰ����0l��M�H�������R��(�C×�T�b�&�:uyW8����*��i�T�Pp6ǠU�~��`&j�IX䋠	��{4��c��:Q|VpJ���W����HX#�U�Tald�Z�F%eb�H��<H�Cq�:���u��`���J�7��FS5�S���Aܠ��N��=�*o�{���r\��p0�i�C��#��ߦRQN�Tm>�"* �׺T�ʮk,C���:��PÜe���C�L�N�H���g�hI���t=�0�3��̈g#��6���i?�yҨ��)���g��<'��j[뢬?���e׿�}�\b���tT��v���1R�<0G���>�g�lT���
�A�_Ԥ�@��ʨ�^���p�y^����R!I��gD9��CE��D�I��Ln��Z;�" ���$���t�(�d��d1�*�}�=��:{�����,���֮��]��j��C\	�,B���o"/
�,(L��Z��56x;���� ��M��DF���r���F��Hv���Dqx�`�®������ ��r5n���SD����{n��=�Q��\�%��)�*�k�Z��ǁ����p�E.,�ݾGwu�+O��L� �z���cD��}��u��D�^ p�|
?l��Q�3����K�1��R�t�1�V���@E-*Z'�SV�mTa8�@���"���g���]*,٨�����UZ����Ru^�	�&�����O[��*�� Қ��Y��`A�Y��M0~�k>�_�b&���ohL��<v;q����ғ��d��ض��-�tr|A�E]>nZG�/g�Ԙd��),���?_G���h���eY�)n �|W��-��Ϡ4�勶�V0 ?��$�>hD8���;��Z�6�v�J����g�/Yg���g�H�q��;��_��C��������P��⁓b����a�Ԝ�q8̫�	��F� :��Z3ӰIe*P�^�Q���Φ��&I�o@[��Rj/���̒J�^�%���#�a$�h���+5�,���h�y��|��C�3��_����P�Gѵ��9���8�������u�6Ɲ��48��P�����ٹ�PS%\�s	���Y4���>�c��"4�|,����u���������� b,���B'�&'����黽����Yi��9�f uI�S�(���U4�l]�l��+��}��K2=�o���Ad1Ǘ�h��2ژ���e��0�s��>><&3��t<!�~�|e�QPTÀ[X]�`��ʲ�\�cD���,�7e��~w{.��i x�b��ߍw+���,�y�R��ciM������̕x��d
1	W\�8�Jb-R��~�i��ڧnWuz�����~�S��\IxD+�V�j�u���r�ݏ�$�wHո��,}�gʴ��0���ƮꝢ���'H��*�T6���3	4��6��ZuIE��٢�\�7�V�T��^s�$
%�y�eW��W.�"����i�5���#�7G#��Wb�h���1��܍d�h�Lvn����Ү�Y��.�l]��ਣ��g6uQ�`�[�Y�I�84B�9A��2[	����٦���#5Ӥ*&��2/�qn���:�X\�m�'�5��K@\h�(�ptF]O�4�\��(���_5��f5h�@v%)�������A��0���0˨V�)N�>pj�uW��1�Rd��y�J���}m@kP�}��;ӟ��}U��C��DJ�y@���Q#-*��e/��l�6~@N]��!.l�N-$�i�8,��]·�b���U������,"�{Epm~[��o����V�*ks>I���������D��$��е
�8����=�p,�zϵ(��)��+�ު1d1�tG�^7b�y��^��%�ܥ�9ش0v�S���*k��Y=][Ȝ鹐�y�H
�9���Qs�p_�U�R?E�?O2�����DǶ�Q���.C��,��J�M��3/�ERJ��z�^;�fUosys�,g��Eσ�7m��i�^w�`]�Ί��ϙL���9��nG�A��Q�c�%�*��ɧ�Lxl_�b����瀱͍��j&���n!o�uP�h�g���ʛ-Pfٌ��s�H�>F9eቒwt`7��� V�̵�w��ۛ�9..�lN��^Ic��7>)�sU�k�!�!����K����O��ّ~PA�?�"��*�ϣa+�Ur��4�	�q0gW�fzd)����h#��T�_��I-02�����fɂ1B��o-}��V��@9���"6�1?4
+��|�I���)������H5��H�A��掂��\�B��k���~�(�?�{�0ɪ��VM����:��E��	�LeKnzٗ��7�؈-_r�4��Af�ScHo5G�k~z��L�}#EEo3���R�� �q*��R�HэtG��!Z7a�M�����X���	dj	�s\��_�hS�d�Ds�v_w�SR�(!W1C|���D�=�>�lx�:B��n�eD�Z���O;�6�\��ρӆC3�ϭ��#���cm�Ta�l�#�V�!����-�S�g)�=%����ۚQ��>2O��=�%���,^F�x�f���nD��0
���d�D=�w��,��(�jR�i�	W#�
�,u�c��C#�}���\D^G!�F��i��h8'a�-�o����Z��{�.6���/�{�ƽ��U
A^����z�ￓ��$B���=7�j����j��L]m���Z��{�#�������헿sV�����u�u� 1����MwȔ�r`�8O���s���:~���)R�w�mh���`uޝ�}Y,hR�/�q�hO<��y��p=q��ϟ�7:M��^�1���S�(�#\c��� �w�4�5�N
�i>�$��y�gOu��ta}��f�13�H��b4��3�MЦّ�j���r`��4|%��q-��5FQ�2B�՝�
�����w��B����.��֢C�*��9}fPQ���L�o2Ev!���`O���^���x�蹡F�!c�#ڻ.�]na��N��h<>����N�t�1B/�(H.�:3�\T:���	aͭ@gչ�s��26�r%3jK��Φ�+��?�-A�g���7Q\�,���ΐ���	��!�Ñ�K2�)�4�rVG���<{�~c�DP+���O�p\�C+^K��T94ǎ���`����5��m㌯oRdG����>��{a�cα�sJ�L���Do��K[�9;���h:O���Qɸ����V�Y><�I��Na���z?O7�B���x[��U㑓_���ϙm�P�މ���1�]U��?�ӡ�cB��D��I�b(��=�����?�9.�9Ee<Z�wWb1xQ[������*X)�xb�|��f��8)�����(��l�҅�>}��&t�������$Ir$�A���!�X�{'w��E9�[��ú�IU� /�T�ܳ�g	�%P���UI"�����T;u�M^7ͧT͝��S�v6�!
W$ ��K^'�[���0��x!�ol�m�F�-����ٺ伆6�T�h���n��{WY"���Y���L��Ч]WI�	�Ĵ��S��6{�Z�z�5]��?R�n5�oGW[�f�m��e��j���?D�XW7;�m��|:s��D�f)����0��I��Y�� �����Q���t���o�U$Y�A��r�����\`����T"jU�=���uLA��ٜ�Z�StR1X���+�-V�u�����7\J�$�s�PO_��I��sv�]L����ٙ|m�)�{��%ϗk2)<R��."�[���ok�E��@�~���l��K	p���K�K(����D��Y�P���kl(�����o~0J�oA�R��Z����+I���ԓuO]�Xx'\f��;꽡�o��q9�,�m*9�I��ä����A'ԒX�1t�旬�"�?���	�����c��`s�m�5��I����Nt�%7<�ȸcp�z�Ъfr4v��tM�q"�1^W�X�0����gz�0I❂]����C�77���N^QRR������4��U������|6R�aa���Aa>��߼fSg�;��M9k�����\R�d��0������?q�(�v'�O-[�"��Ւh�x�!�a��`@�"�}��hd���}�s�t��n�����R��93H`�P����.��#3�s����r��b00ëzJp��Y�r��둄xIZ%�YT��Y�/��+qY
�fY������O(\nY<%��P���v)��|�5��E���^#kEV����[�A8�v������г\�{C ���3��������?����� �@ښ,����Q���)C��:�\9��� ����E�����B��|;��I�q@[��h��X*��;�׊�jh���)c?wÛ�T���p k=?Q��u�2�C
���]��\g�R���d4��ލ+�d�Y��
}��>Őz�F�)B�Hp���?K���/�������5����s_�h,�d�L�{{]������6#�n�0��y��=�χ�ڥk���R'>N�N�Y:�}��C<��3�Ň*(��Q�$�q;�[)���`@��H��E��N���������suX�B7����z�:-M/4z�f���NCe���.��3�Iy����{��Vٛ,��0J����"=���̒):����f�{�N�m�p4���Մ�~��0~m���ZC,-��Ž?q�>�φn�kf���,J�^�q�=L�[ēu���u� ν<�,;SeJt1�������:]���bzѸ�y` Tx')w��c�㐊��*�vez˼�i��#�O�>l�Ǯ��j8��r��38()���4~_;��>�"���{OK�[}��W9*�Qn�W?���!�U��eҳjH	{dW<O�f�1�B�z-~��Zu���������jA�[2����6{���6zv��6I-��4���������Anu��� ,q:��k�/d��dwFy�#�k�\JInT�75o�	���oj��
�Qr��f��d�[b��;��m	^6qڬnP���7d5fI����h���UO�.ac�xNf���@\E�)g�)yt/O�`�ωa�=�9{�aC�σ`bkl��c� P�ȩ�l���Ǹ� �c-܎�������j�ۍ��a�k�#N�^��{:�)8J�g�wg�$VAq�Bț��5�T�\P�c� ,��5:Jڸ"��:���3iY�JL�RE@x��u���M��T8dƳ����΍{X�JG1d"�� �m����R� ��盰�>�Hg\G���*��\\P�
1��!�l��Af���|�70]̕����p�萯Z��L��[kS�+Q¡�����g��A��p6[_���M�d*��F%h�_��z������:.�1y��t5����$��T�ә�#�7]Ҙ8I�@�gJJU%��%��u7�Et��l�e��r���@i�����p,un}Vv�n�/wH]�Ō����xA
]ɽ'���
<V8dC��OĿ���L�:�������j�_ؤQ*k��~���4�{�U�dd/k�Âl��h�? ��e��]��ͤ�P����?�6���w�^�ǟ����g?����a�R�+�l'�܀upD��>�;�#�|I�m��z�v���Ի$�� ��4����'*�y4q�T���	�����9�aiH6a�V'u��]��PL��B���M�q�΍��(����*8g�nd�����q�=}/���B&�2ؗww8(���[�^�(���~[޽}{�_��1����K��J�ВpʲL����1#��*h��bY����e�_	������������l�v��O�/sf��=}@_���m�q�s�Ѡ~J_��I��J^��^�
4�`[��y�n{2��A-r;��QP?|A������(�_�.͜�"����]RJ���vWӣlU���v�}Ԓ�A	��0џ�����8	�]��8���|-�E�L���۲P�|��>����pk��.���)H��9�k����b��@�z>���c�x��m�F�/3ue"G
��W�)�k9�h2��f�/���!3��6��	~��L� ߌA��d�YpG�� �Z][���/MSeT���2m	����7�5�eU}ӹ�s�Ʉ�F����ymtU���&�M�R�E��bu-��GPe��9-��!L뗎���-���a a�p���ļĵƇ��ۯ����q;�?]��v;�/	����y����4��8W�y�
�=�N��e��0�I㩋��T^�����y�#m��R�if��'T��3�~6��7ֵAo!VڄX�(B5~f	`���;��a��A��&d���plb���i���ٜ?��+/�^t��qZ����1S���X��c��[]@���Sm�7�^R�E�#�#5XvM���P�l�x��t"W�2m�ʷ��I}�b����~4&Λ��28BY�G)����.���36�2�'�k��,qLS���	�c�����Sl����{֤�����`Q�ȅ0��@�>K�Ž��%~Qg���y�sjW�g�n ��NB<X�$�۷�$*���g5A�����E�ƀ�q��3I��	�X��vx�"�6�˵wD�m�
��a��n�� �S�O��P�o��8�'�Lw)�X� �yY�{��p��l|Ο��T��kHEU�0fՁ���G?�0]"�;�����[�1
�O�@+Z���&\p���p{h���_�r̬��cm�O���뷱�k��O���	o0�1��x�I��@��:�q$�))3(g�.���%�e+ZGV�'Zk4�P�X�ռLE��L�d�.�L��}��[[j�MZ��7�z�8��<�k����:]?�؛����=�\�:h�� �-Ⴌ�c����X=o���
�n\8�� v�h�Z�z�I��:����9A�߭-Р��PUC6��]뫔�����@9~���9�-=*��;6--��~v�=>�PY�&	��B����c�x����F" �-Q��^��*���m�g�����O>~�����-ZKfgTII>1;�Q~v@>�q-�����>�#��:y~��������WƈL�q	x?
��#�H�O�)+.R7<���?�esp�S�Z�;�{��� �P��o�>Ӓ�ن��6��X��sR[��#��/�0C�x���e༭�M�o晘�l���ky����œ���~?;��^	#���%���N��D:��M�����#���$?1s��j����YiPḱ��A�����T�K��Ms�r� ʇweN ��y�bë��\�9�̝�6d)� ���9�����a��i�P��_��Jf��u�AT�#-K\�Էg�'��_C�� ~8شm|c~��?�{�X�,Ec�Ȼ��Fn��02��/�C��z!�����pc�Z�2���P1�-U�ą��ZW3y����ohM�Jpo�^�=>�ԦD�����!�?O��4q�$iG�P�E�	�E>P�~�����s�[ЄGE�\�e !�zRs�9yӥT�	H��B~̊M_�ږ�s��Z��� �i����$|We}��)s
gџ�/��*l�I�G��I(�3�_�(��=�`�'��蹾�ᱝ0�\*��u�XK�g�ݲ'��yk1����Wk�<:Fj�uK�Q+F��;L�p���d{����D)���C,��L��L�]���*��4��,��rM�RN�5���M��t���Ձ�<Ek��c�U`�S.n,�����P<�m/�K<�'I��C����{�bv ���(�C��Ƶs�i��M'4��;f��C�&kɿ�V]%�;w���r�y���!��/I/2�%(T*�=gtp!5}�y��O�'{ꬮ7"/���� �=n�.��)�(�E�����Fz=�#�inX��]q��>is�ڒ]p�I>���O��x �r�j�k�qU�n�8���Vý^����m�A,���ג��7���qh ��,^�ߺ�h���Xy�x�dR�a&�
�H�@�!a��j=�J{rS��K��2�:9Q5��S�Ow���Ԁ�eD8V��V{����f�-�؋��R�����������ޔ���c�Y��V���	�褍�T����
&7E��������;��2�Ð�]����/ ���@Q�6�r�J�^��Z4�2�y�ve�ؘ�d6�
��A�ƭ��+5=�n@n���79Yn��wO[J@��*J�ꉠ-e����mZ,+xIs?�s���'҄>I����G͆[k��4��������Jn�)�2�Y'�
gi��j�A�����k..,mw������Pm�ς9J eR<<���L]�eS�V	���s�69���I�E0���2�Ku}\����j��^�a`++Jq�����<�q�;H��A�b���-�:��-5�z�,��G�E�	��O���t�4֘���F&���6&�SP�EC���	����&���w?H�:mu�C� �Ȧ��c���������\8}�`ڐ���}.��q^�H�k��i/�
��k�|+_�HM�#�jM��8%���]��&�n�s�T����;Y��#h��#��߸!�6��v��i9�X���@let���^�r:�hM��=��c�����H����k)7>�.qPB!�>�bH��2^������f@#d'ZQQ6�e��b���f��/ZQ�f��G������97+~���c,�m�&��uv�F�ۙ���	Q~�Í�k�m���=�q;+�IGԎ�4�벌K|:��5�؇}l	y�M�8ȥ�K��A�Y���i�0����W���l/��C�S�-�md�� �%T���Nk��Q6���I$aW}�bS�`W������'�*�a�����~�I8|�����`�� �2M���Ym��A��������Y�1���Ӷ�y�$Tu~�ֻiG��}Z�CDVp�1v:��fhki��[�U�K��s�G��N�HW�|�0����O�BU�����O(��W��γ�uq�?4�7������I�.?��7�[m@X���3F`[2��"/���F#+l/����^��X�`*+�,�??*�np�Ť�z�n��kaY��v���xp�G�NȠ����~T.!���߳� ���kd̕����=��wmwu��#����nz\��s�ln\e��F�3?]<G��;a���Γ;��aK�к����(��(+���~f��,�k��i����H��A�E�Ym�Sq��,l�s�=�j�5����F���;��r��능&�p��t�'�f`�%vj"��D/�vo�Х�f>~)�F�{��%�SL:��nR�*���qf_�8\��E�Y��=	�x�x/5�j���(G�3FTdUS��*� O;���2�4ͦ����y��iҵ&n\����}�#��Dw$U�o����[2U�΢�d�x��`�1u+ii:,���i��U��Wo4N���4ټ��0$�6[N�i��z�`V���S��:9��Q����ʸ��$*_4�*�}A�Y��;���k�_��49ۯ��L�ভ|_��ή5��kd�|�u�?A�]\f4��msW���EVˠ]�Lq?��ӟ�J
LB�疜ݧ����7_�ow������n`\R���4~��"���*�����`����l�%�aw��y�eߣ��ꊬ�9A��a�?�����?d��2��b%��*�5յ��<�f)�Ag�I���:�~We�@R����N<�����O�5���>��[mq��e�� Z:�G�R_l��y�uf[6��W��44�N�|��Sb��uQ���9�j�x��o�f�C$Q��Z�E���(b�� ~p0Y�[-�R5��/Q#j\*���s�-�^��֌��GR{�MSW�}$�j��KJSQ*ZSR��2���$�0��y�⦫�Z�j��۳d�iɑ>r�v�ʍ�9�^�\pm��%�������m�ݝ�}�FC�y8$���7㘣��X8�?}�����`j"2�f�n$q����h`DG�0 �j�A��t$���Z܍v����|�������̼.�s��g �۲��{�j�B����|�X��Jm0��P�<�v\��;~u� 辣3�w�;�
U��y��`XI(��{(�b��R��cs��>���. c}AiE��B��3��Է��o��6>$��&Rd7eε�[ۿR����CN�=���=lCMYF\���K��A����N�T�9�-w�F@�����̮y���Ἵ��{�Za�"ۚU6���2�;�6����a�n������߾}c������BIJNu�0='��K%��^ڈ����4�c\f�Z�!~T��t6�������]O��1��Q7�7��b}b����m�zvE�S��h/���:�h���5fޖ�+m3�N୳RaQziZ��l�J�Gg<aU�u��3�M�E��ˠ�!�z���q���3�4���b*Ь��>�=����h�f��	S�������tkv�4Վ�(F뢌��c���V��!I�v�|��+d���C�zۀ(�p��
��Y�(��:�V���[Eɹ�l��۷R:s<s]�o�㡰F���W���*N~l����O���ʟ��O�@L>���ˏ���l`�`A��o��n����?�g�����EϋD��]a����
Z�L;��M��s�(�C�R��Sh�V)0���(~���/ߔ?���D:���h����{���(���ߔ���o��sP���kQ)l�C	��dӫ�ϛ�o�]���c���M���
t���t�sn-'�gu=f�h���u�x�	��nI��G�fF
g���7���s�d�!�Q���q����^ӂ}�ئ3I�!U@y��HH�l��|H;f�e�ػ�p�)x��T)U��f�]@h��?����`f�5�u.��gn�`�~�Sͦ���6�f�K\���^G�Pߑ�n�r-�,��i4��B�\j>A˙�]�p����D�6�R�����z/6�r�o�u��/�>fsq�}8v�\U��gk�F�s���vS���-���1%q���G����g�PZ�j�ӣ�AI�.���'�v7��{�ga�94:�����W�%N�`#�����YSk��=�s�zr�Ũk_\��g����l1m���!���}�����AV��-�w���5Ij�5��&D�2�D�>�N~ס��D���.����u�542ͷ��~�кW���9i�~UU�
R������{@#�p�<Z'K1Z=�S���q`�wׄͰ� 	�@j,c��Or��A�o�r���>�U��N�k�h|����NA��"-3ᚵ8\�[<\�k����i��?�jw?;�/���Y�|D�w�Kٙ�g���.�<�	����hk	��K���Lɹ�.�e}.�Pv������w� qY��9��!b���۞2>q� *`Ƚ��?>q+dZ(OQR�=#�����L���) �0�V��>���H-�L��C6�b��4���&�<��M-�Gɉ������,n�.�AM�k~N�[�eс��AX��[����o2�w*��9��?�;RX����?O��	b)Ӕs����e'�� �3d��|H�I`��k�g�����-cň�뵏�������� &��3"�>��poI@�uz>��ú9�Hfc\/�R�?s�\FzﴢSdǲى[|/��Z��[F�dv�G���Ͻm�;����0ѣ�Yj��mu��� ���=DV��'�`L�5F�b~��!����a��57��-��c��WcGZ��v#n�ц���>�J�v����+G�5D�r>����~�>�l��2�y�}���}>��|r;��x������`'��n�����J�+?�"��[0:_2�8*���Q�I�-1�_7��N�E>
����U��&f�T�*53
��k�������7qs�*`�8:�Ӕ^1�@8�v��Yw�������n���6ʼ(1��GX�`<��#�"����<�v�>�7]�쬊R��l/�9��Tqke��o��&���dS֎Ĉ����V�C�*&^�cB~_�����<6'��c�,�f2����gÑ�#Mq "���k���ꈘ5��7x��u��5�����x�H����%?dJ#^�
�l��^��T�&����_�����{���u�f�tJ"��֩��{>s������X3�p<�ն���?���M��_����_��"$ _�~7L�R̲��K���Q5z�&0�}ϳ�W>Л�V<���Q��a+��ƚ%$����c�ˠi��������ʌ��	�/3Re1+�޼���� �G��ʹ����6̋��.v�;�j�hv�=���"�q.����T���a�� ��Lʌ4������96�S��c�� �Q�]ˏł�q�&�Y��TY�"�2	�*�
��(�U�Ԅ��h�5	�;�<uu6��v@�{��ԫb�H�?c>k�����z>�OH����x!���ݼ��ز�7������M��7ހ|2�<�>L�d8`�Iӳ�a[fp挾X gAE摺��^Uz�!j����l^)�z]��؃�����u��WuQ�E���2'T��\/b�h�Y�9x�j��k�]r�^�kr��Ư�{�/5��q���g�ӻ��U����@�x�9����C�P��.�>kC���ӭhrp1#@uJ\�@z�h�c��Fh�K��dУ��׻�\/��a�P�o���⢿��s��L�z1L?H�'��4{�*)��޶�x`6�F�Hؐ��鴉�����S#�d˒[W��[X�c�Cr�$\��D�Ϝ#���c�{��i�eP[�k�4�w��@I��9ի�X�v1�0�n G(�r���=2D�6�������V�ϑƠSMW��%57�i�m�dzd|fp)ׅ�u%'����R���uU��S#�:4T�D���*�#�3����8�H��UgF&Xg��������c�?���'H�x�N�!n���U<KOVY�o�W�a\4ۆe���U�].׫pOR|����b��\��p����{pqh�p�C {������!�G+�8�\�����	׽�I�}b䰔�������xH�+9�k�6d�������Ջ�YTC��ۆ�!��B�iRv�5Yj������E��aLڛ���p���1�{�� �8pE�s/m��5����vkN��������>�����q9�_�D6��&��N�P�1���d�HKwu�o�2\��qS���#x����x���!�`��"���Pv��WY�J��	׹����Ό3rUI���c/����T��@P�ˋ�P/��faA�`���j���m�� x�B�x�)�R`�y^�~��xKIƁt'�ؼ���y��k{Ǜ��CCg[�8ݖ�,������*�%���F*-S��%䶵�~�BƗ�)��yJ�Gݫ�cjZ�.�bUX��MNE��h7,hxh���_n�Sq��a=��h�l�"ή�yt�ٽ�(�u��b�&�b�K6��<�zцFӇ�R�����tֺ�ڧ�h�G�]]3�N���������}po�`���yr�EE��/_��τu�Aՙ���� 62pV%?��	%�xI{i�b_�ps��=m�X�`����=py�.�Dvf"�����6�����/����eоi&�4�\�'���Ɩy����e������3����	��5}߹��1N*�>6OGM�SJi0�ύ�0��`��� �<ƇbMS\�7=�O��9�0v+1�ikF��s�E��zŠ�Ec��=;�X��	-������ ?Ԓ���I�7�z�ʉ��q;<7��%�I姽��-E
�wY6b�b�yءf�
���`w���6˟�N�:Q��DQ'�BS�r~\�Ai�l�`��n�2�����x���(��7:�f��c����M�<�*����%��Q|�R�c����_���B}����דw�{A:3m��A|`@F�N�䇃n�>��1H�gF�r4�G/au_�Բ���/�jw �~�P�S3�5},�u�������׿��|���X��	��ٔ�t���HF�'.���ze2�%�(�/3R�[
߻�@����HnY5�2���C��A��l�ob܋���&S�Yr�Z��$YWnd�ܥnK��r�򔖳���]�%/ ��8���R'�}���Ɖ���tKzo��Β����	ߍ),~\<S&�Md�5��� ��]��<[l�^�L�,���Y�q�A�LA�,NLt�-�RD���'��(Oo�i=Yt�����y:�~��͔]Y4����"2�٢ȝU�x����&�p_.�Qt�dA�ZYW�/ǉ��H��\6�]�:����R� ΌG�����+!&�ڳSnT$@�>ꐆ��fN���]����3~��~��c�D��l$�:b�u���ڋ\0���P����$$�~�s����u�[�Ã�t��cjMe5��NN�U�'��C��	SL�'�\Ϣ�~�V:�Y���e�P�Np�1�L\�בW�`j_�����}�)?+�y]��O�Z^C��)X���{q��ÿ)������柚s�$�7Wүb����5���V�p� ������-M�����B	1��(iwj�Ĭx �E��P���Q�a��A�9�j1�Sjs������s_4������I����5�<r,��Vc�BΚ��$�u�$���f�;³��ÐT%c1x��y�h<ܱ逮7ԗ��Oo^��:>��Z,�C�J���6\[u�=E�Qؖ6�Ӗ�m�&�Il�:�s.�96�/�e|>l�!���,�}��=��0⼇��3$�n�]nJc�$�ӛi�F����VOs�^�+�s�R6�F|t�B؍;�2�D^�Ce����Lա�qNe�����s�9sPe���k��]	>�+ye����ӳ��!�;��1�.n�ik7=�C����G��x'���h/�)8�Ac����dp�*2য়.珧��Y�߶�N�)�,���;�bϵ:��χL�)D¹�#a!c�A�92{�m�������Gb��Uk�d��\�z��K�����(K6�;dl���."U|�� ��$����"� 	0wZG��q�x*���ޚ��Sȟ���� p���y,�bj���D�M5{�#d(ۄ?_j�M�
������8D�)�	��Z�uɓ�vΚ7���Oi������	�P`?Y�^M�F��c��90�[���w�@����.|d#[�.�IS�~Φ����!5��%q	�,'W��} �,)��w�����z���aga[�0�k�M��Q눙]!�bf��Vk�#o+K�x�l�V�����x���k	��-�D[B�>FDe4hoyg����j�1hw�����_
XL���&�r\{�In-�"�!T��"��0�v$#���31 ��m����Op>���uܮpT\L~q]�@�^s?[�1��V��+)iN�8\��9��q��Q��ىM��H�>��<"S��gs�j䶬o)PM ����T��h��oڈ��@�]i<�-/�	�t�����b6N�FT�i�F���b��XHn�8����M%nS���T�4k.S."��^�:PR�R��=�t�E*;�e�5�1��TWͲ۱F3�������('tP�c���&H���:gVϑ�����P����J�d�v'}G|h��چF�/(����U�6�����}��D�*1v9���s��T�5&��q�uu��~��q���k��#�3q�W~f�́���\�����
�@���8 �ɓ��hU�:�g�3Y.ѴقFW�y�)���:��U���d#x���eR��m�p�ʵt�#��ԔM�k��AC*�
�:�!�S~�W���y��_��^���M���+I����� �/�"�$*["^z��n e��gm��Ҿ��Ϧ�Ң~sQ�/�:�>��Y~�YR���^+��E��UcVervus�.��u~�⢴nm�_�lWo�^��|C��Fv���N"��̓���XMP�ix*ܭ��}�Lc�)d�4��F����=�>��"������^���Y��8��:U�n�[0=�̒&�"	|ɃA3,������UK��=�l\�9߫�N�5k>��}x��Wu����ὤn�����pΒ��}蚆� %��MV���Q�wQ.>QzM��J�MG� e*�?�ZQ������'N�����E	U�2J���k��6�~�M2�,Bَ���Ʃ��'���J|��Zs|{������ ۬ؖǪe-t�φ�����5�8C��c��E&Y�-�Oۑi�K����F�X�������3s|\B���]|��F��h eW�p�<��d��їA�������	��<�M�?�,2��{FrfX�F<귈�̕�^@�q��Y�mDy�:0<��C'p�|c���=[O��t��l��a׍�PY|@�E�2D��Q;���̞����ݾ�����	��ĸ��V���\<��DX�����WF���CbL"�� 8DP��
[��C-%e�]���/'
��cv�c�|�%�z�y̯�b�����1M�)a3D����7qt�yk���rY{�U�g��[�xz�p�,�}������Ɵ-L��F)1궲������Y4� {,{9�j&��[�E�.�Ӓ|H��}ec��V!S���ύ��/���Q���t@n4L�Fa�6�+���.��;}�x��ľ��J�!����'wy8:!۫R!���ʪ�=UC�Ӈmu�+֭�5U�v���� N�rH?7*�2v�-����s���H+ �m�ܴs3D�y�?J��WY�X�0�N)�!Ԓ9�o)@���!�4F�IBO��Q����r�����o���D������-6���P��`�\��͡�T���f��U>������-���)���A��'r��
28� ��d���b�c{Ƭ����
"C�kFF
ag�{e����� �U�$��츒括.��J�l�a��C��e%&���`s�T1��}_K�c�%���/�����q*�ݷq�m��9��������f���v�x�X��.�F��g�qO��q]^�E8�D�7lF����e�`0��5�7݉-A��Լ�O�a�T*��5��3�[麪�w�l��֚�ޯ�[p�B�O�&䚛ܒ}H�p����З����������@s';�g"k�Dۛ�nJ{g��3�8�G��KV��ңu�)��������z��?Ta�'�ط��s��6]K�qm�>g����oJ���oI�QY��T�r~���v�$�|ǡ��v�ÅGm>J�yN� �i�,I������Z:S �Lb�J�/�~Q[����8bY�+��tC]������g9�,yr"�5D�R{�I����0��:��ZzF��j��R�,�����4�U��}_;��=�Y��kEO"��)�mQ���)�{7D��)���N����]t�,����ce�j�F��>�=3@l�*�a^�ks�" K��n�Dè����e�7�!9�Kfz� g�/>��s[g�q�.��XJg5����R��qW%��vl�Z�x]�̓|����K�a�������Ɔ�xcS�$�|H�_r �<�-�gc���=V5*�	���!3	���Ȁc0�'�#����m+u-v�5G4՗�}�k>i$�=�~n�(����Cl,7|P��eɪ��oB�ON �ጴ	���9�t��������� ڈ=�-dp�7]/��������ù�1J#|��c�V��'��7��� �l�̅��}�	�߉��12�h߸3v��t�92Hi��('G50��Is�9����m�2#�gƵ����oLq]*(��Ye��}����e�9v`�G3�)�l����:��&G�QHƙ�*e���=%��K)���-t�03�13Ho��da��%����pM�?1x^�3p��(T���gW�4��M��5 RY�E�Bf��[?�X.���0��X�p��w��sZ#�����
���LєS���,�?Nὢ��ݕ�Bcj!�]]����c�'MM���5N�=;T>x�f��Te��5���,���I�в��&���o�q�s,�=�^jh�Z{%�U��^�jk�duT���h�L8���up���]M��o�z���YN��-�Q~"��.�f֐+�������H����G�0�>�I�0�g�h��72�*GDY�y$��{*��"�؜#��>���ByV�e���p�a����F�<熻���O��b��t��L��]L¨�Z� ��� ~�%<���g�Gb�����ӹڞ\�ªkӍ�,Kynbb�?�u��'���_~��	6��6N���Gl�e��2/y�[W`=
ЗسG��W�?�9��ӧ��#7^Ã55&�ƒ��%Y�ED���(��XC��gMU6C)]67|��<9~���&�����ǽgY�^�q�<��	�i�q�	�)�����~����L��mu�wǼ��*w%=�^�y�?T�g�+E~P�\^	��aa��D:S`�#S��Y_7�P�y��0g��HMs��oh��� ���;9���y#��6zd�����4�O�An���2Qn�kvν���n�".��C���u��"+M��gzT��/՟��8����݅�6&S�2s@#�(<Y���3�����(���(�n2Ŋ��F�X'YڇŔiJ6��(�z7%��P�萴|�k,�-���e��w�WQM�=s(�p��>��,��yROqY�Q���;�qb�`|nd-ԫ �x�����\Ж��Wx����ʴ���Y��0=�
*�ƴ�V�������Bة��/���$�hA@�P���z/)I�R}���U��q�R�Y�)j�4��Xi�q�|�%zW�lx�1���r���^��5Gfs3r�C�r,	{�o���`��[6��:����:�w;�� ��VV{�ά]<�:����k�t֧-�yg���X�3 �]�L��(P���-�]Gd]�$Ωr��J4��IB�!��L�yg4K(Y.k��6�m_��o/,�S���Wc��W-���������}��Mv�q�(�z*�co<��'9D�3�c7��I�����y����J�-�S᤬��JH�WLQڅ1���9q��YĻ�*�j�&r���^z�~]�7U#����9����6�3\�E��Ӊ�.<Hc����?������}Pq �Cٓ	��ϧoy�uх=�X�21by,���u�:S��_Z2fb1;�ߛ�o�LS�(�qݮ?�� �˝�Z;�suq�l����0�29�<5͆�b���%u��lv�3�w!J���{/�����1�Wxϯ�Y���L���h\��y��e)�!���HJ���|�
7m�'}o�2r��b3P��T�K:��g�Z���2 ���C���� ��Z]��0���1�Y=�(����a@�D�'Lr+���FQ@z�S�G}����kPX��G�����!�m�b�'�]m�l���)Ɖ�\nIퟎk�: �Y��'V���}�Oi頛��X�gP�f�N¡Y ��]0�2Ͳ��?,Ynn�tь��}����{宒�����%�{qR�B}��K*�������^�cnZ�eC���%���T�]�M���#0�lg�Z�vIA`��xo_~�e�0���N*N�Y��?�7bӂ���Oc`��J`�y̿K����~����'�IԀ-��t����:={.������17�`_�$�>��ǟ" >Kَx�n������k�Uy��?�xt�*���!9��
�	��4Js�F�Ǩ-U�������4��-��C�_Y�^I��c���!8�C��:�&_�<p;4������x���g鿺*�[���Ycd6�\�lH��ĩ�nq8���&��ϵR܍
�����yω:*[���!�c~,t%�[}��H�2��Q�0�b����Z�F�ߊqMm��LӞ�6��F�)c�ZR�Y�z���D��u�î�}��cbòwMѸsH�g�(nx��=}\NV��K^���u���8��r�#Tm�x�f�$u�era��n(x}� �)�P�FwU�'7��j���Np���^�{[�WK�d�����Z����W�aPf�&�gz�����im�1�`ab�<>�iDpD0@���ߗ�[��y���L�#������� �,L<�{*���Ȫ�EF�k��As�������]%�_�?Y�ib4қo���Ȧ�}I��00�ޔ(��̄2��G`�_ƿ�I����w�[%p����#�`Z@�@%�ydb9�R�LL�����ԫ��w?���ى�@Jؒs�\��3-:����H֚E+���W��b�V��X�p��D�3�C�Q���{��o �~/3;KL���
�l�AL?���o}�E�]����P�4��G`[~���S�%��/W�;�llkb�M m��~���ڷ���UFu���l�f���=�ۧ�7	���~(
h�JիK�ε�]g��F8ES%]W,����7?w�i�k�N��IO
Q������
�.���0�+�k���"�# �Fb�Qd�<E�,Y����6�_��_�d�2M��,q͆A��Y0ÚЀ�yv�Ǫ]���cp:�����l��������%w�,�������lrR�9d�y�ƋKq$^��ƃ���y���m�a��B����]�kn�p�a�Ԁr[�����!�k�*���W6�D>/��z���U���ۉB���<LT��@v���J[���w��c���<�F��2�d��y'��n�=5�]a.k)i)~�X�i�W�L�;�����e؎�"�1"^������X��QP&�k ��U��Ϝ$�l[l\V/{%Ss��z%�^����ے�s�_�&�&�?����x��ET��FvW�����I�8�A*N)�*a���$�
���Y���8cf-o�e�U���&��Ӣ~Z2kI�ځ#�E�I�a�f ]Ǫ��Eq���,\���%x�ʥ��l�V�:�q2�ê��O�ɱ��<�-��������i�x�z5���J�4�s��Vx�;ǊF�!��
,���>�MOʯ�1=(��`zT��mF��)w瓟��u�\~�J���C�R�$�KIj�%)l�	t��Nc�2�R2���D�id����vݤ���?��+'��Cx�X{b�kH�R��u�ܰ������N�a�2�����U�U�,���5�~�S�'�oШ��e�r̖��b~tW�(�"�N}���(���d�7��� �����O�̴���V.4��N�.������:Nlyr�h�a�C���'ao��5�ԥ���U7�ڊǐ&/_�s'�&W+#m�������T�{�)���C�������]j��p�H�9�t<��XMI?�sR3f�@6�l]�8��"��HW�|��]ROܶb�G�Y]Q��J�sjA���p���JN_Df	|�
>ۿ���.m4������qXH��P����b"�ڡP�|V�aHVC\c�xS��Ј(�l��)J���#7���?��C�*fe�U�k�@jb��-wh�D ��@j��e�9��tv���s��#��p��>>ׇ����)߇�}��G���S�I��]׶��Yk1Gr�~�N^�I�#]]�!��Q]�bQ�s8���U8C���{��>�]eM^���8���"7�AR��.p�<�`����B�<̍}�5ͺ.�d�j��E�����'���YҘ��zb�M��X�
����_�V�ŔKqԳ��8��\������ό+������~���?�w��R,�ٰK�5��7�g����t�M�w�./�o~�'mY���8K\�d���
�z*�:�bP��'��s-��U^X��K#b�`�ճ���t[��M�x1>�fO�l1��i�`������/)A�yʉ�T��1����u�����i[����*/����Z#�봮O�a"����gH�w)u�5�x*�eN�HӸ������8��pw?��t(��UA��L�����d�k ����j�����lӿPj���ee3�
\2h1O	?P��,C�|'w��M��J��R�#Pm��t~.�xnܿ9h�8}��q�)�m��]�K�������f���xm47'N{��!���jXԱXWNn`�k��b�e��FW��:�˲}��&ovi�*��U��&�sQ*,牧ć�Q�ha�o��&���	�D��7Yc�,��tlD�fF������S�j+R�jE��-$S=TsĹ����Z��"46��Z����)�����k����0dh����h�ΐ�)V�oEO�Cc/�t���j�y��]r4:bzC[����TR�ԇ���dg�A��UV�t&R��(a�{��̲ٛ��>{�*�ߋ�*��Z��/���E}�Nr<���m�X�&q �(��:��X�Sx��D����쬥�\�ɽ\D�fFG��1�8k'6�>��cs���(0jX	>�! ��ĕ;�}~�T���C���}X�D�T�q��@�A��ns������|���^�/�4PP���Ú�&2<�ږu�W`���^Z�.?�f�������� ��]��-�rW�g`�θ���w%2�k>h��2�a�`�l$����`��qC��2Q1E�WF{e_^}�*��u88���Xo�{۔"�m.)u��)YJt8�v'N�9лX���������Y�Mwc��}��X쇏O��e�y�Uq��t$9��o;���EE����Eж)`4���ܳt#��%�y��Z!���5WAN�v�xe3��E�R���hU��ߥJ�nO�V����Y�M5pƢ�^��1�c��ʢ�()�HǓ��5��>��H��Y:��s�~z��3(���(D�Z��}��q�����ݗ[�$k�!:�8�&�`U���LW���9�����e�Oz^��k<�O�q�ef��S�!ba��9i������ԫ�;��4��x-v�<���&��@:���� ��r��ޗ������z�5��$�'���0#E�����/�����:�0!<n�퍦�������qz�e�8&lT{5�h#�����5�Lt�T�������Q�ӝ���CE�A�\`po�P�!��Ə��!-L�`-��t�ꉍ>�E8>ዧ8���D����7��OMD0މ������`X�`������ډ�=%o�R3�z����[�j#Jr�Hh@�����`^V1�ԅ��Q"q��`�m�߷���x�1����}�}��۷��{X픊sR��^m�d�е���O�ʙ-5u��R�\���l|�^�oRӵ�V쵴��~�|V�	�V+�꥾�71���')�#�a�C��Ol�ڢ�7B��ISLL�O�Q������� ��)�mh����G� 5  ��IDAT	^Sd���F�M �Y\He��6��I���-'��1!�R_�\��S<���R�r��ט��A��+NHϥ�4�Eg�*�k|����:�4G�e�1��L�ϊlP�AI'�5,�JB��M9F�́�q;�t`=wqm�����z����- �������=J=dJ���C�,6���H�(�	�\Dy+HCa�0�L�x����d�>3��f߱y�M���-y����]/���`p
=�s_���~��.�i����G��Vb�Zi� ��1��A$24��b+�*����?��m|a�ʥ)����Ǟ��ڴi ���E�A\'��Q;a����i�m>�����ѕ?s ��ڼ�ɫ�Hp	2��I*\?��KE]��V_��?Pa�aKt���m��Sy����*Û�<j�ǌ��
��ګ�޿��s�>m^��m���x�-�F�����s6��:�Ns�0�����e_GILi����H�h��_�[�?����@c�I�-ʗO����٢	R;]#��/��fJ����^�	���+�G�+�%�Q:~�q�[��ĉ����xi_5%�6���Y�N�˙����]], �;��o��6��(�K�i�>	��2��D�x���d:F&�H�Sb��-��2���TEo�p>q�N�!1Y�g�)�14������0�l�t���(o8�8M�j�p��%��.�|�F��Lq�LL>S���X��|��>%��<k��Xօ����I��E;��ê`@����.��9����E��^�����DzT6$����t����Lb$wj�-�Mۢ��++%�J�/����d�;a/r%e��^�mr�l��������L8��E��F��:����`HЩD�d�5G[����T���qLq��p/=�E��������q�Gx|ٱ�oŴ��r)^�m�/p�_�ڋ)p�P�jl��%��R�� ��R8���j�Zd�7H`w�����JH<<_k=Ã�΍{����iG��Y�����h����$,u��u�����\Q>7�`���HM�5�M��N/��>�M�����:��3�[���>?���C�IZrz��0率Es����.ͨecu��Hl�����3�{�,]zL��K�MJ�kSw���a���CvAd�;
N�Y#K�i��r�DO� �l����(--Z_����q��*��~�1X�+�e���HOaZؘ��o�5Ґ ��4�C&�;I_A::&�XL<q��<�GE���U��k�O�W/�
kV�R�$�"!���k��<o���"XU��Ś����R�=��,����T<8�Pa%
O�J����޽$)/a.�XJ#x�^�l��\�X��ٶo^w��_DÊp��g0]�;�M�+���)s�Y\����*�A���BV$jtDC�H�	�(j �͜���%j'n��頎	s���dZ⦂f�O�)G�tc��}N?�A����^�/ys���7���Ep��7��[sY�=�F�Z��s�|�m����])=�s'g�5pa����g�">#-"�7��%�\��>��=��J6Ѱ�������'�"�}���کn)[��4�]Uq���E�-6c�ٿ&��A��C6(Hў�H1��C�!��agmh
2s�u{ߏ�����A,���S'`Vއg���]��G ��gk�Ȇ�t�v�fmd���[�9 lf�ގ�֬�Q��!�9#��l�K�ci����&&��� u��Ab�(zē�y�C/}�k� �~�,~)�St�������`Gׇ��q�����'T�W������ �F6��t�i��=s�ڪ�NZ���՚0v�lB�mH}��'�O�P_k��]y��S0AO¤�v�M��RC�y��.��$�������u�q�`S��g�X5I�'x>W�x<�Si|��'[sAr���#�*�ʖC�Z�f��cs<.�����)�!]Nu���|O}�m�W9���l��z���7ӕܵ�'�j�.�7a�K(�LoGs/�0"(7��"3��1_#��m��,�ρ�⑬�ރU�>(AӮ�ǋ��a�Z�k=���2�t�j��@<���m1	���;&�]y���XZ�YC"� �*{@�k�k�3�7�x�q�f�*�f�U=]VD�F��	�??���[������`K��霊����ݼa����7T�f]r�ɴQ�Y�` W1���9j�H\����0�ڳ�y�V�Z�L����{!����57�+�����ӛG�A\�_�(�������`j�%P-�'���aS�!�o����]k�� ެ\ܖֳ琝��k�g!t{�w�qp�eR-s��|J��6��u��J@��sww���Tw��pUL����.9��r��4������ڭ�"���V!���i������U�RZX���р��m��K�MO����,���SZ������&��d�¡<��kX�����	6V��8^/wJ��Q���q�M�_�
��ŋ�j%=�"���)pT��=]Yj_��C�"�F�GRK��Jd��ķty�gt�CZ9Q��9�����
g�]���˿j��[s_}��$�������Q��#@]��7�HI�qow����5�X�`�$���I�������:S.�/_�G�ş�n�'ۉ~[B����p���?7��.4#qmrXik�y�����&`:1��m~���u�p���6�������]�J6wv��w*]�A�oE��+	���fVZ�fv��T`b�B�o�<�Z�-��ɥQ�m��>�ΰ7	��^gެ�����luLӺ���%��?�`�T�J)�����i��*л�,(��+Ŗ)z�u�nndZ��l�V��Y';a����(Hm<3�~��g����{�oF0ؾ��tv
��X�ȱ��'��F~�Lai��p�D_+(�
��yӣVm���X+�<��G�[յ�'_ه]`�=7`��t	 ��p�D��*Y�'�a�N �7�0Q	����I��R15�G7�܀�RW�1�0h�cА�S)��s�YbIݣy�k�uy|k>?���T�5��1ڄQ�
�#K��XFYu�9���$��ꃲq7&��ڍ٠�m��1�/���t�F��ʪ�z����xc�x%�5���ᜐ�ݘ\����9���r��$�ȣ������TF��v�l�V1.�,���*94��te�74���J��������^��s9w��t����W'��A����z>��6�|7�P��(3����P;��1o.��8�!��Y���^�*�d6���N�}yj%���BG@�ٷ��	������m
������'q��]��sQ�Y[ܼ2���`�eł�<[a��swS��
���*9b{w(�Hw��>�
R�}�;�g�w�}�J�v�p�9⹦���	�u9�ɘT������-uD��U\�yݾ\�.iHǁ?Uy|����#�R�.�a8�IUת�׈�,�Y�S�@�k-��jXثѺ�yz�3���Um��;��!�?w��w4�f��yNۏǇ���|E��ӾIF.�}SԦSt
]�=�}�;Á.F����)!�Q�~c��X^{�S(�km}�H^�y=i DM����H}M��q�`ɉ
N��~�m$�amgt^� �K�D��P I���-Z+��Sץ[�������Q�������/�pnbg�}�6��QJ)!�i� e�xMa��d5�>_dB�[V��U'���(KZ[��V���f�Vu�yqm��]䎚���Ȓ,�#��]�{M�8�a�3Ŷ�m��n��=qPA� ��"� ƍ�[Ux�)[)J�
����c1gXI�Wf��[�y�"�^�o�A�
������u��׊�z�; B3����%��/[Y��?��C�x ��d���*rb?����'���A�G�B2�p_��[ ,�5�F������Wb�%�X�b$���Q� ��b7��z?d�Up�J�{W�d���O�R�/\W�w0�u�8�� {`�>�i���,?��Lj�]��D�l
[ʜ��I;د`>��Vގ�_���н�#/��}:�q ۵�������0P<)�}&a�!�rܒ��>�~�]~�q���?,E��.�;��D�"u��0�e�*Y9I���p��r4������>�e�M�]�6�fl-c��_���&Z�hJx>w�)�f�)𬡿��A�`Q�+�j0���Z�Ɲ��͙�婸�'�ɹ}a�n����9u*�i6����N����������st�n�.�\�x�x�j+k+[XN��!i&�5�:ϵ̟ĵ���7uU0^8���ڭ�nO �}����6�o˻�]V�p�8Y�J�Rljt�@�Q9�|���-0�\���T�m���O?FF���p���^X������s����&!�B�P��k�D_����O�7�f����b�Ŝ�MHn���� z>�����JC�mnl�Xo��s����b�n�1i��
�P��S�Ӌt
�')�6��a�Ǜ�M��%�?����㚮N8@�y��6�Sd��>~J?,�����
E~�ݧV/1 �/QN��Z��}���~/���EAu�W�����'�8FK��,J!~�z��.�Տ�fS�W.&�T)�hjO�����
�u��Y�ˌ�-z��Xe�~>-*�FM}36��{��fZ].�1��>yr��k�	,��E �\Hӫ��݈����>ˎᄾ�&�z`O�4uEϘ�Խ�<�&�sc�,23�̀l6Tp�`E�<��]������M���{�m��u?cwK;����i���	QU��x�)�����u�^bSQ5�$��.&@�x�{��n�O�yx��<d_#��o��~��~_|~���!s�����M�Ʉv*^�I��*��ľ�����35��b`|�5���o��\�&͊����@�,>!���n<�����3���#&{`���2U\˷o����TXz��Y�k��ÞSZ��m��)(;8�4�瓦Ӱ��7XcȲP�L0G���n�0�lf�����a��E���D6y2�������a�,�|Tew�:�Q��@1����i�K�®�ʎ�h$>߳rz�5q�fAO�%��z̓��.5s/��И�\�jm�����6��ܟn1uM�%|���������GПn"q)�/��V�hF-�B�tSd�^*��x� �T_{=�ʟu���S�x�{\,f�]_��3���m��e�,_���#�)�3�":�/�RO`�E�!'�,K	7�,J[�ܐ����@�B� �cO�)��Ź}R�P:���L1Ϣ�U�I�ua�g%ot��a�w?�9����/[v�6:��;'���ӗ��Fr����*���ڟ5]��<1����ǂ�츯JE��K	6&�N�n?1����{���"5�"j�7iR��]4��"7C������H�Z����
ig�O���z�������J̞�7d7<��������'�E;�����[~$��]6ȴO;7<�z�h(�ؠ^���?�i��a=��0��-��J�.�����"\9'��p=�	`�׊UcPв��ġ'!��f1z%�o!�u�>�F���ե�]���3��&�2��^Mm6uk�d닧k���,j2�f_�/��N�d*nTi�ɦ��=e��P'�i8�+�����^䦌1C�����@
��G
Q�Q�#nW-̢�g?����\2��-���3&7�,eJަ'JL�vy�bR�|�����uRC�J�r����fѥH'����)'��^p�~�2Od����lY�w�G�hm�^b6����"�� ��π����ӖA��e���a���6�����%�^)��Xcl&|6yQ�f����s�����ރ����n��.�q{����fc�iCB<��u�:Y�<s��lBxw���	�p�wm3��f�+�%�5�O�/xN��}��`-,U����E�pW�x��	����x/�X�����~��Q�@�b�7ؠ5�t��r�l.}�w��Ĕv({�[���������l����{�j^>�]���R9n�#�{�`��U!�]�MתlFiF�����|�Yέ��YX]���/�ￌz7�$�B�ڶ�?۵ߩ[�ܯϩ�khG�T'Tz���Hh�p�[E��m��O[��_`$
�]g�P�]��R�Z+	7��,w9�rUV�At���q�o��J1��e̐Ap�q����n��(����,�8���U��Ͳ�16�Z���lnL���\No��0�B�m��+c`˜��i'R`���}���{L�(K
`{���ͷ�_~�;��?�xf&�X/vJB������@*�
oW(�qw�4틦�0�P�W�!h��-d�߼�ύ��Γ���Aim�*���`�]�>�uұ,Z�/��U��Ն�>x
�*a���*�����?�@���x���Qe)uvEÁ���92�����w���=����tR�.�sL���������Il���	���[��C"5w�믾�����Qڢ#�E��V3�[O�S܀q�|�z��ob?5j�^?��C�,�	;�׋�dM79բ3v�2Z����ٻ܍m��_���z�W�F��qõ�t}Ѯ*�	�E��Q�^2W������c���0�2f�j��^��K�ِ.�J/�z����Ew�d`���U�X�OR����.,8��l����	��5��No_�,d,��"��̪H�#J��(�հ�8�7�F;�-���U5��q�<Q�x��
6�n��)��.T�a_�^���?�#.�k=����o[����_q���[��t�9@�~�6۫mc�wU�8J��:�����|�!����|�Y`��j1���M�nZ4�ο�Md�x��<�(O�E
��]b6��.�A�{��ꫯc#c�;$��8�������zl���b]�?�R��_�5��-����)2((ɿ�2�����L�5��k��w����ۧ�I��z�a��!A��t.�8(��:2q��ή��)��&�(Q�q{��"[�5�z�H�N���]V�=�P[l���5�kb�j��"�w����aOS!��OмA�mQ��̙,�E�=hdMw��XsQÉ@��v_�i4��Ϧ{wP_ƾ��* Lsf�)р�����Í闻�]ߗJ���ӑu�j�n`���;a%�P=qH�K��dR�-�N�xl��a|-R��_E@�3e�3�V�1%�ジ�����X��C?gwݣ��i�baFᙶ�-�#���U\�*(;7�c`�w�T�!efMz�$�<Oq_�B�e �Q�W<�Ο߿���6���xV����#2����|z��#}��J���x~Fऊ=՗Ne�5B@C)�k�$K
NBu�^���Np��k���t)_lb�Mɹ��E�W�/)}]�d����j���(��c��d�i3�h`^N�\����|���=l)+�g�HMX�S#��z��^���}�h'��vYk��pN�`#�pܫx�ۡx�2ЀKcWf���7����L���}a��C��ￋ���UQ/��k	�z��7�07=!���}� S�I�S;�p��Ly����VIڟ�����[vѱ)�����d�	r�L0���6��4�Y��_wg���x�~����� ̆JrY^T!h������R
���b3��e���Sj=�\\D�GK��b�=E	q���~'�5�p���<�<�1�Z6A�@���Ӯx��oP�N� �62Y({��נx3N�sNjy.�ﰫ�D��u�A�Rg��w,/m(f���l&��>||��ݲ#v�?
���|M�"6��A"���2X¿�Cv��{U��&.8O[6����p|f`��`�~ձ����3�ٳ�:�p�m�L�@�����Dbp.UbF�NtW;ĤwA��m��u]��X�r��"h6@���B�Tk�A�*=�):�o�w[�AV�a5|�; ��Hm�v���h���!��������Y�a�^�D[��{�0̼�z�a5���D Fј�� "@聆�Y�^q�~��|��)��Coù)��A�l�3���>M�q�p݂
6ŶP�>�R������ �� .k5����1�`۶SA-�?���1�k	��OR���w*N�����ڑ=g��X*���P8����ӣ�蚓�4��r�j_.RohX���)��Q�`�6
6��\(�_F���������2#e&cJw��)�X=i��2�cv�俍��",��C]�mV;
|.�aR�n�˭�3ϝ�Jc=}p|.��i�;DV�L	e��ۿ���r	e��X���:�����E��.=�)�Q���D߲�k|�����T��LB@�1�Y]PT)����<����	��.
�,	^��$|��7�o����r��n/�Fb�'��N��|X�zT�x�*�N��wB�8�8W�Ԁ�&����������m�\�k�(%��c��~�z��m������` %���5<���c`�j[�d�����x0�0�n�s��8 0O�*�q=�1�yA	��{{>H㿷l4���U���N��%F}��p��Ʒd`�վ���E�9�l��lR���RӕU{$x��$N������Ju���}��|[/M��30�����f���㒳WL�#��X]��Km�1T���rYʈ1��:ҕ�������Uc�&"⢮jRQ�T7W���Y�F�j|`q,���]0��sGv2HA���k&Y)ksP�e�.���]�T[�Uԑn�%S���?���ߛ/�����+���ۻ��R�%�_\[�v�8�vsF06Nk�P��+�2p����r�2�̗@G�ཱhd>�n��K��Zm-'��)�WB�����<<�.�ؠ47zh?lPuy�өD�Ͷ(+�	{A������,�ל�_T��`����١�I��ڮ�!�V��t�Yz,_H�k� ���w�Q�f��z�_"��p�9{�MơK�cP���؜��2�iIkp��i���h"p��X�n�����iX�s6ׅ+��x��:����g�J+�e͉HŢ�T�\�2���jx�Zm6��M�|���"֟��V�cMN�^�-U�,��q�q��L���h�{��j�sN7���ܔ(�/�8�x�g��6���5&ya�nj���|�%�{u��n��tΟ娤����[L���@5�벋K"8a��I�]�����#����e�k!X� �ed��6=�6��^vc�F%����5t�����K���6�,͝��]�cC�(+ab�U"�bN�@}ZUle������'2�!�����\� /��&���(�l�5��k�X�/���Ы�#�f,l�����#1�=�{O>dۋ��Ş�C���E�2r���Z��l�H�S\h�E��}j�_�f�E���6ꟺ�]��X�rL���^:���Ս�OŴY�ly�B�K*�]�`���S���љ��D6�6�qJ�>�*qx�(�r�حu6������r�솲��T��p�(�X�nn_�٬nGu=�W���5K����7׼��������u�n:B�{X��xϨC8!� '*� �`���A�V�0��ӧ���Y�2�_0���s�i��(b��Aa�=�씁Ya!<iƅ�7�K~cCbZQ���4��Ih����7ю$9�E#3k�{O���CJ��wλ��9W�<Q��z�7 ������<�0=$������%3�����L߱ #�>�w<�B�S����d����NDK�ÀGv�d7ު[��(dX��P�Xhr �C&����$�c�Nоk����W4�۳��谡�� 8��9\O��ht�6�X �J���C�KN�PN�<�1�.w돇��b��ذZ���8Y~�����EƎO
�5�3��Ø���|�1����|��؉����z��vbw����T��	��:��DUB]Tf[��K����f�����iy�h�����8hl�eiOtV��!�@�=u�sm��$�q`R�gO�ym�j
+�C5�;�
�n����3��r6�v#�6G�T�fuФ��&�⋲Y7�fą{2nv��MU(n�!"WY�?�L1��ǛH��@����`�����E|Avϐ�?�P�?j�����.8k�M���P_ҁt�>̱h�z䍴C���a��
]vR�A�:���o��?|ҬnH��[*��6�b��R/�es��ڶ�F �ȭ�f�{s8~҄�j'�M�x^Q�Dt2�Gd�UB�R�5\�)����ԛ�k��Y�����?��%9�QHZ4�����p8V)V�>�+�oKd�;�.tW��ͫ�Ff�(�� �h8İ16y�1��㬌%~�y�M"d&G���Ģ�<�#��>��͇���q�{T��CJ�J��ðո�a]���\B�*��!(2��Ngf�񾩠u,��H���^M�C[���A��Fad�de��۞����o�C.|b���v��Mu�C2�Rk`g�j�w8�=��ڧmTV1ew)w9���5�N���:^3���Q����Qb�$�A��7�6�.5#�Vq��gU��=j�ڕχ�_��o���Ɏ�J�Ƙ4�|=n$2P�a�	!z�Vb��4Y���XbQ���=�8�R�l.*$��.F��领������������&ZB_�4��l՚b�����gYJXޫ�l-�R�c�AM'c���u��5��>�B!0�y�V����:lrlp�����X]<������R��G�td馋��X4��f��(.���#��`"F^�)���]?�Sp'�/���u��j̹���M��eנZ��w4Sb�(���QNs�F�
���fW����F�7ŭ-s(K���������c�gk ��g-�{�/r/�(9�;k]��6}/qg��r���%9���X�?��l�c\ҜKVg⃚�2�\�ݸ	Z��%�h��kZ��'�s�	�j<z_�t�����Ic�]�WafM�7�pC������^������ߖ�7��9��nU�z,�r�V0d��Hz(/�gW��M#s4©q�Ձ4n�^&���c�8���T����}��c�F'�P.k/�m�rմ=߷�X��L�7[(�x�0 ��6��w�'�:�J3)s�C�$����U���S����F��]�ߛ���c��G�C8C���*��3� �C��oR�d+p��9v��60o\�,c��R��ﾥ�݇��s�c��� �g6�� ��$��M(�S�h�/��uw/\s��Z��*�ۊ�wS�z�%�~���r�4��'��>����ȵ��-J�p��47��S-�"��@�m`n��=��cm��������H�5B��-��.��)�*��~�<e\�,I�lhv9gm8���xT�h��(���w_S欁Wh�e�z�s� ��oO_�}�&1�V�~=2Ƒ���e�L-�~���2?[�ڨ��\�w;5w�`N�B6	o���|������ÒSCn������9E�e��{H�Wd(t�
��}��x˦�w\����h()�6����_H7a����Y_Y*��iX�B�K9K��Q6�e���'��;�usOLg+������	�M�&�Κ�~�,�e��*�X1� ����ÚA�Sey�'�1�>R�!}Ĳ�'kX�X��Y��s����h !As��_]˹�{��)>[��O?��֌�6p�;M��WJY�V�tN�/2t\L��$�U%0���"3��AH���[`�a6�@�d�O�<*Ϟ>-���M��������3�A���~����π��F��&�s�w��|�}h&X.��/��%��@%��>>��{��A�+X�杂���q�b��vǻnІ\�!�Ɖ���X�Ҕ�U=�،,:ܢ����m\[�W_��������睆���3���@������YD����yZ��2g�N	%`�Ą����p�sɕ��7K�����A�SO�4��ݡ�<#�\o��g��˽Q�E��n��Y�y)3��B�����,�Stq0Y��*l����&|>�C�!���`j������?i����(�R��ϧ�X"�Z	_��Џ��y�.�Dʹn�,���xe����Fą|�_/@)h4�ɡ�XĿ����{)��<��v�et�n���>%�9��l*.X'���7���?V�aY��`��b��2��Y�H�G����	���C6ъl���FZ)��B�&1�N��^B��ll-q?}�{ALmmD}	O����l��gO���E�$�6�IuX޽�	� �k6<n�a�!NǊX�Zij�E�7�1��͖<�	�������/��v8D���(�Ŀ'����c�y�IC?����Ա	u�g�|&��)�m��K���t<7��`:)W�I��7���>]�׫�_�#hg�z麰h"K�S����*~I����Rg������ù�?��[�3�+�cվ �����~���"�B�J�]�hJT1Ux��R����H♋���%�D�K-��n��E��Yg>U�����b�F�m$�HU],�p�u��d)�v���z�u� �����>��V���qf�2O���b�*���F��g,��E᱐��-�E|�-躼�g� �H&-e�$<A��{[;l�Re�Ɉ��{���}p��$Tsv���)өx�')t=o��=�Y��k��G�m���ML
�6���	%=�(�G��麰��v��-�����v׌�~�O�3��[v�����>ǎ/Sm�13�K�4���}����1$W*��X�g���a��1;~��gF�����Ԯ�+�ހ�4Z�lf�Z?K�n��(��Z�;$���u��&�mjq�.%Thd�|�Y8�r4佮����V����B1J��vw%���8���?����L��hr!���a��3������;��y���w�{M{Q)i�E��s�g�"`�:�t� ��a�����b���J�䶻ٕP�?P\z�v�Kw��g=��?���!D�R��b�@��7�Tļ�QĦ�hsd֎؟��N������p���kz���G� 3���HUM����d`��m�D^ه%�\��Py�.$�̙�R�w/1b��\8sb�f����8!��Ky.�������i�����I4v_�ad}�p�ߒc��	ܰ�G�BMPY^ pK�h<�shd����HѵݪQ������D���e2�=�HnEa�/��,�}���0Y�vn�D��Z%>#^Rp�n�BG�:s�JA��=��~���0�=-�vni��N|�L�:��B��Ӈhsؽ�4���\0Zږ�KO�9]�s�Sv��=w>�PD���;+(I���n����piX��k��k��'v�q���5l�6���B��Z[��n�Q!���/2r��b�������_��G�����e(�c�^��������!~_�v�i��s��Md�����P�f<M�Wؕ���S̷wwj����ǠL	�G;�)�c�;��\�pЙ�=(���Um�����:5c����<�0l�Tk�>ۨ�[ԅ�8��N���*T����}�4`�Ue�ӹ��I'h���:9L�wY�.�F��`����/^����g0%�l��:j9��k��MR<�u�,�JݻP�	%`�&��>���l��{�WY��և]��Ԭt�RŀxP����}��-��	����������&��M_���YVx��M(0 ��<)>"{�$�9�_�SlX����wi͸33`Sd�MW��������zp�9:e��	Zo��p}�P�qg�Nt����!xS ��.5
̷�1�m�m�|���tW���1�d6�%�6I�Sf������GXM�< '��x��,��s���K=O��R#�K�5S���g�d渎��?�@�=9�g)���i�Ǡ��x���)�^�l�^���+: �b�ؕ6&���%�����g6c�	B��uo8v}�f���'��7q�=�)��"x� ��W������/^�(1hpu��.�MQ���*^Nh�Q�c����6!ei���HC?�c�]�}o9�~��� �g�45rI��W�:6f����,�ur�� ���&5+���(�X��(w�47����3���/_ds+�����R�+��Rxc4�i��E7~�QjQ]�T(�ww,c�\�ww���U*�7�Xh\�`&��6G,����꤉[�x�	��g��[�5g|��^�%�]c���L�b���W���^W�om9d7Urx���H����3��k�t���h{��F>赳���HP�ر�?!SY���J{��c�n&��]�hVp8a<�ɸ�\��$b��]V+�0o3 �����f�4-�:�*�+Wpz'�Ų�F�m}B��Pz2�g&֏&�u(�o�xS���-n<+Q���|�*`Ff��^6�P����J!3�����`d�\�}�O�eC~��s��k���̻�Ae��rKxL�o�344�!���C�5����R��*̎V��Ϝ���:`�~���z]줳0H��s�6�.�qU�jB8`Uéݯ��{!�ll%~�y���(�q$�l�&g?�JZd����|BA���L���d+9@:�� B��(����8k�T���Rl_�vspc�_9��t4���|�HR~�9Wou��Ʋ}u��.��.}32WR�$:�S�~o�a =K	����Pa��.�MOR8���4�(p�f΀\,���G7������QY@�w�[7Y6/uY A�~�f�xc�d��,�4�	b��c<�f]���#˾��d9�Zt U�z���^��%���a9�VSI^g�7�s;Kt���(��ʔֳ(�(�}�9d������pד�QyD�����NA�_�i�u�
hx<y�a���<[��ω1�9gґ�W��T<2"�F�ac���	`'컠Z�M�����JW�NT����۸߸�'�y�n+��C��D���b��Rg��\q,j��M�Pe�*4�Խ�,5;]�b�a>���T���Hu��(܋��S�vRL	��:5Mw�%�N�ࢮB�Į��(�������1.^�yB���M�v�,�=B���=����5M�����l���C���M�2�� ۊ����ڜ��ח��X���!�Z%f1HGI��}�m(N����*��o�r�� ��%e}�w��#@�x�Ic��3);C"�H�BQR�y���^fv�1~x�y��h����������85��[Q�(���݊wh�9y���p��}��]����e��C% ��jpѼ]dn�y �� l/��
�F��V/\�̈́M���FMf�&�/<��n#�RO��c`7z��u���U�c����
�	K����C��7ڡEם�ߓƅ�?���i�_8짳�n�����r���^��� L��G�5D��Z�8XE5 �>��{��)��5�͈�+�n���t#��Ŭ�gQ���H�g�L���A@��R��|��Wc�u�Ր*�g��t�����z�Χ|5��}��r
qW<6�4�P�C�bbsb �v��nI�ߙ2��꨹�����K�rf���S�(�6�)ox{�`!ͱ�lK˃B��i�ԣ.w_����M��h3ITy�3M�þ��,_O	�6�w`H��ρ&'y�!�V&�/\i���G&#{����'�ի��A��p���m���P^፦�n]��ۻ�Qڨm<�T BWl/�U���3��!>�b�Ae#&0�u3�����m���9N�,ߙ��I]�K2�.��rWt]�8ƽ�^���N�D����*�Z��Z����m�g�� *!�!=��Z�R@�k�M�e�,/����6�9���%6XS�g77�ym��9�]��68�>4��OЮ6�R�~b��2��S@v��E��^C1�2���@X�K%�{u9�{}���"�hL�-D�Ў�me�
�AF���.�b����ܴ�3]���YĪO�yh���YЕ%��(K�H�3�C��f�U�ߔS��%�����NQ��Xv��jJa}Se��ϐZ�.�p9c��,V�mCa9=�}�$��ӔN�'3��/���)��d�E��bj�T2���\S��Y{L
K6/VâL�����Ds�]�wG鞁�/v�?����͵tfO�u5���j݈��Az}}�g�I��)-����������w4æ�"'�M�&�څ�!�f_~��m�@7��:o�f�����6�:;5\c�a�6g��:H�8�K�7�ᖓ\}4~>���qL��>⳾y�[��qu5bb|r#�{�8��?�:l4���r���J�����B�O����X��>|���I���As�7�ٓ�Gu��F�-�	c�8��䣧4�]�7�r*`�����^�&����C�'��/g�Kf���))KV|@�^��/T��R�9��� <���.#�΢-���2��w0�	�E`�Qf�S�R��{�]~<B]���?-
�]��@��j�f���S��n����e��L�0��'<Sq������fϕ�˰>�#��S�����`����HK5�S��2��A�%-'��M	8Z���r��R ���Gj��8Mvs��'�n���7�������tNz���;��Ca���{c����"��j�K��%�L`ӝkL�B����\��֌�w=�/�����b,����̒ڸ����[�LJ4B'�x��,�*Q�;���~TOذ}��9�^�~!�?��/囿�����i�ɣ���p������t߃���Ǖ@������{��2t =���Jg��8�9Q%/3�ޟ[�qg;p䰏��F�9V]�O&�\�dD��h޵��o��v�`Y.��5(w�/���b]�+ي)=�H{(1�βL��M5��bx��y��nZ�K.Y��U�,`�]LS�"8-��j>U0vٸ���٨9��n��є�Y�o�UF�;
���}��7�^u��9�Ug��-P�}8\��V�y����5pg�hbB�g�{�)}�%���5W�ì��f����aϧ-���1�v�̀�,��O��M|��q��W�^�R�����Ϋ&Y��D���Y�؅���b�e�*��s�Tj���%p녝�+}�����e����_�9��u;��?7��Z�8�`z�_+�6���*�_g�
�#�#�Ӓ������`�}h<���~�e���_�Z��7�Y������'�'���cܛKV>�$��4G|؈�Bh��u�����|x���Pw�k4,�܌�S��9`2$���j�S$1c2]�خƲUV�m�͗N0��i�6����T�.�e����^}X�����]{���\�I�n�@��]�Ml�5� ���4�"�&y�Ys��[�s�k{v�%48l.�-j����i07�qHuO>8�59�z���T!���%��=y���"�kP�%q��4��<Ņ�Qhӫ�b�,�>�|b��C�$W�<���ܙ���!7��Ce��I�T��C*�Ҿx����sgM�HՈ�����8*�o��#)R�&E�!�ls�!4*����8�1�J3�T�yiǏ��Qz��� 泇L�w�]�p^Nw���J֕��D�r_��뻒S}ь�T��G�ݒ��xF�{'�Q������7>:
�e�i+^i�R��'�t'd|�ʗ	���o��a�~�͟yݠ��� ���͎A)o�(��sG5r�.�Ȉ8�ޡ�Ϻ.0m���O�hl6�3�������pfR�u��aY4�s]�>�u�kI %Ľ������� ���ڔ`���U_<;ۢ��P�3�濐���P�YQ��n����\����]�t�$.�L2p�%��2��O��mb}!��w���m%�jb9����y�/������&��R�?gg��O(=�|Hl22B`R]�8��a�?��}��;�����D}�$1S��Rms��1s]�q�\ͪ��m+̲D�U�T���f����Ec�t%�M/5�א��o� ��a8�S�^\_�0*�]���hT�rR�'�{`��:S�:�m�+iX$"(4��I���n�θ��c�9�.�;�6s ups��o$�k��h�o|F����ld���`,��5�h$%�ˈ�3�E���C�~������R����@L8t�˗_~������4�"��S}-٢��ؔ��@zT���� ������勗���/ʣ�O��n���gR9\�/��V�����p?��B����ϼ�e�����錴�-�PT����k0������h����l�T�J�D��_f��T̨�����0A�_�Li��XpΜ�X/"���挟 x߬������{����Qx�=ţI�x�q�)T�?�z�)$3��]t�,PHǅ��qf��lsdh5#��jg:���9("�.��B
�׆Ї�.?�9�uJ%*o�!̬b"]<��b?�>KEV�'�'%�Ɨ���j�&��h�񉮘��F�S�L)�7.^i2�R����3�E�n��5r�������
b'�BLnͲȰ��6�.J>褶�67��f(El�
+x�K�W����{PE��&K�m3����ʢ�7Y�t	1x��H/��f��1�m/x��<z8͡&O���P��! e��/w�i?^�5Ƥ���'y���g���c�Vm��lF�t�����,�ǆ 
� �[`'J��%{�}n2�h/~]��P!������}R�l4����Tw���3�_d�bL�*i�m����_Iȯj��6`9:�����.}�g�L��X��Ew���B��
��$K�,�{l�&��T� 	��&�z�,���(��qM�
��_]O�Ti�K�MDl���y�q��~��.n[�����xN�V�G��t.�۝/Ev lWQ��!k*��M.�>t:���\��fS�l�z��(Ê�#38��^�Ao����'��Ԭ��˭��B��FUY����m�p��~�����̞��f	8HP�6j)�>�x��Vh,u��rP�������1����M�^/���)�C%�k���`�^��gyo-*�Q��,�a��yԤ����~��|l�nc.� TS�d����
Hh~���������U��@=���:��]i�����'0���~���Q�;��k�U��Cl�����Q����:�1�RM6��Y����jΚ���o�l�(�k	կ���s#a�c�Kf�=�[�@���qb[?�;�5SSi$���$^a2<-;�c�c�D���S��x7j/��9 �qG�������<�8'�r2t�D���J��R�!�ʲ������E�ϒ�<ϒ����� i̗__��q�N')�ܒ�b��ˣ�kBl +��u��e X�|��*<�y�tp;�)CQ�3�����Z����R�f� �����i��Q��	���1�6E��(9��Q��H|�[3�]	a�"c�M4�'�RJ�Q���j��Is��&�*h� ��v�2q�7R�u>���������Y��ZAs���J��)/���M�z���ܿ�aJ�'���d|�K�0��~]��g�V��φz��5@�f�	���۷l.=���m�Co�	 X�-��ޱ�艳��YM�PI�C�4�[�D�$̀b!W�S���Y�Փ�����<(y���ѵ_D;��`��"�L<\	FFKZ����<L�q����_����@j|����T��T����6�H�Klf�6�x�n#۬�(��Xﺰ>�$�'N�Md	x};g��,�M�}��������f���5*Q�8#�8��Sן��d����k��ݐ���@Q�Ǳ=5g��ܐT�J�n�g+��ؤa{A³(K�_�eI�mp�c��׽����A:��o^_�#MM����W�����:�GRrpo���.����<߀4��$[3&� [Z3�kQc�<]���f���#�>"+��ב����$JZ,0)?%n�N��%� ��*��Ǵ�U��9�m����?� ��__��ZȲ��p# F�P�<��w�/�:�vq8�b_o��t�v�
����(�C���k���Uy��>�A�'R��C�o=t�ѥ@��_��_tpt��4��i���1�T�`P�hZsQiG8k�	I3�R-�&;��7�n�e����^���)|bӾY<⒳���o<����������w`�%�HFj��I�/K^$/�(�TڍuF��7�X�U�y�sT.�������(��	�c/�Q]͘ư���Mg0� ���G����o�q�@��m�������0P�� #��(cn�򴩴���Ƹ�8p���,�����v����g����,�<__2�f X*��aX��O�١	�1M�I�s8-2�̶G���������W_1���p�!��`0�\��e��t�����!d���b��fE�A�ޢA6'��bfe���P{�$�Tt6!�Q�IYL��NT��TN��'J|+�Vq�O�	 tT�g�a�yz��B��J�Ð
[`\��H��:����n��:e� �P���De���~����Nl�]�DŅ���ߕ�?�T��O*_|�"�t��@/���˗Ϲ�p���:ʜ�Xd������퀣J��&kV��uV0���nӇ�~稵6K�jIVG!4H1��0x1l���cV�K�5�jcƾ���RfM��3��y,��?g�;[��f�Os]vG�@]r�i'���f�40��M�(:��&̚��@'u*��e`�cJ�cHs���$<��{G'������I�f�m5�H�v�B
��S��=d�J4�I��1��!����u��t��zV �]4AS:dF
[i��w�ҕ�9�eZjCd����t� \�=݊���!v#M���f���<�I�G������P����=�s�_��k���oZ����`���$��Y�aר"uY���+�sw�F9���k����L���6�"��Y�.��Vܶ&I�G��F�a��;��.��:J~�Zv�E���KG�g��{�dR|VV<WU��U ��!�f�9��Gj��,�ϲs�d�Z��ͷY~���Dd'�:���������?�R�3X�����%���&�B�<l҃���� ��m}�Q���?SO�_pN%i�Y�0��J��д(�B��ov��P�v$��J]^��hV/�s�e{�->�m?�&��T���<RO5Y�jR���S�e�ZՄ�/x�I�fq�3��1
�%8k#
�#�qc���$o��I�&Q�ȒX'���P�����/n�Q�ˢiJ�"F3�oe����	@� 4 Z�!T����Ff�����$�X��H2>_��ߤm2���w
b�އ*�)�c�@Z�l��Z��N�4��ʦ>���q�`�o�����x�u�d��������� ��s�ϟ>�pP>�cY��u�Q%��J�a܋���sS�;>��'���C7C���ǖ��!��������~���uX�\��->�` �E�7�$
jʋ��lN�Q!ߡh�Tr|������1(v	���0C�`{�w���tF1�I���I�	�k�Y4��CI��������������tWEtD� ��jGK嫫�`���9t(��=����CWԤ��q�&��N���D(�Ue:> �b�J���d�P\��+vl`9?��PɊ��yeD��V��B�^��ح榳x�x�����Z\,��&`lٷy��M��\Pu�����\-��.�ۛH�!�o��聉h����]�n�˼������4����,;c1u�ZQ��Z����I�nd m3����G��P4��)'|���Of����lP���O�D9�Qٹ��9="ˆ�?�ݬ����=�D'�{Xb�k{n�/�|�a�zٗ�5��=���r<?�I 6��o��A����ޔ��U9����3��_�_�.���o�����J��=����|ï������v#�dx��l1��Ϋ�H�`z����c��0d���7�	�K�/is�A�,`�{x�A[*�!��{��P�l�z���r 6ɽ��)J��NCW</[)���������7�P�z5a!FB�,$h=)��?��
��x)���5���t����C��S�O��w�>�#	��X��|�H��ʺ?�Y���2�'7Ot�~��E��ށ����9�to����E`^��}���3$?�ٟF��M�i�]�4���:WJe �J��=���]w�����׃��������j��GK8�#q���b%M��q\P��4�T[f�^u2�2�+K�j#�,���fLS\pf\�$S��+��D���mLa�
D2ҫ�7k�P��_U���ØD��R#�s��yR2��Jz� 9Dw�n��4iќs�۷(J;)ȫyR28��o�Y�2�4�ayK-��$�>�'M�B�ew��3���)��g1#q�?_�|��!�"��V����C�QH��SŸ�/�B�8���Gтf9����e��<�����������A�i��y;�[ȕ���TKF7n!�#z����[e�O!n����uMK6��>{��\��g����r����t�����0M�qm;�S�H&nu�U^�C����wT[S�;��V��� ��ɗ�LH�8)�L*�,p}ʺ:'�:�,�r*'�}���(3>3,6J�r?u�[|>�e)A벹�ț�kd�����g~�hI���RZn����@)"�s6�aA�w���)�0���t�Eb%|^�d7ӯW�ϕ�K����SY|DOAY���"�OPvVS��%������c�я�V��3�1��RQ�W��a�fB�瘩�I\�(u�=�XJ*f�6eՒM���w:�B�eZ��̼Wa������6����v�F�aޯχ���OW�AaS�^nmX?�<:��%m.�ޔEE)���a���c���o˟��g\{cdop(e�43�b�p9&yw��^[sv�B�Y����Xr�qHz҈�,�I�{�ξ����!�ክ�U1T0�䔇�R2����!z��7��`��af����k��#��j|�/߼���r�&W@(�?X	j?��`p���T߿���^{������~&�OX�G����>0@���æ��g8"v�+�����7Mn�" ;k��T������	���!�M����Yzo�3h��O���P�p�k��ek����H��y��@�e�����eWU��[��rN�x�¶��
$��!A�N�At��<�NJ��0F��7��]���r�w�N�*VbB��VW�� :  6*S,'��H8��x/�s�;�ŧ�ʣ��ga��fD=�+���pF-��茔��"��	xв	�����B���!�\jq���I˧����~\�u��k��I��پ���*P�@
��}@+��(��V%�Z)� ���/2��t�}��b�GyFկ��:�W���s���u�~L���ambew7�|]e�^{^��{pyq��)~3�}Vu��O
@��Ï?��u3�6a���l��q�j/�?���_����/��PڋS��Iv�v'Nx�	�u� �Ǒ���߽�P޽��̖��~��[VT�r�=	(A�&����(���/��=�]tg�!�4�d�Ӑ2S"F���&\Z?~ИiF���m3���8�A)�h���3��ϣbl.��ϕH[�\M)��y0�a8&�h<�. n�xn�U�2u ��֨&O�Y�Vt�hQKB	MgϘ��V�lr��f�/ޠ)nR��2�M�:�T2�&�ˉ����W4�{,o&X���X��ns�PrZ��mJxqrJ�Up��
��f�8�Z7Պ\W�{m�SC���y@SD9~>�O�^=7g��4�����!/+�R�>CC��D�ppM~z�;�������7���9R�Z��E�Spc�ɀFi�f@R�?Kڍ�Me�M�;�s�˸^J��Y�E22z.	{g�z�0�;��hR=�5֟���46w�����˥=)P�^�0Ĵ��P��l�*����~����y� ��	�q>��G�l�n�6�sQ��`�m�F�fӁ����}y��ܬ�2�?��M��c�m���w��r4�pս�B�K�*��{-]	�H�����s'�)CE	�{)��,T:���GL�&��}E������l�潥�x�,�=6�`���]�v�Z��v$�oG��>����s:�Gk@FB��>��V�g����ѯk�3U�?4'�!ʇ�2��F��rҁ���3��s��`�6�|8�F`g�ZAR߆ �Vvִ�ݳ�83�]C�1⃚v�sa�E��T�`D��4n��4�2?s%����Y*��e7��M*|f���Wh�K? �7���z��xԟʻ��qB�Sn���fC��^e9�q�h:blL4CAhR�ӚA���*���-Az��sO*�l�X����|ٿ'���Q�̂���0�3�i"��pswσ܊dW�Q���$j�'\��g��j*����@O���v���c��_�����y����^�� p��~�l���ՔjY�Y��v���Bb<4��1g��z�k-��x.҂m�h\�f���JVV��[����Y���Ɵ���j{6+ι;D�:�Bd���i�X�g��#��.13���aSO�x%���n��3�4N��m�B�CU��p���=eY�ʒ~�������$6�%�X���`���Y)�l�o;�nrK��i����Ũh6T�nˋ�K��P������}��ά��E�/R�@Vfp���G�geYH/����\B�c���ۋ���3��'>�tT�3J��)���~�6 ��J�_hW:�e�v<��Jz��(?���~i��8:�e�ؐ��t�H�~-c�3�ނ	��#�Hdk����UFw�̚�oY��f\X�ō#/�6��f�9�*B(����Ca��S �	�����)T������UzC���|�����GZ�N�Zsz뱂gX�Z:�;>�s�:���W����G^�o��.D�!Q�r,��j��{������q�xآ�@Ѹ<��Lٷ��C'}a$	M �M���P��:��ڥj��8Y�eChї1�t��3��m���|������ ]��ˈ�e���5_��r҇e��y�97�D�{�ʯS7+�R�8$n����6�'&�gG���K�»e	�)���^Ä���Q� �LE��1�h��Q6;�>�AT���0���Tp9�MxQ�D3�+�[ݶ/���N�2RRg�K,8�b����K����#�C��?��rd�ܯ�l�G�����'�4wv}A�B)�{��N1Jo�N��KS�5��KJ�d5��՟Ε����J���1�����'��a��.h=��@
�&J/i�rsc�b���h� Zj�ou�#���Lg�y���4�7wA�ꎙ����}��Wr� �y���~��O|߸N���(]�h!��y�|��oH��-�8�gP�w��b(����jO$�㾜8�o������	6x�q�q(aR��_�z���ua�04U�S��	"��,�.-�yr ՐSf�O� jrWҝ!����b���]���z���P/;�\>�8�6M5��l��q��<�џ���X�,~�c������Fi<�[�	(3��ɀz>�o?_���N"��\~6�Ɉx�	C�*z#��Z!���/��3Wـ��Aؽ� �B�9��6e;n�C�I�u�x�l�M���\��=�)hҕ�w������X�L,w�m����^S���[�ku8�����.�-[#�LϦ� �\�,�`o��V�-x����`��X���H/�˞�։8��t[n��<Շ�~�ݔk��K�O#)>$���__����%r� ���gϢ�\��ׯ�O}��%;��}t�1G��� ��<���5`��gӴS��T5�Ƶ��\\�usuK�`�9��c%2��u��ր�ۋ���ʂ���6F^7�������"p��U�2=�8����u7��I��zŠ#��j���K�L0{�B+8iy���d�ڝ����0pB�*T�b�$F�}}�taL���ĥS�a��Yk�l��j�ۍ;���}7�6K[�W���� �M����\%�;��җ�ҳ�fP9}��!U�b���	���C���%��3�����vI�r4$��گʌv{!�&��9�Ϸ�8G���w���^�} އG`(��}�����R��#}���9t<n�"���mG��"P��ȱ�<!�DOz��	q�f��<<T�P��*i��N|O�D B����q�~��SD�F�#�5~n䆞����Ԥ��nI}��	�e�4K��V�]�뿣�͉�CYM��@:޲\����=�;�#�]�<���؀�&�s�ݩ|Z_���X�{�#�+Ϟ<-�4+��!#�QI_���01�����oI��D��F�i�M�Ӓ�sm�<p���Ȱc$pf� �#����V�B�<At��3��뿠��
�T37G�e�a�Wql�����J���;8�	��X�t"8X������O�Z�@��Νx������(�}���6{v!�m��^xNf�࣮k�4&�s�G�֞<eՀ�;�`�Y8�LD@�n��נ���S�,0_g�JTO���{
]� �Q����;��t#G�C��{��%;�K�l���+�ge�m���=�v�Ӎ���H���p,�T��p� ��N����~� z�9ԬL�7�#q�le�j	�Y�)n��S�eT��RO$�"\H��9:��C���n)�#��F�3H��x:��x�Y<cÃtN���X�?��%f��{�7��Ԣ"r���fp,�:tB�o�� N|p�DVq8�r�i+�[����T1c�$��;Jm�y�.k37�e���=�C�����rW(��?���h>h:�Tfb }���~Q���"����>��Ȳ�ZK������bW�"����!��DB�}?���|�-E��e� '*�J�i^��� ��ei���x���Dk�
�Ŭ�k �/�t8��C���Kwpc��Ox����.�"��$䝃0K�&}`�}[��)f�'�g��0x���D���d)<�9>��l
�W#!��m��^3dH�a1f~�=���h,:���?d@���+R�zjZD3��k��#��m@^�>�!��p}���>/FbI$��Vs4��,�9���w�>���t��e�Ϊ%͎V�!?���:Mj�Z�hɲ��?>�Vܨ��*:�#g��'��{#���8{��(�v+��#�x镲3ɧ���r{Y��ip(˯�}��өb���[�iU&/�w�$���\�%�P��q1�U��c	������=?3��NQ�ز���|.�1�w��@��J~��\\��33�ȼ7Y��;>3��t#��")��V�_��0]�Y�a��@�,<��0Y������eѧu1�%?J{7�n0B
�e���(�w�-��p� � ��Z7�T�}��3 ��Wgk���8ޭ���7ߕGk;��ײp=8���z�M��Ĭ�Ns���������m(d��'i�6'���s��g�5)�����3��ʏ󫈣+]�2t���p c�ܮ��6�`���2�����e�����q���N�u�~�D��Y��=���I������~=01��E���3 �Pv�(�Az&}ӏo��ϧ����X=i��-��W̊��ɫ5��t�~��qu/0�J�_N�����0{�+�8W��vX��fu�ج��2��5��|��N
�e�}�h�Vg�_�lʥt�Wq#��+E)���.���X���+��ԑV��x�&��'H��$�)��8�-��<k����_Z�')<��7Ew22�>1K,� ���OE0D����3�!�V���?��,W��9�d�\�N�x��K{����\ҶX�+���r>+�-���P��W�*O�~���R�ϺRx8p�j�M9���Y&"P�Hh 0K]����r�0?���+L6�P
b� ��)��8�0��a�1���<D&���r�JE)M���FJ�x�!�"�"���Db�߱	�Te�p��ʺ>J]46�m��%_�M/�/��V�. =�����,?%����:��|��N�l5e�E��,
Cpx�~z[���ӣ��E�N~L*�
�ڇ�2���X�L?S�l�W0ޢ�����J�X�ptC�l���D�k�5��!��
	��&�jk�j5�_��f*Ta��v��kU��5�$�K�� ���ա����#��AZƅ4�Ds:�嶛b!rO��> ��P�@�����xJ�_�fx�F��F �Nx������t��@(?�0�t&��)��L�"l���L#x����>2��w9^	�x��/��2ũ[Q�X����`6��%)b]���� �@�TF�Ξif��:uM�I��u	��K�ސNl��ح4�(�A��Ե� YbV=Z;(s��ofI�s}�����͗l,2���!�l<Ċ$%=�h��?}�Ƃ��q�76�	�pw]4A5��Tf��?�85/z�F.~z�jW?K�v/8@�O��!r�C��o8��Ӷ��4S&n�.)W2xW�"�0�/�X��/(y�5��;>�ӷ��cX�@�p*� ޯ��ǈ����>��]�%s.�c^� �J���J����� ��M�9���.�UL"5�9Y,��[���sò)L���M:���S
�<r�Ջ@*��3� �����%���R�����X�������%˩v���#��4m,��.R��_�ݥ�0́D)%tx�<_X���(ZL���HV6��`��ӧO�b�OI�
1<W��V�@Z}*���|;N��j� i﫡�b%�Ab�k�i��{Q����5T do����g3�jܟs�?7D�<s�U�WD�/X�"'uS�75]߰����
��J��/�L�`�C�h�|�O�E]�z`��֠:-�3 Y��`��ki���e� 2u]隣���ƳJF����^`�Iߑ*�F"�nsM��.�%��-}����j�,�G5�+�IW�L
ƈ���R��~��5�SWt��W��Ϟ���7���X����L�v�]VbY��ەTTG�̤f�C4g���^Jp!������|J�̼�ρό�@e����Xf���W��}0���ۘ�:It�M)�J���ҽjY>�-xY��7�����T�п��\~��bs*��Ɍ�t?3�ӇQV��ܥ�T�G��w�������rt뱩ݍ[�8�"�*�i����io��\�%R4����Yw�W�(b�l<_@hb�/2�F��ZZ��Ȣ�č�f]ko���c����F6��[��XJ�����dKwy���s}S��=��\6�����.�.,���~/'H8!�t⼣���s͒ݑ]e0�肩�k.�a d�o|Ko!d�����Zֿ
*������`G���OL+>e����~l����{7j����
�,�ݷ�G����)�9��%�%6��ᥤ.����2�^�1L� A9l9|��Ff'�"�����L���v��)��(eia�SU���)R}���J���K��VL��!�J����8)��H��j��f�7Q�	��iwAO���m��ƭ�:}��6���{�s1���7x\l<ov��!�g�ߛl�;g`��1���K�Y/N�ǛG�|��jR�u�b�1Es]��M_���������m��dƅχ��5*NXX^��LX4�fA�6Ȕ�*dY҆���ڮ�U��e�N�KK��Ǔd�,ivY|$*�(R��N?嵰�@�.F���@�[GP�� ��rs�D��Y���ƞ�����g���t'x�� {���[Q�~�Gf0����}��0*{�Vo�n��8h�%�U��Uɼ���d��\�n�o�s���a=�&�S��2��ϩ���lb8�&ɩ�]�v��x�o`�!Z)L��- T���3�%�|�09�/k�R~��P,H�頳�_�f:`�T�m�2�x����rv�����Ϻ��E4���,80�H(>~����NR��y�sB�7}$N��#�ָ���@�X=�R4����v��ei�����E�0�F���_�	o�܁#1�i̩'җv
\%��"�Rr7�*����[7֤�NI��8�Yj�<J���/a2��bx7F�$�[�i�vV������ä˛�]J����/y�T�:�<7@7���k@'�1"Ld����pee��l߁�N�L� MkR]4g�oAi3O~Y	+X��%:��LF��pB�U���L����c��)~��pPM� `��E�㚁�;�;�Q����pH7�MDt/h^�s⥋^��%��z�a���f.��"���|`�]m0i,4���`�HmG������>Xsh�aW��*�;l������}��S@��tnR ��+�J�X�H%�#)�A)~}+�kh�b����������'1�]&=�ׁ�"�i��My���#�}V�����-a*Q��Y�89�b8��A6Ⱦ�	��'�H���KC��Q�
X��h*����s��/E�ei#q��=�r��m�ƛ�%�˺:ƣ
�7W�\w��鐚�xFs�\o�\0NR��Y���i�ޝ�:fS-��l��X��^��V�y�0s<6"тZ�ϖ��p��A��8%��
V�W�,��rf����5������U��R�@��SH,��.���sN�.%H�$���/�@�� �/h5�f��XXeL[4)f5�B�w#H%���9�N�#~�?�� ���v��0C	�����FV�����?���Ebm|�y��xFjtL��vM	����½�Gy�r��_-,0��Ti��K���?�JŽ�3ŊG��I�.��<��mGضD5�go$��~���19�Gf��{a��������zj�j���>����ә�k�j�n���@�ဓ�6[�����Wt�#��sy�KWߚA�{k��zԡ�
��:���T�pQ�"��uwY�7Yͻ�w���q��?�ڷ�����C���ҽi2�������� 9/�������^�uQy�R<	��%&b斋�+��){��м/2�e��½�W�]=����'~L%�9ic���=��),R�I�Z6㳗R�	}]� �@���b��q��7:րK��3�C|����j�@G��7���Z ���8����:ʢ#ӈ�0D,�~����FY��E��x��������C���x�,��G�n�������o&y��`s+#`���9�q�T�ɚ����_|Ů�N|0[�����y�����j�2���#�8T랛u����ǝ���Yf�%.`̡����c^��9�_?HD���N�pә�!���U���L� (&A����6|���<�f^o[��/1�Y1�3�l��.����;0��fh?4��*���}#ڵ��B]���\,����ӟ���i�I����}�iz�����G/)S�y���:�`N"�k,�"1q`��>��^����w{t�'��)ˇ�t���υL�,<\o��Y�0FC�n�����Ɇ�'���6��|xS��¬c��Xi��ʂ��v�� �ˇݧ2cl�ѩ�FP�Z*�����A����Ä�Ⱦ����+�1���,�Q���gg��ٽ��������i��x:V�� {lP��FA���d(�ݶ�Y�ǉ�41��������ݭ�ҹ9�fw�V�uo��뺚�}%ㇿ�Pǃ6�(��o�a<��բf��T�|w�'��ѐ���(�%�|ntؑ�o�����t4�qa�:�{�q�`�	er�7�CY9�qAl6&����i�{�P*�kzT%F�|%vF6l�'Ա�)�}H��m(��:���ji�rM]�\�P��|w��n�dW�m��0����݌t�L�(���&pȋ���)fW�{H��!����(E1��(�Gԃ��˅�����ٺ^/T��Am�~F�zv�Ǹ�8y��g��N�C(�/��:e����e �����j:�s� w�(��H�E��f|A��z,��٢������׻�x�3���]W��J��`9��:G4ů"�I�������ẩG��_K��u��Z	�Ӂ��m���ch��psh�˃�">-�cn�v�xx��nF�����h=]i�K{}��k�]Rg|�JH\k&���ذndCI5#]�ac��3��z���#)��A���*^;�붼-�^.1���D(��R0�{�B�\W�!U�<���2�SN٘��:�P	t@��>���x�����"�NM �X�H�(�:35��"�Ɋ������H/������g}�K�@0&�u�oxv�7IY�9Z/�^Y�U}����E��73��-)�r�^��'�RqQ����o_�����).�qӒ�>�"�R�wu�jiJ1e��-)XL�
����,�l�&Y6d0�$e6M�������L��q��z����b,M&����Y�#�+�J`\s�ŚL�A�ڮ(-&ޑ>��b�$"{��!�s"�'�a��sp1nz��Ō��S[�"]������]]tf���Q!�G��oK��?c���R�`'��qH8@�����VD�w]�Z��
%��p���0���	f:��H��h(�)��<th�&fH˕�63�C>��@�~�$T	��+�S@��xh�U�Y�RG�ƙ8�<�����I�nQ�����3���x��-��h׃��)o�gM~�J��T�JR��[��'�m�!?p[�%F)L)�e��(0��}�]�	��D&�Ũ|��P�S'm?�^�W'lƜ�>�V&l|]-����˧�F�� Z��(�2%�/��أAv[/�)����4v)R�?�2�s{T{��M�Z��F��W��q�ċ{P����e��!�����m�[m�ϽdV�4�*��3�"�7��e*4W�ጃ�or�D|�f���x�@�MpD��q�0|s���pY�}��^_�	&齎����� �z��������J�pă�Y�r~�+�w*��|�Ek�辎]�߼���Myj���FW��)i(��4]b�5����$�������Iy��%����p��նߡ��ʲ�*U��O(����P����x����͢M&B�P��CǮ�SRZ����A������t�M�K��G��.*'hc�@�Sj�,�$c*\s�"���f�S����X��Z�+�)]s���%S�o&�/�.�G܂�4&���L��V�q��FsF�`�ٷ���R"�s�b\?7�6��i͋s���@�f�,�&x·;�x//��d �葴��xt|ޥ�ƌ�� ��x�8I+�5�-�ğiC!��<�ys.��dш�4�F6�]-9�βvA��.3>��R3�6�a$�s�g�u�������,?��M���D�~�i6b�U���0.�������x;Ѿd܅HI,�6���"��<�$p��Hn6����N��7E��z�u�j�.�1��0�w�dY�8n2@���z%@h\K�Շ���
���I匠5P�e��g/J�"Ll���a���7,�}a��C�r��n�B� ����Z�Y���x�]������^������aF�5ծ/<�ߣC��ɼ&�f쏎�jO�I�����:Y�r�L�"��soO�) �-
��
�E�>��cC��C�����ư��,u�8�Z�'<<��Y{P{VՑξ�r��E�7k՛ ���vsw��u �`H�yM7���Bo�>W>$<O.��Hh&�z8���{�~}��F �vD2�(M(�񳽰�R4�����w�����l�l��/�L����\E-�ک��㸡��E&�s)�SK��C!OЬ�����?�KQs�	��`��K����v�y�K����d����g�k9�o�Ȣ����A����l�\�Ϛ��s�9	8׊�9З��Ǵ�����l��i�U��X��'C���,�zǤ:���}�>�I|��x}Oi����O�r�?k�!
���)X��d��d�_������?��P�k�4�"�/ƿ�e����f����InvL�xw1�)��]t�z���̇d�s����S�=�0��=�� ��P�W���t�i�V���@0 o��cq�wblT�֙b���s��o�Z��� ��=�������E?�( M7�m?R�U{���f���bi�������F��$��0�{��e)"�sl����^�/�q�� kl*��μ��6Z�1�Y+6�I�O^�,����7�'��%�gF�$��T��'�ܪ�i�
e(�s-e�e�?߈�WЫ�i�#����Rjf
�^-T�ϩS�E��6�k3c7?�)�C�)�" k����[B,{n&s�	8��-�)X�2��s -��-.�ES�Ą�"�js���գ1���G��C����QQ/4x�K�B7(�[�s�:��d��`˩�7�g�l��=��4q���kɿ+�I#�����
�G�|6����/� ����e��<�e��[/�A`OQ�ܮ��xw�cҦ=�Qچ�׎�����f�T}����l�1�K���_���tNH��;��eG|;]��W�t+ ����	��l�Gp	#@�z���R�Ė�\�-ϳ������8Z��g���7�b�?�����_S��/�s��?�'3�5��=��T�<r��?�*����� ��Ȉ ���+OETn�I�͇�~�ČX�(�pT�M�2�9G'���r3�+�Ģ=�LTY�V��6�K@H}4@bp���W���﻽ֱF��['*�A�R�֯�1����Xa�Ҏ$�O��D�l\M���(�⳺�aU�5;ż�1�,?�k��ס��>����Fj�"��Pt���ף�����ۗ�O�gO����H����81r�Ղ,���I�g�6��Hy�Ͽd�P-Ӄ"	U�asHƌ;��oERC#J�턹ڊ[�B$�(�Ej��c?t�6��3��Ҁ->(�z��TJ�ҙ+h��|�b![6���R�ڃ`o�A�%F0��r =q�m��%�f�w^ڋ������;��}�(����X�q�#��9>)C|��� �a����2��t7ۮ��{O6C( Ŵҍ�E���|���,��d��o^��Pb!�~���E��̌6���4�����i�C'�R�$_.2㺾�fe��䭙3�ߎ�[����ķ�׃�2�a�Pc��l�y�~[|u��mr�l� o#�*>�fJ���ǡ&���+��H��7sӐy�SU?���� ��_�Z��\ͥ]J��]r��lW�'���3CW��a���Θg���~��L~��fR���G�Ž��2v������e-�R| �{���x�r=��,��x��}LHTRk�hw��׌t�r�v�b1����A�U�7@��A�C��]��R����e��ץ���X��e@m����=������fiTq������9���6j�8����8L�"#���6:`U�3:���Qdx�?*����JL�|�K%BPY3B3��oN����	����u"f����5]��`pާ����[�����-�X<��kg��n�w%@���Mr�
�P����o��M
ŘF�A�'q�.�b�O�ţW��ͬ�̹U2�ŧ�?�RN�(�f"���	H u�J�0���2נ�X��&MVw� yE�Kh��x���d6���W�Rh�y�[@k��$H&�AP�RY�e�"S���e�.�� sB��y��n�Kh��f���6L�K.��RrM����hvjn-uM��.�����P��Jw�j�Ce���i�WS��Qq����}v��ɭQw%TK��RU������{⊪r�}M6����<���a�dm�?X���6����}�G�����Mr�RSr��_����Գ�0k�%�����W�����1��p� �7E��MC�Y"N=�*�$�"�P�A��S���]�c��TJb^��K��$p�w ��w�6Մ�"��5�V���rgxި"��2GwH�n@!���g��W�)d�=E��ГlDy��C�N4�J��!Y$��Q�iߧf=uj�z�e�ػ(`G	W�����PޜQs�k��z�� 
˗Ǵ#~Q^�q_{����3�QӅ���Kh��&�藥�q6�$aL���=���=z�-�&+Ö.jTk��zY�(�LjH��KXc)9�P�e��>�+u��v�'�,����%��0	�5s静�U��o��_q�庾�s���|��XeR��(?^�Pi��]I�a�1IB�;)������xy[vc]�1K�y~x�jI_~$�� �f��/�{<��/�9�Wf1'�K�j�y�1��肋d[��t�B�{/1�#����YZ	:X�3����44��#��	C��w���H��_�L5�j�}�Q�$uC �&'�.=g<Z�i��PY����m�M���iOb�3GެMx�[��/�iRFj��z"��� h�p�r��)�$���G��S`���*�&��KB��jHuu���~$o2��R5�.�B��k��ur��FLh[�W�1��/<�|�g����^4�����T��QK�_A�����\@������?wW�Ǽ�;I�����n��5�O��� +^�%��&�ٝs=�4�P�GC�o�~��t�:����.�ڰe�_�Di"�	��㭇T�H�Z���� ����֦b���L����چ��[qoG��א�a�������H|�,i�y�%05�����P� Z�}�������������=��5�zE�R����.j��W�	r���Sv+�,,ؾ�K�0�)J�6�Y1�g��s�U�N\\L</�7 7'�p�/�do�z"�J�{�F�bX�M��m!��B�,��+�*2��!R۴y�ʑ��!�	(��\2��Z��7�7y��[��t����.��u��zu���e����Y�5���t���}P�z����E!���q�^KIg�x��ۆ����R��qΛ�͗�&_藯������">�
4>��`լ6�֑Uʫ�k?ls,�B ��a5!�����B`=��j ��E�OҼl���bZlϧ\�Y�u:ͱG&Z�Q�_�fVe@���/������0	(�pX�\�7M�b$��>WȍY���x���������7��U'w�P������ԜS6�����I�G��� :�������ǯj6��d�X��s���;�"�ؿ�4��r��E��1�� 	*�;�T:?��xHC�z�#8��˂&�/����٠���|�#ٞ�91�^5Q�EI�Ʃ��O���X0�v��.*���\ov���^�$>?0+����q�z�\���kb���F�K	6��ȠBQ��Y���i�1����"��Y!���ZT��_ڲ��;��ݠ�i��X�ᘪ��ә�����{U�s�싗�_@�	�>O������5����Q�.�0���{�Jpo!2�3����]bddඓA��$hhn���
�M�*5�-� ��{͈[����.�<���{���vQ��jX�K�6!��\{�q����K���z �y�1Qd���XkN<ܔ��o�-.��c��o5�o�v����-���d�qȇ��?�^jV�}0n�pof�d�SV$�v�5�֘�K���Jk�?�2����r/�����C
{0���EeH��_zG�Mz�lR�"�Cp�B�'���u3w53�����������@�]�ӟ�ěg�FS�p��ͼ���ہ�^���P>�|�){f��7%Et��}����чz�V��6�zA���)�3Kah=?��EB!
B6��QXw�f &M,��{ ��1�c��ٓNMT�h�k��YN�%�Q�P0�\���.��MQ����I�J����UvG�]bh��L�R����]��_k �������D��`�j�m�-󒽯R>oq�
l���������	�o��V��9���=HHĺ
�F��Y:���?��8P	Xʰb~�Y�wK�����9v��F����߮���+��l����'z����O�\~�O�Ĭԙj\���� ��ӄ۝���%��	���I����D �3�듧����ʱ�@���EV�2>i�OQ}���򾹖�&k�R?H�k�+՟��T$a��p!�l�l�s��7
KK=/�a�x	��c�<�Ouk�UOl��YNn'K�'�Px- ���@����[�w����������Hy�:T�)ӵ^|���A��A��׍_s~fbŚ��k�S��N٭G[Ķ�w̎�9��w�����@u^<�k���a#%�ི�<��`2�6早A��.U�1�o��7>g��C�W�'�(3�P��YN�`S�����ט�u]�}���rkQ:�[�������w�����|�W�Z)^�y;}x�1f�u?����:��}��+>�RO����x����r������n���E�"�7)��l�\�E�#P�yI����Qohc�}������HKv��%˾T2;$�������S�������������Ì����;�/���۲Y��ڳ�1$݄�O� ���R����O�~���8��εT��+�p��~���w�0uR���������Qyk�.��F�M[&�=w��bJD��8^�Cה<��.�����W� ��b��cu�n߀�>�k���a���f�s!h@n �8

/%O?�@��E�h��g�4{
N�{�pm��(62��FR��P�x��C�'�$�.U�,[4�{k&No�O�dĥI����M����9QvִJ�c��`�ts�Z��`�K�.���_f��X,yYJ��K��u�bė��E���׿�*��.6���L	8� �CO����oT�\b��v��5�89Ŵ@c�b�	2d��F��)�T�G�h遒�N��>��PL�La{b��V�.:�`JXw�SESfO.㗸�pNW#�	�o��Ω]�ϥ��,V!лHܓ���̏W`=����U�н� ��P�0>������I�Cd]��������+M��������'i�-�\WX�#���O��j/!�3K!���n���ϺJ���6���F��|Ef'%��$7Cq?�{��F�6� A���iez�8(}NJ�'��gvIw�G�]�L�&%�.2�?mo�I���/� ���z!�x��_5<w�4�]��b�e\TD�,�ȪjNTG	"�mQSE�O�T�7�`;��ـR��7j������j���A[�|��&�y9ǆ�[h#8��
�u�r"W�+�ԃĽ2�2U���>ȳ����}=�jü0)h���61�&,�8e����O0$'��8!*3�'3�[�Uv��
�]s���b�EriyHu#=��^'!�ԝy��8��Gg����UD���m����Q�D2��*��Z��;�zx�⨮��=�h�(��Ś���1���$V*}��û{����}���R~ݼ(����yph����\�>����zKM�YE��<P�^�Z�6�I-7G�SH��7)
�Ա���zA�0g�?���q@@k7�_�(OR�?<��#�2|N$���6��o�K�=-���>��3)e�(�����"��a�`�!�������z��E���jD�(v]׬�z���q-啷z͈�ħ���3D�/�5��A�yZ\c���E;�M�8��K�8mH��`b(��z�K��ZkVY�OC���!�mum�+�M�/�e��dԞ,aH�ȷ�O�֚e�ˠ_=��������B�|��ݷLp����'E�(���eG ,"CSt��?�Ʌ4�1��T�&}�6879C��.���.��n���g���(Ȑ�ȁ�X���&i,���	Z���E2��	{�Hx�ۿ�[<߽}�̑ɳ�S�ȱ�7X�v��oƴ��n����q��B[�P9���%BWxP�x@2�!*x�ž 0�0�����]# %����Uf����\�������{������\�����=p�?�h �ID�����ޮ�5���,�	Ӌ�/�	�N8�xў���lQs��	#ڍL�Xs�0K��%����#Hk	�e6��@�g��++l�HF�"7,�v9�R!���c�s|�@�k&O�Ѫ���c���W뫏<9�7�����=���6��8�&���
RE*�i�zu��.�#VG���kz��ì]B	��?`V.�[�kҌ`TVe��w���|=�������F��)���*��c"�"��혛�L/�7JgjR����W��(@�0<3�󪊐�j��	'<0&ͯ�3T�橘i%�nn�����O[��G�'}$Ԧ�(Qon�QA,����>=��������?G_{�e�p��x�7n���R��3e���m��;o����n�-Op�(zb?*�-��QP���ܟB�@Q3�z�Qڹ����iQbL|��4�!I����m����B���<�dތ��cDp0:��i@��yWx���"��^d�̍`��ߚ�[k�<�1=�N��sx�OOSޝ3��ws�1��A�Ar��*jO$9��'�fTW��	�*����K\9�b�-��}���f���mQW��sܸ1����i��ά��NL�*|�
xL�xe���(�߮���iG^����E�<������m����Z�xɅ������"af�K�i?̙�k��"˫�G�5�{+�!�#I�=KD�e��'z9��R�A�~���#*���=�^9���E/p�pR�A��v���"t�BP~�6��Y>��"w�ǁ�]$�@������OT�T�2dYfx�-�x|Ц9���C�J�7�Զ�~�r
�&�}ǚu�+G�7x?:� 9�#
�1�u!l�^��BB"n�R~���x�����TQ54���RP�� O�O�K`��p]���h?D��rS��&�8�^ρ���>�1\/n�MVɵ�Re�'�׹��p}d���k�\�z�����+L���%��ѮG���E	w����!j�Ѭ{�]i#��<.���n�P�${:d�����9(�"�W���>̎h�?j,��R��A�ˊ2�ڨ�JL��!��C5�1�>�z��o!*j�1�E���t�rÆX,�����o��S����=���c�c�ӠT������y���d8���yֆ���Au�%9��m�f��e�E�U��D�p���˯gb��?�����-�g55õ�UPۢ<���4����}
�)�N�]�C~n�Q`\?eS�gqlkE1�h*��S��')WK�k()&�A��;��'�C�����N�K�C�7�Q�U�ȵ	�5CR��L�7����ً}�1��:�ⓖ��xf���6�Y/��x�?{X�\4wKz�ħ�0��������$�d����/��ϒ�[��>U�iP��)�����!��B���z.��k���,�0	�a���׷�ފ��69�xZE?`6Q�Q��q��t�!����:3u1֏�\
Έ��H�bͣ"h�h	I�4k9��5�ǔΐ���I/{�x�gS]�y���I�J�i����kR��;X��h!;tl��Oo��FI�R11��6 NR�k�7��>�}�M���ℵz�>4?O9�'-��Zz�le�0N�M�m&g����mdʿ��`�B9�׊m-�gQk_�Ǜ��.iSx�өSGMʶ��-�#�Kf9�NN`�����R�[l2�T���>tJ�c$h����aO�X��-�=6�?B��g��R��s0�d2 �d}�� �7�)���a}/o��UΐF��ǨLB5������0���X���f2&�XŴ��;2�
Akr��H��Xn�JHd�����T~�	��{7����K��
FQH��x���ah%�����������_��M��s�߮�*��"]���z�&W����\�;�Cy �x��R����ٌ��oj��	�[F(ƔMK3��a��ʮ��#�>);%���£�OQK��k�vI��(\�C���EB�d)×��/��և폺�ѫY�{S�-#J�emz5uiYjwŖ���n��b:Q�%�G)�܋�'aP��\��H[9TUt��Xk�wc%�/�Q��{�!� �:���2�� XA�������x�E��}����e��͢jc�|gZK���׽���u�l��~���%�C͎z\�T��e;vm����:��Ld�! �=O�?�qaCpw��?n)�Z�e�����k���|���w�m�w�ަ�v$8�
-��<5:����.�bPo�11HB*��%'�/.뜧{q�Nso?��?�R��(c���^���5����
,�������q9*��������"�,Dh�2��L�\���� �bb@ۼ��F��1�pG񮭐�ŵ."�E���"ٷ�s��-�6���v����jq�)Y;�<���Y*�����(�Bh
{�*�e��l+y��\r�ԫ�k�I��E�[��� �?)+�eD}aj����T�N!]�B��M/E=\ƅ��#���.A�M ��ĺ�Z|�1m�R
���P�{��O"�d�;%"��a���q���:�NX\%<����JQ�#z�bِ^�ɴښ9���Qn,3�~?�=���6����W�'�ɈgQFކ�uah$��{������%�~�)��_?�Z>��!<�i������˧���:�sM�Z��*y�=G��hG�����W�ӄr����\e��$"��혌�LT�	@�M�����4j��wX7q���7t���Ȥ�.�S!1c��k~�h�����<( >!�yē��G�)qx't��l�Qಚ��zd5>��c���mXp����a�<*��Ȭz�l��몽��=���6�N����~`�0x�F��	�d��q�Nb	$���W-*3���Ȑj�&������ژ:�o1ӱ}۴���AB2i��B0<.)3="��qdI��=�m.���$E�/�Ԗ&�[�����ROB�ά�T��e�&�
(�
��8��v���I� ���̶�-])�{��!������W�S��]����Rn��E�7L���U��'6'4Bipugz�V��\t�(��,b�d"��IN"�$���&5� ]����~���X|��������Lr���,2�d����+5S��fm�;�D)�(E���G�g�Ͷ�{ml��3J����M��Ya�uY�y����"���?o����#m�*���Ak3G%��t8t�}�jg�����Ϗ�Tߤw�;2;N�#��QG/Z�lS���17��0�!D������D�E1n���E�#���`�y 
�S	F}Ɲ��&s�d>/<v�H�[�zR6�aC�
2�LC
.��(����k���@X�7�a|����j�����,-�l"�I'�����t����T����"~6u��D��DAG��N�}�E_M˼#�@b�O��kL�k�[j��|Ԓ�)X���S�ӧ�"�xd�`�э�Ԙ��[)�W���ј)NL,��ԉ�
k������	^V�
��VI�^Vh��>�J�P5�������%==�'$|f�<��&�a��&����Cy���HX�d��E�r��&�k����!��I�����fyP�A��W,^<²ޗG�a2�f�6Dv��v{�җJU�|��.Z������]����'|ӜԮ�֡�v&��aJ�C���4J��]���w�b~�Ys�7ôa�>s�+B�r�C�!!#B	��K���Ab�8�^��| 邎���^�����a�I`��Ebz��VFs�Q���q�

�~���e끺'� ���{>�/�&Ы!���[i�Z^�9�������7)�+����9L��d��og�M=��i������Sm�O�������cf
1!� �{�p��ކ���}̺�,��$o�0o]3Q�G��[z8Q�&�ױW\Ų��@��Ȇ>�G����Z�c�^��Q�Br��&1�5�4�
V4&Ɯ�y��G,�Q^&�i5�2���_��~�	�Z=��ez��oi��ab����[�X�6�	���WxE(I�m���Q�����*{, h�F�	����`��gb뚘�a�[���Qdь8Xg����)ֆ#+^[�&�Z��b^��h��3��"�JzIg�圴�p��91֪�d!?<��nY�`i�vngUka���ݻĝ	��
����ib���v�k#S�Q"v`>Je?q��jW-�}�|4��`�����n9�X���o��/<�W�,,�W��ݞ�_ϒ���â���D� ������8�Ǘ�U�]χms'���������:�+<&���u�L�EYHf��#%�o��|��e�u5���*81�R��;c�Zf�:�9�JtL�F��^ҧ�G��(��<�j���ť�"��X�_r��{���� `,wҋ����ʹ��JV��!�j�;x��5�L�!�������:���5�C-�ͬ�e��n��<Ϭp��da 3�!�?�yb����o��p�5���)����=m�(�-)���:����wU�5x��II�d���V'eҫ�^?���b,:�E�2�W[~�~ %ѫ=���^���z��yU~zMH�1�O�(<�������/ϟ�>���z�G�Le�Em�.<WT0R*s�<öם�c>⒙y*�Y�tI��[�
�^����~ȉÊ��뻵g����y����ᑚG����;�4~"�Ag�c�l�����y&��v�E���0���Pi�֎��w�YH��7I���x���X�P�1HnB~W�!`�^�R��ݫ���i��K3�u��׈]"����ۤ�Pݦġ2b�a5�����BW��N<p�?3��x��)��)2�Ƴ�Ӧ��k��ш��k�!Y����4έ�=��KG����@�˗�Klfױc��H�2�e8�̂��
в�G�1P� ��p�X"�ޏ!��!y|�)Y#��^ۺأ�G4gb
���x�/�x�F��ſ�3��>�䫲�N6Y�&���ʎ�|E���ݺ0Չ�h���x�Q��ڮ/����9A^�x�j[���}FyW)-9w�������,J��m07ܱ�{�^�.� �p�w�6I��i F|fW�*�>�Z\��O�B�-=�i��@�cmC���o%ӿ2{�-c��C���_v/��{�*�)����H��O�R��������]:M*�޼mS����&�N~���>>�W��)y��5�����{���+����x���k�12(o���Km����i�cc�ZLY��(Q�Z�$t'y<>�=Fؿ��q�삃$�+2�rk3W�dc�	�~��<���]�γSɡK����G2 ���j[��8����'b��Z��aO��&e�̆L<x�9	�̼aDoS*&�*��z|���;���s�n��Ѕ��T!������5�BO������W֛M�0��U��r\�`�Dx8%�va"�Љ�mZ5*hD�rƶߒ�wz�<]�)����c��<�'�K�+F��G� >Q`��R��Wӯ愼�w��n�c9eY+�(k�On��\#Q����č�R崔�kjN?��̥1t��j�Ք�������UV��ǩN�=�j�ǈ���}-Z��IQ��jT��D(2�w�G�{�����>0jبT�~L`�2iQ�x�ݝҝN�I�R����83_�+��s�$�/���d�"�Q/�6Lh�k���&x;Ӈ0ː�ENچz�������]y�=��a��nw.��R�dR��:W�}n�k
Y����~�B��ɼ^��Qs��
�8�)�,�գ�]z�yq8�E�u75�x����I��14lM��M��݇d���%Ń��#%x�R�][���)����׻z���@C������ol�Ñ"`t>|�D����A�l�Y�rK��9��0u�@0Tz����֬��k�S��e`��\\��^��|,mG;�CĤ#�s�,�n�E����d��Q�
�cL�1����YQ̤��l:R�w����eqB��3Y*m�;�K����珄����k�h2�%tׇ����n��m������G����G_y���Y��G��)�f_�6TN]/�?K��[����bj��nZd���|�}�T��΋j�q=Q��t8�b�!��}'�;C�P0��L'��Τ�X�I8S�}X��I l
2�*xTT��Z��S����Fx�P
�u�����/�h8Yf�;g�G�VowƟ�2C�e�,�Zz�����r
��":KW�R�v��92#���J�L�g̗���zT�kd��,����+��	0n
{p� )�Z��WjѪ��&���0�X�(�W��Ȥ�47���S}�u揊T:�B��{2xs����k�Eob�و��Sf�}P1fv�!��N�C��Ug���t���l�kWⳉ�>dN!<�K��I{+�-�ٶ/�����dkp���f(J���c8<x�u�褻͕އ��{�������O�&	�k������潞���-]~�Y0�w�n��NL����s�аZo��G����x���Uǵ���N<��Fԛ�,pВ� c��ߑ�9[1�Z�1^6.��7����Z�o����N�9�Bwr���,w�I�i֋��8�o6�s)fR��5��9x1�K��U���:���hh�Q���w��d�t��Р,)t�W���%m�ȕsx��L���1��{4'�Z�^ -\����
k�h/��;oLE��\v{e�;U�]Û��=���<�s�.��
��K�H6��@2n�W���ȺB�z!��8��$���s��Z�\��T�Jq	F�J�5&�u��*f�CiJ4�ue��2UF	���q}XnM�J��o���F���>j�qS���P��=��'�֩�hO�u�]�(Gđ['�7{����O}�����*�Y�@�w]3�A��C<�2��Q�0��N'
��`���E��볔��z�u�+[ZR����{��k��H���wlh�I��z���MS
��w		aYϏ�\���%�#��ɚe�˦�[����"#7q�\�����n����xK��$��&��1^z�6q�ߤi9��n�ߡ�������]Vz�;���|����"n����_��c�a4q +Ku)��V�R��^_����	xl�� �Ql�P��fa��-����u��DVR����7�%��󙸠[������}�Sg��`�өꑶP��Hz�Xl�OO���Cr>�dG���\c��w���~|�>K�C��O��AD�%�+�z^g�w�!�$���n����p��Ѕ��xf���� N ��d�n��\0��̈��ez���)��L�^h��M)����.�#�r�!>)��}�U=�5Ƕ�Qц����^��R4��L�fٰp�P��B�
� �ްn'^7����5��ZArܩ;��[t'��{��B�t?�~4Y{z��i��?�遼I�8�Z�*]�D��(�v�l��L>��3�|���H*U���F�7N~�7v�q�S��-r]��I$n���]/�u�Ԉ>�8�b�z��ZQ�����u�ſ���،e%1��OT�Y���o2�F��(� `����,���+��fu�k������$r�B��-4+�l�U����m���)X�1>�l���Ñt6��L2t29�p�5ؤ�`��:�C��+"�|WR�r���Y0�Oj��+��^�gׁ��5��G�:����/�5	mg܅��nB���k�	BW�'[;�Z�%���aT)8�%���CtDާ�zSrK�b��cqM}`�9�u-�*MM|&�:�1�"������d���f�5��ض�r�ї+���[kFGZ�1Bx�B�l�1�ƴ}��e�?�+�ݰ^ؕ��1x�Hy�i������O� wK^ߡ�D_�/"4�!��s�r2��ٕ7I=N���d���R,8z��KI;��=4]�B%��9���H�J�~~��?�!56灲�C9cw�*4�!�N�%¬��Ha<@�\�g�_�Z����O���}�q��q��-��T�Z�*�<��ŐE`v{�nݕ���d��GW����oW��*хaǵ�N�;�p�\�f3��s5��!���q�7�cˉ!����>��ck�DhB�K��w�
�FDr|J��j���8D�od�Q6����	�$_D-=-R(X=���w22���=R�=��k��Z_�*O����G���6��L��	 ����ct:��:�iCp���dI��������\�f�3�c�l��>VA|�W�6<�V��PF8M��8�NVwǲq�6��v�g�M�[+VK���U���3��׼�H�{џ��5������l������X�d���2���h
ňutQW�_�X���B{~�'�9�m����QM�0�nl7���*�	͞x�s��=Y���Wx��=��F�+3Z�����3�T̼�u�!��13c�	o�F-]������bv{ge�c������s:�j٩7�M�:���p+��5 xh���X5 �^;���3Zqǫ�#
9{ܢ
Q���
R�<F�da��,��:��b�c����y@�w�z�a�&�6$�B���1 $pm�&_�Z��x��L���T� o��來zXW+�$�R+��Ą�����Ze��v]��rqǬr[��YK�3���"�7�`��Ե�5�u��B�a$M{�M�<��ͷ�5�w�h��:)�4]�D���ee��	�r�q3lsa�+>��d;a�.��:aGx����ڿn�~��F��hL͡=]��ucm�Rn"r �r�]�'N�u͌�=��8�bK2��@�{s5�"���,*[]���`ׅ�r�4`«m�Ko"1C=[�2�.��[r6��{�x<.�K�U�LЖ�J�̍��Rd��z��#3�cq)Z��\1�/�X�7���b�vB8&6�^��>�Fӱ�9Wя|`P������PnaL� *�0o��o�m���c���툟�����(�m<��&L�	þ���w\c��V�����K�y:�<�m5�1���+���A���Xc�i�eС�u�҃���%�ǣ��$�*�`��~�f(�#�C�/�^�D1���S�0�3� �}� m�����@�f�^����A0��SJh4�iY:&�n�9���
/퇤�Y�e���%��tT�2�svy`�.��c�дb$��>_w	��tb'�7��h^#�EzB���|�-�r����1�֘�ޣ�OR�n�D���)��K�"B'�v!ls�ݓ�u4���d�)V�V�ǣB:z��/c	�5+)���g��x��V�@�f�>K�܀m+�֐��[I=T鄁T����ϟ�|��
��\ϻ�މ^�&��Ã=�v1N�uw�*LbB�k�/�E^S'��2@�q��1(07��%=�ݰ�:��>X��.�8�U-�C��s�AJ"�{�X�p�6��� m�|����K-gb��a��m&t�J��)m�W�\��8%���zz��r����nRo��q�"*עT�ˈ馌9z�S�y;8�8<�Y�йr)�{�[n|̽�#�ab�b�8�M��eU�A�M�'\�����ņ���2�w��U�آ�9+��aD�.EP�X	��:;	�~�1�/���)<��k0_'���}�2�Z�������K�����)�������kCK��C��c�U+��ޥ>�׆��7Fj#J���M����f6t���"�T�t�˭�tux/�t���	Ց�_�������λ��&MBySuc�y]kے�:q��m �E��6=^��d������τ�j<�nL�bh��H�
�����<�����}C�G2�)�L�|����đ���9t���.�"I8�C����&���I�ɋ�`�X�=�RJ2�5��3�a�>�;0�e��U>���p�mS�	5�1���XZ.�4�ʈ�pO��1��d+���^s�m�'�&y�ز���H����Ty�Jp1�C�����)��� zܱ��P����t&�3�>��֔XeD|:|ݔ���J�RP��8V&D3�##�z�mX�rUm9�Ϝ��1-EI�1�C����X���%yG.H�� ���{�nWn���e��/����ׇ�A���Q��S�{����;�tr[��+�NYԨX�H��>�M?��o{��	�P���� ���ڠЋA]�4���g0�_[¿E+z颶C7jb�7���*'��� �������٥�������Y�#B�i��'O�|��M�V3�i���*(3!�2k}�)\m�K�lk[�G�!)�M}S��(5Nc��i]lC2�������&��W�^���;����&�	<E>��:��T��A�*����l5b�B�l�:�W7�1��"3A๥�u����l<�O2���І����+7����Ĉ�u���5�-�=-�A:��.!��u�(�cn��.�\1mؤq�F�q���Rfr�6AE��-��t*Y�iМ��l�+l6�v2\��[�q� iNzԗ-�{_�u~���Z*>[]�5a�4i�5n�Q�\~e�hWjh��¿xdh_�/Z����P	��/Ɖ�#���R�w��Ӓ��b�1Ɉ��a�
�p�l��8����9!�9��>�:�c��C1ׯ]���`gʚ��"��;0��x�;$W�tR�y�4�Q$w���t9}�@���ٕ�߰jf�k�g�a��#���^��_>[��F���lx����`��2��g�ۇ�U��*����c=Y�0=�^	9�.=ĈPJU������®�w)�։��怄ln!\�)3�V-r2��\+N�:��P$�;AY�JFg�M��S��x�����18�ı�$�����ɪ d�8 eD�0|gaB��yT�I��e{?��_�����=�"6a��\���+����}|0���t,'�S�~�/Qe�m���]�۪[sבa�~dr���O��<r߽�Ȳ�>�� �`����}��2�mDkh���~I7}�B�Q�ԯ���ͣԤXM�6j�M�i� r1f�p�hL��!C�IŃ�����
�����V{p����
��3ؔGi�><̹��� ����IB��x�I�o��#X����0Jx�7����'�:K?�B;�j��A�g;�)�F��������ϰ�'Iz3����}@�4�����׿�t�{I��񟳫Q�y��,�䂱J����Ԙ�RwT�f�rOob��QX�N%�U{@�`����<`�]I��2�N><nj��|ΤM�cF�'k�5�[;q;fRe��f{|��I ����n����������*���ڳc��q�h5}b馻Q��6G,a��p6�Pu�������ݓ^�Ο����t0XCI�q�=��1+��:M*{�2~���F1_��tU��]��x -�3�B������/�#ǁ�1���_��/�E ��B�z[���P� }��4�M0��M� �k� 3ac#˥E�P*]Ĉ�2��y����+-�fw�9����KՆ��*^�K}"8�!�P�l��
��K��06�7��TA]��|�kÑ ����	��)�[��}��l���76�ZR������ܘl��x-�����#C�6<Ѩ�>oF�֫gn�A)�zCu�r&�����ӛ0�Q�-�_�{�~�4�c���leQ�}M�~���f���������)@�}��]�b�s�Zb����	�� ��'��v]WѲ�� .ˎ��T�2De�t�W��KO�-Y�%�%�j)�䌌Nd��u�吷����~�g� \�ظ6Z��)jï��rȕ>�\Mڙ��Yk�	����D�K_�a�b��s��	�j�'��A��^����`Ōs�Cj��5E�� ��±t��5���Z�vq��������c�Om+
{\�,�Nt���in��\.���Z_�5��ɼ�h����!�}�����MUs@�옢N� E�u?5<�^4)�	a{C���r�fۆ�'=:�`���P��g����&L�gB^L��U:�zW!v����'�C}�?���A��J��	��]jY�T��m���d�܌)������2��E��H��$�'2�a�{���S�n��ύ��>U�R��0�;5�s�������߼}Ì�9� ��3�}Z,��6$Ȉ��|��s�>@4xo�F1&3�0_op�bl���ZUI��p<����3:��Ɗ
���lP�D�D�q��^�uSHi��Wo��;F�A��sx���<��_xGxB��k��v�Ǚ��=�E35�X�ޕ����z�XP�LA�k}�V�O�{J���=̨rJ��gl��*��t�(P���nA�qP��0�CUW��9ƌ���{��R9G}=a�q���unFH���98�����w}�d��4�_=]=�2����<@SB���E/�ڷx�ɵ�[]R���ېv]v����L�q���0&+1���A[\��'��p��iN
O�o����r��zĂ!SNJK$���H���`�W���[�k��)��=D頽���H^�2�-�s�ު,��ֶ,�o��t��{(R���d8�y���Ƶ|@�Ǐ�B"F�k~�W>/a�ά�R�dV��8�(]�e��Ǩ+_������/o���U!�b�\��f,1k�
nJ BR9<ҧ�mil���X瞆�s�>�W���0���_%�Ъ�r�����3��")�m��KI��;�2�"���'G(.A��#��.
C/�քܥ�t<w��������P5M�A�6�zo'��}3^0Z_��1_GDk8�e�GtN��if�t]i��}�'ʩ�����/�}��6r{䥛p���u%{��Ӱ��UY-+NB`۝����UQ+/Y5�Z���Z��2�ݮ*xq�5#�y�^hت���X���2��W�&�Z�y�ox�!��v����5���׮��]K�^�h'lT�6��Bķ�i��T�")����M�H�S��Yaz�_놮KU����B�l}0�bd����B�	�f���V�-��'^b5�qwI!襙X��Ε�g=s�k�,{�S��z�[���rͽ�gU	���\����~��^��{@��Z�=���*Y��+L!�T؃��c��Y�{�����cVW-�f�qnd�Xco�&���'i��jM�.���n��j�ǡ�,��yq�ޮ6r�(H��h�&�ލ�G�_�i�b�����H�ݙ�EԪ]�5��"����%T2�q�M���z������
m��eÃ9ӓZv�8�t����&���usy��঄�����F�I���Sp�f�����V1x�8|P݅�)\Ւ6��w�[��{#Z~�漾�z*%j��.�v�[���񵤭���35ú�ق�R���Jq�7-}3`�t�ځ�\�t��i�QWM�P��a� �K�����s����P���?%��I�/��j)�-;X�cg���� nF�ͥ�^D��U�jI�t��X@���z�k��!@,ρ^�Quף4��^��w�Z��q�,O7߱��2�z�58�zc��`c5�S����6��c���V���y�K�֣�'��!JJ{a�X3��3�+JR�Q���`�RtY��JWxQ��N��+�%�0`�BA!�j����4#aHܰ׺t&|M��Mm6�9���o�{eK8�����H�#k���U��g6���� m����Y�`dT Ѡ�Ɖ��r��N�Hv	+�.�0DC�cm�G����K&���_u(̍��	���VZa���s�����i���F��;������&d�']��z'�jK\S��Rգ�2�J� w�b���u����l����1�E�4�qw��Zy��%]���	6v
%,,LP�@EjY ��10�I�!��=K���GKf�a#7�%Swݧ�HQ-�����mǬ�=Q���I#�n�����"z��qx�2���e'Ԥ�<Q	�tS�i�6[FveEO+�ioϏcn?~t�����d��D�A�B%ЧO_��a�M�K9��aR�)�|*|q>��ؒc��OѶ�ɒX��s9/l+m!od{�n�B�v�������#0�jm�Jhg�㮅��+ªM�"��$1gR����K:V�?��ڍ����\�BW.5-�-^nm��OQ�X�������n.R�=q&?��э��Hh�穵mOڜcF���xNvົ�����ۿ�����R����3����M�fBhP9�XC?'G���`D�Λ���rK5�C��W�H%�Na�=1��x���q��\�}�}��.��)�9<����q�?��S�IT�I����8�����nz2ؒ�?��*�g�ø�뷭�dc
��P�l����i�]��^�tRbǳBi�3W�νvA��3�Gj���+�?f���A�,�|�*�L��+6���o��Ǐqfн��@�rwX��O�o����B�>9��Ww��W<XBy͊%jpM�D��2i��j!fl�i�])�ҎA�B9n#�l~OO?��#a7V��F0��羼��h���)\3��{�q�o�0� ��̒�g5����{<�G���H#_p`}=��	�/aC�[%�1M�l;��)޲��/���{��rhڂ9I�b?/1PwK8$v\ԗlҚ!��&�i��ԏY���(
�KY���{`��봷��a���d����Mîʖ�\��V�l	y���W���:u�n[�ƞ�'�,,,���X�}�)�Uq8Ǉ�,s��
�r(�:�u��i�N�!"�>����k��s���-��C�ҕ�0���,oz�}-�3Q�E��Cū��nA��p�{��XCR��b����F5z������?V�|�󼮢8�#��My�В�T�o*9�qh�%wD%����5'i�S�szd��(YSB����EF�Ɋ`D(�8��}��ڋ�����s�D�<�Z�x�Y�䵊��u8*�஧ւ�aSe
X��OY�N&C/��R~�i�gYKE��i3��ν3��I�~��A��N#+�`�Ia��&P,���M����q�������GF�"̶Z#+���VTQ���G�Y
H���^�y���F�60��x]iB��׻Ĕ߻��5
Cʪ�D�j��!�Y�#�l�~'JVI�7��1�KP[���<#W���������o��ŉ/+hI��XL�t��6b�\�4t����c��׊�cnG�1�ɦh�ֱ��P�3���gY��kI��KiZư��O�Pr=t��w��`/�\b*u���#���ߑ����czh��6弸�I�����ׅ0Zz<��v�m����g�ٞ�����r����%qm>�Z�,>2��0Ɠ��q� ��Ac�:��=�;c<�*TI@�?�m߬�~�M�f��^�v��^�`�8�5ε���9���Y{/��Ү�w5b�sY�z���<*�b���[�ǟ��z�"�zͪh<@�8�=�S�e�ě�N;�"������?��a���a�;�aD_M{e��
�6Q߆�f���4W/K�'8yA�xf�H֝�vwxj)��T|��kˋ�Cdx�x��I�#�h=-����$ �~]���6چ�LT.y��s.>7Pki��D�q��_��jh��Rq��1����ky`�6�{I�ys���N���hq[mztWC#��	�j1�ֶR1���.��3CE���ġAQ��y���S��	�sa�9=Rc�>(qOOo��L�f?~�P �4���~G�-G��t�+� �])"���a�$��K�1�f��.R0�����2��tY-�]kҭn�>����f�ΰ�/�=e�=YC���Vw���Cd���,�eVCG%�b��ʲ�5��xhqb.�V����T�;(I|U��5�����5�H��}����+C�_m�7���k`�;"x�V�|�XF9Gw�)�,->$�,�f�o�G	�����9b�¡��c	�|U��S���^-���˼�K��c(����x8�oq�6	WG�dH��q��=O���z��z||�/�C@�����J�Ǝ�]7$�� i<�z�T�6!��f길����4�Xt��=��z6Y� O­����00��Pinު����^PP�0'�]B��oY�%3̤���E�n�B&����c���k,�^�Z��Y�$����Qk�6�#�,�<��3�2�IB��[���0Zg�p��B���+Ӧ�^���Շ]j�b\����g� T���k�S����A�|2��nJQ�ʸ����n��QJkJ@g�g����O?�P־��E��>3�Y��fJm�^pM-х'@�~N��	�^�>�d����)�	�Ɍk1Y~�	�Mb��Ҽ=-?����l ��d2���ރ���}n�Y׌�-v��r��ƈ���3�*�1&��F�^[�m2��	û£��.����V�?HإS�,�����L�����wޖ����:o�!����}���"�y��di�Ξ��Vb�U��a޻���r��`�@�� ���?G�{h�>1�zd���]�Z ��^��x�n��4}_uT�	;����E���)^�s��ㇻ��%�xT�G)s��Y���E}Oc��s���9�'Kԡ1�?���%�ЁHZخ
IH&$�{�p�N�����M��FB�㇏����0ce��RV;_�
�:NͿ���t����ߑ'�*�5��/(O�&.��p�o�9ޭݗ�����=���ZA�r�:��Ґ��o��rVޜ/�Z�s��EW,�\�	�c�ƒ:�Mh�ɕ�6����f6�{o�#TG���03���X��F�1���(��
�5�f�ZȞ
��v����Ε	���:T1c&�&��`L�AHla�۷s��πt?8ٝ`�&��%`��;ER��/��; \G�4���e��.�\{N䜺� =cy4���=�]z�+�9�i�S��m���N�y��킔Dl�%�Lȷ� �ê��;hY��@Fq���Y�c|�E�����0�c��6�3�Bz������X�S%V:���2��}��{6�#<�{ó�?�|�P"|�Cl<񙕵r-��4⡷�2��}��B��{iq��:�SjtP���5�o��j[_����rN�l��z�ޕ1[�#l�r.��������Ŕ��=���~wwx�q��'����x���#�P��z�2�M�BQpQ�hL'�Ug��<�B��i;Ԭ�zZcA�"c��}kw�[hBbB߽}��»��t��Cie({y��ǣ��Sb���M�	w&��V 'W�	�VVRʧ$�hۮ�ɐu��=6��G�D�19�!�+�Hʥ&=�Ge�Y6����Â���f�u%�<[Cʰq�|���U���v0�ȑ�=+߃�8�E��=Rx�y��{�A8Xo�W����ujwR!�{}���L����O����8�g��X��V?l�q�H�zdP�?���Q�����k�?��ShD�f~>��ꔴkڱ4�b(��~O��	`]l�H sqVc?����a蠫@���{ƨ�}�+��V�E�����/hW���q^����/���8�ZUB^8X�YFv���ܭ��!�dB���P~QW�x�t�ꙺ��y��e���!m�y�Ү���7w�BQ��]qQ�L�{�C�]w����>($:����\�.)/��z�  ��&O1cR�B~O^DܠXx��9{�Ж��*�r�
w�l� {]�����5�7�?!6F
�kٳ1Ó�Y��d�	H�Q�*���9������ڬ$�E���b����ř���¨[����`%v&y�6��J���UnpV{Q�$8���'ݲ	�)��~�k�
q9�)8w��2�N����~K��v��g��a���t�t�L���_g_xR�N� �����v��W9�N�{���{`n(�3nF�O��؝��� fIcڧ��0��,�(��+�`�Zv�#�e����X��?��f�����q�f�3�3ߑ%>������i�f
��?Ǿ��}"�D�lkuY�5��)����dT,bL6�nü��ߩd12����m��Օ�[\���F��:��v5�7$sg�^5��E�VZS))����Ә��-KK�r��+U@=#!�W���z-�c���z9�"�4h�PIὒ��4���B��؋naMD�#�Z��͜���d�����8�k��3�Φ�PH!VHY;�b�m1S�T)7O�h�ߛ����~�����4dy��/$����������Z[���(kiQY����R�����megWDȤcЛ"����4S#��@K��d�v�c:�sf;(d�g���l�'��2��g�y���-���xP��%��ı�������}�hG�Yx�U��^;�Z�h����k�����u%ik�P|���9X���~c���C�Q�a�/�0O"9�8�{�0��c.�9�H�e�d�����d
��1�NBkk�A�Ib;�CVu�*M^�0"�����݂�Z$(ݴ_��Uc�ڿ���L>w�W�'�/6���G��1�*FzgL�2��Ċ^ik�7�'a#!b�Oc-~fCi��O�4:7	��zQ�x��GvwׅІnƉ�T/�'�mVqǞ[xl!�<%^8ٵJ��#��m��@U8Zء�_Xs��.�$��9���P���T-˫y�5D��N9!��8�B��x<R!�� 9��@-�Q��St}_���ɿ��\��E�6eR�J�؜0��F������K�N�nqϵY�����5/|������x�sj�f���u|��5���e�D�w����i4�v����@���b��q��j���Oq_��M��C��4X���Eoj��uQ��U�*�8�����G��c��۞h(�ȉ���:>�:�w�Hɝ��#e�Ae��E�@�f(����c�DϹ?������f�2�j��5�
1/8T����w��S�Y���-��u����-����K��-Vi�=:~��ih��W�������Л���p�&���y%7[;�J����%��a��n���X|3� ��R4�d�����~|QS�Z�����91TׯW����s�1To��l�[f4ݣ��VٛqF�z�z���p�w��>�o]�\p���ȴN������K'�w�a�Z@�0�d���VE�k��(e<s�P��-	���͋�x���V����)�ww:�oJF�:֖	2�"���}�;��_�4������}z!��9	郕ɠ!KIɘ�@�n�K��8V\S�<��ZFp�m�y (P���a}�0�
P���%�޼y���ے���WәT*^E/��-�W�R���v5�
����}��뫅� �W�z����tN�c��Sf;��3�%�����n$�;�C������k�k�{���&��L�c.������pеrBY:��D;�C�V��&D��eD�m��W���_/A�����ʖ�`Z��*��*�6#�eUHKYdD�@C��>Mm���u�+�Iok؝H -�|~Sا~��I̺;\�����`�X�r�����&��zbe�[��I$n���}�~Nqwv�!���On����=�G�����8(�_���5��p�a]c����B:�*i��>�n}]��B>܍%+��\�y�4l�M�n\7��}�š�7��־"��2�5'���>�T\7�h�zt]I�Ͻ�|`����V��k�Z�,|6��'��M�$�Q'<�i'{	�6,����T��S�7���L�?D�Ǹ>�u>I��mЭ��OuŰם��a�Ē�6��Sm5�i�N8R��se�-H6�.�J\��~��F�4�/��U>�A�����Se֗�T/��.Uq|����-��M��Э�����j跮��qI��I^.�`D�ŜU��y(�2�\@Y�+׵��86\��
���w��w%���Q3�;�٬6.T_:��}Є�H��
z<��y�5Y(Ā{m*74+|_C+�!>�X��K&�w��,��?���\9c>�%n�Rf��sS��F�s��~T��u�pSGY������7�a��
D��|��h6�S�%^k�Ja���a����P~ؑ3�T_yF2��n���t�TU"4rR�x�twJ�-:lN��D,.8��Op38��4����*%Y�\����!��P�ߌ:�F�Q�#x������nL�SVS��û�ιޣU�U�����5
�
����[�}��4͆���s�퓟�g�|��_�� :*�(�0ts����_�Ҷ}�{ۻ��{�Ta��i�ڤ6���H=�mx�F&��щ���Qr�}X2W�]���
��#��+�z����2t)e-�::���E9/�f���9*4�gɎ�>��<%}B��A�L��75�,����YF��
guA��iO�A�Y�W�|*']�h�ؚ%`~jmsa������� ��;�+T�����9�g��V>m�|��b��8�aw�ʻ]�ۇ1��D����Z�Y��+���d{�~�^�|�q&����z�`!XFO�2�W�����6�{��-��ޅB?��9ڌ�Ӽ�(��B�������Ͽ�g�S����/�$�L��m"��ʪ�#hs���<������!5����4�U���������}����Qd�Iz�.p���汣ȷ��MZaH?~�{�>J�$���iG�:Q$�1��V˛�"j"�fM�n�l�"�)"��2eL����B��|*)������*���~3�b~�/]��@�62��o�Q��j@�ƃ$� cl2��%������	�i��IE���Eڈg�;��_�Jya��u���H���ޙ�y�5s$ZmQ�ՙT�w�QH��,u�m�UNp�0���txd�ґ$�X��G^,�"��Ncf��<��]��q������޾��)��8�y�#bv��1Fn[���"]$�ύ
Z7^k$���z�j*ma�p��:1Yϯ���/��j���F�I�R���nWF��~�1ĵt��*��=��c���YMԜ�v��5I�4RuC� ��/�	���6�a��7�F��)��b1����.��<[7�ks5GQ=%\h��}>O1O%u���P�����䔢��:-�;p��3���K�\{Q,��]��p�p���sx欻'��xg�VE3��X�6���6ڃ�L�]왧��,�=YJ�ɳ�����e�[��_/=U%�Zl���������x��/�&�d�GS���eҐJ��d|]Yq\�Rp����ʆWC�r����9�U�i�Tl�q�ֈ=�=�E��M��e�Kqݱ�'�+2�R[,dz��X���6��Ќ�$��Օ������y��uvJ����|���u4њ����Bi��<�`�5`�O\64A�w�}�k���hU=� F߮�e|R�MB���N�as`C��Q����HQ�]���]�&�p���ZU�`�1��?�&>�g��n�HCJ��S���zZG]�L`�a̟�(��nYy��T{3XcWxW'�Ipw���e����k�5�n�-4
6/��~,n׌�@[8��n0���Ѽ���
�u����
�ob>�*@	~;F%%�Z�+��9Ao5q���U?�i��H
�!���_%�qv�v6:pa=�W�D��^��0�7��M��F��>[���mkj�t�7���~�N��R/,7QgP]������2(��7�^i�&*=`�dH��Vf֭�]u�T����q-իY��^	��!i{�0�e�eRU�3�V�"f��>���'n�����!� 媝�	�:";YJB^x{)���1Ύ�P2l�1Tf��rC?�g!���^����ㅺit*}P�!9�s�5���}���w�v�T(p�:Ӭ����!�\.9���p��]s�q� ��7�i�g7o��!V��e��@0���t�>�)<��\���K��2m6.�==�VV������������%��8\�;y�(�dRjJ��Y��$�Ǻ���6�t<�dY�rH�կ)L��9(Y�5��͎B���X�=Z&2�B[2/,�\f̛!�%�NM�n��v���:��!��1�tJn*0 U�Θa{�X?�K}=�!7�X�O���Q8l����Ï�~{�~�}O������6�x�6��e�m`�#�?J#)����1����5��Ef0����'&ssm��x�F�='V3�^�	hэh�!/NrQI��Z��=/�f��Ъ��|P���^����F}��,��v��E��Z��}�vЬ�����[骖:lZ�R\�D�b$7����l���a^��Ù\�TP�{O"���Fԡ,<J��v�XpF��}��z��E`U���9[K���q���6'������1Ϣ�e��k���ȋl�#2W����ʹ��ʫ��BS��=zm�u�J#�����h��wKd7�9���v�xG���� ��͊"Q�:Q�XT��i�$���Ö�JY���eJA���1
�M�7�{o�YW!?�_ÈU����H6������oe���bL_��	����	�R1˯�Ε}�!ǂ��<����~�/.�Ph�Ev�"�-m'�x����R�^`�f�Ș����W���b��b=ٵ�3:3Ί�.�
��y�+%�$=�^ߑ=U�/�kp.gr-qW���*���7����}z̬1^�%f�p��-��3�M"�K�8�"�S<=j޹p\7���%��L���2����a{�����6�Wz��ֆ��k��:���i5<�Q�SЋU߫�Ԓ�|�W�i+�3A�E��������`�c�9�l�����>����O�&[,��gH!��̹IĦ�*�=Lqb�F�! ��	K����\�U�y�~��8.+u,Z/k`�I'�1��j����:8�cDyd��.�]qk&X���AM���\���쟖R����H1�����u�*�I4/�k��}��E�h����O[��!M�S	�>��6A�fX\���В�T���A�{S�c���w����MD�2��.�!I���(�L�أ�Ѳq������Xlͨ�.��B]S|����&o[؁Ę�Zt6�+�7����4�P��֌}��8��3gy� |�O���U0���!!C΁)1Q��_����5��ֵ��ŵ���j^�n ���TBh�؇i$1p�$��ưW�=���������d�kR�o���ZֱT&���nu:�UZO��7��."R��a,�#7-+�xHY��B�!�lr�#u��k�#P��ō��na셭[L�;Dh���Io�(�eY%k���a���vgH]�ϊ�Je��r�(
~H�&J;�vn�\9ن�nҫuG�1+j/�9j�`��ʁac�.�q���:d��G�H8_�fĝU��(~�}A��M�ԏ��H��K'>�K��4��[�%B%4Jzy�[U讐���6�
�*#nc\�F|_z-��Gͤ��15�w�����9�=��ѳ��5 �����5U4�4�$�fk�i�):!�$����r����7���:�U�*�1I�դ�X��1V����z�V(p���.H�Ŧ ������� ��a��AI
�(!�L���߃[D����̈́QU�9�ŐsU֬�6�nӖ������OJJE��kp�,�����IWܚ�Ʃ���ېP��@N��7{�[��x�������1�dp��þ
�8afm�0���0�4���:��'�4>5�7�^c�歹�Z#�i�v�ɚ��岦����mM�U�*�p�%Yh���-chЊ"�����P92��f��b��a�a�zkc����G8$��MO�X���{;q�\Uv}kJ��eۄ�k�˿iqӑ4ٞ�^s~�+�*K��06آ��yΌ��q(/R�������r��'3�>�������-����ʼ����b
���O9.�Y���3!o̵��� ���
[g��4��>�((���S�9������=�榲�$6�6��ņ�uͦ����M�
k�}�f����B�����ӳ����ن�&U��XYm��5��x��(7��m����e�{��1z�*.L-z_^�S�=�c,a�>�����-�uG^��G���a��Y����s��5e��_4M�5�/�#0Wu�}�Z�]D�Y�� ��a ����܊p��&�F�w�2!��U��Kx����"��K��Ѐ�r�H%C~n��-�w��.��G/�G���_�iM`k?��xm����I��O�8��!��poT;[������t�1�k-��r��Z��u��H�)��<���Q^@�1�q$dd�ƴZ[C*kFT<Hg����Zр�C���L�t�iڶ	���{@>.Ul�Y�L2lF|R��' �>�}�v�����Ơ���:�	pOI�B�ȫ0�����/�!�y��D_�� �qz��c<1ASQ���f�U_�et�Ч!�c�Ә��ء k�G&����>��q).�/K���,�c���5�QV�ZPG�:����F~b�?(+����6q=(���x��5u�2M'w�rҡ��+��vUC@γC�6YaX��Y�Х�5g*ս���Gi4{��	QYkRS��Z!8O�FF�]
�<ilUq���"��g�O쪬<���p��p?��
�~��pwR��wi0�,��3�C���ݜ{w�Ad�u�4t���w�0�|>}�|���I!�ݒ��}�P�/����C����QZ�\�47<`�?�jx��麉�(�����ZY8��>[)ª�!E2��lN�Wzk��4�ɬa�W�lW3�IN
��v��;��:1Z��=.c1�O�*7�2  ��IDAT�I	gݗ&𧁧R���0z��L�n�~�F&b�~�y��Lq�7�(#<��J|n&�_o�����2г��2c�
�8:�p1������#m���"w�4$�o;n�/#q\��W�6��7r#���7����a��&��s��N*��0�A�G�c�q>��g*he�ɍ=l���H��F��gaC*�bR`<�)�FU����K��u��ڷ�خ�l�:al�q�Y1�'������"�E�_�h������8�k@n��8�	�>fn�bCj���N�Q��"T�t����z��d�x�u�0����f3������%�l���Wp'[�=R�s��W�%�^��v�	7#���;��0>s@5�+����J��9h�]�����'�9�,d��x�7�\ϔ�<ǜv�}%���5Hc[�̚��^:���Yp\�U��;e����p�_+,z!�׺�嫇��L���X�<A����6 ��X�>�{�T��ǲ.�Di������.�ME��±�]vv�U��f�!嵆�����k5#NVc�7�r$���z|��)�����a
��XP��˓�b�E�^K�n1c�{��u� ��}u��3�]���<x�=�%����9�Ð���K�EU�̚��l<W��a�����Gf���aW�&Ɂ��i_�2ޘ����
^c�P!#{������Z���e��ƺ���1.wgRUz�{͙�Ƕ��,JN�of&��e�U�+ܕ��>���`����W����/�Z�<'��Φ..a��cp�:��p�d��N�b!e]skޏ�.������y��5+�&��!�,��4�:]]	y�r�i\�ɶ{>���Kn�=���u �e����x��揼��y-Z4K�ć�Ȋ���XkGE���ll��P&yRu�>��R��MM�&P�@-����%�� n��4�P��N�g5����"CX����)*�>�)л�6ɘY,�fL|���M"߁�x-tL�t���=�	o�M��Ħ���r�� �c�>�+�cx!.4zD7��\H�E�Y�(ocH�wFh4\�Rd�!L��.Խ�!�1��u�z�����ڷ�f�JқQ��\;Үkӎ�\U��v��2�ֶ� b��#�U�9z�	�(������g�����Â;�b3�@�5
\�f��$Ù��N�<6/��_Iȿ�nMB�cЋR%��	}?���2�Ӎ5���n'c7G�g])�7��KZY��4K�j�8�����XP�nUVњ���k��K�+��4���G���T�m]ˋ94+�V��=�$n&�����i�7~����V�Bm��\�m�c%21&E��wڤ�u(�X0>��p����<-�O$��J��p�0�.�>���`$��͒<| ���0�3U����3Uo0�j���-Z�N�\!�z���=x(/��<��>M��Cφ��m�>;�Ƴ��e���	u�}���t�/�ӀP��m�^���;k>y��Exw��`�v	�
�@&x>ǁ�1��^<
�| �T�㏯.D�zS[�0S��!�#������r�z����x�aLN�=喓�.�6�-eω�93��>I]ҫ�I�s��:xzO��|Pl��qx~�ؖ�Nʜ� �����:R��>��ub�>�(�8b�+�A]�1���cn����`�� Zܺ�D��8��p����n�7H�Z���C�2�uBX=�Z?/�j[o5#Gf��ݼ0��}��i���ڝ׉>�kC��.�I���t�e8ZCϵz�2�7Y�w������6�]z��q<����xNh+�P�D���M����sYB����~��w��N�H]�ۄAkQ��T�����$�"x�t��BW���g�� F��At���5�'�+�*x�#1��Mw�Tl�E^��ۉ�8,��f`lHC�3B�k�#0�녛���ND�c�$R���������5�cN�z�u���em<R&؍ɭ*8��HgM�B^�m'究�9D���1a���K�}QYbTN]��5W�o'�J(E�h��CtR����voHO1>-��:���u�"#�v��0ϠȆ�n�m��h��S��r�H��y�t]�'��J>;�p�s�*��-miCc��c=l�Ԩ��AX �]���M�T�6�V�F�=�Z�z��l�/��1}Ͱ�qgH�xC���^�0T~YU�	x�+y�_xy�:]]:��`]t��[Wr���d�dR���݉��?��p��JaF6h� B��s<%�p�x�G��'�YQj�!���Ώ�=��bL&a��5)~�^O�kU��#���Lp��V�N���C�8.FM��X2��w�׮zC�*f�F%]�V�1�!�7Dh�1�<ᥘ���v�hAa� ŵYQs8P��^na\�q`�3(��!�mܹϱ�V�à�n&.W�G�p����+�t�5�dmн�.��ޠ]_!�K꘰@c��\;'����Q�a���{q�8b�gŽ��(�̍{c�*qV�.�F�� X��Q"���+�;�$��f!�g/^%�=)�O�],�`��%J�[Ke�zTe�3�%�ۅ�~,�El���2��~{َ�1�BEX�E�gz��7X�_�<yįc���wn�0g��^�����%C�I����fVk&2�m;%ld�l� ��î���h<�������d5����$Gf{*�bC���",,������Z3��K����N����@G_�.n��|;���I��Jщ����F�je�L-�{E9����̯y����N�sgo�{���8�1����Y��e�����m��������>��>�����f]��gQM��^X�i_7@���j�m�U��Q*_�;�Z���z�!܋�7j�{�������"y����!g ګ�?)b}�U��UF�*/��!ͧ��ck�� ��wf�}�M��A /xʪ;+h�Lp�2܍�NcF
<���{W��۝Gk�7�eu+.��x�A�ג�9�@J7@�A3%�u�X�jX'[��c:E+6XZ�;Q�����i������a��g/�S/���H��:��S$�񸸙Ų�UF�AThg�����!�1,ǝ�k�>�D�.�%V�������$}�&�r���1AEC���^��mO�>�BC�������	RQBi���~�^���󅽚�e:T����)G���p�gV���h�02z�H�ﬤ彲
��ۭ�9�][�z��S���1����b<�+����G)���0�����3��팷�v�XA��Y����H��kF�U������|�����5��7�N��󚞰&�d�z�e�� �ˀ7!#����Z�G�o���yV�����A����+���pv�vM<�J��s�"��n1��@-��CN��t�#�9�!�58��Om0����)^I^x}������m�c��W��k�E9ؗkI�"OLV�=��������q�5���E�+�N�r'�p]�L_&m�M�מ���gx}�F�5�j��޴&���F����r����h=�fa�f2�aj�)D{�(�鶫� �Y�2UK?��^$~���e_�y�3܉eu5i��Xj�ƀ^N�u�>j5R���f�apCo��W�!g�ƀa"�}-w��mԻ�|�ӆB�deא���0���J�Y�����>/��tfy���G���8�ː� �'׻M5����}'�g%�9��Y��dF��65v1~�ޝ5�g9(�F)��{|��⌹�*Χ�$�u�<_v7p�x��y��� .wې�\���.�M�������0%v�V"kt*��s����	�(*p	�.����F3v�-:p+�0'�4��ܘD#�f�w�I��p3���d���J��Z������wԦR1<��lz푘����v�f^�$i���6��]1��#_Dљ�]����׼{W]`�P<��t�y��j-�"|Bx�zZ�/R,�K$b�:�4�ȋ<lx]WT��P2ۧ�9�Y�5u^�]�Xb[#MO�a�3�.S�z�3��� s�h��0 W�T-�#*�z_�W�9��Ė��]�A) �אF�L�ة��+\zivdf<!l��K8$B��s��Q�rc����A�O0����=1d��4�y{[��Q�6��F���O�Aw���k�S�����!t?��9C�Zq����R\�V�⫲Q7&�y�{��ʻx?�k5:��8�&�zTƿ��aF)��.����fCq3|��R}*r�Wş��M�Uӗ=�=>��A��<��	R�p�����U;I�y7��1�FQ�M<�.��E�o��#)L�[h�_Vvf���>t���/b�����x����TŚ��{�i�(��x�t��k/�s<�jц��%�A5�ә�w ��CX�*e&>� ^1W��7������>�cx�g��(]և���]%vL,D"T�cOh�TR�t��5BI&ov*S�%[��V��T6�G��e�ƭ�gΖ�4f�6F�=s����'�Y�/C-���2�偶~��t5z�����Pp�F��d�I�u��������t�U8��4(�nM���C6Y�L�9_��;�UO;������z䇳�I���p�7)�Tl��:�7+�SwQ���膕�]ʽ��S?a_��F���Y$���2]r��_�`տ�RMU�����(o�G����/,j���?iБO�l@^K���Z �;�N}M:����rH1P��xw�]���:�M֞��LIȹ��$���|��Yd9E��b�">�����,~d}�G1;B45]ݜkR��G[Dȕ���x>V�)７���b��=�n I�'͑5�"���`ڸ��Ŧ����M-����Ur�I��pL[��q�;�r�b�4qc�ߌ��1Rg6$��b�����SP ��p��=ZT`���N0�z:�	n�h��y>�R�O�t1�	ͦ��q��i�O���	/,�u.(Mb��C��!|2C�/��:i�f<�pΞ��f�]>)���N)�6r��F�z}h���+@��n6�2�h�=�;l�dwu�N9��e�[MB����f� q݄�R"؆�S��tn��?����ʃ����Q����i�����RHL��ӓ�C��;�	K�	�!۪��"I�w�G1��~�'�CD.�h��B�gPO�X-4R�����G	����	����"���v����e��������w�^)u��/G��x`��@� A^H��\a����L��6�n�D1q*�F�D�X�O?�l��47w�|'�?˦����W�1�O����<���c���D�"}�g�w��߉�0FT�	�J3�}��〷�G8��M�
�:��r�`�	L[33�����o�H�$l*]XP��Uįm������E�f�	��L�u�L���M;�L]�N ~�nM0��DA#b���u�p�G�������R;��AL��b��s�M����=xpk� ?j�#��@�g�0I;�v-1٦��'(M����8>������5���h��;��MP�Ă�����l�E�xB��T8@�1�t�1ȭ��� ������'�{Nx�x�>FӡF�����-BUE�#� )�V�|��`����X�f�8O�p/��E�v��E�?��Q����f�s���#�[6�ys�6�A[��zX誅�^$l������q�@)9����^��t�	��ɪ�h$�j�u�
�.EE�(��9Qm��kD(���$ޟ�fd&��y�}�q4Л- {��#���-Ռ*mP���Ml詡�OX���wj�*�Ǔ�}�7�hgޡ��!�z`�Vd��j�lE)��p���~�K��(�5��d_σOcJ�ٌ����L9?�{^+J{�@�Տ������bh R�!ve�1N��D�>H�V�fS'�a��@������{Vq��$e2]�q~�|@����ц��XDĔ�Af%;Zy��y�͹��S����0����Vv9_���٨�|���S�.vh%〳�h��X��ٜD������kRĢ�����*�1���_Ս���K�qz?٦"6<�y�6A�҃��$��ya ��/�]V�6��y�@̴��}Lc�������S=��ؘ��f�US���& e@�h�w��>]"2A�-ǑTC��;�T�HkN��nȉ���R�C�3�� u�徺�:9@P�� q_,�.��{M̸�&��5PKjw{T8��M��t��m3WǻEڂY�nL!�*�������4��l� Iќy��7T5��ڥB�ۃ!�Jb��!׀e�o��l+�ӎ���v��0
e�����͈�`b�&�s��m�vtϝK�3?�|��s���3	��I��#:��B�a������Ĕ��Jz��ɢt���"���1�M(��!�,�/<��c^��b��ĒyBk�t�dβ���Aw6v;��	������`��:Y�S�ObJӋ]�����&�d�K��ן�����S���ژ���)V+=�D�����?g�F/jk�dtb���"M������a��@*l��b��T�����^���$��"��Q}gI�����N)%���Κ8�I@�Y��p8�w�M�az�Q�խQt�c��p� RدJ���r�$63RM���?ޛ��^��?p��5v�EWn����j�. TgP�	 Nϴr�����{��G����L��v�Y͢�d�N�Y�`���\U�{��-L�nOL�H/�	�l�&R 3]WTD�C5����c!��9�4IHDW`���_d�P���v��+��F��+�p`b�p��o ��N���θ�"�r�NG��Y6w{ӟ.MDӽ�������1���ʖ���tϻ{�,�m>�bL+�7چ��Kz[�to�]���3�<��NW�%�!:����@#o��{t|âzѝ�b�fEυ��#5I��y����K����M�`�#�Ct,M#��#��^��f@2yb��\h�����>������ҭ�Rc��c;*���ӥ� �3�#�JOz�?H$ulHr�rI=/�*89��;�����K6�i&
;����N+���`b.յ&�6���$����c�V[�lni�F��U�3��ȇ�F�����{#R�>�J l�x����ղ��0�����>��0C%L�M���ت,���'A��xx��h�$�Ig2Khl�`��K[�\�`�X��b��;�H����`�)���yp~o�=�Nr���N�<A++)@�M�(N���lܠ�*u�:�K	?�QQ}�6�4i�dg�邩����q�1c�������DE�y襠_H��C�7xR�@�i��w�Nt�y�+<�q�l�OQO�{آO���N~���>��Ϭ�|O;��! d/,5�B������;�Ko�ҟ,,���p3bl0]s� r�úA���1��@,-���p�uK��Q�H��'"+�5�C�~����x! �� �TPp�Db7j�w��e2�ƙDŗ������͝�X��� &h�ϒ�v�f������4̃�3�w�.��Y�d���S��	�q416|ﶽln��dL�� ��rPR�x�ܝ'��
�̨�ci�10��mf�us�R�N��Dj��9	��n�!�rѵ�7�+L7��@�̷� ��3j\�$�#�ﶕf��$Q�g�Y�����A���&��<Y'"�#X�d�1���S#i脰D�Y=p�g�S�$�o��N����g��B�Ung;�@DW�_k�_��6�σ���Q��_�<?Γ����.�Ё�nK���+���-���L=BUEH�[��g�\���LR"!^%��.'����'`�`%K��l��< (DH1E{p���l���Z���C������Cc�m]�{�>�v>~���0b���y��㉁���^��~�r~��f�%���6ez��ٳ�a�OM��%ĒH&�*Q�?�gQ��ھ����q��^��&+�_ڕ�9 ۜ�4�-Ggc�Ϥ�BV����q�_$!���+Uԟt"�!�M�jQ.����%�#���!a�1]��qF5�6�z3��v`�k�:B��"po�6H��D�%��2.�δ�FOv�Z���Ү��a5�OD�)u�dJa�pg����A��ۻ�	~CWD�@�3V`]��i$�Q���mW^Bql�����cq>})��L�-bZ����m����\���30��&�,�H
S�[����Z��Z����a"��8�0��>K���,�9��I��"�6��_k��k`R�\6;k���_�RH����:U�c|PՅL|i�%�$Q	��3JC��E���ee�G���'�a���4 >�c ���]S����߲��������Ԣ;���CK�������G��>��PE�;�\b����}1��5�buJ;�̼��8�T3˞M��Nc淢Q��P[��BR��0�VJ�6U=v��{���;�U�sN
�����q�fR��@�����NU#�/p�ֶ4�I3�T�R3R��܏�90y�1l��"~_�B}�Y�ҍJu�>� ��������2Qz8��t�V<X����v�/�׿�e,�oe���������yM&�^�L�d�M�F�xc�s���ǐ��a�&~����?�aP}�m|�H��o��D���d��iLP�>2?Z��cvP�&z>�s×f�ȱ���j�1Y��)�4��J���8y�y)�'��09U��7@*�z�Ӿ��!��h���U-2��g_�g�᱓�|�ޚ��6�|r�q�vы6��v�,a���J9i�ĔΙ��+E��bzc���@�9(��E��e�̆�I�4��S|�_����,d-��s�4��)���7��6�w�X�o3r�xJ㛞��|ǌ�I�K��{�4p M Ou�8�1�飴����u��>������$�r�s���i^1���:���U���4�_S.�JҸĴ����Y'$x:<�%YDD��RP��C�LE�l��B�>�x����N�d�A�ؚbo�}���x&*P�����Ɠ~�4E�v;��0G�jV�Ad52�r�2	��0c����Ǌ�s����75�@.����}y2�h�@�6x�/�`��B���~����&��d�ai ��d���F��w�Q/]���i>ۀ��hFX��G��!`�ý->ӗLnx���b� ��C�`�8Ur��,��E���Vك�D�r� ���P��{�夻ޑ9��ޓ��BY�jͳD;��6�{C�v� G�D\���`�>!�g;�p`�ub�:�>��;�ۀ����?���,�,	��!�8��Tل Ф +tC���N��DTz6����Y��&S/D��
��#�ț&7&�V��}tqA��c���Kx���b9b<�=�;�s��2�����������+������7��������n
�����kRk�����:�m@s��g��2w�̂Xk,�lR1��X���4�.�C���k�8&������@�i@N�46�ݒIUadv�jT�>	Ŧ���[ R�)�l�=4΃��Wa]��h@�oTi2��|�C_b%���?�������d�fH�HR`
�~ro�$Y����N�{�@��&R��wTkzr�(�ɂ\P���Dk����f�sҡ�ƚ�q�?��lOY3�5��g\�}�ϗt��"%
�0.Ztx�8p2���m$Ŵ�DV�d����|�_��W������/�
:c�g�2֤n��nK�����E��%�Q���8�|0���Xǌwv6�x�00	^0��?g�|:�o���_�w�������˿��f%4[{����H:�kp~V7J�E�T��a�;a��t]�����������Xw7��v.%�Cx�g�G���D�a��˓��f�qi�>�c�'��c��_L���?D6~f��œ�������lS��ꙟ~�����?)�	��Ӏ�����d��!�5Ʈ؁N����{j=����L����%?�\w��RV$�������;Ğ��G ��)�^l� 
�جʕ"̏>!���s�8K�jb)�dS9�d#�'6|8�؎��`�,����G۔`�H��;3�O���v6ٸ� ���_��+�/<0�!t�GlQ�����~Q�Q_\xG��Iz0U��+�@Sv�=�D�运I�4r$�u:��|]Rt�d��Q�-��QWu ���z�=�m��U5Ei��k"�t�  Qw|1p�Y���NH�6�1�A�|�f\b&4��f;@
#y��Y5���y�,>�4� Ԭ�#�'�܉��l���!hOl���".��i6�G�;VU���H���B5h�9X-T5�c�7M�g�NyV+�k�8f_xM�B�ϼΎ-(�NO7�}I���0ie� %z�]6���I�@��8�;p�>����:/��_���;o1��͓�I��Z&�G���荥�F5$9ۙ��Dw5�AI�7�^{���vѢJ���6�&Ʊ���F�t�	��q�E�̏?~��b`K���[T�B�rG~��#V�"D�E��?�Ov@��+Qh8[��~�`"��fL�8�<�mV��T�`z;�h�x���T����ķ/jy@����r�q8ɑkƼn4��,V�yO=�us�ЊI	-(�-q	�UG7�9���.~4k�m�KbάS�v���"y��������es5���ޯ޽Z���'��HP��C:oa�%����u�׌��xSMy HY�F���6��M�H�3�%E�˃:���,Z]��d�9��$-��ӡ�<�F��0��t��j���*@��`����p�\�Rs��E���c�J��$���k0��{5OC�+*���2�L��A�����q��Y�|�b�����H̡Lq�,|-�`����9��a��;T�/���Z��/�#���� Rb�Hb��*%ܚ{��X�+@
%+��-H�;��x� �s�!��G�j)��)�����b$>�'9N�rT��M\V�E3aƈA˝�@Ҹ��:�Im@�n.�Fħ������.F���>�]�r�c���l�
}*]]rR��R :�;cGd/��^69� �Pdb(�C�^Z\`kQ���^bՍ�33;=�.����:M�w��%��gb�o����S�Md�l��ID!'�F��`�:{ c�"��p��l���A���ӳJ>����1�/"�Ѿ�I����xP�)b�)lE3��&��DU�aO[b�Ѣ����X�W�s
5M�󢙖l�8�=�)��4���X��zW,��уC�C�F�G�ݯ�2��
�{���I�ݵ���%H^:N�[��%�m��0Pk�ٞ1�ɲ`���w%](��Ү	�Ķ�?���	H�DS���^_n��i�#xF��5�� :���:ݜt`�H-anWjv��i����礉�h0?'_q	�&��O8�l ���|v�]N6�юBP��,�KR���I�N6��OWV�6Mi�Ae�P�	��=�l��s��T��޴��e��,��dfQE'�]a���qԲ���g�A��fa
$�a��~�P�O0���*���ō�Y�lN�Å���q�]�I��)x�t�>�`$�(n<��؎�8�	�뵣�������%���##���V�L�v�p0�}L|�Wo���G��Ǩ}�>�A�8T�)�8��/Zj����KU9J�x<&�fZD_}^p��njJxP��;5�'񝎕�VGě�:���Y�p}Qi���F�!8]`V7'a�f�[<�mgKE� @��&z�"��8���i�K�/�I/����?��z` i�@�T�VY ������*�hDF�zF\�:�0��p�M����/��FM��"�r3Q�C�= RZ��Z�7��&Ou2#}�.���}�4�E���}��.MZxM�6�f�� �}��U�<N�hd'����󠍃Y'���h@-�Ɔ�$�Q=���B����98��vPi ����P�EwP�m�0eL":����b�����ߋ>�2v����� �2~�|G������i�0`�Ht'8z3�lV�d��v�������>�g1�
36Iu��ީ`'A�{�1��,<�n�v�����m>�T��Jz�x��Ŭ�-�~.-���0-�P| �3Fc��и9��Ɠa��;����5� `�H��w��I7?�=�{β��>����c�K����`dAEj��n��T�����G��g&Jl�o�;oܹ�Ã�����K�5�g���EQ96����P�Z<;%v��p�޽#ϓ�ӓ=�7e֣��������W�k�s�c�{�Pi��l a)0VtO�`��ͭ�"Аѳg���8-��0��yhJ���x|D$����h!Gٍ�U.�;4�6��ܔ��!VgD�`�]jw��頣�����b�<�S��a�07���߶���I�x4w)M� ���X %���16%��A��0!�"Z�RЮ���;�0Ə�+��ݫ��� ��VB��ł��q�b������.�n���,�A
N!.^��9���;r�x�V�ް���{m�	�z�xt�P����2���A�)�Y�񁹀�kp}�`�e�i�g�*��G3yz�A�,=�����_�x���*WQ�M��{�s�K��E7�5�8���G�ͤ�a��t�S]5tܐ�I�I*���O���4��e��,������2���������.ҳ@�ZX<�3��S��:;Ȟu����j/���-?N;��ٛ�O �y�01�Dݎoo�}��3����,&b_�6�T
`�.>�K/����b����CmL�������7���?2zۼX\w��K)��qs0�z���n�����>]��Ϸ�p�9�c�C�Q� `U �:�
q=r�8R���&iy���f��˓�ؾ37[�xs M���Y�P���yۡN X��ac$J\���Y�Kp�D�mi~B��5�~D4s�� x]�m���3��Q��`���V����+洺_�^�A��1���$��ōߧ/�Wk�ȓ�v�&a K���*$��~a#��SA<Jv�k�F��@�w�6�0d1��A'� @s�l%(����_1�R�����،�榢��1xEę��.��4+\�	T1��,�����m�60!�~K@O#d�$�175v��E���Z���W��BM�ک�g��9h+�pe@
qv2���}���X9� J����m����\q)nV�fR�@����ޥ�|��w��codT�`%�h��D����|�86E	�#�BkǗb��.Ʒ������E�â�`Tb�#����s*�`�c��z���d�h1�Ɣ�L���	A8���Ul��^P;�/_�Q@�z��ȃY�\��$����,��!��
�z:����0��G�tF���>X�_�N��WY�m'�YRQcӊ7n�x�� �	�J�{���#]u�'�gT0߄��7�z�]���jw-3�&c�c0E�w ��U���->����1�g�A&�%��R�����#�g q	���oR�F��JF�HL�s�4v�X �6485,-./����	{/2J�	C�筒7���K�F)`�# �Q����y��(���Gm0L3g\�J-|�@st~��K�T_��
+��w���:NХ��c[ո�x�.7T1���<a�Օ�?��@�xP�T7һ}AR�����U�j����epOA�I��SO�x�,]ش�sK�/�K�L��|9ɤ�'��i�r�dM�~�n1�x�Hu�1 �F�|H�"e���n|(�4�(Vuou<6�b��bv�.CW�!a�d�M��MQ��)�M�͞),@�O�s�d�J�D|�L��I,��b *y��x��#˜��� 	fzL�R��}n�p�]�?�% ��bFJ%R�R�@:���
���A/�7ڀn_z�dg��g��Ydb�����h�;U;���ݬfA;�NS
�FY��~���/~�?��+���GZ��実��P�oi��@:���U�\���>�\�wI߉��Y�M(�m�)S��	#�;��Ǔ�$�g���D?��O&�}YI!���T��O����%fך9�!�.F(�B����Y�j�[�l�hN�Ic��J�c�w����)������-���=�:��'w' e�k@Sټl[�?���&h���ӞKm��zCq\p���1<c�}Ľ��~�J�{^:ލ��q�c��p���4�9��R�n1cά�#��P<�
�=��8ݬ,b�L��'�)��,|�s��_kI�4�󄟫���Y�O��U���f�O��u��%���C�p��MA_�m\��7��F-�{0K��-�k�X;�{�b�+i�t@Z�M<y�Ѭ#5"0�>��l�����M�\'飙]���JB����a��j��-�5dV��x~TFꢽ� ;P�T֙��6���K$]�6�T����5[(��"&ZŸ�5�~�����Yu�Q�쏏��{̉Gc�����|�r��8����=[�b�Q�j��w�����؁7�&�vԏ�YpƎ"�� ��<�� ��I�|��z�&���c0�i2#�,����p7/�ğ�`;C_6�`�gF*aѳ��pE���_@�����2�� _x���6	����IM mm�!+l 47r�-iL�X���:E{�9lP�l@��vf�.�6���9� Rv�P_�������N2�e3H�Z�Q<]���|�h��n�\s3�!0v0�l^_#�� ���1�K����m��r�����t��e=tQ�+y�נxiik3	��qE��Ů�t��~[?04�'1`����RQDs��¸z�o�P��)�E�A�;�)����n5��	���[�z��(��Dݥ�8X%Jt{��\5`�,�ߕSN�fp�]����,pu�0�q�*
\�ħ�a 5�ɨN��KtW]�Xۅj!l8��c|��P��Q;�S�2+r��&�btӒ4�=�F���oǞt�$��*�h��Z��fx66&i�h��Λ\B/0Ҿ��u��~���j1l��x�q���c@f[.���OyG��p�G�5?�6���%u��v�����:�(�8��I��̶�l�$e߮�)�9� ����`d`��?�M��?�_O��ȶ��>UDxi4�c4���<~j�����-3z��]L���sН���}n�g@��|����8K[b�۾\���zk����\���'�$�iy���F�;7��8j�SG��fZ����([ؚB�I�D-3���:�?�3�����~ڷ4n��|^scs�~�e�<�')s� �a�>³m��%@��v1������?��5ƣ� �;�6�Шv�<G`y�B��u�O����#�σ4J�����	PM䆈>U/���	�˨�	}�٢zȽ��#m�3�rq�)H>�Jl�Ew�C,��飃hX�OdnD?wSl������6a�Q���{��< �t	 G�>*��8~���׀�gI[ly�V!
���D�v��:>��l=#8�8G��{6�v8��\j�y�nF&J���>Z�M#+���0'��,���a3����e�O�v��O�B�6?;;�\�J��mH�~	DGc#��HGj�X�S��6�Jn��?�����z��
�T9����JC��C�C�]�4Jβ�sm�21��i`���ڄʎ������|�U�-���:wo�]��m�> �ȅhA�Q-�q����댯��Ɓ�/ ��wp� ��rI���#�����;b�}�Fuv�p1�����d�b�,�`��j�������g,L$�3��<������"_���J3�΁��AYx�u����9���^=c4�9��Ճ�W,��um���+`;b������ƿo�GW���st�oQ9G&8e6ډ���fC��Lm�����[e��uw�ͯ�(� hj1 �>���8`�q���<a8r�<�E;�o:���Z_qb:(�`��XyL�ܔ�8 �ʢ�2.�e��cp��!#�]���������[���^�7��V]�@K� f_n���f��e\�&k?5�<��,E�:�Ц(�F���rB����la���mV��\
*�Y{�~��9�=���u���Aԁ�sj�y���_�~��8v�9�}i�\&h>o����t �wW����<zǋ�Z�
]��qu����&Z\����G4�L`��7ճ��Y�C�Թ��E6n�S��29��G�L�g��[�lj��Jٷ~4p�pY���[6��MX�`�I�͒�n*���t��Z�.�M>7_�Y��)�VL�w�o�|o���;���M�r�Pl`��U!{g��/��&[far$o<a���:��n�� Ew�zYL��Zb1^�n�Fе��׎,�>7�M���C�ɀY���mp�*�9�����t'�M�jac)����@j��B�r�a^��{�ͦ���{��R�{eڞ�Zw��ڤ�\�^�EGd8콺�z�`~d�G�!��I�� �7��D��u����aB��قwDS+��0�C���=���H��%&�EK߼����E��:+��ƨw��%��#�z�#V&�R�F��<A���R�9�E|��@�؊۞zTz�u�{�-.}�4�5i���i� ������޿2�����?���>/��-%��[�D�$>|���x�� K�p�9�@4~�^�X�� ��~��=/1R��	P��ԘW���n��,V��ڱ�&W�e�4	�د��e'�Os��7�3�����B�� �Xw�`}��5�ՉP 
��&m>F�62п+�Cx���Y1�4���]ǅ`$*G���td=hG��*���f7^L�i�.���h�~׋ξ8h��Ş�aE)6?�kǎ�	@:�4�~�*+-�j��O�<W:0�ة��f�طE/��yv	Qn����c�ʌ���.vL�<ҭ�&��Pq�U�V�PeȮl��)r�]����:�m�������+��G_t�T�a�����K � �O=�0d��x��f�� @Sd��u�3S�9v</�qNxD�w�}89�Z,�՘���C�c���h1�e�fX����������c��Gq!b��m��<)���p��*�4��# ��x}�����$&Lы+��B8�4�
>?�G���q=gz�Y�a�g��+H�Vi��c�xr��^�Ϳ��u�7�=�>��H�JŁ؋j�M6��`%�;	"}��{��f@��M�=� 1�dKWA@	�3��������Rp�kB�[%��s�	2r�Qⳝ?_z6��7c^����v"Fs(�Ntט}DP���5��WQQ0��4L�֢��=O8 uy���(��2�̀�K(�wd��Ζ
C�<��;��#�����zJz6�����C�3�������{����T�h����TO%.��&�F�z�^%�Z7_xf�D����.�h~��K��o�|3������>��q��zv�0�0�{��`Z"C�i�-���F�>Yܥ����+��Ƀ�f�R��d[SH�%�GfJǼ�<3KH�Z�d��ß�WJ�z��w���q����Dk�;�Y�]����'{�l¸��߻���9=�JT�)�'2�N�+����#��O��,UMw|�,7�{��J�{zjY��0j���Z�=Yb�Z��܃чa��$���a�XI�P7��Lc�G@����ٛ��1�����=�^+��k�R��Ō�J�:�X)�P� �'����H@�Ӹ��'O���8���D�1aF!�Ii���D;�kb֠#��ti;�-I՛�UI*QA) d��B"�Ӑ�Vٍ�{��w��zz��u��@�TYp���|���l�{<��X_3X���V��߫���X�]7i�S��΀�Pnwţ����2��M�A�P�����5��{����j<�]I���f��F:n4��Z��g\1S�G�mAk:1}{P���%�r�'$Lц[��� �@���v�~iY&��0)�@����.�U/!|�>/Ɠ�DQ��3Ҹ����V�O7(1 &Gd�3-	�-1��{�u>ivH�t"���F�R��8�J�ܳ��q��גkt�c����i�>U�+a�K�+v�k��%�u���ˁU�rca�@o �z\�O���4�J��}��]-��:N6����ź���"��9�6Aه�	�� �c(y#�Лv��Ƅ����4k�i�s�]ڵ'�^fU��F�����,��A[1Vj��B�Ǖׁ��X���K����v�����Ez���d-�W>\���sK'��4��D=ᖯ��5�x�Tt�7�u�tI<��NbG���@��4�}�vO�y�Vg����f���w�ڷYڮc;#un���}j�X��t�ˮ�l��[��ݳg�ɍu��
q��@m4k=18.�\���hZ�3��?B?������G�GXD�8�:#�X�w����^�؊�x:!��,6��1�K���Z-�[̴�cvYҸ�����������i�<^�׈ۭ���6 �����QL2�WP��%���]�@�a�
s�'��c�3�=C �#91�⟔��:Ê��1"%?�<�n�,ј4��z�e5��~��R�ž�~e`K@܁p��Zߤ�lu=���
u�Ł�A� � ��'j�:�
�a8І���z,��"ѯcvj�;Ϣ�`�1�l��ll�(��w�^�8j���=��C2Cb��Ʃ�=�~�c���zO@
���ryL�Qױ�Ī�%ɓT�S�d�U�����n�x��e�[Ǿjמ�Q����.�xk��(�0v�Ζ��E$�.�tv}�'�c�׵��&J?�$���Ym�Ā����LE'*�}P5���L�bv�b"����-~
��q{�;� ����{��ؾ�^w������$���;�U�5�46i�,�8�����r����Gwǡw�M}�s<~  �Ծ����N\��?��-m���e�n��i����`fRa!�*`�3�$�* ��w|�R�踿]��ڬ�ݖ��xi�u�z�k�KJ�`�I/��]�"���¯��cA.�k�@P�Ϧ;�a���1n$��AT��z��/�čc��& ������6��?�	l�$�����ՁI�8��dկ��8S ���t�X���k��Q�/��ՏetO�W^�
~�\��R� r��p�;�����M�Sd%
r�?��N⥃@ѻ�ٔ�t�:@�j���)9���$�w*�����w��GZ�)]t�y���!1��ë9f��J	���i��֋G��(���F0��/ǵ�Ղ�t���6��E@
���
u,��D���nG���2I= �zH֚��`G��W�滭�A�����G�X���-���+������&�a9Xb0�=5q���s��ݐ&�ף�D��$J]G�@f���Q �jD�$��Z�����KA-h��ͬ�荙����=7�9�"aS��(��̀ H����w��{Q`����<����y�^_�$��5����<�wJ}��T~�����籗��A���D����@ʛ���H�Dן��~W�S���H�\�y�����z�����Lf�O/�k:�X�pr������\Dq�F�M�� U��� c��GRE8���@���&F�
M��h�7��x#�L�ņ�
L���<�~19!�d��.� ީ�����E�L@��^�d���c�Z�8���z��I�d�#��X8B-��YGRJ�D=,<���X�b���z����fOe�Q�ՍVC¹j`2}� �"q����[�:���GuE\��~�>@����EşW wI�t]^��w��L B*�y��Ӂ��Yy�n@���̋@�\��l_w[�1�sSQ��V�|cA'��E6�қ��j^R�Fi>�|5̺6fY!77&j��A�93N����{�\*MǬw�k�� ��%�k�'W��m�ړ�i��A�=�O
�&*�F�y���q����9�l	/�K����$�y�Ǐ�[J#��%1恋��5�:Mc ��	"��{P�%P��f��8�4�;"�SL?�+w6����#�žb��|�s�U���D�����`:YlQ���gi$�޸�۴��1�B��H�U`�ԯ�l�+���Jg���;L"�-�0$�1�[��X�L����b�M��z��&���[��ӳ�T9��&P��r\���z@���V_�{�"8�@��'�qDǺXc��e��&��H����War�@��� !8�v��=�dI���J��θ덉n̠Ӌλ�&�_g�k��n���!�C���ȕe�Y�����u�n�-y|q;�l��B;�{�U��I�##!@s����m "sd0��@��� ��wg�Kki�d�j��=ð2<'3͉��-ň�4����� g:���6�To����9���� ���w]b�׋�y��J���4b֋�?Iu�?��q.�nG|Y�-&��ᦟ8���T��� ]2#��DE��Å�1�
�$����Ã2Le#�s1�9<^ǲ-J�j�U�x�PxS��?�:%�E�f�\R6W�y"�.�1��!�v�Y�l~�Pl��r1.��Z����Z۱�g�N�h�L��̝�.���'�-W���ا���%u>(q1�V��R���z.�_ �f�O%"[X��h���=0�"a�4#]`؜><���c�3�k̮���q(�ބ�e��9��Iw�)��o���yw���6�y&�N�q؃`d�>���3�,��`M$M�����溢$;җ�+.��a��\���j��P�,VF�e�r��b��]��� D��+����})MN2z�@�L�&�(�3��qw���5Ճ� ��l�L>�-�\LV�fj;>-KbS�H�)�|�$Q(2�Rkc��}n�fD4r E[���_�瘞���Q*��+�e[�<�P=�L�@T+�+��:�D9�ˮY[b<q0�����T�P��4]"j�[mA�(a�]�O���6-���9l�A[v�W�i%K}ܺM�#�Y��e�HS�ϓ� �Ya�6��Z<冲}�]=k�.�Z�y��{�N���zk�	猖����_��Q�����@�AȄ�� ��, �[��f����3#%�R)��d� Z#�@4l��!U�A�QM��"�I��+��O����i�ACT*Z�Y_�#�:IY����I��	��C�ω�,Et��;-��Er�].�' ,>9�~�`oL�)�X��Ƭ���a��<Yu��P��E�n�����X��u_��O`�e�p��P�q6	f���o�!QcM9�b�Lm�Z�#%HJ��O\� ��,1�/��,��������3�-6��o	�`5���/X'MX	QD�^�u���D )�#�}
�al��l���%Ϣ��O�cٓho@�hb=�*�.������\��V��CHR�D�k��� ҶI4w�w�$RM����ig[k���XN�ٮ2'g�)�Ӳ��^����C#ӫ9\c�Ne�Ff�cq�ꢀ�M�&}�j��PƋ[1��vI��N�\�,�ҕY7���tSU��X�hX��)���D�����%�K�>R��AU�TQ/	=E3��7@}�����4^��|�[��b���#���R�=oLUＨW� ~<&��ę���C�D]�xR�tڝ��}Y��e`�����y��hC-d�� 1O�n9�����íD�� F[�I\\&U#�r`.�zSm_��U+.L�"�F�ܬo���ͱp�İ0$S�%L�D)t�5��`�S�X���cR�DMn���!IB�~��lRDS1:����^�����hX�T�p�?�	��}���$u��!)غ�[�Y�i�� :Ƈ��Gg�� 13�V2H�N�$�[��{� �����������:Lk�%6�����b ��W̱�iE��B�� �����b6�����PxH1��yt�x��v13���Qi�@�:/��Q�hZ�n�J-L�I]úF S�����/G�E�A�3��I�5\["�-@��y֗�-�D����$n6���	��eu���Ԣ1xf��z�UkW<X|6[dL�V)��ժo&�-�d�U��-v���F�8s�%�=��F��G��*�%���*�k�:0�ثfۍ�2(.�G�D|X0���[1[k:�k3Ь��o�[�=.����54o�s_
�Az�QY�6W� ��gS�����wi�$oDD�.v0?ސ:�����+|d����a�j�{�� ��8�}r�E�4��^/j�L"��%���/�'�us�k0c[����g���7d�ۊ�c�� �n���߾��u��Պ�f�Ƌ�YpR)lV0���G��X� ]M�����1�礛r�7��MXg�����<��l�����tL�~dӽC�	�`���S�q!jz_V�2[lԄ�(ڇi�7���']�b��^Y��]{��m����e������!����r�������h�5 �HZ|�;���6f�����]�&���T�V~ڝ����Y#=ZyY�]�\�nq�,#�I)L���Z&�EAG����{\J�Ȅ��x)iPz&��1e� 5L��@�Ƞ�46�_����\���dS;E��8�4�e�\Nr��J"0�����t ���URq����:Fvz���Wm}��:�Nn�ld�G�T�,.t�^ց^��e�ը?�S]�	W���2.�+�ƀ+J��i�������x~Cɾ���� �]+7�Y��*&�[]�Ǵ�����y۽���>��llPE(I���E�O� ;���c9��me��u����{#�2�A��\�0�*@�mg������ы��`���Nt6����������|d`���Ed��>���'����M�>W�zrd��ű�b`�6�V��'2u������?XT��W�M,Z79҄ �>�QW��ޞE��>���`���T/�Q�������zz1 7�H�:��g�VYad����ԏ �43��N���ʀ�:AxF���(����4ϦUK��U��{�Ć\ש�Oc$���<��1�od
s�RM5�&ߏ6�����f�@��Ԇ �o��A#��@*���q��|���1� �EK
��-�y ���(��; S(Nc�SmkvK�n�����Q�/�l|'�����ėnW+��im6.��4���`1Z�ƛ���A�c|R��T'�<�dc)l����n��iq��:�@X���P	�z\�՘��@��<����]j� ���x��7��6ߕbv�[`Z��4n����� �������B�v4XE3��U����/
����˛ �ag@V�Ӏ�UW�����u�Ii�4c)����  �:#�v؉*�>`��� sR�;���rf;�<2�H�Oq?�St�g��/�l�yE�u�Ha'�]�ە��@8�A�+����T�6"Ոm��t�� @��B�ӹ/w4f5B?_�1/D`��Ls���ؙ�$���%�cs��ݣ�8%��uc���7K�	y<_�9�b���S���Uey^@{}9�ߵ�ї�Qo,�k��H����:vyK�+�����;�� #���&������.1ŨK�p�Y&���h���ĺ'�𬖐wLT�o�b��V�,�U��T�1/����B��9`:n&
�"}+a7ٙJf��ibjʔh#��o� �	��j�� >&V��쎬M�:B��nf�AT&8;�t@:�xA������6Q]j�w��"+���f��= Zy�ٟ�E6�̘~¸FJ����!���"��<KEI��(lg6��e��s#Oʑ(�/�ž��
�®r�Ko��Q�˥^�^w�c��fyU`�Xn�o9N�n2�Ae"����81bg�q�)�>e�@���0U���j�}A4&$f�TS�a�)Q��2أN�X®�PO�]�5�X��P%��e`(X �b���V�uf�b����|�LX�KƆ��nu5.�8H}�o(er�R��#�Ob��X�:���TR��I��u��@h����m۸7Ɵ��5M�M��a�
��7L2�Y��q�S
j2k̂$��ɫ�O$�la��'�.H�@���N�dq���{����*���Z�%��:�s���� J�w)�k�����9XI�h��?��,����?��(�BdW&�rT�P�r`�A �>�����d�Ǧ6���c�4`	�=qd;U�������� 5�,l<�ۢ_6f�hx�M `�>���|��vF���:�za2��c�X̠�50����2�%�����\㇊�Ip�R�t%co��Ԋ��(�`�+-� ��5^�j�ƇHҐ;v`�1�U =���(R��u�y"��S�,��?���3�ϋ}���������ؽ A\��_���k�\�
��ʭL5�����@ �nN����d�T"�؆��ŀ�v�K ����j��*D@et�R����'?�_�7nb�ڊ:h���"���pl`^�:烲���H���ǉm�6���!p6
{ƽ&-l�F��2+U��vuKd�`�	#��kc*3�n��(W��J�Kmb&şL�N5`��
�K��}3� ��x��vaV��AC1�h}L+b�2�U���?��0t��&��w�@z0 �t���M���S�o*�c��+���e�A$oۃ+�f�`��S�	�M���a �F�N��H1�lb5	P]<�;�;N��TU̫�6���,�ؓw0
gw��>&�'�O��M��&����!���3�ƌ�:#Z�И�k�9�j�r���#����� ��<�A6�p�b���-���Y�5��/� 3)��'��<�b{I�6��b�'툷6Y];J��e�8��D�L� x؍g�O5�otD7!Q:���&��iB恽Z��Bd0�T���X�����p��e��\�o��=�>k�^
�Evn���~�i'�5�+N ɂs"��l`���&N�Ln�C��a����KFk �EA�Z���sR-2IO�+ƾ[��վ����@|��p�D0ƄO}�l��q�giy	}+���4Gq
����)�+x氐�f��7�L��+T��=k��V�k��՚z��e��"{�u�̲��H�U�8��L��b26��,E/Z�V[�J�����ԑ-0NЩ.���Ǵ�c�%3B��'�fl����03�5Vߔ�,,�_ї�ɼ�\8�S�l�g��藍e��ĈV{��1���S.`��F
�oԸ�	���)����ph]��jjR��dr��6r�2~կ�� ج�NMM�Ǩ�k/>ѐ�'郓虡th��Y����IT"�X�诀�/���К�?M��6\+?j�#���t 9U�]����t2���
�з�}b?B��ؖY_�8~�e��q��X���c'�Sx�� ���b�?�+z�a��N�-/�0&�{���et����0�}��L5�T|۾�%N�x���;̓%�����0i�S�Q��5�
(u;Ϩ�I�l��#�+�D�]��᢭!�X��~�X�|���Iеgd@ ]�',�<�m�c�� ��l�W�"��i��Vq0qp.�7�?�6D���z��@���@�%��+�F�"i�>m?�G�_,�����-[H��KLxE ���Z�z��-�[��7%����1O����P�`lIa�Lv���N-ww��,�R����ׯ�ą��W[���ͯUl��"��D�R�z�+�bA�U3Q7R9\q�����}�L�����<|�\����f��HW���x\>�7�{���l���C�� |����J	&,KhG0\�o������ٕ��]]d�DSK' ��#z�?q4�q����8�}�
ڴ��-�}����T�@�����#��@�4�0����{���C{� ���^PD�*����YE� SW[#�0* }�Ol��X�����+���%I ��^kT���c_����o�=h�t�ۀ������g���0w�v:\a��%��k}�������,�j��>�����c���3w�<O���1�P_}&��$�̫���&b�1��I<� P�h�x�C����tA&H`B�sLA����YU��HP`Z��?/"�;����N��5V�� 5�ݭ�z���7K�4����Q�yށ}d��N��S�d���G�Q,:vXd�y�C��Tb��G]�+�j��><׼���]�د�K�E���<��B���]�b�#���l�6A�4" oQ����Z�e����b
��d�kx�4XpL�7�eyk�t�p�P�=�+>�@���vn���f:���fP���ÖQ�<^d��մ#�$���WRl�����)D{����� �N�m� �c�;�7��6y�LFś�~.`���e�wtA�!P�?c~(L�D�;��3]�)�Tk���qn���^E�k��zn������:+Ee�s��|X�f� ���\�@�XT&3iS)NU`�H�J�H5��=�>�F	�撴�V~	��\^�/)Ww�m�^x��Mt��^�(&2V�e�tc��`7�)<(Z������������O���w��w���NK)i Krٙ���Np��뒮�SC��%@Z'oӵN��1j8�L�PJ�ګAl�Bװ�������9���q�Q��b��%�R�^�@�n�T䋦�fſ�N�[��Q�C���8��G������
^�>�);���z�0I�w�IF���<��H�X��bt�S�_}��I�J�f�E�ʡ��|`�|�Y6ը�Ѽi�6��Dc6Q�]|G;��ｱ�"�5���S]���`�z������U��:�Jla����u�8�`,����0#}|(�������Ǐ��Ǐ�ݻ�I�e�����������K��c1�������+�aw�e*�:�N�
p�w��Y��ű �r�x�I�V`�~�8^��o%V��t<�R"��!b�G�Hծ�WaK�Lo��u6�T̳��#�aU��b�<���h�;뱂�X�}m�\`�Ffi�	��~o�
V@Ҥ�e,��YNl
��#WŝzyAO:2}ZaF�!��8Oc��^����~D�������W�P�^PFL�V���7G�h1��Y,y|x(���˗/Ogf�^^gf�ylt�,����O�/�RtM;b�"��z쇴���`�
��<1�Q�h�k�.�'w���'��(�[
�1vއ+��w�5�:�(�Bġ=��i�k`¡��1�L`���Ġ����N���FuҧWs���.s��գC�FO1���� #���r�:˱Ks@B?3`�&U��͋n��1��ԶK5]���:��Z�,/2���)����3�bX�$�����	�T,B������G����):��L��ȞŃ���Y{80�i ܟ���i.O����O˗ϟίϞ�ޔ��]<?
�X�,��'Ì҆{2��^����Ϲ�����X�1 jJz�I�8�DxԸ��˦��L�.Պ?���_��^�Yw�[nۦ����5np��s`N�g��g#��pa2���>#op�+(�4�LWq����S��@9���p=[?�^Dc ,R��u��6�%����Z�l�Â3M4�F�H������� ���F�`�e�
�-�$��N�>ߟ����~}W���{��ޝ����G֓�K0���~��P$I�0�|y�R��d))�W��כ�󺲏+|/�o���{�V"�����h��8���,�mɥb|5)�/��?�{<�<=}.��3f������fD�w���R2�-=�	�{������<aխ��I�`��f�Sm���(����	ȑޡ'Gc�kѵ��#�lb�ˑ��eA8G@Y'��*7R޴��tV@�/��������]��xJu^�O����h�0J�Ԇ��U��2�F$��O��X8�`7�R��#�UG�<��N����yޗ����u�O�EtQћDq��Uo kzS��s�������Z�?��p~��|�����/?���3�~�V/�Q��Њ1fi5�VVa̼���o��Q��������K��o��,�k�Ȫ���Y"�F�b���&����(b�r�O,��i�I�X��)��3�O�M٤��,�Va�[�E��h�.��/v���-I�n�@�������̐S��g��S���߼�X�z���&5nЛF�Sm���ꗻ4��=,��h8N[z��[c�@Pk�Zg��q1k`c��u���j��f�H���Kðͼ��N{�K�Ekf�:>H%����s��Z�:#o��={}o�ڀ�Pbx~=0����Qz����N�Tv��|��
 �ޑ�+$�j��<�\h~��j|��k:ˈ�[���ec�]J�\^��{���o�� S�e��w�Ow�1	��)J���:����|����.���S��"�ܰ���N�� ;�u�.Fg�p)����v	�TL��v+�l�٣{q�j�|�x�iK
Њ9]-�V]q��L�A1��6 ʾ�׏�t����5�P8���|�M��A��Z#�@kw�k�n��ʶ��l��`-)[h�}!�$����|�Usvc��Z����#% ���}9�+%&J/��>6~�9B^bi��ؑ�r���Xl��~h�������l�I�<c�]a�:Rp�x��� �u�V���Δ̡ļ��@���L�x� �������,w
������Z�����~k[/�݋ķI1���
�:3Z����HV�������|�IC���	�����N����w��T���Z'�t�:#��$���'	\��K��Teӎ��8]Ms��?w!^,L���ј�TY����g�d&����H�g})��~��'��f�ة~Y^[n�Pz{��u"�Ӈ�0��ꀯ�.΋sR$t����=' ���Z#�"|�E[ د�# �x��k�6��{)��k�0#k��1�G���V�&����x��u׀���F=�n#�됨��V��B��g)=
6�!c�9�(��Fm��ȬPu�v�c��CH �uw��DJ������3�|�� �މh��	,[��&n������oqߦ|���\u]��}�7�P�B�E�I*�k8����l���RR��_�<��3r��2�B+\���GߍV�[����-�A^V[Sd�B��1C@�Y;-e��J��6Ľz�X�EQ�J���K�i�[UȥF>ېv��ԙ=��iz�ݘ�z뮻3�]
�s�7��N���C\:����3x�;��;O�H2�g�H��O��MS� �T"��#L�ޢ|�����Xh�K�� �*Q �>��|>2���� �"6�<g���~sV;�@�g�#��E�%ߡ�*e�X�ԼH_W;��?c�|��n�&{�v��o}�pG{5�1�zQQ3���R%��^� �[VD�0稟�o�wN,rw���{��#g�{�L�4��K6��<��bT�������1�����R�����,�53��A�v#[s���u�5�ì 9'Pt��3��4�]�C �E:�G��V������w�'��/w^���o����/T���˟�߷c����;���}c�^����©�34�3Q~�,T����<��T=��0�ċ/�a�ɞ7 ^�-��O�{<�KKl�?c��i���7��q���� 4~@�o�m�2�f`�� �[��-0uf}2P�	�n�'>���K�����������Z6�c�<������T��U~�v�V|��?�{�����֗�At�3K"<1�;}'%'���,�+y�4��j��1����#�n��T���M�����	���Yd�K��a��3R���4�޳��n��16͠��1��x���{D����l�l�վ��=ՠ)\���=�}[䄅�$\��.��k�������H8�N4~{N (^ Q}�wO˹t{���1��XLZ۲�.V6J�& �=Տ箚�ӡ�q�o�b�@��z�a+m�	w�;�xg���d��d��V��#����H�#'0���F����H{��K�������v�\���u�� ��A�#�@��WL���'j�d��\_���(��u"�@U�J<у��O���\����~z{f�?o�v�|3)�w鴿r���� �3���﻿�Ʊo��62hs	�_�=�*��墊�jn�<~�K"�k7��5{���F�=,���^�ȼ�`�A�Z{8����&_O��A��"D�:��l�����u�K��u�z����/��y�����>�Tx"��S���h!M٫j��� �ob;^�[K��������M��q� ��j??w��wT�Ћԕ��3�H��||�z^�W]�o�	\���ֹ[�M��=HJ�z�Ku�ާ=���}�����+�{%`(������:������F�>L[ɠ�״#C�YO���t���9&RHF G7��z�	Yn�i������EZֺ{�K�z�x���^\d2��(o�#�I�������*����3"�g`����,Ë����Q�)c���x�q��^b��:���G�O�;C���D��'���e�u�{ĝ펯�}�����땍��� ��D��L]�i�_���@sq�]�Z�n{|������|o5z3@}��U���������o�p5��7A!�d}j�\�7��n�6CJ�g��x��bq�5p0�k�߻�rvy���;g�%��5F���"����rS�D��o�!�k"�"e ����o~ΘU�]"1��=�\��1�AB�T]�/��$�u�XVe�}���ۄb\��u{��}�gQ*_��rc҇W �,]��ۖ8���+5 B3��'��JT���ZK�����B/ׁ����
��ˠX��=�o��}��^�V��@Ò]��Y�1d���ϫ�
�� ��g�H�I�C����8� h ����='��ߚ_��s��,�Jo��u�TzpM?��A�ʛ��<<������Zf�ߦ	up�]� �����AͿ䚦9�_G'�駺ү޸!�^˝�ҳG*����.�eN�����'q,�.�{f	�g�<�Rz��ۗ�E`�s�͞�F��R�6v�T/q�o]��"_���B�\���ϼ'��uz�:g���w����c���۸P�EY�l|��`4n���6	��������iF}�gp���fX_���2j�q=]�hAڈ�N�f�a]�K�w/·
����}����W�0�m����Ok��{����W��c�ϗ:+�JI߁h\���ێ �����~����p�����D�M����z\�m� �r�+k=P��&q� ��@�ǟ�Hl׳�_f�9�m����X���IW,7��zU��t�[�_��O�T�	���O�p�j_�\Z�V�Ǥ��=}���ce �<� r/�0�sV �1�S� �{���2������ė�P�$�&Ӫ�~�o�|Q�(k@o������r=��r\'�����`�kF�ϱ��
[�' ��ͨ��/���Q�f�Ժ���V��W*6�q߃���������!T:Nw�mF�z�� ��ҭI���\,}燿�֛���ј	�uF׺��c����=z�A�ZUl���>��|�&ܲ#	�zl�s�3�?sz����F�^���沺�Yʛڑ�W��i���h��a�D[�~�I�NI���[�= ��u�{��=���5@��O�֒/��>���4Ɇk��R�Y}��ڼ.���Ձ��reQ26�֮�~��MKR��K,4g0�`�\�n���F�a��M)�㵀���b�z��&�%]��ѹ�(��nD#���D�c��o�绦'��]���r��Q�~���r�,�>D���y�b���a��s���mW4�c`Y�S��8\3D̉m"я�����w��,�{��@Q����`�-7� ��g�w�:]�k���(~T�D����G �U����ts���{�z���A��-&A~��Kf�u%~�Qu�;�() �����z[㠻1���}r��15�s���y_b�#]�7�7*��X��~"���1����)~�i+끴������%&�븆�&[
`�тF����q}����͆�����:G�%���~�ZL�1�(��l��ؾ�WcQ�(4�Z%�t��CJn���>����%����F��1@Z�j$�c�[4c�r�m�}$��Rz=��ރ�t�E�@o����&V̷�ib)�Z�DCtY��c_���6� \W5��y4n�.l�wP�c����7���55K�#�R-6���V�k�s4����6 E��@j�����ط�K��Z�2�`�uBB��^��y�v?���R��b/�m�h'�]e�%��w�5V~~�
H��z�^�.��{�]�ޗ�u&�������}��6��ۺ�������Wm!��|����s*������o,#M�'��M��p� �W�8�J)����N"�%�-��u�թg�=H^S�X�ݿ\&X�@�/���ҳ_k��A���n;�����.U+�9j��%]�
���$���ܷ�* ��k��7�r�0�y>��\�<��ّ����"��8�4y�ёX�2��k�t�[����І[��t���փ���.�hz���n-ݲ���2�����]��Z}0�os�	@M��u��Kt���/��k��O7��6����"�����2���;h+Q�5�e�`�n)�c�΋okp���V�[@t��8!	�/r��~�U�Ri|Ǜ'�K����)�a�]��7n���@�I��zᘗ ׭j�-"r���@���ko�t�6y_x�׀ӵN�N׮���^[^�[z�j�ƃ���\��}3Ϧ�����'2�[ڧgz(/j�v���z����A�&���x}Em��    IEND�B`�PK
     #{dZ��� �� /   images/7b19d218-2217-455d-9a43-b73a208c2c5c.png�PNG

   IHDR   d  �   9s8�  0�iCCPICC Profile  x��||eE���6�ѫt�q�"�����ٰD�ݐd�b	!��l#[`a�.  m�"M�(E�HS�. � MP����ܙ;�w�������w��L;s���;�%ɾc�,�3��$s�-�<��Ǟ{UWz%���K6Jt���-]]	~���{,i��G�i����g����a~���a����_:`���'�}�s��Dc���!z��G��xrzS����
:�jKf����d�:�Ë&ɪ]�i�=<�2���м����3�Θ�$�A"ɬ9���>�Ɯ;����I2��E�ó�dm����}F�5k���6)�L\R��~��.Ӻ���nU�2֜�ff����[��78<4�M�$%Ӵ)KӁsY���L�M�M=Mف����n�ٻG�e�'+�iIW��d��-��N�˒f�J���֎�5��׭�Y�`2���P2�l�4�]�3�M�^�����gI�Ԯ�� T'~{\ˁs1�Y�ѶE{oR,���g�����u����C�f/��@����jM$=	�Bos��;}l���-!����b�$I�`�!������d��c��$k��$��@�y�S��������������)�9�%ɵ�m�ɓɫ��6l� vmاaY���6<��ڨ5Fe���:d�e��]����G_<��1��sژ'�n6v��+��s�wĸV�x�y+�v�MV^��C�LX�;�<Va�+�:c�?�ֹ�]���~�z����rͳ�Zk��������:����i�m����w����~a�/\�aۆ�耍����M��ț�n6c�7p�c��_L�x[�_j����O8cˁ���국��f�/o�����iv��k�}�/��u�|~�8X�Q{���Nݮ�ӷ��C;���_;�岉��>:�;�<y�]���~���t����ԍ�Zw[�}i����O���5{��k�7���ߞ�w��o���)3���f>��}���y��_����^�xs�p���]v�w�:����>��#78���s���vܣ'�w⸓.8����O;��	g����g�t�%�u���Oν���]���W^~�{������|r�S�����r�W�ܺ�����o��󮻮����N|��<<���?^���lz��g|n�秼8��^���]_�ፉo���x�����^�тO��_�?����ڕ\�|���pݨG6��3p�{�ye�A��w�J3W����*7W�^���[��5�Ys�Z�}�:����z^��>�p��&l��&{l�x�S7���W_nL���MZ���լ��ns���������=���7�x�XY���כ�-l�v[5�~�vޱ{����������^8麶;w~l�K������n�!;w�2w�q]��vo�+�+O�j�.����=��/���7_�֊���޺�}��͘3�p���3����{�~WϹ}�C���O�W]�ɢ���/����Z���c>c�%߹��������#�Q����ѳ�Y|�����q?<��.��U'^{�/N����N�|�����?9��3�8�Գ~�c�>�C�=��_��?�`���h�O�^<��/�x�֗�}E�\��U�|�Օkֽv������冎w����C7/�ղ[�����κ��;����~s�o���߽|�w�{���������~�؃?t��w���G��g���������'>�������̎��n������^���F�<�o+�����������vx}�o.}��^����<��'�����>��Ã����n���c��_���a��Fm:�Q���Yc�{����ݱ҂��]����U�d��V;~���8u��ֺb�׹g���{q���0z��7�z�6�}��7;a�K�������Ҹ�Mh�r���n��6�|�'7����[�ro�x�{��-���JfU��v|u���A�زӔ�}�e��C[O���kv���Gwy���]+_���ީ�N���{^�6f���'�����W~����ӷ��{l�&�dm3�����x��C��{�~�Ϲ{�S�^_����٢�Ż/�}�A�����:��e���{�*�m~8;���ݏ����>�S�=���w��p�9�铞;��S^:��察���>��3�;���>�чgp��~x�G���@�%}���.��%���ν��+��򰫎��q??��3����+���w\�����M�����o�ආ�+w����~��o�;w�]�]�w��Y�ιo���>0�����!��c9�ѓ�x�c�?������'yj��s����������em|~�ƾ����x�ٗ��ݯ������?.{���/~�7�x�ތ��ݿ��ƿV|�����m>��x�'�$:�%�5Lj8���Q{��{�}��1?��7��m��+����U6Z����V�r��V?s���<�K׾v��ֽ�����+�_�x�&6]��M�?S�ŭw����O8g��zh뗷�x����m�X��+��˲�ٙ�"q��Uݣ5�ؿm���cvXw�	;�u�̘����I���z�?M~�}��7��t�޹tʏ����\��	���L?b���͞��⛛|K~{J߬��?}�+n����3�����7�>�o�9��m��������?|���.^��%���_?(9x�e㿣���C�]r�I�_r��G>~�kG7�ޱ�/�k9��=~0p�ܓ�|�)�N���CO;�G�~�ǜy�Y��踳O<�sO?����~r��_x�E����G.��e?���+����ّ??���9�ڳ���/.���n��������7��WO��̭�����o���?�͊;G�n�]��W�g�{W�o�}�����������w<rˣ7���]���O\���<���O�磟9�/�?{�s�����x�{/��i/���K_���;���?����o���Vo���޷�}��w��w�n|������~壷>��'� rX8��< �8!I&�+�jŊ��N��]e��X��I�J�s�I�����I2�KI"�a��g�ly0�j9.͹�g�G��1����Ã���צ�L?h�C'�Y<���Z�ޕv�8IF`��'�utT=`M�?���iI2p�{�14��V��@���u�5x� ��������������v`�dc����ߍW��U!pS�0�0{��_�+p|zT/^'����gԅx����xm��7z{�~o�~��ܿ�~��W�zF?�W�3&w�ok��9�v2�@���z�3��i/VJ������hq�>�[�P�Bp�OH%8�����/���� \�������p�e
Ҝ.p�j���|��n]	��Š�o��?If�����W[2%iǘ���|�|�En����&��[S�p,D�2�:�L8�=Ȁ�Au��z�c8���!O��e���7�} �s�;�5-�:��g��?�?�2�\�M#V���+i��A��"N��tm�Aw���$%30����@f$#:W������S�7i�D�� ����?�!� s?�4�@;��J�8�-��SX����e��|�I|�?o:��1� $�)sd���2���K���gA�qs������l��g��A�s�"��m��j�R��������;����2<k�9���9C��/�?���?<kpQu`v���м����������ۧ���:ch�������޶I�ƞ�E����Uf���N��$sՁFL=�����������8�����e��JO���m}��;�zzۺ�'��vv�M�n۳h� ��:z��;�v�u�uU�'O�n���tOn��k����=��mJo�q���E�ա�:	K�ӿ�kx~S�u���Ý���7���|]}�{v�aܝ��zv�6N����Ll�i�k�~��J�(�[OW[kowKGޭcZ'�6;���Z'u�j�5�eƤUkk�k��j��Z��e��2ejwgKG�^m��z���ٗ�i�q϶�����ImS�:�����abwKo��)}]S{z�'v�y���6�TİgGGD��=ugz�Si^Rm�v�����܊ί��D�ڊ�\48�z�Т�A"���k�fk��?oF5?��Ξ*�e5�Xm��a�����)�J�L����=���Y���H�A�;ZZw��!?:��)=nW~3��sw7d�������.�8�����3��z �jc3���s���]F0u������Ӷ۴6K�qjWo{'���	c���S�4�T�2eZ�Ķ�>ld����I=U�E<����og:��JOKgW�S
��n��d���I������������#��i��fZ����A?�c��V�2���'[�F�
+a�ҽ�U�jt�W���^U�ƅIU�����~�������8���R-2�YiҊ�����~�f��k�q����O�����2��~�	f��ʚf�[�O0�
Q1Qz��8(���8:���'%�JM��=����&2�9�Ei)h�V)�T���c�e�k<�R��<2Z�Hוl�����AGͳ*�]��(4�M%�2����*�)�s]iMs�Y4�q����u�r+5�`�Iiy5n�E�م�Y-�)�@g�٪�%�#�%�_������Ό��Ԡ<F�J�J��X�05e��T�B�)����U%�%�1rנ�*Nf$3T/�i%C8ľS�v�Y��̬#�J�F�-6bY�܎>K�MX�6�1�HJ�H�U��&�2l�p�4[��M-5�$*���NA�� �Ժ#��e�F���ƪ�fRn����I�2G.�R�H��
<P�C�G%�Lf��5!�$��j�x�י��5��56��@���0�)l�8�z�k��~��R�Sk+p
��Q�:��Ƥ�ր�{� ��)�T�[��^G0��$��e�TY�#f��p0ZV��dXOp�T�9��@H7�R)�F+s�u���I)@�����r�
$�tMH:�z��mKx��ž�K@�p�D�G�%���ʩ�%]C��T�
ǲ�Gs�Q6+SN�����~*���L���p�8w�9iwRA#�5f��	%�AX���K�uRKK�uk3if=�Fa���K��*\U��y��#2���"�'����&�q4�xMl�i���'~D�T���@+G�$ͬ'������ ���B�%�ZU8|,ܣ%ͬ'�/����;�m��>�"���N���a�dA�t����,U�YUX�ι�:�^��#��0�	`��FA�֕�0�j�:~(+L	��CU�q	Q��u�Dq,����p���?CGQ�h������?�>�����=PH�?C�_�?�*L���ʩE��;�:��*J���+58��Iޖ��	�LC�d/n6�FC��� \��_1�?�$U��N)"�(�4����@���#&��I]�)U�6�2�)p
P{سդ�������z��� ��
�C����{*qR�JM1�T�� �42�U�hB�TJ*t��b5,���h;0�\��Z�F���*p�Z�!�:�t�jx		,��a�`�FT`)��| �#$9bFhf���Q�ë�R��%ͬ'$ia9Eq˒$�TFp\W��a�_G�,Q��$�#�Ru怈�HS5�@)���76�R�Zҹ 2�,�R:J����4��pE���$"��(���p�_G���r��>��P����j�PX��zB�n�w��0#�8y���(�؎$�'�0��C
cB�"�R�iA3R�z�0	�o� $CZ�f̠�p�v�u�!p}�5�#݃[� �Z(|���	x�a�����G��j ,*J�d1����%!�B,a9�8�]E钬!Be��'&���2� h�LI�gD`E��Q����.8 9�([����
�Ԡ�O"e*O%� ��d:EG��e:PFX�i�s�a
���X!�F$�.}0�P�9e,��c}G�U!(kd�FƁ�C&������ܭ�#�i��)�%�j���QĎ��8 ��A�=9X�/ WS���wD<Eg9X�?	��=�ȭ�;

� ,���{���P �K��x�@*�@� Dq��<+֋l�>Y�R�g�C���	r�W �b���A`��SN���D૘+��()���@�vd)*�������� ��)���BN<YuT�Рd�Ry��Dq�jd8��)2��(J9��*3*�0#I�p�BW�,�(���)�T�j2�3G�tQ ��W��(�G,U��bV!����?C �A"�/�-wE�k�b��d�qF p�d�>0� 5����%�*V(��F�RR�wK�;�O��g� "wnX4�T��R��1+���[0��+#sQ��+p���W�@(�"ׁsd��Y�G&+��x�(@ #C^N³!X��
�W��3"��yXE�3tP��U��)����������TE���U%�R)�g�	�����
�е��=�T ,�ܣL��(��q��5 aԹGC�F���pl�{,:
�r�F�s:P�I�-�J������Pmi8a8��Sa���f%=�bIU��gR���TH�>����mZ�6��"���'��DO^�[���"�g�[����� ��(q�Q�3
v�%��(��:��eU�b`���� 	E>��C��YVG.z"�d 䒪3���u�3����w�(���Ѯ~(]-����YVK.zr��T�#+�����jmy�񫥴�CH)ὔs͚`z%+-'�@��`(�%���%�	;��e��ؓ���M�@�=m��=Y�(4�� �1�p�䝡�����KL$J�����մ(u^2@��)�T���2r`K���fN�3.d;��\�I:~$=��@�{�~��*�5z��t�S�V��9�jڧ.q�q���s��"�	U6��eSY���}�eS��)�f�)0�iKzFϔR�I �`��J�+S���@ rZ6�D�ŠU~8��L#��� -���/!o�ی��-[Pi�ϴq��2�Ig��D\���j�yY��y ���%=#A���i��Ǩ"CePڧ,�q�������T3��%
�SOU�5�& ����kAu*�Жt���U���dÆd��	dwH�H��Z=�Z�QIy*�Q0�&+���%^3���q�yBR��w*qpNz�KӘ��`S���K2��Pt��A�����OQ�_S�q�z�(iNV�M�$&H	��1
WlDO	� ��L�Qqr�Ty
��H���cJ��D�7��(�J�¸K�0�0�
=Ed�?'���4��\������`t�L%(9�qZ˭��P�3���� �!����U�'�g��g��=�}�f�P���L�H�EO[�f�����J�r���0�(sy�@���Y�t<�aj�9EV�

M��)���r=YfiNF�G�A�c��KI���I����U�HV��q�Tw�u�J'WyOn4��(K�cOzPĀ%H��H�)a��\�,���B֨W��j��J
o���Y���+�g�łzl��i�S�`���p�����e��}Ҝ��g�'��	�h
���.
�V�;r�p�6��fȊ���,3��	�
���~��C����2+�QT��/zR%�S>'Ҹ~H�����V ��* ����J	�J^�o�O���(��;�×t�R��ۢ'E�T@[2*S�(�I�"�0���#f�̸���P>MZ=DOU�3n�����:=Z�甔��2?�Isfy��V���<�8z�{R�R����K�?�ׄ��ZP}Or 1:F��q�TR��cq����A*0��W�e`��SGeR5��%�z䚹�^=�.iĞP�Y�F��SN�9�O�}~ڛ }̃7K]D�H}��J���(!��P�	 ń�"]D"l�dIt��Đg�(Rq�Q\d�V�ʒ�BfX[
���1����)\�t�����vȅQ.H�o�,�Ӕ��� ���'J�����)[�
MȨX.�#(�ڼgF�L�9�x��=�|�t=��BBz�������&�bR���a��F��q��PyM
�i��!�	I��F����pʤ���<O=	�iQr�q�����N(���)�)���Y&�
27�dqѮB7?���%C���
۳����ڭ�O�[��Mb�rÕMVm�n�y��Ӽ��c�y�u�yfF�~�mD�Ȫ��]:���EP� ���!������&z�Dw�4E�j�������.�=�o���Cs��1���s�.l�6��3�r�VYrIR�\�����$��uH����!��-�G:^�g\DR���ݓWJ:^M7��+i�Ƚ礥��@�x���8�Z�*����ע��b6�K��缔���$2c�tňx��G{�UѩOZ�	��2�-����Ll�HCT�=�����jEh1:��N�|T��2�EhE`t��������9�@��9^ZB��rFO�s[�/�uG��J@�@��Μ��;��?1��N=���%u��RbǫSzt�Zm�]x+��At����n��A� �����,�W�7;���D�I��'qX��E��}+��n
�:W#�V�zU~��x��|H�HԎ�~rAѵM/�@��٬���Đo�n�1�I�9?��x^�$�Z�6�df�r��B�疛�k�I�
z��0������9�L�d<�D��Gb�\�	"o58='��|7�e���,#_$] �����ߦ�3"�d�9��7$��V�$�~�5Г%��*52�Y�u�6�p����,_B� ���U�nЄn��x�Q䭈�~��":Jߍ*z9�SIתa�<�$��|~!��f�i�Pf<)����s��]�kuY�$N%t�����Bb�0y�I-�9�)�r^�?^�V���Ҧ*��X.3�^��`��ZA�����r�_�s��z�Z��yu~������a�s]�ru��_A�xA7a�v�㕩7H�D~�#'�)4]��ym�g��iH�Ck��Y�n2o��o��S(RɜW��H|84�TOB�r��(Z�V#�
$g~�ty]z^�_�r��MV� 	�)��&�F�DM�9'�nN�y�5�\!�N�<
��<	��K* 3HV&��|Λ�f�ji	��6���r�Z%z�@ʠ%�J���7����I
���`o�\+�_�� �K����V1(�w��/�$�c��"ZAx�J2+F��+ϋ�٠.ጵ��S9�k=/9k�j�)�u� (�t�d^��N&2?B�+���
}��a��;F:Mu���v�c�tN�:��PQ&���E� �˱��@������q/�\x���>P+saϓ�z�D��܏�è�U3��PH��IN�]�[\�g��=L��K�)q��0�g�,�"��|	�X�j��_I����\�X�\+�i�z�5{O 2�^�"��­	�2V��~��� �e�_:�˯��7�y�,d�ݵ��D��e�C���r�*@�6tC����C9�*0DAfE�������'����ޠ�{2]|��I�HH��
�L���{��/�� p Y�ܤ�j�N!�d�y��t��n2��0L���u [ɘ�![|΂yO����������0Z"���D��x��0�W��đ����0p�և[�ڛ4'o�<bfl���OhE��yC�@��Z�'��1�GC�8
��{.FW��-0�7�HN�7��Uy_�#��Ⱦ�C:������EuӬ yȬ8��a8D�'��&�V�}��d�0}7�9��1�#	���p~ǰ�=o�a�՟0���1CF��/���{�2{�~܈ahZ�Ρ�2�Z��1��7&�T|���6�WO��er�Y<���_ʲ0��>BrJB��"��xx���ӄ���[`(��a
S!i���+)��H�׳�a���%G���$6ă�D�)Y�D��8A�q#��p�ޭ�L�ԑ���[`��F�{؁��WD�i$�QyI�g�y��g>nR&�]7�����Na96+��n=o�0X:��v�]<� 恷�0Xm�r��y3�yC��T�%|�IY�1t�� �t�6�,b��=�a��>��F�\[�#$��I��ﱧ�BR�UP���h���-0��2��T��c1��[r�S�1kU1�i��R��I���1}އ$��U�5���ɽS �¹�"�z#����,���eIoC"b����Z:pR���E#$���J��] x�*"��y=�T������[`,'�E�	gA7e3�[`,�ER#汧�F�'D �O�;�֟E�0��4��U����ED�� w�n\i)�-0]m�NL�B��)��F��X��_*��AF#�_xCY�&z��-0�>�f�e����GɈa����̼��TH��AF��2���T�j_ޗȈa$2'�}���|��g2b$����&�t����0HWT*�$���1��a\��x�g�"#������0U���x��H�UэPYNbX��2b�n�R�Rg���0�"������K
�y�)�O�%9J����YDC�\�NC7�9D#	q�@j���F��
�xT��XЇ�a��yX$\E8!����1"w�- m�:�ce1��Oɛ@Zx�9��FRu1LL���I�fàՆq�����~܈a�¸D���G����d�0hաbZ�:ݤ�k��R�nP�2�𵷋�a0��A Ï(�㐊FR���`��i�3�[`��S���5ؼJ�x����JB��`��U�0��/sOʀ�1�J��-0ZC�H���С�i=o�a��m`���%�>��������-�'��W�u(�[`�����w�i�k
*bŘ�ABk��MK_�P�(�Wo�
*�}*=��511}ZW�����*b�L�+�����n��T�0���+}���	0��uZ1�E�U�;���>`�y�(�{�!z݁��>�Q�(�[�ިXx����1���?�ʐK��k�y�`AA� |�Qt���Y�0��3�a�*t=bEwȳ� |ȧ:��Q�F�9}(�=F�1�k}~���xo�ȭx�F�3�!X��Ǫ�a�e!��A�@�P�V� �����҆ڕ��ޗ�A�p��V|mEG�+}D媠}p+��a���ح�礦˙��FY�@א��R��ۦ���D�=�?71��k�{���)�C�atV$m��R+��:b
�,�&�&���ǩ:bڭwx��T���WG�黩�s�9i����a�d�^B^�C�<>��h�SAPT��"���k�x���`��l��?�À�{��X�Ky݉F#��O�#���5D�"|2K�T 9=�p��`
�Y<��O�Hn�`
��%@g��@執�a0��nE+���Iz^��FCS���B�J��a�
5��M~M��sވa0E𓚤Zu�Y:bLa}�Hw��,��5DC_�ࡄ�¹�}~�#�q�گ�(N����y7T3<���lz�c"���)'?�:���8d"�A�

Co�2C�R¸�Ak�{����5�bW�G��5T$	�E]��-�뺉�Z�Ã��89o�a���!�׀��͛�a�5���-OZ���Z=ޡ'����%��1�� a�n����/��a{5�C��X@Z_G4��W���W0o"���~oàU�:�!�/H�k�&bËg�=4T������pև(�:i"�!��^ʇ�� �L�0`Pa�z� ^7à5�>�X�¸:�L�0��Z�;��ri��Ɛ����4�<7À�P�pB*?,�[`����-��GHz��kL&b��3���6X<��g&b�{Á��C��x�D�PP!'�q5�k�&b0dv�CӰc��#�1�e� ��]<\��+11��Z!���b#o�a� ���z�J2��[`C�)�Y��z��o�0�M�c f�&�k��+ۈa,}Q^�fC}�����1P�!��.Z��f=o�a�V�<�����]�����{Ɲ3�!7����E1��a�p��`0�c�����Bɹ��l�0"!B
̛��/����0����o����(��2�����xa	��q��_o�0��*�W�����<o�a,U�Āj^�ع�b#���)��R�y%���җn�7@��Oڈa0��
2@*��5R1��uK��wA��<o�a�G%����K�d��-b�3��ᰃ�4�x�-0����n:⃔<&���%�;pt�͇qrPao�XCߐ�I�t֕�r��Xz�x���[��Iϲ��w�Z,]��֥��Rw�$�_�Q���d   	pHYs  %  %IR$�   �eXIfII*     (           >       F   i�    N       %     %      �    R  �    ~  ��    x       ASCII   Screenshot�lK  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:exif="http://ns.adobe.com/exif/1.0/">
         <exif:PixelYDimension>1662</exif:PixelYDimension>
         <exif:PixelXDimension>338</exif:PixelXDimension>
         <exif:UserComment>Screenshot</exif:UserComment>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
���%  ��IDATx�t�wsd�y�y�gH��+��Ֆݤ�5ÝU�P����kc���~�Մ���H턺�M�a����*
ޤϼ���yϹ@��l�@e޼����S����+
���P*�B�Z���~�F��W�e�7�y���A(����{��9����g���O��W�X̟���o��~���>�ߧ�^i?��5�S��B�\	�lƙ�%d�o6�g��nh�l?�)�Z��1��;�O)�K�VSSS�d4��תzϟ]�z�>�Կ�ݞ��h�3�U�Vt���is ��MOO�iS�F�f7⚴� n��� ��y9�p](��}����}�<!�ߧ�S@��$���{���g�~e#�$�
�7 �0.��H�,�
�������~�`3==z�������~��+������R�:�F��n���b���C�!���/���������011!��e�r���I�I �/0�����R4�q�H��S$C|��I?	� �� �kN?�n��a����䟉C lŸ�V��C��Y6��X1`7�(�L�&''�1�͚N{������VWW�~�ޥ���5��+�r�t:��>�����밷�J��������)�E���O�[B�	Ћo|�u�D- 7�H	xIL����_TB/5�6��u�^�V71��tO�r
�)���d�9���~��E���咉Y�nǈuR�?<<�s�./���NDv&��B���?����WXYY̝МX��T� ���o�����mX_ꍉ�{�)�N��,�Ά��#-�an�ۡ�j@P��diE3
���=�W��"�������u:m�=a��j��ʟ����gÈ���#�FNC ���j-�f���Pww����01Y�Ŝ�qb����P0j�2 p�߱��0$�H��)[/ϫ�R�+:�����0�����f�ik���?�1\�r5�������&�`���q\� ����ógk�Љ0k�<cn��c������B��Yϔd��k�F=��Q2��UJ\����QR�6@� F�L���]1��!���Y#����O��wR"grr*,//��㣰�jSԉ�  	�����ܬ��3��a~~^����ֵsssZ�ٳg��Wv��p X��:��⚙[�v�����OLN������%{o�^��3�������i��8(9Q q�X�~�
�� �`�K�+aqqQTztd�l�=�1 i~vND���?ί��77eI�9�`@r���0ʘ���כ�,�k�	 �~m�� ��� З�����W�k�%��`����S[�Rx��w� <Ar?� Y���W��UX{�,|�����\������Ξ]5.�gm}�Ν[[���Ja��>��}+R�U��>:�$�j�8��Xgݮ�+�bq�5�Z-��5�ɥ7�h����,�P�h�����t���-!�ڨj!+&
�X����]����e�ՍZV@=�i��6����ٙ���m��SS�09?a�Z�1D0(����`��0$��f�Z-k�z��Q�+Q��o�fC?++g� �}6��jќ�p�bx�b]߁8X���C�g2�1B���e��ph�8bтtK
s���"�ܬ�D�C�"8�u�)�)�@�:��Dٌ�鴻:_g�ͩɦ )��{X,20�t�ʕЙ��A/_�4��� P�RG�j�ڂ��07LO7��W._�s�!#[ό���߻'N��_�ҷ/��e��@��@�Hy��D�Q�3��%��M�A��lƲdO�$����K����@뜰�1QeE���A�:��b��:�����G����¢�uh��m��)�3rH�N�6P���h��"�c<y�D�2�ƀ�	0�˻�����A�о��vwvEm��R�[�ˍ�F��[3q�L�mr��7��3�+1b�C�Ǧ�^oJ1vQCq�H�����a�D"��GY�9��M����2{S�s�("�gH1 *������ϟ��7V\6�5�+u��ã�8*9��a_�Al����C7!]�OfL2�6��$�rg6wj�Ȃ�QPX	���Š��h_��W�dY�6��Xל[]�&����E�>�{e�?�7����^�a�(JL���-]�rL@Ƥ�z�Ϣ%M����ɓ���o�#�C�j�b׈��7r-�n��S&��-,�cqQ���gl�:�b���P�錾E�a���Ǿ�D<a�E 3����~s�U�HD4j�.���E�h��b�0��c^3���c76��Lb>�'���x��^���KN���M����ٰo� �����p�r��2 @be<c��#����� ��!�5��{��ލ��#}�XA�E�,'b�bn�P����f�l�1eg<wg�C`D�d��j��dW�BxDw:]�^|�����ƾ����.�9��"I��8��(��R�i��UbMڗa1��E�L�C�\�����}���h ��(��-8���|�p��w �=!?�b�`l��ŋ���Ʉ����1����_H!��$&�PD�DKt��P����r�x
ݬ�?����qʚVWW%����{��T Q �{���80��̭Ȋ2�ʞy`�#��H��~i���G#ʰI�r�*�O�l���MmЧ�3Ƃ!k��sm���3�g��`߃��������08;3z�q(�cf Ϝ0�xl���jz��ޮ �?!��e q)AkkϤO�Pj�G}��w���� pNj�K�.�	�������YKY!{�H@���5t�!��� J��`�ez`b���`��/A"V���q�GI&2:���.�ƒ�p	�� brS�d3�(�y �OX�iJ�e
�������ϝ%q����lCnV.��I�;4��,LΠq�r�<t���Q,�g���eYNl���=C�ŋ�Ddw�����gr_8�G��Qs� ���/��3�_�M(��!���(�Ơ":����n����s�$���'��)���x�k����p�K����{* �������w���h!����s�9Q$�B$�1�L�υ)�tɼ)K6��ƽ�Y +����y��C�� ,./���1ſ��J���1q�%l�b/x.z����B$pHh�H�8�q���Dt�,�D�"Q�T��{���B�z�߉!"�L/�O,�Z�,�@��.y�?ZZ��*a	�ƴ�<��ttӁ�� �,$�������_w�i ET���&�/L�`�/��(Ul�ݚ��Zqy
U�]8E�nH���[�1�`���H����(Ii��M�㔮w"z�2x�������x��������I�H����0	 �v���H2��Q����\0Q��)�(�s
)�hp���&�� �3uD,��ˤPA��������r��u��{z����}���ׯ�� �r��S��a�`SljwoO��XGW��]4�����l���d_�<���ϠT7�l��L,�o�N����t�3Q��YB�m�����\ r�&�TAӐ�.��س���MU�ݴ���D� e ɻT����!�zt���b����Ƒ�]�b�|]�|A��������u�`(�n�t�6�����(����e |���)�eCʖ�ݿ��_�����bc#� �#�|��~O�êa[1y6�x���ل: vJ�7V���7�x×2qH�B/ ;�r�V�S��S��ו���X�>l�3A���W5�`�X��B��3%���I65�ӦW)�!0M��6ͺB���X��9x��[)�nO���gW��^
?��Q�X�n�;$ipCr(�8�=N�t岛��cPHx��<z�8�5~ ��$�*�ΐ�:�N�.�5O�<Ud�?�+N6cV�K�Ք�ȩJi����N���J�ŀ{,�T�G`��XX���!E������D�8%��5<��(��H�&�*7G_���2��{ ˈ�@�������;�H6����p��j�z����)d1g�Čm��O��e�t~�嗹8@�H�Oz����ښ8�?�P��K%z��@*I���eC����w�
8k�FM���	�_��ڂ�x�5��@ �p=y�+DI�xۈ��K<}��!`#�X+�4��-�6I��l����D�֑�!璲�[1%�A�Ŝ�HČ[�r��]���0k@^4j�׀��W�j �]]=gb�g��L�	��u,��s�w(��u�]������s
@b�o��:><R����T�]�8��hbṉ��m���Ŭ!{w7��XWL?�2R�E3n
� ��k�{ ��UWܕŸ�ҭ�,G��z�tL��5�Y5�Ƌ��I)i��zAN�1+g{�#pW�������$�5`@aq���B'�޾<Վ�)��Ƥ<�ho:e����O��ggf�u�m,��|E\� �]s�3�!d����=یQ�){�7�|�{  � �?�DA,�'�=�h2����%��#���BO��Ϟ]�ߵzU2ߨ�dԵkW÷�~k�~G:T{@�,�7
�q�L"�9y��.��?#�x/,M����v횸B�h��ȓp��'"�D��/(��ܒ�үU��Z,R���]�.Y����Ʊ|<����{f�C�����+�VM��^"�h�MJ�"�-S���p�ٳ��" ��Ec��/Dg�8EؿX1e�J�Ư�5���8��4�UP��@%J}��n�� ��I]��d#V��!Y6�67?k"�%��������Q`R�O�sh끈��1���^�0�-(j��޸�4-	�T���_O��ˀxy��P�Ke�M��cC��ޮ����f��@�x�$u<��Ő z��LT�����pw?RaP��!�Z��e���Y:���sCI�&�R7����@��e�2f2�DWa�% {}�e,��������JWd �D")0(X+�Y>�������X{���ck��� �1f���ʣ�f�cEL��ɋ<��گ�(���c�π�պ�f(ׅ�}U� �ub�����2

� 7Wb8RXY���3a�LU�ب���0<��6��#2;	A(\���Wo�sAf�YT+f^�}��P�ô�P�+׺LkއS ^�d��Yu��<�Z��Y1|eģ5JAx�Ϟ>�5�6L|c� �@ �f"����ѣ�yб������7��R!^�4��1ȅ�L��(%���P��c:�X�B��F��g{�,,��MG�c�� �T�K��"ڠ����?�x'�4 #U�4F�`ld� e�LW=~�<\0����+F"� z.2��p����k�E�#7���|���-"$� 0�B�R�2���
q:�o�\�����Q[�	D�	��p����!��0����N���!)�U�ߊY�dM�8�9d��Ҋg 톄7X��{���
`!RH��H�1^�����>�j�&i�7�k�������pG����3/󩅚Yep�Д����O�<����(#�4d!R=߰'�� a8�d���+�ޚ�2 ��@2/[:*���AĀ� �˗.�[�nI
�{�%��r<��>N�
"�(�sf���+Ix(�!��Mq! xt�6`x�m{g[����-�E�"2`�w�}W���=��5B,袉R�Ħ�l�y�jǳ~��OHRa2�R-��H��s_h���:�����#J�&J�HfOG �PD-Nݵ�W�����H��� ��z���e�bأ%"-��d�nˊ�rѪ�G�7"���R�0���F|��*̟rH!�����.������h�����X�X���� d`�ݸqS���������!F)$��6v,DVc�'���b3":]����Ѩ�b+���2�����^�m�^S΂��D,\���w� >6�w�}'��B5˧�22��
n��z�psRD�j�{�b������@@O�bs��'	P�R�!Q�S��.�X��R�h�����9�T�X�5$�q��}��1J�8�F�Ǩ���G2Ѡd�T�}��X�Q�= &&k��G��҄u1��P���}/s��Hr�o+�b�ā�j��8�F�(��b�E�$��.6��|��P�v�����ޫq ;y�	$𣠡qg�I���>��t�B���T��_�Q����X�������ǥ����ū�	��%3Y=�'>��]�R�����_� �@۹s���s�6o�T�/%eH�"J�ݿ+'%�#JWl��(D����vd��Km�X|`��j�����w�M�`T{<�ᡂ�k֍�c�T��\�{��h����zݣ�OMD^�v[�=�2e"�{�QE�7��:���y��I7��6{O�r�1�bVN��%�ć�t���1*Cda��(Q��1�#P7�q�LS�>n���<u6�|�Y�w�(�[
��X�[�u����,��=�>�=���S�(�k `tÉ�2���B�qN�)7q�rp�g�cA��TP�QĞ?�補�	�����ML�{+�W�R],T�%N�.r������S/�%eBOv�h8g�ɻy�fx�b]I|�(�#9%ĮG�<� DGt������t)?��'J|<��#�<Q�� ����zD ��Y)w��7���)w�F������ˉ-K�#�@�W6z?�!^��Ck/�ߐ�T����q�'�t��d�\ �_mz��@"\�r]�Wq1Ux�;R_�g�^��y�h�0H�-���w0�"���%Ʀ�-���;,��SF�ޑ)}Ҳ'���Q1���|���TI��rB�������� ���f����u�xp
?��Se�؄C��͉YY�hø�\�3�����EW{"��W�D8_om��񒥆����Yqׄփ����´��x���O��B�{�cx�S�X�`�'8m�K� ����v�PJj��E�.R(��/c�lQ�gg�z�@�A�b�����fdy�Q���q\�~����d!&���s ޻ﾧr~��ߛQA�c@�e�M�+D}��+��;���N�3��dBW�#ѓDxa��?_�|�Mx���M,�#T�Djq����� ��(���5Ǵ���Id��Hj��B����f�&馈����T3�D���3��8[����?w�lTjn�C9�CU�{>ً�r z\���#�G*P�-����tbRU�/_�
��V�������&|%�NGQ%�ٟ��#�<8�H0@e�V���.b
uC ��>x>��3�q%JG��olo��X�F�rl��dN�lI�g�I����	Q�*�]�ES\P,��`���J?D��P�
��x�I_�&o�>!Ԡt��LSj|ɿ��hK_�z.Y38B�C�������ڱ��.�
  �?7�w̪��?��v�Y#���ס9�O�?>�jt�fjo�X����r.����� vMm�SƄQAo�O�,����O�)��?�ڌ���W���i����H��/#JB�=W��6M�M*�5���֒:�����r1:K��%�SV�΢����~%R��$�}�o���V/t��p��=����wE�� �IG��B�^>k[���H��= �{]X=���T}��f�C����*�΄��n(�L����C����+.���Q��hP��!d� ���%"�U#�%C>ݦqcoߌ�I���q��s��l4�" ZLo��H���2?djrB�����U5���TT8��{Ks�p��m�	#ْ���M8傽�3�'��=�,PP�[険��w���r���I[��8 ���H�TE���#Q噅��2@�H�*�?���Z��pbꦊG���gR|A"}��;�U`��8�g�;Jm�ʭ�P�X��1�:|#"J��؈x�dA�ʿ僈!�r��b�I!�+F�w��� ��d*> �HE��۷r��T��*�r����\��萡�+Y��)@PӾ����x��X~���S"�gYA�yA��3y�y�@Fg���LZ����,Cn(���GO"烅V�޵Z���hi�;>'>�A�����z��I��T�ԿFH�tM�G9_�rM����J,n�➒L�8��/�J���ã	!����s����W�U���)"���ɘ�������r[[{.���������6+f*|��w��Ç�m������M���s������bu�B冐A�{+oa��B��	㪙��"���L�U!4C�[�-����aoǬ�U3��M�-I�:�AT*kV'�ًu��jF<��������eEIE���Μ��(vI�L4�S����&�$��H!�RqT��7 MNM��:&��k����g�^G����r *b�
���W��p�7�p�bf�����y�и휙��aŵ�弊^�����cؚq�@4ܥ�E=�9���g�h�x��wLy�ߢ����:����+�/U+�L���5�^�������"K�Fu�9 g�6@L�1!��\�!��,�;�߿��p[[[�L�`P��U@qP�-"��bY֏�v�#�$B٘�7nݔ���_��/!����#Y3�ؖ�%��
�Lfnl�D��;ъ����
@z����j.��~Ĺ}��i��&�fz�15-qI] �8��&8��SQ]��J�L�]�jI���Q�s���(J���k
�ye�RX{�L50�p�����)�c,�P,g��	�"T�@��%�+���+����f��wR�B���y�?ܹ#�q���\>S^'j���&"�h�����Ϗ�5E�!r�\C4$�����1��YT���!�b��>���#lˏ�a�0�ҙ,7���nGa���Ԕ��` Һ��H��S��'��|���z��5��N?ִ��˞:���ce�"
(�&s��>+A�Al/�#�<�b��(z�0*�\����٭���?|����2��7��*Y��pL��typڤ�jeh)J^j=:l�b��]ZxN��2q�}��z���o�����H2����x��CҼp����b���O��Չ� ������R�������I��I�r��Tyr�[
x�;xB��k����OA���b�O>�Ĩ��p��u��(P�Fg�D�ɗ\�b�v�P^�G~�N4�czF�G�j�M:	 *�H1_��4�,.�WR��<z���R�q�Ç���Ad�?�`̺�8jѡň����6<1�J�n[�ƍ�Ѿ$ �;����H�I�.@�"â�p=\B<o�,����Dc��'��X��@A �
ѥ���ѽ�B��L&,2���ԧ�������+	Z�/�R���hـw����( �䱟=}�����eq��/������'&g$ǹ'b�Pz�.Z�9NQkQ�E�<|�P��ԟK�.+�8E���A��˯����
AU�(����BS/��NʎHNI��A�P7�%kĶ"�J�?�I��[�J �pq��333!���mI�d
�	kC��� ~`w�'��Y&^�O]o&G6O�u�3:
 �!V0��M��#ߝ�J/x%�[Gp)�g %���eh��l'GB=��KsZ�@�"
y�˵���^�8z�6�ݱ�!���ǚ�s��qP;�x��q(�)I�!�����e};�44g�]�iґ��*�y����@�{�~^k�RWa�'e�K�JD�;t!�6Y����8������	.*��� 9�օ�����VN
�"�}�QQ9l�D�jiy^�QG@Y�\&:�/���96nE<��S��!�Ì9�ݖ���ޖ�C�M��J��I�F6�ĲW/�v_LU��a4�׃��MJdU���M�x����|-��
}�؎�y�DH�V�>SЛ='��(�K�/y�=�_�cE2Q���ߪ���䓏?�"�(�ʎ���A(�`��Ca@�tsFE���Z�{��8�MD�Sy���'^v�(~>l��Y���*�O�Z����ѡO������JŔg�&�9�p��+揠�[��2jF��"#1���g��(."��v2an�De�hp���2���ئS��8ZY�-:�'RX ��։�X�a�%�"r������TgE��ֆBț���z�-�6^��*LO3J2=[Gc`�Ox
�M��M*�*�^P柾�ڋ��fOj�AȅX�eD��ҀR=cb1����s�@���\ژTE��	�I��Yo(y�v"��3��.��|��ɔC������U��J����{&i��ΈMɑ���i^ӊ�B�� �а�+Z�X����~�3�>��h1T�B><�/��R KE)BMlB��o;;:n�H�6}q��E)O�$��E�G2��3c�װ!��Ԅ��G1y�M[�B!�-s_��p����5��n1��*���
8���* ��F�0H�b�c�$�I���F5{9>��$B
c9wӱ��ۦ�ѯ��W&��P�����J�P�=e*�=�{�*�9��)Ku!F\B)l ��-u�h.z��A����7d�C�=V�4���0������vh*��b��V�����0�1��o�'$�pf�4��խ�@t%�	iJ�f��f���V�9�N���3�s�\h��]��a�P%�/�z�/i�نX��(ℱG�Dl���U'E���KW�h��e����X��T�Q��]Y�,���/?R�Bg�Q��w�F�[����,�'�H�8���g�,}��>K��3K._��� �C�c�����0�޻']	@h4�厬��ޚN!�Z�j�8�m3���8����'C6��"��cxɞ����l�5&�94�'(��a"�X�y�J�(�Z-����+2#Sʕ�ǭ�7U
�l�+>��Sq���H���j�F����)q�][�1g�>�π���> �J�k�u��US��35%�����I�;��`�bQ����4J�,:��pp%ZTT!..-(��g`���l�����d�1'Ί�
�e�����K�F���?��Z�v����Ӏ�<�82s� >P�^e�pǮm�X!fBP��IsCP���s�Hi�D���Q�yy�l `�j�WRwE	?���L����xaVR���$b �!��
����}�ԇ2�pGj���X(*.��l֮����Q�s,�Z��p�!,7D��-������i�sR-�<��(W����*�jiK#X	�1��zd3�ǿ�7���B�tE�ñ#kH�L���Ϥ��uT����\�?ڱɾcA 淿�'��aq8	dAu<�I�CC׎$>��oK�cU��{q��ݝ~�)��n8����pfA�Z�����xޚF4�����MD�[	�}�Ǵ��:�M�Q�A�6����y�����O�Q���)F�B��{R��9ߞ)�#S�d��)��u�F%��=�{�u���[�5�F�� ��]�}��L?ͪ5��Gm��
IB~���W�\���3/�S�rET�C�X6}`��*��&� �h�?�P TH����s���� ����Uc�(�k=z$���4�!!N(�E��B�y�U��łە������]q?�E��"�����C����J��1�bx^�p �	j��lo(@|�cB����i�F�(K�y�&��q�QO�<��ȿ�Z�Qi�du�PP,}��+"�iL���Q��%�B���� QXV*Q�y���dA���/�I�e�_}���L5�wx ���j'9F�3�ڝG�P����1��7a0��f)#�'�B��ʅ�*�1�Ǳ��D)S�CU9s�ٻﾣ�A�^��~��˚!���/�["LB�͸��0��^��W��Z��X��U8yi�SzR�h��P&��}܁����#q4Ā��Nk����f¥�F�%t�X�P܇,K�PDq�q<�WV�b4�yp1kR��!��ycM��H\�,+S�
���3g���\�b��TKh����= �7�-���A>Hy�6~^�����1�k�9T�8�����' ����Y��hB�A��@,��Ԑɂ�L�g�F(j$��lM���pN[5�Q�io]ʝ�-�N�M�0"�w�;�@�d��i߈����K�0� 0���58��ѯ�`�p�H�vQ��z,�%x��B@l�Ƒ��Գ@������/�@/BK�jP�m1A�~���0���d⺷�z[���G*~�=�Bg<� �AD����\ȕ�`T���u!���R���o߾>��SQ(���i�4��z���=��+g�63r"#�ܚwo���{���3%�: 8�0��*��_��93K^}ЦF�}zC�e�<+(֏`�E��I�t����1Z�����ű���5�j�ƕ?.����U��(C2vs�q��(ޭ���8oP�LL$	x�i"�Xp�������ˍ)������S����,�&��JP�:?pg��aȜE��4gC�`=3/�C��^@����bD/�i�i�ٺ���� �k�n(�"��\�\�;zr�TFU��e�ʍ�����v1BlG���B��Vy�K��z(
�9���>z�O|��pc��>�ţ�U�a�g\oq/�mE�m���7�:5`�ؓ��0���ſU2�����N�eL��sG�3D�����6ۓ�T��h䳳��LWyթ�/�#��s@jr�j�>qʱ���E�В�`��R�tAȋ@hj���RG\Y)J&+�������r��Q�$o4�$���� R����DJ<�2��ը q�@��"�1�S��r�L�K�W�Q|��?�I��4U:�Ue�w~�14�G�=I�b�C (e�P����a���?|[<$�����|�b�k��>�k���Y���I���j�&��wzw��y�Sِ�7c$�G�z���.�p~5Z^�s������*�]>D�,����z��P_�/l23=+dj\�!jSs��xY�#��)���8�]� �\U��}zvvU�����3����b��s��hA#��3�\DS?�WK���&]+��<�	Y,*�i��e�a  J�AP6{ �a�%��P*[&���TOhfva6���1�O��4�u�^�)����q!�hT�1Wa����g������p�#"l#i@> �~�g��|d�j��J�Q��\���iq�w�NH�a>b�oۂ)����4c qQ�;��ߛ�p �H��y*�0ġSh�D$lL �`? `߸y���Uש1��B)�m�4��n�{~(A�S��J:ڢ��Ou�Yb��4;;��ý(V��e�*���A�D���{�נ0
�yr��x�x�
��3\.�Í�>���5��'_���d����w��T#R� bP�*���b�C��< ƍ7L�����h�`�|�����8�z�d2�  �Q��)���]'[bޖd�]{��y!��'�����嫗��Ֆ,$5��y�����a�`���Ռf7߹C"륒]�s �R$�u��Q�)���������<l����\�hn�����[�n��?�\�M�	P`wOx���SH�P �ԨQ @�ģ���NÛ��x�(a�=�6�����D�:�*.q����J;�~�0J5c(b͕��$o�����A��-?���<�y�ܓ�Ha^ӄ8C�`�!eɊ�Ќ:<9\��h��"�4v6��U�:�<���z��a���23Ow�ÇO���T���ޡQ�9[k/L��4����K2q��³�k����3
�=;~&ca1Nz����$v4��ņ�$�p�L�=�����N���-�V|iׅ�����/�_I�<��X�|f~Q�|��a.[r,ød�~V�`?�rfn!/��v��j4z��Κ"\gx?ʤ����C���R��GD�K�$ON�5X�`�P�"�yxpO���޶tWC������Q�"Q.�$	�r��=y�����~���ݻ�@X=>j��k�B��{��#Ǆ��8IgRqTC��GSS��~�v9z:0�By�<���- {��mQ>�W��!lv��`�"Y1$WT��b݇�5��jΆ��������sa�9gD���:�ɸ"�����t4�4hmjʇ�������``;0�a�P!x��\�=a��C"���1X� �B��o�Bsg{ꔶ���
eK�Gvɒ�� !�b����ƱTr_~�:�g0��7r	��~��X�.�t�e2y��7oi�o�\�Q4_�D!���[�ҵ���9#Y&A�7�v miq��0���X�@��ڔu�Ӳt�&��x�`O�EW�NL@]41��)CGz>��(�ux8��HB>R��ߥI��h���Q�<u妘V��6���"��F��%�VUD��~�d}�8eƳX���W��L�Q��Sؚ�At��������`�*3@[֢�ݞFq��+��u�/�E��ܗ��Ȅ�1c�-Y6:�������Xքc��	=#{!����#\�^JS�T%C����]M�M���[~@M�0�����;���V�%��7�L)�S99<���L���@�XR��;���Bɦ����|�A[��Q�\��9���Dhzgr�01k:^iG�=���x�Ǡ`�P�ѡ�� ��ǀx��w���T�����9d4f5ҸG��͏��{cS�;O(��+�`Y��V�4O����gC(X�.I�����Ayhɱ�bq䇎����x��^��1��o"�ϖ��Y�*>L>�1
�4U�"�;B� 24 ؔ5Vu����!Oȸw��Nh�k������]9O�uA� 0/��0��'up �"�Y٫��� �	{<7��C)dv'+.���Y/���4��c���vm?8�H�t0�����Xlǖ>��y�R���I)�Pd9�DN��3��rL�#V��r�>=�2�yr>�	c���"%5`&�0����#�Hڰ`"����ȡ��2��Y�:�̀퓪_���L��P����߹s���R�a���3��5�\���T37Q	F��K���:̧���='�h������9�_1�#�w{�n�0%E��^>�3���}/]��[��9?A��{��2(KQG�9���(�@�<~�T�C/bb&���[��AU)IW0��Y�@' L?��}�̄D�'�#��}���Ԩ/�ͫA��qp��#}����ȿ�T��|˴k�(N�rc"�1X
v��ɫN���c�'p�_�/Ao����G��a�H7����2��8�J9?��Q�	;i��B���·���_�E�2B�H iZ���6����o���A�5�ׯ��vO�_��FT$g��L�p �I,Ϧ���!L��A�O�
W�>N��pxO�Z/o��P�� �F�ii�qx%'L8Χ5���p p�`X���'�X/�x:t?���{��r~Iz�n���R�䔟~�g�"3�6�^29>�G����a�c!�M��F�?x�
By��?�y�K�ǁ��X�R~���R�y���˯�T��Vg0B6�&5�U"{!M�Nsx9֔F�G���c"1�:�d����8�1�)��S��NU!?� ���S���SMS~:�-�C�Lj��������R/���xz��v�X5�MO�a�������3��Xa������J���n{˰=+�@�z1�����/r ���Q:�s�Oq�r���顯��&$ܔ�}xt�<ap���?�R��N�1d4b4Vj��,�a���)�F �Þ���:\�S 8����<�A<��{ 7|*�w�Y$pX��U������U��f�g�!��P�S��H��̀�sr��U񒦶!�YF q嶩�hö�+T�h���v?I�N�pbc �GKL늵aXP�����s�J�I�����c��C�?d�'O?0q��|M�|Ճ����d����3�ʘz#,.W.X�M2��y�t,Sb;{�a*�X1��A���'��x&�;H�������?RN�߃߈bge|��VE�`��&�������Z^@���?�ՕN�
	:"v�C|?����������c{�
j�
�Ӝ.�:���������T�r��m��i�.!? ��K�t8����å�#M)�������ё�70�	��~��89uR����[��R%%���$��Ѵ�hz�j�B���+O�%����n���$�o{����/��WR��ߎ��7oݒ��NH�JfN#�t�$�r��K�Q�ra`>��GAy�ss
�4��4yl�(G�r-Er���?����41���KG�a�<%%y�5)]�F,󉥘�XJ?��bkT����F��׏?Ϯ��f�9�����4�f�b�!jw3%^SFo&�C���Ek�ǀ1ỹ���31gY �=^ɂ�j:Δ�	 �0v��e�nD���Y&k|`ʟ�S�e+�1��O{ÚJ"Q�{+~�-�
�!�q,�k~*VP�U���`�L�L�C�/_��s��D~�L%�}@AԽ�^~v��O��\&{�'���i�;�7��W���߰�|.�7~�DE#)2��6 �Q?��:ܤ`AB*W�6�Ή�(��yP)�Ks��-�U���@b6��0�W�����	\�\7$�p�G���Tl{f����9�i����7��A׏���b0���P�eË�C��^�����(՜�a~���@����� e�NF�u0�~X�G�?1鐟t(�8���Q��U���μ�˽t�3qg�^l�����TBa�;5�m�"j�%� R	E}��ǲH�S�~=/�q,#E������8r�D���^I�8WDی�0����d�r;���z�98�x�����hu�ǝh@܉x#���<��u$���oR�kv����d������s���^-W�Ir�=�6�V��'O�1%5��_���i�h?Ü���
���*��8�x�l���.d� ��C�
����|	��9Vẃ󈬧�&*R:�Dʁ�f/���f�2(��fǄ�A���?k{B48�ٳ�Ⲇq����T�� 3�DME�o4��/<ΨH�c ~�<���ݽ#C� n���X?z S����t�	���z���d�CRo7l�؅^�We���(��ŘΞ�P
T�"�X+P�~��%�^�B�FGS�0>��o�FPp_bY���U\T.������l�i�='�|"6�<�P��JU+�#'��7p�䴧�u�Y�.ʥ��}C��g�D$�I�҉��$�`�v"�8 X�[�q�z1"������o��N���*B�0�{.N��L��#�V�8��T���({���  Ԟ��1K)��3D޿�,(s��^��)�D���T£�F��5B��� �HB�l�/�����|j��`
�D��~I�ȍlr#�-�#}��cn�]�N��ў����Q���:��@~�Έ�ڦV���n�{Ko��F;��{�I�+1!6�ӄC�횕�0Hj�X�Œ�`��cJr�v)s��m���Ac��	�Z���`�n�%G��'�Fo� 	�8z�*|8��u��Y�L�I�r���Ǵ������n��3�AF:�7/x��j�Rz]/��{��z ��(i�NU�&]�9'~��A�!�?ͅ䓭s�����T��ls����id7"��A���ʆ���~�sE��w�����s�U�8G�ٓ��p�N{6�����#&�MEi�4G�a�l��i��P{�(�<G�cn��M�t �A��1b��p�}�`Nr`Oj���=2���^Ҝȁ��1��)��,�oU�R�;qoD}��:�t�>����_f��6v6�0<�	����7A@
����Q��)������ |��Е�*:w~2�kYG�����)�y#���������� �(�ſ��d�%�)�~�#�Z����\��9�ju�8�����o�ƳY/���|V��G����*�Y�(���X�u�.Sh��;��")U���b�ח�>l��
x�x��Ԓm�
��!#{�Yu��*��!
��~���o����w:���L�V������Yq ��  dAi�8�l#׽�!o�������������[Y���,�Ap�t*�=�HM����:MhM��i̘��ׯ��QV'A�t�EE������Ux)�gi�n���K'�3�����,�L�l�'�����R^3�.�YN|��产X�U���O�P5�)���R��F(AI���U�Ky�$�w��1�h;m�`�zs�%�l�r�TH+�[@#�ѩ8�s=K2>���CP��G����ى[��􅘯\�����T���*f�uF�?zC3���|��ION1y6�5��Mg��<>,���}�
?,ޝ��w@�g�8y��������+�%����YB�B!XU�`�Tپ!�L���y0�jp���� M��B�f >�֞(�%v��cDi�)�`�#ǳ2;�i��~�� W������,̫7��ZP� �}�]�O�o,Do����G�������@X��p��e!L�.GbLD�F�{��ώ��4�%��B�����?�3f)�I�����.�) ? �#�P@��l��Z�"?O�# �CR���~(�&[�[�؎�~�I�w^�R&W��@�Cy��{�)�݋S��t��ťF�#��P�[:�w Q��P?8����k�zQ}#D��1������>����<��eᐂqJJ�<�0Z�7(�7Gj�
&;�o���,�L�6�����-{�3��+h��O��;ԧ���H ���7Z%�V=�0uƹ]��� I	�X|�{�u�D�#`&7�C ��/�&�?�����Q��@�B<z{�w�[f 5�W�&���)l*�&���ܐ&�AD���ܑ��d" ����P|#t�r)�W�@�g�����G~���J��:�M��Ea�����hQ-i�-�IS$�rZI�$"��������*I�Є=i�TO�,���9l�D�f������^&� 0���j�*��<�vz!5H�0f�ъT@��Z���r�b�@�u��=�������C~V	H�fv�ƊTވ'��{~w͞�qD{u��B �*�;^^�d��œ�3,^Gvs~��M:[ӡ���$��y�I����P����t��g����1�I�BFt�)p*1�T��_�3ߗcE=D��4�u�rz�W4�#'���=�>�ݩs�Q��v�1P^|ǐ5F�P�L�Z[��y �k�X�gWW��~����{�jMc��,Oҏ���?���A�):�Ͼw��۪�e�I(Dh9�A.C��8^��0n��Y��W� �o���$��cM��Py^ޑՋ����|�������@J�| �G��{ò�WE?G��C<��Z��q{G1K�6���>Q�/>�����Y��h����Lr,>�6�i4���ӜR���y,(y���FmPoYJv�d!�
%���z���lqO�=�hb�r���{N�D�QJ"��Ǎ���$� b��$�.Fc*��׿�g���YX9\����Y�x8�⃨�an6�.AߨG������-�˷�&Ș�;�4U�|�.XYݘ�1;�(�f$�^O�x~�7ި��b]���it��y�:5 �kg�[�H�ˏԟ�|�mx&��i(M�4�H�š/<=[���j	�OD$��b�,b�q@��)zP �m��;�}-$�Vn�h�i<ՌǡuOM���W�]�x�qM	�
4�Y��>D����pp�uV�X��v�C?Sf������h:�4N�\��s�7S.F%B��=l�ZZ�8S��G
�`a*�)E�(� �gŚa1n�����{���E#�UI>c�a�2R�e�Y��UJᓏ?`��{��с�϶������~���O�̝�S	�ah칭����F�G��a܉"&��J^�]����q ���B�����k~��Ο_� �ơ3���8G%q\�O*T�GG"zLw�����~B� k�Yb׮�ɳ��x���a=0C�s0�0�P�n\�L�<[͈����D]�S�pv(���F�`-�e���譲2DN��P<Wa{��O����.�W��r�"s�ΔjB��C"
��8�:Ey�ǈ��ٺ>���q�{G$s�Y�߃8e�4��mm�l�D3�	9��\	��$�f��w��H�����OM�N�#(��I6���iE��ڲ��H�_KD�B2<g�QG��^>�EG�&b�����8ٳSt����-�i��9Xk,��0����7�n����kEg/���B|�����p5��S���r����%��|�ng7���ۨ�g��#�Ux"�����F�0�6<x�bC+�2�A�#�_���S��|�b�x���k/����9�>���R�����Ţ!؍#�Ҍu�?]�($R�L4�J��S�8/��,�Z������~^�&�jN��+E��Ғ�Gd`k�O�a����:�e�
Q���N�P߽q&2�M:e'�!�"�E�d��}�3�8)��ޒ؄�1�iO�@�� ��}���j#����A��2�ʊ�f!�|�Ӥq�x��cM�1�@�5��#�Z��Xe��TS
Ċ��>m�2�4��D�6��Y�X�z֑�������A:(JD�^7�<�U��Ӫ���Ѐ3�P��(0H7^:'6|�^Ws�~(Eӱ͏��6=�B��M�����H�U��7��ɐ@°O8���T�TG>}jjFHK4��lc)�s�Ė�q+S�c[1i�m?x�� ~޶M3��C �*��I;�bl�i�T:)g��|���W�~�bQ�2%��sR�=/wX:p��|�R9
��KZ��KqR�y�⤲�n+�ݰFjF�N�v�6�?\�GN�
��8�B8��R,��MCJ��^x&�T}�U7����$�E��:����X�qQ:��'��cCL��gojJ�{�lͻ�H���JE Ka	��N%�G���Hn�z�s��a�so(�C�%�0Ԍɋ��+W��ڣ���<} j;W��JWc%!T���2D��=�e�=�WZ�<Z��ҖAfk�y<, e?77��� J�8#S��&�	D!c�fu�΋=z�A���*u0;-c�C��i��9D��V7�LxyW������h�S0�mK&�8�}�&��՗_�.��Ce>�- ��'����ԁ���|a2U���ot�v������u�O,6e��C���_4�2'T�>�"K�/~�����]P��=u��^�����)�dq���b(����jЉ��zL-�^(��P�~S㧒ŋ�"�Ʌ�̡�n�6H ��>H�1�[�75��A�:���b>�ZOX{�7�dN�P�<)�Om�>�O���Q Z�����+��]^�tvy�O*H�Uv��͇U�Ÿ�b�]lǒV�|�Z�"�=!\=(1�_5 b=AXU34�/���a=�%`�dS�Zd�a\_�O%5r|�DRn$m�:�C7�I�(�u�2uQ��!����a$�dT7��¿�6����]>�,��+Ȳ�pJ�jޡ#c��x����9��J������/�C�F6���hm|�N��N�C7Qϕ�8VY��*R��ͦ��������n��/s�\��~�I�Q����L�(Ɓn��:C�2{%�p:�gb�h�� ���0���$RQ�9(�%�賒��t��W�	�DުʢV���Z�X-%M؄v(/aN���ޅ�}�~�O)�sYkg�e�f��S.!:�W�.��c�J���ێ�q�;�I@L��Ұ�8y�w�����<ܣh�q���8h�J�G��X�>�X��R4Q�	1�Q�����YU�^�'��r�RɨQ�OSM�O�8=�4��[6�Q�T/&�C���ZF�Τ���x�h�[�c��Gc?#���8Aw�Rk�Qt�µIjrPD`
0j�EDZ�w[���45�&������)�T�n(
ϢB�̑BP��L�8�GU! ��#���x��D��8�ӓTň�R�o*YIM�.G�j���%��*��=╅��'� w����ǉt!;rt�`����9m������	�l����- ��H-F ���T?�C�����A�B|�O����|�JYl��XO1��ˑk���̜�aՓ���+�c�ѯ��â�1�^wI"Q��Iu�����\�8�K`|iƲ:���\�	�y� f�J.U��'91=��u���bDXp�D�H�$!˧y���sW�Y~�obo�ꙅ4 7ł\L��8��-I���{�s��Թq�6~c`�C�(�"J,J���rH'�$�����E�A4.��Gt�
��N��E쥂�A�2-��o��Q�>�C���q!	��zKN�A:��9!��B>�0W��8��/ǡc����q4 h�h�a�\�1�3��2��p��t+�!bĐ�P�ȹ��|�0/8p�qDH�#)�qa��u��
9窍-�.�����(s����l��(�l
��O�M�.F�|h�n>������#��rwE�dr��r<�:�W
.2��Q!���ܙ�H=����F�uS,`(FG����{�pR��S����W�O���.����b�N�`��"�S��Qju�iN8�!�7�*�ur2�ʣ,ϚU5@�)M�D����Q<.QM9v\�#����ƈ�4�����T����I��eD�-�,��#��rѩ�R�J;�g��q���5�sTp+i��0��A4�X�&%��d��|�R.�+���2}{2����L��Բ LSsQ�_'b��0{����~�\�霋8,�O���n6�Iuы��+68�� ��%3����d�Rı�f\r�k��P��`��2�ݔ��,��6[*��Q�xr~ր��!�8s�@���;��[�2�M�<�jMJB� ��Tm��yb��룘ױ��8�O�m��#I\�T(��[l=e���^w�AjŨ����%Y)�_���yv�aw����K
��=�j�m�q��#,7�M�Y��c?��3�K�}�������Fy�T/>�+�G����7.�b�^�H�>�#��@�,ˣ ���yM��8�S,�	㓂����~D� :��)GҥZ��J"��눙UK��t_HzF�Ǜ��(�jM1�BX֍#"���KĲQ^達y&1�gΞ�Ę�R��tbM�%�=xDw�y��tF4����ˣT|�r�?���8u� d���*r!�.����٣�>�}��,W��u��m`!,�Q{ۆ�M|���?S<�ON-�u&��>:9�M�� (��Ũ`	�Z�H�L�����B@	�tԏ�X������M���;����O����$�5��T /�� 5�0)y7T:u^�뙔��NN�so��;k�J%)m�t��'q<>�<�9��j!�����|����(J1���J�����^�8Ώ�(K��R,���j�zf���r;ܘ��>�Ps�C��ygR��"��S��l(��� �գC�����Ƀ*|
[Q��8�E�,��&>�A�#�M���Mބ����P�lDg�Tj�P������ Y��VH�'�ݏ��(��
�vj1j����x�V�t�9��e�8?w@('%�+�c���uMR%F�A)��{���hO�(�y�N�b����A�@����+�c	Յ�(E5�!o1��)�MX�{PR=,Q؝�}}���Tc��X���n��ϗ�\�(,���(F5m(5_��Wj�C�e)�xRz�ɧA.6 2רe�뺂��z��he�w~�r�6�l�9��z/[�h������z�5U;������81�cB�Hytf�Ձ�&�ԻPt�{b��?b(c��L]	k�X_t�ۃ� ��m��(G$�*��7�H�7�s)G~GE�Xڔ3��\Z Sv�<�0�%��2�3�i+�^2 �Y҉%G�GvO�A�#�p����|��/��!n�k ��x��1�]�M22�]D�*�*x� �NEי�}۱���u���n�H5�
�U<�NH}+��1�g���N�XYiP�h��k�w�5v��S/e�?�9��Ee�x ���{�"��-Q��b�4��I��}�U�z�>דC��))q���" �+Q��򖷁w��E��S���V��%
�$R��.f_dIp|R:�!��&oWp�u�LT����E9襋�e��$O����8C�G��>�3���P*�"}h����#P�bO>'�)�F}�������˄b%h2�u�m:��"(������p��9m�jD�/nF�3{���ҏ	0��?&(\O�=�	�K0^��R� �T2�K�����n�R}?�f��@.�'��Ѧ�Xn�h�ٽo*��[j٣�8���d]�c��`���_�^ih���Zbab���81O:b�F�7�By������Z
Tn��US�&sG��l'����0u+e;���)8��2t�N˞y 1S��{~�ӧ�#��}�A�3�\���W<�[��~�I.��!1z|4�A�0^8^����熼�~^�X�4~xpC�n���wT�4􁡈A�Z�,G#�z̡�_I����'[�~��|��)oj_)��X8R�iD�7�:�뀊� dAQԳr�
�z�K�aWӠ��y
P�U6g�=<ؕ����� ���zc��p�����+�����~�����bt0�3䝏�r�j����^�'��0R�zfz³���!#Syk��$�t��)t��Gٜ�;�sF����d�{�aKMMH�t���MK_�Ϥr#)�}���������k,sd�q
y_�<���ʀ�qEt��u����y-X�j%f2co޸�Gi�쎐\�x���t0���r�/����^=������cýX����a/�m�ұQ'2�n�K2��z�:1/.M^wG�e%8��i
Ay���Ǯ�f)��Vq��^�8ܺuM%<h�<����ڵ+����Ҏƒ�_|n�xV��Ұ�'�UjJuN�4A�F�/6츣�_�8q�^��8�
�L��|�6�4��@��nK\yaI���hP��7ߺ®�Sv�4@e2tl�^���qˌD��yΒ!����b���@�nw0̳z�A�����~�䄇8b��P��|����H��!0�Ϻv��:�@4K:}�BJ�uvyA���T�G��̲�Eͩ�OL�'bx�"�M	+F%Eb�b>)+��T�j_s���A��g��=&����XM�3q����5�T5�xͬ*��GD�P���YP�u�qM(3�����`]QnI�֡,�I���	��V�&d�L2�0�2t& rw�fʺ�בy�r$�����:Z��k>?��ci�i���\]Z.����u�d<|�Q�J0���	9ч�ǡc�[^Y�)������.����+D4�-p�
�㈔����g����tzjү�a)��,Mf>��ry�Gq���2�����o@R�FK���L��R)���T:*���w5b���z��d�P@m��**�V��R�)TB5;uP�bC�@V��+��b�%��nt��"랬%�G<>>����r�ʔ�7�no)�7�U���J1�hJ,1�U%��h�W@�m{���38�G��G�T�C8A���cs|�DD�8�c�hC�'�܎I�0fc�6Ⱥ�3�0GG��v�Q<�=~�D�dL�k2�]�>�=(7��k���O�G�M���2�
`�WX���䧩t)Q�����]�NfW �E�(EG4�u\���>�,*��$��qO�����e<Ƒv��{���y���b4`���%D���s�O��#gfbn 7@���l3<Y�*�W.���^<o��M���a��x$����`L�Z�,ǈ�,)�F�S~}�j�g�=/6��m��fJ��u�2�(J96�g�Dm�0u��oV]̓���Kx�����`�a���x!�ŋ�,��x�]Iʜw�_�\�����i=0J�Y��ٙ04��?a�"p��I��b�N�'ad4L/i�Z[�9:*K*��i�����%�!.�q�
5�<��3jx��w¥k�E}>ý�c�Ut�jq������������������ZPn_|��q�81�1�� 0�
B��?�Q]c�m&��O���P��V{�����V�g��8ɱ4��h ���[�:�B��Q�z�Xv��f�S;�S�j,J"��Qu
B�z�|t,�#A:���t
�j*}��D���1�i�S����|�x�j5/�ݑ2��2{��A>��G)�4oc�ǣ�Y>j��J|�����y�f���G��GtO�Ϲw�^̗��I��c{i����S>�1�(}�7�3W���Y���J�1T�(2����bE�C=1����RU����v��¼Dia�nj�Z)L3�!���O��>c�Ӕ������s)=����구�b<��S�'�Xy�0#9��w4*{B,�$DP1y�CH���h �ӏ)%������A?F��Ĭe�؎���ɔP��;wD9L^#�����#�e�@�T�|�����PX3:�>z"ЈC��9���]�tJ���=�6����=oa�h�hDF#l�z�*H`����aX__��u���Q[C�@}Cp����@lMS�X]���@�,c!A1�
��Gf����0�NS����8��	��p�i�tcA22k.���T�d�"�i�ǋNGL��2���$�X>��ЉD��z�؂�%\��J>3�o)�#mp�b�������P-H�C������F.eR�3j*�/����6UO��iN��-[F�+�h�M'�fnO��::�@e�lMIɳ�5q�`��J)/�!�=��g⥁��ZҌ
�k����[���!�U�2\X()��Bqd��7
�5�ik'&z�ށJB�����
�t��aL){����?�@�N_ll f�߸~SG��5Q�e����ǰ��əH�Q\a!5�#kҌ
,/��:��~VV�˟p1}(�bgo_3��~�=��85c@���� <x�T�|7���K""�*׎h��
��gT�!�@�SHHe9��#$Q1]K��W�cӾ
�Ǟ�&!�{2˜=p/޸��=ӂ���P\�Z�2��zw!�i��4߰-6�b��G�-�!������Wr��2��6f(Y�1�^o�TU��K>1th��?��WΞ�u4C�������_�"�x�Nxnb	�
%δ��3��{�,N_����.1�nd��B���˕�t��(�3�������~^�>\��U���e?Sо�f�#�� R�z�}�F2?(<���h�s�Ȓ���V���?�1Ί�_:�	��?ƏY�kb²y�ۦP�D�S��A�VT#�J��g���1�Y͠��<��ta��+U��(T�g��D�ߺuC�QN�"s����[��vk�,����!���F�uO�������O�{p�yfי�͡�V�B!�� ��&;wK#��3K��`���[���n���NlF`�DΨTN7�;����n��� ��������ٛ1��u�o���mStey1|{Kb��#��Uök�"BcTR(�b���NoDTBT�c%<|�Xe�-������z���8&����\�[�-�y$�G���WT��|:��s�g�6E��D-ka;�e5���*:L��+4S�[XB�OA��ƚ�����08l>eb$�{p7L�1��f�f�f,��rPatxhT7�5b�����t�ظ�0j˶�A��m�Ėe�Ǆf�4�Ҍ�|SZ��zر�/�s��7|���~8��@=�
l��]��\4~�M2�?���j���V����p���8��%SJ���0pD�yajH�3s!�ZN���|�P�<�ytU�6�; �l)�+���F�V6�V%`Ak�1�d��)��̟�nԢɌ�[,s ^�ˌW�]3a��h�d2�>�_9X��\J��@f[1�T�aO:��טG�A"R��4g���	ᘿv�eGJ6�T���� �ad�tŒZ�}t9��.����G�h~�VoN�E��+�m::pnu/pþ����ͺ"�۷�I���\i��p��7�w�l� �1����>������ճg�2i��˦T����9�g�y�s�^��~!{E�1;;�B((]`�J��5�P)���l��@�*�u!�:�} K�D	���,9> ���܉ ��~�|C$2N����	�٘-v��I-_Gx�"Y.����Z}!Ac�0	�LJFn��8���vH�Pt	���w�?
ׯ��	ڍ�ÿ�7�'��������C݌Đ��x��I[�ez-,Ǝ��ZW��i�nZ���}/�(������p����{�{_��ǟ|bI�n*��Q�zY�
nF�]W#+�oQS�����a*��zͼ/-��Z��+�l���G0���O�ugD+Hh�����)���|�Hj"�!'^EgT#lf#9Ul>���$`�r[\Q����8�I3acNҚJY�~67jB} "�?ܯ�m��$J̔?s�X9��r�rq��P����)r*�����F�!e�8�v��$!��#3��ͪ�1�q}�'�WWkZ`և[�$�AX�j�ـ�q����T*��J[�:W�RfK��(��\7���ZV����[.�9�!枹�&	9���1����N�G���#c!��}Nj	l&�t���ƒmJUfjr����Q<c��ٳy��J�5[����ܹ�)D��VI:E=�E��w>j~�l~H�v�/]��N��<7?���z����6�W Q��X7�Ұ'?�M� rT|#�-E�GǬu�D+��|�4U�@�'�;�ߔ$���Ʀ�X���<���S�-�L���?�(�L h	 ��Q�=�U�Ʀ����|�+��vL����H�d�"1�� :J������ƂrHn@b��q�I� E��a���E)����A7SȂ���LQ?��O��������?�/é��L�A� ���C��6�:���nr�Ty[PV)�T'+�G1�]�"aG^g#��1I���qQ	Uu��&dq)/S:�9����1�<��?�i  cǗ#�X:�5]KP@�%�Fk�~�fS�R]vѰ�Bj~g3���k ]��>��4���lJ�L�Ӭ�d�k4t0�D�, %����.}�Y+
X�nd e��z�g��v�A�,,��YY&�6$4t !�)�*ab|�����'
|���֟���Ǵ[�-p�L}ZXS��/M��)��rY�G�\�g66�0�[�?��a�0o����<t���X5�MKw��	m��ڢ���\'l�V @�ot�bP6Ӕ��e����-�q22�(��8hQO�L�>�e�f� �i�d�ڼiz"E��G6;������j���/�	33S2)����ɿAO808jA����-�G���'��t��Q���%�5cIi!W�ν���V���e�8����p���H��u5�����8��̖�l���T_m1����<v섈WF�,��5����mˀ��;<�/�,1)���Q��ɰ�~0Ts����!�+����H�9����p!�{���ʚJ���zػk�I��v���&}�n>��Ǔ����޼u':0&ǎ����dfh~zN��ܙ���r��|�[�ߖ�$C���Q�E��<�9�w���U�B���S��+W4ǈ	z��Y[̂��>ۈ;����̌�-H��6����k������(�|V+��en5{��h��=~	f�����!
Zc��Ld�#������77µ�W�)C�̲����];T�X��θ��Q���d�\.��¡C�u�@Ob��7\a���}����_=<��N��R�w�ȑH3&�6�vlt$r��zzT�Z�o��*�|���~m\Z��Z��fL�cv8�����<0dڼ_f�(H@R2�522�葟�ϫT��ߩ8��D�>�v/̈��e��� �q5���9�L�Pm?���6�.J��[��{�����,E�������:eu���H�{P��g3��0m���V�z�L�	'����
,<z�R���t;���姦�%SQ����V���\&fZ	L��*|.�u:�Tc��o���+�.$3=������e��0�:3;'à�L�=�HR�k7	�e���F@E1�P%`�ص�j���4��)^�T*&.�8<�T�P�&����:=0�2>�l����u�����%~��φ�Nm��;2Җ��jAע��l�}^T��XtS��^�������-��m�	�x%����ɓ�Tp$� :$��7	��/_()��ہ�����n�a+
F�p�+F*�\~\�+�G�y��z�PC�����ٳK�.�Y����l$u;�N���5މ%F6$��e�E�'�ȇ�g��P��;!�̶Ɏv<���=lW��DYQ�.�V��k����6���'�����RZ��0*�9PZ3+$ev�\�&HΝ;�ȇ���������֡��>�͇���,��R����q1C�)f;|�w����I3��2�E	�x&9>�M�g���g�ӟQ,fz�LQݶ��:d�DyD�B�ح����&c|�!�
	������5P�T�k6�z�]�t>"ͽpV�-���S�&s�%����V���8���=z��!��-����ߗ	,\�!�����>ᯡ7�c�D�C��oߦ<Hbő茛�g���W��{�.�R�,�����0e?#	O�SF�(�:3��z3$*8�Хp��Q�Z���Q	�V�Wl]�,�\�H��x���r0�[Z->;�MH�&_�vټ��M��Wi�E5��7u}�lw�w�4<��ia3�='Y���^�ܾ�(���^Y����*̦L��-��FH�H<��zS�{�� %(yN5�e>k���� �!JBb׮:eW�]~��K�#����Bo�L��BSJ�O-�����|�>Qq��9��[J1i4�8��0�\Q_�k��B�a����̏��*M����(kA.����ĕшk��҆l���T��~� ��{w���H\�E��nO{yI m���踅��ʲ����r�z	���A��aS�d�bP���[��`D`�%�l�#��a��=��8�J� �D!���W�Tm�!ϔp*�����N�M����I�oܸ�>�6w�,ü-dZ5��JV�3�o8�13i��Æ�r��5�*�К�&y���(�3����=3�S��6��z�X����5K�-[�n���]�`����ȕ��n�"c�G�T(���Ǉ�}�JB*�~�&"#�b�fN��D��|��O`���#����E�з��J�ݻ?��^9����ou@H���#��q�琉����b!��ɵ�6�@(�����^j��'��?��S��0�T�	<\TyE3��Eh\90=�z@���Wכ{b˳��ڑ��;I�������z��^��T����I3�EC����RDSo4z	t�@����LrҢ���Q�ՉS��U;$�R�5�.����1�1���k�����J�h��29 ��4 %ZY��px�ZP���&�f�6%�y�0��"��߉�h��w���hkˑ<�5x�O�L��0D�����{�<�8VMohj���R:�E�"M6�n�{�(>[��KP�#U�E=���)G|�.F��9�':EP/�� 	�Z��ʪ�#	�M�?nkG4����b8`\ZU�VXYZK�������?�|iTP!ăA@�@D/|;�i�d&D>��><']�B�&��y�T��?T�#憬��T�m��c����سxؚ��1i@E�eb?˧�й�����U���%���]G$q�=S�H� R�,zr�/f���e��9t�px��u�AV����[�Zh4���..U�ЅW�n��/���=L	t"�eD��Y'~�|V�F����{[@K��kk�2,D���|T���8�l?����V3*DL�����W�
�.^�w��)�3�V�W�'H��~&�sjŧ{��v0^:}ZU_�'aO��YV[a��\jyn�E��q<������Vc�SRR���Ȕ�#��� �N�f�<��3�Aʆ"���qRʀ���9�tj8���~���f6�T`S�V���V�Dp5�Y�3�w����3�U�����yĶg�.��K0Ծ��tUڂU���tj1d�о^��'�
�0��{̊s�CXw�౦�N�?$��	e'<�q�)6�E�C�����!ª���**�֪>�OR��H�Q�H�U��f�q`ǵ��#�[;˷zܳR��On��2f���q�7)1V6i��af���a��frNٟ�j���ܶ]�6��fT�⦺������a(�]��C�\���J$�_>����c^�H���\��䓲&��)���~��G7dHξ�l�6�7��(��GL�@���84r����?�קB/(��o 7'�̒�n�I���:cE"�����(p����)�M!�#�����S7f؍EA�jq����:@7ڷTz�-�CFb�2�.]�T�{�o��w�牪���q��Bɵ0 y�v(�)�:��W�������+g\�A>��b�䷿��ݖ1-��@]����~���T�?�^�GX���9���x�r��&�O��㺃 :V���W��R�ҩ�~�KeV���e)��Z�7-��%�;�����Ő걎r���m9�Ro����5i��o��>	���߈�	�<��t�ٽ�p�x�B�Ǐ���'
Y=	�]g�'o�:�B�tZ:�_]�(�Wa�#�ȑXJx{A��S�#�M��،Z�)�D@�z�L-�29�.J��C��CH՘�R��_�Á�xK��I��n3� �N�0,�"�rc���H0��aC|Ī��fQ�YY��:�~A��Y��/��o8�X�SG%g�FJ?{������>��i	R�����;u�D�o���8�z��p��qs���1�WR��d���m�|�+{������߆3g��e[��}������}��pĜ4K �q�FrK�b���:�������m3q7����z$x�kz^ ܇�������>��/D�#ڝ%��A�/�Zd��w&�����" ��F��e��o۹�%&��tl�Q8�)�:=(��9��]��̆�;�'9��s���
co�:�Ν3�O��w����<�s�m�Z�%j��aͮ��Y�fr�����ۊ��T*99R�B��54��`@���4N^�概|��w�M����2<4��]�D�WOr��1�N�����	}� �'U\�DP8s��m�DA�Z|X�9�0�!1�6j��JN��y�!K��We�>��I�=)?g#��H|�3Fdcs#Һ�ʂ��S�0D�5�y���f�[fw�<�{���_�);p8�<{N�Y�DI:KB��"��gΆsg_�+�ϦB�ʹ��w���Q������HGP�O���5s�͟=��k�v�^1�[�h�����9E�>֝UB�p�3���:���yU��|bfG�"���I�B���F��$̷������DH>�?��ޘ��:[��^ٙ�D�H� 8c�k�%gE��U�L��.ڝ���|�����Ri \�r#�U���ᚙX4�)(��Z�|��8E�;*��}]���e�WT'K�������������X'4Ge�Ν;zY�2�E�7N�yYP�'O�*BLyuuC84:�X 6�⡦�]Y��0Qp�������[�K�К�#0b�24�,�czwՂ�+w$����	������2r^�"r"-N;�F2p�H�fO
�T�Μ&`m_ɂ){��rea�B��Po}"�W����l�ێ�t�^Y��,
�{g��f=�F����D�>�Mc��֒0�XKY�@�c�> �Ϥ0A�gl�/j��z��K_��d�))m���̟h��A/���Qϐ  ���v�u/���u�Zcw����zb�G5i���v2D:U�Wr�f�����f�9�P}��o�u�ٜ酧�sF°݊9:N�6|f���"��`eI~
�/�C[��KG+˥+f�������#������ӧO�$R�k�������Ӄ9z���R �3}�}φ�A�=H��F�5Rx�(���q�4�*�F�%�kd���=��s�#7}Nj�>�������2'j&�\���i �o�^��gs�Yp����`��@k��E�z�(�,BN�BsQ#	t+��h��P}�md�!��ȃQ��+�(Z���|�N�>���'?�������G@���f~�� @������Y^]r	��
,$��cy�*�Df7�nQ�y7�DZ�h�0I�v� ���&�r��8;��J��@m�I��t��*�t"�-�k
����� ���搳�8����`;̎��:#\ϩol��@F ;��AJn�3ā���a�Q���$
����!4	P%�BG�y���dN)�pp���9levN%����^P����z�9;\�6�Iԭ��6�g#}�W#�0m����d{��,8��gy�|���H��<g�OB*�
��nyK A.3碧Ol�50��� {MQ��EnZ�.H*���cԢ$�r`ݐ�,�,R�L2i>;t"���5Cc� p���SK�#,��$�bڶ}TO�I��Y��̡�r��]�-n�tpJd����9$�ΘW�3�p$�e3[��5��T���Q�$�D�v�Ӭ��
��ea��q&׼�MSbY����([�1�l �!�����a�ўH�q]����]/�W�TT����cn0WRHF?��39,������ʼ>�/3�|a^�a$�lԉ�&��vE��R]H��6���Y;�)Ao��l4&`I��5�0����%	>?�%�J(���'�D���:t
�?h�����e-�@�s�}�L������ㅛ��z#lJ]�M��w ?����뫵�ȁ'%�$��&��Nۉ#1O^2��`�E�&4<6��G?n��,�:�}�bJ�3�A�l�.^�`�΢���6^�ȑ
��}{��|L=}���9Wș����XT�	��h[�'yCu������?�zyP������q�p����[�БC�~�~��0k*�on����QA� �Y��x��N��T����3�B:6�ÞD^}b���f`��Aj��8�d;��D�G���zVމr��N?6T������&W�.R�����r�=Y����|t�T
!�۬������^{U�Q6�&�d�,�������%>SQ�ߠ0'Q�L1���):�'|������_�\?v4<�P���_�QE�֭�Q/�-a��j�_���0�{HrA�p��%�Z�y׫�$���&����`(ȋ�^K#��z�#4����|]7���r���g�n������ 	Ǣ~�VA�E���CJ%y-,�&NHP�F�ـ=� q���Ts�}^\N�Ç�\�)	���������$���{W��xͲ��;-Y���O���|C3��r0��C�_�B$�)�8)Ⱏ>���]U�)�xyd%�`N��?1Ŭ��g���jQ���@���V���Y?���׺P�qrO�eJtW^���9�D4E7�Įي�Q��>��f���	�l�:���b��7���];5���1]��Ǐ�g�b~����p��d�'F���A��'ɶYPn�ܵ5L�zX�lz�n�.��SQ�R�b8�ƶ�ο�Ţľ��޳g_�/�r���gN�E��h��'"Y�0y�+$&}Byn]B��;�"%!X�n|�Y�m�ZL�&s��
u�?�[>#�/���!=�����PJIW�+Ƶ�q��qhǹE�,^w��la���nȫ��&�	q�����~;)L1s�K�ᓶ��	4$��G b<�!�����.d��@/�����m����/.�O>�Ğ�����'�Փ'�#q�ŋ�d�&�~���o���;
O������
��:d���1��F��M�)a�9��0وNR�6'��B.�����T���,1.��D�r�;�J�e7'wMD]�EMAu ����K�VTE�6D��?~�s1�:x |���2	8�=�h�J�D@����5պM�.>��~��脝�gv[��P`&I�-��}����I��Ɉܮ�;�N���@*�'}a��t���f�&ë�N�Aѓwb�cef����rرP��NۃnrB�/���~3f�lDXly��ہ��Г�.bˇ���h�5��:��-����퍜���$�v�صW�D{4��՟.�!f�DowS����M�I6���|qU��g���)��{�7����B�8;0&���K+c����7n
x�}�v�X�]�F��ᣇ�F�D���ů_����RtP�������xX�Ϲt���M3�9�2�7j� B+y{O��@��pk!��AH��t$N�|$m�H -lN]�S[O~��0���*Ӄ�n�`�by��Ji�S�9նO�������.Ӱ^_�d\AT�!Mf�½������UA���EH���ۏu�0{ ��X߾;ܾ�4<zz=����m���V�[{��Ec��N����̈́�v'�7C@��޺uCu�m���-"kFނ�y�-�g<z�<�	W�t3ܴ@Rɍ�A�i/[�Q�O3Z�T&�\cieEEW�6`%"*�Td��Vun�ر-)SC$�3��}֒�O+�����ZOm�E�6'��v4�?&"�ݮ�l��`�Ʒ�rn��U�����7{@	B[�N9� ���D7�چBjj\���r�EB7<��ei��l&��� �{�n(o�;各5ԋύw�1\C��-8�t��q�g���m8���[H$��:����#Nz+Va��Di��"�A�aN�� �
�X�X���^�À)%��*P-�o���W���D�N����Y���IHIt��y��Z����e���^��nW�U�E�Iؘ[wnhc���҃]��?�LC�26R�����H8�-�o�6#�o��������e�h�j�}D�<k	g��@�|���p����gD=S�$zT;U����aˡh@u��n����2�tչ5]�������ʪ֢l���z`��錞�e;�U*�_�7$���Q�%�U���O:� RF�&z�_��6N���S����;$fѩ�1�J<N-��2�!B�������h�-yjy��n�[���ݒ�xl�S�[j-�38����67��>[��(�����ʴ�� �G�{�5Ad]	t ���tG���(¥�����"�̍���l3�������E�t�B�w;����oޕȔ�-x��)$y���>\"�g��$sT`;�v���ł2mg1X�Os:Y�z��B����3@��rc�䤢7jW�Q/~�ĉ02^	�͟z>~��2퉨���1�T�Ep�|l6�Az�ϜSDR��5'Wr�0�I(%�UQ�+<{��Q�J#>?��7{} �M��U�/y�9�N��#�����y�$�N\�����E��7���T�A�_l�N�ܱ}��O��Vv�O��pR<$sF�M�5�]���D�����򻗢��3S/]��k^}2���-X��בk0�IY��_M�`͈�,N�����)��_�5փEP�\��lޞ�.=��jY��P�댳�7 �憳���u(�3N���g��k�:�L�5Q��|�7��-�����Jd���8�83����7i��Q��m	��-,�ں� %u	�>�����J�΄��y?�28�HI��l���������{SϞZT��=>s��L7q3`;%��e"��Um�`!�D�Ad�-��%Ε��8_6I�k�OR��As81a�(?�XP��萸L��Ll5������X	����3Y*,F ^Ƒ�N'�ðpDL,�
���GN����s��_��_�_|>��c-t���o�!��'�.|uS>����D�:yJ'�������>��ɓ�Qi�q�S����O��%	�s瞙���5%J��THĸ�]V��p{���uM����3J�hdtT������j�F� ��K��J�ԤM�\t�
>�~F5�x�Yk��L�{Ԇ\�ć^:`��5$����8���x�:+^YehdT7�b�)=~��#�$-�@_)���Yu	��'h���Q!Ů�>a��4���}J�u���)����*��cz�� 8B��N��������Z�3D��r���P�@�i3c�l
�y��.��Lͳq�œb�!}D�?f��A�x�N�O�(�B�fc�%)bÎ��3g�ʌ��=]n��kJ��^�C�Q���ڬ��8N=�n��Y�c��FQ�b��Ͻ����Tg�gc]��d Ԏl�C'�����'�:����*W@�����C�4A&>�k� j�����+S��,��E�DTZ�ߌ�-�Y#0TZ1'�ɚ�CDȩ~����]_0�F��D� "K>��`�6Z�Ul��Ƌ�2���$@C��� 慲�6%�#���T��X���E�D�;���4},l�sx�,����'N����2�8u�%%o7�|�?�ף$�Yן��|	961�����9aq�ج/��2L��N�)k�X�&�`�|Ms}S���t��lg\*��Dm�I`�-����Bĝ�D��+?�U�k%V�ki��ڕ+������� �HG ���f��TȽ09���ı�c#�]���5,�a0�� �M]�p@�_|&���N�n�-�}�:l'��8�dȝ�s�cx���z�w�9�8fֆ1�,x]n'����ᙙ�;���������
�ю�O��q�u�5C�@��~S�_�'�C�f��qțG�\|u*��[���S^� 8��r����㊝1uȻ���z��6��"�!݄&<���ܚ(��/m\����|1��s�	�g���m�'�S�?aЅ� @�[�n�M�m���/���G}
X"���7�юlv{�����kq���h�I]�7����\c����9L�^Lű���,*�"�a��	?���,y�Nr���Bu�ç�Cr�����oVj@��4�u}}Z�SD�*1�ZQWtG�,[LL��@B���3[���k�6��u�-Zlv3���uK��NI����3p��˯�?�h�|S�@�e˝����g����4��y��M	/M@q�~�P@A	@O=�j�@�lKcJ��}B��K��Mi��\���x��|)�;ک���ީKYdd�#�fÇ�A��� e�T*%?��St��m�L��z��wyO��2W�зnH'��%��p�`�٘s���-���?r$%Ȑ_KG��	y�R�i�qh�V�ʥ�Fm��f&`�چ��ɘ�e��+��ڍ���I�S7箓e7�-(�:�%w����C�?#��Ug�8�C(����m� ��k>��YS��	E����s�$ө��`=|(,;&?�F�ɨƆyO��T�=|6�������-�޺Ɋ6�'i��|���)���Vϝk��`aZ�3�H>�� ���/
Z}ue#\�v]�3zd��?��	3���`�CN�0���e��΁ba�>�E��a�drǤP���2W���P��y��rK��`sS܆5�h����&}��?7e��CՉ�Tf��vi�"$s1bcXra����^��M�9bji[p[����@A�����zѱ����S���5��hF�e��2;�V�3��"��k�Y!�U�o��Z`�m�F,�X�L�d����� �ܳk�mD�,)����������p��U]�};��/g�d=`v���_���G}�l�՗_Ӝ�̓�a6m7�L!�ڴ%�]W�#�h�)�#��Io�HK�xx����x�M���
W�7z	ԁ�t=�fۍ��;��%x�BथK��J ���,-
�:L�x|$X3����9��D�PNk1F-�=���C(�q��s@,�s֘%�_|��}�4�N{��e%�(�1X�ƭP��cZ
[{���:�3��ݻs�e��\ ��#�X�Җ��42<(��i�Y� *�� <��K�y��f�0'�ĹBׯ���UR���O�=뮶�ͪD�2�Q%y�7�L�.ܒU�-8��u"��(��/�xYQ֘c�1�xQ���z��g"r��M=X+U?#�̘*)���^���s�|��m!8xD�S�f��-�4����e�@� ,'l�\�A��ԥ8�O�>���8yB�����R�K���U2�U����)��`3Q���҃G���4��NE�� ���y.�LO����f$��:�Q,*:>mS_��6T)ljV����5���Խ��R���EyGև�A�^v�jG{�F^��C�u^�u�M.�y����^u��99z%�N���e�ˉˡ�r�Rl:���ǎ)˽y��~br�|�}����|4 5N" ��$c�3�r�G����ơ���1��O�(�, �g4"t'2Įiaª�]r�8��-�5~դ���F�D���r�>9t3Z[I�Q� ��;�߫ȊM�Hͅd�iu��Aj]u�J�9@vh���2L?#�x9��&v(��fZzpƚA���j#�֦�*��y��/�l��l�7���*��^��D�	GN�|�QrJ%�@
��*�1�����ko�Y���Ĕ�����@УÃ�Y[[��R��"�w�9�A�s>��/����=f=[���~g���t������,IPt�f[�&bt]u����sջ�c��E��=�ܪ�k�=����b/�r���m �Y~����dZ�R��@�:�@+�.C��)A�������yCv�E��,�+>LѲZ���i���>�ĉ�A�(��(�1�� � lH����U<+'9	�D!I�^}��t�F.6����VW��tr� ��	�ǟ� �'GI�$�"��{4NN�P���7��J�E>�/MiY�e�z��E�'�o�ů�b��wĝ�
jP�C��rG�A�o� 7��Ih�W�i���9-r�2�pZlHB�F@��S+(|Pa0 ����-�K�,�`&�((�p�Yʮ�f6]Z��F��S��@ՀM�Ɔ��X��W���0��W�FScE�#r9&����%`KT<1l�z�[֝�iE̗3������a��?�[�F����O�3�	�è[-U��v�ĈN��l���}z� u��M��S*��P�n|���G��"�80���c���:��`9��|7�Ee�1��bNkқ�+LuLD���Uu�k&�A���g��sr�kHP���r`N$�Ѣ �;C+�SKQ��y
���9X)-�Da�uI��E���CCZ�Uшe�d���q`�8�U*9�����^�̙�D0À�!{I� Շe����a�+�U�(W'XY6_���4=��?~���%�R"�SF�-���'��S/�
?��_h�;@��t�}T�y���Qa`��γh}�9A~�!I���`Y��M-4�8�DzC��Į��k��J
L�E.N7<��%���\[r��	�B���8�d9�\ nVr[�h�SQ�I��E 0�Y�	�Cʯ����U۰��z���{Nk76,n,����ŢK�;r��Ȳx�e]�+�DCw�ݕI�{ϭ8z䨐�!��qiN1�Ʉr�l�����F���Q]��܎!KE�KG��P����F��?_��i/6�Ky�P�o�S	<2v�&$�I�L$��q�iYKz5�x���%M��J���\viml,INT�3s֯��3�1h>�F}��Í;42���n�_:�S��������20	�3SX,�e��� +D�t��Ԍ�!h�@���R��l���"f&Q��	��\R#����3��;�S�p��������8JR� ���fcS�EdAbK��LzTc����� @_����fI�̡�u��CR[�_�����g�7׏䆯�eIy9]������:���l�@�D��pJ4mk7fuyM���r:eNQ��W2�o���]�.#��	���;o��g03>T֯�����аc��rG�. ��OY�8����"6/a� �IF�y������Zn'��z�m�UG�"�Q~�ji���ZCo0���7c��u�|ʁ�#��:Uio�
\ݏ�gFΖ�Hß����+*�0��/xyiJ	���P9���'����a%YQUS���9����ݾ{[������-����&mPj�#�@�X�����Y���8z0�濎�!�Mbt�'�b�l�3��l&��_rrP��[�����8�dR�9߽6X���P���ǲT,���Z��M�U/0ʅ�Q�8��,�9\���i%i$�����">)�؟kݒ�fYhs�l��k��v���kW����ɫ�we�tn�T�j7��?�^�\�r%LM?��BmGC7�#���pFs���?����ܣ�����Y��w�M��9ɑ^vscQ'���Oߞی	8Wml*��ϒ����6��t��.FznV�A�	��Jt��nD�H7��RY�
m��� H�QQ��W�iY@h���o�OY��'�U�P|8���Vo������-|��j�O(�7��F����t�-&:�MNUv�@�;5wZ�N2$�<�\���S)Ü0�N����s* Ҝkv:"�-.�rqA&X5���o�����Ci_#�v=�-7�uÄ�~��/�,�N�)>]��z���&*#�jY��N2���I&�ySX���=���6}����6�:���H�R�-�����o�D@v�>�#{չ�	&���`f
��J�_��OH�Dk�]k����ZS�t�Y��왩]a����mA�f����ٸx$��mW�T��+	�.	k�n�{c���bW��������5!M�Uws�PNѥpoMף�&D���^#m�C[2A�`'� �XRdT���Ke3لj�'�.�� 
;_��-[���Ed�rHem���Pb��a	e�\Լ��p���A9}e�9���jL�g�7P�ry�L�h.b+��RI&bh�����ID�ڨo�_�u��JR�lS��dj��������s]�s�D�O���DQ�ވ"�C�M|�*u'�I�� vK&a��:22	��s1b{CR��=r�`�Z��u�U�WVEY������<�M���l�e���t>��F�[ͨ7�����RR�v�lx����R��	�'�ia�0Oj/��f�e�Pʻ.�CAS�2es6#ysG}���X�S����<�W)+�\]_Sv�4��tjO�s����p{��oc��0������."7+9�������U�|��˗ͬ?R��2��Q���iVh�P~�׷/�b�V���*��O8�A]��9G7���v1ϱ��պ������dםT��i�\��o7����R�Ļ�Ҝ8�UYܻw(���V;�qM'?Ģ;zT�4��`��17�K_)_���b����F��䔍?q�4��֭{2%���5��N߻O>%��w���UR�\���NpP�:�(ʹ��@O������.Bw��Ƌ��<KL@��TL�z1m]U� �h��H/w�����'����������^�jg&�	����#�p*j�7��y͎�A�կ���Dm&�ga�~��߅_��*����?������҄�����{�|����֏?�$|j��O~�S�U�V��;�� 5Bz�$��G�2�i�ic�>%ib%`�#хNǵV���r�=ԉz��t�:-��ShK�V���4&%,� �M[���Q9�Z��~1]@M��w����([�I�["9���W���	��9��8�]w@���r���^_^��y������V�Q,#1΀L�TH�$$�I�~ �r�6e|@����w�:t ��2���E�Y���p٩���x{6�����ѷ���=J?'��$���,��r^�T��l���ɾ!�`1=wsm)��iY��v�Y<N��m�J�8U��	=Y�n�����<I���u������ח��f
Q.��6����h&��CI�$m�s^C����l�/�P�P]���~��H�r��~�-U}V�7r�ڈ_�FN��FZp�e����]�'��w1����s�X����ӽ)��x$H�'��R�^�(���l?�Y�}���@I��/��@�(�|As�]�Q�A�IT�K�������`b���hS���$�,:9�+�����=0��>O�7�8�
a�0%v���������[�o)	��^����� a /��,#���@ȌCT,����lQ����݆u��e��OHW������0�}���0-��=`C'j�'
;�o9u�cJ�=޲U�_P<~��E��w��#�@C�$�hB��y����N+N�ü�W���ܒ@q�%��nN�M�ܴnS%a^�\����^~��-��p��Eoq����@�zXn���J���j�8D��Lݹ};�r�L�|.��/u�����N��k9��eՈ���KϤ�?�ֱ��ș"���ٔ�(f�TU ^fZ�Oӽ�'��j;!Ջ�<ܗ�g�{�媲��(���|#����ʈ!`�v옔i���(YAݾ�bv2uBL��d�����s��~EY}Rm[���)��|_��8LK ��ӧU�Y��VK5�FNI�駟)�z�7�1% !8`�U�K'O��X_o�j�J�vBiJ5�n�q9��8�&	�I~�!T(hx��?���{���h2��Dg���Ӌ��s`{�^b�Ad%�v��4�S��>i�/�p��/6�eƃ����l%�����s:QR]�f{�2'Lg�G?�����&$C�����ً~�{��^x38��=#���__���o��I�p�ԋ>�M��w?PO\%�bI���\^�ЦB�3�}�����>rG�bJ�V�I�ZXjU��V{|Z2�(�F`k+s6�wO�XΠ�qfk����Ǹ:LF�H�:5پB���2���ⱓ5��7e� 3����iF�|LV��S9%^A�_~)�M���揟	����K/��'�oiE�Y��3/�������~�.7�ŅRXx��75c�,b+
؋P�����C�O� ��V��mb���Q5�k��f�� ��q�-������j��� �VO�;�8�\�P�	g3��"S�7�d�F-@}�}PJ�?	��<@�&U�''���ݩ�W8���9�;!{!�%������"۴'��HHb���F��XgK���M�"��?R�șB��@>���C���^W��7��W2vx��肋�9uI�N��R�C1f�W�����U?�]���TQ�(mQI%�VH�z��ܽ�7F�+E��TlۦTB��|���N*��:#��!��8+AuR)� u�fHD�|�ں#KT^��vSQ�z?������a�k+
�Q�~���] &������I�K14j?��T{�9Z�8�S�z����g��TvQ�8���C��ƜECpZ؍MU�}a��c���:@x����j#�Hx��5�t\K�[S�lfJ>ty��Dl�p��:�C�����Q�ᠸM��D��H�%>�lZx"�&�qf�,./��bQX�D���aKQW�M�"�h0a�9�8r��G?��K�ơ~~r�(b���G<,/�9u��C{�|���eY�E�]���w��^�^�ߑ�G��3��*�s���H�ڻ庢MBf�@d�r��0OH�½�Ŀi�@T%�|^��ߙ���Jw܇$�V�A�IIxe��Ռi�C���rkF�FE|M����S��"���T�)K�l%^.��eL87���DD �ON��{v�lb*xH���P�%��0��D9⾵g_1_Gy���^Ӏ)��-V��x�;�9*dd�K����	�i<��k�l���M^��'ԫ=	$x8�Ç�`��D��&���e����P�C8��PFI̥�F;[\'��44�P �
l'׉+z��q�J&|�W�
.��U���p�&@0# ��T���]�0uAc�Е9���q2�y�w�r��q�n���ί�?���Iņ�Mߛ���\�)�4~κ
ȭ�]��\{0��IJE>��u֊�23w��U\H��(	�u�f�lv���=������]z�Y���.��H�����m��"fJ���xs�+��E�J8�I���>�Д��M6F'�2��^@LiC�M���2���PS۶��%Z#���ӏ�W%�lI,���S������zVA��eߢ�6s�-�e`�c�W���P-�:�F6��Q��g�ܵ3LK�oA����~/g�hdx<J}�s$$�_E��;�I=zr��x�}�cfyG�g�@�ݎD5��ԅ���r�T\3x�E���#}�&n��Lےec^<�g��0EÖ�'vO=K��"
��f��?َ�
W��yo��D�@�+�3E��a&jn6L�����B��t����͛a����e�<���lؿwG����~�{Im�>bNxL�٘P*����q��U+�έ+*͜�8�Y&�2�޵�f��������J:�%��9����Xߌ$�^����E�t&�%�Ő���c�ָ����>�.��G��4���])�a��\�7��)-� u�J@���YR���A�\0�kLÚ�%4'�U~�]��0-�M{dr��1U߁t���G����������N���q��s;�y�-����i��%�C�v������ �����1�o���rL7��,��AΔ���aL�軫aA5�-r�C��e�
�m4]e'�<p	�k��O>$�^�g�N5�?a�������,��k��'"�D-{�C���v^$,�����	XkY�X1#
}���*���H�4���S�*b�OK諸�?.{����8�(��g^o�)z����]er�N�8e���Ls��{0Q}�C��Z}QJ�U{gpÜtz>RE�v{ �|T�fʗ?c�9����+^��	�o�~]��%�)16���bÖZ��@��:#�	�1�a��� ��Iv�5�@y�Ŕ��%����[p 1asߠ�[�����J�q�U������F	4 n�ޔd)?���.�ѵ�~��0I�v=��?����y�o'���6��
�Tp�7L��;�{�*��C��т&� LG^�m+H�x�gL��\37����b�k�ԉćy��)�]'Ά�~V�6�����m��nB��3 ��P/ǱJ�R�y3-8pgڌ�@��N[�����$B�T	V���f�`m
DVA��b'���ڭq��N좹0rUy�#GN�5�s�ݵӿW_�g�妏�qFS�#��*[g���*�W�f���7l7 �nL�=#��c��l�����b���x��,���|�,���Oj9���զ]�o���Аw4~�}q�d�����Ǖtj�%ѐ��!WD�
{���
:"�O�!]�4��i��3�hAf�9q�`�a }>���|u:i1�b��H�)nd�5��Rš�0ag�`��,��ȏ�hutG2�h��'3.���}.���}^;j��k�9�cAQ����>V�aU�Y[tiUU%��a"ء�3�XJAUI1�-�ګ*w;"=�|4�v�f��N=��$Yu�ےy*�ʒU'�I!_,�ה�B�z]?�%��1�q�uM�GI��ʶp�a�@�0�q����}-������E�p�]o�,�VPBa�XL4��j2�э8'�&�k038qrߖs�0�ֽ�A���vn$u�~��,��J�`��E�q"�,0��wM�p�?$�$��k^*J�[��z�%*E�7�+�5�z8G8\,9_5�y���I,��n�W���Ph�pɖJ��O+b򩨼&v��ح�� E�_؂#A�Q�ϱ���ۅ~I�kYԖ��6����F����s� 3	X��V���Ƶ���Ʊc�*(�r�}Q�=U�ڣ�eͤMckzJ����5���󨹞|﷼y��U�Ai�q�FP�"s56/�ї�Jݳ!~&��[X��qt^W]<gj�~�����!�ނ��I$�Į�3;�W��^ɚ�'T<%Md���9	ɩ��OL�wT9ئ�`���6Re�����t#�伉�&�m����:]r�2"��#�qUDnc�Iar��;�Xl�G�
Ж�A��c=HH��xN~ :��lꅾ���rxj�	������i��pG~��Y����l��X���a`F4��re�D��d�� � s(�(]t%7���M'�p���_=��P*���Q��A�쨏K���]S���Y���B7'��ԅ7��x�M�}�v�T3$���z�	�ygmq����I*щ�a����HK����lܸ�GG@�.H�z���kɊ�<%SRb�4�#���t\�QH�\1,Uk�Y���N[���ZW!�qe拾Iy0�����0��zQS��$?|�3��z8� ��\6P�zh[�>�J��Bbf�T�qf�$�{q�mjw�|�چ��,�c�-�u&���4�ޮf�],��H|��$|kB�D��Ej�z�h�~��f���
��v�W.	яo�#DP1v����VÌyE�>���ؐ��>��D!��3��f8Ô��-U�&�_� ('��5�:\�.��X� �5n7�
���F�9���8p�*��\6D"��G��y}���eͱ3R���2��Q��X7�7�������m|W��3���O���إ����E}2+������mA��a�:N�p����Ӊ�y}��!��Q+%�,{Ϟ�"=��/k�`}mY;�T�e�;��Jߠ� �>&����k}��7�����IQ�j3�c�rg��� ��@��dm.�U�Π�C$��F�-.�(-��u.WTU�pؘ7�3a�cAx_����!�O?���r��v��`G�݌�j7���gX��K���L���̖CT�KPFUޮ��-.��,(��f���\V�fc}E�DQ��SU=�m!Acqv��f��=Q]��C��.?����AC��p��Q�;MM=Q����K�$WA��
1*6�R����y���&	��;��>mV���5����&`b��`��i1Vͯ��5�����k!�2N\�`8�p�;�CV�	>�^Kf�6Dq�G� ;�}�~��{$BU"H����\*��  @L��5)�#G�)z���)���â%u׮|���w��n�i{j���L�K���	@b��-������ͅ�=���8|W���LՄ���>�(�U>��Z뉩���7��@�KP��8?փ��W����y������u��'	����ߢn���u�@��^��ֆh~!�C1d�f+YtL�݈��{w͎�*�����^
��a(%L���G���}��_U��"�LN7��K'�*}f����kN04J$����Kd\�Si��3�=�a9�:}�j�d�!���>x(�%��v�w�K+�!qJ1}v�=ñS���QW�F�e�>׎�X��J���	-��e7��;����E�%Y������Sw��Llo:�V�C��J��5.�)j�0?|_�@E�L��H'KGprl�����+4m$N�
����zU����>o�RиY
�h�v�Nq��!_[���y�Q��M��YELc�*>��Q��f

:p���2�� 6�@$m~o}Ӊl:���MY����� i��o�m���9fn�ڦ��������75��)L"+j[�5R����:}l5N\��ƾ�Q�n6����[�M�X۰��:�& u�O/E,���4�9��@�0�FՕ���O���/���ߔ��VTt�G��e�(��1]U	�Ͼ"�=��b|bW�l}�r� �
}f�Ɯ6)�3~����V�s���N }��Y�5"a��^-�W��p����e�Z��l�t#��S]ZD!,�/h�}G�����_�W�#�Z9D����	�G��8uV,�]�n�ە狉0p°$P��c;�'����.�ױ|���=�v}�k�Veo�dDX�vΓ��$���{���ҥ�4{��%�%�c��Աѷ��
׮^�ii�/���X���cH^SK9��_��ZUdH.E~ѵ��42,�<�������@K��H(�P���C,_�P-�a(��Ą6�*��6O�(��#P�H�V�#"WR�J
��etI���o�q�0W����5ۉ#�Ţ���y�~�b҂#aa� �PrdN���i^
n�|Q�8�����3ܹsWa-��ӥ��D��F��[(��8��ͺ"����M�i��!�L����JvM���UZ��0��>�\QD�>s^����n���xO���gR��ϋXC	"��:�ŶY�d�H��B����T�,�&�x��|!�td"�vU�vM���BمX�2,�=n��6U���^�[�_T��B� ��b����kX3W��y�E)�:E��Y��X �ʊ��9I��SU�+
BR5�Rc❧���Ui��PZ�E��<G�oE(�@B�I��@�
���9����~ex�>:�Q`@�:��vSxF�/�LhL�"�m$cw��Fe���^7J�#a:�d��t����ĭp���ܸf�,�h8�	�@hǦ	��|�H.
��T��-��nz���x1��H	&�cu-����	ϳ&���8L#����N��SO��d������=r�Bg�PH�N�0���WW���:�kɬA���e��g'��\�DA���1�k/4��s9��I��ŭeϿ�n:�I�'O*&=��зRЍ��vT��i�����H�NH����݊�<��ڑ��I�c�XK�+�[Jђ�Ƕ���x9G��A�3xy�j�n��)���?8v���˱@y�ĉ�01���m�: $�� #0�(R�>}��%'6��:^e޽kG��=ba9yLqW��`��#�v���a�f�M����X6��;U"�|��+��B�B��\����3
����R�^��%mÌ�N����w����|���'�w"�g�_�ue�~��^�������-ju�V��خ�(n�_^����Ț���ɉp��I�(k�������^9|����o���G�a���=���?�X�num%�o�'GDg�~뼝�R��/��r�{**�=󲸹|�5<nܸ.^��h�rN7C�Dw��q�ɪ��-�K��������z�~���4�WA�����	�ץ��t�ժ_N�ƀb��E�}��uy����M$>z����#�ѳk/&Q��yHj@��;͎N�өGfg;�MG��r=�7<2n޺!24����>���~�;oi���
���$�#)�0���	Kbɑ<�/�`Bln2���\W�_��v �ȥ|��k:DT `����@t��@��=�V�y�@S����PӴ֢�^�g�A��EK%	��umH"
��Ԯ!Nkt� �%�gfZ�<_��r�┱!| ��wd����@́V�}��������d-(�=����}���~�M����R~������aZt�nؕ�������s����߻�|�M�������ۚ���Er�?�(�@�D�ލaP�������pY����]���\AA]IG#V��4�fӧ��4�5�̳R���e�G��vR�^�.Ay���q�Û�e+��f��A��>%?�(���)��Μ^�N;u,2~G��^����cGUf (X�fYs�#���}�yط�	��|Y�l��Uk~>C2�dƥK��V�o�y��-5���D�:u-���1C��a8���v�IQ���H�P����&Q	���	h�Tf_�{=~�Ă��g��f�Du��r+<���Q��'�lIб#�^ީ�;��Z�}ϔ`��z�RȲ�?`:�@�_׃q��q������j]�?3��ˢ+nU�K�.
E��3B_��@����l�gs��#	%��V��R3�Dg�UVA߄S/yX*����!~�{�W���_�*�M�ץ�������+{�<�b%6�9a����TM*�p��FF���A��a���-���cGZt�����Bᆶ��;͎3��\���E�ĩ'4���eqv��쑠q�=f_�]
����>*?�g�$M���O�,s����̂�5@�L�D8���oh<m���U��1j���`7��@�� ��B%����d�ͣ9�ɓH�:WV�ڃ�h@4�d\�Ň~(�`�=$��Bi]7K�e����գ�#+7?��3�Ȱ��~١�I	��+Hd�\!,!��*@`,!b����p�5�K��zGH@�!���b�B1\w����d���hqi�B����ڈ���A����7�Uc�!OX�n�}yI��g���A�p�oݺ����B�5!�L��~n&�	^*�2��L
s�m�T}�l]`��0O"f �r���;��b$�N���2I�KB��,n�c���Jt-����\G3bg1?t�ঢ���`?��Ca��]�����?�vP�'���[?���T��~���1�d��OW�/~���#h��+8�����P�O{D�����
Oũh�A��{@{���r��>�B�Åz���9N{tdL_���%w���y��s��O��t��m9�5��%��/�H�F~�RO���]Z��G�P�Dtm�գx��/�d�+���&�)�.;4\�Qݙ�sϦ5=D�y�bx�J3�O��ap��GO�����M�Mq����O�D8���̎؅m��s�Th:�5-_ea$�O6�Z]
��!M�I�6��ۉ"��)��c,	��U�Ǭ��>��|�S���4��<"/�m�k�B^�K$��e�f|#�;���k&Ae��)�4#E,7�AD�)��D�m���]+�3s�,Sm��� �����g�Qs���'>G� BM9]��-� l�#� ��֮�Cɵ�W!DG�%)!�~�X���v&�(�Sl;���,	Q��5�k���A�p�fS��Zw���QQu����#6�|F�60$mD#�b��@ 8Q�V�Q�ٚ�+p�1W����AY*L#K%�ܧ��r~�G݈�Y��#ݸC�:.Y�s�Nԏ�nPK�Hԇ��R���x����]�ѣ{��ݹs\}|�J
�`��*��8a%~dfv.<�'8x����p�tI-؊J-M1Ul��!ۆJa�n�&���}���325�ܾ}K4���gG��Q�l�h>�N���p8����H�Ӱ�G앳�q�l�O/��']�X8[I�P=�֗�B��mVQ�2�u Q��0�*��o�
�]y�1�Qm�⌸�Ԥ��xS���Y�#�hayi^W]��;«�^���N?����N/���֞����n	'��1�|�;����4?���f��5	�6��Ս�(g�C�ڟ>y��A��?��L$]K���͈!���i<y�޹�o~�����'��i.�q�L�_�n�*-Uz	퉈�>h��t�V���(�CwޒLƩr�<��LDa� �"��� gzfJ>��M�W����q��e����?p0?�9�D�]"ŶL�!$cӰt�>�h�>�����pТ)"�n��3�T?�geD��n۶�p��~����|�j7Ys��eS
IY�?Y6��{ vڸQO����е#����d��mgϝs���p#��)��I�{瞝�k��K�u8��h��á��p�q���eQ�Ty�uex@#:?�CQ*��a5����p�Wg	���O�)�EU�=R�A�jI��KN��Үs*gf��t�}�m�x;�F�A�'�|cr�v��$<�LG�A[����ǎH+?���������(VR�������mρ����͆v�@�����0��f��~
?FYg���Ӛ s��Q��f�&�(�l�]�&�����)DE�0��	�t�|����C2�����CR����8a5��;NO?��Y���$��<����������&�T-�GƠ������*���L&�2/xPW�Av+n�{B��|E{��V��q"�u�P��5-T���z(R:՛Np��h>�M���}>�t��y�|lܼ��%Q����͛�����;&�������ɨ�t��U�0`��3���*���G?P���ǟ
�J$�ĕ�Q���mc����^G!��bU:AM&���t��v�S��LQ�E���/4����G�`)�)��Ȇr
>x<����X\>߶�zY���Ν�Lb��0d-�ܝ;w��8(�^=�%�����ǁ��yX[��K ��U�~����pއV09�$��n�7�9��>>7���k�n����ۑ��ԩS�F�շ��������z�r�){�=2�T�Y�%��ej��h�0rV���L�q �	>�wfR9P�u#�'%~]�1�-,����,y��'N(<DP�����e&-�%88`6z����%L���in�yx���e���g¹s��-X�I��Ѿ�s�Ϻ~�9�q3���80h�}媅ާ�o� +��NVN�
_4鰙���~G&�\�}�%���ޅh��={��0N�o����ݻ�����h��r����M�8� ��U#�rA>��$i�V�V��2�Lt�lF!o�����S��O�&���+)Ab��g/ �j'�t��n*!I"x���~��_����f����1:y�X@���՛ͷϣH����fԪ��k�n�kd�ν��Y�$7��� _|�m�AM�޿W�I�Dd����ѱ�鍚�Ub�5�l�e�1�u�D$��]A�C*嬦SSs��T��C��#)����o�L��ݓj�5[=Z��%��&��%�[�=�Wg��DF&�Q2�!�t鶦|G����qs��
��m��֛*�(�ܾu3ܲh��#)�0)u{i^� �&�&tE�:L\���N:|��Ө�\R���!�Pb�5l�IaN�� �lzf6|bQ���)�gQ��0\����&(�r:<x��մȵZ����y��GT*a���}�4�����_r]ٕ��	�$@�,��R�L/�4���^3�]�dk���V���r,��b����3û9�}�}	����23��{��{�>�,�!~��������{��]sE�E���df�Ʋ<�n���Jg����C�'�����4ڼ���|FzW� ��� R~k{W����
��0�c��掤�i	,�3!,������e�2:tK�YA=������4g��T
�<����81]�?R���i�3��!� �f�\�v��5]\�z��:��%Q�!p�/��_�|�؊ך�R�Y�tk�� 	��t'��J58dr'A��K��=����,���Dw�E�e'&�U�҈긑����YU�v�j� d�-J��B�)�0�LJ�P�9*\sC�avv;�����KN�"�����I�?�F�=���z;��R�'�	.
$Ԝ�����{]u�j�S����0DgX�Y��:]����ú2˻���|�k*�c�9I"�)W$�����ի��4������- 98�׿e�%܃���=I<zA4����>,W؄<�])�bJ��a��-<�b�Ç��5T�9:N�1�N'� �����-�X�����Y�Y�=�@�+��sR4�3�nwnC'h&#�)�ć�Ӎ�[��}��@�։V|öi���CO�>�v��Sjdww���S3�d��n�[#����"SQ�gICÖ�Z\Wi:h�|Z�H�_8RC���jz[�\ ý�8T��T<m�d
�LK�d��"�7�uv�-�&�u������8ڑxf��ƿAr�J���u��cIg9z�4�T*,�dyɁ55���, �����+�{��%Ye��[��~֝F(�y9*�M�KPWl�����	7��v�"B����/�������L@3-�P��sQ^(���Z���ͩ��ɳ-u��$G�]��Q^LpS�D�㇗D2g�t|c�����2�șs(fіz��A'�GH`q[Z�����	��+�gԂ��7�N��WFJ�Ý�	�����'��Fu�t́ ��1!� 3�J�SF��pp?M����- ��<?��k�u¹	��(A]eOk�#9��X�Q��MP�Ѥ�{1R ����c2P;�X�A�wFN�c��s:�nʓ�{ӾF�L��*U:���������1Kd��͛±���[[���7k��
�k'[�!��Ym�+�+�;�,U��?��2-�ڤ�|^
ϓ��jMҏxgfJ�����iNCj
�@��ϗu�ZШ�@���'E��*M�u���L5>����i.Py���43�;R]>Q�Ѵ m����.N���;>s�d+�ֿwv��0�dhH��!��D���ډ��$+��4�����N�6��{�1�̬�Q�H���ɉpsZ�ۍ�k�ye��E�d�	�W�>�:���U��vt�!:0��8e�M@��sa�iRWi��ө������P��]x��Y-�� (.���X�(UC!�jgcSI<��4���8�E��g�ϴ�<<w�0���aWղ��9i��xp��l1 �<�=����E/Q?�����G%=ά!9,m����LR�u�Q;q�C�S�`������B����eWmxE%��Om�u���E�z^���B>|�@�F��A,�Q�N/ڱ;�����:���K�.k-p��ZE��˶)�� �b�},uU�1f�hr'c1� ���gH���g>R��E��}���AƭVUQ��[�qL��s3ke'���N�d�c��3D�M�i�`nZToΚ����Z�=;9Ͳy4�>}Zt�;5=�%�*ʩ���>3wA�׎(��z�RKl:�U\b�Lp��$4��[����X�T\_��G� ���?p�$��h׵�h���T.g�XG��G�88��}y#�4�sbw�i��%�Ƀ��^���ÚT���N�R����ݒ1a�¤�T	4�a¼�f��C:f�"���iF�Q2&2���;|���֨�z��{�a�����]un�i� ���.�*C�<�RPwxK�T����-:Rme%P��j �	�	�Z�̣E}GE=�=o"�zАj��[4�d�'O�V}^�����CAZ<��d��H��^F���]�ˡZ
��zx5n���y9���q??r0�J��ŷN�n�T���鍜%yqxo�w"\�xᬮ�e*�9,l ���	=�|�;wa4�an4�P2_���ɗ�E/Ϳ2o���eUKlAP��Q�J�n�B�XCt$��ak|���]��� ����'������bS�y�a�cq <���0Hy�8�?~��2���mJ�A��g4���t>]�~M fH(�޿{Ӥ`�>|��@ې�s�8VM߁�GzJW���2i��6����鿿25����W�\�u<�o�S'�K-��Z\�S-c0����8��(�˻�ڛ{x�&^�=r�ד��+;Tɸ�R�$������q�Ą%y}$_���:Ԑ�`"��$Fq3�$4�&�y����B���	9B��u�9x��4��VP(��IpP��)�h���i"�@l��G���~�$����:�O�~�E!�?�㧺��?�Y�|劣�5���Z7�w�r�Z�B��?���C�<�8=�Ϝ.�g�-��q.`�U��(�q���ݰ���3�tFy���+!0�-o��A�����u�A B�4�R�MJ�G���QC1L�������f����R�#�i*J��{�<��)u������zn���7�H������X�a@h�I�o2�m�j�{�����
��T����A�ӤTN����^���%-��'r��>�T�2���@���Ғs���a�x�G>o�B�q�I}h��� �M��8�Q�o6�9�6�3�qU��Dۈ��F��k�򸊊��H�:�?w�t��-ϵL�j�ʜ&D���:C�� [�+��^7�x%�Z�g�%�+J*?y*�^ߔz!���:����1��E$���_�2��+�D�'Meb���!o����Q_H_~��l	��"}�F�S�ɜWW�*K�{��Fy%��b`%?KA��.�*�y*�tO���n����pҚ��6���rL�� ��U��<EN³ @��~�j뵸����𖧑"(�4ۨϧ�>�P:�l�Y;��$�����gSǌ���M㫇����� վn���ɟB�}�&�ל͂���xn~Ʉ஦�ANP�͘p�B��fWQ�}8��y����~�^we�U�u��!\sa4r�X2ߢ���X�9�|.բs��|l+ϺzvU�C�Ɂ��>�N�����c�EA�G��`x� �[�<Bb8�=w������v����7B�`7�Wr�.\8/�9P��`��\}�)g�����;i{���Ѥd��\:t��E��hͧ�������^��4�� �o~����{�p��t��C%0�׫��m�����m��4�WR�#��O�<
��K��=-8����6�x�&PR�t��w��c��C'�'UC�� ��s��7���RI
 ˥�?𸊖65@��hʅ�UY�ޘ��I0���G��ePAp�����>-Bx�����Ͽn	��ͷNbO]���	��+��!0�Mf��=x�*�F:p�pzi�ɖ����Pc#V1�"=�l��Ի��e�nܸfц
E�/��Z%Yrc9S]	9�:�sT 2�T��P��ʽ}��Q�6�7���P*�b�M�ۂA������P��P�f���`��E!>�ۛ�>�*�E�����7�5�g΀V�k0{J� �SP{Ϟ��hϴ�������{AB�d��4�����=M[p�X�)� ��w�9SO��p��Ӂc���%4�9м�~�y�@̃�+_�Y#�>�s#Wu��kR�J�����Zuqy�*�>�IZ=�,���NTS�F�^G����y� gw����b���#i#�y1t/��m�*�-,B�H�+�,���{�ʝ��B[<
uQ)Y��5�2:�>?g���IArqY�p|
Xإw�~G�d��߉��R>x���.�%d��AC�j����@�X?u2W�`��F���Z���^7`�I���5����Q�����`�+@n��vp(>w��ʕ��0���a�xgNM~N$12����u�Fإ���;J���)W�	?���'K��������(��
�F�(������R�E��(l`�',v �B{3�?�7iZ�͓�i�.�&��`��NJ���b���0�CY
�ջ�&o���5�g�8RxD��7�|��B27�K�Z��A���1;lY � ��W�f���v-hQy�� H��-b�ZKS���I	�N� 1)�Gs��K th��v��Z�53���H9��������G�ff@{���U���YEJ)�v�3��jj&��&�MPȀa"��|�K���{��^�d��Rqm���y�{�ܥ���Ȼ��P-����J/;�S�k	�\v�.*�/�F���^����l)§\�~t�沩 ٜ&��L�F��r s^��y�UE˵�EF��8%��#��tp���}^�p-m�?ƚ�,��3������@/�FPpHK�I&�ϐJ��H)E,6C�p�� @�Ũ*�l���=��A]C��ӷ�&pN��Qvjԧ����$�����M߈�t� �����Z8	��g?��a����a}𣫚,���c��@�#8?�����a��@�Esj.���YQe�c��^g�4�q�PoL9�F��81��?�x	OAgm�r&Q��<)�w�f��*�3�>z�kߒg���E
Q,6��;��G�Y�ݶ�L2���7��	�9��;�\T���Gu������1��_��|~�ڽ���.ؾR8͙�����Ϊwc2��K�k��;�������'I���3>S��;r�ŷ�%G �!�AA �OMz��3A�/�-(�_b�������(k��y���N1�(佉=�mҚ�fZ�AB�B]9�	�Wu���d�8�Jk�][��3�"�2I��i��u�4�|+mm�� �-������<�v�,�8<�Ξ?������ǏS�>g}{[��/"�1�淿��G�s�b��n�K�|B��I>�՘K���Ry�,��vlmt�`��_z�C�Jy�:U��r�����N�(����U�0�JG��ύ������OjyR�*��52@͙.�g�^˛z��W�k� ��1���%Z��Ղ�`H`{@��b���%ҿ�h�TV��R�6��J4���UQ��!������i"�o��Ƽ�gf�ү��o ]O��������:�hK���μ{* !D�À��e�I&R�n������n|^�N�O ���c%:�������/ҷ����?��2�7�<ely��-xF�W���?�v�!�f8 mpH���cAXkb2u��Oݜ ��͠%g0���T$,_�Fx���x$G���16�c��~S�D�^wX?s�H>�Ac_�-��P0�T�gL�L�VK�Dm�5����ҕ+�r������b�94�פ��T��^?����	 T#�:z�D�[p��g����t���>n�������β�&�K�P�����f2Q�\��#'�����������,1dj�sY�<�D���uA�V����X�}}P�d�������*��.���
�+R��5uO��ǰ�w&һxP���I�܁����>;���MSߧ���_J�����=Rv����\��'ω5�v9J��yEp��*�ؼ b`;����z��ͨ�@1x��eע�/t
4��l�|�����m!��	���ٿ���Q'����ש�f.�A�!��-,��;fO��sWϹ����ډ���Q�9e_H,�c5�LE����!��n���؈]|r��NE�O�A��s]e���(�H.�sjC���H,��G���0�ZH�
�Qѥ����W�
=��@n����m0�χ�����єk�t,,�f���C�1!:{)�Ŏ���L%x���-�.ᇙ^@j���`?
N�q�G�ş��Xe�J��#n�����e#�պ����2ȸ2�|�!���%����I�A�?gB |	A����
(iq�{Z<n��7Ŕkl�F��IE1�$3�yl�墿���Q��3�x�R5
Z4UsH[q�S�f��B~���I�U��.n��^,���H�*�c��A׮gB��M�ꌄ��$�8,��Z��x:Vnj0���Ъ:�ȞR�lssc^c��4A�G�7����$͈eG�!v�+W�����w����C�uĂ��R�"#Վpp Z\}��߼y���I�W)ЉD�<���>�j��y��^��w:�>�L ��Qڣ���;�4�|ڎ�k��z%������n^���e�M�7�7�B�)�����n�;>	Ȁ�e������7w�߰*��L*��ֆv��2��.[�#Gh.䜰YTL��t�'�>?� FVE��u�q ���(1��4�x�m�2�b_kR�Dd	�ɚ�¦���L� ���/� ��J���PΫv�-�A��J��^�ҧ�\.��y�ˏvZ�� Xc|6����L�0u������?��f`o�5m6��	[\z[�Q�	`g��T�F�v�܊���H}�6�����4{Й�Z35Mək�����R�(�B�&�NQ'Z�*�����X�F�q���- �&�G����>rH�]{s���)��1ԣ9>ǤݸqK��������������0����eknK�5���zѬ#�^�+��t���?�m�h9(�}KAY��U�Pܙ3'-8�-m`Q񻪝������Q�z��)g�t�\�� �y��9�L`�Á�u�3Ft�T�;w�t/�q\�O?�4���h�u�'�t4��W��4�X��s��Qe���no�mkNȥKu�X`��/]zG�I�>}d��"@�m�_N������~��i����;{F���<�;�p��^��?T��kL�͌ax��J[b���+�����z�X�u0t��Oc[Ї
���k+����=3����C*RW�_~�5Ҁ<r��R�P�rTq{i�سr`)����Q�Ǌ3�r� c��w�E|���qɧw#���	9}�zQ��P��6U0I]P�!9��_}`��A�H�B����5{������ 3���!2�������l�M�'.=z\ �O?��l�ց<��8z�l �I����v3�o�G�8:�ߩ��`��bK�g�o�n�������	lc��抖J#���đ~ДΝ=����C��9��H
b&U���x��� ��h[���x���;�˩��N�m�߿�n�v��s�&�Fx�Y]�q
I��1���'���8�~�+��]���9	d*[Ї��fP�C����?N'N�Jx��n	܁���	,W�}I�kb;Nۊm��n;�6|p�x4. �E�a)��qI��\��'A�1Ѝ�a�X�n�HO�<�I;����N�dd���I�c�f�>�/�".�qzbj�bxYT��c��}�����?�ې��E��~�P�fFNMވ��H,W\_�{Ho|g�x�Q��	_�|����b�I�CZY��J���c'<;~���[`��#�8��<:�M:�D*	F���X�(ஔ�q?(P�ݩ��)6��9��a�4�Lʝ�_�i�v_�H�"�ƌ�?����W�1ޱS����//��@K��4�D�[����խ;߇+</)%�%�c^mÄCS��T��\Ť����wӣ���w�iz���J]�����/�'M���)�0�3�e���Z�)�8�z�!��u��4}�6ֶ�����Z�����E�k�+%���qI1]��m	���M���p:��ʈ�j%��1gC9��I�K�LN�>�,���O�v�'�ǈn;굻�Ŭ@��Q�/�������sH�:~��'���E�� �)	���uy/gO��j#�Y͹�5Z�!O�ۻ��:|{R.dY����Mu��,+��W���>��3�isc�N�s9�^����#J�3�� t�ѮC}��@5�r��sQ�4����A/�dr�zE&?�O��&����T������GS���S�z�ۢ�`-�JD��i�k*洮����� ��3[p!����Ddf1�Җ~�6jdj౽���dF��$�};�R_t�פ������3r���n�{��Z3���5�+"��,�ᘼ\Sj���띳���Y�n�O=~�T�\�v��$X͛�Y��B�Gb���|�4�J����GՐEv+���>wؔ�X���\���)E��ݤ��@m\�I��X�[R7-�cIP��޽�F�A8����5�W��1�{ocہh�&}v�jOX��,�JqH������ǿ����ߧ{�t��{J�|��ע��VQ�8h�/@�����:j�ц�$9:��`�ٌs�U�+�&.-v��嫊qn޸)8�'�jJ�����ϨY�)�X7l�w�}��}"�B���'���R/�ߚ|x�"������f57|EY�=5]z�:�lSp�]�%[�.]���]�6큔7wr�)@h�k�d2o���W2�$������4S21/�������,7��~à`�� �X^�K��.�ZX������<�/S�<����v�}�F���mKMΈ8�.�>FZ��PF�1��d�G;s�IhU��6�����Du6�4~�QMm�o-,18�����\�=��N���*�2ZYiҸ�a�i��{#�F�$�����y�>�P�%x�3�Q�����jw�N0��a-�H՜��5�E8\ֱ�B�o꫻�T�K*s��Y���Y�������1նϙ�h�u:~b��¡t�Ԫ�>�������J�Ƶb��5�[��a����j���qM�c�h��6�۔m%=g[��~�J��gϺi�U�)[��'RN��x����lH��@�>��{
SJD�JG��O����H=����4DQS���e(>o�$�읶(@t��S��d~��(1T&-�!�1�	/�葚c �w��yE��fVS\"��Κ6��\Р���J�ʼ�]ض�����ɳ�=� Mel�������pц�hkTT!{�(��{�*�Ǐ=���,j�͟�u�uv�H�T?�80�j{�#uǿA�$��)s�!E D�6��	? ����M�ĀEb`�Y]P�4P�? ����W"@�X_e,��ٞ���=�_�*�C^nTR�����WX2��i��4����9yc��t7�����7�w�6���U�:P���T_�ISS��N��a�`��rDi���m!G|ښ�.�[ڣ����H��
4�B�����&5�ܦ:}1m5�E�?����ZP�<���B���$!K!�͍ϙi�&����6�����������r5�˭���O׵!&��գ����%E��^���L8"����k����Z�զ��p�h�����YP5yp���MgO���tcc[�;���8l���lP[}�=��#aٔ�U�M�T?q�~۽Gث�ǩ�D6B�8{ޖ&D$�!��w�&�J&x��F��ؑ�}Q�W�~������s��j��K��ao���i�3y#�K鑟Q�@���Y\F3Ȼ�H߅�_�᪌=���+t���%z�RI���)��^u�z��6��ѭM��S�HX��I��T�K;����w��[�ӘS���,;bA�nE��c����S�Xj�;P'�w��b��~p��  zIDAT���YZ���$6�L�#��5;@�}E@;����i؟����Grm�@N��[�aR��=�l�Dڨh](����3+��G�0<�z�Gt��!��7�_	��hx����;ҟ�-o��V�Vb����Rr�k�~��rZ��ZԐ���P�Am~8�ʦ�^4b�~���������#	OC�ۺ'@�4�(p��w84A�w��B��n���.�J�a伺1a���醴/^�N�j������������kgX������5����n�8��)�K9����{��M���ǋ�)��T�9��PW�#G	 ;��4ov:v��V������H}i�l�g�r�uw��z�l���'ц�4a@m� �i?��lC���\`N�������_��A"2[dی1���@�,^׫W�>Bv�5��6����-�_?�MY�^͌�e��(ݾ}Cx�a� �j�P2���v?��یy���,�L��������<Y��)j����SD�w,��w�Պ�YaԳAW|�ŒJt�Vb�B��V����K�
���>������w۞X���P�T,�5�uWEy�H3�;�H;�LOhzz�
\Ռ�{&�/�Zէ���}�;�ҩ��+p��O�T0G` �Ra��qyx�\����j>T�t��
�vwwSu:�Hy�2ϋ	��s'Sg�v��;������~8�Ǐ�ɀ�������hJ����'������V�L/�h��C������ZFq�Ng3h��m?�yT�*otb��d����]�w}t^�6�no#����N�3��f�Gl�$?~�6vQ��ܒS�ɾC����gO���)� H���!��J]���ޯ����t�ѭ�3��{��/v5L[�����{�呶4/˄�?J�ע�S˝m2	M��c��L=&����Rr>M�}�u�X$�������gD[����*�U0Eӣy��t5鳬��}g��NoWE�cսb��Euq��D��(T��z�aߋٲ$�f�gt��+���#]�Ce���V�H
�gd`ɤ���+��6S���$�3A|�)UK8��[��>,��p��$�Мۺ<,�h���9��y�N,���*�Z#8_��D(z��U�{�H�'�hK�jA��o�6g�NǊ蕐(�%A��|�r���<���SwFR/�VM��, ���f�ˠۨ9��O�)�`?(���1����^�d�	s^��U��`�����N�t�WD�v?�Q5l1���m�oj���b��ʪa_�:o_���(�1!��?(�\�<R�U�Pɤ�jF�+��]2f'%-�^tQ�7�/9��:��7f$���E$��}��|p�[���aPIN���'��N����g�$j6mdGEj��\WxZ�H�^z��"lo���́8�;E�ԛ-G:�� p��(S�1��$G�,��C��Ҥ���9a5&��嫴t`�;�*S��[���P`�Hɐtur4�~���NV-`�]
��Y�}���lorjO^�1D�'���in�~g*���rzl���[����<҇X^��I���`(�o1\�{ΏB� �%���nG	M��"v��~NК�k�.ܖ�U�QD�^95�`[�@�r__����aT���܏%#���B��D���E�R�t��ܗ�'��Ȇ�)\!8L��e�����v�\�!�>�'Ͼ�ܿ�e�8�&�6d�w��z��źs!��EM���Q*�3�ӀB��n1�(���^
S���t� �{��Ն�)�*�[.;G�;�hދ�P�ks� *`SX�A��asZ8�n�T�7�l ���#y}�v_P��_{���]?)E��5M���-xug�����^�$��M@Y����N�EN�<�R9xq������?R�gb��q����>��M��Inc�!H�/�x�����&*�==���'����|-C�L���gO�)��G��>NZ�#L������]�ا�$��G��tK&����-���f�;� ���;��U����q?7.�Ո��Iwx����HX�q0��f�'�`�����5#�U��99�t���rn߾��?tp!�%�0J���,z�����F��j��!��#NXt�Xx82��ʞ�?����?�/�����7���)����i,\ۼ ��c���E.�ni)���>"�Lqu�k1UC��N!J�@�����|h��i �b6��`1N9��MԌ�Pc�:����_�rrl���*C ��ş<{�,��dy�`���-���Q���BT'�X�"�jq���1̌?��d�1XL¤d{�RJ���O���?��)9F�ŗ�����1�S�����ܑ�C�3 ��SȢ�a���~��݇ϴ��(��(������U����(<�˵�4�l�ӠIG~��w��1��YP|k��꨻Z����5?���Ӵ_�m�q��O_lo�&A�pvx.��ǎ�P/.��$������$[�8Y�4a��)c��}LEY�GT]�v��BJ�p$�G�țM�@@v|�=�Q$����ZzB�#�0j�G��<�a��8Y����$Ѹ����ple�8�Ɇ1�H�;6!�E� N������9�33:�pj�����ť5m.��
0^v�E�	1gJ��u����k�j��;@���V�	�Q��k��{���*�xl��HN"�&�w�7��N"�@�]H'\A�7���#����cg	�t�q�����o,�6�_�(���"i<4�&.#9��ԛLl�D4=�;�3��՟���y�J�t^D�/�"K��wr*R�(�1�ӷ��]��/��)���>�Gɣ�3���Q�����p�ɽ��xnh����zC�d�R�H�|��r=Ng=1>T��~eČ�8�o��&��>o*�B�ݼ�#G�,��% !���TNԗ���,<#��I� �����8=��,�5�j!�hQ�zo< ga�i��1��%�6�R��詶�i��&og]��D��R��w�b79t�a:=����q��
B��	C�/�Z��^TNv�;�]e*��� ��z���}6`�%�<7��/X-xy�$�) ���)hL�mll��55Uo�K��Ҿ$�歛��5�Sk ������84� JjbϢ�,��/�ԧ���w�o�J3��g�����G='����y�&Բ�!4 ���TQ����T���щ�}�����PRi�A�oq��\��j>e���;uՋE��l�� H���qH("��N�����참:���S�%�/i'��}^H||N�4�M�dcX<%}�y[[�Mnʨ*�=��Q�#x5m�B�����~������4\���CS�;�PJ�ՈQ�n���Pk*	/�&���*Pu��n�Ȇ��6!�xo��<):��fx�$Hh�T`�+��� X�nϯRS��unj
 D�i7��%��ǇW�s#R3vrT��u^�9��/�m���]��TI���&��F�D�U  D�:�J8dgRM�t����Y�԰���������\«z�4+26�2cN����SI=IS1��bM��#�
i_P�����d� ��_qC��E`��X��}��z�<��9=�ܕ��|j�\eN�� W�i��4zA<�c���"͈��+$EzZd�M"�0�G93iY5�<v)����R�Læ�}�8����ӥJ_W�J��5gN�>�/�i�7x&y�d�q��`�]O���m*G�I���b�As��+�H팂���GH�qJ�v�!������(<��:g�-(���K!ޗ�q2��\+Ԝ�4�a��ڜae�� Hw�j��B�m@�>�>��J��b�����n������'����Fm:O&���r=%�B�TcXL��]���)��T��U�Q��%��r��2����u/��q�{6�ެ;@B���W9�^TVJsz�8"'�}�����I�C��OUI;̂�wN���T�	OHT�Zw�DmAL:cow���S�U��0_!����E�vP�����c=TFkdr~U�έ�G�c�F�P���j:E��!�k@!�{�LQ���]���gZ�������	'�B�[���%ي��d+^I�'o����gX.ܼ�F�I1�!��WE��q�Nռ��8<���h�E��MƱ�X�J,$�N�T�Z��c�S&B�h�n���@�Y.=E���v.u��|9V���YkL#��v)�,1�@u`�#'Qȵ�ܓɺMs#2��4���}@1�V`���}�8�V�z��Δ�%eDv��1ڭ��# K�ގ������xQ�0�I��a�V�u��>#��7_#���2i�U�|^�R0�j���WU�����25Hn;.}��v����T�(�MC;�&�������}����{@�1�>�Z�f�I��ѯ��*�W���f�\94ŨTu��˳��d0,�7�h�~C4�;���d;�>��R����><�f�vdv���sHl�0�o)�B^�NVY�Z�(�k�_�)oC�����>q��`sK������X��"Cರ�k��Q��\*�W�,��8�U7���%#ٮR�h빂6�*T�MSR������� ��fU'�a��?2ԍ�~�u� F��Z�Fͥ���ۣ/�����A�Z,1N�=�ז0��N����ٰ;����p�s5��t�A�l-�=�dk@�н�i�A*L�2�n�~Pq��K����lS�k��Q�W*m~��4K~�R�?r�B��&�kǨ�}p�OM}�[G��w0�(��WFu�i�ƾ��Ѥ'��Zi���=��E�}��4�'M'1:�I�( ᆧSt�)��m�h:u)<3�e<��騘q�W]p�f�b\��R~Cz5�1�<�� r�c�U3�qD�KʟQ�^�Gu<��ǤP�?�e��,E
��ԉ�t<(n�AjJM��T�P����)�S/���*��g���S_�i)6M���c䈎�c_*X����)�7���)6^��zK��**OݙF$:>�?s��G1�+����B(D�c�N��d�I��8�<A֊��dx.��r�甔�̓\�m�t?0�AU�H=��.]N��>Ô�]d�BL�9[ �ȃ�JMpTk�ϩ�m�mkj�(��N���$����NK�(��u��.�*bjpiv�/����ڌ�����>��y[���H:�J]AW�A-�:�~��@��o$��T�8	W�C$���P�#�f!�'0�5�����"�t$z�tyq>֢*�n�4���h7KSU�@���T�D�0?
@���^�.{qf�|��C2;���{�	CՓ5�Q���C �#�#�
�	���NK%T�X��-���Y|�Lz?�0/�M��>�(z�3]����It#	��"şp>�Уwy���QS�x��I�:�K)E]�=�R��c���d��;:�^!A`����A��	��8�[��6��:6w��C�Hc���T=2���qF�pc�n!KN 3���Z������*b��rsK")�L�խF<�im�A�M�&�f����U�=r=#�>� �4�'�=�`9s�c�L0=����Ź��yӧ��@�R�E�
-�']�J�:AV��k�!�!�����<��9����MI��X�����? �4�#���j�}w�졨�e.$�2���N��aFjf��Q���IN%�r8�G�(�N��%{�p����H1ͬ�S�^����>\[}#�Z�!��Z
���½PU����L//�ۅ�vd"颹���+�S�D����&��6L��n:s�l�,N�X�!���E��"���ժnH$�v��v㐓��Ͽ%�FM�'SIG��>��ލ% ����d�h
Rڜ'G�z#�ǎϥ=����V8�yyA�"$E)t%�)~�z����7�Ƒ��i�x�{s�B�3ڛϤ��m�`5M���I2qf�.
	�$A��F9*���2��&��Ec�����O{ǹ�rp"@Y����Mg&��?}�4�:�x|Ig����rH�E���hH�aC�#"XN{��]���\r�.
_��7�*�֪]�G�L�� ��h����Iԃ�|L��|4ZV�q��8�ЁP�c���p]8u��	KXhtE�>�4����=�l*�uѬ`uy-�*�rd��!\3�Zj�������i�|��1/Nj��g�8CD�=Q�P�'�rbݴ��Ciފ��Ѩ�M`B��%��~UT�H&���?�~���34�I��3i���AmQG� /� ����=��i\�I)�˽������^:rD3���꣮ͩsVЙB=Rf&8��H/m�\��H�v��D~�$omy�],�[C �,ɫ{���"�qT�g�p||�4��a���ȋ��-	9 d1�@��J�� �3�?����ReI�K-ƖrQ�v{�ݻ�K����k+[���͖����i�ݲsm9�{$��?}.'�U�J�!(�fO�EQn�5�ݣɯЍ��:�Vp�hE����0	�=��9h�=T������� �3�TF ��8]إA GA�	�v	`�0J�V��q<j�����"y�WQ�\�.�z�=��У�>x�x"5��#��ҳ�6�mz��xh��=Se|��H'x0zB p��b�1uz��	���Z�ʠI6f��TN�&}~< ����ۏ��6�@�&&p�e�xzᲾu��> �*�O=��?j��]�WHc'U�v���}eԡ��L�ϰ[g��=�\m6E���h4�̪h\m`GÓ���R�:
B�N�Io�uQ�B�Pm��!ahM�25��=�x�!M��e�[W��+i������ԁ`A���,6�4N �w�kjj>:�� �a�����+� 4�P��յ���*�Q���ĴT2:���bY�.rQ �6�U��ZGQ�[�ʕ"�S���\1z�X�\���y$u�&P�d���Vӻ��=�b�4�N]d=�O<+Ȍ/]���z>��pc�x��f��m�#�+��o��)��rJ>��#y7Hl��2���h�ul�Tp{�'&͸�G�D޾};}��?�S�c��fϊ�E�Y8m�9�Ҩi�9\6���|G�0s�Ν<%g������G�2#�>;�� r�3q�ʺ.�z�sKl1��T��J�#�fx�m�~]	�/�L
8�.^�4r��hG�8�t"��_�d���Y|Eʳs��S�p�t<�9>x�c}Tc�=�䨣�P�^�\ ��_����ء+%��\��- ����_��l��Q�ƀK6��g��~>��G��ބ� ��P��-v%$r64xrQ��5�.���Z��h6��\�v��h���Sw��(��Fݦ�N�؂�B½V\��Ulb7/:�k/Ȍ�1��H���g������`iC23�V���կϰ ^oF��z�����p�e-��Y�gؗ�"�F��������s��,�n�mq ����+4a��sT%�����lîc����OV���>�E���Al8Ϙk<\W@s���Z�8�����f��IfIyA)�V��z0T�[�t���v�_����5_���!Y|F=74�B���*���p�ӄ�V����� !C���,>��;7ų�n�SyN8�e�����9y9@(8�4���|Զ7� ���D��[o�%)F�w^tN�j�î�+l��{����5dMm~��M��6���_})0�����O�Q�S����n| �K��pKT@�y�`��=�#�@s3rMi|\��M!��yGHF(e�;Q���L��5	�O@��
��0�����*�dQ@�sm����4�\�F$�{夡6ܙp>�R�9u5�}$����n�_q�<�Lwp�p��[�|�nw�P���J�<�M�!�
!����_̓�&QT�\��b��V��˗�uά�9����S��A*�� �<z9�fB�Q7l>�￿kq[lne��끷ű���\��i�nnaV짨I�MAxx1���������< �,6 o��8 ��iN�����ذ����9��@��I,8'���ӄ�,�`��L|�!�0��9+g��F$3Ȣ�{s�AW)y�%���a'pל�Ш���CM�s&� 5L����pN������:xF�)e�Lz)2H!�"\E�v������M��V�}�����l�5i��$�a9*�3�(?xV6������J3�õ<��ϼ�S�b�|'6�N0��q���>�Nw��w���m|n"���S�J�OvD��CR��	2����)���ka�ƮRl��hNӂ�0	���3 �BC6�����8\Y�$Z¨�)yeS�W&�A9�,��O1��O(^y����CѕK*[���m$��ƖlB*���=UF�j�B�2��a�p�Y�K��Ǌ4�Z�4MtE�Fk3��I��@�S�=�|=��\�������]��Fog5;��r���-1����;���T�V�|���4&'|��׊�����K��\c� 3�j�FGS^���%࣏>��������˗ӭ�7�� �$F@-���
Y�N�a��$_8�L�E8a��o����%���Q���g8��AC];��Dס��g�l����kb���n�e|��\�W*��������F�Օg(ї�h) �!�:��XF�i�/�a�W�H΄o��/�g�qd{UרENlہp���i���t�6����8}괌�][lN�@��S����O�ܧ�����<���٧Ϝ��l�)_\^Կ��k���u�%ZX2�~*��u2��28 Yp�S؆v�i�u�{�^z`�|��$kJ��]`���,����^l?������A	�_�w�*M��_&Uf�Y�HKӼ���Q/CS�����Wp���B� ~(�\��6�����v�*r�KRLZ���x@�\`N&�[0/��Ġ^������Цw�!�lC�<��`S�ښI�sO���q�,�-�In����l��^��io�-�rI�,���q��p�1�LBm��	CC�?��(�Q���Ι�C�J8+Q�b�(*k�R���x:H���tq���2Q:�A��#H�nv��т?~%�����=y�Q��|ԓ'��EqMM��ĺ��Ǥ��d�m��g�ׄ}��{:��m�Q��s�E�UR���L��]�/�	ʪΌ4��i�(<<(�S��ɷn�*&z�||��>�"�^�ԍH��{!���Ɔ8��>��)�GJm&0� Ţ�Kn�I+�c���e��A�ΐ8��^*�V��}���IH���h��(bG�H��&N~�SP�i��Rx�h&N%S7�}� �{	��yz�I��腖	��M��c���Ę�i�4�qTy����W����M���g��R}���pz�T���f�i���E'}���-[�b�!'�N���Ot�y���g[u��Բ��O�Q*��E
��{꼧���W��eXII0��o�������8��@}CI�!c�LTj�[���~�YL�?��ʩ�H��h��Nز6���2*��{�u�,\FU<Q��������cӽz8�Y����N�8!|M��	q�o��`U�
s�e7}����0$ �Dzp1�"�ܖ
a�Ο?��;?#��+A��J]�$&��ht\dj/�*t{�n$�,��-Er�����+ޒ�ͣ���l®���4��'�H�d�Nbc�Q�׾�N��@�sUH�d�K�*c㼯pd���'-õ��&�:�y�h����}w��*�m��������Iơ�(����p2L��P_�0j���@\�ԑ.!�駟�k׮�������X	C�$qp� $������7n(�ŽxHUjq&�A~8H�K�<0����}�$����H�����`�3�g��DGӜWW�<|���"?y�4�r�< ��T�6�~~��w��5PϷ���p��������ZGs8����7������$���>(^�G�C�J��-��հ'+�8J�|/cL�x�13�M��g�#���ykK�|��D���� Di���ϖ�x�7���&�R&��-��[�)ԀJM�Yr	��
h.)��V���$*�'�h�8m�NhE�g�xF�9�K�bC��d/��M���0i�(��Ln#\my�\ڧ�ȹՄӴ�#��{J��c�6����[�	��?�$�k�����	�-F�S�s}P�ۍq|�1�����k��7�rZ8x:�q��`:mۊA�P[���f��j1�7�dL�6�7�!��0T�3�Ϥ��%c�r��Y�!ۓ���s��y�vٔw.]�b�d4H|�d� *����9����7�o$�T�5��$Į<}�l�q�1ب$�M8q���d������I���\��W�H��$����_}-��
�Z;���`?�"�K�R�+��I�������D�S�CB�Y���W_}��L�9�EP��-\QT�Z�#[�=�X���sF��G7�M�io���M��p|]+�� �ǵ�Niׄ��/J�����3ʯD-87r&M���GJ"t(�G��7�^Hu����,<�|of�cPc�Q��nJ����&�Py���85�e3�Xd
~��_�yv��7|a��첻�[�t%q��=  '${0|�����F��'��!,h^�Mpv8gt�c#�z��[����'��d���ϊ8h/�����i�?�X*��o�}��ܠ�z�+�:y���$�H*����䑷G��:N���I�;�M��A�Q�>��]�!$���}|\]�N�7������K:�>�e�PK��|-@��bF:��&#|���3��Y3"�*v�UF�~`�pH8��l�`K�ௗ�މ�=T3��өre,^�w&`W�\��RWo9c�!,)��PY��}^�#[�S]yQ�#ܜ��$aH%7�^e�	9A����O{ܺs[z��YU������@A���=�e�sɕ�9/G��=�&Q�$}��>���؋�<���-�Z����r�9�˵X����͝���W�"U�O�6ւX<HR�,��J>��<�=�{��.ƾ 6��Q��?��2�B�-�/I���v4o޺^лR��P�*�x=nZ�Ň�4p`.�͛7�J*w��K�Y 6M���7��I��2�p���Q�Eu��SfՌ2^؋y���D�:�qVS����9�$A��3�k���L�cF(r��0����1�H--֜&�ʅ0R��Au�6ɕ�}����T0�������ϻ�+i�1�0��W�*�4C��K{&�e��
<�=B��c�=�^� D�C����>}�Lj��L�dʧ<{����&7b0���Q���h�ʌ�D��=|�H�#�O��{Y>pP�N*���� G��g'wռ;�.3�3�?�Uڞ��<��'�\9tPD0�·Mc8��8&����ܿ\��=a����س����8r�qv�/k�d���sX��U�6X���c�%&��2YT;�I0|/^T�N#�ۙ�H������s��9)Q��bE�*�t�T^��M����%O%mEFU�מ$$���#?��BЉ}��f��a��DANC6�"��!Ӏ���#u�!�-\6#WEmO��?q�-Ҫ����iDKH��)�Kl6�����(���W��2i�ِnEW�t����~�=n&y$)�M��6cU�AI��&��d<�-{���{�h��Ұ-�V��������!��qc!s��թmw����tR���s݌3��us}|0��@D���5�ϙ���k��D�,����#4+�Ÿ9����YR
��N,��k9}�y�pmlEn���#��r��!{��i4�{������	��F{0	��D���E�(��z j$�� v�	��~��N�,C٨EI�l�1�i�+c_��'��a�����.��X�qPo���g$5�`����T��p:����6#M��U˚�'u=N<P���;�R}I������u���A��盌�`s'H�G���&���y�̞Qt�z�4P'��kE�ή�Du���O>�D�AFU|�0����]\��,��Z�u�BF� ��-.�t�q��kZ����w@9OWoؕ>'AH��<[�f���"���C �P��h23�˝-ԼzZ�+��{���1�}9,@��r�K�s7�fP�;����A��Ov@�Ī	W6�R ���ے���=�u`.�<'=��vv>It$~��۷�Ҍd�	�N�����;�	/�F�z[1��A����Kj6�+-����IWQ{����pG9�
֎�Ho�H�����%K���[��U��-�A�f��س��^�!GG.I=sz�Nm�(��N3(̠h���.J�)�d�ƙMf�p��A�nn��N��&R��zSS�������M�Un�����%R�����U�͹����,<���==7���cE-��:���%5Iˤ�<��Y������2�����k������ٴjt�ζ�!v��՚>��|f'�Ae�h��DѠ]�X��̅d;���q�s�ޚ�]�M۶�NfyDk�I�'��c9X�����%zq2����H���c|d� ���u
���AT,*m]*XӼz6TJA�膌h׉W��9O��Ls�Y���7W�Sbt!I7�0l�w�'��}�⹂=R���!9.�'���8IO�7�fA�r�I� h��Ӿ�!�S�Tb��u�+�+�9�l��p��-Nx֑��S�J�ãv�|M��J�J)�h�X�q.��۽�\�0mǹ��s�[�h)���a��TI��]D�<uVL��*Αr�z�L���E�p�}m
=w� ���'e�H���Il��k{HM�����њ��q��`���~c��r�X�x8!It�����+Z ��b�9Y}�'+����!e�<PʝQ��X��*��=F�"��WH��?4�z��	�ؿF�9`�WK�JJ~j����uD%UN^,��a@��5�ɬ7HKƛ�f�Pq�R�頨�n0�B]?�l�%��n�u�'#̀b��q-��ی��N3��q���
�[�)l�5�ǌ+A)]��@Z����jFZ�� x��H�l���ٵp��z:����Y�B8_��E����Ɓ��l����gz�'R첳���"v��E|Y~�X�a�F#��Pp�&�O�zm]�{����H7�w�u1�ǜ�N_���q�`&#Y��C2(
)7�t nc�"s���k���U與8�|q�4��t:F]L� �L���;�v{˯I G���`�ݟ���\��<[Nڐ�����IA�V��|gFp1����h4~b�(��.�y{�zrrXA+T��jg(��H�H�:�d��=�sz(b$O;���Dj��xcS�#�� �R*7�"aWp)9�dQՏa��4����q.���h
�!��7�p� }V��쑰lI�R�x��$��) }"OhE����KA���=�I�0��M�G���8���B;�֋��f�2�]��Jo���/��o�ԋ�\Rb_�-i��FHDA%��N���S�\��t��a�r�����M�ίB�G٘k�|�4�������"Lm�H^^����Zz����5�*��X��u�.�S0):[{�|i^�L�G�niaob��k�6?��Tw8/
�K�ǳb?P����ic[�A��s[�j#�: �j�������H������.ʾá-*��x�Ç'rMِL��8�Uu��U`f�>x���y<3'���������;�4?�@�4`&R���͠����sH�A'x���i�R�B�t2�Y��C�)`����L{�v1�̳�I�4�v��*�y5q.8d��gL�7���ćy��+y��K��h�������Y�.^L����n_��>���ͫ&�)AE�h,>7��s�����͐��V��I\ޏ�˜��{�~��m�PrL( LSR����O� ���@mSD�����.3��N��c��h5�p�=sN��i����`e�]����[�YKE�}VS��ozo�
F*6Ա7}B,���Ey�ė��\����)$�]%V�xs��((�T	��֑�==�&6�Oj�t¼'$mqeQ@�ۦwŨ`�G�9�kN��/��f �X��ex�:��<�Y\|O|��=}&I�K��Q�]�}r�=sr�%�j�]q��Ncc�~��Ps�j��ŷ.:�M �1�d	��<�X�
e�xn����3R[RW�Z�{�&0G��C��t��Yi��3'I��if�p��f���0N���~��t@�"6�l��5����� sJ��s����d~�{�︱�2�S�^Q5N%�+N�(�l�޽򮮅Z:q��e�/ⴡ�H$��	@�������pb� 
h�3 bNx��'�\9�E -�ݲ6��ao8��z��N�s���`�-
EM}*��0@�۷n�4�|��J�q����~��󵪁�S :|�<D�l�}��]�0�nbG���G������3X��G��z��zˣ�I�y㺻�A|������n�=�z��{���O�M�ͷ_�+�^ѽ<y���ܩ�(-��%���8/[w��!	q�
dC�\27���ި�
������>Nb7◮�i���>����O~�S�����=��U�Gt6}��_���rp[�#�7gt<�Bb�?�G)��L����%�(N�5�i�x�â��B��u�E��&:)�4�&ɦ ֙� ��93c����>�  a,� �5��5!��8帹)��yr��ٵq>nݺ)!'euEBG.������[�\�e��^0�9fm��"R���ꪬb;J����q6F�ZH�S����8"O�!��J����B�O�{](7�w:=ى��C�ҽ����0��,0^��̙�EC�L�zEF8��E���wGa�Vp���G�H�G��L|��Lr��zk*ե@����;qx-A*����Δ�$�*6j-=�F"ٵJ�o�����=��C���)ӷ������溛���YI�͢^z�L��a����&w�.�f�u�f�O|���7�ҳ9�L�����'�n{&)�a ��h�}!�.)s����$)�m:�/)�^�9��p1�`N�&�Ta�Q�J��8B��5}��HjlS{]ѐ�L�h��������G|`��%�i[q��9�rsџ�ڕ=2U�]ٍfUx��l4�쫬�rZՒ�:�֞��b_`�y��x�����Q��	5�#I֗.�Kё76�@�o�9 lN7�#]n脲PM���J� ���.���p�����,"��o������?ӂ	Nc38ul�3�J��&�--4^Yb�-�a�@�����ƍ�z^�[�BR�s�"Ђ��¯mx�홝|l���@���'��x%�}�k'�7�F�BP�4z�S7�:6*�kBL��gQ4� .óHѩ���R/T9�D�ݖt���, ?O��r{�7*w�N[l�W�:R+������ը���ن�l�wD-��'�r/9������6��+a���qo�(���K��?ԏ{�ɟL�l�����辰aK������F�ðc�p[�?R����_UczCVY���kt%x���L�K--B��߸�>���鬸�2��(R3?�E#��c���˺6�1�ln��x�|�;<�y�Ҩ7Tʪ�+�*.M"����*�jѻ�*���s��U)��x���1h�����
Olg{���;;y'�e4��}T?��%'w&>��L�h����F$�\��OJ��K�>�U1��y}$	)Y��$����S|B�ѣ�1-����^U����G͜S�k�I1����yGۋ�/�@��%K�Z❸îEƕH��+��]}O�� �RT��{0�>�%�A�Aoee&������� ���g��箭y�C���f#��.TtNC�{�M���N-V���H�hxv<u�k�S��M�0�\4GTm!2l�D��m���.X,�_�&M�� �Q��u��6��u����E ��M��o�oJz�,�p6Ժ��%���ۗ�m�{�:k�*=�=v��/�-7�,�;w�9.�%���!�]��eù#ힹ���c>

g��wO(�N�D�gA]5͢M�����|'�r���-����h;�j8�TJ1!��p�|N|͙����2�\�&1�Hp3}���j2�:h' Fkl�=4Q7i�<_�Bՠ&�]=z�D�������m��PO����ay���$�u�㫯�V2��l���)�<�uX`��N��.�u��6������=�3�zMν�>|"}���ҵ��ub����*ZG͑�%{ґ�*�5�l��pb�;K��fy#�HF�M����8�}��M��3��y�JӒ�,ۻ2T��T��pЇ豦ւyuJ����Z��*�M ^���m�����0>�vqiA���9�O���C��C}.Xvhg��o ;f�w�����Vb��؁b�ٗ������ٰ5��~�$���u�p�p��#l��ZÜz��º!,>�\8!��:4M�����(ƃ�#p�IKωs)�M+k(�^��]�~CN݃���.�*�O�)�v��Q/]�f�͑#A��?tu��S��͡�Q,^N�Q8R��$��r����s�`����;õ���|�i�%<)�(:c�r�P.��h̉���\�oW����\v4�6A�-�>�r�lr�~gr�p{�`���,�O�\�4�_X���@��;����"2W���s.�O���3�泧�I�>t����Q$���m{�RH����J�Ϛ�����N�f6[��}Y�'д�`�_��xdK-msJ���'[�����A6�"�B"�xUcf�`��F�BO����Ltt��w��U���.�iő��7�B�J�������4�-eK9��!s� 7N)���
�0e��x>�\���ǜq�(.)RE���	'?�T�8�,�� -�n"ej2]]�g�;�-�;��`�0��35)X�3Sρ��x��l؜B��E%̓3C]ELwͦ�� w�U���� �If� 4�0Q�<h���ްWl@v��AP�7�� ����~����KaT�Z��7'���(�v��Y��q�b4��E�OY��ثgl�n�(N�g��'�[��A�6	 u�Be�k���a�.��R���*�*(�_�	ł��x�'�������zŖ�
�����}�88��XjJ��^�~�3�M��o���W4"8���b2���7��?�R�T�Q%�������L��5a|`Q2�.��p�*!@���q������I�;ܼn�k��M�S	�[�+rd��@��0�-_�A�ƒQ��,^�w��ݘY��x|����	!4���K�Еv}<,��8�^*��1|���A���|6�U�*�ٸ�{��m������S'��6o��UL��e�i>JH87C����,*A_'X��dj��~WYZ��)b�) �n�H��9�]k˂�{z=Ɩ�D��\�.���`wg]��S+�ή����e�1[k�Y3u�Zi~�I���g�@�0�:�4��{R�f�._9+��> �>�Z�i{nj-�U�
��+�7Ri;=�K��a�X#��"9a�~[�Z��ڽq\I3��x�l/�i��N��آ9:�o\s������uB�{1k��$���ܢ�#�K=a��'��yb�6�A�9,�apW1jl�����NH��cS��&���`Sh��X�cKi��R������뼺�������?��ȝ�=1��f��������93���}�5sR��J�J��}vG_�
�������gϜM�N[ƺJK����[R��ϊ:�nB���ك�w54rcmC�Ña@>g%یlC�9pa���
���ć���gC����(ꉈwu�ג@��B�:��tz���\B~$ے"w����,>��jp��z�o��Z����Pr>�,w�4��QO��Lh��w��5l#�7��8���	f��z�����G���~l�n��r��ܻ�@���˞	ʊ98&5uG%m0]�+�R���ͺ�<���߈Ld&B��{����eG��:���E7j�N_7������L��������|H���U����D���aqG�z��ё�؆���������\����?M_��$���w�}cj���X�#���~�D�.��u�f��m��8�����W���k�Ν[ⅼl��<%G��[n����3� ��onx����n�ϝ�%}�888#[��Z���`
p\v��i�J�k%����r
P0��vѻ��QaޤinaIFV����"��u��F쵽ae8��W�;�-"հ���#�-/_>W �ꀱ�������_�E���_�B����<�ٵ5���E=���׾5�q1�_����N?�u�:���j���`�q���XҨ��>�D5�e����Z��k��ܷ�����&���TQ�Kʮ9@lQ�O!R�Ӆ��N��uv��zUWz���<�"!	C�����1�N��I�����|I�G�������*N��v�;1��n�A� @h�hIw��d����yϽ��o�@���^{��z�:�:6�WD�3GeW���U�s���Ā�fr�b3"��b�^aӣ��$�MR���(���g�&�"j<3<�3g�v۔c����j�6�yR�+<�Υ��	��|��O��Y`��YW�w6���j*�$�;��I��vv��_����=�D^�yM bcv�7�hw-/i�P5�[�_�Jr��B:~�pV������ޅ��&1ʎ�6�K�HN�8 5��ڇ��lKww��6$H�T%pf:v�ί�p�uGjwy{�Z���T��8��$¾qsU2,�ѧj�Z;]�.,�0$|F�i6��� ��g�B�t�2�`��Y�,vs��N���qz�_~�g �q�e-��Ӵ��>��gA�97w�׳��y�������y1��ܓ��#8���C��Ս���M���/�������ͣ�j��
����^V���9�j�)/�ڇ�^L��F���r��O����V�\ͻ�Γ/�#v����'l�����&8�{��T.����/2��q|yv�UMZ��gtJh!f�V��Dh#�pF���8���9i#�Ct|������@P���I	���H��>I�!)��j>����_��<!f����=��8���z8����i�F� �be�J:��yU�Q?ۂ�������B���׾����L��~=}��SЈ�D ֳM�ti:�Q����QƩ( �ȁ���5�Y�i}�Mo����8�e5��d7��X��>R���˧_��O�����47����h�d��G���Sgi�������O��"kk�ɧ.���y��x��x!��=�#Yj�=�=�����N��ޗ�Ȣf�nfv>]�b8cN�h�N�A_I_�U���C�n���g�C�<�^�7��߼b�7?��lW�dU�o��Bz񥗅3���c"E�����~>TR�̙^z5;�<��1\l�4o���y�[x垍>rUe#Л��Z��P&6��EG�ƃ�aB��M�FXv�J��s1��撒5����$.�����4U�L11��ӿ˺wWF�, ����/��s�U:n����N���sMW8�7sI#�j A�%��q��^d6V�n��\�G��=��^^��,�粇DPz+{I���W��@�04����)�HT>�϶e#�Hfs��E	'pT������蠍�i�;iK^��+J#�.�4�������~�b��koO^	C�)aC�;�.���5'�1�O��[�P)��^oC� 3.bY���v&�]�TL�.l?�P��3O>����~�wrq��&!������H��vs�����9#T��xO������0Y"^�[��I ]C�pR#�/_KG����_��r)�����9sS��ЧN��w���G�B��eݺ�f�X��65ǫ-�)�,+T~�(�ې�2��3&e�����Q��4M`v�jP�^��{4��R�^`� �*��&j+�2�!O����s �D��f0Ⱦc��)���I|����[�;]^^4���'r���E�"���-�0���t4�Q9B���~�����.%���sS&��7�j�����O����*=��/������\�ҡEC��?pi]H���z:u�Io~5����yeg�ֽ5�S	��S�!�3�^V��)Z& �Q*~�H��?� Oi1��j@q^HJ�h�Ե,��`]L�Jm��7U�[�NU�S9\���o*�� w��i��t3���x�ߧ鹑�'F�7�C���a� m��ż�d �e��X�[�֕��]��"�
�w�y/=���g��m��mar-a�������'�Ns�3Ug�aM��Q��O#�Q��~;SE�]ؐ�(&��?��ڲMcF�q��G�t��~�ݬh�ٮ��>�(����8M�X�����Tvq��]��(u��ϟ�|](4|�~�����-#�4�z��k����.�3�y\�+xoY�N}��X'.fնF���|��(�4����8�	*���ګ����A��h�z�����X(�-��~��kJ����tV��}�s�^*����L��a�ޒ'�ĺ�
�e�x��T��@=���Ta�qkm�-b��7^��x�,*�5�f�呤M��ThSQQ���:I���X���M�s����度�q��.�_I���w���)��/|!=��s2�����t������i�}��i&K����WY�}�z����d��I#N8�7���\��!�r`�v ֙��~);����';	��{�=~�l)93b�	����]�� it��a&�^�n�Z'��S��mDd{�
�߆D
�&>�����8|��^<ʧ���ZH��}���=PT[��՗6�~���=LEm����Ϟ��AR��H�A�y��SD�z����hޟ=1�}�w��_����a)�T��B������Uf��=G����y��ϪB�d3�ŗ~�N��ռ��]z��3�<v�f`��#�s$>*�m��dUF��>w��f*k�\e���/�o���n��+�p�b�0�
���G?65u����!4@��1���qSJx9t�]G�����D>)Y��L�$5�����#��M���֙��4S�Uռ���ڣG�9:*�|��9�;�~���4(x�1�q���u�y�]vd�$5o���{l�/��2E�މ{�DI�5��_������U�vm*61��#����'*
��� ��Y�} 盳c�{Y�?!)���&��b"���pY[ۛ ��.�/������cGus��^U)�:�^�b�i��ܝ~%K]gbR�-�9O4���h�v>X�*�t�ұ{�W.�s+��o��N昨7Tj��/}%}��ǔ&���}/��ץ"���re�����jD��Le^��d���Dpԣ~��\��WO���� 1��⛢��ů�9}�U���ݪP�\� ��S"ٔ�{�[���7�-)%o��$SSm����ʨw��JZS[qR�UN
�}��4��,b�q�p{�>掜.*��Q�������`xj�Ȗ��f��q'!�d���b�X�dSi�/�߭Z�I��:��x7��ގ�0��~,���_~Y��g.2�.4����n�����CF ����R�b�qG�<�j���>�	q��m�8�+�ӵ�g�r�
��|�.y�F�14�n<VZ7f�$��w�&�T^95z�Pl��b[�����$4CU��z~��r`@e\��u39�/�4>��u�0k�8xSw�$A!�\���I'�\��*leWui��E!������K�G�c�*����n�-�΢2��i�fO��l��)�./l(ǅ�ԔAh9�9�ٹ�#�v�َ�)_�j�;Wx�|_���Y4"kl�~��l���FNO�`������i���k��3x:� Q5�،��-k�%Ŭ�����ݫڸ='D�Q�����W��=�|�sOʆ\�|U����P�o��N��#�K�K�Ig3ϼ������)�| ʅ�=���UU�rJJ"ٽ�~��AJ{��i�:ɿ�����;ޥ�W%���,d���OF���t�׷$�ׯh��k ԰��^5M4FKE��mF=() �n;	�zn�v�a�9О�J�߶aZ�
l�J�1O�o�9M�-H'�Ŝ��y�>�`z�D���N���p���ƠF�O�,My�IWЯRBnH��׽o-h�K��j��f
�Y�o
�j��RE����Moբ�tͥ|�.X�:�.��H�`�w����裏+��^���
g3q�� ��Z���~Q�}��׾�I �!˻fʾ�P9�,�Z}��d���B^��^5r��t]� T�Zȼ���;�v�,��|(�������kO��占��`���Ni(�KW���J�S�d��69��@��l��|���pY$pZ��Ͽ�m�?�3o��BvC6ϲ9�sם�"5��0��ݔ�1�0P#F���<���a�T׳*k; J<?����!��4f
�<C��v�H�g�䝷n'�2�B���A�/�Ҷ�|]YǑ������ZבGj�l~��GU�?����H/H���Y���彲Pl��mt�����/9G�O�gdcs����B��1?���2H�fm�aVm���� Z-������=;=�S�����/�g��S	�M���Oq�(���f�ī�&���4
=Ć�?C��0���X3����+�k<��y'��B�ǔ��Y����:��)`��d N'����T����Ϳ�=^z�e�| Ck�j��:�=ɽAٓ;�MY^X�����g9ZV�s��PCaTϠ�O=������H� �Vl�Z��f���q�Q&g�eCٌ�����i�қ�G�Yx'� ^&�Fj4xo�֨T��=vyI 1q���r�*�ɕ�=L�9 ?G���B�ڸ;�09)�I�&@e��$�2w�qb,*v�jH}p]x߱+����|⊶AhhJ���	<*6���7��y8g��,��,t
�vr2;ׯd�.c*=�������埾�^y�%B1�$;������.\�y~�l�3����<&p7v� ����D2��!����YqH�YP�k����(���rhӇM
Q�|ĈɄ�]�y�\��@��>D�⯽qC:<�.�ay�I]�{qʈ�I^�5��Og���̌b�(-hH�^���v�;48��=��x�sUS�:�F���5�SD��.?��C�mP�T� L�/��^�ɋ�^)�'���2�P�L�q���o�� ,y�9em��EU�u��HB`b�P�˱Aw/+U�E����Դ��#�l+�����'c���[��	Ժ�f��H��!��3�9h��^!]o���L�Y��Ii���x�8w���g�{��� T-������6niW������;꺑oh�n��	i��o}K(j�4j�h4��&�n�!�-`�N�|@�TЙd3x {S�k�s4:ن��7�V�OV�8c��;>!q@H��+�ӱ�1�;��.ZvI�`��=��}+m�E^��ZZ�N�0؄Xd^,��䯺=������`�/Xֹ%�L���e �)���1��Z���$�>6�nB��axE���hW�^J�m�@ǽ�����\p�=u�1�Aj� @���/n�r~6�V
��%C)"�8=��h�+)3��r�-�a�|�g-W��f��p}V*�159m�]N�w��D��XHp�4�QqY�j�4/E�"�G��͢'��Ǣ�^������5Eg���9�G�BO6Ӈ�SC ���B$58�W�ʍfK�U��F�K���x��z8obKe`ZӠP�𞬹f��N��=��x^~f7�sg�B#pF�yB���+����%�Y�|�9F����Dvw��8d�2"_"Y�HS�)7�6l�4B�͋A�#h��G��E���X*��KblqyH�kH�2[6o:�<
E��9eؒ�I9�&��7��nN�~Z�&>�J�����VxW�5�H����8ZvEńK|A�"*È������� �VF8������r�����MK���0�6ڷQ�Ua*�n��ڏ�6��ٙY��XW>��]G�:/�=����J��&x6�����5���=r�Ps�($	�ـ�ѓZ�MԼ��u�8R
��vD�m�`� �������Ԇ�a����c�2��'��3�{mH��`"l�����9;����]�Pޟm�ة�u���M��8x�\�`XP�AO6����~��RgY9!�RD�N�g�*�Wm����j�ɟ)p�$�H�е\A�st�H��'��G?91���7+ra���-��M� J���:�5���&�8+v� </:Ɣ�A����3K�%ӳ&\�J�lZ���q�)~���jT%�j��i:$yI����YJp��ά�DhM�������3s�)�6�c�`q�����Os�@��E�&�G�jZ����<��fvcNhH�ɓ�˰��*�<'�FT�f]�m���$���M�hbC����V�B`|):q�5�"���̾ʞ�z�,�.���bhQY��2�]̟a4��"�߳����V�΋$f�w@^��2���Y��p��~v��H�_`f
em*�����@C�m�[���h��,�V��� �L΁��0�&$�N�K�b`�B��c�t���i2�"�)�(𫨟�H�a#�.y6�
���A�r��T3/�u��U���CRK��ˆqM#X+}N�ا��@:���Re|�~ޑ��G���|����暢n��Ն��R�\s�h���+��(�7?�8�?D�Gr,F?��O����ny�'/�OG��"���	H�䭿�
�m�[��RO��s�}\�=��]^8ҹ6Eƺl��,yF�.F2QO�W�uwRܤ�A��Rxnj�(G2� "yIlX�b =��m����6]���ިf�X��^E"��r�tgR@�M]G�F�fÏ���6،g���I�jW�=T�R6X ��l�/���ᗻ������z��8��k��U��d�����߉�Qa�`��uv���q[���U�r���/О��2�����3�= ?}�דtF��ɓ3>�}���<ڔm��1ݟl )N"��1�� c~���v%8m�!�PBa{�7l��h��#�r�k� 5V�j��n�����]�H��؄�9�$�#O�������u��!� �G��f��t$�S�����G�x��wk-��fH�+��{�%<��M��2���Άp��C���B�zF�P)�!�����o�a�_��O�%�Ϟ���HF��sx����C��w�dh6J�{�r{+��2fd7>9����Ʋ�+ҙ���H�eQ09cҊ����h�����x2_�$�tPU�S�\^<K��hs#=c|v�`z�}�jq�M���^�~F�A�8p/rʐx�������������kZ��Y�zW���R#���C��0��R��k�G��kC�l�ۣ��Ȯ=�F��]T9#�5P��ZbQ�,\�ʎ�:��r�����Rk���q�gZ���-��^5��^����q�:�%�+G����}A-�߀&$��n�[�1����{�/�������H]�N���i{e;�fg{ۇ�,9�_�����$aC�sJ��w��7R:�MZ ;�0��?�6;~�� �^���N�e��֋qRa�wސ���L�p4�#m�׉i;{�����lז5R1�PsG��|�i�jzvZ�\i�6E�eۻTA��mv���2�� �Ɵ4��F�Pc8!���*J&�ŽAHb�����j�80v,���|JN�_�g���-E�s��?�0b4�k�>&�SD2�� �����a��H8mB�4uBj��٨��	����:gb�Դ���v�Mmm���T�L��\Aw�)X��Ń�M+, �o`�\7T_ ���t�
XP�A؛��XR渭!/NXF C����`pJ��k$�</�b���mm2]�l����~���u	{p]���qb�F4#{0ǰ�)Ù�y���N�6�������0fsɓ�l�@/V���U�g�"J4NOI��߶��ㆴᚢf�|���]��!�N���]�|���m��m�!=\�"��]V��m�NnF'�2<�)|W���QU,<)���^��(����]��J�	@��iTjSj���*>9;�T%��C#�4/p���H���g��@ᡞɼ1�*�S�4,������SY�ƖCj���F`{����%�� �3�z8�[cG+L�Mb�/h<�$QAc�[�sy�I�@߭&.cw�7t⢮��1X$5d:�P�/OS��R�X}#b���r��k��6��p?5d��M���m��"?�F6h�77�U5�S�)A�o ��B������M>�p��s]�2�Ե���,d 1X��򉊋�ρ��mJ�)��V���I����э����u�^��7�?t�yf�P��Y(����=�.��,���g�����Ą�
+v-G�R�������2Ww0��}��mh��*zYļ�&�:�w�����Ĝv�4��(��76o{�J�܏MA��ݽm��zR�M	M*�]bRji��a��#�O��tBJ����p���w81YD"nz;4��$��;�_0�5��}%��;Ө얌�
NM�;jE�n�Ԉ��q��iP��h�f~�E��h���X����q�7��q�Q"j6�R2�{��֟���>�J*��(�-���7���fώ�D�2L�/F[�~ii!V��3ڀ8Q�����; =�i����Мu4"g��`�����-�~�
^ר��(\�CΗk���"U���������ѭ;�j����CQ�hZ�ں��(V���=�Th6��Q�F���3�9{����5v����E"�]�q�+�o��|%�g�i�z6�@G�|���$w�m&��?yD���Ysx�
���j=r��qvAً�A�n�M�Pgv���6���d��r*f�#u�(0�$٘ �]��5/����C�瓺z��`�G��īa}v7z7*#��mx����Wll7d��t^��f��� ���5��>{2�l� $5��Q��IMQc�T%.,%6��m�0VVAd�9�J��L���y�}�A�Z�ъ�4:ޡ��60IX��<<��0�D6I;Udf"륂�p�	x��wD��i�Y�PC��l��4(m�ٛB��(8�H�؛� �2����I��֝;%�6������ AW���7מ��d8�sb�i8�W� rL�vNK�;����"p�5����坔���G?�sh ���մriE�+6�g��Ϥ�Fz/M:%@�W���F���}A�#�{ާ^:H��S_ �G�p�����Q}X6Ed�RCVGfXD6���,іt{]�skÈk���4�&�f�$6A6e��}�9�p�2�g����F��m7��eH^�)����*[�n�I	h$:V5�s]�ɚa7x�M߁�
���)���6�Z��mf3=��#:�*ߪU���R6cR'��Qw^�9���c���T�4&>��Ӣ�
|��<��s��T��[�[��>��+�!�H��w��Б�������C���o����&��Jc���
9襉�ImK2��/�inn�G�N�ԅl5:�	�\���Q*�?����*Y8�lR|�g��4�ܚ7y~�IYfc�\�w|��Al��?��z��U��u�$�ϘX��ߍ����n�"��U�$��c�[ؓhn��mڼ�Kl��0D�����mw5��b�^�ͫ�D��ZP
��.m+�ܑ�P��n��k�+����$�*f��1r5��w=5�Q;B��>�j=սMM�"�ü~�w�pqEj�����G�e��b����6��ʠ���U��Ơ�j�����j��8	�&�T� �������0u�'=��ea���ţ̽ex0s; >J�I�|���Ȣ#}e2����-��t�X�FUb.�/�ܪ��Os�g�G����R�+(���Y�mM�1N�N'�� �N��G'�'J����L��j=�ZU��}�i�P��.74&�8�=��� m�?�� ��D�x� ��7��h����NvÆ�t"-���܋Z�f�*�!��Ѡ7*��RY��{5�JuD�Px� �o�QGWKj��Г�����R�]-*�\�Fs���5Yh�J(�Yi�(�Յ'��>f���!�S�jgcC����g�t�����<\m������u��N���i�Ջj-mûrJP�a\Q���YX�z���z�4jf��:6�1$��5��LN��}��N-��}y��h8:U�J�|�v7�7��v����5(�V%$�~Y��`U�6#�F��چ���i+A�CxN��/��|}y�����,ÊGjO��=yH[��)���s�.b׶���P��In��R�D@f��4*�b�yVbK]���{c�U%��F� �)Oɪ���^��F.�p4V��5������O����_4�0�$c���S��(�e9p���w���[r�q����AE�2L�BW)�8�3n��i9�p�{��嘬����J�t�sD�8"hk�Ɉ���o4���)�jH�X|FN3m؁����ưu+ �b̷�@���/Y��У��W�9%;�='������g���`�H�3P����:�h�z�����j�:X���.���~�F�����*1��Aa��7��
D����da�'��n�2Ζ���>'(R�:�>�.�_}����e���u�O	��������";v�}_3��X���"(i*x��U�+�\�6U����nLG��6��V���,��s���k�/OPJJ�k�y��	��w}6	P	M*ܞYu4l˄��M�{=�_�0Q95^���d�Gs8�^W1�{"Q��ؠW���pb���m;����K^�lVO�mT��S� 8d�m�­�����M�te�v|@�I��'��4��V(���(#�B����"~l�-R�]ؾ}�дwl�d��@.��~7�r��R�%��}a�����Q� �5q6ʱ ׽��>�� �;a��m�>��Z}{�H��	��Uގ��M���u�D��~,��\�E��z�>Xxd�t�Z�G��[�M7£���Hd/���B�4To�P��x7٬�3�z�+$n-iTѸ��pz�9�=TQ����p�tp3�36��Y�n�V��ꧥ�O�Ƒ��@���@��nM��#�"2_��py9PI^�1�a�6
�=����T���o���WPYt�d�ʚ�-}��ʍfur��#�: ���޶׾w��D߽f�2�q�r�cݚ���Z�g����*4w�!w:6w��W 8>���`>9{Y�F=���M��Ƣ��rM=��d�����-b奆#�u8Ђu����+}�B����9p+j�dc�9
�/�Qc٩��:���)�)��� Y�@�8h�Z����"�t*�@��	)*�OQe��i���b��c�7ڕAj�m�q���	�����J���ӕ7��j�o�*�� �f�-qh6ʒo}?��Xr�}Fa]E��N��T��H�X[uO�S�96����*���F��1V��-�B�Z�99ʊ\�fmdT1.8ݮ��r��Sk�#T��oH�����=�(�l'�6ia��wD�mSЌ�!�;FZ����|�,���Y-�F�v��hY#�y6�R��1�6�6$��֤!w6��J�GG��M����&���k檛�6�P)|�`د��P��p$�MsqU�7F̎�u{QZ�T�2��6��~��ؔ8)�&�J�YM�����y��ݪy��UF!g�{PZ;ND�"����
���L�傶��"����@i��yK܅�Hfy49��H���ć�	充��Q �؋�m�����j�T&�~�}��0�SR�)�i��I��G��*�}TD��F2��UU7��{���<�._�,����;h�|�i��&1�J
�{�֌����B�/fy����փ��	�(�Bhz���G���Zt��&��s]@%��C�,��>x:u�T~���P6����>>c�h؎�ߔ�mz����P�����oR���N��'� �5kj�xR���L����=N�	{
�J�T.x=5Q�.�l�a}3R���RޮWO���/�\�ɴ^�V -�~������ee�LIZ)�~��'���q�hd�c�A�	غͨ�Z��>w���~U�K����D����u����mSw]��� ,3ސAe���"�M�k���7&<�ؤHQ���'|R�~�sMj�3ڳ����[�'���2D�$�1��������>���'5[�6�OT��}��X�˚{<��'�==w�cC�߷���pWKF��_�Ro,T}C����lc��=�kۛRu�-����]O�F������~i�}C>�;�!��]~Ԗ��΢��z��5�SW��������7�����t���3��<i�aޯ�M���cI"������̦|䆘�{]�oH��d|���-w9�e��rI�r_4�=x�o�%�鄌b����Z�S��G�3@2�>S�_ڲE��^F�ُ=%��R��z<r�k�X�(�X%�Dc/Ζ��ޯg��'��U������O�mu�;�J�¹���I���*^�c�FUb�Q�޽�>�iS>vC"Zϫ�?�DDa�٨Ƌ4��|;���f�Ft�5�kσ�Q�s�2������L�~�������z�#��q��;0ݿ���|��	i�b�۔E�?�}�anĝ���y�RQ�Oe���[������������8e�����>�l�M5��;]��<������	]1X�Bi�    IEND�B`�PK
     #{dZF�i~�  �  /   images/85e66502-362d-4a26-afcd-97fbc4859675.png�PNG

   IHDR  �  �   �lC   sRGB ���    IDATx^�y�o�U߹�������$��$YÓml����ӡCU�ؖ��bl�iL7Ch��!@H��ҡ����Օ�*����ƃl��,����7�������]l� ���٪�{~g�:{��k�9^�   @ h0���m�i�   @ p^� �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   <TU��tYE����^��}�w!�   @��J�����s�Ҵ�1˒��䞝��_�t)��(���EQ��8veY�eEeU��M��$��yQ����CKK��6�%?�}���v?����|���   �<����}�K���f?�mw����˭V+���]�v��p�i��s��%x%|��4s���E���(��^��q����o<}�ռ����o��+� �W 2@ ��_��[���r��p4��<��N�'q�z�~�eY����n\u���E��(rE��5�k��*��*w.*�8n��[U�$���<�'���Ao����>�W��}K�����K@ �  p@���_�-��o�Uu�sѠ(�YQT�4I�0��W9�+W����]7����v�-�y�$�Ue����$)�$��0.�"^XXpG�������?�.��	 x�|F��   |I��_�g4�LQV��Ey�fi⽲R���\�f��v{.��������q���E��o�����)�Aq�ī������������ر����7��!��K@�b!�   @�/H����O�]W��8]��&ij�Zye�[bZ�\�W1���ή��]9WV�%����%ᬟ��z)���j�+��?�}��C?F5�_Є�s@ �  �	������sQ�3�V۵���b_yA"�G+D
Sp*<�BcUY���=7�\QN��*�g�6x|��g���������������/��g�   <�~�g��ue���v'U%	^��Z)^	� �+W���Gn�?t���%��*��ƉD���UY������i������O,-.��7��۞zN��8!/����! @ x�D�ϟO666������8_�Y��>���O�x>��\��\��-�4���]�WB$�$b%x�vw]�Ԥ�]Y.IcWv�ݨ�q��eY�i��ǎ͏�-��Mo���=g4^�F��;�ۇ   @�Y#���oM��]�g�������J++�[�9�F�ϟW2��t:�{����?�c���'��:�v��z�8��,��r����4sY��7��w��ļ�u�1_���t+��^��Kb7����Ve�����r��v�E�o�c���]�۰�9�   |�Ο?��Z{�E�B�f��|���v#�W�|>���N9���۝͕7r������,͞|������yy��j�ť�:q������ͦ���c��N�m7�繉_��*�-ސ�vX�:M�s�,M��`��xÉ���~�~G�~��@ �@���mok/,LW�i��ҕ���������#��d�L糹sլ��~`^Y[;�@��w�4��iֺt���.J�?�y~c�j�+++i\{x}H��\
e������W�{������!
m�	l���u]�!xzu�.S�n�[�r�/z���G�-�Zs��J.@ �������[�&Y�����;����,�LƓ��S7�F�ao6����Y�n��w���7�tz+��kUU]lg�Ս͍WW.:[�r��vkG����g�4�{+�Z�+��=�ԓ&�����t:���N�c���^>�k�@b�9�����۝��go>��7��/T���}� ��wv�KY�2n�Y̋WN���E�����^\\\*�����gY�&�I����\�����x4�~o�$�t�8�tUV����v��\�ӽ<dۛ�������!��u'p}@ � ��D��ߛ-�^tn<y�x<���h��py\��W]���p4����|��4s�O����;n<�Q�$�����y��Y֊WVV�����ʻ;�͝�f��Ӂ���=��&t�VW��+W���UkPȮޗ�������u4q"�����G��P���O�'O�x���w��k_�ڃ��4���~A^��q{����׍��o~�'��������f����jd|
ש%���-t�uUI��p��I�<����ʭ�rqi!�J�,�r0X�vB��v�p4,v:��u��^w���t��j}���>2��W�vze>ɟ^YY}2I��<o���gS���������@l^�   <	�{�ə���O�:�����[���O�E���4����b����իW-�LUN�V��&әtC)�!�mY�q�jۿWWVܑ��\UQ
AHL���g��w���-,�x<v�V�b|���v:9P$    IDAT� �,�G*[潻����W�D��=s��ͭ�������*yra���ӹZ���v��x�b�WY�<o���'d}<��{�wskkmoo��Ҭ5���Z�&I�U�p8r�N'�9�Y+�]�rcGiQ�&���[\Z,u\_�ݎ�����ڪ���,��,���1#�Q����m�M���T��f��oQ�J������l:�������M/}�ՙ^+++&���tʅ�������Ǐ�g��~���=L[�F����WVv���S��������r��v���ne����Y��?��y>LӢ�nz�����"�����S8o_�`?`n	� �{�ϟ�wv�3���;z�h�e�c�?�x��z$����M�3w��I��[ZZr�/_��]��������q)A<s�<�.q�O��y�&TC��Y�0w�.^t[��nqa�zݎ˲�'��J^e�� �l�
˵+.�Jl�����dmm��G�9��N����s�X���Ӂ^���t �4�İ~oν$.uh�����H�n��EY�Y[}j>�(�>��葅�ړ�Ї�/�����|珟�p��?�r��=�����MA�k;�'�ټ����Ι�i�R�v�]�}�����6�����b)����d:���=7��}��JFVJܪn�l>7a[�2&��d�Y�SQ��N�k���iZ������knuu�mnn�����j����ZeY��.�:u*�Wݓ<�Z�i����c���h����`�O&�X'&��p�ot�`�߳�$z��,�*.}���z d�>�=.{ݞ	q�S�Ntɋܼκv��c݋^�^�T����^Y�f��dF������q��[��tsyiy���+I�&i�'}˹h���o��t#���V+ݟN'�s��R�jR��EQ,�ǎ�>��.T���է?��ꮻ�:��x�y-������'@ �+I���#�N���J����`�8����v'��/ݰ�?t+�+��j��d	��dj�Q�P�C�+W����b)���[_d����|,׬�E+K����{衇,�aia�v��CJ�0��z���Xh��Z����y>��������[��x��)�,��y�/�()#W�
�H�Ԏ;�.�.��\�Ib�9˲T�7L�����uUmggǴױcG.�v�m����~�o��7>o�x^^�����t��zW����p����mi�eY��u�ťXbLVb͋��)�a�H�*�@B�o��ޣՏ��p�9��� ��ܒ�˵u�؛/������$�f���î���rww�l�[n>�cms�b�����>[;��������ŋ�3E��F�$A<�ڶ�|��m����4-�BטO�q�nǭV�&�=h��4I��`�����d<��ՙ�E)�E��_���q^�Y^j=���3l��������ի� ��q�^��N�]����:�{0��u�45�����X���E��w�� b���G���&��/�L�3�3����ask�?v,�\�u_�~�V¹:3�S}?�ά����5�8P�&q,���VҠ"Q����'��L���8��ι�(�v�4fY�RG��h��neq_���v%{eYΒ���&�YUӪ��ը*�$)��h�P��~�·��jg�_--mU�����_�����B�! <D��{o����Ϝ>��˗�������z����z��:�Lb���敥�E��ZN�1�淽=w��	7�L�Q������l�Ξ��u{}?�ƾ�B��n��]�$6��G?j!K��n<�V��U���+��%�� �噕Ksߣ�>�>�яh��G��[�P�2���\�H,�l^��j��+	N�ҿ�$��컍����M���������}����^�����:��ox�w|����ϼ���[�ο�|t�䅤��^�ۍ^2�L���y�W�A��i�;*�x��1w���|}}=�`�v�3�닲��8)KW�Q�>�QF�3�*a&���ֶ��4m�BQ�����ڪ��ԋ+]C/}F-P��RBp4�'TF(&����г#*���ʵ5Ź;��㏧G�������1x��5���WU�T�T�������b�V����G4���s{ �7��Ua�RK�ʴٶB���ʕ+q0p㑭������ʲ�}H��M���<y¶d���IH�c��Z&����3��*P�P��J��mmm;�b��tڱ>�(�r0Xt��[��G��>��������7
�7�?���l�8�@u���o�k�>���@�ϴ(�W}�ղ^~%��{1�5'�q)��i��$I�V�m�{8�b#AL
�`W?�z�� ك^��E��;-�n�e��f�ҖP�Ӗ�N-���R���T�����.ky��#'�Γ$��I:K��*��b�JG�r[�N�ZU�[�Ngc>��D�w{�'ՓD�^���YM�v:�|ҞTyޟo���[����?��-���ב��� �U��c��ϴ_z�ԍ?�����{{��c��</�K�/��hT�:uC|���k��ֵ�aG֎�G}�bs�ɕ�G����op����m��`��;q�;v�w��[���o���3<��g�ǎ��jrE�$�(���L�8�����9y~'#9�z�x�����"�S�i���j��	��<���8���)���x�}��h4.
�P���W��y.�q��W�*}ӽ���[����|V;�Y��W\�J��������t�k⸽v�ʕ�<���9�;����<�&_���M��nG�EbdT�;-#P@��R���a��y*Q���WJ�J�9�f�.�L}/cԿ�ʑ�V������[X�l�*��L�x���Ϋ�q�J˪���"�2F������g�'�\�����^�V� 1���'�k����� �%�������t:��H��</�Y��(��(��|�Y���]C�Q�~�@Mxű	u��ޞR�-��*�Y֭�Mc"�<�z�$�CL����l1	Z_3=h�	2O�^z`k��X����~��?\bN�	��Hp*�ٲS���ړeY��Jh�aO��G��b��s�(k����C1W��_���`b���n�+�mca.Ea���A<��e�g�I<�LM���m���8��j�!,�� <�v<��Q�*�g�@Vxz�_,X�N�mJ:e�ZhJ���N;�X0���]n<m���n��'IR��z�,}<Y��6��T�N��}��B˶�|\�����z�(�~ͦ���w�\�W��a�n�&Y֚��^U�$��dY{;˲Kq�\���b��,'q+�fU<rU9q�V���s�<Ϧs��ؼ��/�D�����f�w������,N_�4����s�>�%�{ݽ�ޫ1���r��g��[����h��o;v��w//���ڵ��3goi%iZ��?�_z�u��	w��E����*���s��Y��Oژ�9L���S�np�z�8y���nqq��r�6����2~֘�'Zv���K���nr����D'��#��o�:dSC�vU(O(�Ue�����p�������[���e���c�^������ǡ�	M���Nq�ߧ��.�(��2�����C�;������������/{��O�Վz/�������|�D���t�<[K����=��mnn��j�o˲4Ue��gϖ/�˕x���(��mw�w�~���cy׹s���R�j���Tq���}��]��v���f�Ф.�'�p��U˪��g�O<n��.Zy>%����4��������n0X�Ѕ#G��	�bd,�ǂ�͓�U���塔���SV�`�`���p_�&�e@P>��o%h��{�Kصfa��T�~�C�qQU�,�$yu��{-�����VJj���DĪ�Al$̵h����HyFm���
f��ĸ݃��:8\qOzpB����c����Z��(�Oq��u�j����ġ�E}�~���g�<�A$�����-�������B ����>$����ޣ>�Ng�]\\��]��P�Oy��¶��}�]�`P�Z��]}m��X��7�`��a���[������	b߄�y�g� 
B����ص�5��xњ�G`>��Q�Ċc���R5HB���w�w�b(I�c6�u�{~��\}�lc�\�O��^���L��u�waQw�(R=�:^�`1P{������󂰮���Y�{t�����Tv�ݓ,K-c:����d�¦{�#��e�x�4M��E�4汋�.r�8���$ُ�h/��^�ZmM����*�QU�q�W�عj��8je��s���y�-�E�ϊ,˪��A�yUe{ډ��I5�v4��c������*M-77��8]�<y�ZY�*�~�����~xn��|�����'/��/�G����y�`���')�x�j%����N@�e�V�B��l�E�l^鼩Y:�#v���,?������z~llͳjEek6�f����:�v5m������|�1.�k�M&݃{o�'Q��~�錿@D�8�g��c��=��iԚ��Yke����i�<�R�·j�X5!���������[U�5�Z���Im���޷v�I�R�w�q����+��;���R�����(��s�>]��U>���"��O�������ޥ���}��_\�����0���[��l�����ܑ#G˳g�Ə?��m�klO����[M�nnm���������ܹ;�r?,ϯsG���J��]w��Į�Q�V�Ú�m�w>s�V�}�c��;n�����7g�O%��خq̋l��k~����ˢ,��͍�7~�7,o��U9�v)��[اnL�'Kg;d�6Ԏ�0k�K;̃镩����Nݍ7���[�'���?�귾�>����W��_1�{����d2�vV;�ѵ��8N_q���{����$�B���q��m��f�2�������-w�q�����*��N�(vS�T�˵~���9���P���x��q++��ĉ��Ť��j]���/_�l���_���K��K�/�Օ�R������|�ķ���N�nu�J�^{u���V?&�%:��[�Cj�=;�!Ճ��]	3�W�^�I��ջ恬's��lIgϰ��m
���o�V['���-.zqP����gW��z���G�j�Y��D���e�=�M��o]O��5�Щ��{}�Aܒb�l[Ư���Z9︾\��8`�;KP��ыm[�>#Y\$���������@��{�9xsCY�0�����^�\�O��h�h4��}j�S�/!����(a��� �O�6(�&x�vc��z#a*���lץ��y�5��Ff#zA*{V?*VZ�݉�^���>FK�J�hů���P�Z��}ɓ��B3����W5��^�o{�칲�K ����ņ��[5��mmm����g1pIl�9O�&�_��oj!8I���Bb��kaKݟ�]��w <_%�j���p�/��6�\������a1��e[��EL�_��'+��Tj��}�cгE�_p��O���Z��a0;�b#��L�DY�}B�j�\����Q���;��p��v�T�bk�S�0�:�Oת&�i^�y�β|6���N[�e^z�}���X6yQv�=ݺN��z��W��'I<�YY�8N���W�m��2/s��)�ٝV��Y��iEQ�ɪ��4ɪ�|j�5�Nm����J|�ԒoK��~'OY�dU�đ��(ɋ<+�"��?�1P*�Q�Ω�S�F�%U���W��_h9��/�Y�¶؝i��/�K9`�|>��H�V��,J��2b�<��yYUc�dY:�NgC�[Wj�5�Og�B;�v1�N�Y�M#�&�y1��,�#7��|��'�M�v[;�U���·z�n�]>�fUU�V�vUN�]Ͷ��Z���u����nlT�kk�����������(�����ҝ[[����;�\���?��C"^�(6~�����v�l��*���ޮ%liӘ)�A�Z|�Ue�sy��qKZ;z�yv5�v�}w׋_l�Y�l���	�v�l���~��x�V�A��:tя���_ph�_V[*U��P���z׻��K�]n�~^x������o���wm�o�՜�-
�|��_�x�	�q�j>��oz�7��{���?��|���
^��� ����%�I�:�:�.m�YYy�'_���q_+k�yɋ_�:y�Dz뭷�흝R��&MGj�g�%Eɨ�=�ʋ�.I��ڲ�!���r8�Wɶ��c�T�,T��f�<��4W��_�'k�D����i�[�u�%��cǎY����j*������7�x{s˟�����߿��d8&�wv��U�����20����`���i6��}� ��B-�}�\n���0�G��n��~���3�;��*[�eR��8���ݛD�ڥ6�-v����7ݣ<�>�IIj�u���g(�3}F��8H��is��{R�G��Y�ф��&�Z-�Z�r-�B��/���9t�~|=n�D`�	����WՁ<�p�1�����&s��b��$]j?����D�v�YɄ
	M	b��a��~���e�j~��*_��B�{BK��b���bD��gDqc�~�@1�ynI�O��Z|�m�+Ժz�7Q�P�C��r(��=�~�d5%k����=3�=���B�>^9,n�s�4qFaa�(�a��O%�la�nY��`#6I$�-$�u����F��]���v��vdG�NH\Rey�N'�΍���ښ���l�]��P!3z��;]�۠�,���*,�$��@��ؑ�m��@-�F/y����A��g4��ł�F���P�y��Z��,w���Y������Z��=��6�S��z��[+ܬ�yf��~K�'�J�q�s��K�kl�c���|Ȕc�M��g�:���F\|R��r��d@��q��󂗫��河��cٵ�#I�E�Ï�4K�{9 t�zqe����um�H�W�D^��|6׎�A������(�?�N&�Y�a��R�9�N�$�4ǖJ~�L�~gS�d�����vi�g�i�)YK�Zy��U��gu�^,��t:1��������9��J��J���*�~�j�QX^]��4=�6��ŕ��Mr@��Y����ͭ�B���Hĩ�L'6��eY�'�����f�r����</�QU���t6�t:��l6.�bE�$��8�6����h8��,i�:Y<��I�����D�@t�n��St��ߚN�?t����n��E�Gܤ�+^����c�{��^w���R��Vn���ډ������S����#��$�._��n:}�yx��N���n��X��q�9�ͭǇ�{Y�ƒ�=����[-���V��a��9*���>�H6v���/��S娢P������'Vh>�g�.v�~�ؿ�Nfx�un��H�$��ċ�;~ꧾ�;X�������k~���
�_��_�>��ϦKKK�s{�<�W��u���x4������0��VN����KV22��K���"/�*!��5���K�M�u{�-�����hT�J��<y����N��iG�N^��e+��c6m������(h ��B�Y� �H���e��zo��;ku:-y}�;�t_J\�
H�OM��M7���8���V|��&MF*q&Q�kx�n�A59�^,����%�D�y�Fc[�x��� &t:����'i��������=�A Jh�E}�{�0�6.~ҲrjÑ�z�R��)�L���D����*��� �T>E�v�s�G�c�uj�x8�IT"�DW��ja�'d�S�A��jF��%�)��(W��@<_`A�{��K�x!`q�
��g���l���-��V��]ha�#�*�d6	\]C�ӄaq0���������U��M�g���t?����'4h�$��=�~�֓���0n\�n<��^�kBTv'&�d�ŗ�/�Rۃ���p�P��4�Wx�~g���Z��N>��8f�~qbBV���~�� �k�P'o(�Cu(}�H�B�BF�ۈ�x�{��_���O�p|��-O��I�+a<�aW%������a��g�o�w�W?��{v*��V�~���|�^��>��/��4x���Vq��{_�ӿ�;����[���� �-��(��*�}��d��^�܅�	�-}i$%�&u�?���^�_����E�����?�j��Yy����yĪ���u�P��{���P���;��Õ\�;��kB�����eu��o�d�agF�ճ&�	�pz���摐��2��v�mI���)+�:q
�    IDAT����Y��z��W=O�N�Sja�C��c&,p%���aGF�=~A�j�&ZN�w���7>�� ��~��>1J�� ���\����V^�r�Ǳ��5����Va&��v����;kA���S�N���-s�h���!ۓ��!J�ʗ�;)�Jz��*��vR�zE9��}v���4����I��2/˲�&���ӓ�d�����V|��[�����;v��{�k^S./-ǿ������cv�k��B��ɓ����Vk���f��h�ꩧܙ�g��ή;v⸅4Y;j����oq����������OBQ� <�����w��ͦ��9�<WoW�}�zhṵ�e�h+T�*��/��/���.�s�.a;;�^>�Z�Z�_�@��x�FXP�vy�k���{��SU��������������7��q�ϩ�}���M��^�S����֢,�-=�ą�������������a�N���$�bN4�����D�]m�?��S*� �mm� ����z-�q���d237�ԗŲ��YH4@���Q�s�����Ah����Y�vJ��g��ì��O?�t|��q���W,NW_͛�Y�����+p7��(��2��	sm�j{[�;?H��M7�d"[<�:��f�'O�D	m�	���4��B��o��ګ��ݑ�O�l٠���'�6�מUMn��U��~�^^���Ԏ�&�ڳj����:T!�����i��U�&L4����щN���$�x&�U��ϼV��ZE���յڛ�aZ$�dGj��>����(Kk�a��[[�N��ˤ{��).K}�'3- �	-1����O�Q���D����q�^o�=�v�L�:��EJ��'�N׽�>m�V"��	�d��V�u���G6MZ�2�{��	���݀|n:
ێ�y��Z�*�#����l��*�����8� ��=�0�á3j�1��5���:$�� �,|C���	���>R_h�!��d�SH��5+5���	�S�|�1��pr�eJ��|ȅy�����v4�{���[����N�_���eĞ���h�@m�݅�L��+���/T{u������Ņyլԟ<��4c�,�<�/��������3Ʊ��L���El��:���Ś���K^T/���v��ߛw���K�Mg>!5xHâ���!�%xyU�%��aW(0��;"&tK+8X��z͹1��'[(QY_�k�Ì�B(�v]W���˗/�Yc�8����cA�	�^xK��yAs���b��
[�XZ�{	�4�T�<�د�Xc����;����x��ֳv_jvtM�lX�����}~'G�-�k�)O�2�g�JI�*�?A�����gX���C���ة1G���X��իW܊��,1+ɕ�"�8�Z���Q��i���D�M/�23vU�Z(�[�}�-KKK3��j\�t;�B�&��U����s7�xS)�����;݋^t�����L4��\<��Wd��SO?es�^�B�ҷ�rf���:9a���ٛM�j����v@E��y�t���k׮����W����ܧ�>#�>X�C�hüb��`W���z�v�~���=�ȣf�g}�=��{] �:$�����P,�5��-�9��gϤ���!�?�O��~����;�ę���`U%}���ϗ�)�S�����篏��ߺ�����)}������%3i%��U{ȴ���>g+)J��	�?H��I.CN�$�V��gӀ������L���(,�O�B$��+w���vwwsy�%x�W��͍�:)Ǘ��Jy!�3LD�xJմ��
�taKO�S��&ۦLӃ�^�/-Kwd��m�ol��+T����ow�.]2���J��r(;��VĵU���ζ=L���[lҳ�ʺh��*��cڠ�Й�^���:x�o��%�����Sf�AK����,�����R1����@����1�A�g��C<��,����%{���?�~"H�7m��*���`[Mcl�EV�� ��PIh�y�b][�C����<��{�h��P��A?�#�~j��@U�Bp�n��X��~>���7[��4��w����-O��c�v�b���Z=��}/��A?��M"Iό�B�>�0��޳n�
e�v�dbq��;�B<��U��S�E���=E�'��:�Z�n��A�t�-7Y��{˽w��o���DK�|���$̐8�I�����{|���[��x������>��L
����gܷ< ����`������ɮ�����/�� d���:d���{Y�7��u���/���b^�_�%b8|�]Z{�$��,���z�+g�>a�ě����}�R�����z%ԭ�h&��%�h��Wي-0�0"�OϺ��: İ�!o���%�󃒑֤�;���(bK,��� sbԡ�U������^{�C|y�M|�bB�l�{��d/�b���5,D��Z�ڡ@��BK,�B�d�I9�l�\Ϟ����|L�2�C��Ⱦ������Ʊ-f�i��k�{��3�{ް���B��V�Ǣ��0�Td��[B�G��6�~����#�X!/�|8N_��>�ּ�
]p�^�m\�p�k�n6��If
���׳��������h�Q����B��Z��L���C�|�����A�$�l8�4g�z����bg:��
)[_?��O�~؝8��������?���VsW�3g��m�/v����'��+��M�	^�5��O��PL{njի늙�;	�GyĽ�k_i�Q���^���L,��r�n���,��������D��x���^]����=�P9P���a^��E�9�*y�˳7�U���SO�Ν����u��|�7h!2�#���v�&D���n��҉�_���~i��uC��}E�*4��O���._��޻���O���&v?�яzO��оjPTb��?aF����m�۵�&��A^��M-�g2)��q�j�q���O>�d);��FK������@��'6���ñy�?� t����ȑ#��1ඍ<�"�J~[Y]�%�����GH����uْ�5c�˙�|���cs�V�a�NBW[�2\m�ϡb@%h��J��o4������&�u��䁓a�_6�E����U�	$}� ��������y�*�V�I:��%0��+�V{/���D��K����\��O�yh�~����v^`��ĵ<@��~����=�uHB�h� ��lb0qh����:	}a�ǻ�W�P�,5�(���O��!�A��{��V�ru&��!�q���r�?��>F+�;�\�pѼ���b���Ja7:NZ	�����먅����F��lL���^�5�t���'ݹs�,3X"M�y��	[T|��pǏ��lYM��{̾��J}�c�?�^w����>�s
T�DL�uY1�Iμhӳ�����?N>L�{�CB�8Y�ϡ�-]���S���>�W��X��ｧ?�0��PB,�y�,9�{4�ת=�A�A޶syX��K�:���{���[�_(�v
j���g8�ə�X��xe=!��J~�P��~�8����x3C�v}�p��}�u�"�\^z����m[_���P'�p8�~/�u�{��Q虰�x�"���������4O���q`�Z*t_�����R�E��q0a�g�3��� (C�Ex��(=bX������{}^]�Ǉ��~{�5O�:�]Wv��7����ٝo�	Lg��U�C�tȑJ��H�w!�"��汷�z2��K���£�5��>��':��%�`U홗�A�����M��V�Sdi<���Nz���C�B>,<��N)��3�ɤ.��żBq,��Լe�6�� &�ލSm��ص�)m�o	�v�]��/�X(���}��ti��$��*g�d2��:"������{�|����㛿������>����,�W�^�m\;�U��F}�X]h�����X���7���7�t�U[q��/������~���_�2i�[�<���۰z�`�o-)ܞo�{#;�Ї>�~�߾ׄ�6�j�Y���K=�>�~�-�Ü)[Ҏ�W�WYy�K�.���U9�W���e�ݶg"�)�nA<�O�#G��+��O�r���������}�3�������9�umƕ��?}�K_�-o�ѷ/�G������Y^�:�V{JVS����2�+W.[�ݰ�J�@�z�݌\�x���gY���w��]�%�]�pa��'��x�қ�$���y~tssS"֎��jz8Z��:�,��z���g�ɤUO�*7��	��`�K�	m#�D	��%��[�a�P��젆�'BH(I�I���Q�v�A��_�X�G�'ݿVg�:��]uf�	��}���b�>�&�:s]"��V�y���P�A�Q��W����4��j�ı�C�_��g��#�����?4X�3�U�2���mnnF]'l����8�Y������^�x(G��B̪<���t���AI"L�f��2�s�}�ٕ�<��Ӗ�xmc�^D�ٽ�:�O��"L��<���9�V	����j�dC��hP����:�m�{�%����}i7Dm�HW|�&�n�5� y/����c���>C����c��� ��#���؋�����v�Z��=�.zo�����a:~B����@��P�j��'zI���e�!FU�B}�Ŕ��W��{O]�:x������۝��A��a+7� vW
	W�'�{>�Vs��>Z�;2E]ø�&�V�]�2�����>�&������Xz�v4��D� �LI�݋0Ä�yur��s+��4��r�>a3��p�R�0 M�����-�\^�:V\ai�CLX։MV�^������8n��8��]{0}ȄّF�"[��"�	ֳb��"(̹��i��{aK[������"&�b����	�ד
���l�j��]?\���y5�(�T��؂E|½(����y�1�:�w��g���%��b��*(��i���f�ĲU��Y�hŪKR:�u��V��|�,_������l!�z�v�Be�R#ǂl_s�v�R�6�h�Q�v�4~*LO}l㴅:ڂ�	1ǡ�;���J����٭vv5H�8��}�Q;h�[����}؜E��j�x$����I���/%*Q��~�aw��Y����n��vw�����׼���D�e�0N�/������~�m���*=�q�r`��-�x�=�!�浢t�=����_��<�
��s������Wi~������S'�������ߖw���x�Z�j���㥅E��`�MyXu5��̦/}�P���������{_p���~�m��͵�s{-�A�w]�|�o�����s��N�k�?�'2{��[a��^W�^�%�|�5��t�n�����|6�t�8��v{���������?���ċ�;�����t�TU������f�7����^4��u�8�M���E�����z�`�*3����A����Ǣ����m� j�nirz�
M<�� �B �8��S1�*�&C� ��!`�=�}�Q;eM�C̪���VW��:���I�<��=��^M+k�7�z��~��hҐX���nw���Į�lR�>�O�w��V~в�k��Q
=xv��%`���0����Y��z�V���c�g��e��M}�Ŋ����y�ud����i��`{�δ����I�[����������I�\�SB�&��Hu}��{����'9L
a�>q�Z���ާ�k�6�S�	L|e?��:��W�~�[��~��WF��
�I�y��(�'~���u�و8��$J}�}��ڢ�+�T�m�r��bA��[�V.��6[���n���o��be���Bu���-��Wu�{8�1�>��Y�v��������o�9�'���q$�VO�Y�CW�]����L�#�h���u_��2u���xӻڙ_`�e^��`������O�����S	�̨M���)��3�m����K`"ӄ��5Aja^h�f[���F(QX߷��m���01�1�!8�9����=�S��	��&�r}R�����;�q>\���5���WL�O��]�L<�Ƕ�1(�"��ɍ�$�:�ل���P.J�5����B��a{c�A�G��x�=q-\+�j����#T��p�:�Zs�v�B��ƌP?��-KK$�)��V�u�;�o"�s���*{O�r_$Z}_�C�B�����>B������IY�܃0[8�B����ϗٹ]}-YUX*��\UL���iU�E�ƨ�W��Y��zs��c�Y����7���-������p�b�yV	��!&;�����I��m�m��n�ɓn2��յ5����k�í�`%��
 A��m��c>�w����`P/f�ck!Hv����.x5��I�-
O���w��-�|%�~e���
�/���e!����w�����ʝ?����?��}����p����1d��0ֆ�����p�/{�ݿ�W��M�u�ó��}��ߝ<��7�y~�|>����;�$�s<���vm��m��򖷸����v��g{{[A�*�*~����o��gΞ)O�8?��c��ŋ�nͲ4�?y���x�����?﫡?^j��K�������v����l�X��EQ�M�7�ey�,������"/��"��y�)��2L�U�X+��v��C�a���i�mKiwo�\Z\�A4��CB�hH:��D׬=F�B��-�C��X�~n�o"$L��]H��u�t�zr���ղAP�e�֓�ek��3��$�=*=3�M���b2UZh{g;V�j�X�O�Q	9y��`���W;8�N���E��vS�r4Y&t'vh���U�Y\$�4X��tm�l0���>�Ė���� |������/1?|`G*o��uyֻv���)i�S2�&U]��>�5ē^�����MVqDO�)q�W�PuA}��ש������u��~��{�������~'���kK��vj����$�c��y@���rnIo�F8�D���xl�Fؒ<��jQd���'l�}�~����Raj:�N��A�!(����Hq�:�Ӌ6ُ���[�WI��vG��Y��$%�~N��Wo��Br_����ra�~nq�
��L���l�m�y�$��*�;��hѣ�$}o��u�q�>�Ӯ�
�[t�� ���'a��L�䅟/�e�H��ض{
��2����I=��8� ��sۉ�$iz�.�-�/T��$Ϻ$�a!*n�zM����PBc�� �C�Cr���-*�m�N%FB؅��ק� ���uBN�<���M�-����� ��m�R/���z�^�g>P�[�����`���y}5���vT}�B/,`��aa�� tCIɰ���,��-���Ƌ� q�*E�C�܏Ma�/�؄E���ױֲ%�ݺ�Gإs��{�1�w8Bl�?�����0���b��m�3%��l:�-X��>Y�v]W>x;u�V6.���RK�Yj�<��z�!�0P"�5+'�q�ۿ�;lN��?��n4�q_�9ݗ�=������U̶Xh��SM��yr}���=z����X(���w���'���ͻ��='�ˇ?�Aw��;�j�Bj&:l��N�rԵ��\Z��s?�c?f���w,��6������p|�-�?C�V�Sc����?�G6�������t�����:��q_�u_����5;t������Znye�<}����[���B~�W~������'��}yQ���r9/�Ţ(�W�\�
�sébſ,,.)���0(F����[�F����+���X��{~+���_�ۭͥ��O��.}oQ��>_���k�]�]*�Fky�w8^j����n�+�j0�'K�8Y呢(��l1���i��̦�SyY���|1/򥲬:q)%��v�ݲ��|��n�b��(N���IT��lނynɚƓq)qy�,�������E�|4ZT�V��Z�R��G{L��v*��7��y~�[Ž�����i�qQ���h�/.,��N�D�&)/��@����Bb�2L@u��	a�VP�.[d��:�p��yO5�k^k�ߟ�Uonn	���>}U����H�V������5��3��    IDAT�'q)�Q��r����Wv�&����PX���������C���Dq�ڵ����kfξ�ުM���jwz���A��h�0��T�<�E���u(4�q\{�ԗ�_[�{{�୦�� �<��3}]��`啔=X-�y�7�v�<�q	Y��2yu��B���O������N���_�
[�����(��{SMt���bM����]ً��*J�a�G_1#71��>dM�W�i�V��uBdJ��RR����	� �\�����v$~��
�
e��!��x*�e"N�]��>�6�	�i��za��p�������DT�(�B�%�ڢ��A��8��5��mϺǐ�瓖�(�t/���0�@�Fa���0����Wտ�3�1�۲�P�-�<�V�d��|��Õ!4.�8n	Ͱ�o�_��D�-@+�~�?G����U����S%�+xB%����X�m��_B%To�/NB2�Ć~�qG��}�̓;�}�{<Ǯ�Q6�*a����-���*�s_&R	����R�������&������~�����
B��c�M�-��sѱ�Z{���}թ�
���1t�`��
�FJQ��$��h4����ߍ&&/׈�Q�DAЈ��RTC�u�N��w���^�1��gC���H��O�n5c�5�?���?�^sɱ�l6߁<����ٽ��z��&�=��#�o{��s�w�� �f<�p��N�ѱQ:15mA�ˎ�S{�ҩ[��xF��������իג�����hFU�s�)'��������dcp�@�ə�m6�PnUGf�H���BQ�e2w�Z�dC�.��2f�?�	x�5dKQ���_�4�;��A��O=Ų�ۮ��� _��ivv�9�X[q��}���d|��ѥW�� ��W}M�Z{_�Kc�K9�$��J��7=3����պ�kQ�C	��Ɨ/W�o=�'xS_�����j��-�c�:2qe����՞��뺻�����^��n�6@���'��|��5?�.tw��F�U��뚓��.�N�w�$���4YM��Q�t]JiX��Wk�M�>�,g�h4�l6��Y�@K�`R���9�#@�D��X���P��q�����bҾˑ�H��._�w㔟D�%��}q�j��"�ʫ&&T�=b&��_��3��9ڶ�`�
*��2�t��LX��� b�1�N~��Ȕ� �
�
��e(�4㈇�l@i4N�^��b2D�m,� 2 �Ť�4�$� �RRF�ͳ�u�ܸ��cLm����:�&��-�[E��j(8!��UI�B��4a��bF��`��ƙ ��d�)I�?�ĵE�`����4�x-�/C���hA��s�[@��m�C�T��H��3)��{�^0�1�7�j�Uin���4A>��eH�� (��2���t�v�@�
�@j#�(|��Sݔ�4~�����B[�c|�H9�`]:��<m��(��s�����y�9�ŏ���}pT�d3��1� ��	I�c|��h�D�qS�a�(��~,����t	��8�+QV�RiFcZ"�X����J�D�ؘBd��.� �
p�9�om����l�:�	�9�S������z�(6�z��i���'JC�?㬆S6A��q~�5��p�q�Ԙ�?4�a��v����u�i��6�1�$À� L�8�(ж\��0� H �A;�e쬢���l+<X��h�s;g�F~�,�_�CqLZ����qM� �q^Y���	��ctw�V�t�e�q0㡇�#G��=ŵ��##��Yͩ��"+��t�t��={h���F��h��M����bz��J�����K)O����t򺵆&�m�m��"�#߳4P�{z��=�^�Bi���KH�g~����xqN�tw����_y=z�G8z��fh��1z|�ڼi3-[B7������b�r���[N�r�Uk޴m�6S��m���c���7��߈�dU�ă�r�� �N������l�ru�֭*_(�X��+�i�����$��>u��r[`L��уC����8���d�߼ꪫ������{������f��k���������\=z�YN��QRq<�墿=T� dP��=��W(��$I���f�\G'�II��q2�l6� X�CݵZ�����g�z�-d2�����r�V�N��,b�@���ӎE���l�hGʹ����� �X@D:�X꤈Ns7*ȳҢ\e�C��p��3�Wn�X��-}�%��w���>𹙼��j�|!��i"j�c�57`G��׆�E�Z\��ڂf#�:��ϒ|%�(���B�, &4\�N�E�Wu<ϒ9�ET��q���ǿa��ŝ�`Ҩ�@e6����-+������]�\���(T1ϝ�,��Dlq_�-�	w���g"����\��GD8�iS���Z��+Y�!����=Fď�
��(Ѹe�
�)�8��c�D��9�Fc�a���d$3"����i�(p*���%׾��t�i�!� h��J$Nl�4���a	(��J�u C�7��l���9�XXę����� [�k��� ��gqQ/�4W����~�,��q�Fi�4[ިP&�`�o��I��D��Kj#���H8��]Ÿ��K� xI&ׂ{��5�^�wzj�����8O��=6�=njp��Þ����(:E�1�97�g��A5@\ L� r��Z�A#������Y�j~+ �-�F�nV �s�B��]R���1Q��5�y�E��!ٯ���	K�2��v�c% Pn�9v,Aej~����gG*8۷og�P�(� M���3u� w�t�z�V�Ɲw�[�M��o�Hh�f|ڸq3)H�q��E����}���E�֭����tp�`�B��(.x6ca�!#C��7@���P�M��rn5�ez�H�ϲ·��|`���_�?[p
 ��4148@_���<O�q�t�_7L#'�Eψ#�522��_�������2ww��/��u�֫�8�K�����SSp= ���1��B��.��M��P�
`�Tv��]]��T*N���-ǡ/._��;۶m[���;���/�P�8::����"ʋ(�R�LV�� J
Q��@�p\��]�rǂFcyWO�x����LO�J��oƥ��2J -\��I�Y7�7VC@Q^�� T�v�(k��9�f&Il8�
�#)d𘮀�]@/k�FaZk�X�#�ŋ��n@V�۬�:�[C�(0@8�"%���V��j-��s����� `�c� �X �hS
-Q�d�l�BA�jsw-���=�.JU�����p3ޙ2!<nȈ�!��H��\��ɴ((����51(��b9��/�Z�,�	E;�P6��1�e"ͦ9�|�d�h�<�����Xd�0~�I�ֵ-�"�(��9c����I�8.RD�>���+i|�!H�����(����������=�,WfWY��&d l�� �6�� ����� o���Ie�c�l�	J�d���pі{#���Lx��"P�ӮX8��[�U� qA;R�o�L���Vj_�����>E%� fӍϯ��G��Ǎj5�@Yʃda�L�v�9v8���R�䜰�Y8�ss�,�%t(�|N�8��3�+�W �P`	3vlL������N�c��F��Q����T*\��U��7�g�mb���B7��8�.F2�.]'��	+�&���@޶m7�	�1�8!��a`{y��?y�A�=�u�Y���*R.\{�K΢rw�ܹ�9��>8ppl�F�ڽ����~��d$:��q��=̩�O��Rd))�r�Vn����m����ˈ﷾y�]������"��Q�_^i$��Ҷ��4hAMD}�#�Ҙ�������$��Ȯ|�6L�t�?���"��CC\�=2<Dw�yk��t����u4�b^4�a&��}�}���q�Ҁ��A0w�B��$�."rr�N�ayy^X��
�B�b�
�e��w���U��v:�x���������=<�HaB�!��֪�Î�>_,���7��xa������	JT�����=�W͹'N$�^�h��T�����@e]W��f�,U��hl��HGCI�i�9��F�!6;
��A�aA�6E#���ʂ)IP,�E�)����@���)�d8�*)]pC����6c��l���V��*�qQb�j2��pÂF��q%�U,�~�"#rjd����>�V��*_[&��
^h |&j~(����8.2���!�q[�-Q��h/�%�!I����av�%�`9G���2iRP%Qi -5���}����	�ߓ�$w�s��Y!dx����f��qlt�;;�R\����I,� 7 �5 �E��w��!�g,� 6bo��.B'B
�p<����,w�4z��g��p>�7�C����lIQ����(�dQ-ʐ�NH�؇���".��8?�A�3���a�n��G
Y4�Q� \h&�2c��X��}�1��QN��@Q-٭�0�Ծ�Z�����Z 9KC�2�UDI���
���9�:� �2�!6��
�%��.6��YD�%c�6��4�`�̩�L�g�E�h.$�yD8,RH	�e�z�y�Y�L�ų�j����1.N���t\3�
Md����p��8@���m�-7��E+���[���-�m�Pi�����B��؆Zţ�-[N5M���ݻw���]Pl��:��s8�g��I�~��'�������v�߰��(�=u��-*gU�PgZx�9��wҚU+�l/׮������Ym�<ԑ ���j]�����]GO��e;��A_��[�?��C{��}6ҎFK|tt�~��d�\ֹ�M�Sf\����0:�a�ݰ�pw��Y�H�qS����W���|��۶m32P/���4|���홙����l�a�����3HR�����ڲ�T����s�qN���Too/��喯����%K�T�X�K��]�F���)um.W���o}��p��]v,��B#��R�=�玌Ī��7�f�K�j��u2I=ȇaҕ���j���h*9�"j\)��Ѩ�SJCQ��fɀK�<��5�x�Ş��6�	�.B0�ZL`[�WC��].R+2�zl�ִҙ��� �� dtr�+$�2��t��&H�!J&�a���/�I��  ���J�� �T�s��m�"�6���cQ��#�.86"���p'�(�yƈ$��(q@���/�R,�(�Ĺ�8�B�aY�/�J��D@ �� ��jժ��2"|L�`�R��I�d'�b�k�"��ַzٰ�I�ǭB3�8Hq �Q"k(�d��3�upF� �*ԘΉVZM"���}ʽ��6�� c|�o-� �{dZٶ��)�2ET��)�b��Y����Փ���L{z��J�ml��1��8l� j�41��F+d�Fb�����@�����2�H{�Z�q] �8�D��N`
#��d$��x��~�(�:�n�� �A������q� hp?3���p4}�q��W�_�0���$�viKmlcim��L�z.�a ���F��?CxN}Vw������y�F��Ғ �?��r�ѱڷ?��g��̰�U+��nQl޲���>�%���ldd�Ќ.�)^��كw��H8�b9��5�WQ>zGJLW�)� S
,M14�-Ow|�Nz��YK:�IwG�;�L���,2e�K�Dq��O���5�\��433E����l�Y�����N���@��?>u��8ԥr	u's�֟�t�蛶m{��/Ԣ���Pg�T���&"Q�N� a����}���������	��k_��ڻw�i(�G�g�f�Z��]�v�=�o�b>�1�r����o5nng�X�c�����t��ܩ�(���W
i&�t �t>��b�2��
��Q�YiECav+W�DQԭ�����(sss^�\V�>�2B��dy(�0i\�,8³��2�Y�GS�g�!I!�r�'NS�h�%������i��E�������sM�� ��\ +�OI4`D�-�}n�NX�ܷ�_��q��U� ��yJ���F�`�s�x��Q��c���x�ϋ���������E�
�m�/��[I�\�iD`:�=m�е���hc?���*X�*�����t7$`-o��N(�_|�.,�?���1c���Rpi�Ϙv��.�4��5�[�_�"L��k�����P_D��&Jk�D��k�'n��%8��4���j
�&&(�H�[��]��4���mw�l/�Pc+l�A��ka�j�j�Dl�����7��}��ڗ8r<���&]�n;\�	� c������Md eB�0��#�I-�A��f�c��9�ڰi�}�1�s �����K+W��@G����G�+���}���QM
na��k���?�7�m����a�y
��/�⢺��:mKg ^pxW�\���Q[n!l�w�7���B�������w�G���o�k�f���v����j�?ae��k�m�1�P������M9��j?~�Q:p`?m`����/�2=�ē�y�YNA��S�[صq�7��uo��B-p��~����v�|l������8*�Zz�zzzZ!�r�S�ի��G��-o�C�2�Su�}�� h*�	�^ !ɒ�͑��g��ɹ���������r/��;��X�c��� �?��O{�n�����; ��b�����x٬�9.:,��sc{A�\�\/St2�@	���>�SCNJK�T�8F[�|���4M{�8�@_'���G+X�Ez�6�E[�B��P�"b���z�j#ij:�IT�F��i͙�3��ߦ([�#Bq&�(IT�6lT���,`�st��h?(9,�,������3��H[�֒:�-����"@��ٔ��n���DG���RR���k�[K��k�g���g�0 �c3���yxo~a��m\�_�ؗ\� �g�����ب78��,���)�^�߳6mp� C]��m�L =h{�$(��wbS�hfl�5�5)�o�J%Π�8��#VUD(5p��G=6y� ��d��+�3�\4����F�d/��7@��b^�D�\�t��5�p��}��,\�p��]�S(�՘�n���X�N���B��m4��طs���@KPC����=s��e�p���~�X��r�͠c��N>)���{= _�s��@^|��t�w�Ӻb�Jڽk7��/����Ɨ�s�x�}�z�Z��ҫV�a��p���-Y����yp���d̶�CD����{�T,���U'�)�o�Ŝ^��YѦG-�b�� ��#�0�͍t�%���� ��{��}Z�b5�un�t�k^M߿���8:��O���e�^���P����N�z[W��˶m;�B������Tp����]�f�r���GC����vz+��ԛ6n�ӳ3�E��b��:��}A
ixx8DǛ���(�����<����f���ڵ��/���u�;��X�c���#��<K(��=D�w����g�755���\�U���T� �=�O���A�G���8�Z��(*&��Nt<D)��qܣ�.%Z��Q��Q1
#�+f�|	�h�R{�-WR@$�yH�-��s#� ;����q����J9VN��=є6;�X|��X!t�F�� AC�k�9�à���*�%Ϥ�m�N|�����l�8N�CY�)��7	������~�Y93\8;0q��J�v�,�5���p  0o���Y�BX��42]tX�"B|���-_�����ՑF�WtŲ�,;>0�� ��&��s��x	g��0l��e���kQ�,Ks���#tM3v�0-��_�K�j7���+���Z�.���Ǳ�C�d�5W("�8��7�@��R�B}Fmڴ	:��������e�����w���vÆ�t��ws��W^I��w�	P~���� ���o}�;��_
=��NZ:���8aJê�k����:ۂ<�v�C�����G ���u)�DS    IDAT)Xù�����>�Y��,3	Z��=Oэ7}�9��
-�Kk,�D2�ٿ|_���|�Y��Y
���^u�JVg���_�+�/��O�qjg7��x�>�e,�-�#���uۙ�Nz�+�����s����gsa8s����Q��p��A�~�RQC�#�y�fDmibb�=թ�i�����⊕+�|>�jqh����D�Xxd����f3�ޡ3Ȕ��۱@��ǰ @��w��˻��{{�R��LNN:��7P�9i�f
�DU*�!j@��#
�7�Bܤ�
Ji���&ITNSg�qh��8K4�t=�I!���8U&�!�V� �FҤ}�U��"�)&�k��1�$	��G �C�ܵ�-q%Gl"��:X:�I�k�Z�	V�F��-K*�e�L�֤�h�h�0f
,v�2��Dy��2
��{n���h�k@?� f ɼ\�� ����6S>�\���h�f8�F�(�e��'�VQ`��X�l���"�U��­�يV�s�Y�]�[�'�08��]�/ 7
4��g"`.��Ç��A$���/((���x�RQ]�2^kÁ�����-�n�M7��^�*����D�W^�Jo��}��g�I7�f��������_��8j~�9����w���n������z#�$%n<�gQ<j
5yP	������qt�Tȷ�hL�����xl�e�F���� ����t���7h�n��rP�����Dt��+��o�S2�}�O9Ҽ07G�~��p��. u�v��I33��8�����Ü�B ��p���㴗����,�u�]�_�N�j����x�[��/I!;�a����i�ӸB�5XT����{�n]�ꢾ�^�A���zn\.i��?66��\ד�^z�!u��:�X�c��~x6~��' ��MW�\ũ�Bov6U==�E�g|�O��a&� ��E�<_봜*���@F�Z'�9�l��a6���0���N}Ju6b���Z�$ ���m��������B�0E��`D��t�4%0��#��{�U��qc��.hh!XY�����R���B8�`�B#��~V!]my4�x�2JN��v):Et�z�oF7J۵u�3w�h[�h$��r�����#�x� C��4th&�^&�!���C��C$i���Y.B;~b
tJ=42�N�z��׮����Ϡ���raa�n_��ӧ?�i.�:�sSC������g>��֎L�l�@�s�}ͭ�`Oњ5�(��wP��v�	K�f|��xbGw����)��"�����raG�5��TjT*wӾ����چ��q���ӚD��N�X�b������ p�*x~O?m+����w�#S�_���1Rx�n�}���d��o��������e��ٿv]�/<8 ޅ���u�r�w� �{zj���{�r�����484����#:�#<<�����5%7��}����c9�����9D�t,б�z��"4����7���Nw�s~݋"���mz��4]��������n�*����䂉�U9��0��g
n�Y˸����~1�υQ�#'�d2��8��:N�J9����ϓD�w�DY�y��h���Q�j��d}��G�<��Q��6��Z-��a����8�>Q�t���i��u'I�$l4���?����.;iԛ�|!�L-��xs����޾�l�pх�L�K���'v�B�� �ڻo/�4׭[G��'��:��x�I�g��/у<�Ō7n�Nk���z���MR*�^ ^r�A�q����R�C{�즮R��"�� ��B�¶���V����nŊ̥�(��hph�����1�5�FŃ�ö���q����۷r��hX�4��;��;\pרU����FG�i�[hnn����hvf�c� Ƞ�p�j>��]e�?8x���z����x��''������(ʙց �kxOU"~.�^4#<���0�|���s�kpp0���R�uNPJ���|1�����^�tW�郲�:�X�c��:��-�\r�%~�1������w�K�8t萪իt���>�����˖-�cG�ѓ;w1W-tQ̶dl��NLpdzݺ�h�S{ό������L��E�+WQ6��/���H�E���}��RW�D9p�S���a�F�W	�2�_C���s|�j�A������̖�cѭ)
��X�	�Vi6������^8�8i����uk�Ү'�����Z�n-_(I�̴�5�p ��_�HM>�G�n����B��Z=�+����f#2GDs�פ76n�DK��ӑC\�
PD�!@����Р�`�RJ9sD�wV�X~�R�[���������;�X�c��:�X�g��ygo�rpd��s�9w]� =��cMPW.��B�'�[�j5<p�*�ˎ!`�Dr!�5;3K+W��Ch����Rf��OP3@S L�e+Vrњh�t���?����Y�`ux�(l������h�_���2>���v�~����[��+^执�Kb���y��㼆�`��I�j�ϱ�߿��}��J�֮����;�q���Q�����<c?t8Gt|o�Ÿ�
��������޲m۶�g�o��{Ϲh���?�~ff�=����C��bQ�*�h힘��7�󱣓4�t��$���/hӦ���ΝL�.�(l�gs�=��7
ݟ|!�n<�u~ӱ@�t,б@��9,��׽�ӳ3���.\;<<J;v<�*S�|�+�>�Аb��-��G~đ�+V2g���+WҡC����b�
zj�S��h�4==�T��"�;�l9��zZE���� ��8`��o����(��Pk��*<�Fi b�n>�z=��+W���Uֹ)wT�����O�t�!���\>�z�+V��O��'Y��𡃬Q���`����d��&����B�h�z6_���w��m����������W�f/�I�3=�M5+�@��\�<�
�W�a�8>�vD�ќ�W��5H����uk�B�-v�Z�AW������(ow��:�X�c��:�X�y���/9�-)9��7��g~�J��6m�{�<�@Q[���ffgi͚5r���㓓x�FG��ѣ\�p�l���@�^d��]��I�hB�,��h:vl��8����/N5��LdW�9DiA�(��8��Q^J]��E�����0��t42x½5Ňk7�>�z��^�:�"�VْFCT�X*��� ]p������!Z�g}�ۙ�EtB~��A�0rlF�$	�l&�5�q�\jA�ֹ��;^�~�9�{��-���zsm��z��u����^��x�ez~a�/��!�a��("�`�ׄ��Ç>x55M���➞noph(�������|�|޶m��Ǳ��U�t,б@�t,���׾�m�j�����wu=��N�P�@70���?�>1=�����L���	����[����P��r�*:z�e�9.2����.[F�b���"Œp ��`�!:|� �8���A��ǠwQ
�ʋ	tXſ9\ʭ�xk�]��e�˝ۚߴGk9H��f&x�#����q��B��󐑧��~ں�T�ȇ�;����:1�l~���8���<k��f5,7�ynFa���\���n9~|�7_Ā�Fwvvr}�2wea�FJu�i���5����j:�ܗ���I�,,�ѣ�X��Z��͸��K����>���΢;d��4Տ�Z��׾��h��:�X�c��:�X�c����^|��/��?���V>��Cܵ����tOO�B��U�z���!��՝�v�I�Nb�U�92D���8�T��Ӭ���+"�˖-���"��"͏�C�2��]�x�t��e�l���L�4�3��/(SS3�����)N��\���!m�ٴ�6�MG?uTO��9l���*ZF�Li@�������t��E�]M�8Nc�#l#l8���~��i8}}��T,~����_�^�����_��V��,,� ���U��� 4guu��.��e����Ao��'Og�徾�����w����7��Z��C�=���\܉�>��vggt,б@�t,`-�K.��T*���+�t���q��8��GG���!�{�}���hϞ=�!2��p���Gi�I'���,Dȑ����z����4+@$V,]:N��L��!~-�)x�)9r��8���~����	 �^Sdւ����:3�	`I2�̀���.=zl���������"x��k���Ip7�!̞�m�r��Vڟ�uu���.��`?�W����A�she7�]��q�С�����NDw�F���G��o;es��s�7���7������=���.�V�n��(�=H�5�MZ�~�\�����Gs�s4;7G�&'��뱐�e�]����52:�,
*��]CCŗ���؉�v���:�X�c��:x�-���ι�����\r��AWػw�[�Dm��8�����]w}�^v��ȣ�p����4�t��t�u��׼�5tםw��ի����c۷ӎǟ��O9�v��E#cc�X#�be/�y�)7���"iBG'�0ow����pV��sx-45=���u��p4x�l��8��ǧ�o��[x�7��F�1P3��y0�,����MͶo�/���E�T�e˗�`� =���T�����jFW�D���d���0">���F#��}� �7�j�^Ԁ��??459���V��a�>�}�Zoi���ņ��;�Оr s�B#�a�W��J����}�����n�JK�.����ۺ�����7�y�y�v,б@�t,б�/�.y��o����7���C�so�0�w�������y�]t�%�Г;��s�9�u�f^����W/��v��I�~ի8Bz�7����}ڸi37�cJ@������lk�$ǔq=��k/��� �W@o{���e�4pw�]�<�ڡj�A_���|M=��� n]� ����jQ�L�/�D�$�D�YxtϽ��+9����n#�!.���M�:>�:�Y��gx�5���^6��]
���o�-�7�<?�xq�[o��w��£�ssK�MP�����	A���ϸ����@����	��"R_��u__���W/��E���������5��e���w����Od��;�X�c��:�X�y��+~�����������W^y�ɬ��c�կ~�~�w~�@�D��J�J]]%V^@��(*�� �*$������G�j�z�z��~G	�X��~��F��6��J�đ�~�8���Ѿ]��J�UT���5������o�����?�
	 � ˠ1@< ��<VhX��J�`���eI� ��l�˿�1AM E���}/�n����TUDo��`�f��z�Y?K�j���YN9������Z���M_��m��9��^{m���[?s|�}33ӿ�Fq'��Tƥf�(�ъ�/z˩[X:x��/,�./��A�D�5��������?��O~�\n���|�X�������Nǵ��Y��c��:�X�c�_X\�ҳ~wpx���7����RB���_�J�����733���l6�tl�47S@����`)2l?|�A����X����^P$h~v�V�]K��܄� �̀)F_7�#�1ww���#�&(�o˒�L��������\
D{ҭ�~�~��G���tȖ9sp��ܘ˟�R�1 .su��͘��j�#� ��ۻ�������G>�a�H4u�6M3��wV��Y� ����3>�)ͺ~����t钛�,Y���o�����ߛ���h�V/�H����I�F#�(Lȵ��1�]�����cG9- /inn�2~�&''������}����_�%�} ��}wp`����w��_�y�s�t,б@�<�8��3~������|�o.��Bu�豸Z�y_�ڭ������RWw72�t޹g�$U~�aZ�|�ؾ�^��8z{�ofY�C��Be��L�z{�h~n����|�#�Bi ��tx�l��"�ۮ��x���B�����(�P3^���۾~;M9�Q_�Mњ髶���@j� ��f��
:�sx�>��������W�����Y�"_����,y�����Ӕje�����)�=@�vhp �S���w��׽��_�y`����>⮿������WU���A���i��г�W�
^x�"N?�tb��;�#>??�r ��"\~�gқ��&ڻoo��_����Ǳ�%_���}��W����گ-MS禛nR���*533�tuu9N�Xu���L#��O�Ɖ��|a��m[,�I���߶��&���Z�Ժ�b1�{�I�V�W}��ժ3���$�T*9�|�I�57�.�Q�8��f� �l6��� �r���D���D��?lA.h���*��
Z:�F5\Q��)���2��1U��ņ��J8�a6�n;v6�L����������������I�5�hNe�9}J����J7u�<���{���6��y?���tV�ɻ4Ǡ��~+�v� ������k�1z�јH�����8'���۳TZH���ڟ��{־��p?�����t�n��Z"�����MOO�����g���^�w�Qq�o���7]N���_l��Ӊ�!����ްasǎ�M7�d���s��W�gj���S���3>�;v<�&��fgl��o��3�km�oέ?��_���t�M �ɽx�>��W\�p�m�����:��X��g����ĥ�^�C��#G&��������~���g>�Y��e/cU��/����X?u�q���op�ђ�KX��?��
�>r�������t-_��x�'k��Xk���ː���*<�����O�'���J Z��a�����~�V��_`�+���{_қ��\�Vpl��Cm�8���� ��K/~�$�G��@n�
:GD�z�J�n�#G��׿~[86:��F�z՛����C�y�8������N-,�Uk�Dk_;�B;���
X"� ������-[���E3�3t��16�� A��\�����Y}�i�х]�����}�ݕ�=��R������C�Ї��� �^s�5��<::�lߞU�穱1Wek%�����y���*�Ӛz�8���@��n��r�v�$MpS*�IWW7t�u3lROW�`���T�V%RJ�<1P��
��@t_6�u�A��j�f�k�z���C��`6�71NC�2��͐�Q�I�(W�^#hdr�\6
r�L�l��q"����3:�b��L6u\G�@g<��~�[�R�������(vc�F�����92I���AS�������0RH�tuw����j�%��=W��ϟ�ku��2(8�z�����So4�B>}C'�"?N%��y��d2*�b�/���7��X!�����2�r��(L�z{���
H�2<?b���Tx��AS�ge���N�֍F#�}?�V"��
yt�I
�B��J�$�i�FhONi�Xk�7����8n��e'MS�����\�Y(7͸���D�4��0
��J\�&�Oy��� [,���^��J)��V�Q�vK� ���7�͸P�QGn�Ď�p�f��l6i4Q.WH���8*�bS�I��^�ѩ��>D�1_�$��^)כ���q�Ui�T�B��n��ƈ����-]�����̶<c,9��\�j7Ց�S�M�ȅ 7~��
%!�㩔��s����K#/B~\���$�x�`�*�B'ՔSrh� 91��u�$r<����x&�lj�HD�x��b�9�G1��D�r�a��e�Y�Z.��2~�fq�4�x�(�x|a�<�G�����2��8��0�>[=��0�Q�����H�4B
�J\��Un����x�^�g=?Ci��b��ԫ���0Iu��|^�bc��Iy�
�X&�~�i:�������|>
�(I�8q]7�=RJaHi3�4�q�8�I.�m�1��u�</�y:D��	��DI��J{��?v]�T'�#�s5��U*m����A*4���O[���p�$q��*G"Q�	"S�����:ѩ	RyG�_yY    IDAT1R���qL�Ps�i���K=�`����T��Џ�J2Ik?�M��|�� ��"l��l�O��Z��eSE|����X�Mgg�i�\�{��XJ6h�,=����������y���,�8�%[�����_t�E���aOo���S��[���m��LLжm�8+�r�
�����yƙ��#�pQ��@?=�k'}�;ߡUkVӉ�i���e��(���Dx� �*\D��С�n �J�c�-�0kpL��!`�`n ��u3v��d����n�� �f��N<״`���em�p��h���P+z�������e�v���@]@qZOw7U��yM�9���SS
�����]����Ë.��je�w�w��G?�����o�������s�s�A�C�������N�֭[ǭ���╯$��R��fff�/^c����l� �7n̝}��4>>^߻�����S�?���[�Թ_�x�r~v��5�L&Ӻ�l��D��l��r�y ��֔Uq��X.m����j���\.��0�fg#���F��]|�X�q�a��@1bΚ'Wh��uY�8Z��j�h���2$פ  �\N�Y_�����wvvF{^FA����G�K��(8��А���c� �I�BŤpt1AZ�D���Z���ˉ�X+������/&&"�k�}B��[�������f��`(p��?F!������rڴ8�`�G�/~#������,lR���$���/�4 %���n~~^�㞛�S�&#���V�� X��86�cBDS�\�`c�؟|�{ �{����wao��|&x�'t������u>�W�8u86�L�&W)]�U)h�v�d����Ts�uh"&1����mp�`\'������a�P,h��;Ʊ�A��1�1�(��I���	���-'ͤ	�&�W��9fi\'�>�3�����m&pI�{�a&_�V�o�(e|
F��$ &
*�X��F
萟�4�}�u'��y��p,D5\קuևN�p��㷉r=7FL�]tH�ٶ�<�0�	�P�+|f��0�1`[&m3/b���O��<'�B����PJ��"/F9�݊�Ɨ�V�q�T� �_���Z���DkTO[Qy�2�1gAMp)Ld�0�����>��+���1�kP�V�k|B��,���Sȵ:)� ;��|�pjI���Y������)��B�)�k�/��8!k�z�BU;�m��|H!E��'G�p>S 0;�M��8~����(�v=�n�WEe����	�P�DǾ�����DgQ?�G��Lv%I{'��A0&��h&�uS�N�&iC5�r�:��䪦Gn��;I�LRUW��<'��V1 y�P���0���i��@��M|�Q�����F#��siVt����رR��ۛ"��� ,«�����T���K/9`L�A�'����_�r�韾D�r�&'��W\A�B��
��Ɨ��đ#�i�&��룹�yھc;7d@���D1sz��-23�7M4Gr1v�ϑ�ё!�A��0�����Y��kR\�v�=���w�N�ٻH�0��v^j��_<���6YG�״�!��Sb
�e�]��ׅ��c<g�o��
P������驩x``��N'��>�Ğ�^���x���o{����<��Z��v�Nܨ7�Z�Ω���q	�$[�T����16������=:1���D�a�Mؿx��1�^������=�:E��r����~%M	�o�$ �]�.'%]��|7����ӛ���.�s��(���cjvf1�Pk�cp䴧�'�Vk>�En:� �Y��a@�S8o����yH�R7[#����A�ׅjN��B�@a1�����10aca�uXb���\c�(�  I= �b��2����3$SG�@
��:q��z��TIl��� n������>����>r�g����Q�i���q. �A"b�Q3 S\�ѣGi�ʕ|. �x@�8R �x pM��j����T�9�罰P���0p<�1��ax� R�;�'�/:���{�X�`W��{�,^�"B�}�5��8�o^��q�����)C� �s�9Z�>h|?�!�n��Q��g������ ֑�-M�����#�+.�2l3�d%ep\X�-%�3�c���up��
�]���[�W1����=���&ZT"���{���7D*��k�fjR�a�l�g��g�r �Rw�Zx��\�_��M�L�y��l�$�ϠOY,9j �r]�qj����{CV  �ύ�h���8:�+��U��&�\� �1΃�S�9Ž�����:�N��-pfEB��u����E!� E<a�u]��u+���'�2S���-x�xqƪR�Y|az�'�)χ���ր���(����4���
qAsN,~�hvg����MA-mPܛ���u�����0o�;>�D��	ǘ���|����1pM���g�JF��i�H�i���XX��H����Q�^E���|>�	�?w�=W��\��<�C�qJ�~r���N�8���")Ju���G�JE)"�C��D�$ҩn(r���T�(�%i������8Z���$qY��٬��l-��r�J%��d2Ŧ�9�_U������ew�u^}��'h�m��C��
"���'m��8L޸d�R=;;��G]{�����#~q�m�1��Z�K_�RZ�d�׽;n�ˀa�`�Y�|9
�鶯�Ɲ��qm��R:����U �\`�5��WC��������`�Q�`
��x��L濖J�)qd�\�b�m9��-_���wP3�����Dy�)f.��(`k��(r�?�v�"#�-�4�t���N���Ut���;�Q������6p��R���P�(�es\�P�˗��4=�"��l��ڿ���U��w7�pyF����C�v���.��:��3���.�s�=�M��{w���ƀ���zsa~!�ROLLx� ������!ꈭ^oh 'Dp\�Q�����I�D̿�A7xfz�#f�yv���!Z�h4�v��M�p#��a��[�Th`p�$&3�#�!n>^�:� �Xx�� Z�Y�!@�  ��7@"?�k������:G��m&o��y#�h�F���@�����+B�����Qg��I����(��<!b;�} 86b�?�M$7��X�(@���x�s�B'dx�: ��a�Z����ʈ΂��4~�- �b�,� v"�D���7��Qk�e��Qk{�X�%v��
:�3Z� �����"���`rCd�͘�t�ᨑ7�3�|\�7QM�"���Y�)���G�6�@ �A��<y��k�aq���d����&Ƴ���\@��=5�Qx[8^&��� M���OaC��#g�1��s;���@���%�3�� ���X|��j�v�bW�[~���CZb�/�0� �p��1>d1n �˜�~⶛jd~$R��$�v>1�d9� m{�0�����Z�3��`��-��B!�?���3
C[�#�A�C��:"�fnr[c��?s/���p=�^!� ����DtΤ�J�����c�b��=���NII$�S��Ea|ǟ�>�XA�}O̀iRr,� ��8&[rη�n�)�vc�\������pk�|x���F&+�`��e�`�x�A�Ü[�Umƥ�Y��Z����3�6s��x�1k�#g�Z�_���e���6���=�S1��ԅR�4�r�US]]]�V�*JAڈC�z�X8�����|N7�D;�Hx�Nk*'��0���zEu�uq'Q��䲹j5��F�V�sٺ��CGU,�&ݦD	�MW9L@�Zk�?��Q�1�U�J3���0H����UiQ������I�D�S.�I&`�T*E�%^&��bɇs�IR?L0���Qty�$��r�
�"8�����􇆆y]��;�eN/��g��Gx��K7���N��c�	��u'����iz�ǏҺu'�S��r
4�����]�H��^�k��ݻok�/c�)��e�켉5�H�Y]]dM��!��%�혊�2����:��4�[�1�]�Z����Et�8c�4_��$�'�8ñ�S4��N�y`��6�Hg�c�9p`?gI��������n�˥�����֭=��/���6Po�ᓽ�Jp�\��j�ޥc�!%��y���*���)���e�_N?��}��餓O��[Oc0e#�J  �u�Vo�~&^d�ZC��J�0���p� �k�׌)��8�� ਏD������J��f`fE>���(�@�pG-�e�gB�&����)]���	nnn6P<DXP�%�� =bDD�9������T<���"��Q���QE�Ϥ6L*Z"yv�jE���_|�S���We� 6�"��#��1��F|Z�g���<pD4��"�!�G�# E8w�i�#׆�`�/S�Ώ�q5�R��Ga��op�v&�ց���q]x���A�rL ؖcpKö�R؜��&����^��/Q�Z��)S�	 @����G���Y���"`�Hv=�l�S@��l���:;�n�k���׀q
�ՠ=ʅs���	�b�c�&�3�]a�f�'��Ǒ���s�#���#�^���xA �R���3#Nn&Y���$�+��+�hk��b"�ߓ}��D([��ǒ�n߷L��o~�G *�,ƥ<O�D�1��x-��a8��z�ڑo*2�g�����d�-O~'`��ff��xk%��~�G�ni�H[�O��=m�^��aGc>��yv��4��g��e2|���sC	2�R��,��xN�csD��5)�Q.,��L��`˽�h�DO��Y0QM��V�S�~8��~qdUz��Ⱦ|�s�(m�z��L�9�Uh#��k �F��g�eC���K���xʹ	��Q`�/F��$�/�L�I�fƺ�k��u9Z���PC�!dXN
Ͻu� ��,�0;�1��e'������p��j:k�r���l?M������#�)i�-7�'&5P������`��u`_x�ڝ5�Q �{�4�a�5�y�L6C
���?��b͓��������3����L�4��$MsP*�g�F"����M[�����]�����]�d	ϝ���?Ӧ��	��U�V�w�^�^�@�����N?��.�	E�������"e`���S{����e�\�"l[�2�M�Lp�k�8��F���{�����4q��薵�X��v�3��k���$�]��81&�������^.t[�j�����,نc��.�,�����Sp���qw��ozݶm��Ǽ`��Fih?C�y��f>177�J�qLf���GyD��p�)���3����ן1�ݴq�/�8� 6��̴j6���hÄ�h4b��x�\nh6�
A.�Eڇ9���3��J���L� 8�W� %ȼK���r��O���D�o��5x�.G�lAJ��	���nY�\��h�/��-�R��SƜ�C�� I~Rm:���^���P�S�QD+ ��"� E� I�pUmO��x��p����
�pē&Hh�4��V�v������x-�@"�8WL�f�4(��JTGƎ'-��0>�lp�+�PNÀ�������i����j�ٴbl=Ԟ�22؏���/�͢�ץ�-`�� �x��8�k�3�k�M�{��X�5cc�A��r4�'<<lP�Hg|ԏ�D�'m�^`�=�����0�#v�')V�vP�}D(DBj� ̀���<F��o��D�e�2�C�Q0���#��ޤ�o���4��b�t9���sԓ��R{�K;9�͸�n�QW.�8��Y
�r�s ��A���Y�J��3<l��4R� ^ĕ����|��Q�W8>���S#mڈ;-[�=���ϗBy����&Y~&��R%r�V�OT�!���3;�XF�8���iv��rx���07ro�8aG�5� 6D,�c�T3���T+�l��P<��|��&cc����aZ�(�1S�%������1��v�q&Y��SC�O�3�!i�g��e� �<W�a���# ��2ob54* p��tXz�����`=0��3�U�'��uq��
�ǜ��sЈ�
�\��533e��c�|��|�Fb����	����5%v�6��ƸGƖ�a��8(l� �KH�	�9W����5܀��8ˆ��q�p��Pr�ɼg��mI�~�^3�Z|�e���d�l�2g�,w�t3N��`����!T���1@������	�q1����"������Pxbjʇ����XX.w�?K��w��UA��T�Hm�X�=�0w��#M���M߻�ڴi� ���:������]���@6��D�D���=��ъ��Z������)�hkO|�������r�w``������&�Ʈ�n���Z(��2c�k�:H�c��~�L� 6lhQ&�?��zz�[����P#�,	Е����\6o��������,��Ol۶�S�zA /��O-�����'�f^�*Յ" ��^ea>��8�w���-[�z�7m�`����zU.�tOO�BԴ��wZ!b�IX��� ��ˍ�dc��M�� ��*�yR�d�������HE!O��� a��1�0�W ��m���Z��6(aDCp�"�� P �.<���H��2�0�u�5&_��?�\�VL&�CHD�D7[��2�.G���v��#E(_�Vc/U"	�� E	D\m�!��,�uM�!�"O�(�G��ky�dBC-��/�t~-��+[p�#�-�2��H.���-;��5��O���"	���`��`
[��L4 @�/�v�04���"���f���� ��-)H���,� Y�`#�_*q��D��Z�Ţ����ȍ \�`���ļ]K��}�"�i�'��� r�X�%�K�>gM�T :"�<����8yѱEY�d|�u�)���:~�J�b���f��@���������0-N������G 	�*�-ֹ�g����m�D��B���8���م�ŒC�y�yq�P�}��m<C�{0��K\djsݚwL���T(T��[,�g�����)<3Zl�[�qq.����#����0N�M��{�t)��g����1C��g6�e�)�1��8Ѽ�[�,�n�<�� �/��gF��b"��$��(�E-@�g�(�1(�4.��费>����������ɺcǵ\/� Aqh��Fˉ�G{��y���2�8�:V�Q�)x�H����1�����4�uDB8�L��0u�=Cd�D�����1=5ej&x�4��m��α�� ��
��}~�(�����^�]��i{�#�E=��F+��G�:��f�5<��Χ��ź����(���� cj||;�w<��0(�}���� �������h�L/
%��m=u+8x��ȶ�z*�������AI��dp�h�;�����r�:^���(q��ӷ�����l�Moo?}�#JP)��mE�-M��mm#T��.��-�+�
۞�
�$�O�[�����vev�<����K:15E�J2���e�=�z�%�.w߲m�6+���K~^� ������̆���7Q��(�ʾ���4�''������s=�."� ���l�������
*<�x� �	
�.Q^�Zٺ}1���bB�F>Q��h���T�D!�1 i��ǖ�?&�V��V��,�g�|Z�"��V�E�T��4�]89�b�D���k��X� f
f��*@�6���n�C�*�:�#6f�d���V�(Y"�]���t�Pc����Ij�������MմQw�M��ߘ4%2�E�B<S3��V���U,J� (�s��5`R����H	v�	q?$j�c�|�V����ʌ�;�K�'������s��7&L�����B������VH%=�O"r1�{�N�����Xf�    IDATB,��(>�B�g�h�g@�����.(����Lt�<�o{om�u�w�sΝ�\�j��Je��ɒ,��ellc���lpҋ��:��������0���Â`��4s�n�-![�JCI5��7�������w%�4�ut$�wת���w�����9�����!Z�\��%��,�ƚ]��_ǵu�ְ��3��b��l�!>�}��:*�x����v�k�8=m���?�u%�z�_�gL���ř��ƚ����B�(ˆ�AV�Xh��x�htp��[�2�ɭ[��UH��b4n���݅r��2��V�g��r�B�u\�DQ��[�J�xǄ�4-2��&�v��VKs���wu�
�*�hz_�ww��(�3q�+ޗ���~]�L^b��Rӊ�tm�@��/��/�X}��_�C1���9]#~ݖ�;�q]:c����s�����6-�qAnBRYl���ן8$�^seu��]����\�(�ğWj�牸���\���r1w7�=�Ŭ DO����O����Ҹ��N�t|��GA�>n�g5V�G,vEF�Q|��ƍ;xq->W�8��\z����wB&��̜�g�1���I�'��>�P�U���;\q+����~��*��:b�J�˦1�9xi)�|����㧭�Þ�{�̸q�}����y�P�%n�B";|vl�n�i�{�X���J4}�+����K.�������̣�M����Y�#Wm3P�9Pׂ��vm�ύ(95_�<W�Ţ�m��?������>S�]��)���4�}h��Arr'����c�l�Q,S�������c�?���֞|z�<����"��Mo��ܵkwPZ2�{H������ڵs��+.�^y���s��;�y΋�yx�2�[
��W��=}v��?w�uE�_"q�]8w�%�p���̊���J����T�&W0өS�L�3~Sh�d�TJ)��#˃6M�fEP`8�V��bj(P�IG��C/�rsj~Y�ˇ�����rŜ6�h�Y	R�0=Z�y5�Oi��#զ�D��}�.r��۴v�:N	f����(��V�.d�y��sT/#3��XNPv(���P����ɧe�ln�k��E��h6fu�*=V,s�IȬ楕5�dŭ���]��x���A9�r�1����������[\���[�YTu<.�􀈮)]˧�mk�^�	��B��z�^�~��9L4+\|`YPX9��"I)��m�8�]�?D��Bښ�-���~��J��/
�!��8[�8�U�o��[��<��-h�a][|K��J��͢�nA��syϏS�x]uYr|1�~u���a:-��D���/�������E¢̞1�ϺHt�eT1�b�����K���/0���,���R��a�VH]G���HG1눻�L��޾O��^��}���P��]'���-s�:���<������%���� ����2��[\ ��Pב_#Q��	���[���5�1���-�����[p�~�.����N4x
9�>���B���7��s������]�;W��4g��S�E�ZL��7(,��(Ztyl�_�f�/.�bI����#=��nH\tLΕ�ciTs����vw���W1S����;�:�F�v�Q�<�s��S?m��<ϡ*�mGf��ֵ�{A�V�	gϝ���'xb o<n�����PZ��1�4Nhg��p�j�Z���yRsd������g��}�tұ��&$eT��-���W������V�l��=��˯0�{��m�S-�&C�������y��A_��<����n�)?~�D�b�$�/��rOYh!)��m������4��ʠ���y��m�z�w�����0ޙ�����l�����y�tD�9�M�o���w���/��̀�h����-����ѣ�ʩŃ��׿���W����,��e�3��{�}�鲱�iX�2�?z���t{��w�y�_=�\�|�W�����_���ܹ'o_]]}O�߿!I��|�w��ևgΜn��1Bzue%��-Z� ׄ*����:�)��y�t-��DdLe-�0��y(ߪ_(�W9I�wܺ�?'���V��V$JH�ߛ���u��ض�����$z��r_4��օc��~�Y@]���r6�SZo4Q�z���*�ӑX�m��d�*�*��L�T�;�(ʭd�J�����+A���z��>�>yF�.?�-�LX�[��>��K����e�s�GD?�迬IK�ī^�O���=�5�㼸m���'M���)Mރ*KȆ�\r�%��A���8y���*�r��I;V�ww�q*��ϭ�jC���C�����u-�t���-��z��t�J}��c�����H��E|00��]w�e�P�G�����o���ͳ-G�^ѻ%�-�n�T?e��XYO��˭7�a�<wC$�~��ȥˏ>#��ŋKVvS�0	�����t���N���D��5�Ā����lg��tK�k"ָ�z9w�\�=Pu#qZ��,״G-��,iхE���?l�j�]Y[�q�������[e�"��P�ndSq�}���1�{~�1�{�_�.$}^���fv#&"� )�?.�ݲ�g
���c3��VMw)����j{��8WO���0�Ϸ��Z\f�`tK�ϑjӯcbޯ�����/'���5�~���&�]!�Ϫ/����ͤ��B?,�]��n*�%I�q�DڄU>�=,}xK7;�-e��s�廇�bj"&#���e,c�Tt�YW-0ls��2շTBV�w��k�\�.L�j��w��5^22�F�M�E4 h<d4�	07E���-p��Ȼ{r��i�F/�ɬ]�nx������lP��_��_�ڟs���oxc8�ȱ��s����%��n�a�,���9�H��W�'��_~��$���+C�XD�x�8ȝi��=vL!���^e���?;V/�]�$�}2�ٝ�
{^[\�(��6�{���?��ٳ�L���-P
�I�.|��3�Cl�nV�P���8��-���n��3da���f����h�"�gΜ�D�gϮ�������F��?�S?��χ�}�6^�[N��'?�sמz������H��������I���0I���5-�Dɱ���/>\{8�.8��{7��5a���a�]q[����Ed���ߊ5���mY&�m'�m�̳��k�����!l+J�\ʠY^<�I}LB�D���Y�K_M�ԕ��v�[	b�-}��X\�U�_՟�]��ͭ�:Y}'�#��[���J�z����D4�O�V���$��#p�d���rks2l��E�ڗ���Jɧ}�1�zɟ�3]hB��dM�-��Z�����6q��r�>��ֶĨ&p�����+M֞{W��{��J�K J(>|�xk��
\Ǡ�H�Q��OA=����A�M����ک����];�,ؤ/��������Շ��رc��k����74����W_m����u-������>�*�z@�I"Y�ݷp��-V�Pb���������ĉ��z���UjG�� �-}��-����xL��U�S��D����4�%@�b�_���zU �c�=n�-�g,ǭ�D����8�=�����gu�zi,_s�k�g?��h�EƔ�w�6�g3�yh��3$f���x�G��9x������*�#x�q��е5kSׅ��z�)w��O�K��S���+���Y�kUף[������a��/��@�"��ח���+wAr�>+����9�~�ˈ��8�A�,�b�J�T��9_$�x��r˦��ntA�F�p��Q�Zs�)���lkm�v�&��n������v�h���d�,�\�eY�\�Zƞ�R�����wOI-�1?�^&fʬ.�'^ގ���y��l�Me%�������J�/
�w�ww�p��s�,��h��f�w-���\F�De�Q���������3%��+n�ǌ,�J2�R`�L��l(c!�~���E}|h�V�ŏ�TϬ����D��?C< ��[t݈s>�ls܉rk�� LҢAh[([<I���ؖ�Wm���s�ȑ+�G>�1[�J��������ݻ$�����P����s� K{���"Ӝ�*k�t꙯y���C=������4�[Y���C��tW�,Gץ�UG���E��i	N�'��>�q�6!!<�򅖿�\��'??@<���w��Y܁���rUd�ܹ��H�c�V~�QΝ?o��Z��ۖ9ix�K�_��oz��]�z��_J�g��s��	^��`���w����{�ћ���5!)�O�9=����ȟz�D�܄�V3_]Yk�"w˜Z�����s����mq[سw�=0v��m=D�ä_���utA��~��٘Gtl+�t���0��ߴ���EAY�l<BU�	ãFu�e����)�ᴽ�U����շ4�F�mD�4������?o�kb���Z��ru�Ь[�����/��>K���IQ�cYQ*�L��Ԕ	d��S0�Y�إ m���+z�[@[�e�B�2�`��'M�B��C��A��i��,�:w	<Mb�c��$:�Fc���$��a�F�-k����\L<�T������Xu7�Ճ��-gsm�F���Rol�*}�t.zp��ڲ���6ӹ�U_��ﾵ���B�>�1����B���ks�(���{'��t,v}��r=���d�}I�~���]�-��&tg���-Ϻ�}�X�j�}=Pe�ѢD����>��1���g�9eX)-�vߔ���`Ό����o�~Կ�[�����~���c��Ų�G�)�Zch����:�.��~�]/>��^׻�CYc|��=	C-F��,��eT?-�vi�w�d�/�Bom���*5-]���ţ����t?s�kQ��_w��_k����_OT���Vh�ъ]����]�.-~n�0��2�_��_Ǥy���S�Oٱk����RbR�Ʈ�=#�"�s�J�y�ͫ�[g���X������b�|�����x���Q��8u����xf�4�,�ʲ����,c������k���8Ǩe�m��e��vsA-~��t��Q^_:�]�:O��L��j'Kb.�~*;O�����y4BlY�yQ��>6�-�_Z�=@��CY
ܷT"L�������߹��]
�O��_��an��E�풕eԶ��w�,[GL%g���4`z�]����oy��m?򑏆V�T9�{���������l.���v�cc(n*;�����8h�Sc1��={���n������<��I4�)h9�Ceឿ�;,�φ�ϪX�eA��J6u���+�r�x���䘃~hk���o�x��&x'-�.v��f>�#���������ʵ�N���fS~�������y�a��WVqe�Ю�ⱔ��'Ӽ��d�׾�+��[n��g���o�����u�EQ$?��?����tsw���N�h>�/[^^V-k�:4N�<m��*��A�o߾T�.�h5h6�ۖ~Zf3��Z}�0�OexX�[ܾ��)����+�X�ȷl��oc�\�2?;M��ߖ,��o2P̬����m���m:^��%�c4!�L���3�U�y���/.E���M�p�ҍ�	��#�tg�����JKC�V�M�zx�LP�Rtt�ɳ�^HL��w��Y���=$��rV�D��G�}�p�t~�6��N��[=�f�MaY%�eD?5���W�b���hb� ��b�Wgm���r+�=��C��=mY<�\�>^�iV���1S߲@�
]�v����tO!�~�Y����b.��#�V6q�?�'V�[Y��>�#����,	:F�'4�x5=O��[�n��1�!/�ǭg�[�����-�-s|z�.���\zJ�L���U�������l���w����d��>���2�w�P�:o/� ������l��(la��Ec��I�.M�:o-�t�8{}F��u�Jz_�k��0;���zW�bm�O��$77���5BN�ܭJ�V�������HzO�D����t�� � >�7]�z�o��ѱ���ެ,w��ir�����J���u�רm�x�0W�zk��9T;z-.n7��}kS���:�/���b,u��()c���ÕZ�w/?����<�?�,���{n,��4��v��RV�3~kn�sG}�p���v1�~-��J���w���_ϲ���]e>�HǦs�N���̌��Ug0P�$���W�,,鿮)7.�*�1Y�Y�g��OB�}��[�=�(Q��P�����:��������zF%]�����rn;�V�3�����������t|���|r�t��n�U�ٹ��P����Y[�Yi��9��O�3KZ���2�>�S��{��{�/��/�˚+b�c��M��o����S���ǎ=jnO�8a.�_w�vm�ܙ�<(;pLK�3?��q��w�������J)X���\�]��?;7?�����'�`SY��m��o�wLp+��|�uW��ƶ/&v�}w���V�=�o���H�շ�j�
��~�~(��_����>��%v�X���m�w���ݘ"�>��c�#G�h�|�+�����>����c�R���Zx�� ?��C����{�-/�\�5�W�{��z���|T̮�������R��������0�RS�&���U�}�4��u��2_�X�(�[Q��)�*�`](^>�� �"�*5I�e�Ge�������v��*>�!��h�T=YK��W)���IB���Mě�d 0�[�q��+E��]�eZqp!f[��V�nz�cY|9������ĩJx��}�qUQ�Zݕ�n���kR�O{0�����������z."eM�skD���#�݇N�:���\}O���w�"L�S�׶m�zl�Q��]�W?��ǥv$�\���19}����Xsk�D�Y��̬�����=h˅��)����o.Z4��X�����#e$�]+ed��׮����������MO��aV��,��6��d]�z�Sx��q�_ҷ�}�-cb�������������x?DN޿[�l��}��g��v~�]�:�()=����`�N�[�c��6����u�t�Y}�m��,8�O�m��_�>���/�|�s۾m�xLtf�*ŋ3�w=����פ/6&���ʷ�}��"B��x�r�"��5�1�5�������{T}�nZ�E���ݶ��1K�����H,v���v}1��k����Ԏ׽��"��*2�Y�4O���c��zdA�]9�ta,k��]q��|>r�]۶p*s��X���L1�9[�-г&����Js�Q,���E�Q�y���r'Fj+Ι�O�ˊt1B_���ǭ�z��e���ЖAȪX%��A��h�p��]v�+IgJ�[�p���p�ˌ���UHA߿�Х6��H�+͛�o�>;��ra��[����>gצx��L��o���Í~���1��M;���E������X��ҁ�zq�c-�*^�by��U�+�#ǂM+�}����oyk���Q ۹kwx�{�>��o�Rw��Kh+�	^ϝ�u�b8�WX��Rp���*��`8��J�R�=���&S��X)���=�n	����޳�Q-�6���z�ŹK��qn�"V9q�=5;��z�d8s��Y����f��I�k�T�3�0����[�Q���������}��i��M�d����3���1���:v�t]�-�ma><z���;�x�/\v����]�x������>������D�����|���y>ؚ$�ֵ��-�V{g��q��j_s�̙}�Q>��f�$�|Q�������j_��&�D�~BJ���U��:[�M1�0�c�v<���fi�Jː�f�e@�D���z�J�p6n�mr�"&Ib�T�S��`�2��o��o���I[	ŵ�V���^�%<��^>==ee;� ��2&~�1��8!7-3��Le�¦�$Z�R�����=`���|�����ҫ��*����"l0����.�Ԧ/ZJ_QY���D�T�u�\ ��ܢ��Ē�������N�*׹�N?]�4������_�
��Rȥ%`�I�
@��׫q�7���?X9j%��5W�+i���I��ܚ�|;�?kQ�V.W�TM-V>ڜ��"fr�N�?��2�22t�q���%��JZ�<��U��7`    IDATTn���Ϯ�mj�Yב/�4��t����
�o��W����%|�`�����-�.8M$�/Ll�\���LG߲T	m���Բ�j��s��Z+�Q
G_x�;	{��uح�~-y�=-���;*x����˒�c�M�/����r��Z�!�uݮ�B;W^f���Js��LT��r��S�^�g�p�W���'��Ɉ�v�"��>-�yOx��q����[��=U�,}V��JQ@NZ��Zf��M�g��-v����8~�E�Ħ���� ������[s�[�\H{NaϦ1�H��c�JVef��R��4s_���](c;���}>>1��3S��+Ziշ�b�.In�йĒ�Q��q_q�\�T��*�s����x��C�?_�y�js��w�*�[n��3���g_�ճ��Z��.���~�2팜8q���(F�=�Y���xl1�h���_��E�D�}{�~�z�)5�D�������jO�%1�]I�᧟>m�
e�P���Xڴ�R����<^�ʫ�G?�1����C�,����D�3NCtG��TL���������v��@m��{���u�]oB^�x�F���ʬ�ʼ��6Y��ϚK��OYNc��ʲ-���R |S�zLA:Sڦ���.��������X [\�yp�3Ӓ��}R���c�.�ߋ��;v�P�"+r�{p~~���dY6����R�v_�Cs�v%4����͵�Si��m����?���ɽ�����JR��n���0K�E�|�C�����g�N���v�V���ۣf��o%���l,v{����b�_3^��vw�����P�TuMUsL�Z�r�h�[��r�V�+U���*=����l�҅�A2�k�U="�Ys���A%s�o6���v��EI�{�)�`�(t�0J�T�]G���<��N��rJ����~���ٙ�p��G��pmu�7;7�k�Z�S����z�z��F���;�3K����W�͢9hLgâP��~6B��!�.�%�(���Mͦ]�tVdYZ���os�Y�=�7���!��hk�Z��Z�D?C����T���d��L6���,�K}���$n�m�E�^S��Z�_;6��+.^�1@���r7MG�Q��3i�\���v�Y�	!\ظ�m�/q���e�;�N:��H�iVdô�]+���x���'�����NTF9曵ҟ�\�������e�$mE�ɽ/I�F�!A;lE�%�Dk�Qk�'ma�T.�)��B2�b*a:	IgT�Z�4�������C3Q)�����*�1����ǅJ(ҤH�������E:�U9���H�z��f:*���]�!��D�I��yG��H��DU�:���*��Q��jTѐ	%^�#+u�hC�CR��onnvf��J~�o�[k%�Wyo��%DTe�R絚��?̛�F*�[�4�����t��d���_[���1m���T�d�XZ^����Q�������^�A����/ŢU���8s�-�T��,`���x�w$�=��]E<��d���[��n#z/�����ʨ�q�R{�W9>6/a=�F�B�|����YbU��h�����Z��E�[�Է/R|����g��"�틴r!���H� /���
�%t�kf�S��Ō�a�(S������S�r�
@��/�|QMT�ڂ�$��(��՘��|2�2���1��lĩ�]��2��U� ��g�Jx㦅l���L�4'n�3�ڥ(w�<���[\	k����)$H�}��+�+r��w#��}^�O�$f�P���0a�;T�R{��X�/w��r�K��K������I�ƝΘ�ͅ�D��(�+�/|�N���bi�o���[_p��?�Z�-���k��淄}�C�{���G~4|�_~��r?�9ou�ˊ���<ށPW}��w�ɧ�UW�+�&�o���4כ�W1�����r�kn1��0�w�L�>��C���,#����z�^��\f]g�[\�)fE��&��j��:�(x�i�k�4h�������'�?)���S���U��V����t�33�U���}�7!o{�m��ɓ6�g�>m.�^_s����W_���#������A|!ޏ����g�2�E/ˏ=�Qb~��wz&��;��~=z�ɽ��29q�D�w��bω㏝ܻ���x��<�m[����,,,$3�����l��a}}6�gݹ�͛�p1mw;��^�gA�f;Z)��Zì(�Z04�Qa���ۑ!�F���lT���QZ�2���,ϳ�ʾi����?��,I�N��I�I���`��nt{��Զ�,l��}7K$��bX$�0
i�$Y�5�Ծ���wҐ֗�i�e�D��̋Q#M2��V��h8H��<i��m���n��4EF��K�d�b�z�Pw&E2i>e���1�HeW�[���lŔy�3��|���X�!�Z���&�^o����N��.B��w{Y�lHh%덙X�:�LO�.\�E"J��4Z�d4� ��{�-[��p(�?HF&�m����,���2X�!���E�,�ZtiG��!����p*
��l�3*
mq����Fh�[���t�h�������ŋ:[�Xv�Xj��D��d���G�53-r:�{f�-w�L��~�h�t�ϺQ�����/�Q[��KHsq*��t�jӫ=����dnn>/���̒�U������S��-��/��|�-Զ��<���|�`�e�RX�]��[V(�z}��R�iG��ve��B�!6�ev�}.�eE�^�LX����"�\t���--����:K��3K��<������3q7/�|XI�T"5����u^�.ow��~b�����*�)�YY�c��8M��l���]8	0����|Q�EF�1�).'��o�����w��ѱ���+���nw�b�\4���Y�]f��T��/���B���}�Yxc�t��{�'��O}<,��ąg�I�!Z~�2-f�3e�u�F�����*\��d��7����d����e�XU:���I���?l�2>�=�}+G�{Z���G/���KOܭgѵc�)���~����z6�g?l����G�ѳ_����y�������r���j�r˚����ͥ���B�$�����w������G��ӧ��33z���ַ����v�{������y��x�[x����J@���>u{*!=y {���O�<��b)��o�������W�������g��$�7_SS���D�~v�SI��Nd����嶗4��DBϿ���As�w�~S���%��	�ì1j$��K�a��v�pJ�R�Qxˏ M��m��Qn�)L4�R�i���6�JJK3���a���(��`;4څ�Ң�F��I�&�`�Hv�T��|=M^�I^���F�ݖ�F�r��e͞�Di��eIQ��F�H��aV$i֐?��xQH|g�^��j�[�Ѱ����I��y��,It���&m=o��A�!SY��`�i{O"��ng�~���(&��N�Lq�
�]���	]�l��eh�A�tY�A?&����Z�WC������V���Q�{�Vk+��?�ti�|8F���r��q>k)�C"Z�����+++���֬��ڜ��MW�Wr	�&h�|ii����&Syي���\�Vo���P���2L@��g���F�,��@cZ�����m����t&"Ʈ3��	��kA�
$m7lZ�7���X���GAJr����&�jv�-�L^�e����n��y�]�������n���De0�������ܜ��ښY'�Bx����ŃvBe��L�)�9%V� �b����D�V���������K�zr]+V�bM��%#���mneNbY�u�X��b��X-S�(�ۑg�e���윶m���7������-($���{�7������D�ЅeB�G1�R���׭p��m�f.b��#�̟��'��+�:j�_���C1�����^�A���p�����}��,��g��M�T{�V�����v)��d#�A�ԯ�F+�&�g<���q��������}�ex�s�r4��ۭ�hϞ=���Р���/��Ū{�ϟ�%����o
������	;2]��w�z�u�{�����o��o9��~A�>�0i
/f�z�m���=��{ｉ��x.�5�p�	����h�>>��_J\�KlOMM%SS��qv��DB[�~�%�h����������]3L���R6��|C]�e��Q�XR�����,�����2c��~+�VZ��YMi(9g$1��Y?�5�ͩV�8BY�sY�cE�tFi���F��9Z��@���N�Ք!\�7d5MBtm�ﷳ,I�a��2�����3�)Kvik4�Gj<iHi#+�Q��p%��6��U�\"4E�oL#�jn4̟<kFf�`�W���oj)�M �#��l���M�h�-�!���Ĳ���#%]n4ZM���5[9�#�Czmu��$>��/qZ�L��F��^��W,��&(�b86ܧ������eY�Z���ж��q����%��2P
��>��J�
6�3��,����Se��q�]�$
c��,�+�N/�^�		�I7���S��A��A�SFf�{'O��u��� �M�"���I�k�ko�+wԎ��]�E�d>	%�w��ږ��9գXnM�q���b�2��Rc�ٴ����Y[hH�*+���'X�Q���Y���K�:4X[Z��=�~̖��B,�b��2���.3T�[���K�T�1Ӊ^^���sS�+�Cش.�VQ��y;�Yrԯ~���·}�Ï�؏[�	��w�w�O~����>:��g�ڷt���6X �,�s���'�G^qUx�G��W_c�ִ����W����+`ӊN(Vd���ea.�>u2��;?�� ���Z��8F2g��C���[�&���?�n�d����?�X=�_��"x�w⽤��fc�m۶�.�]�w�~i�ݻ��c玖,�1�b���T�~-d}_[]��[ػ{����u_�����}qϳ���"�4|qrK(��	)�[��LN���znn.�p��ff&Y^^���ED"��^O��e�Y"{�7�(�,�E�P�z�DZGb�ݞ�PK6�ҫ�\cؐ��|*�a�)����5���a��I�2њv�4���$n˟!M$^����iV�O���L�vai@���I2�Y<.=��,��D+w1,�"-����FSA��6����E֐WI�$�|F�Q�h��� �L�O���?=J�$#�:OFr�)�&Fy���F��,�xC=�KE��Fy��;-�6�C�Hd4O%�ͣ]���TO.��6
wh�xW�g��N�L��9�m��Zn�V;�wM�6��^U4�?׬�E!��R[��+K~�~G�o6��jhA�m�~LAְ �F�w{=�<�z�*��,m��ޏA}QM�W��/��"._Om�JJ��Z�P��xͩ�k�K�xK���#��U������1wo3*�y�cY�c ��P
U/�`ŌJ��R�����=~&0G�qN^sk1��\
T<����`bq����������yY���AVͅ�9�ұ� �����[Au�O},u\����ĜҪv��m��B��ԗ�M+�Q�����L�hbw���L�h�W[1�_L��W�Vۮ	D��=��7���_��ό�`|�?���+��+�yے��S�fyy��S)O�*�������^z�p���a���K/��W��e��
��Y�𷴆�����fg���b�rլ�e�������Z^]1V���K��⢴d����v����=iݵk~�b��5�}f�e�9��i(@[����-[t����ez����[�ϟO=�����ss�z0ݹsWسw��{o�{��t�M�Ợ��"�4@�� `��o^_�r�� ���cǽɃFWY�gf.$�����YI��Q:̥��F���J��n"a.WQY���F����y�dyޒC�D{c4��4key!���Y֐ی�HՎ���yt�ɂ���3-d��"���h�����9��N���.Ƚ�(�NQm	a�3Yċ����V�6�E1jgY#S�Y#k���Ei-�YCޝqA1*F΍"	�"�a��n��._�X������E����n4tN�"�(�߬,�E���F.%�C��E_�I�GA���-�Y��g4*�L*!�6<�hH,G?v3s)��m
�Y.i��Ǣ�%����3k����L:?��JL�}1P�yL�!Dw���K��*�y�]���mk�,:F}ʟY/	fw���}��&�=��D�e�?O��J@�ݚ���,-�(������ܪM��ĸ��������g�tt,�빞/\��>��qc���yc���,����Y��O���`;	Z�^HT�8y�����2!��X��Ñ����F+8x0�Y3\q�	^�:"���t�`P��O<Z�,,]���U��ҫc���U,5F�ې�����I���/�R����Ltm�T�.zM�>+z�����Ȧ0Vi�4���T�;vl...��~?]���6����v-e�������/y��ʵS�{da~��w���ۺ�����߁�}!�@ /m�sp뭷�>�`�u��dv�T���;����\�0���C�-���ES�M٪��Q����������Nw:�N�f�kk+E����F�ΨH�`4T�4[�a�ʲ��e�N������ز|�!i'IҒp�F�BgMY��C�@˙W��a���(�I�����N��6_k}R��{U�L�6���~�f�E_[����huZ�zɵF��̈�V�/��F���ʉ*���ʤ��%��\Z䴚��F���7)����c��C�����;��\37���͚܌n'�!A���e6s�T���(�t�0��h%DJm1��MJ��6�r�_;
��<��.�������]H�>s�����p�}X壿��o��oYnc��J�+��'O��z ;vl7Qy����کhay|�*��Z�W	�+��*�˜�7�� �"?�D�hm� ;73mVj�%7/�|(�E��7f�.˖�b-k��T%�_�w�]e�(+�>C�*���}.�;Yh�fw�����O�puu%]__;s��e�^z�%�>==�SSS���(��Ԃ��E0  @��"0�2dM�u_����ѣG�S�N%r�{r�ېķ��h���5�66�(E�OYȓv�K�B��4Y���a�-���[BG�|a4�
�Y���e����9�*_���&ic�����z�n5���.Q�1�%�+Ko����7�l�|aG�F鋮L2J{���l�j���Q>ZN��B��<�&�p��G������������;[��u_}�QГ ����g?k����[͂}��-��|�e�ܾm����b
1�?���v�5W)�:�3V|�K)Hqx&�hZ��?y��p��y�V�ܻ�k���EA�Y�cA������T��?���T�Ĭ��hi�15��<���Yܦ/x�rb)�
�0�g_���F���K��^wM#I�����+�\�o��g���w���u-?�� x�O��@ ��s���ߞnݺ5ݻ�Br����R@ʃ��;��h�,e��ߞ��yb�ư�]����������O>�R��9|�p���YY���˂`E,�"M�^�CE���!�l�p߶}G���=�|�[���/�ܻ������=���',�,/��ki�$h�2��r%��,�^@GbYrUA�n�5_��(l߶#|�S�����%
�ͬqh<cų2�����<Gt��Y;�y��;�<�///M�޵{Y[?����_�����_�� ���8*  @ ��������{���n��Щӧ�%ac}��w�ގ|vϝ?�n�m�kz����S��b~c�;���۶{b���;w����[P����Z@J��������}����\�"�NO�v��D�W�p[���W�KKLO&嘮O%{�����%�'K[��]׳��@:�&}}�~���.�=S�|����p���e��=�u^��[���~��i���܋������   �$	��������_�8r����_��U�ۻg�e8}���H�_	�X0�JG&_��S�l����հeqф�`X�F��4�ڳ��Y\-G��y���~��)�E�J�zF�f�ҠT~�[g��*�    IDATj��dM�o����\*���������p��3e��{.nc��zvj�I���p�`�W�a~a�iQ�n����?�����w���/�ہ��   @��H������W]��z�C׭����ΝS�B� �VW��U1�H���U��zؽg���]^]5�l	������7�(!W�Ç���W�]��Z^�R����φ�U��lԡ�̻R�Y�X����{�*KJ��Є�$x�_��J%������r��!V'tW��Z��gա��i�V_/PQ�1K���U����|zz:�ۍյ���}�g?�����Cޗ���9A �  �$������o���o����OR�������ť�&t���Ξ=g��JC�������׭8�\c��-[�����0=�<�i��W����L +�Ī���*A���_>fg�Cwc�,m�f��Byn�+K��TS���&d��bK</n�~��;�;.�٫�X��ڜ�/��O�ޤ�߽�]l#�B"*��\�y�7ff���­��z�[���?��[��'_�./�Q�  @ ���n}�?�����oݺ�Q����|J��;�7..-����}��s�,{�
+(���ʊ��X��gf�ov}m�R��:��ewP��ѫ���7}N>���h�Vda-����ga떅���b�˗W�T��$xU2\i┗Y�n�Πlk��EB�_+7=ZŷO�w컱����1K�_�^g� JK�hq�J3��g� �o�2�ڠ��,���)Z�:�N������}�9������xѽ�/�!�  @ x!|��o��[o}��R��;u꤉ə�١�J��W��ٳVnqq�	_���+a����l8�B���&�UiM��
�������*�m~�f5�-`M���O�$�ܱ]%��w�I+c83�kn-C����"�ʠ\�r��O�U�)����󰺺fyx%�%f�Y��[>�`gkW~�zy%>�_���w����V��f�|�����s�������������_�q�R�@�~)��  @ /yoy�W|�[������]�p�� �����K�_�Ғ�W��KKK��V�rO�~ڄ���\.�;��}{������lu���j�ʯz]Pel�hdV�ق�Ҥkk+�����V�|s�`&��>a���� [n��(�3��>�)��h4T�m۷������lY���7T-p�}��n�
v�G�T�^�D"W��d����1����9s͐E��(+m[����H�
ߡK/��k_{�7���/����   @�eE�n�q�Uo����?��|fkž�]�v+�lz��/�*�� �������رc��,ʰc�sc8q�tX��l���|qێ��뇯��׆�ьAl*���1KC�ŋ���T�N��}��y���	W//\ZY�X$Eѐ����t����LMO��K˩�_�,lyu��V�6�[�����^~�,����:���,�Ibnr���~*��Rw���y|ǎ�ǁ=���-��������b��   ��	�y��c�u��~m�H���l�v����,��t�;����ì�L����Ç+����C�n�ݳgw8t���c���ի���!m���7�l���DLG&���'±G6�;�����z�^黛�2��,��(7��<�����ư�pvv������Eq����͚�{��-��t�z���T�����\KץJ	<5�����F����m�ۑ#G��?��O�D�Ab�����4�   �痀������6��_�m����o9w�l��
���E����7�w�u״ґ)PMY��p�5ׄ�����f�ݻ���j��۝�p��W�$m�?�	LY[�/K£�	O=y��|lc���j3�"�,K��n�͏V�W)���ݓ�z����RC�U���W]����;���}���15��;b�}�!x��x�i@ � ^��������־+�^<��n�}!�+���z^�o��q��?/1��Z���뙛��e�5����m
b���a��u�
O�$3WY|'�<Ν=ڭ�X��rk��@�C��m�:V|B�w��zP���Q>�*�U׿����[��|�ϗ~f�/�߄   @�eH@n_��Ow:s;��͡(�>���I��nwv˖��F�ۘ��O�a�ܽrT�L�4�0;;�GE�k���c�nZ�~5�[��<��p�������Rò��,�2�ʏ�)a[�3��6��lҿWAnY�>t�-��ķ��[���pH��SB�~�i �   ��+�:�pfjaa~feem�Ә:�5�WdIv�����<��4�23;�j���VVV:�Q�P���������5Zf��J�5�����1�[䣘w7SڱAh�ZV4BAn�\n��|�%�Ub��[�"�h��y����W>��w����r�/��_=�@ ���H��o�=}��Ls}��f�/O-,l���jLu��Ő���$y����W�$�)w�v{�̿��X&X��f#_��=�"
Z��U*2�+��!��exdo^xB?%��A���)�B8x��Ƕ����}�{�������z�޿+)>@ � �E�(����Dcjj����ص�����<==s��tzf&��VtBb��A?��E��3�m��e1�������������d�xD���[��J_w�u�`˖���w,1H� ����   |���{������ݛ.,-�`��y����r�Z��3(��4����҅��qA>��Ao\B���U�wg0���hI�b����*�ɏ8\w�������<�����/ۡ��  @ x!	|��?7����Ϟ>�}����NMO���ZtI0��,p-���Z�V�W�Wi��%_�~�?.8!��\dٕ�D�����v:����_y蛿������R���R-��   �-�����ei����K�0˲#�vG&�4W��4�;���I�6�4���X����+Q,Q+믂�$j%��RК`�b�=���{�^���ݻ�<p���|�C/Z85����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@���� ��E   IDAT�u@ �   ��	�go^J�a�    IEND�B`�PK
     #{dZ�  ��  /   images/b13518ba-21c5-4f60-a735-1d8041d11d7b.png�PNG

   IHDR  �  �   �lC   	pHYs  �  ��+  �MIDATx���	�m�}��}��g��{�M|��$Se;�58��Īb;M�D�#"���v�N�&�ӊr`'�؉I��h�6���7�[���R"QI��||��<�i���k�s/i.,:���Q�;���k��^��   �#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   om�����^��f�m#�  �I�z���'�X+���~����������޼u+�0��mc�6��<�~���~���7~�����_ϊ"�ײ�gk���ol���٬��'�|���[B�  �
��_���֭�'��_o���t>����Ai�6O��㬪�&��\�W�7R���e?kB��7򪪎���h�յ�?��ß���?��z3|Y^  ����3��÷n��=G��?d!�鵽��ˬ,�UQ��~��/��d��8��:�ě�Mo�x�����<o۶ʲ^����,��(&����x���������7ڿ?���"�  |����?Z��;����U������*�z�q��ZM�/�(��i=��Y��]�[P�BUՙ�ۙ}��{=���Q�������e��%^  �ߦ����_<<����B��Ъ(���An��Q�BS/�'c%�\�������g����Z�/ϋ,﩮7􊢲/���~���e��!���oVWV������4���?��K"�  �6����g�I��Bm�����r��i�[�m���c����d��,����&+�V]��U[�i������Mn�lgw�/)���+fs���   �M�鬧����l�x�f^P-��=���IUƐ��zv��k�)��~�Z�f��z���|6��,/  �o��yV7US4e�_��N�k�xo�f_h��w����(­�H���ח�*$K(}8y�V��������?����w~�w��W3|A^  �߬��SO[[[Źs��~��Z�_�{��j�r^ͳ�*��,s���WB^U�n���+vn���7�W��!�?{���Л��vM]��.�f�wX�^��Ex  ���~���W�d�lw688�Q�$7��}�/6O=�6�[��/��h���'�_|Zӈ�f��jl������ܞຩ�����tBl����\�?TM������}�������i4�o5���<�g���  ૞��2�qcp��-6k�hi���7KK�j2���٬͛���;�o=�}�lv�eg���O��;*bț�ݫ�z�כe����ŵ�W��GI�-�N&��l4���J9�g���Tڛ��I���4'���ݪ��S!�/  ���҅���F9m�ނ��ۺ~��ҷ��m�մ�-�֓��e�����6ͥg�����Q1)�v0�NV,�Κ�n4W��djwSIC���r���x�A�7y V�}cϰ���r�DB�zz�5F����+��mz���	^  �U����h��=ɧ���7V���l6����b�r�͎����?8�c+�;�yu����a�w2�~�Eэ�n��ӯ��e�gYӕ��aV��{Ku��泬Q�-GY^�ƶ���e���nz�}��ƃpS���|���/�?���a������~����ֻ�y���t�Ak]������o�u�|p����}4���Ν;���J~|tT-�,[+j����ٶi�)��O���G��۫�������������� ��zO=���p�����������Yx=g_XrU���fVգ��g�����h)+������;��㦗�%�|���R�n>>>��,{(D(��g��d�z�S�͛�߰�:��h�ݽs'[__˪6��ka;+����`=�ا0����j�ťKK�d2��~问}���2�&�Q^�����������������?���]���d*���������|X@A����V!7;::�,���Y;h�4�hgw�Y�X���[ߡ!���5'��KK���Q��<�=�ю��μ��t���qc0|�v���yu��w�굳g7�E�]U��+�i�=���eo2  ����|$?�^yxm��3�#��Ł�a���8Wa�J���PU(�1�KK�����zV5[B�ܡ���d�[8��1ΖF�L�������y�Ӫ^[������R������WYD%3�^ӫ���-om���g7S�qv����|ns���������7��n�������|4���5��᰹y�f�՜I޲�Ww=������ǳ�<�̿���;;��~�e���U=����0{lavTE�_�rn�B��<�u�x����o�7�픃�0����7�m��;�ͼ����{zt�է���}t|��{���+n�f�Zb�֒{B;�Zj֚S�nf�i�!
�O������w>�?{���,�fmu����W�.]��F���2���=*��~Y�>s���t2}՚�;�^{+���v������?�Co���G���|Ŏ������-�׍s��(p׿y������ �Uɮ����K��z��n�X]]����Umn����a~<g��;�p0���72��f�o���e�̮���77�fw������t��-#e���m����3�̠̠���x�^��/�ij\.b@+B[x�p�����:W��`0X�498<x��>���[h�S�ᰜy]�L/��n�����ן�f���W��=�y��f(�+p�c�Gu��?����_�/~%+zW���گ���?����
���_��}����Ɲ;w>�5�K��G� �l������Z;�3gΔ�q&�
h�.--��յ��T�«����V�d2����t_�gZ��s��l'k�ժ��$�Cm��N��d�^�\E�����~�M�w��W��oŶ��lln4v���Z�y���奕\j�TV�uo�w���R���}�\][Y�Lf�kCA^�~ǖ�YYY�4)I���>j�{u|���vs; ���+���|}^ǉ�u �k~��U��wfٷ|�F��o��������r��g�Ｕ�8� h4$s||�����sc[/;��t۶ǡ�B��|�(�;�|;���֠_nU��`0(�Ӊ���F���͢>:ڷͳ�\��yW�T7n�h�\��~���m���w/�G?�TK  �Y���w�,���eQ�X�X�'��ں]iu9-<SL&�ll�T�Ӫ@����׽�=��욮lyw�N����=����:��gh�#��J�_��g[��5���RM�{���@��!4�5����$�-�F��|f�?���eZ^�"������^�>V���������G���+������~��o�r�Fѿ�����ǰ���S��~������=�ؿ���W������/��W5��'h4�;[����S?rtx��1��
�]--/����}����m��6��VWV^UF����ª6�?�ZS�h�hXB�p�Zm�����ڛ7ox�T�nU�=���j�PJ_k��k�hH#WX�ίC��󐫲��`�߼y�_K���F?�@�{ܾ}�T��}���p���̛�4���>G?����M�[��,[8��ݾ>�5$b�QP��������8�?��t����W�ּ�9ф�^�W�W����U�3��|���,��6�Ѱ|��K���K��Ȟ�yĥ�b��`��]����l2�����F����ʹ]��a}V
��x����^���\˥u�����}�Y���
���+�-�Ϧ3��j8�5�8���:i�Ț8a�ƙ3�5`*�3k�Nl�ۊ�����ʲ��n�g�O�����R�{�r�k'�{�Y1����,��vЯ�㶱�^O���Z�\����hu���[i76v��͵v{��OP �����|d�����G~��۷�N���e���{[�w�据�*��u֯+���]��:�+�Z����]��>�E���;�߱���?OZSX�(U��/��<罯*wPi�����j��2�84���k��B���v�]V]��}/�pup�k
嚦�~����C�����V�]}]��������Q�E��X��4gp�k���v��C���ã��3��J���<}�����\���O����y��?���S��o?�C�+�C�n2i����|����F�@͙�3�ŋ�K�.U�Ԛ�3u׫��6�m�VϓVYCi[9����L��;;���ʒG��\;H�`����]�T@�Nt��h����Y�����zB*s0���gtwwW=���;;;�B�\�v��p��x�k���
h����C����*���Y;0tz�܂�����F��i,
�^/��@��kGU�����`�֚'H���k}�Ν|�B��>[G�Ϝ=�ˡ`�K=��/ߧ!�|پ�ϧ �kk�������Sdt#���¿
�=��z��6Z��g�u�v���z�ɵ<
졆����=�s��]k%?`���sv����j.U��L�c}�R��`�@�7j�2��<=���.ʰKס��N8�\�g�`�l]'�<����`0��e�G���@R�I�!�o��m���������>_9��`��U������s�e������F"b+=<QGډ����!�g>yx�����NB3[�֖�f9(��ر��=;�G���|��k��5�����e1<��I3,g��R5NڪZ�ٲzy��S/�G�q�������j{ܠ	��SO}[���_l<a�,��S---��AL��޽��2A����E�f���k�%&���� g�����<�ݹ}ǯ���|d״��N��K��9ш���ƙuz�wKu�Z�!�4qF�N�3��[U���m�>���`>�t-*u��=�N=����da�v]�N{�e��"�&�e������&��=�vͶ$��/�K�o��'�}�G�ҳD��^����??x�\��eǫܾt�^u�?���?=�Gkk����zr$�o��o�X �l8�2���zGU��e ��-���V�a�S��A��]�����*�Τk���_~��L��
R����B�Zg�A�a����0�]�ND߳X�֭��0�H�'}O;�>�!����I���r'a'�eP�;�?Ph*�8�^z�=������X_W�To��n;z��R��}?$�,[��(��k���^%���F��}��K�E3��o�;��Z`��n����u�C7���f�jh
��E=�
�)@��˗}�=�&�{�%�@[��D�i��R��Myhi�g��^��w���ݬ�y� l�:M��tOu|�����˯�@�F���Nj
�
�z?��n�����C;��$�Z^� l���9�󕕕j6�ض��ZFՖ�a4��}��z����~Zμ��^��*G�5�����f`�W�Jhp�g���h�{��m����=��^[-p�R��o/ڄ�L���_���g,������}v�zٿ��wf�K5;�~���	N-
�e@^*����Vi��7F��c�KCv�f����9��a�m~�6�~�k�{�5w�^{�~u�a���~�[�o&֒�l#�hTU��ܚ�ڰ���a]j�<�loo���Gk[&�@ڭ?���zO<��/q���nj�V��ƍ�����u��n���3�@�åAs����u��n���Z�S�O!uem-�X��D]�Bn��묮g77��x����]쭏f��A뽬z��ŋ��۷ny�,�گE����5�����zO�O�m�kr����놏~߻{����/�>#yu���K].�Ƕ��pWGX�#©��Թ�^���,u)�������{~V&Q����fŲ�'��w��?�goa�c�7<z������]�z�+��ї�������>d[j��C����=���{��^�x��֑zG�m�S�_��Q�廟x�Y���jc�Li�sptx��d��F'�tjV� ��"s������]�
C��rM���7|Y��^[{]L=|+ .�F]]]�҅���Ǟ�\|����{Ҵs(��z�L���<��*kM���li�d�i��v PY��·|��>{yjv	m�M����ܢ�[�u�U�hZD�յ��a�k�c8Uֲ�T����g��k�(��u���~'�zC]o��4��;	xT��J6��p�<��f˰���TC��Zh�ȧ^S��������I#O!6,˒�Nx]T]�<��'>�P��O���V^����(�$��캣6���u!��R�]om��t潣��k��^ʢ�W/�zx�84塾V�x}����C�I㦊�a;.���^�]���>0�����s��A��N�<՘�9�xJ'E�(`����5=[1�K���ė�i�x/��[�;�1dǓ���dg�N?~z=���!Z��A����9􂍖�ΝG*=��X��h��sȢQ��|ړe?�>��n.=�/�uh,�2"���_���7~��Q�n�O4z��1�ʇ�>ի�QjD�+���5�T�f�����S0W-�혽#;0���C���-ˁm�[����+k;�Gv��7yy�ֵ]Aډ��qoП�2u ���Zi�~V��Ю��6j���NG��p�N�#}�fi��V^c��jk�Y[�/�9�\�5�/�hϞ�i�Od�<��/<�{=������+��ͭſ��m�[+C�>��p2Q�'�A�l��(;����l�7�G�����Vϛ���k�<����ʪ~�X&�7�~�o{�:7>��������Ǜ�l����ύf�v:��G����ht���~��X��pҋ�-��h���p6��ً?�u��N��`6��{����?[���Sf�|� }��>��n�\�ˑ}�}�A;��b��I�ŗ�d���������x��Zí�z����hmۨ$���~mڶ����rQ.���ӷs���Å���j6��&���Q~�Ν�������U��6�p7�s�nJ��;�~�[_���^}]�eG�@������B�v���]�����|��9s6{���|�j�������ݺIDm�vm�lvəL��S�׫/h�s����ڮ�S�R��������>��x��"L8����c/��K��E#���d:�k|虾sw+{���s�������}zx�c���{޾tns4<>�ٰ����_�C���;,��-�>����c�|,;�|~�����^���4̬�������{��M!:5�E6�����A���w_So�BV������ܹ���x�h'�x��B��4��;/����[���u�V~���|��f�;2��~��������W_������e��m�.8���
��S�������=�+��@��]�5��z��c�a��\=��bn�Ƣ�>Q��Ϫl���S!H�A�⁨��X⯧��%�ݖE� �4�љQ��/˼5�P�����5T���3)+P�US��H���=���4���e�<-��q�׿��O�iOX��
�)��=X��逬Ю�S5Tt�����i�S`����i��ZFՆ�v��P=�gϞ�bi�Fr�?!ؗ^+��p���S�J�6�u�co!�~3�����Z�:�����"LK�]�^ �稆��2��y��We
�ڟ�?��F�C�Z�J�!�嫞�ڷ�\w�wz�PH��^S�[ˣ�t����Ν[�?Z�0�I�ˢ��5�-U���w��i����8P��֥:����M�N�~����'��¾����kT>��z�QZOZz���ԃ?����qR�+������,)��i<ݐҺM_�>�I���t��Ok|g�����wSǹ���⢥�'�R���p���7��gZ���(��k
��?�T8g|��S%Q^w��֫�le�f�sϏ�&\<_k��4�G��8<��Tk�㣱̮2+���C���lZ�hZ;i�u��m�FC���X�J��X��f�5\������E�����Vu�m��]4��� ��7+zŴ�TX��	4o���IQՅ-�h0��~����m�ׅ�O��DY��U~��l�h������lP���t�����>泽�-��R��
{�fسw��jM�YQ���O{sk�i�򺢢�E��X��W��04����h�Q6�-�,��iE�0U6�-��zM3�UYU̧����Ӄ��W�Zc��G���p�{VG�dz<:��e���j�.�k3=�`e8��{��[�ɏ}�G���U��ٱ1��u��'[�v���hǃ5��z2k�̦7��q�Z��Rê��6���6�O֨�k��Փ���onY�>w��M���n$֟q��N짞���������_k����^�u�kUϩ�q��V�����Pݨ��o��M?oZv��aP��t�޶�c�Zh�{�nv��,��
������<��*?��`�e
�:����xٮ�:g��E_ޢ���Mm�x�E�z���}��z\7Ξ�nߺ�Y���x�UU�!�|3�΁�,�|�M;�Z��;��5][ԃ��8{�Wl]ݭ����[؛x5݇������+�����[�ް����ի�߱���M�����������wd�{{����ZX~�v�#�����ga�|e�/��[�HK��:���Tb~���1}��,�>`�R��h��T���Y�'�.6?�?�kR镕����������677K]ptq��������vqU�TX�0H�M7j����S����Р���̃��o
M�����Gٚ-�BT�I.L`��TI���g?�Y�W�/^�ϧr�Tޡ�l��B�&<�PaU?S�d�u�����{�z�=oZF��omoś��x�����3-�NZ
�
���!7M����&-��kZ���4��'I=�
�!��_W7;�eW����b�ƻi�$�ƞY}O�@a��'?���z�0%]�_ײ�w��Z/��C��ֳnrX���~�����k4����������P>��׋�/��AK��Z�z_��<��%۞��b�y�D��7x/���?��;K��!�R���*_'MzPx�Ի�&AW �6PcR�e<����Zư���XU�ƕ�᳅�ƍ����.i�FL��"9�7s�O����ÁOѣJ�~1Q�@���s}�.6�Imw,[񩆴�n(��z�t�֍��M$a��d��QjP�z��ު/��'�6�dFǺ7�bX�bϏ���+)dO|_������Ko��Q�آϛ�#�2���S/`i�0,�2z�U��������N�q&[�����u2_K:6��X��r���~F����#D�0к�s\܆���:7��L�Pu��F��ױ�-��3m�,�M�S��7\�9)��d/�-��tПv������>�dYx�)T����y�r;���Ըj�6T)���C����׫����M�&S�J߮{����as�������(�y8����U�3�FeQ�m�͛��p4·j��m}��W��GiT��.�Ւ]!�H�땦Z�W����h6(f����}֨��<p.��T~6�k?��+?77����%��R�u*��x�-Ν~ޝ�f��Tg�:�����sQ���S������Jĩ��t���ʶ��>�ܶ��ř�a�Y�)W�M3�Mgc;O�'��ض˼�+&���^�e�l�_���z�/�ǣ�5(ʢ���{��Y�������ѽ��?��O���e{�Q]����w�����.zCUYD��>��Ғ��};g�!��\���S.\��y����^��5��k�^����ϛ��s�ƞc�{�pX��g����Fo���y$^=���o�G�y3���^�L޳����ɾ�unq_��o�-�[�����7*���5��|ue��r�w|�������OngoAoj�|�r��ϖv�>��s/<q�?���w?p������)Xz��s�=��d�Чq��i��6��mٙ���ÃR?��N�
mv�kbU�`��;MLG� �a؞����d�Q�a��]���	�NB�:
�*�Po�B�vv�"hH[?�״ךF��J.�Ë�K�`j���Ԕ"^�z��������=�-����(������P��=�}�%�:�ؓ��)���7̾�B���O�vN�y�M�EP�8�R�n
�
C�����S�{��K�hi[�$�C�v�N��Zn]L��T��?u1�����n�e$C[�TG
@Z}ch�xAN��0uJX~}�<����Sϥߐfj�*�{*O�.볅p£�h��!M��7��xE3Fh�J����z+���*�IR�E�JU!P�YW���S��^�>�k_��r�n�X#�ϥ}Oˣ��'>�Ҷ���G����}ݶ���Xʱ�lZ�cR�zZ��� ����x��:}b�:LA.�:���C����ɔ�:٧}�P�<�}�R��|�>=N\Z.�ꩌ���v�´�8�[�z�f*9]Ýz����}(�ظX&���y�k�}R=4�N���X��+K
���I7���9��,��./��xcdK==�KqtF�S*��c!��7.�K��^�D����s���-6�I�%Yz�:��X^�b�o�f�^D��,����Ư��zzuG�F���ì)�b�$s%���^˩�;�}�º������b��m�v��Ξ�����֫�R��w� o,��[��*��B�.b�Ow�k�N����t.��~�T�Mׂ,��~Vewڷ�N|�2�1��l�:bA�K�4�����`����:ɨ�>���j�������u���f�I3�����a*�C*J��d�=U������c�k�����,Ko��q��U��a��x`�U������Mq5���;��^��]�x!�Y��ͫ^�wo{�;kf��I8�z�Y�O*k�WN��F�:����Ѡ���M��,�_g�č���`8���P _]9�8ZZ���Uu�W>\�����ny���gׯ��]�t�υZ���\��G���%+���צ8���F�λ>JcǺ��Օ5o��u^ZU�({��>b�O��l:	�A�á���h�%\�EG���(�k�2�*�;;�'-���k��H�����~Ly�U�V��LI���|�C����õ��?e>���/ފu�oj�={�_7�?�����~��X-��W^�[��+WF�����I;س�=��b���������^}�U�@���Z,־������v TK�`k�jԍ7
ӈ����
m:�h����NT^{p��'Le�9�d����ð�@�)mj��F��ի�� �_��_�/�wIAp����on߾�ꤳ���l��<�
,�f��p���^�u���{T��.��,$[8V/oO"�㐲z�ԛ���iBv,��$�n���t���l}^����B��G������^�rٗMR�j(�X
u���+�� R���3g������X�����&�=(:3���P��4oy�3�G'f
�j��B^����Z�\�ԯ�z�x������FL�M�O4ڏ���룿� ������w�?�������Б���O�Q��C�V�b������GK�<�k��'�T^����E�~Fvq'l&���z�N�k�nݺ���Cxn����~��/o�Xd�E����^�12�]id$� �3MMW��8,��o�0�=*S	ʪי��>��O���X��آ|�,A�?g���m�!�67N��_����;�&�Tc�?���-4����,�t�JB ���I'j/�-zHO.��B��h0��JJ���F����:�<.w��zī���˗z�㴈Y
{��)���n�u��E� �2W��y<���������a��b1�H��K%L~��p���4��k�}|6��)��eѺ�q���T���ŹK�����0b���c���˴��频2����/\�ؤR��˫�]�p���:I���oW�#PM8g�͘޹1�&�w�Ӻ	�V�aw�O´�E#�v��U�S��Q���Sǂ~���<�@���.��E��okk����M�/4��?R��W�d�̦�ڰs���/\���l{�:Q��^O����ԍ���;NoiT�,�Y��̏���}�d<�o��g%��j�	K��O��_�z�l�-Νj�k�L������fב�xcVQ�#�;l�u��u���z�y�JSs�/a_׺����Y��GZ��Ml����"�~�4��api���i2����ꩴk�N25�l����gWy��Q��&3?G�q���0����p�ѳ�׿w�xo��0��s��ѵ�	�65켬�U몪C��v�����������c6fH�����5�pi�/J�|�N!�z�eo�4H��^��zx��.t�y��c#,���s�=?�iƲ�虧���7��~�/��_����h���>��3ӷʃ)����䓟���ő�����|���M���ֿ����y��K٧?���I����e��~��ϫ��o��ڥP�Y^8w^;V�D�"�^�Z� ��cvrZդ�
=vQ�4��.�z�ّ��y��FAHñꎿq��~+_�Bq�����P�·n�Ց���5�t�bx^ʃz�;==������A�N�]x��<$y}�}���yo���*��^z�j��w��B�-k�=p*�*d|�3�Y\���w�ν������|���}����2��L��؂��Q�Z=�['f���-2.��^/��Y�լ^�F� ꤥe�t+��b8�O�#��7��sj��� �gv4�3]�p��r�pL�'�xh�r1�ً3>�Z�";o�]aL'B�z����t�J!��g�3:��*F�?�s/��.��t�K��ԷeхFu��	9Wl�$�Y.�K����RxJ�o��ç����׼�A�������!�pTOp�e3<h�`ɾ��g>��VￖA_W��BR
���F�P�P_�q���<��t1�{�����m��c-C(�Q���_Lg��n����~�>�,4'=�����l��3�Ts߯�p���4�3-�.�jx�ѕ0u��{���=�E�C׋��`��K@�����|��=?��m��c3��bq:��^BzG}��8cI*Yx�>$�~����I�j*�H=�u� �=���i���Ϟҏ�w�X����R�tSlz�r}�E���
q^��=Qy~�?����S$*X�a��T��4����Ǜ{�h�s�=��T���|
}�~��Ҕ��g��pt����w�Zibi�OU�כ{-c��=�&�fִ��I�V�M���Z���k<�s�]�
f�Hh��-�f؎t2�ci���j�_ͨ��kD�=��o�/����E��⥋�vwv�5uD�>O���J�q����l:��Ԩ�yR��m˘�ȕy��`uQ���d7.{��ꈽV(��4�̭x]�����!���5�u}Ӄ�,�g��G^�����+޸�y߽�UǛ��>K�ܷ�,\�.}��롞�����SE�횽`4�ٹ��������7G:w���F#���/���r���k{gVJ��f8��`׆�����ً3	���06d{�8�T��A�Щ��R�F*����m;Cb	�ɱ~rJ�
���rx�p�_�z��{VD��p�iHei���ק�e_���ܧt�3�}��;:U����-Cͮ_�~fk�����~Ys�?������ޮ]o��S��-���c�Go~�����a�#7�ي��ȏ��o�����|�{�����~�����r����	Uh�<������?����}eeէ��2\�'v ���,-[эB�]��l�W�����g��qc�ñz��*��_{�5�F3.�e<�)�gO��	���l�+u����������K4w�nXe��'�L�a�U��"��vB�3l���VQнs��7����D��"p������&����ʕ+ޣ��jY=p�ƺ����P���~�EH���u�ࠡ���ʕ�f~!TN7�h��6R]�JO��/�^�>K�Գ�^j���>������	7ˇz���.���^��[��Q,IH�d�*gi���$݀wzhT�A�vP`T�������FF�6&�&�����Zq�:秧��z߲��^�k���C7���}��M�}W�j�ÂZw�X������������v=�j�脪m������?�r���'�𰩐���ը��_�{��|t�(C��5�vo�K���k�w|�wf��ԧ|��τ*���|U�<��:�ҷǁ-����X&���򗁇�����׋"�i��,�b���i'��*,��������2z��wn�2hY}z��Q�-b��A1����.zX�8$�����4|���p�Hurm,MHe�ϰ_Ws�	��o��A
ۗ��O�/��7��S?�z@��Y���`�u7n��r�´��!4��+�����kR�a���e���4�P
ӄ׉=�gR(^T@�龃8CJ8O�Q�S��xc_��s��M=�>:�@��ZE�(5H�݃��h�F����'.f�y��hAZ���L���=�鳝�?R������Ϝz�&���|��\S�h�3��59��O�a(�����5�n;�>w�\������������^X�[�}-�X��q��~7��xՊ}�p�I��q��Z�"�J���z�z�LGz���G@|��ҬG�S����z�0R5H�:���uGjB�sii�ܵk���Y����4�Nh���;/j���P��_�p1��qM*�Pǆz��������zGr�P����a��뭪j�����凉5P��>^V]�j����S�p�mm�񹺺�S�.����,N�Y�V�Zeuޤ�����554�c9R�ao�ޢ� ��P/�OE\g:/dm�q�"���{:�∠OY��|����ݿ����>�n�/n�tՁ���'�I���,�L�*�X��,����ܡi5Ká��h����:���7������?Q)w�=s���������G��}�7��Doz�m}nƏ�}�W���~���!��������T��=Ԇo4�9�0�؅m�\�@��ӆ�?�`�mۑ|m���O�����?���_nYtݍ76�j����o�1[�o�s�ӟ��B�O�a���`��RM���6�,����*�ܠ�����3)��K��K#�D�p*�A��f�~
G�~�L�a�j�����`w7���Uk/����x���ih�[�
H
��_{�C��O?���"�}��E��իW��vҁ���2�J{�$���e�^�س���V�~fgw'�\�'b��zb�5���B�.n�q&�4��!�4���~#K��N��>���u���ށӼ��Y�C��j�o�����x��dšv��?��gRo�/_�����c�z35|�ى/����Uk0�f�{[۱qΗU�&��u��K�M)k��'΅Ϫ@�j��Y�l�xhR�Nd���>ָ~<�춳��
�j�h���mg}F�tՇ���Ϸ���������~�Cpy�ԍ�M(�2��.�v�[��������l�{����	�a�C���,5:���Lge�Sc�Kl�j?W�O�A�]�z���q�muˀ�}Ɗ�E�b�/zC�,	U�����J_K�P?��rS�9�3����5>�|����tꦴ�,3�4"�P��YM(og�p\�a.C��h}{�y�/.,��gQ����c8�}���X����4A
Ⱦn�U޷sk*7й������Zg��4�C�}/�Cݡ�����9�{qyb@nJ@Ky����|5�Z�x�T��9γP����ң���K�TF�3��ЋJP�y*�ᓐ{�(Ќ�G_�Gקra[N��Z�
�i"��$�4�����W���9�O-K�<i$���ף�<��4�}Ҳ�O���у�⾘k=����NN��^���WG�-�p4����`�e�-�g��<=�Yy�*N�XW��k���j����+xC|3O��׍83�bV#}v����h�^K���E�S�c]'t��2�U�����qM�fi��u��Z�\YZUO�ȇ�/��Ӎ�>\7��w�F��5��7Z�䲋�/�yH�#���R�'�x����C�fo��:m�E�z������]�[��R��A��A��2�"��)�z�/�Eqj��GC���5+ܯoN�ſi�*n����=
~3o�d
N9i*�C�_�5��]޻w��lZC�o�.G��e�E��j�R�ؚ�W���ε�v����Gٛ�+x��������s�,;�������}���?����{����6w�wsk}����
a�5�B����co�?�ܳ�|i��5�5�c����v6Z=c;�߱�',����0֑ܳ�~!����[����(ֶ���ۆ~�.�8:8z������Ajg�l���@7����Oeѝ����'�t'��Q�eRo�����&�p�V�p�=��$���n�X�Z���}�{��:9�"�C�
7�9�ހ���z��\:j�_e$zʚN��fUua�,��߱���I�xN-�B�[�8N����G7��	���Ah�ۅQ!k�J1K��i�R���xײk}�b���,����~|�Z�D=�a�ǞA]$��6�LH:�O�g5$���f�:�?�֝�N�YR�`?>�yb'���O�##�;�y���t���UϹ_��w4#���W����?�����y�k׮�6���_�p��n�)h�E�X�Z�:�Ʃ��������K//jm�}��>��؋��*�Ϸ�h���𶎴}`�yE�OAZ_�y��"��k:��=��P�H�[�8N���R{�d�7��{�E��rORR@��>�������_|�?tv�Y���,(��~{33�%](�$o���z�:��=��n6I�e��Lә� �z���)���>N�A���\K{�5c(ܲ��+B�.O����S�ԥeN�M?5�N��Ƀa3rě�⍘�7@�ϖ~�V�4L�T|��7��M#X�҂<�P7�S֧fr�O�Զ��K�4Yq�C��������>O�/ͪ#xT���,_��'��T[��C��5�?�����e~��{����>_�nu�}?N�φ�ºN�Bi*¸��?_o:��=���p��#�c)Zӆ^>�Vp<^�ӝ��mo˿��ɍk�Ҩ���_��ë��ڷ����~|죊a��8c��w��i�K/�^l�?�dȽ��_.�}P"M'Z���F;��7͢�(��сT�i��;��>��:DO��9�gc�Ǘ��y�]3,5*yШl]Hӈ���z�h����/�����|({��+a۝*�K7��c;���i(c��ڥ�@�y��W�˛t�kR�R�q���ٺ/��TB���E�|c��j�ziQ�U����<Ue���6���+���"�T��#z�mg0ibGђ�����*Ubf׿fue�{Օ�V�W�V�J��k�����7�ƙ3��.ՙq����or��ޏ��ŋ/>���^�����m�ǋ����x��t6_y�w�~��G�o㓺x��kʦ?6?r�T9�.�ڡ~��{s������^�oݼ�Cۡ�/��/=x��?������M�8�w��������>��[�������n��d,�fG�M3�P����d�����v�<6���Ps�.ښ=}t��]��T�g��q���"�y�t(�̠Q��h���4����ׯg�iX������0�n:Jw�~zY2��.�:�]����$�rx�}O@���v)��O\�w=��+�t=M�[�k��O����Y�LS�LgS�S}������'�&�/�v�j�8���T{�S���9#�g��Q��eA�M��3�%~�p5����lt�F��EXW���*9� mM��j��6�Xc�;j[g:�鳫�F����ۗe>���#�� ��w��i��i�ܯ�k��y8<0���c]����=�y��w)ܕ����'̉��I��q��t��͍z��0�����я����O��=�xͨ�m�7S�k��.L������y��G�%�	�7�~zXI�?��N�8��=z^FT��S}M=����iĬ���@U�i��>ǵE�~��:�����=����pmxl�����&4:�z���
�!�����|رi7�itf%ֶ���cT�S=���{�^��x�b�:N�;֠���)H���ѣm�3,�^��ӽih5�ϼ������E��Eu��A]�4�v
G^�Tᩄ�t"�w��".��J_�<_�y���5�>�2�(k��IH��P�J���T!=-�d�����5�8O���+��Ѣ�$�<��W�MC����z�oh?Uc6�]��[,ch���NǺע�0�|qæ���m^/�A���&3��5��\���m�q���� ��X���Fc�Z6�W��C�چ�75�2<;��Ž)�<��G1 �M��.� v2�LQ��ԙ�$��r���X�s���<�h�)�)0i]�b�Yz�����G#gi&���5&�z�����T�WqE�K��e<��X{�������T�f0	3�.�K�(�+��G��]��ty�z��Nu��k��
]>�X��J8�S=��>����9�#�?�i�w�t�ZwGǇ>z��a�L��8O�(����f�qX��X��s����<ͦq���]t�f��ͼZ������0�r�6�ꉍ��$<��/V���c6��//�(boq/K�C�s?��|9Z��ry��m��M�]}���=�?��зյ��iT2<�`���|d������7}߯H��{�'�_���?`;�v��g�LU����l�޽m�iF#�^�������T�r�����_�������������p�m���g>�3
��p8ؾx��g677�l]�/���5��K�|�I]������W�u�褅��[[[�wxttk��[�W��~��j�1o��֒:?W�u[��Dtv6��_5��u;���oG�f֎Sv�|�.TM�]�K����-�X�(U��'�褭�����of���N��¥f��k�U�_������^�S����u;����/����&����`�T릇�4��y^���i��b���x\��G���4_f�}��{��������X��3u����p"�g'���:��p�+��]��G~a]ZY��>�oo��i7�ז�~,޼h����Lei(=�(�Z�<x��-�I�5��4Zjz�����BO8���}�s=���T?���O���2��u���ڜ=s&WӉKӔ��['�]�z��ᑇ�6>�lo��C4M�Bp��M���M;�o�Os�څ�. �d��4�K�����z��N� ji����q:�0r2YLI��LAV�5a���������
�?��0�F�Z�i��zKfވI� u|��8�z���>����v�0s����Z�aj�P��!i����� za=��Ƃ��nj�ǯ��c9�Ɩ9�$�@?�!?I�G��i��R-������x(�Q'=�1>v[�'�N��W)�����H�L�������n�Ұy����j�/�ZOa֚c�)<�z���	��r��R/a�=5�Ҕw�O�i��<�_U�Ǜh�0k�b�t�����Yf��<�Sk:.�?+h��~�È��Ã\TG굚�}������}�Nx�Of�9BC���������4��0�@��F��p�r,'�73k6��;6��z�4B5�fa�����"L���W�x܄2�����l���\�;�1͋PJ��~SW�1�z8}�U��*uO�}JSօ0\���|݌,���^w��H�lј\^.c����W�Q#n��řw¬0����E�|
���J'���1�*��qs��㾌��fu��7���8E���7�@Ϯ�[���p�\����9{��}����p�"�i],��4�G{��7���ł��{��L���N��i�[����ec;�i���{���Y�㩝W���wըn��w�W$�N��7O����[��*��:ǫ~R]�z5�76*��~������S�h]]�
 ?��~2�ƫ��s���/��ľ}�~࣭��AܟxS�e�?�{�f�_���3�.��������N�v���R�4˳^�ԫ�%���|�-�����;F4�rɂ�Y;�k=^��|:#;I��gRǓ��(8ߤ�n�y(�b�!r�7��ԓ�z|��Z�:ع�PQ�H�S��YMOǉ�!>�z��O?�XA^�_�~N_��B�=�i�m=�U�r��Z����h��YY[���4g���X�^X`,tr�3a����·>R��*��kě2�8�Yx2X��-�"ΙY�i��~a�J�c��TU�Qp��$D�gni��fP�k*&��$���AM�wY7E�gS��w��w����u]� �O�K-�z�Ğ��?��\ܬ�j��v�T�&H
����B�����wa��T�aL(5>��PW'Sť'���>O?d!�P�BT�6,]�ROc�b,M�������M=��җ�����O���0�9iz�4[F�S;�����S��y���,�\��
��{ol�u�	�Ϲ�o����T�R�ed�m�8�1�M1V��h���p��A��?:��#��+���S`A��*
n(O�O��Yʔrz���;�a�^�Z{�{^�6`)�vq��~������[k}�[Pq�c3V����j@�ʼU��)�}����~�6����U�	g99�¡M����<i8���2{�q|�Ț7^ x5�TC�]1�J�Z��J��Q�ٲ�b�`X��F�~_�)������)7@Pˁk!����W�f���֊�/�}�~U�7���0P�Ds�ה9�[�f-..p 	X<����R|�ڞ*q4s��pf�	1�:x�G� 4�xv��]&��!����mܧޯ��80�5� �h�U�g��'́��y���e;O�Q[���*��yJ)�R|!Q��R%8�34�N�h��	�؋�T�-�xn����&"O���%SiN�89Wrڕ�Z}��Ca���8.�\�����V�&T�G���=H�2fRWZ���"1�%�%P��W(ϗ$�c_t�!�ײ�,���I<8��'f�ֈ�����s��Q�.��K^����9������׆�7I�=�w&_����y��uF���L)@~��Qs�˿�y��_�ܳ�xP}�?ŋ��ܜ[Y]�w'K�^��U]��k�"}@F�+m ��z׻�y�q�T.._��n��[��X��o'�h���آ��Y����;�^_���M�y�봉���:GR��Y��~# +Z	L6��bm��@�c/;�@�W{�L�#
δ�P���mӵ�;�ori\�p�*[*-լ_�O�sJ�u�zI8�}�ɨW��p='�Ђ�j>�%��%�[���$S�
&|�z�V ���>��"*lkvs���f�͘����1J2�3,/-��+,ZK��t�\ ",��q8��v4����B#Z�W=����lxNP�7�c�kA�/�V�҂8���)WM�	�0�l���ޮQ��PN����E�*U���Rx9����I
����$!iF2��y����z�-��qQo���c�
_)�7N��w/^�Xr�q�zp�<��S=�
\5��EK�Q���^�7����=P��h��*�@�� ��Ӱ��2�z��>O@����ڔ_�Y�xx6U�k}f6�cƱVyse�7�<sMfU�]U��rQ�QC�")7�V��R&�����PVVy�{{ݒ6���}5�f�(��V3I.1<YH^��oD��ŋ����{���~�O?uV�\�'���H2>뵰1��D{\��dH�E����H:E�1 t�6�g���~i��!N�uK1'��H�e�~����$&{~�xMlDӪ�p����J
*�x���.��3K�M���ø�{�`��Z6�d fHN��8�X��aH�(���;5��'N��H �ن\��/<��P_"�=�0���4[IA�4�W/릆0{��W1UϬx��F����5\Z�Z� 	�(�?��=��P�]��RM�?�� y�)�o�M7'�6��3�����K�X� E����>��瀤gx������S��U+7<z��/sw�=�ȱq�:(cZ�{i��D;/�M9�䄍�̙3 �0�����ş�&�a�fD`��4���N��z�w���A�UX�cڞ��s�>��D��\Q�6�0>pdm�Vwas��4/:�w�Y�������px����8���6�$�F��]�E�C�+@�hH�����h`�D����n����]C�܋(P7�e̘��Qšm�*N"�����3�"�b����ӵBV���A�t;�!mqin����k��H{67?9k�� �ܺƋm��yjX��e�
�W�.���no�y�,��ڹ����>�hU
��Z�,j��i	�xS����hcɳ	O3��V:A� �S��z�8�륅XU�M��G��X��V[�=�5M�2h4^�K�
�|H���~?�<R�0/����qQ�׌M{qe��r��Z�s�9�
x5��@T�'�'�K}�Oi U`�T6Q��@�ЄD}��1��Q8)$����+h��Ӫ�A�

J�p\���{vRr�(�CP�����\�v[��Ā��}K�G<|�m��u��e�(rB8�D �/�T��}"�1��+c�G(�������<��~��kA�/�zww��8 � ��c�vm�s�����m���R&�i�$4��5/�F _x�1O�|B�ի���D����]dp	�ױ��q�x�ɲ��5m ��$j8I��0����A��y��x���uդR�A,����zr�l�������3A]������b�&�ӧO��	����F��u@��U�ڒ�¼w_H?�5S�����M��,�_$����_��z��Z"�@���}!�\�N��{�����|�ڿ_�^���R�W��R6~yV����؀���*s��V���Κ�H���ws�w��ǡ�UN���-����Q�U��}�{�S��8{/M�������&�]��h@�a���Ewms�';����>��rg��A�n�:
�I�ץԞk��fڦ��|"��P]?4x��S�������	� ��׮��^�����L=������ţQvSa�L���(IeY���9������~M��A�D>7Q:b���O?����d:t�l3mj���O@�����yD�r2�C�UȢ�\g~ց���ȱQ�H�q�Z�v�[�+���,�'��m.0��A=�hL��Jf��A����U�1�����G�d�xʂl��#��� R
��C�� A7P�8��*g��݃@|Պ[b�*jx�)(>���Q�)�
�4/��$ԹTR���z&��(���q��^��3x�po����7���V2� �;xmk��Yl�x߃GN�pm��l����S�����m���C�&G�$&ڀ�I�{fwo���(�V��~w����`��-W�	-���RP���1�?�+�O��G%�E��mP�$?���:<G_i&\�+ҨB�״�����)�� 9\�ܫ�TC�Zښ�9�m�"��ɒ�۾�w~ 밖�N��R(��Q�'�\TP�k�6���q�kԾ�A�C1�v�Ǌxnc.*����JZ��Ӓd�R°�`�5��̫�.}��3�T(c��$�:I�D�5�V(㟍e�O#?�r�c|ćK��Y���b,
,5)K�4���F�^#�>��{���o�u�O�n�D׃��~����ί� �v�ZZk�z�>�$��q���c:�Я5`���=_*��ǣ5�A����[�O��T�|B�*������f����>V�B��]>�:�ޭ�k�)��? 0G�F#6����#�0��'Yr�ԉ����|������^ॉѦ��L�҃_���2P	mtA277k!����F�?����g>���CG�"@\KWo6B{���%�6m��U�*����������F�����C��C���- �hԊ��W��=��Z>7�$����Vo؟#�ݡ�F+�1��M�����*mlmZ�;^��Ԯ!0����?��Jy	$�j����ı�ʍ	�3u�����̳�`ۋʋ�&#��j�2� �>{\A''��r@�^��Yz!u/�B���׶Z��$Ud�����q��+��A���1�@Ze�'87x�
j"�9��X�,W:hv:�86~,�ic��Ƴx;E
��y "�AW�
�X".�$$���|��7��4
�@F�u�W.�A���M|�������^��d�W��5�L=˚��*�(��Ew"]0�*�&X���Ox�h��c���6M\Ԍ}���"'ꥮ��YEI��2�ArU�P��(�
^5ζ�%����a�!��Y|��5vz�lRJ��T���T������'���0D���;��@�4�T�t�hw��\�П�:�=���t|Gx��q�M�-d<f�8:>���^o���S�c,`���	E$�����z{{YɑքG Z}��)����no��9X>n��fN%A1�ʲ��7��zI��ƀ7���z��W�0Hh&26N�9�x���2�Z�t�*h����O�ד�ÇLg� ��,Giؘ"���7��8���駍BY`n<���+��V��͐��Jz����x~��/�$aR]Q��C������f'�-�޹�����/8��W�+�R/z�ɖu��%����M��c��x$C�s�a��������P��|c7NF�;9��G���#�?L��ܠ�� o�lE44�Ӟ��4�z��<���j$H>������?�y~�>�gX�-d� ��(`1���{�'�x|���g�ɂ�h`�O۴Mۗl�?l��v=_{ee%
77�B`{�ZE-M]���a�k�i��27C#C�h:�V�z|�6:T㙣E{�֐9�z���(���QgfF4]=���e�j�Є����K�߱���{RLtq]��|4�c勢i$.6����0t�g��$���^ˇK���PY�;３�� `u�G�z������W�{���G\+{��6��^$�b��r{O�r���hm5�7.��Ǐ�=����޴ܭ~7��ZXє~���E�i�ޛ"�n�i&|ܘ���E��M��5�T%��r��U{���%�Z)n���eR_G"����ꨣe�Fy.�R����'�D����d-|�:Ԟ��Rm���V�D�e߈W��/ޣ��%+����.��0��=*��8v�'����%Ƌ&l+e���&�<�LY���c_$+��|vf�-����}I`��d����Zjzݤ�__/'?i��Ѡ}ǥ֋��4=���c\�Ӧ2��$���]��&HE�Y���@=����k�C��1��)dp�_��G1���9���] 	*�-�Js���s�uVr�J�n�V<'K2�im�vH'+�:�T���~�+F�P�X	$ �q���@�̮�|~+Ip_���`{ߗ��
$�W5�	ߙ;n��<���lH�y�|����%���G�Diw岔��1�#ǎ�PZ�Wx?��G�?�Б<�F�}����RR�b�8A���h��v3�:�"��h{{�^�|�B�Q"�i�DI`�����Z�S��K�]��3��N۴}�/��F�aj"W �{�#������4��v;�ȣ�jQ��jP�D���4��f�x�4BW�¨�j�e���w�Ȯ�]�
�B[+M�f��y:�����8ɤ8N���f"�6JD��\���L�&R�̒:�E��R�(!�y:4I�	�0i����c�^q��bS� �?��<��D�#O	�d�J�aɳ�u�� �i�a�z�������Ϩd���{��r5T�K��a��߃r�a�)�W9�J����þ�ɹzg������&C��vv�����G��֝���p���k�����xDcӺb_�9�H�
�7c�"_]�DP{��T���o���(�o �N��">���e�� To\�`4������jVc������SC��B��;���l�#t4o(�3p\�C�'@wDt0��Ƽu�-�-ơ�|��ﯠW���oL�p�+�c�_ ҌK�3J�wv{{t,{�葬3Ӊ��q��NExƬF��=n�|�I���#<��#e%�mI�f�*ԫ�^��pv}��$�8����"g��<^-�˰fxO4',B]��`�8�>2!�B�Ъs��%FUA�z{5�
;*s
*K(���w�h <��n;c>��O0=f{k�����c�s\�7���=}��gb�hҮ_�}ŀc��&�p�E�1�������l7*��L$��\�����h�9L"��h����g�=�E��q���p�] kk
x�mڦ��l���%�n����)���s���kbǱc��mnn�,����l�vhi��qL�?�#?�����dY�L�L���<ws��Vi�] �8O�w@I�5{�'��'LYa��(zߊ���+��M;&���I�V�d��N���95N� ��z�y�mUjO5���t�Da �� ��=p.�vW ����*l8��MTu�o+F_��y��H?��F)�����.���@r2D,��d+�M��ـ�����������_�@X�/�j�T"�S_;�;\)K�i!_�/�<i?�,Ss� I%8ǔO�d5�$���p�cP����CN���@nk��*��Gu.��uy<$��R�$I�'�
sR,���,xԹO���'rĪ:�h:�g,U�f���T R�U9D4��10;$��x�Rڷ�-���B?�m���������due=�x�"VgΜ�P*�D��p/@��C��Jǁ���U)emY�4"����e�Ī�U@�$�~�M��RH\ ��}?)=�q�y��Z������ �˹T�u�]�����zn�F�4�ZÉ�7�W��fr���:d�~"���z��;;7��+A��o���RTL�Wx%��ׄH��x�@����y�,�ŅE^8�Ñ�ag���Y�ow�gqJ�O�T�q�^�l�v����{>iڦmڦ���%<�����'��� �?򑏄33O�<�t:��ʕ+���af��F@���Z9�n!IH{R�y�&���h����y���!Whk9B�u�1Hw�`Z���'8��h��K�}6_l��}[��dpH�0i���z2��s��q�{�/���忭��
}V��R�Jd�M
>c�������GQH�L����򯪅�U��M���{�Y	���+y�*� �E�G ���&���b
MH�e)3\g�<;��z��ӱp��Vm�jiaX�_^�D�ܹ�mH�E;�e-ẻ��+��:p��.�]2f*�pFCn x�b�G�\ˮm^��33�S�.]Ƶ����ozӷ�'�|J0��܌}�+��9�H����� �r�[�������fsk���x�����%#��^��_��m�C?�GQ)A��O��g^��������FB�<�|r!��]&���)T�_�M����*k�?��sЭ�-��:$`�9dp��`<���l��"BR����=�(
�f��ǎ���+�4i�4!���T~qE� u��Mv��ǂb������-����n�^/.1k�ӦY�6ɂKɚ�J�M۴M۴}�5�_2>��ݾ?�@P�����~��v~>
�4��ZŹ��ER� �I��(&�8SX��$�r��+Ж8���6%u���%iڦ�/v�����5�����*��, �V�%t�R��UU�jR8N���B}h4��}��ta�I��]��C���(9�LJ�Z/?��u�����r�	p5W��v���k4�����8 p�/$Y/	\ P�;��LiD�sYq᪳����B.�[y���,s`�2'W�D� �tc��ӄr��Ѭ��!۳�Ι��6����ٶ���� js�s��5�j�.���Y��Ck�'�4;r�HY��Lx���kR.�*ka	d��Ɋ����k�+��o�)O���{��� �K�4�'�uf�|֊,[�ȨL�/;l��E���4h�Z���t��,A=�E�g��;�Q�y��*`(���Xƞ���uC�HZ�V�-�	�dRW=��;�w�ANj'VI�����K3�>ml��nw��e���sڦmڦmھ6��U7�Q�G�]����{{+��x��B��a�!(:����0�� ���$�5�¬!�S�a�v�՛��~-I��h<��d�HҬA��V�5�]��:�Z�?' 
�IH�[G��p ��� �qq��#�:"aL�w�����zc���I�$K�9�m���:�"P5-���yJW1���q����}�v>�z�VcD�������C��ĕ+-�?�я2��e�v�������+)<d�o}�160����Rh�Ɇ�ï7=��Vp�Aj�)UP4
PJ�>��suE�,�0����0�zj�p���������O<�Ε�U~/��wp+Z �~�'��v��zю&��� hϟ?��4K �
�f�y��F��P0���Y�����6��`�=�������^�VnV�6� � �gZ,�9�g�2��ymɺ����|��������mڦmڦm�^�T8���1+ ��m��[���V�ٺvm������U����lnn�����q���Xcn�+�1���ϡ�ҵL3@8x��,�뙹��/��k}�aMe$��+�&,i���'(^^�_K}�y��Y_%��+@��p9v�^#�_F�W��ޛ��z4�wg��,����K�
	G��((+��8.�2���vv����@����%0-�b���/ԍ����ڤ�r�r��d�CyYS4+�9�^X�w��:�D�2�|�R�^[3�c�mڦmڦmڦm�^�V|���}�<����$g��V���G��%�c��I�a��*�@:� l(����Kc�&K!�`��{gsWېs��8�(�@` 1a�aa]�0)�	�@��U%�PD���TCp- pV�`LJ?��Ja��"E)��t�'O��'��R��oy����x�ݽ=���3'�L ΁�-��iѿ�k�Z�N<��[i�V��S��-.�(ٺ����Y?xZ�\ ��i ����I���S�H5ʮF�F��h4:�jՓ`ZNxڦmڦmڦm�n@;r�p������ՠ[���EA���!R/�'�T���W���k sx�9�V��-�0gF��X3)��vK:�j�2���ag�T�)�$5H�q�9k|��yի_m����C�7�3�`R�������۝�&�K v�S>q�����5��λ^��i�z������4WT,��y����FvPo�����z;�%��P�IM�P��l����^w_*���������:�5s��id�gΞ�gn�ńdU�;E��z��^3m�6m�6m�6m�vZ�ߍ�q�r��q���3����C��7QP����iϰ�W=�3 ��5I3
�/�+%�A%Ș��:ۢ1�A�_So)� F�U<03mT�t�V��6����a+�	�mY7;4�N�\�x�)�9=�W�q����DD��\���e�˄;��Ue�F�in��V~��q��A(�xt��"6d]d�c�:�0�뵬?e�vg4��Ur�F� Kf/�a���p�g�&x(�?g���ft�1�}k#��Ԓ��<�B ���c�w~�w2TT������(�C�gnx�޴M۴M۴M۴��l�F#��fan�m\�
��m��,vqa��wQU����"C���l.]��U�\c�E�<�a��`u:���/'jI$<1��B�!��VM��c]a_�"��1 $�U��:�&�8��zmlVʢ�w�e�3�A�l,�� j��
Y��V�̄��^:�p?�_Pp��´Z3�zb�����3�N�@!��^��4��KK1�d6��KQP�xx�a�)�������c���`GG�X��^��9��)��P<���滿�{���
�q�
?������o8⟶i��i��i���m8k����<��"�v	{[�^��VWW��_��+9����0/���20Mg��1Ph8��`6���J���[���'����\a�e�G `G���?c���Wo�W-�r�}��<��7W �*oq�YH��Z����2��f���d����E�y�9�~�����%p��'�z
E:p�ؼ�+������ݯoxB�c׺ɬ���8�qݍ�#������������g>��;��;���/�������of-����1}o�ߝ�i��i��i�����^j5[�oo�DR��~׭��;;�%�y�Qs��q����j��a�ᔪ���yU�(mE��V�o�E�,��T�ջ��2�CA*ə�M|�߭��5��P�Kx;.F"��	5EPD}��ad4+���*�*�N���\ ?x��/]6���O���~��x`�;���������=#��j����Z1?��?nG�8|)����V\��"T���A�!�q�hL}����q��� ]�x6<�2ommE���������r��?�Q�]����f#�zx�mڦmڦmڦ�4�a�ު]���%��{=�v� �6Sڭᗛ��������[o��<�ȣ��;�2��>dN����~��桇6�[�,www͡��r�|�<˼׵�$�PU|il�Ĭ/}]U_�&�F��L* ��m�\b����J�}��e�H�"|9�R8��L�%��@�:#z���w��W|�����{}�s!�,5�����h����Be8N�ݲ=���ަ~^YyI�/�FQ���$��A?�D�ԙ��"2�.]�dn>y�Y?�n���Xn��6xp����d�������W�q�=���ɡ�`�����}�#?�#�fڦmڦmڦmڦ�ElQN��������7~��̩ӷ�q����>ko��Ns��%s�=�`Ł׼�5�1�|yì>D�������ҧ�~ƈ�C�^՜=���d������h�=���M�r����(,�@T)FzN.˿��x��^���9_������	`A�P��J5��nW|:��h�^툽���]���~����e\�2ʋ��M޼z��@���6 kp�����8�z~~�����7&�����8�F�1�F������?f.L������Q�� T+�e �]q�������������.�?��ٯ���"zoynn�7{��������i��i��i��i{[�v�e�QT��3�щf&l��4s��?�v3�0o��n�B�C�~������l���w@@����0�6���{˙[,"yҬ\��0R8�sЦ 3g%�;���.{�����	J�E�7
"�B��,//���Cfkk�A���q��V���Ѣ�V�[�n乺�`�^k@ �Ԩf������������+��#�T^����"�H@�t���pr]-��t�.�ƣ]��ŋ���\��a7��d��w)=Y��Y� g�z�x�	���d,rgbp�,;��q�b_�������A�ַ�5��w�L�G�QLV���o��_���y��߾9�䝶i��i��i���e�4#���.�3���/��G���UfgQ4K��By
�՟�V�=�o|���É�'�'>�I��3g���>Ips��&K�ɃI���B��eު,��D��J|�a bz^e��V���HS�]��.���P<�"����D��{�C�>���R���;z�$�=�,V@ w0L�����.�Q����C��0��Ȥ�c3���l�%Yz�̙����ho{�ۀ�?�ۿ�o?5j���?����e�}Q�Ui�~�Ϯ�[N��j�I� 8����"H���o������T��w�ü���ݠ��g�~�Ի������uu
z�mڦmڦmڦ��hY�Y�'�h<�!�z��F������-��̃~��梦�7��>VC'c����?~����_ ������g��z�����g��0��X�m��ƃI�"��<}tO �<�ʫWg�Z��t��Xa�˅q�czXkskSj#�^�l�k�����4�{�ሿ/5 +@/J#2�������X"*��vw�\/.̳Q�vh������fL#��:���p�G�`g��6[u��//�d�+��ԙ[~������Ǘ۽ �[�9����`;M��v��t���3�td����x�	3ә1�k���ORG��pk�
�E�N~�{�c���������y��3k��^����O��/���;��$�K�K����hwvv Ob����΀������h\�/fg��a�o�����ϱy�n�������J��u��N��o�w
��������^������}�_P�vw7��d�u��Ís@�^�O>VL���h_��V�=�m��������t�	l��Y��~��S8�jfLo㪸t ^GYh:���z�U9w�>*���>O��E��{��0[��K��iѵ��z����њ�a�9�����hHj��ꅼ^/�z����r�2_���Ö�����2Q��y��KE�y��w��sh�;��bo��E'��܎�������U<���r��^Z���"��[�������yΙŭ�/noO�s��%��^��i��kw�w�q���/4�qo�<�y�7��͋����>�h��ާ6�����/h�E�]\=���Η;'�W����`�g!�����-o����w+�qڦmھLK�6�666�G>�s��haq���O?m����o�&� \xi���������k�N���g�⅋���#�i>���ʹ�s��Es��1�i�>/� ��@C�^ XN&&�t��{0�K����+ڰOnom�1�-u|� �k��s{}u4`5���gt�R}.g@�k�1�x�m:�U�7�Q��D@:�Cf������C���
>�ŋ���������zO�T���"��}��������F�c�kA�'�lX謧�z�+o��EI��������Ц�A�����$�x�+^�������W�^�i������������t��/��/�_IGľ�]���v�뗂��[���������ǵ0L�͠�|���׋t�i����<Ӯ�� m,̴¼��84����1d�Q�b�g�� �3�f��:2v�AZD�*���=��� z�~�zH����d4v���|a}�Y�n���M0��lgm1HF}�3��[[��"&qmi�QO�Im.k���PM�0��64��$M��Y/�"qE֠��k�G�h�X5�9$�FY��i-���!B:�a�h�l��(�p?���z����[2��۬����A��2�2d�f͠�����Z��}���m���`�G�fv;��㒃�m�5�$ٲ4��^o�7�)�-�&����'����3W���Dt���bqa!�wM��8L�4c#��(�<��	}�F�a������\�������KÂΗ��+���lw�b���Wy-�>,�tدS_���y\U��O�-ƃ�1Y"E�0Ɲgɂ�6W�Q�4�,��F����$��|�
I��.���$B��<�Ie(@��0}˟��x0�G�Vkv|����-�[��(g��|8���|6恭����`� CӞ:�������Ռ3��|��t?��1��i2�h85�[a��H��cu�l,�������|�
m�,��5����0]R���K�gR��V!-u[�[B@3yȖu.rA���l�(4p㽝K�G����R�4����3�]2�ji��(��]A�R����-�{���b3�$�t^��@7��F��:om�Cyuz��hp�,����c�^�qR��i��sp�`C���U�M�&޵��p?��S���O�?���`<l)蚨�AP���B�6nϴ�Ao��?�I^�~ż>f���i�]
��4�\�d�cW��9ͅ�����&��&��wRG/Ҙ
��"�\� ���h�c$�$G"���m;�R�2?��r�����:��r\��y�Pk�X������/sIÁ�@h�D�+�Zq��	�V�|J�����p�4��"*"����z����ѧ�s>�9ײpdsפ��
�F��>��A�_4�u�)?��f�h�w���v133��bic� ��yc�����"3m/I��6 ��7�԰��K���ѥ����ի�����x钹��/g��ɓ'���ڥ˗�˿��8Y�}�ɧ�ͧOq��׳�s��8�/#\}��ߥuE��)��M\SE`��+J�6�Af��^ڪ�n������V�_����S �I2.ύ�`�E!<�g�>���׾����r��ss�K��v���m�ms�lҿs�q��̧���y�����K�^����d�4{6%.M"�HK ������{�=�gΜaj���a���o6k��L��v�xx�� w:x�<�N�!�뮻:��w_�~����g���^�|��-�?���F�b�V�!�`�Ή͙:����BN��I���w��Gx���)���Υ��=������3��:�F�6�$�6dK�Iy�i�KA��O�1�@n(^k����6>C��8��[I�� ��cIdU�{���l���k��$����^pv�a�:	 26 )e�~-��I4�9�n��I�-����_��A�pyD:ρo�����W�`�ࡢEa�&��������������v��V��,~b��:�/�N+`с�4�3�����軝]!��wlv{�{7-B����� �D�?����D�A����KKK������8���EP*�$����s繿ѧ��K�'�=6]<[�M�h�~�|n;X�gX�9����С���@��
�^J�!!*p�,^�E�������p}�v�?�Cc���z��
��A]�����y�=S0$�ȩظ.� ��;��˚��紌!ԝO1������u�Ι�./?���s��S>�XQ 3
EK2�}D����,�E�R�ف����#��z�c\3�(�ņQH6	�t����v!C�!VW XR��*�^���H�	�UƮU�o%!��w"�Kx����M�;��>�V���q����=��{��Z����0�����>^��P�%�@=nX}���� O���N&�X�0n$4�ҧ9z'�ЗQE:�E6b���v||�k?��%�^�cر�h!���qGh*G.���2n�Xs��A�K�z��f�̍���,a�a[l�X{�����H���"�_��L��I�R�8?�!���.L)ػY��;�Lc�*�<Ip�YlȺ����lX$6��p�$�l��c���8��5���`��]�A<�o�F�x��yt0ۉF��}*�Ρs�#:�����A�5%�!�Q��g4TpIl0�������"��MC&�U�y�`Ȱm��K�l���4y�mlt
Z{Du��JCX?���;��$��E<'�kfgyo:{����?Kkl�5g��C��z�!�O���������sV1���rv}�{<}��we��jf�}����H��M���礼F^��*p��ʹ&^��oz ������+#<e�a~����e�?��.���u�����7 iMxь{,>{����#��-��{�W�~����o>��Su�#�/�]Y9�I �>���ُ�<m64c $�ر!��k��O��y�7��^?��8`I�Q�a��e����.�!4�|���c�XDǏh�^\YY�{aq�n��|� -��nw��A�-�'jHN�y@���M:�k�jt�N�1O<:��Š�7���s�a��������F��; P�z�I
@Ӱ�� � �0�p�Cyk�3	��?�+&,��L�΅�gee��'�X�>��>y�$@�
���@�gP�@ ���W|����Bf$���2�Zw4!-��y 7	$�t"4&��è�,R�w��'C�~��b�v}�0WUYX�S�N������<ȶ�2s�,a�
x*a�Є1M�l���NCGZ�@ߣ~fapȝ`cv�'��~��C����q%D#��
��� �j�s�^<��~�s��ˆ
�o3�����<O9��
��
``(d�;��k��܏�V�y諘� :�I� !��@����HYF G�%B�5q��G������xt��y�-Ƌd�f_k��X���ɞ���Ɵ��s�8kXN^�}��Zr_U�QMn��13-IƮx�C������M(��F �Ȁ����.5�5A���!B���윜�Z��\�!�I��}��?@�|m#VP���c�6+e@�Z�� ˎw��<Ɇ.�x}9�ת��2S��n�28B�1����u��0�� 0TbN
a(����uG ����^���/F_b.��B�T�r�x�����I��(��U@3r�)V��D�C���H-{�`
��"5f�$c[�n�����@�0?�G��r�$�8����7��| ���c#O >ݧe�Y�2�)�TΊbS��?K#}$s�ף<�S�z�^��z͑����5���;x�# YA���a"ศ�E+%=
2��B2v��h@ڤa��qV�XV�l7�g;�GA/�h�؏~Ϧ&����7�����EA����ԏ[u2�>k��x�[��Gt1Yܳ�6�t4/�o����<�;�w������]���n�^K�`77�9P�ɘ��{���ٳ�>]�z�����H@;rD���?�c�c|ƍ�@�s��ڤ,���}(�T;SO-�:�/7&��M�qTUR���6�և\���j&���<�+�ت�X)r,N�G�-ɯ�<�!�׉�4�Z�] ZM��sϞ�O<���]Z� vaXb�.��
J�����8f�o=~�Xc}}��Mi,ߘ���7��0.������i&�%�qZ�"�Q�i� (Y��_��כ7��������'>i^����[&�`�7lԨ~��'�@K�@�ho�q�wZ�JZ���<����(j�4�����Z�bW����x8�mr4 ٓ�Ѐ���bp�+��4�
b��O?�#��l52�I�/�\U�@�%H^�vw�|�x�����.o\f�,D�l˱2��!  ,�R��ǃ�6X�^[��f��|_�`{05�w:l^ j��ƕ���x�с��x�f�yx�|���7�Z,U[�r�p��=*�y��Zl� ���޴��ҭ���4��5`BC��@߁7
�Bǰ��3��Zx�A�{�H���4aPXCA� q� �N�� B=Z
0�k��W�Qo7�	_MP2���ߘ�z��ClL�s�8�x&X��'aM��Z�Fϋ���,��zb��W3�pX�^w���M��H�x�방J��ȏ�L��% ���G#X�7�	�ɆC��F��k=}A��ê�彼�P��_k�Ðs�ʐ�)������B
Ð_�5W�1�3A����s���/#>Y���To�c�)�E�az�(�<oU\��R�G�aFɲ.�3KZ�q�uB��-���p���ƞ����� �:k\*�q���|������@]������E�Șlh�!�?B�Ք�J����1ck����иM`��Ӌ������g}R�<�&8�r{��a�����Y?��5i.hߋ�RCFrؓ�O:�=�5`	�{ų��Ղ#PG2�\�7����C_k�8퇎D�I�9j� p�g�s�&q��EF�D7�)�v��X'5Z��Ԏ��1����� �����F�����(�8�zX���#��Gq0�PuT��x��1��*f�D@������_�)JV�%���8d�kd�ө ֋� ��̎�#^oi�,.-Z�*���egI�ތx����>�{t����6�9��w��|��YJ�)D�`t�!�L[G
�޸Qo��ɸ�b0��q�>�j1��=8.M��w�٘V��mJ�	9���VhTErUb�Z::=MZ[$�-�4	 ����w� y�3m�^m�u�mxi	��(��}��q�'�In^�d�~7m~߸��K��u �5޿���$��!��U�<���� �mgn3W6�r���ŋ2�i<#B�v�PyO�w`P�92?6y��+Q4o0J_`U��5��>``�j�#���g�t�~까cꭅ�������LQ�<l����}z��	c��GX�(��HU]ȗẰ�<K�����#�nnn43�i\�|�s��̍n/���Yh�{�����4�gi�@�9rđ�d|�A^�������
���ln��6vnx��3������B�xq�!6�~��^?b�# ̅F �(a�#c��ᖧ�J�V�>����Kvd�a@�99وxP���,Z\\b�&!c�lA��޽q�m���k��l,p��{{2��m: ���z� B��]�x�ݼ������� �9"�@��_zW�yx�`�U/��~`�!�f�n�l�t
�	�QO&�N�Ä	�ǧ\<�ܕ���a1PBHQ��B¿	_�xO��>mBBQ�˔���{��K�6�{{6)|G3Y� �ց�x_(9G-K� ���Y.i����7��A2���1�7���+�?�G`��0���X� &A�~�sQ0
@�F��͚=@�!�y�o\k�h�{��!r>�W6�r.��פm8�/�p���GáU{�&�,�F1Z�#���+Eס�RZ��?� �zo�W�&���=K�����t�\��	�W��x��d��9�)��?3��p=�dM��ܩw�@�>���>Y[�9�E	>s��n��AC�'8���E
d�Z���:'����C�xpX�=x�x�1j��'p���@|�1kdf��gãBk��]��~�0�}+�^(J ����2�z�qǳ<���"��r�aʚ7p�� �X�}�=���v�: U5݄�[��O�+U�5ӑ����y0�	8Z	������5?�4,\3��ǥU1��<�l�����U��k}> ������_^�+^�!���꽩��k�衆��8��gI��Ep˱��蜥~���1� ]"vBݡ�v�9��H*Ŧ��Q�D�z_M��q�s����BV�5�#f��}���|�DP��j+�Vi�������P�8r#³~�I4C�����؇��]�s�2ٺ}I ce�^9Fd�Q�N�eH�h�E`�u6Lx����.�"�X�9l�y�is�@��#G���,��+tz�J��"oQ�A�}��L��b��Q��t���me-�2�4��P�Pl����[[Li �	�*�ߣ����xʹ��r�z~�ە��hT��!`�3��}>u�����c��s�Xlx8�1�}ǜ�_���Ml�--.�940�~��U�����������'wx���p�܇i�|�����ٞ>}�}�s����Ϙ��1?񶷙������ʯ����|��쮗�c7�P,�P;rԬ,����M�l{g'"K:�B�A�٤ͮ���g, ,��st���e���C�[Q��������:���V�わf�)��R�J�8��&�� Ā�Z��n*�N������)_�D��M�=R}8��^�!{�ěpd�p	�T ��'T�}�C�9���u�U��N�8��U�=�0@�Z|���CP���N��
�AA�C��Ӽ�c1@bX<x>mx�=o	��>�G@��i�\q��
0����<�lL�YP�+6"zQ�e����1'�~��/���+��fv~�&�"�% S��5�]#�S��s6X�K��x�I6V˝��xh?ʑ���=� T�YZr�b�x��\-��C�ǧ�TDe�5�[� 5�DF�|��T-=�������)�}M�!����k���2J}X��y�EZ<���RYH�A�Cך=�`ת����yO�P%*\N~�;jlc���-R# ��f�N0���Q��r������1`� ��t��}���Q�W>������O��}(�B��N�Ay�j�gؠ#����Q>���3q�QH@&Vk_�;|F �$t�8D2�`Pσ���X��6rm{zf0�aXc���K�~�^/���ue�5R�)I�x~�~]ӱ�g�(��3�^0"u�$j��x��Oq�1��%���3�R�F�g�x~�D���7��� '��B�
=/���4�&�r]�����k��+��S�Z���1��` �b�3�C����W��=��7D�E {�#Xs�{c�-�(�xZ�^1�ZFف���X��l�C��QF�Ұ�x����n�Aǘ/��"#�Gu����Tg��k��<�k7��α�s)��}����0Y���JTC�kV��!���vK��З�%�9?F|B/�K=��2(G�3�\��NO`�>�è�v�v$^��5/^Hh>А�h�y��yL>�䓼?��n?��Cf<�X�;z���'>��-H|%Ɍ�����u,-��s�8��(�	�xM����7���0���.�	0�����x���uLuΔ%�%�!k�_�5AN4���Kd8It{
8B�����w�����55Z��1���M?��^��E��l��ߋN�rj���3<������S�z�/��i��uҿ����4_g�Po��wޚ\��?�أ�����Dw��e�m��'N0�����s����`���Ǐ=�E8:q�x���\c�@-�À�{.'l������̌�8D��3i:���@�
k>6�Q�U#�r��<b�-����}]A_X]o �����]A�Q��L����3JdC���%`�Ԍȇ�q|,���<���p�jL��z:*��S�	�����҆0��a�e��z�>{�Փ���+x\}2Ρ?u�d�k���IڃWB7,L�[[	<���/' ׬�E�sQ��*/��Uk��3Α eY����?ހ�My�F?a���3�{�~��Q�[�L�%VpB�I����C8Tiy��A�y�Q:���r֠���ە���q�{�MC�U�n@,ZJ�*�Aiz# �H~Sn`y|6i1�Ǎ�c5��`I�k�O!Fx���X<��x��%�����&���_/2��)H#4��Ŵ�o�7[oXӚ��%W�t�x壟|l�:�7�}��h��f��Q��_���3l�G�N�Z�|�fʹ/�&�h2SDt��$I�C�m�!�=X�VW+��C�����B�� �
��1��o<Vh��b�]^�z?��s^����C����{�����Hx�<Z3-�v4�������Y�}>��Ng��[�D;�D!3�0Wz���*��x�E�En����p�
��1���Ft�(�K�z��y�k4�����՜	MRE�9�jV�4�9jk��.�D\Y�؋�Q�����ku���dQ���/�*	˨C�F�Q���eJ.�+je�dh�1����(%Ʊ(WtJ����j���N��砋�{O(-��b����5Y���f��G�L�Oi��lfy.��zG�א�Z�U;b�W_� <!r~�⳸V|7�E�@��Z��R#�hA��$�ܿRh}���F�R� .��!u� �9];�?{�9�#ĝΌ�P�Y���@a%uc���,����>�����A��p)��d����j$��K<p܃$��xԗO���E��(%�d�1m&ί�T6�[B���ɹO��}J��x�D�c�̻�}�<D�80���i�w��R�����}��5�T*�;���>t�Y^Ye��N�ZpXw��ř�_~�ˍ�v~m^�y�f��������&�yZ~���f��f7�n�����1���� ���^�:������sL���p�<�i1�v��1CG�)'����Mu3d/2�"�V�n|m��c�k�
 h����:4,�h��W7/����?��c㳊��4a�ƛ�,�)���)���ɒ��\����1Ǘ���7*H�����@M<)��K��� ��}���I�+�EiJ�П�L>������.�[*�L2���J�j��� ����'�N��s(h�ϋ��RfjF�^��5��ϊ���U��hD��R>,�UA�$�L6'L\�D���$�XǇ&n)�C��Ӿ�kF���@��#G��������c�?��$�u�|�O��=�z�)&��¸pc��/j��L����:�X�9����[q�V�A5�X��(��+������c^��p�Gd��g��|���l򘇡H�
�\���e>�`��~U�㓓g�<�}��ϱQ�X�s���B�����D�C���?U��q�י
Aߟ������g�G`�ycO����^��>,��<�ћ���+��B��y�LE�[][+6�I?Z>�F;rO�H�V�Xc��U%�V�(�R~V�������L���]3�؀R�q��,�7 tS^~�Z�B����T�u�u|��\S
S�^x���f�{�J��1��G^��.9	?���:��֘G�+��tL�8f�	���~�<k<���%�����\�� ��Ɛ�[���N����t�@_I?����O$�!�T��>7��9��N�0qXS�����5�?�cpm	Q�5 1���?/U�i��$WxjH%��ΧhB1�O�e�_gf��*L�����h���N|�-��i���n��SH"�dnѳ���Xx���G�!@˞[�̧�/H}�-G-DՄQa��uV���'ޓp,�ه��D:�G�r]+�a�%���Ս`�)`x�só���%?�=�D������B84%���&�����#!n�؆sB I�5�)EM�J �ɧ�6ozӷ�X�؂:����������j���S7���:�g��C��xѨ��o�/����������������Nh�,�DQ� �C�ڼ��bc�����m�ݦ`2Z�����o>��d��9!Yլ�Z�^	�ҁ���x�W��j*�P���E���ˇ˞�
 �b��h�X6Sސ� -����w �� b�a��|�[��*i���h�A�y˽/.�����bZZ�h�縩gS75I\�L6�yo{�ht]^.(�_�ԛ��`�Ӊ�g�D���
{�G�r��f��M�?��[|\��h�ե���5�\�g�,����V7�j�_(i	J�����`<�*��SS���]d�P�00"�]�*�k	u�O�k��E%��E��@�s0�0�k>k}��	7h;;ԫ6���{:q�w��5��\��A?a�`!.AwMh]r�m60����f�Ú���iҕ���X�[�/	oT�虋�g1	�M�!D�̈U'Z���8d��D�]�i�&�2ܻR=0�E�r���d�~P��c���������14J�$,7ә+���1L�3<�S�l�}�P����:?G���\k�w˝�HOǉ���x�l�<�crf���!���S�kb$���ض}x�(ý��f�����))ʓ��f��Z5d��H>c<���������U��YC�r�	�-Y۴�uz��'B��iUri�s��K2�����ӥ&;�^u��á�|1�R��8C�u	kV�g^�N(�`�kQ/���ѵ��^�+��p�tY��d��m�$S�+��j�hc���ń�5'amo��8˫+޸_+4�ǥqt��i��j�,GI����*�P�-}�<�d�>����^K��e?�g�QE���Â0(��wN 2��P���?�Ix�e�ܧ��z�=�Ja���P��S��Z��^���>�{�4�����dRjX<��tF�sS�0�,󟛌cyv�S������92 z��]�rT���:I�V(Fܐ��fJg��t,���G�N9K�n��%�B�9�P�=Ĩ���c/��;�=����{^A{�.+2��;;7�����5�NϮ��O14ni՛7T���^�@�B<���l-����~��+� ��>/%w�ڕ�:���׮]�P3P�mR��B�N�&����3�������ҍ#N��.9��L=092�
�e){#6���۶����>\��5QB�a8��������ذs��%`��\V����E7dp�^$� h*�~}�����$�P�fݣ�1��a"ϫ�P����#�aJ�P"�����.XlPJ�蠖�(�E��e�3I �>dY�$����W��zPԋ��|i(�������6r<�8�"V��	��'�{�Ƀ�r,��OgE����5�ᩱ7�
����.�5�+�Ǉ��-��8 ��4��sĸ�|yC�l�!����:�=�<~��9w�\Y��p�"��{�5����x�D��-B%�K$�ʍ�z���`C=�:��ӈ��1\Y�
�]7_�!��瓟מ;Ϟk=�
����������צ>Ήs��Qy:�5���9�1cR�'�\�R~O�O�����B�Rt���7\q��.���<�xi��+ր7�1����))�O�i���av��5G.W�7�0�����oJɸ_�/+:x�~��$)P7Q��0�)��1����t��f����s��.4}��*�iJ���dMd��dK�>���R�jH�r]�� Y5|�Z����s�9j��a��E~=P��2}:�4�M@��$HM��1�&,U�ᵮ�-W:�C<n5Z�k��T���gS�o���k>��J�$���Gc�V�ʋ|��I��a��s,�h�Q�z)15��Z���1X1��4J���G�2���
O�icO�K� B�8����9
�u}WN���(�DS��Tv�:@upy�4��J�W/v�@R���/�A�i�N<��_w�d"j���l�v��DI�݀�_ĪB����9��*7V%>�nE�xK�40���f2��B��D��Ct��S�?v�8�s��^�� ��D�^���-�� �~>�خ _�6�7������a�� ���G>⣉M^�M ��=�_�`9$���I���k���.ƧN�4���KV�|1�������n���{�{ݸ���t��M7�Po�gghb��Ď��2O����X���$3�\��Δ�#���ox�Y���;l`���|��&u���,<*:���3b�0�ϳ~��\�!��'|����6Nd|���u��o�t�K �7���A�~����'b������*�׷j���\,��� �I�@��b"���<�Ǽ����-@	7�u�^�t�����k�b��Ϟ=Ǜ�t[�,,,��e'PjX�3& 
��>sXݘLh�pے'ڨM��h���`���ƘH �d< +���>��~�S�2�~��͓O>���M����`b��c�F���~��864��) �b� _��� T�}���7g%�q{���뮻�k���.�5�q��O0�����X$J������@�Te��TYU�� 偉'�i�D�*?R7=���������_zȱ0"ԅ^����fD��c��c�Y+H�5+��gq���g��W��|�3�0�FF���E�y��]f�O��>���rB胛����R���z�M� ׀cb\����csC�I�x�T�t��I����xV�*�}5ք'�������/��"��I4��Q
U�P�����@�ȅ�����N��Q��Z�
&{�=�I��jx*�Q���J��MT���R�f�D2�W��0>�9U���AW�7H��h�?/��pDΕQ0�G�S^UH)�:X��,�j��I���j s�>ӨIDA�gB�R�ҫ���k��Aׁ*����^uQ�)�3��y�_�}��P�I8 Y9`q�4��?q2�kyY4G�����&�Z��~��&�iu�PiTT0K��ͽ���س
-J3�=D�ulk���&��L�Y"QՄT��1	�S+�Q��Ј�zu��[�~B5 �j51`����o����W�L������NB3j �'ޟa����զ���"M�D0P���;����8��.�%1D�2��=#
����sV^��g<������/�Y��a��C@�셽'�(ϩ9?L� p����QN���?���E�O������߿�?��7���Kx�p�����@��_P'�H��o�W_���Z�z�
���Y�/\�����9G$?ilL�O�&����^���������u�0�{��8L�_�1��p8Tﳀ��6EGT+$t�Kle�p#��x�`� ě�J���������ڻ�`K����}۽/�6sf�H3#����1`;T*��+q9e��xpbʮJ�R~�S�J"�S�cRv9T��<$�)I�Jv\+8�.$@�F3Bs=��w���Y��Z�ϞAرAF^�~TS3:�}�������_6I���{��F�(s&���a��8���0���a+l���۱ٞ��> 6��{b��n�歛Y&Yi��QV�s+J�������]�^���V|o��n���T(�HY����w18�f5�����H���B�M	u���B��+.:w�j�a�&qYE��vP	��=��(,��7L�񫻩W�.Ӎ��@��O��O�'q�z�u|�FO�es	�X7�9i0����A%\ڌ�����P��o�-H�X�]�+	�NQ����׾��/�(qQ|��P�CRzO=��=�X����Q�c���ey�m��}�x�Q��H�h�A�[��q���N��ޕ�¥:=.��l���}*|j��I��������r�d�4���b5��kW�^��y��V�U�ǟ��!D�6�szm㈼ʫ���D�Wx��%n��8��mc:�(d���_���q�msz}b]r�/�#��������o�@��P����'��N¤P��D���Q�8���_ۚ���Jʰ8��Q�`�?;Au�q����a�/D�>��(k|�zo�������^�j�����9�5R��5Ρ�"|f<cȉ=l���mD?�Bw��".��18��:�~w��W��ܨ�����'.����Ha�k��	��A^Y��Ik,�ҮD#s�b1t'�)��� ��0���y��hn���u|�lp��Շ	ҧW���Y����~�ɔ�՘�m��>�醚v?a�&aZ���~̶�1HǳQ8a�.=����.�ק�d���=�'�q��:����8��w|��iK�xf�7,(3	5��o�b���+<Q׵v�S��,L��,�!��X�fl7hϡ��B�M����~X�ھo��|��]A	Wa�N,g�0�����﫧�B�,~u��
��ڏ�*@�}�>U?'�Nm4uj������7�_�,��,�������C��i��/���KBs{��YX�9e1�����+��>����h��6��>��o]���	y���[������W�_X���8�U�B��o��o������E;�������v;��#o|xr||R]}�Z�w��=��#v&G7�b_�v-,p3{�ʷ��%b;o�!T0�x�'�&?ѭ����M��ߋg���$��V�M$N4�a��͉by���#:���pIW;��$�+��w]V���έ۾,!�f�w��f�k~�i4�U�6R>����?S�#E~2@�[���8
����&�u�|�c�'
q������ڵ�����O���Ʊ^2^Ҋ��C��?�}��&�(pi$*��h���0��u�.����t�)N��t[z�*S�k��/�W���v	ͷZ��م�f���;����U�����kqYbݯՈ�ѹX��Y�`#�a������̿��/���)����$�K�V��m�a�G��Jxz�1��ѳ8j����s'�m���;��f�F����\u�1��筧t�K6�c���I}�׊�NP��jT&~_�P{z��x������QJ}_'
���Y�'�'^j$^:�����#n��)GC�X��B���z������kmW�J?�~�V!j�l�ĭ�Iۗ­�����uЕ	_�1^s��rt��~L�5� �I|�[��QX^;�6��a��Q�8���*�T���g��/��q�7��h���w|�t�_��Wm��VWr����~\����
U�K�ǺY=��J�\���|A�m+�YP�?^jå߻�Ą�C,X�ϧ���KM\�;n�qR��3�S��׿���	�^�0�2^�������,��k��ɨ���6'��	A[�$E+�Q(����]�D�ޚ��:SmwC����N�Õ_?� �K�
&:A����:)��{�	����}����NmUѹ����k��ܷ�������&��F8I��궟�����g�e�����o���Va4�*|m�V���߾���K�H��⹍�V6jj�5;GvuQ?��e5��ˍ��Q��+���_�v9~>Զ[��>��_>{��đa����o#���J�J??gik	�٧?�i�9�֚s�z�q4^����H���Di)M�k/~{舢��W5�����?I���p�|��qYg?���J�]��?��٧��Ӷ/}�+_����C V)���}�{~[�Iq��}�o|���c�=Z��G������k������(<����}�Cϲ�M�|�۸��ov;��x��Kn��v.5�.nܼ٩�W�0��g��;l�èH�T�pcQ{�:��㊣(~���/����T�ee�8���K���j� ���Ku:��;���D��h����m�`�	_����F؁i'/čtZ���:��%B�lv�uџ̓@�W�]l5S����~��jQ9\>�߷��!�fd����HΨ�AO�.�Q:�OU8��L��񠬃�nK�~��^7L����G>��=���
q�u��ӈk���;aM�����G?��ȪɊ#)�Y��`CMX���C<p�v��%�z�N$�c�Y��б"�-���]uP?�p���&�EK�Xbhю-�%���A9v���+����򸽈B`�ֿ�����˄�g%��������Q?�+^���}�k�����'�~U<t�n��)������so'�s�:k����/�(�������]W(�}��k��H�^/���>�w<Q�s����r�F�%v�3��t���~7Lڌۛu/	�~/�hœX=7�S�{���[Q���_�x�������p�>>�8�_�xrq��G����:��Y�"g��1�m-�7�vs��i�镝X��T������5��2���.�dJ�� �ݷ�J�0u�N"l�B�Ȫj^��V�~����X��pU.�N��+�8���u���f���8��&��_lۧ}�_gmW���ye>���C�z,�?�~͎e(��K�k�FI5w����G�?��e�N���z���s��z�|G�����.��D,m�}��_J2��-\ݸq�����:k���[��	F7�~��/?�;�}��7����|O�n[�����0�\�K�}/~M�C�O����ZP�銭x�3�;�3b��xB`'����u�d�	�~���tl�����#����o�ۇϮ���Z���m���-���(\a��sm��F?������>c}v�Ä��H'V�Gw�u���J���Ս����apeN�t;�o�d�����^�GO��a��N��_��N���|W��� �9�>|?�K"��ŉ�z��O{����{��瞳<��.�T
��zx�K��l7��W���X��O�a��7<���#�l����R�4|7�����=ӳ�	~����GݎlV懻�z��u��{g�κ���_pgT=��oy��߾�Π�n��v;��ѱɰ~��`��A�ѥ�tR���Ck�X��3����3���+���bH�*���āp	�VG5bV���Iq�-J| �NM�a�/�]8�*����~)?��
���(�}=��=j���X����tg�����C�o��\<��ã�"�ek#�Z
�7��y��%�FY�vq<sWA�0��wa�ð���~k�
5���QH� �}tae�*�[�!.˻�ڹ@T�	|��G*�}MJ��f�5~�KV�?f7���g����X��YvZ�z��O?CK��;:��>d'���<(b��٪U���W��ͅp��mS�������ݦ�k'��o;-����2�-����t���3���tYX�l�^���u@�I�'��뱆 ��|Zo@��e8?0a;�_�m��9�Fu������?s��q=�6�#�q$9�X���_�X�<փ;c��ڡ���=j��Ȩ.���&��x����c���'�|I����5�Ш66^Yp��mxX��/ �;��+Q:Pk�����o{nqd1Qm�z���"����x99��oN����҆Ǥ�s�7n�qW�M[�N�89H��ަx_��V΋0ڼb�S�~���B�����9���W^�e�E��.�s�+8ƓG-媰鶞�?�='���kX���JWشA�^��*�JR�y�C	�ܼ}[�MO�$t		ǉ.|N��3߯=��awY\)��xa�+w��k�����,�j������-d侖U���������9ƓC?9��P£���s��Bk�5`'���_���'���"�����l�����>��1ǽ�O=���o~�y{\���d(�&i��,,�_�eN/�t#�r���1t�p��3g���g�f�:�\�j<�3��XC�f�_�|<�5��~���x���u����l��n��N*�1B-$�ՀuׅQ��N�����awhWW$O���ҥ���8�� �/��
��~~O�Gc5�&��	��Є�xU)t\^e�{�h���b46!�z���%���v�q�6sk ��"�^�ڦCP��������89�������=���g_N���Ν?�}򓟴En�\y���ߺb�ݸm��u�z�۱_a^�F]��{��x����|~�Z���5;Ij���'�=��������?��r�t�ҽp�����rY6��h�h�|UN����b9������[��Mpr|\�xPk�5�������؊�]��S&Tq=��J�.���<�a���$��Ƨbw�f�ee�W}�{�C����ۻ�~^��X�=2����ޯ�v1CK���V��[��_���Sj�ո�i�d�2@�vҭ��K\^���d:�6G�g��j9o���6�����j�엫Q?ZU���{������=0w<��g��s}8g�V�P�»m���]��]������G������g6٥۫�^��#��)��Y���Ёw���u��ns��r�}s�Qȴأ]ޛgC�t����\t�tv��[M��P�z��/�`�ˢ(��:/��֤�Z�ݸ/W���.���fv��
����n��Z��s���sl�~�/:_=�Ka����&{�2�a:�A8���+w7��ڮz�1�ܗ��������{�
�m��e^��^ݷ�Qv�XW�Ct��{�{���O��4u�����d�w�y3r�o�Q˺n_���7���˄
�]_�l1���myy��.�iF�۶��Z�-��c�%i�M�s[�)��ځ�����)�8~�p���\�B]�t���k�{
ݩm�.���ʦ��6��f�U���sҷ�~z��}u[�|e�I�r�6�Rn����D�4�֭���U��8���V�
�%ZN�\��ں�lӑ���2!�z�N؊�PF�󋹖���2L6�|۳"��"N6s�"�Մi�2T�:!����:��J��þ�SA�t�Hc<8꽉�G�P�џdn+��&;'Y�iX.9�WOV2�\C�+b��w߷�XcYJ<AQPW@��k'���khue�ãN��Xb;�n�����N�4qٿ��R�_~��otZ.z�GӴ�)�E&Vǫ.N�����9�6�P��x�g��#�;��m[�+�,�k�E����Ix��]t�`�p�/��WQ�N����&G٢z��u(�1,
�A��F��<�Y����h����5����2�Ez��߼��m����zrզ��)&��Pc��������v.��cc�>}�ʕ�CYAZp�5��|���mW��1hB����j� ���
��o��久\D�fX��������bw�x�J��uk�廑�uS�S<y8�p��H^|��v5S��:�~��k�yVΕ�?��/�Q�mԵ�Օ�7om�ǉ�9��A�=kߠA+���wV��P��N��>���bv݆]�s��bH}v�J��mđ�XZ{����޻Tq?����~�-}�����N�on\�Q�Y��u�{�*-��>
]]|y�*����3��^Љ�v���t�^���h�X5��W�ޯ�������p��i���}�z|W���~������A#�ָc�O>�����>��ޜ/�W�݃���+��F��.ٿ��_��o�;���b�L�ut�oo����v�۹*�O�2��ڭb����,'Kk�1����n�Xխʹi�0T�O�m��Ա�I��k���}�_w-]�^��o�ѹ�k�7}�[����I����̒;{s7���;8T�Dd�������h|���R�������G��������]�����"�W*��65��K���������;(�y�.��a/i��L�[t�c�Ř����g��#��t_��v�.��q����NW�|T���lk�P�/lDi\�ŉI.�P��'�z����	^�Nd�.����_t���G�ښڨ]>��4���b(}�U�ʝĭW�n�pa����:.��k�~9r[VZ�>�M˾Q���'j��.]QY̗E,;p��N��	�;ؓX����aU�ǵ��YQ����n��c�bY�j�O�����Z�O�����k6�{����ޫ]l�'��R"-u�ޜ���wM
s���׸ڣ� ��wvv�PW�祫C��s!��'���_z.��~2�p���=��ea(��$D�,O�����O�w�"��զ��uA���ɷn��B@/6��ʙ��:�������η��}p�ݢs�>�o-K�M5����RW<�Η�0m��F�����u{�x2�δC)�MDW����=�7�����t�UG��h|zX�dT���bH��]��?������tuz���8<����h�]�!;��,C��pE�}>����@,w��g�TB��c�4_�s|1�Rl�ڇR����U�£�s�����O�։�檌tR�=r}K�q=
W�2�\���N��6��*��	���n%���S'$��7����+a�ɲ��m�K(i���aۉ��"LH/6>���#�����EE�G��<��<X?��ڹYy����v�����Z�?����5	���wf��_Ȟ��3ٿ���NN����ٽ�'��O4��;ww���٫>�~?��ת{��~�z�3 x7~�#����s����t�����.���=�^x���~�7�}�����������Q�r�~����0���==���������r���Q:wy���{�
z��F�:_��!����5��纄��3�&�۲ZW�;$�j�e�rUI��=Q�;�c�]���ծ,4L��
{>.+��]2T�'��k��a���i�B��Jwpw�л�cK�V.���$W�X�}��z�[]����d�k[Ml��\���
�{�;�B��+��t�����$/J��h ZA�DJw@q�w\��P��]�-���Vwi_OQ3`�:ުdF��F�ҥB��:���w�Jg����ۧ�L��#�K�\���� ��
������+�J�'��w����ʍ{�j��G��V��B��=����ۋK��m�y�1b���ྈ��6l=x�E�鎳�7j{;�]�*B��fY��������vqt�ӥ^]
W�רj�y�H�ڧ��x�x_�碑$M��"6�_jԺ���G���iif�V�f����l�����E�ԥR{*�Pē_.��H�a��OG�����+���<􁮺�ٷ��*l��z�G嬃�m㪈sA6�6�m����|~lK��whX$f��b��%o?ү�6?��U�K�|���(p\�&���q��>�k�N�ز�_����݆l��b}��&!�ْՍ_�T��q�3V��(�J�b�����$��ĞĪu�I�-�au��P��+u�%���*�IY��^��
ܾ�&p�a�K�Ha�
ue#������t���m�UO�'n�EuTR3�9��f���m�.�]����¯��j�0��t�pdeV�WX�m�k�s�X�������O��F>,��rN���dT��tqq�̓�w/m#˝_a�Ug����C�{>�����PN�%7n\�>���eozӣ��>�1[����jm���߷]x���+��^A������R�����A����S����~���	���N�>�x��/|!w;����S�Ϗ�����s�C���n�w���[[���x�O�i>��s��A*WP�g��|� �j5ܮF���}誒kex��ܞ�.����&|�`����c�o�������}�`]��Ua�γQQOTR�~��i1,V�z��Tg�ue��p�V�p������d<�pR/�l���Φ#�k��>湝w����Z��.�Rٍ'Ũ�U�ʔ�d\k�߅��p��KK]����G���0��0p�L��²;�k�l�Bh����T�֥򢛸�ȿf�/�� �#-�H�Ze8��ؿna���a4�;�����h��.��z}U�#գ�hv��UY���Q�r����e�.,S���J�p]���H�ޛ���"��ӑ�׶�m�Ӡ���0z�j�Z�=�<�g7ڇ9���+cYHh5���Ia~b�:���F�5�Q�؛��g�C=��6Z�m�FC5ҥ������?9��nv'�����>P�=�����gvm�{<ֈ�&�N�d��Zy�r�� �s���R��Z�.P���.$��F��YgW����Y(Q}�͏9��c'z�v����=����O/ok�͕�V��̴*�,*�k͵�:�(/WK?)�Y����9.���vm�r7�t��W5�U�����3,m���}���;*�aҵ��j�׭T�°/KhZ����	����׼uQR����lXX(U���;�"����FWU�b{Q���~~gw��#[-�J0��:���~�C*E�W��[�I��`gM�+?~y�k���RT�T��*�6?�GV��'��K��g���� �{n�A��o/�dW-NN���#�>��3����Z'�O�:]��|�w~�^���V��<��4��>�����+���F���
~�Bm�,��c�>{�����}��
�͛7��.��}'�>��(T��'yY����'�]��O���F���F�<�����y�k5um���R5E;���ג�������U��u��v��R���^jb+�R
�e��[�B��Ë>w���+{������Ǻ�?�uV��V������
T]�)'e5ҤH�6��f�ە�J�U���ͺ��u�6�r�3˭��;`6���ד���J�^� ƅ6ݗ;@ꅪ��r�kH�R@�{?���!��r<�-gt�`��6���dU�����v=+	���mA_W��
�Z6���v1ua���/TۨI='��b�,l�˼
���^O�`p�L�Z�B�W�%���Z�ki.��T�e�HR��.7�Ye\_,������)
kU�z�[�B�0��9,�k�]��vto|�;ռǉs.�BI�}r���[\���j[��}�ф1?�V�x�!�BW���-�$��;wl�1��j�"I���bxNH��]W�ߋ�=���ua�طe�ʥ��h$�VԴ��:X赳mJ?�����Qͽ�*}ow�����8ʯ�U���F�7�j����0*j���6:���etUN1�Y+��Nq�`���2���g�6t[���okͭ����~Jj�m�X�3v�Ѯ�z���MV�
u񾋎o�=��T5Y�z����DfdԜj�˰*_:����ኇ�C�'���'�d/|{�/����2�*���0ʝYK6��2�v�����U����ݣ����v��:. 3L��	m7z�vw����fy���m+X~��+'�&����6l�m�阌g��sV\�t)�x�~-M�d�0/��p�6�C�{b���'�_�Ǎ����w@��;8�B�����˭���bq��L�Y��NQ�swBP�����U*�즩������U!R���o����k����z��%�Je3*;����|�����Ε.�V\�Y6�|���D�9G��x�\�)���=ϱ��U���_��>�Z���򱆖G�������wO�P�Ne�/�.�+�Vlt`;��*Ս�V�w騮���8��Ġ�:k��w;�;zL�	m��7z�Ʈ@
�Zz��?��4qb�O�6z\�8?�
���n]��l:���?r���e%%K��X��2o�1����/�>��2��5�b����r�T��B���Cªk��J�����:Z���/�+�k�g^��䶹$��ȺE��c��hq���d�Z��t�l[jw����ͱ�a''�]�¸B��&�gu���_:�N6t�7o�*���7�������m�����wAN�.�w0t�Љ��}��J�G�_-a� ���1.��R��[?�����Z�����6�#��M@��ˡ�%֥�:p?2�Kh2�JKT������e�c�m�Fb��]���;G��´�O��}yS][�DkZu��bi��z���5�k�����+jwם9���n<�;��w:��N'�;9:�"H�4/ �%�����3r�����?U<��ӹC��������b:��߼9�U����٬)��	�:7���:�t�|��M&�������Éf�������-���jݪ�{ѭ�z�v����M\�i�]][#�E���{U+���~�Ye䂷�na��*�f����42�:���Z�C��W	mm"Ug+�V]V �]*/�T��jՏ4�%eM�k]�rq\�>�I �݉���g��Y��[��
M�T9L����dT��B��y�W���ڿ��/6K��|����ȯ/m��*���b9�e'֍dVN-�kVd�꤭�⭕�_�S��M|�|���Z�t��4��N��ltZe
�S���*����M3ȭz<�mVوB�F'U�������DA~ݿ«~N����	)�k_�*i���9=�z�P�Y��k��@�b>��=޾�C���Z"�zl_�۬�䶢/3_z����muӮ���ӎwX�_/W��r�o�^\-n{g+{�{�Ӻ�^��p�����^���4�m���>o����E'��Yx I�ʁ�Q2d�����[��:���-�իWs��k*Rِ·��u2P�՚�.�۔@%�X�Y��g˝i��c ���j�m�s.g��F�3���w���~AŮcfGu/���S��e��KW�ɸR�t�q=j]��J�Q�
�#tv�_���Mf��h�����j�jJ��ʅ5���e��W�h|�n��%�;�7���%��U�}�%�G�ܾsх����ڭ�;w�&詎G^��e��ٞ٤?mZ������I��A#�]X��Y�}���������g�J�U�۵��_����_���bP���В1tɇ�PUrR�~��F��R�f�-������s��I=*��/���1��{����q췽�Ym�vN6FV�� ��}����=ԣU�^����}�}�{���U�� @B6�����'�xBu�ťK7�+W���ҥKZN�����=�_�q�G�o\t��ֻ;�`ݮf���/�NQnXU�ޅ���h����u��뾿�:,Ha�.�� ����y���f���}��u��E����r��[8���W}˳���ѱ���F��a�X+a��de����ۡ�����Y�^|����P�j�52}��K�����N�ܹ�}�}�w�����o{��܏}<{"� �W����|D�j�����8��S���?�ښ�vaq_��Z����Y�����^�Z�Vd��tb�RT2bەZ�S���>�h���CDVՓXFP�J}ٰ���n�{o�f��X����5[��:;�g�=Y5o�~nj��C�a���k�v���i����'�O����1��6iN^z������l>����N�'�щ���Wj����  �&UU9���z�ﻇ���r�:��ՉJ��^-^�C����EGf��X?�.��q�Wן�ާ���U���7C�Tm����O��u`P���ʸ[}�:RX?�vm�42ۆ��OCl~��q�f��G��ʆ���5^�p�կ}5{��Kٵk�*u�p' '�����٫�  �&��}u�����J7�U^�eЭx�,m$�:A�e�.��DFg�5��j����2�( WUjg�0��;�����uU��)��j����\�=88��Z�������B�V�S�՟�<��a��F�r�~���k��_��ް��ݵdu�͸�y�{��s�}�v����M������:���U[?O�  �I�zy�ח�syk6-�_�2����=����UX�x2��+�b��jzm���:�e�l[}�߁A�q헶�ä0��R���؊���6�*�H�:GĖj�E]4��N��E���ܲjy�1��:e��yb=�Cp�#���6�¹�����*[eP���uϻ�N'ŭ�7�w���w\�~��X� ^  �T�e=�͔L��]1��u�ڱ�""5��0*�ynm1����-�����*�5�©"�:,�!~�<���6�,�u�����\��K����[���w�G�m�؅j�_�<(�n.�z�XJ�Gg��|�/��������Ϊ��\X��������5��*��k�e�n�{ӛ����UNX/  xMra���W�+��В�.���ɤZN�6«�`
��ԯ��[�#�e
��@}qmB۪�~�}a�׺�s��yc��_Y*[�պ?g�l��kCɄ��(����0q���8<��ϙ�]�ޠ�_�dݯ-c�ZY�������%�7jt�J|���Vh�ʾoK~ےӵ��w��������n��ˏ��-_�߻�^��  �5i4?����ߛU��k�^(��>غ�W-]hti�q�֤���[��j���(����hh+���U-5�;;��Ivxtd+��!HV�-�l��C���о�86C��l�e�Ȧ�6j?Z����Z�p�.t_kwZ�d�5+�]>{�Lwr2/6WZ���N���;Ē�\�~��S���1��G���w���B�V�[,���b��"[�J�r<�74��({5#� �פэ�n�x�_���_��|օ��;;��X�E^�p�J���j��{���P��~�+OW_��-�?�U��=��}����p��jaU6�+G��C�-Y�YX���*��Bo�0�M��"m;�W��teղ���[���!cF/�?Ѳ�UuG��Ԏ�]$4k�V5�[��j'V( �0^�r	�f+��'��mݯ-�<���VMS(�7��m���s�����j�*F�  �I}꩓����o���'�5��v^?{�֝w�{��ᡋ��I�jڲ�o\����hl�4M����|a�pU��nm��&���I���8�,vP���;�uZЂ�������CnKǮ��᝻�����+�����qպ����z��o�p����7=U��Ϻ����ϯeYw�e�Z���h��������t��۬o��UUu
���c�=6�~�����?}�Uۅ�OC�  �YO>i!��O<��ŵ߫�˟�;{��~������mU��Jn޸�����y晙r�xRg/�t=��̭NV�7ͪ�h����Z�ί̦%����*��a��H�3��ժlBAX�x�GV\[�n��K>�-�������j�TZ�򥋿��{���/��ɫ�[�
�  �����~����o����?qt|��.�~�}�Ѿ�Oܟ�������'몢����c������\X�U[lmo�m�~�
�y�}V���eEy�㰺]-={�j�7�]4b�FtZp��ߡ[�Bs�vvv���>p��d��  ���w����'������mko�߯�w�}��.y��駟�w�t{gw�p!W+�������Z��N�[�:�3�(�Vck���:,����wJ�����b̀~_u��z4d�u���md8��\ݎ��WF��<��"�  leG���O|#˿����ݭ��㽝��]2}t{k�m[[����x]Y�g����z<�N�˦�jc-Ȳ*�4�ۏ+�u]������R���&��|A]�}�v��ڲY6j�[�6c���ޗ�u�t��E�  �.B��Q���Ͼy���'F]wg��w~k:����j?��������_w���z�jh�]5�Cז��Jf����%���ٺ�¥-Q����E#*-a����V>Q���Y5M�T�bk6{v�/^���   �z��d�B�Y8��>���?\]�p�>:��ݹ�X6f��}���s��Z�u����e��y6�N�f��J�ٵb����K��:�땅\?��N��_<�]Y�����lo��l���gxY^  �?��a��O�z����z�֢i�Z�L��>�v�FE�/gp!�V9ú͖��|���z����4q�~W+���$6��+{(;���C����~�����/��  �=R��G?�o�m_�ON��x<.��R�V�$h�Zۭ��A_�hnݏ�f���P�n�ZݸR�-F�g����#��V�Oo�^w����u���  �}жu]�#���B�vb.׶k�f���]��[(�6
��l�}��P�տ5QM����il4Woom���Z,��s�ۑ�9�"�  |��=�r����^E�   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   ��� ���=ׅA    IEND�B`�PK
     #{dZt��n� n� /   images/c750f18a-9432-41e6-a6ed-179e28bc29f6.png�PNG

   IHDR  �  �   �  0�iCCPICC Profile  x��||eU���4�K�ҹġIr=g��3�0D���d���B&3�F�� J�6H���U)RD��tA@@i�Ҥ���}�>;p�{�{_ s��Y�������M����/X0gT5I��[4�=ybuϽ����j2���l�l�?�pAKWWG����ٟ�O���f+���Yw��$iX�_1�`������.Z@�ĳ���~��a,��D�r���'�7q<�ݭ�S�d`���!Iƭ�?�ha��������sA
z���w�Ag��3�dUH$�5g��!��јs��>7I���xV���=��f��[��&�I�K
:߯��uZ�ؽ�RƚS��L��uRu�Y�����m��d�6ei:0c.kb5֔i������);�u����:{��l�tE2-�JX"���'U�)~YҌW�Yb�ڑ�&��M2+L��w8J�m�&�+p���	���@2#��\��,���5x���o�k9c.�8K0�vh�M�����,<h���_�txh��E�h�`�}�@���'!Y�m���|��_z2�%������v�EIҶ9w�m��$��$Y��ض�N���N��� ��)�J�����������i�y����������ÆU6o�5��phÙ�5<�����Ge���:l�壞]���F_:��1��sƘ'�n:v��+��c�wԸW�h�y+�f����x�-W��ʏWX�����X��v�z�j-�ݺ�^��5�Z�5�\�k~�ցk}����[�u�Z�����{u�ÿ�ᗮޠm�?mx�F�lt��{o2f��6����=��q��-�-no<�˭�O�ݖgm5��v[��͵��������v�4�nީ�^����9�/��]�O��9j=�t٩�w}m���qh�w>��g�\>���&�}��ڵ�}����η�n�պ����z^�6a��=��s��S���o����}����;�6���l֑�ٯq��9�����C<3����o����6X��u=�;kv�ky���s����{_?᱓�?y�)��z�gu�g�朙�t��:/|���_��u/}ⲫ�8��}~�r̈́k?���~~��1��]o�����|����u����{��'?x�Cxt�.z�wO5=s�=��S^���ޯN��n����ķw~G���?�~��G�~��S�bE�W��h��(�v%%5�6\?j�QG�zs���>c^{�u�ݴ�����|K��U�_��ՎX��5��y�Z׬}�:����^_����pˍv�x�Moz�f?����+�ɗ�4�i˖��m=k������������jO|�����C� ��5�zzc��m�~��e;l��.;u����9��֋']�v�.�O~y�w�1v�M:d��S�N=�����~�w�������=���G{�������o�}���a�)}3�.�y�o�>n��]��5s����濵���Un��i�Kv;p�.=��C�:t��o����=w��G�rT�hq����y�������N��K���ם��S�;��ӯXv�?����<דּ�>������s�>������hᏇ/:��.Y𓹗�\��e/�抵�l��ë>��㟍��r�:�mv��?�7���q�7��b薅�<��cn;��s���k~��_���G�z淯���=����}����^x���=��#���]������.}��'~��<⩅O��̴?�?�ӟ�s�>��_�a�ǽ4��ѯ���J����z�����ߘ���[K�>���s׻Ͽ��?7�`���������>y~�w�'�jأ��Q��:fԻ��F�4f֘��9n�qw��`�v����ݕ嫜�ꉫ����k\��kݲ���<��K������6�����I�-����S[���q6ܲi������>�.���۝�����n��}����5����j�+�U�ۯ���w�vG�S��S�����o=uҏڮ��7�����ww�tl���)�St��������<m��-����>{�����꛿��?~��}��o�o6�6c�`�̡Y�g=t�~��Ü{�>=��ko��-j[�ǒ�|�	K�;��Cn?��o���_��͎dG���1��{��w�����;�֓����'?s��p�˧���3���;g�w��gp·?��������.���O~��"��O���]���n���+N��諎������Ӯ9�ڋ����~�����MO���/^���|��oo��r�:����[�&�k�߶��{Ϸ�uߜ��<�߃s~7��A��ѿ?�ѓ;��?��ӟ<��{갧?3�O��N��n���|����~q������{�ѿ����������/}��7��u�������#����7���õ>��/�q�'3>%$ё�0y�aR�����g�=�����4���د��y����Y����W�p��*�]�U/X����Y��5/[뺵o_�u�^�o므|u�)/�d٦7o�lu�[7������n���m^�����mڮybm�������旈k�m�^��y��u��v��:;m���zGˌ����>��_����o����&���=:�N���[���ݳe�iӏ���=���{�����-�5�o�>�����w�xh�ə��zq�[C��ڜM�6��i~ׂ�>b�E�.�Œ��Ao����������_r�)G.?ꎣ�8��c�[��	�'���yҞ�8y�)�O=�CO�����8�ǜy�Yǝ}�9����sO>��ϼ��|�Ew\|�%��ɓ��q������^qΕ'^u��G���w͉מv�9�����p͍7�t��w��[~��'o}��n��7�|�W�z�]�;���=�޻�}��?��Ox�����C����;�������ǯy�'/���O����gN�ӱ���#�;��#�r�G��ݗN|��W.��e����]{��}��7�zk�w�G�;��{�{�޿��7}p�������۟��ӏV 9,��Y^�2I&�+�zŊ��In �]y��X�ƁI�J�r�I�����/I2��I"�a��G�lu0Ǫ9.͹�g�[��1������Ã����&˧����,�wc�}�J;�]�$#��j��::��&��F�$����{_3�m��u�:�����W���u�� ��};0{�^o����+r�����)E�=�?�Ư�8>=���z^�3�b����F�6���������_��S����|=���+����;���^���h;s�{�
L�K҇���������%�����Rp�8d��-q�~!8�'�������}�[ ��@����I�ecv��2��	iN���V�c>�~��Y�b���E�$�A�¿Sѫ-���c�V���E��"7R߈l��R�ԭ��D8�en~&�v��d@ݠ:�\��1�K�����T�2r�����>��9�ƚc����܉��rO.æ+l�4�ɠ	|D'Q{��ɠ;�F}��CCsI�K 3�����e~��ɛ4J�OM�i�����D�9���?�I��f�K���s��)�Jad�H��J>Ӈ$�ğ7��6�s �m��9��|_�P���Bг�ۺ�S�_���c���3��B� K�9Y�w���j�Z�Lj�i�n���]ml��tΜjk���}��͟W���5��:0�xQuh����s�?��������SZFv�1�p��`���Jkw[KoۤjcO��jg��*3��n/�����@#�����������Sm�����ѲWc��}�䎶�I�}=�m]���pS;��&w��U�a��i��u�S���ۺ��ݓ'��7Vz[�'����O�����6��ڸgs�Т��PV��%��_�5<���:�������
�Xe���޽��0�.�m=�V�L��_&�����c�Yc%N����������#��1�R���cq}��:Y�ъ��2cҪ�5�5ci5Km-S�2�X�2�����}�I}�S����ҴڸW[Ocez����}�z�Z�0����}ꔾ��==�;�<SebN�bث��"�Ꞻ��4/�60����Smn��WBI�Vm�Y.�Q=ph�� LS�5S�5^�7���|kgO�ղk�6w�0G���J۔I�sW�N�i����,��p�� ŉ-��a��{۔�+�������uLkice�v�O�D�♋�}=�^�����9uj�#��Zz[w��i�}Z���8�����}�1F��)X�E*Z�2�sb[w6�K{[Ǥ���"����ҷ�Vo������)ib��w����$��t������	id�s����T3-G�Qɠ�1~J+k��\����i#L���k�^ӪQ��ǫV�O�*V�¤������a?Y�[�VFd�qn�`�Ƭ4iEUY�M}?V3BI�5ոVFq���LY]�U�~a����LUeM3�-�'�L���(��~��ha���L��b���IU������Q�Z*YZұز�5�	a��B�X���J6Bc
��Ѡ��Y���m�Y�Ѧ��P�BFEG��ܹ����9�,ȸ�Ry��Ŏ�f���F�ʤ��7Y�����BǬ�f��g�3�lUԌ���ɒ�/Zp�f�N_gF�vjP�D%S%�X,^��2LB�X���k�Ӫ����k�X'3���괒!bߩq;�<u�zf�x%�d�q��,SnG�'�&,t�ɘf$%e��*��ki6n�v�-dꦖBFgj��SO[jݑI�2C#hK�
cU[3)�d�uؤP�#n�V�XF(�!ѣ�l&3R嚐q�[f�d�B��L���|���Ab Ў�W��f[=��5�j��j)穵8�LèI��	Vc�hk@p�=jJؔC�X���s�#�V�T�t���3ȆA8-�IE2�'8y*r��a��Z�{���9�:B� ʤ Xʍ�E��@9df�&$w=c�%<F��b_
��% h8"��Ba��B�T�����KY*l�c��9� ��)'�j��E?�L�q̎�� [&qPB�W�;��4�;�����d���d� ,RK��:���º5��4�� [
�0DHÍ�%
kf���ּ��yF^���[XGF�ь8h�&�z��]��?"w*H���T��#t�f�`cF]�p��@i�ƒC�*>�ђf���Z����j�6�C	]`�P�`uذY� B�pR�`M�*���*,D��o~/��B�
��YT� E�JK��N�L?������*ظ���S�:f�8F�PV8d�?Ο���J4��J��NW�v�G�TR	I�($���#����a���� �T��x�x~@��_�?����$oKl��T�!~��
�e
�!UCH.������掟[�*�X��E� M�YO�L S
���ʤ�����ai��8�=��j�F�x�bh=�_G��X�!AG��=�8�
\��F*]O�_�ʪ�L4�R*%:�q��C�u��J.Hi-t#E@b8[��A�g5���K�0qR�h#*�mj>��1#�
�����(��U`)���f��4�����eI�d*#8����0�#\��(RUǑa�:s@DV��A������Y)L-�\ ����j)��i	A�s��l�"�fkLW��X��#���O9Kx����VTV�H(,if=�I��;H\��W�<LTUplG���X	��!�1!��W�a�ȴ��)X=~��q��R �!-K3f�Q8Z;�:�8�����	�����T�]->Gb�<Ӱ_K���#�a5 �J���� �����p!��L订tI��2�
�ǂHL��A��V�$k�3"�"_�(�XC@��U�-�tbn{j��'�2�'�Y�NK2��#�I�ӌ2(#,�4�9�0}G�Y#�i�>�I�֜�
�]챾#���52S#�@�!G~W�|D�V���4yE
��^����(bG]vD� Ԟ,����@��;"�"�3�� T����G�V��f r��S�=DNxI(��%�c<J��g��C �8d�
�E�X�,c�Ȍ3�!Ht��v�+�p������� �G�)���O"�Ü�w���T	y i;�SVǉ�w�PC�GP�����XMY!'�,���:*	KhP2a��Da���52���
�ft%��E����F��$g�h�+F�LU��t��N�G5
���J:�� �q�+�S�#�*Rl1��u����#�� �I���"	�5i�TS��8#8r2J���w
�Z��g+��[�r))Ȼ%՝�g�����;7,�S�CV��蘕t��E�-B�ȕ��(�{��8���+Z �U���92J�,�#��K�\���!/�����ci٫���dq��<�"ˈ:(R�*v���g�W	Qc�GDd��C�xŪ��q���3��U@yKf�t]�Z]�G* ��l�Q��Qb��8L�{��  �0�ܣ!]��RXA8��=i9`#�9(�$�X%K�JN�`�6�4�0�Q�)�0W�K���q����*y��3���e*$UY�k��6-yEr@���E�'/�Q	�R��3�Z��SO 	�S�8ר��ԒsEz��
pU�Ҳ*r�
���Uu��"�p�!_�,�#=z2 rIՙLH�:zB��YVI�;W����hW?����LQi�,�%=9e�j��U��L�h��<���R��!���^ʹfM0������U �B0����Sp�焝Sϲzr�I���&�[ 슞6E����@� @��S8l���|�[��%&%D�V�Ef�jZ�:/�P�e�SHq9���ef3����YS��$?��XC ݅=J��S�t�� ��y:�)S+��|5�S�8̸OlN���Z��*�L����\a�>E��)��b3���%=�gJ��$ y0U�e� 
~��)�H`  9-S"�b�*?�
�J���UX��Bl�ʗ��7�m�X�׌�-����΁g�8�Oդ3V�T"��|_J5ɼ,��<�A�p���������T�cT��2(�S�x͸OE�{�}S�P��˩�*�Q�YXJص�:�q
hK:�t�׌*A�A�aC����;$z$[S-��T-Ȩ��<�(B�`z��W�ȸ�<!)F�;�88'��iLaw�)�r�%�m�M(�A� q��srK���䯩䋸B=q�4'+�&E����+6���O�es^�腨89h���a}�p��1�Gb�ěD	QL�CaܥS�K�M��"�/�Br���.�͉@���e0:j����8���BZ(�WK�_���C�r�*�ܳ��sSŞоT3W(Fz	c&}$ᢧ-s�EO���v%`9MVj�S���x�
��j��,S:�0�Ŝ"+s�&P��N��W��,�4'#ۣ� i	���˥$E���$�P��*T$�W׸Z�;º\����'7��S���'=(b����$��0Xz�Z��G[!kԈ+TK5�x%�7�C�,�Q��3
�b�=�R��4ͩK�f�}8Ah�
zJ�����>iNS�3��܄_4RN@z+l���O8W�Wm3dEyOC�V�W�FR��t?��!�T��n����(*K�=����)�i\
?$YIςPT+��Q��|~GB��o%/��'Pa�e�OY�����
:O)J�mѓ�H*�-��~���S�e�z���Sf��vi(�&����*�7L��S}���sJ�td����9��� o+M�xx=M���=��m)����%ϟ�k��rD-��'���?#����z*	��Ա�L@�F� �S��2�ZU���2�e���
=r�\O	���e�4bO(�v#�g�)��ڧx�>?�M�>����."I�>�x%J�m�Uc(��b�e�."6Q�$:D�hbȳf�8�(.2F�UeIU!3�-��r��I��.wP�T]COK�����(�ʷa��iʂ�HM ���%z�A}ᇔ-a�&dT,����Hm�3�X��t<a��wQ�L���f!!=B��{��P�E�[1��srðOw#�\��OC���&��4��ㄤFV��{RI8e�e��pW����޴(9ƸO��p@'��Ru���a�?�,E���e��hW���_tv�������\��YԿh����g�~��&�a���&�60�ڼ�]�i����<κ�<3#z���fd���.�Wm�"(k�A���DS�=m��F�"a�yOZH_���̞?ܷK�ܡ9K�����9�6V���y��3�,�$)J.I�u������:$����AqG��/"/�3.")�P�D��I�+%���N��4���s���
G�	N�@{T�s�tBrOr�kQ�J1����s^ʋdn~�����
�bD�Vѣ=ת�ԅ'��V���xΖjp�j`&6_��*��Z������"���ka'Y�*nf�"�"0:��VpOJ@��D���/-!�[9���9��y^F����[%�Q �bgN���
Z���I���\Ⓔ�`)���)=�w�6�.<���� :�|\I7Y�٠T�I	[�I��+�N�X����ړ8,��"E�o|7x���D�|�*?�j���y��X$j�K?���ڦ�T ��lVӅ�ub�7D7И�$���f<�p�p�g�y23~9\J!�s��µ
�$�=��S�R�x�SʜA�p2�d"��#1i.������nk��ʲ|\K��/�.�z��T�oSЅ��
�ΜB���B+s�c���ɒWZ��߬ĺI�s^����z�/!g�w���*I7hB7�p��(�V�a�He��F��ש�k�0]�y��m>?�N��4s�3��k	F���.ʵ���y��qG���V!1H���ޜ��W9���Q+F�{iSF`,�y/Xn0^x������x9�/�ca��=���n�:�vG�cR��0׹�g�:�
Я }���0t�����$l"�֑����l�6��e��4��5S�,r7��Z�7D�L�)�dΫ�a$>�d*�'�]�mf-B��L�3�M��.=��/c�K�&+H�ϋ��x^�_�r�&����l7'�<�t�U'j��f���%��$+t{>��M3o��OrxaO^f��r��d e�I��k�BԊ���$�?OJr0�7Y��t�/Ge��h�yU~+��;Ox�б�e� �I��#@��ņ�lP�p�Z��D������o5�ҁ޺q �Q:^2/�?A'�����ij�>��0A�#��:��n;�1m:'S�f�(����"g�	��Xa�] ��q�EC��	`�	�؏_o�����If�m"�k���aTު�WO($}�$'�.��-��3���������8�u�3H�K�B��a�o���/���ɃLM�g,wQ��4~�Ț�' �q�g�P��R+�R�Y|B ò�/����@�ԏ���U2���LN"��2�!L�j�w S�!�x�͡�k� ���]�yE^|u��e�daoPz�=�.>��$P���nd����=����l` 8�,�Fn���G�v2���x^�q�IN7��@��|�:����d�ې->g��'�I��Har��a-�Rxs�Vi<o�a�+�d�H���[`�z��-H�M����c136gl�'�"����[��`-�����#�!P��=��x�����_$���Ъ����pd_ގ![�Bk��"���iV�<dV�E�0�
�ړByA��>�GC2l��ܜ�{��E�s8�c؈ិ�0��O���!����GC��k���M
?n�04��K�PoZ����f��H*>y��`�ګ'��29�,�y���/eY�J!9%�~o�P�	�H��i��e�-0�A�0�)��4��F���JA$���Y�0T^���#��~�Aw"��,�E"S������p�I�V@�A�HLe�-0�x#�=�@�H��+"��4�_����$�3������37)������r��P����W��7b,�y�J��.�n ��[`�6`9څ�d�������i*����,ƍ:���d:�Zd1|�����0BF��y#�A�-����@���SD!)�*(y�D�`��FP����@*�㱈F�-9�)����*�Ǎ�4�)��$f���>�C]�����y���)�T��h�~����j�L鲤�!1�T��k�8)a��"���y���. �O�мJ*��]H���-0����"􄳠����-0��"����SD#�"���ҝQ��"bZNx��J��""��r���R7�������z'&`!AS��z#��r���	��� #��/���,N�
=��~��s�Ҳ�MK�d�0���Cf�WK*$�� #���jH�}�L�/�Kd�0���AKp���31ր�AjH:{�[`���*{B�r��R�0��a<�3_��HB
~op�*�@�e<o�a$��F�,'1���X1i�L)
^���[`L�y�	Rz�̥����'Œ�����,"��x�R���I�"����t ���T���LF#I~i<��`,�C�0p�<,�"��Y�k��;��6Hﱲ�Fҧ�M ����RF#��&�Oh�$}3�?��a�jø��ae��?n�0ha\"�{�#���g2b���1-H�nR�5D�V�C7(�_}���E�0�B� �����qHE#)��k�\�Ӵ�ۙ�-0��)�@�l^�r��Ak_@%!�c�`�*bEϗ�'e��L�����n�R�|�PT�����0h�60���E�M��ME�V�����+�:��-0��}�I�;�4��51�b�� ��5D覥�U��a��7��>��e�����>��ɂ�`��1�B���Kc{Ni��g*bzt��>e��L�:��F�"�*�~\A���Qݽ����Wi�㨈a�-~oT,���|�FQ�xeȥ������Q�� j>�(����,bE�H��sR�1��;�Y`>�S����(x#���>��ی۵>�@zg�7R�V�|#�Q�t�,I��cU�0вP��Y e�A��a �{U�wiC�JE�H�K��}8Pp+���#����>	�rU�>���t�0��B�V�sR��L�y��r�kH�L���mSGC�"�����ߟ��Fõ����z����!u�0:+�6�����I1�~H�z��`��T1��;<�Sa�_���#����T��9Ĝ����u�0�2_/!��S��a4� (*Vx����5D��t`0�q6Sޟ�a�ǽ�k,� ǥ��D���xՀ�Ɋ���"��{>��d*���U8ވa0��,Aѧu�?��a0����3�� ���[t�0�By��]�$=/�y#��)T�U��G�
�at�0`�M�&?��K�9o�0�"�IMR�:�,1��>k�;�wC��"��/T�PBC�܌�>���8P��k��	��� S�����G6��1�h���n��Ve|2àU���7_��{)a�à5�=M�DњW�+���*�ޢ�L��u�DC���Az������0�����k�`��M�0Ԛ^���'��x�DC��Гh�a���k��Z}�0t��OAy��Y�0����!p, ��#��a�+���+�7CUO���a�*}ܐ���5h1��ų�����F��̃S8
���{�4�CX/�C~
X��C&b0��y@=V����a�|B,Sa\j
&b�T�wW�N^�4��Fc���npaǀL���a�P(}8!���-0}����@�#$=��5&1���VNJ���31�=���N��!rx�c"�C(�������5G12;�i�1�p��ڲg���..J�ڕ���z��Ga����0`�a�t[=o�Y�-0�!ǔy�,�P=�l�7b��1 �I�5�וm�0��(/t��>I_��ㅍ(����R-�J����0H+C�e�{��l�.�y����=��Ґ��`�٢��RӰy�_}0���FC��s!�����6b�!�����	�[`K_n�7ρB�l��x�EC��}������Nů7b�d�+D���c���0�*�ab@5/_��?o���	�Dz�˼��xc�K7�
����'m�0��f �T�����:��o� MW���0���P��ǥo2��1���p�A|p<���gB7��AJ؈a���8����89����a��o���{:�H��F9o�a,=D����@��g��ۻh-��ņV�R�x�;I����Q	�/�   	pHYs  %  %IR$�   �eXIfII*     (           >       F   i�    N       %     %      �    �  �    �  ��    x       ASCII   Screenshot�j�Z  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:exif="http://ns.adobe.com/exif/1.0/">
         <exif:PixelYDimension>1018</exif:PixelYDimension>
         <exif:PixelXDimension>1430</exif:PixelXDimension>
         <exif:UserComment>Screenshot</exif:UserComment>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
�v�  ��IDATx���$9�&�������iqo���νw��o���������.��*"3�+� �if����D�g����H����"Ȕ)S��P���IɺO��Ӎ4�3f��dʔi���7J�9T@�L��'�j�/�����{	����>�t�'�2����%��Lg3��p9����%m��T��̹�����t��1|׷�-��>���ʲ��o��s��9��nT��5�듸�j���e���́��y����W�[m�����S[?&���]	׵�p ��;����{����{{{����N��bd-7Ӧ��2eʴQ�Wܿ�9�U8�Ko�L7��������/a���2e�t�D ����qJ7�%�@��Ι���u�u�wd�t���d2��dR��@iK��fpyy	gggpv~^��x��/�M�Zkk�րb��Zk� ��N�Z���+@���_���cҮlW7njS|�g	�=��&kAZ��nX.���!�����>Lm�ڶE�r�����-�kI��P�3�"��ɚi5���͓Ъ}�����<V	��s�S,#ڌ��)ӇNm������^��+؀��v��Q9J"S�k$��+��1���<�p�F�y�}���p���M���*���fO�L�6C
�t����޾=�7o^CY�Q���`2��t:�Y9%�`1py�a�W�2 �j!���|��21�����ٗ��]�*�y�uP��.��; Ѧ��ha]Id��՘�.a:���;x��&�1ܻw ��{�������q�������j���L�2m�l�wM�-la�5��G��HO"�&eʴY���R�{Zp�>N<�~��mGNxJ�6��)��Ƀ�b4.x�/ѫ�R���r���p�� �g����;mkk����`�����2e�t��,��s89yG���նi���Q:	x�).������gڛ��hP�0���Z�x�.I���,�!u�Ν�ArJ�ǭW���ɤ��鷸~᧸����i�6�i��5��/�5_�>�lf�t%��r�L����J���=�xذ�"I�E\lM���[��)ӦH�����4�&�Zp� ,�{ݬmU߫���B��@�c��N���&S�5���GQ�*�2��d'�� tqyI^����0ϫ�E!��Ng������p��=��ݭ~���.x���r�L�J���������/?�L�ɘz`ww'�_<1,�X��M�~K�T��ۃ���|ڒǆD��Ɩ�g�$/v�M�����i��x�8㨿I�\�ctLk�fS��Ǳ����,gf�4e`9��f����+�-����:֔���kY�]���Ṕ�%�&n'�4B1��^�<~𡭆�e[�8�)22eZ�7a�	Χ�����K���IQ��</0**kUF?���Ua��K�ٸh���߃�{�mooC�ߏ�a���C2e�*�:̙�s�c\�������-���g�y8����4G��)��"VI$ռ�:~2O*�xF7���ނ��C88���sl�O2eZ���s���W|�ů���۷�; �»wS�)H�(Ȁ����Y9��X��������*��0:���_�}�^i��F�k��u�����u�w��s�kjq��a��M�_޻�Ҹ�Ϊ�9��3��5�	�6KX�t���c���	��������|�n_�´�B�'K T�\\���$}N8��=r]�k���e̆�T]�~�;��чK�OF٦��y���.���y0����2��"���+%��g-�����s�f�t5/�K��=��>8'�#�2�!ǲ������Fx?�j��z0�T��=%'�������3�� ��2���+�*���@e_��Z�G�E��<%e�Zɰ������ل75��8P�qL����vY\B��O���yMnmo�\�)S�Ť������t9�''�C�[y;���l�a$|JGY)/e�S���^(n�t��ϭ�4���n���k6���u��]x�m��ܮ�:�TȠ{*���H��ׇ�VW ˗��e�$�{ L��5��!��'E`�m?~h��Zuw}�3�k%����*�a��Y9mS�N�=�L�+�m-��	=�%�K�Ks��g�.�1�(4�-z�{���Xm�~00{�г(x+���H���C��n���<~��ާPS�Yȡo���1Yiw~1�D�2��)ӕ	���W��c�9�Ȼ����;8o!.)�i�8��(��RP�=�C���7���􄼖1�=���2]3��=�����Z�����������<�s��ɚ�_x0�* �1%C��A����>.w��$(���mG�H����a�Ճ2��)SJ�mB����s�_\\���#x��%��>�:A�A ��$�`�d�Rx��o�lDw���B<�k�_��t=g޵��7�Zl���wTxO����KA@¹fG�R��xLM77�=��6OY"�t���-5�r>�	Z�yGKp� ��,�6`���m�@fI��ֆ}~�W@mWo��y`k�h~��L��j՗��oH�W���4�#������.6��©���a(^�'��I���1�y4��^#��=��Pb���1���(d��DE/k��w���s�YX̘r�L�!���g��.<{������^��2��i`������c8�Ga9�E!
ꄞ�����C����ڜs�fʴNBOe_��x���V��݅��!�$�� �����XpZ��M��eT���z1�2A~2�8�bO��-��Q~�|��sywo2}�tݲ�{�߮��֓��.v.3A�B��R�����p~~NE�&��$���ԋ���T�"�RЃ�����4(��1�r�1��F"�`��W�t���)k��Xވ�c ��4�_7H]=��DN2|��+B4^���h��EXδ!�j�"��1����x(~��V�T~Ɨ,�;�G��@��;�O���=At�m�%����ߔ����ay��b��d��\>TK��i<�� 8��X�a�Q(D�e�,Do&�>�|h&2���s�Q�Lk%�⁇sP ��%G#xc�Z'-vK����Y���k�o�0�z� ,�3ɔ�Jd��QJaGF+aT.j�o�7�<(��P�=%FS;��T$�y1廓S����ɘ�#����a�953e�Nrr󭦖����g�T�R��e�NF�T����߅�`���s�,,�;�X���2�)mc�%߮wV���<}������t}�)�z)_�|/c��27_�:S�Ŕ��L!d~%y��)����c*���%F�^�ecλ6 qN��I.�u��R�I-Qcn]ˢ���2���"��6Iv�~3���Z�@8���8#%��>|T}ܪ�8��]j�L�2��pN�1�z���P����,��bW�Z^���=lL�������p0������>��ɔ)���_�NO��~��J�D�yk{�R}����.X���9nQ��&^sS�����3�$�69�!S�VЕ�OOSx�q��^�xQ�`��tz���wn�"�81/z�7P�i1X�)��I�r�vQ�qD�]Nn��V��t�ɍ-�ɤ�)�f)˙��R�,��Q�R�Z��S�������~ţ$�]��,���mL�Z\�����;9.�A��$��y�	f�����l6��N�縍a���N&紭�3��Ɉ����Tc�男��uS'ݤwz�im�L�n?10<�)����%��B�qޯ�ů`�ja�>*Cƶ�*b�L�S���n�X�L�L"gV�c��EEoC�R� �����IQK�>�pc0W��V��s�R��[��lۃ�5�)
��Zt�>W��m�1S��E�VM��F̾y�^�x���X�� �G �(�eI=��H�����y�y�!���{�������&���e�<�7OW�PROd�n�G5�;�����f/�ykB�L�,g�&R��w�?5&e�r�둹�,���*خh[��e��U�%��X���26�C��-��_�_P���� �/�9�k���cl����9c@��E�9�� *�蹄yQ/.9E.Β��kb�!�G^���V�L��иX8#�'�\��Аnh-|32�,���8ZX�����y�fʴ���/�6�Na:���2F`q����
�����<�8ѳ�G��3�/E�^d� �E�]ꋙ��A���J�����3�ɴ�u͝C�1,C0����s1���?��#F�Y@c\�M���ݛp����(�_��(�x�gXAY��sy���d����/y幮���\}���*S��S�3m��Cs+c�*
��*3���O:�V�T6-��i�}]E��(vξ5Pl����S��Dn�V����j2.q�0oQk*hK�U��C�������l��x:��h�Ǖ�6��(�7��}w�P����p����q�x�9�2�$I8��T�ߘ?��q֭��rwu��?�x��x\�B�{\�"ARhPY1�`fʔi1���&�S�ns��38~�����>#:�c6�:C��:�1�`%E�ڀ�����G ����/+9��Ӝc�����M�)�?�r:�Tx��:�8����x���3T�}�{C2�r@�������:?Њ׋���y2�� �d��T{�+Lvȸ�<�)�z(˙6C�l�]E^" ރ�0nd� ���"����M�{���lb5�5��l�tn��yx,>�(�m�MYa��h��NF]��E�<f��u���<��=�C+�W��^�k�F��:��z��%SOX����ɴٖ���9Wa5bfNH�)&>�2��v��b�5��8�@>L6��s�&9\m�{g���S�t
��z����  v6���[z�[�|��8O��Pu��K+]�U�n�Q6���o]��ј�c�j�p�a*�<�)5�)��g]�L�5@�0D`��y��� u�S_�
/^� /e^��x<ETh�ͩ��k�nE+f������Ƽ����2�1
u:�b��h���u�쥜i��L!�<=C�>�s��gr���Pْl�����J���j蒗��~ͳ$_1iƍ���\�����i��]F�=`���hopc��6�-膕5�UHE}J�h8�'0��7ʷV)e�;۰���~��#Ɔ����{��USO��"��,����ym J�e�~�v���*�he�* �����*�Hd|Ҽ�����)�bbf�o�X~���$�CY�bdF `�+<��U�D���K]W�i�� ��l�<W���[��i���&�~ω�f��Y�Iv�q��}�r%/s��>+'� r9Q�,��}��}�F�8c`0�.0��(��]��Dΐ�T�=D%P�6>(9��6� �q�;G�2`���<�^+@sYZu,Dkܦ�q�LXδ���us�t�Oi����_9�����G�mH�����<�%������~���Bi����鳏�����+���xש5$rE����,E�aJ���k�ޘ�o���Af�}#��]!�^��kz�۵�)��,���⅟"�#ʫ�����ex�"�-�%���@�V�ϴޫKdI�3�&�[��F��T;�����}x��q��X�V`����x�M���:vW�n*�2��w''���k����Hz$��O��#WG�G�4���@4���_�i[����˽+�gM�Nm���m�.�gm�ɸ�1����2}����L!T�;	's�:ߤB������\c�o�������V�}�f���>����j;���l5�l奴-R{��
N�pCE��(o�Ͼh�_e���7V��/�j}�$F#��n[�齑i�*1�/M��o�r��L	�AbD0�HR�'��MfC��P���j38;?���7p~~Jk�`�g^�@� �r�x���]'TH��^����6��.��mC�`�<`٦�������_���K��&~�J�m����s��]�(rc�
F"ο��ǣK2� ����K2>�Q�'�@#��~ۂz�z��%�X��z�F4�9#F�[�癖���_,��3�gi#T(_-�d(��(˙��,�<�W\-%�A$�Ya��݋l���r���m��T��U���,���S9�8�^H�؃���Y�BφQ%���q.6[Π��簷�W)w��Ec�͛��]�Rt�f�E�־?��V�������t�(�W��������D�T�#�<�M`V}��ih��3J@���[؝�ѲjV~L�.�Mt�{G�8���wGpt��Z�/(�*�wxood���4�l�9�Ć��� �RZ��o���/`8p^�%���c��&4I��QĘ�'a� (����B E���K\l�#�r��j�8p1��[ ���d����Eٔns�[p��� b����0�����m�u�~I�CEv
[áO�e�qL�ڰ��~�ei�����8�G����I�l�3e�NX�t�<�^ʩw���S5�@�Lu��S^6�p��<�WЂ��}�S%�h뽙:::b������3x����Pu�C �)c�"�4�ܤt�_���b�����&�k3�S.!��6�ؑ,٨,���a���ۦ���7 �z؄��
�Z:�	t�MX�A -Лz3���)ݮfZ������~߻J����l�E�F/��d
�^�"��� �K^�I��Ģ��z_bni2^U}��f�V���\�z���]�����"�͛hf-��@yͧ9r��3_��iI'�%���x�5�g>߼ڵ���60,y=��u3�F$�[Wc��`���﹔2S4Ƙz����J�ʍ��]+4&S�L�>@��r��/��'d�"���h(7��G26����<�,J�1.}�
A� �M��w���~XQzB�[I�+
�{{��Bܣ����ul����MO�����R����;,��X���F���?:�{cP���BE�h5�s�*}��1���V����zF�K���)\ �D��#�8���a�����rpj�	R@�Ci/./���װ���]�F6T���bK<����M_t��p}oh�Б�w�9'���/r:�	j|���Z��!�3z�M@���q@Y��9�	|����#�l�������3�y'Vs�v`�����%=�D�y�Mdo�֥�*�羀q�?'�)d�H�⧱��X$�����?��o͛�:?���c �nE���V@�Ϯ	��Q^�sDO |�^��N'Zs	H� ���.�>���hFy�Bu|Q}|J�wnl >$��)r����ӕe��HXδr��[��2I%�칼i��] xBJ�\�8oC��9U����c�S��J��������4_~�%��U�Vj"�B7�C��F�~�@fXa�PW [QK�:Gj��S@mVA�c���v��Xp/!z1v�����CQ�W�� ��Bh��U�!cO=�?s��n�
O�Lڌ` >�������^
j2
h�N{*E �Z�e�#'''�����C%����u*�b��?�^3�'@CA���{G^��}�����F��^��f�v�[�m�]xe��<�S���$��r��HA?71߶��A���.�~cB�~>�6�ɝ��5*�dL����C�[�"��q�G��6�y[Nh�2�.`�����S���	���c��ʦ=
�0��n�i�އ�'��鮓ދ��R�Є��c	Χ^��z^?C�A���~p~*L��h��t�#B����$IȄtc�ȒtW�#S��Q�3m��+����Bd����iޢ�����k�)u��ӹ�.Ϲ\fe�O,2���� &��y�X��PT$V8�Cc��j���+��������,GmY��xӨ�юڽ괄B�ޡߔx�-�~����9]�Ӆ"�@��}�Җ��P��l��Z�U)��I� ��y���Mۢ�9Mc�څ��~��%�mχ�( .S	�w���
��2l�n�@�7�	�\�T�4�u�̺�j�� ��m���m&>�,:���,2X������i3$�l��rI��3/K7�g�F���P�*�XƱ?s�u܁��y�\�����"b6��<�횀��6��z�^X� y��´S��!��3��h�Q�!�)�,
�^2L�N�Q8ޒR�S�ߧ{˻<���ڛ"�w53e�HRe��>)˙6B�} �2��\΢�j�XOe���STȢ��$E��i��ʟ�s�Ǔ1�loC��W�Q��s��	��`�i8��Q����}��$�z����m�eb��.�|�i��_�*�݂��i5/P�J��K�l��/��`�) E�k~��n�{�s�Eٌ���K�߿���(`Y�T����^��.�߁䜴�Z.S��'�.^��[��s��5Bo����fЩG�d�&��HB�Ò�2z" ds/'wݞ�u�%B�<..<�>�Q��خ׍�����vdX6s�t]�r�5���'�������p�i�e$�@aLoQ`�N)�q�3� ����z���ȣyƅ���e>��V��y�q.� �ީu��EL���6�M����U��¹7�?2�?��r��'���T��Q �D-0�,��H�#���
E='iQ�o1c����pz���)v�xS�s����TS�|�i��9�h��HZ��:����/	�d�]�(�����+VRlѮ2�oy{=��t�����Z�s[z`r���/��
�O�+�m�c`4����B�k �7m���v����_3]/�R��p^� �<�!�G�[/D?LB��g�N�0�\D�p_�z�;*�G���Z��]��d
9��� �dm���S�_��;���gS���(W2���6`��|a'3����$�5,��C��7�0�wp=y��a-do�s�ꬍd��QԞ#~��9}���S�3m�B�һ�dΥ�)%��;Wç�����kD���t��Pә7����%�k�T4D���(��\�����ҁ�B���^���/$�z����-�ޗD��x5�]�oXZt���p�,E��Mjع����J�������HT�S��U*���Rc�z�����2-R���y8�咞k�݁��&�+�xV�6��,:��,Nk�e�቙�\+� '�I	�ed��˚>?>�=���&��~|턹Rmy��6x���O�Ok�#�*@���<��B�������q�����O�,'9�9�C}u^g}��T[7�$e����膢G�Ƀn`�a�ϊ�_���C�����w���-��%)���"�~\��-��������3��~����<��B��g1��Oۖ)�j���L�N�%9�<x�$�i�p�Bd!/Vw����w��h�l�B\Y��{����l鼤*O]�u]���tF��%o{{��J�	�N�����W���������M�v¹�4�o�չ8qha�i�r������}�Y㐆Ǌ�1����-.Uӷ�{
�O�z�Ae�*�,�*�M9�0�uQ�eI@Q��@�"�(`����^���~�4���n�+��Vo[|�f`��Y�9@�m�5��r�K>�H��ז��9F��H�-%`]$�w�k^�|p��|@`��$b�^&}� K��,�g�X����a^-�<^pI����e�q��k(}#y6��f	��p��� ٦�Y���ѕ�vQ���v�^��Z�
Tk���y���# �"�9G�
!^R����󈭮c���)�>��of� ���#V�u<��6gH��^��ű?��1(o�����Z$K�קϰ�QQO�W��V�`0$pAg�+ŵGEd�[���L�@5�9nl9��)��������q״��uX�������͒���Y(І����y������Y����s��9ba \l�c�p��LY��J�Sb�yg�Xz%��3Ğ��&�^�	�*���O���o&���>:�d/����N��D �抡y��0�<���t�ۅ
O��@�~Pd���M4=�yb��WV����y��Rdk�aߚ�$��R����7�o���p�풟�}(��{����n����֒����e�y*�D�[�����Gx�e�ʘ�J:e}Y�D8��<·A���@�&��W��d82�ϙ�[������G��뽷��v�eI"��;�.U�:�o`0B��yJix�^k�ugX5:����\N� 9�Q��A�dyP�~�@��p9SU˥�����`р^�j������D�1����]?a�?�Eֳj�����q���-�uL�{w��(�tj�w�#�7D��<��6H��]hX��{��?+����.Zz׺6���nܰ�G����X��>�p�1�~��[ܼ�V���ߜk���\��$�o�3U��q]�]d�(���h�u����"kHc�H*C��q��x9�����;�[8����DCk=�uD�c�wwwa��������[���ɢ-ka�;OX�tM��Ϋb� �r��;,�f�U��ԕ���Ly����w���Jٳ8��t)*&�лpZ	�T,g<�(�E���)<w���zE9�JSק1�=���GX-�P�<tS`Y@X �Y@�Dp��r���O��Cc�E��+E��A�Ϋѧ�8���<���5p�����x2�%�TY�Zu��
��ȮD) iT����1�^˪�~�u�F�[�����eP�C��zO����^��L��
��2�c(��)�s��ǐS~�[�N_�w6���mX��<M�����yg�?��/,3mX���{o��V��h��F�ʐyOo>h}/�F���,�c	[	����y��o�����<g.���(�4�1X��_���q� ��2��s�oZ;��M�����2���f�"4�~�໙3&n�ԭ�>�̭� ��
y<�7 �]�X��_89�&�')��n�m�����J�1f�����dH7��%�߹�n_�x�|�|k\~�e�M�X{���L����x�JWG�����E���M�'�y\z�^�g �IG5jMC^�x�@�>�B������͘��+��Z����v�J��
gg�py9�ѳ��gggprrB����!�����lmo�)d�)S�,g��J�w,�twz�nb�U�<���E�|���F�����E���hK���cj��!�cy1��AZ��@g�A�����*Bt��|����E��|�|�Ʃ�^�guߵaƺy�wGH���'�W4�N�P�X�m�o��eW�����F�/��?u8"mD������KyѮN�.��<埛�s}&�-[F�2�)<� x5�3U�E�׳ޏ{}/�C���DN@���L����G`,�dA%�~K���7r��(������41M�����S�YX��C�q`e����#���7�����<�f`"�5 �-����GI�y�
.&#���kz���@r\+�{�x��~0M�ޝ��N���c��aū��[2Vxmg@�ۍ�z��L�½���=�)�h.�������~�ɍ�h��I���$�;�0	@��qʴ�ԟ_�0��D ��=b-{����Q:�f���yoh���J_���.ԴVن��*d��5�aϛi�*C�Eh����~�� N�p@�ol�F �R�໤����	�VX�M࡙n/I��%� �!zl��9y��N�ݻw����G�`��1�/�0�����?��,g�v��BWo8X|�QBQ^�3]7YΑ� ��&T!����m,�qh�e�W��N Y9��ݮ� �w���02��^y���H�~;�-��:��o�萛��տ�m��u�M�M�k��Ň�7�N���t��<Mm0
�n�ԍ(u�2����u�����g_5�zP88>� ��)Wj9s^W�[b�q�A~;��3vRL�{����NR[�Q���4��ɪ�� ��:E��$݊�S4����E�b�0&�繛��Q���6����Af���֦v0\���/>׏����~&�:oYD����2���A�.Hi/	�bHp��C2X И�~4Ĳ���i�z��0�	�N'����h���Yi�l��ti�f�sW��sX����[[C�+��s�A�=�v�wh���l� ���><~��?/_����^�=������`o�[P��1�)��E�������p��ol'ELU��$xLcdpt~�K��Ӎ+T�Ϻ�l�#�u�+}�4I�!�����7���a������;@quG�P�p`����������$b�x�r���������&�����^\�x�D[��~lw���Vр�R=�F#x��5�p^ܻw�{{K<�rn�:��z)˙6B$���,{��N�yP�	�0�|jj�*B�1n�E!߸p 	ۗ܆e���(!~��u��;����A'	����v%O�Xd`�T������I�	�u *Ҽ��(�Q��~���R��n�ndt;�w/9̓��M7������ ��[M��vi66�n�X�ݦ�]#����n�pm0��"�ᛕ�Ъ.�Nl��J� �S�P�q�z�8g*~ݫYX��L \��(($�����xiR \���HGt{�;j�o��|cjR��@����z�����5m5ꀫ͹�϶�{��O*�~�-1ŀ�B�	U�K�n7/t��J�ַ��[��B��;�;T$�������kY��4D#t�/b�� �� &b�:c^���A�]�{0C��ޢ�X�j8Pb�QG��s�s�R|n�=���S��><|���z��|�ׯ��a1~xy��� �8%`.��g�����Qu���x��Qɘ2�^!�y���Ny�K��@�ف�Pic�y��m�ܔ�9�f=k��Bf��mk�
���cI�c!���*[P�d:�"�u��:�/�HS[�b�L懖���t�I�%+P���1���ܵ�X�f�V�H��k�-�!�a���8��u����"��N���2�o��r��%�NB�2e�Q�M,�6��� ���ܢ����jAEϓR���:�-wse��+u<�c:�;��N�9�4>ȽS�k@uK[�](Q�Ms��1Z����CY�Ԟ��6?!9� �i�=�R�����~����~�(\� lH"`�ya豴���R�%�H;����}�@�4�'��P� �:E�b�=�k�w�4�� �(��GN���Ԧ[���+�"t)��e".ʾiC�VN���z�6z��?������8�x�sm) �u��1�H�{�6�^22Tv�ݦX!$x�|��?��E`to��+�z�|R�&[�뎊ޛϟ�U��G�a�ر�������X	�!c�ݿ< �y`�sw��ϩ+���U)}�N�� ����������"�F�/\*�//ilN(E���[���۷�������?���;w�	З�p~~^}艞���):�L���E���
I��8ؼiK�$��8�m�<�q-h �ו
Cx�6�ѩ7~�uH�# ����@p|� Q=�K[7503��Z�fӳտ���/��ge���9�m�rӆE�L �B�M�/n�St��\�x�/���L�*�S祟����J/�C��=�u'�LM����֚���!$	�6�Lz��̔�����h�� 2{�%���\�R�s��K߻Zb�X�w(5P+JU�4%`���!W��y�t�G���D�| ��I�^� ;0*j������{�H�ª�unc�j�9'u�w��,���9�F����)�_z!9��MH5fs|�:	�{��0�l�J�+��ei\[���6*��?$���S�ǣ����;��K���)�c6�cH ��bj��IOU�u�q��
�Q|�|�MW����uȶ���>����M�@xV�U�th�UoܰTs�Lc��l:���_ �I��Y9\.�0`�������NSN�V��%haZy�dnQX>�~��r��$h����L �Լ\y�o��_S5��=���+��}Ji�����ՍkK�g����3x��	<|�ȥ��(+E��3=���1���#�0�LuNo ��?�(������iα�@g���#����}x��)����;�z���#Ќ�����w�m���lcq�,Uϵ�]�*s�xF������Q�u}�]T��!ƅ���N�悀��[rSQ�m4n���(b]�p�t*A��f�����$�3��`"��m�a2u z���>#m*��ƺ���S����ʶW?��L��Ds���y�0G��~��@����H��$s.p�Lw�2���.��=(R�=���$����k�d}���2�DBE�VJz�X�T�	�*/��kdQ����\	��k	
��<��/Ӊw�X��p�*2�=0��PHN���ئ�
?�'�|'> �xۀ���y�"i�$@��L#?�����/#��K-#��V�ܨ���{}�G{�t�Nh9�x�i3�q��Y��Nm�����mYFPaEí `y<�+��0�X����z/3����\�L)ͻ����I8T�u^#oj��^���Jz{�IQ��XW�=6Bm��&й�81F�֣�s�ٯ���Fٮ�.w�yT���3
�h�
nO+i/�����mV�q�&�7L�>pr������T�x~�m�^A��¦)�ĳ�j�y�!�*y�ћA[�������Gp���6��㏞=�½{�\�ܢ��`?9��?���j�"@2N��ނ��e�ey�����=8ؿGmA�g�P>;?���xw��哓��S�==���s:�Rl�����.�u2�0���=��'zx��m-T��=���}bt��:׊��<��S�q:w0L4/K*�ͅA�h�łk������\��d��tI����ܰaMp�{!Ƒ��I�5'�8'���y��ɱR��;�(���e`�%�������LI��8���c���P���չ)�v��y,#�a^�;[��v�W��#Ë&*%�� F�c��ߠ�p�y:x%�z��zAخQj��Blڇk�������%	!O�)�L��6�淼)E�����8˟����r���0��<'� m�z�p����D�ϰo����X��ʎ���T������I�4ܢ�+��(g8FTF��~�$}�F{c�:�����S[��KG,� 2��6��_-(�ƃ��j��Y�"�ͫ�{��jpY���=K��3��!s�Fǉ`��.�n�:��u��rb�C���n[��;`�x	�7[w�����h��"g`a8��ǘ��zn.�W�cB�	����4�s�Ǵ�:�N�����w�=�&�xgwz�{�w� <|H2�z*��'���Gp��C"�G3"E��vN?x�j�R�\"�P�vv���ѣG�12^^\��7o��/�ůϩ���89=�T���� �:���!�-!/��+�n
��;&�6�(�"�FFgj�K���r\V��fˡ3^s4Ϗ���u4��s5U(�)M �ItQ���e6��9w&�EQ*�.c�#oo�$��1d+X�z��a:h�;88��׮oW�LX� (LvF]N���\.)��%�[W%�����[R���X�A
�f`�i��,�&�t�zH�60vy�P�鑃W��v�
�Vp#�q�|X7͛;֡�:l����Ѣ�-�Gz� ���<.�� �M�U��U��u�>�J�N�I?7Q+��[7����w�P�m4�
c힑�Jl�ߊD�5��v�m��y\;����z��u
ejX�E�:��\
e�(�kP /ga<��5�:�l�u2�m�Lu�L�6���D&(�b��×���#�(���-�HG� D Z��:y��S5�Kk-K���ȏ���A@G�iC��m�Vؤx��MK�w�t�����#�fJ�>-F�cm$�#��jZ��`�j2���<iG�sw{�R�# �2����_|���o\_r񾃃J9��x�����dYB�+y��Z1��G}_������qqb��������\��a����a��=����pt|������{5��2��N>�6�.�x�9���w��u��z�]��_�~�~�^����d]��T�lhe�Qa�wٯGf�@V���)�ij��F�sk$�L��x����0�V��l<�㻺�8�N�Nᗟ���	�������56��(�f� 2�[a�LOq~~F"�@�y��@(O�`�r
^��%!�eKn��C�����!ԔdTNE�̙?^�f�4���౬o�D�i2ϕ��t����.VA
	n�;t{�
hz�(��-ϠX�� ^��s�Q�)�0� |��c�Vk3�� یi����٣X��kml��M���y<޸�W�~?M��5Q�>I���Dg5�<(����(*�;�b[0�lxͯ0�{��n��m�NXC�y������m�{M��`��'�g|�+�
V�y�m�����v��C�*��C��`;�����- s�ٞ7��(����ث�U:�V�̈́d̽O��o��Ms�=�Q)���M k�U��/t�>��=]��K�3� =|�J���<����U�����W_·��۰��*"�!�MwZ��L�1�u��c����z��l�3�h��a~�3`.���!������bt	�'�X~��5<���qVBqyQ�q�$D�%zT�.X��2T�dmD�&���.��`������a,�X+%����?�\(\~��y��e˲=�r��{'*�����m|d�2���yS��&S��Hd���Y�M`�~��)c�����!-��/�)����Ы�r�y>l���&f*a�Ff�y�޽{�޾���be����b=�hH�-��1 �r�9M��Jn���<�'��<���D!�q��z��9�3��`ɼ�� �p-�ïE`UcD'���\�a齱���VDw����GE�zN)*�r$@��)/C��Sk��rAz�N&S
7�b9�����kY����T@�pNEW� G�1V�4�c^�s6꼡5���%���,�{
���9��M��mma�-J������a�+\v���l
�me����a]_y�Q��Ҹ���5�� �pۻ5�p��	���j�Lw���ܣ<��z��M�@��[z��&<^�V�d6�%抴�׾gh��	|�B�/�)�a���a�\�
W ��ʥ棛ƹ���20�k0�\�1��M�����CJy���}2���_~�E���J�����[f��](>9�L���Mkd9󾑵u)��2P����l�������3��sp�b��eL�1s)2Ɠy�yc��j\J�� �[��f޴_u��u���zX4�����dsYK�SY>d%e9�m���f�>�t�x��F�D��eF�@G���3ʠ������C��GQ�'��P�!��^/=7}�Y��C�$�>��DE�E-��`=�����O����)�w�|5,O�.��m%���hr�X�X-�ͼ Q<��H	�T�b����չ��F�N�i��>� L�p�:J�)��̜������N�P�A�u>՜6�sY�5J*1��"�JP
HC}���M�TJ��$)�b��z��q
\��T��窶�z\Q���������-���\�[(���� V)S>ca�}~y�g�!�8#O��;({	���G�W��>������G�����hU��҆B�^<K�=�j@��'���S)�	T�>벾�G�N����%3g{�'�p��g3pz�]޾񂻿RK.
����)�@�7��*0F
[��w2W(ƥ���m�Fߦ��M�7����Y�4���wP; ����d[�_'�o�(��ic}&��% V [�@��t6���%��{��x��$�A}�+��s�@��״^�.�z����n��{�&�Ѵ	8L�h���Ab�v��Ƃ���V�0�N�Bc���ô�����o~�}�)����(/`��-*���<����&���#���趫�_����}�����6����m�w��?��ׯx��q�۷ǕL3��.D�?�n��֦)�ܗ���r�.Ջܕ�o� ͽ���(:��^�x/|:ǰ��6�_�=_s��0��C~o�rt#�i�J����H&���� �2��(�\n:��T��<8;;��ӻ�B^dZ�ߒ� ӝ�,�U�!.��K?`u��s���X�$(�����^ϙ>D�q*3����d�J������XQ,S κ�ݥ���@E,�bf�p��+�)����D R׳h��ۖh�,�1�}"�MaU_���q��;�ٚ9�⌇�Y�t
#8 ��u�U?OƗ�}4�"��(�{}ϛH�����1��(�
3��%�xL��N�q�y(=��U���G���Y�wv���τڳ����v<�d`y꼙��O%W=>-#p��L�0�B{1���ޣq��q��Ŕ�� o��[�s���3�z��i�J�5;���P���z}�����{�H�M���K���:���ie�L���D�׺;�a����ޞ�J��0R�[�$Sʉ���Yj� 0����T�'�,��9�?����0�
�.a�c�{�0d�[�8��$�l[t&Y�����~M<�Jp5Nջ�[�?r���Y��#�y�����ф���0W�)Wn4i��gb�A>��yi�H,�5.xe֮�@�Ծaq1���l]҈�����ߥ���@��V�އ�� �V����:�9�0ƴX|#<X~����w��o~�5ݐ�?y�s*�Ԙ�>7�/���TzH���ƺ�'~����^}�?>|@2�)8�Q�����Gr��R3X��^�ӑO�m����k���5��$���[Z��"~��������6�7#`Y�M�L��,���4���3�u�ѵ(�{$wbD���ǾEނ)$�4����
!S��R��A&7g�Znm�}4�������7GN�9��c�_ZN���]�,�!ҋy���߽;!�5���LF��U�l�o���lT��i��d�y$ 18�N�Oɥ��W:��V
]�RC�Yע)z��gQ��mw7�1�ܝ�Y��+�4`���OpwL�dY���  �`k<x@���U�B���i�P�HA´=�wT���D�霼�1�"
��m�,�ܚ�ጟ�+�H
D�O���F� a����-����g�{X�܃�}R�zJ�S!��xT��kI�e��Rf�h���	O��]�
1�E���a��~�\��1�a��a�L0ȑ�'��˻��/�]�N��S$bG+�{����WO�d��mL�BAN]˨u|1���Na<�gw�w�#�4�����m�m�O,E�V��B|\�����{��ƫN�W�O>-�::�P�p�o�	��yߕ�4��*'���,�^���ܒ�Lz=^[J�q˲/��)�lď۔��J�މ�$qRF���(�J��G����&�~OT�-�O�٨��iޱ1`�+�(� ߓ�O���?������alo���>y-c��%ԑM�R��5ԥ����!|����G�(��/����.�kP&9yw�1����Fl��W�d�5 �1uv��E�_�_�����h9c��D�Ik!ϩsK�>)��C�-�sr$:�_L����oyN緆���cNLs�"�X~,\?i��ɫ��`@��{v0ʴ	��A�l�9RJ�jN`�.1bA?ԛ�^.���Q�o=�Э������[8==�\��Y�nZ��Q��H�KA��ʔ�摀ĥ�:����"Ȉ�i���$�����eZ�ܵ=V����Yp�>�ܐ�<f��l���-�`�SD�K� �u�!�9�Ш��V��=���y$x;+�b0%��9%)'�dL�PI���T�q�hvwv)�ћ#��� 򣽽=:���3s�-��WrѠR�*EwT)#�>E���E�CO��	��T�~�I+�d�������ɔ
���4�s�<�'R!��=* �v��_���ȩ�H�_8@҅��ކ���s��Kc�Z�]d���+��)� ����+g�P�cy2��sߧ�� y�Ai���Wu�z�(�t��|jV��+�KER`Y@ȣ)���˪�ǈ��B� |�Īi�������ؖ���/>5����>G��6�z��vt-�T���Ze@|�<L�y����n�^�2�?G7T{BS�˸��;�1�հ��M0hV�G�qcS@��w�����gl�br��V���Z6O����-�a4I�)��1��0�d/��bOeIu�y�qM�u��o�����
���Hq�cp 9�u��{��w�e�������]�pǈ*���~�w�������1<�x���3� G]MO	`���Ӊ��Ҟ̾����W�J�#� a,�]&��F��`,�H#I���� �1���n�,�EN���c?�h<����
�q� ~S���/$����&�����&����;�}0�{�K#S�L�õ 03�d�����[MdH0��!����+���C�`�s��P�H�^�3��h�[Eλt��Ң�3V�-���5ƹ�X��Iѹ��+���(nW�X��9Ί��0�4�, `���J-��5Zˆ���.V�b(��7���[x��U���"�BE	s)޿� Tt���y�ys�?������޳�Ͼ �
������a���:��^�|o���Y%Q�[�ϊ�E0��������������+z2�Q��:���g�U�:�g#@+���Q����#K�ht���h���X��#�[:pZ�9��v�6
�	��z�{:�o�GÜ���ǟ�A��S�¥m�Y��Db睊�#��v8��{=�E��.Q��ү��_K{�� ˤ3X��:9C;T�1��Zļ�$}P 1\a%h�]F�}�jlØ7~v�<+c��Z� WX��ǉ�u:Q֣��i3�G�{�a\0��ݧ�rn�>�ǯ��Aa�Մ�Q����ਕ��b�gɡ����Pjx6����P��og�g��r֭���l�N�t�Zc��6�C���10�*�B���[4�\��6Fݿ>��c���G���O�`��{VI+�P�E�TGd^ǲ���mn��tj�Z/�{���v>���J&zL����+���4}��s���K�sP�ڪ�o�l+cvs�P�)gt�y�Juc-��n�S�h�.ݘD���~|YI��9�0�B�)E�a�1�mk8��XO�G����s.(e��YA 2:!/~2�\�ո�Q���K�q���v{G���d�tur�-g���k��q}y�"�H�<!�m\�픁�;@,U]L��/0'�d<)X�:i�� ��C�<Ty����C`�B}(x<��"��:(
�U�	pf(B 3V�U�q�8L��I�/����j~rפ����2bPA���#z�?�w�ć,[��݃?���T��L��!�m���Q>�'�ҴS7M��䭃i*��;����8���g�ǟ|B�*	��6�o)U�	��P�$�^�G(V
.~}�3�����~���פ� !����?�O?�D�D�{8�b���裏\n����F�-Pё��ɔ>�ވ����^����&k}AG$*�6�Ə�Z�4���S��:�F�Kd\���W�1G#��䢏���kt㫶�[{*�g~�@����q1�q�T͈ֆ���5�MJP��c��I�`@!�Ƅ����s;Sb��	X��-����'2�mX��y�QR�2m��؁l�:d��]����ϱQ��W��U�.ʥ\}�Ӓ�֐x��,GG
���󛌺�;n5�l��ZK_��NO�h�D����!bj��:���6���~��^l�s�w��8�6���j�|��|��G�Z�?zϞ=��S$���Xr��XS���t^����B�F6<�o� n�᫩m[���m9w0��`0#����A%#݇��������f=V�1���W>�+}R ��."/�Q�U�����[����ƎLr=Iu:�&F'.#H��."��za��}���т��jz�.��Ȫ��:х�-}�L����y������8�i1> �����X��&�;�����
ש+��2�f�X���O2�|{���/����0�8�XNT
��[ң�{Y�Pټb[k��p�<C��;�䟝��p��
w�v
Ct�z_r���8�ó��E�'��ǌ�#F�C_\|�����Rh'V��w�j�U
'��;�������<I�+=vD�����������lU
��C2�a�
��8�V�'��1�]�=T`��1yJ㳞���������Ͽ�Ͽ�D���/�;z�Pn17^Vm��I�,O),�����L��(+2F���/~عZ�n�������SP=�`�5	�r`�(���<R����Bh��8p�����J()���Ltf��L������대�y+eKؠ��d.3�f B���B�D|����Q
��������G@� D頻A� �i��L�l<��<�	8�}�0���r�X�����n0���z:��:��H�f�����<��b.TT�[�n=q��K8>:��~N�J�Lu{ջ�����N�7Wi 'r���* �y��yM|����mx��1|�՗���~K (�� 7 l�W�U��M��� ��������
L��ZH}İ
  ��15�MG��粋��RR,Z��(Op��6<>�d�]ʹ���_�y3���{ձEc�x�§�(�X��"��Y; ��VzP0:�~\D,�-�ػq9��@���� eQ��Tci��ʃ}�y��8s���+�^��-��wc�}$�a�"�`c,�@��ϔ���q�-㊷:�e4�NON��?�_\�q~���+e�<e`��Q��haVMd�!h�ynƣK��*ڢp�U([�2�t2�_��y�+ ҫSvC�4�i�S�X��c_M���W�ԄeT��=�먶ϰr{���W����J���)4����z���x���0_Wߑ7a��ӧO��/��/>�>��s��O+���+�RK�?$E ��Q�<#/�p�~u�y������{W#SO(���8~w/~����<x��bt�g���LaZ�'�V���7ګ��z.�r�>�Erp ���	~��o)>z ���s�������R_�u�o���O��׿��}_Tφ�G�[[����[h|y��1��~`6���g���l�ؚmK۪'�J)�� ���S")G���e|gwuݐ�A8f�Ӝ��n�����F�S�|u7��}j����6�P�"/{}�x�@d�GE�8`��BC���Iy�Y�6��I;�>hjWܖp�<񞚤��8݆ ���uQ pCQ+�I`}N�țU���,����Bó�>�Q�]��9cN��X w��T�mww����sO�W��{�H�8�h�y���� _�ƻ�~�ƅ�5�y8�/��&J�aT�q�a�"zvw��ѓ�p�����)��p0�d����ة��ŋV�3Ƃ��q`���[;"n(�p��lt*�t�{�<Q�w�X�1,�0�`��]+�������MϠ��Q;��z����%����_�wI��9Wr��o���;����J&����%�W(�̂2�-5��{��Kl0l��yTJ�PqcN��k���Iq_�-�T㻿=�6E�={��"ذ�2���(K"�<���K����B�V�1P]p�rN{6�*I;�H��2�]ˌ���R$�ԕK�X�^I�Q��P��&tFs��%-F˵"��Ϝie`���Bo@��{wrR	�S�a]�"K¾���@��G�2!�1��N��iF�P��� �)m�N0-+�1;�mNِ{\u~����E��a�GJ�����8G��J���q� �E���-{��R�<��W���������������X����?������޽��o�$oQ
�!T2=$��R �d�m ٟ���E���!*Sz���-�}̡�F���ļن����8�'d�=��ہ�����a����������|����&��F��J�q
?������������M荍�y5��c�w�(�T���1�Z׊����V�$A:X@(eÆ�T)�	��fRy7y;��8�z���÷���?����0w�/��B�S���T��y��UL�y�ٶ�1|� }D��Y1 I/�����*_;��	`R�\�Q���x{`�iM�"�� q��^y2�Lh{Ckk�(�M|5
����$���-����E�w�}!��{n������7�Z4���`�v0��N`����瓰u��u;��ydG/C7P��2����R�15�M��/�MޝF��i�BO4Tk*��dx���K��O>��<yL�߳�>"9��/��H%�F*z�̅�N���aE�����_\����xA[bk���p�]./F��G�68�c�
�R-���~.B
�8ńI��Y���J�K�(z)��7� 0��aDFP��O��˸.s�|�-�)l���?a������v96GM��|�^�u;�$9ei�i�N�!�-�m�W���2:,<|���#�0�z��̺S���4fl���2s���g�����l���]Q�Y���Db{� R?f��F�WH�;��W�{�����I(ϑ�HX��ċ:� �����zZ}X��{��U�����L�6M���)�	A���%�7@0�&(�VB%����Aeb<��I��Ћ�'z&�`�4Hf��\R�5���hS?��ȉi$��Z� �� �T�E��R,ހ��l}��)�O�>�O>����k�Q��z��!�Ō@iT�^�!=&���[����������4�9�Ơ���`ovP�n7�w2�V�1��yx�^�R(1*Lؽ�Rv�Aa�g:���B���gx��1<|pH�.��O?�ϟ?'/ �����w�?�c>��A��7KX�Ao�Ϫ�q(r1�-Vb�]z���Gh�*PG�g��-�>��7�'T �4AL�@���#%߹q����b�J6>7�ۗ�^�Ͽ�L���l䎒�1��'D]T�ʶn���{�`�޶�:��2)�#e���Bz�e!�B[{��-���؈w8+��
,Zn��E퀢a��d3��� ���a�|�~��`z���N�j�?RÅ��ُ�� �uU6{E��e)� ߘx;GӈGeK{�G���؎��O�\N;8����F���Tk�}�1�W�`�k���A��ԅܴ&���q<���׿���J�F�/>����[���H�*�h�,TM� {��L�q��ֱ
ᯥ����`p��9��#�7��`������H5����D`�y�"ȋ�����م�Jq���})R	��,��[���ۇ�B�)KMu��(�̂�����b[	��G%=/�x�VȝQ~�;����^���`�r5��秤Ϣ���;�у�`9�zuzB�]QdL]����S_��}���<�\���t�O(�-�\��;D��`J2��xl��A7���*S��t���t���S�}�s,#��M�Uwʑ$S�o1q(�<�qƂ}�Wn��ⅰP��:=��A�A�L�6M!��V",�5x���3P���W3��c �?:9j����V�8�6o��D�Us2�z��=6Uޣ����U�Nt�!�Οܣ.C�I�����KqN���������������K�1<sK*t���!��bJl�w��G�agg�@�9�����;ג�4�4���T�sl�r�C &y�Tς�.�����`�C�߽�{�k��!�Ȋg�A&�{�"�T��_V�7��7$���xD�-/�>��� ���������������l�x�戊b�&*00<�(h�`�����`V)S[[�!]K-������d�H� �JS
B�;א�HX�D|D��ņ	�#������ޯ���%��Ɛ	E��OHqH���sȭ���
&�ݦx��D.��).�K7�!u.�z����^8x�������g�X��%ց�=q�S�N@H)���� }ӵ�mԡ+�����A,�6.n'Gk/h�-��K1��-���� ���G�Q3�ijB�����Eʆ���#>i�P��͵��n�d`�B��S�(\/dƵ��q������$PS�����a���z��,�x���T赌�毾��Z'�H��]�M(�LSt��1$ۍ>&J�y|L]��;0�@I1Tpj���\*�(�麐��d>Loe�3�a\�
�K�ؒ����S����*H���p��!fe=��e��=Ȑ���BY��F'�'�~J��&�������q��,����#JW��*�f���S�6Z��'�����h�R:�_��~���2:6L\�3�;?;�sKu.��"�3�G�Zo/]�d��A��H���u��jn�<�UXpkbX^��y�Xd�rkʴ�2-Ek�\�<)~�r*����y$��\4�8�Z&��}��Q�o1� ��/NH9ǅ�慄MѼ��R$�l�i����X25PSN�R)�D�}SN`5=)����$\�[
�����FJ�9��d�����T����8%Dь��w��QT
G������!�j"������J�}���=�O?��B]�[�E
���5����p�Y��{�@J���]��ַ�;��`ǥ"TJZ�^�x#�����P@T�50������6��s�H�,����n�x|��#8��$��蝍����~��Gx��%�%��6�F����z���[;����k8}�
&zp���2@��z?�,��eߥ�)�g�����d`y:�D^\��vWRa.�9���)z�SJ )h&�0�L�=��¼Q@B����ȨX
y#�
����&^��	s<��������I1��{P����:9�{��{	�!}�SH�yg��]#�/�PB���� �H�c���,\��~�$�rC_6�2txoE��N�����U��1�q�T^��t��P�C���uAIN�T�o䩄����zb�US�H�A��4��߫w��k?~L�b��}�ń՜�G(���]ƒ#:�ć{ 1�Ze�o���ޅ��\��W__~E�g=�X��%}�e涄�����ш<��-�Z��/.��"���lL2��l��45+����(��3���t���X8���nC��Ep�c'øZт���c]L��w����!�fCB���qm�����h<�R?}�����W2v��o����j��\�3�C��z����Yw��_x���jB�e�]J�vov����^��~Fy��S����'\gІ(/��Q��P��}؏(o�F�Ȫ��ݓz"���!�#�M��L�>D���DLg ��hh�Z5���ћ9-�ݡ,�R*}��3�Ӊy�]�0\Y�	´�E������G��>ׇE��MB儼[\x�~�(�Ra�bB�XT�P��Lw�P*1!�^�x�A�|�����,�,͞��Tze�.-���ք�{(sx�<y��<y��xB��4��O�����g��<�A�+��uP���Z���)-����VJ��-���D����J��1����pՀ�A҃�Ϣ�2�v��\��Ћ=��x��!<z��Ǉ+Z����W_�?������������7��O����GJ{�`5�?���������g�~F�'�������Ϩ���!$�'��� �S�"S��	��HAv����W{/�7)�8F��a���*��>�ٱ�^�9�U� .x�ǣqa��g6
p��7P
����uE	�-\������l��נ�5l��k�U���@nt\ {�B�\�\��K�W�!�+���]@�`��\������i�����3'����@q��sf��A���U}��D
�����#���a�Dim �fEK��͢��kaȵ�����4x��D�	��I/� �����1�QM�5R�+�9[�1��.H��5�ٳ�.]B��~��i~f��Q!̈�6�ڍ���P�'�UD)����ˋK�wp�Vm�����ߒ�ي'l! �q� �N<-B���,�Ŗ�np��QsV}G��7GG��W �R[�8B��e*�6�#�Q��k�y���i:Og�C)�2�dp�� �����
�NB c����}j��Pd�dBQP�S�aD*���˧�)Ņ����k(�|�e�VC��Ͽ����z�����蘮��dYϏ���
�j^����cj��)��8��P��׏W�$waB�d��?�ŀ� ���u<���}b��{˽����<��}�hx|/2���1���P��fZ@iW9py�ћ#/w����N��m�2�6��򭠺��!�(��g)V^��jy�cIVT m3�	 W#�m�&�=�m�u��EcZ���{��2W�F� �
�(W�ŕ�_�Ja:$�p,ֆ`4I��Q9:~�h\:E=A�/R����3�鴮倌B �~ئ��>��w���R) %G�dTh��BR�+���>��g�o��O?����`�+z}p���	�e 8[�
6��НL��A��l&�$`���w��Ge���ƥ*�Wt0MƤ�b�*��B�믿���w��?�����T��1�g��������|
�|�1y2�Xz��%E��Ǘ���a �X�wJZ�9�B�bdy����t��ԻG`K��/5�$m����4siE][�+�i�!C��F�3���C
�ã��O�9�}�GC��E�(��O�w��a���O�+`d
.)O[��E��p2�ڍ�uS@���
�m����gW*͊?& 2Q�ej���|�+�Y�����ߔF&�X���sf.w:�lh2� 5�k��r�)0�#�S�a��8)(+��)�ً���(��]ۅ�O���d>��q�ɔiw�;�����Y_�S�Y� ��`�(�J�n�j Z���[��(���;�]2ɑ���М�� K��td֭�9�293�8)�3JJ+���Z�4�x-��ׯ^����<���41?�2�Հ�w�8΁_rj�4�7���sg�i�$�`���h���0��~�2�b��	mK�8��c�|1�Fa��i��^�RE�yF�p���˵
H�q�!������>��������>L�ƹ}/*Y�"�P��8::&���>���E�w�<�{���o/_��?���_���$������j��s�QW�~��܇G�����|�w����W�1ʘm�DŢ���eL2����j�3�
�By$�A`ad��ɓ�Hg
������z�ɰ�<���{�溮,Kl����D��<�))'ef��îꮊpD���?�?�mG�wUw;�a���2SʔR�H��88`���޽>k��=��EJ��dB �p�sϰ��k��H�Q����Q�d�_c@Îi1�����E/a�e��3[�(���ۡ����D���۬kz��}E��1��o���~43qOHjܮh�Dd��>�B�5������ϯ���f4�W�:io׾��*���vj���K���d���^�G��Z�"
�#@�;Y��s����WѺ��>k�F��EEk��%�(j�Q�%�a"�Ü��Z�mh�+��v�=5��f��h�F5��a��z/�8Vt�A
� FkOo�l�9�����l���kk˾�H%�켶�
IP!8~
��:��f6�� �]�诂YGM�T��M���B_����R�)�c�!��q�]��3�OSk� -Mm{��O��s��۶�i׼�hN"#ўh_��NBYъ�ade�gEFQU����Da�C��7[��+˫p�#�r��q�!���Ρ�*M���:"�Q
`��_��/�.C)�-f9E��[���
m�@UxΑ�j�����%�|�@b�D�nN��i���s瘪�` �l޽q�Pnǀ��3I�s�ӃI���%p���ׅ��8-�y���hD`�?{��%�}�a�Wt��R��G��p��8�]�6��n��XR��	����drnn08i�^KU�槞 �2 i�5�BA)��/�u_J��*W��d�+ ��f�EZ���H�~Oʿ�o"
r�[,]c��� ��I /-u���Q�+v�Gʄ.����xJm�V�{[8����_תAY53�2bnw�� ��֠�{����>Ũh��u�mʨ��3s4�z���B�3;:�u�ot�1[^�)j$��Q��!�׎�
;`��_�_��߾,����a�-rg��ٴ��.��f�������U�OO���}TY��4f z�n��}cs]�-67X4w~nN���U�w�����1:6F�;�=_��*��2V�в�}�����h�y�gmR��'��q~��#����G{ h���A>�^W��
m�����"��>�$�~d�P&<�[�o��ǎc�Aw�RM\�>&p[������cb�I��k~���F`�v�r���P����yQK"���ĈO�bA��u��趫���mj[+��V�kK�/&.��� ��i�ߏ֙�]�~;��^�i0�U~|m��Cޤ����Fy�F����++�杙���e ���זM���@����TF�|�D ���^NA�����:q?U��H�m�x��K�u�h0�1��2A[_WG	�,���!��i�ZFS V�_2��)B�̓��Y��k`�lJ�������͊� ͑�2��}�Y��>k�"cZS��R{�z�@�p�� Ym��`� �����^� �;{���O��ё1���Na��BnA�.y-�Ϋh|��E]�����9���)I�g��ȵ���Kpv���w�d>v�%2nߺ-����g���A��Q�����a��=$s� ���[(~Vh����-7�{D�\,���,�'�ס �P�ڀ�7)��P��r_���"��M�^�
@����rK��`{Ɩ]@�E<z-��k��s@�t���9TIf�fB>lA��}l� n��{@���� ���F �����F�|p
{
�ڱg����i*��wf�-/-����F���FÞ`k.�nz@��h�����V����G�t��KL�R��M������s�� \�k��RR*P�����
��mlj;����=����L�V��b����"y�A�_ڋ,�I�ć���[�s=i1m���0�i1���YSY�|�!�u̩tL��W�1��%$VW��L!�����;o�-G�; �AO�Α>wε �k������c���u�~�:�!�f��7�s����U h�Q6=�)��h����po�����8��g���_�J~�������8�>����`"�t��aH}X1�2�~@����ק��d	�������:pЁn�e:Vq�w/`"�?wNΝ?��"������lz�����6��i �ͷ�2�c�/l�ޞ0w{z�|ox >0����N�7	��Q�8�-��ֶ�d"g����D�0>;_^�_��]�ܮ[T��#���*�jdCI8��X!P ��X3Q<��
?ݶo�3H?�ӼϔzI���U��H����7�#�Ѭ�3�.Je4UU�vS�?�k��{�m�b�U�#�/�Ra�G�z��;~��[E��h���]���O��Zڰ/2������(�F�p��&�0�o�I����ŏ�=�U����U��ݪז3�Y�d5��t��a� ���*�$ci���1,~���qm j�`IZ�x�>�ӤŘ�{�P����S�f�\�WL��ӭ����<�h~�����-���֗�J"ռ��)���t�:��P& `:[����������)�9*n|�:qR�}�]���M����<z��˱cG��`�=��?0��Tr�}�ث8F38ңM|�#��+iy��j�6n����~�.�"�`�`��u��%��';���Y0X
��:3֥ǭZ��vh<�»��Dv��Q�];���;~}�~��w�2*\Q詓���:o���ϴ+��;���\�,�����m@ȋ.S~���"�[|��RAÚ����r�����Vk���T��҆�0������>��������$��&��Rާ�Y�	Ae��ς�>{YV��v��;�95k%���:?^���j���VNBpT�R���o �3�w�L+!C��������K��y��.E$Z��. �/�ҋ��v�`HΥ��4�=��"ԉ���`kЦ����(��,Ղ�ng�> ~�� h�\aQ:�>��ܹ���{����dhxį	iybٳ)��ٺ_W`��y1;�L�ݽ-�o�b�;0vQ�YS����� (��<y�� 1d�L&`4���~t�{����w7����I��z�yQ�M�ݻ��~n� ���B���VY�B=g�y�-����Q�a-0�Ώ��ʺ�k�zz\���[�������;2>>&���5�{< ֒5w���p�]{��>c�S��p9��i�N��'��p��X� V�H]�tokq�pkL+'@�Nd2I�4���G�oޞ��/�l�<��f�x�5)�2�nW��\2+�&a6ngL�`kF%�#�'l(n�|wA�n�W�l�w���Ɗ�2_��6�^�K��)��O�����bXV��ZTh��I�,��yr���!����dM#����̂�dm�n�]P�[���,*80��y�n���5��m����`i�H]\���"�n������Ș���G[� (�� �� ՙ�[��͡���<�R+�R|�v0k+�n2�����k�b�~�t��F6�l���3��ȕ?��Ǐ��#�j��R�E
��e��ط|���X.�B��p^�J�oM��X6���	̃��Z�Hل �-E��"=���Z$�H_ #������ݘ (�`��(�P�pe���qMc���M�8��x�|�y�r�K�[ߪ�ƸAr}"i�N(��f ;���H�_J���kC���}<��J��C;-kl	X�����r0��s�z(#(- �mS[Ι���B��]�Aݨ�C� �Fr�i��,��^�ա2�K������ӱ��^��SO���F�J�(�j2A�4�2�$�3����hi�X�4���w������<��^P�U@Y�E�v�m�>���f��E�`h�����*#SI5@J�����ԗ�{ӂK�����^��i�
�C�
r��`$�Z�A��٩=>�(���i�gzf��7��ٴ�F�$�TP���8{�A u�/�J�r�7��?��k�u�a�<�xH���͑�a9xp��"�l0�?y"�n��̟����,����.ȹs���#���/O�<���	�w���J���3�y��V�o7-𚷗�������`� �������6\�^?<\��FoO�ȳ�s���3��y�cZVV�T�ll��,R�������pxx�li�t`��B�.��P����'��ǭ��Sc��@78���8=��5��.���JR���2P�X��E�q/-�B���FN8f���ض~�h���L�\�5Oם$+����r��G�g ��۞]�ްV�q�@vQ;�=,�7�ʶ��0Sa?�n��ʑ��y��e�Cm���e�l-{E��gwe1�g����i��"�l� &h�U+���ژ��4�L/-�f`H�u��m yF�{ʖ�tll
608��G�bnpV��b'�����x��)����ɨsP��� �W񺹩g^U+Zt-�-� 8�V��l��	_h�2z�k��:ݿa8m2,w��笍��S���?dq9���"ZR���Fj
���P�w��|��R)����~��i\ZZd�+؈�X  ����ɟ>�\<x �&I��/�* �Q�o�%�x���N"����i`������M􃞩}��Y�>2@��E�s�8��9�&W�V�����\�  m���Ir@�����u�ے��5ܗ���ulq�BQ���b���L�D�����N�ծ �`:����4��%2$���ˮmZ\-��R0�X��A�J�Y{=�IO=��y��c�������ys��U�h�6��nQ��饲5XA ,/뮄l)k�#�Lyn u��r��1�<��W����:"����0ƊVy�	��Yꃸ�_c`k��j(�h �vV�e�D�e]߳��`���k�Y\X�յU��-����g
�{���fYqM"K~3�D�����@t�u�1���jC+������劜>sF���x��T��{�� 
��,�ˍ7����`9��g��x81A@y��#�/� ��`��(���ѣ�����_��_q��a��?�I����<z4�>��2�� +�Ơ1�K���2_s����+��BF�3���+���pFP�����	ƾ��3@V\#���<��R��СCr��b�9r主�ôQAZ���sq}ѿ;��. ?��k<y���|s]�<Y�$t���-f84٧������u'����ۊ�������3[����5;����u=��<Ȝ��j��|�IV�x���Z�zf�K �_'JN���$���/.���`t��h�x�3p�-�*M{#���3{}�X=d��;2:�e1�0�~k�'��[������dqi�����*��Hڿ���]�[����2��o��~HK��C�4c s��Q��T`?ll��^�3u��3������w�-� ���>8vH�f�%%�V��1�`{�ڎ�S}��t�1�߲;�p���;�|;ճ\����#��z����ޓ����0 qˡcg!bqtn��.�f�������w��lwb�{+��k&�&��G���\c�(��jT�ʎG�]J�a�x]�cp��@~��2=3Kg��F4` �e��p1����@�M���-D��ֹ�p<� L���~��w��9<"����w��]�Lg0��)�M��:����{�%P'�G�r�S��^�?�j�3c��\�=�����n�i��iEK��	�ŝ�c�0��v�<O��S�1�K_K:c�E	��mH��;6:�b� ��E��B�V4 �UB�.�۞\f��?����`Pq��.���0���ܿ�޳~� ���w7_�lQ��ӎ�x� ��d+�����Z�+�4U�֕�W�p��WI�'Ψ�{-�c8nܸ�F0�m���"����!?:<L�~�E�h��n�q�ٴs�g���B�`�C�	A ��k�֫jJ� ˹������zE�������P��N��4�o>Q��t�$�+�v�εh��;w���2���� Z0�n���P~�D�(����B�@1���� (���J�7X� �U�A����$�+������V��C�m@��`��J��kkҚ�f���]?VaC�3�����no�k>��"��O�?���Z���S���(��Ј�o�����;Ȉ3y%��W�n��u�sǂH�����_����Tu�Y$��Hq,�Ź0C�����Eg�?�_��E �x����F�������kB�*������#r��nvj����.�ɠ�^)X����P�[?���O-�'�{�:^l1�ß�%��ւ��B�څ?���b�\.֭���@��r���+��B��l����u�.���[�I�8�m�����ڜI��v�h�fΎ�M���}����-�Gk|B�k�7�3gx���5Y���B��KH��}­���pƼ���
��ԁ�!��f��E�vph�y�C3Y�R�m��x`9;��<#'4�O�>%�߾,o��l�$�Z\C;��q��Z|Ҭ#�`��B���S�I�k��g� m��p=��#U�_˴�=u��2 �����ɓd�o%B�z�q� �1
�,�FK�7�����R16�Vk�M��ͣ���@����ø4pF�1b2E��N�<��@ѝ�Q���_��F|Z_P�1�8���V�j�����Z1���_qK�5*�5�<������	���~d ��:~D�U(��]�%���ˬM�Bq��*.<.�{8b���W������0G�Q�T��٘�ϻ��R�kqi},1�_;�U��΢=�mFt����krNd.���(]^cP����itZ���d�)��-T\J�^,/-q�|��q��u F��˙ӧ����E�玸=�ɟ��G�󟿔�%Yi.;�>%��I��.�އ���oȴ1��v��,Vw�\�|YN�����L�j؂�I��l�=��g�o�o1֑�u���r��M��#�Άp{`Cf�fejrJ�ܽ#�?a��X( ���.QC�����젉	�=��{���=��B��\����4؜��4k#$(Q c�):G�~��!ˑ���Y�.4�ossս�����i4פ��Np%Ϫ,����Щ�Y�x�L<��陇�Fs}~���\�gg96��T�ʾ,[_@0tq�Ǥe��jߝ�p^U��Ν�Z�C��nC_F������v���� ~]�9Z�aM+����eܻ}��Zօ�X�7���ż)^��m넭9E@J����{֊���F�5m{����G�ۺ�E���	c�H�<��� �����5�_T�,����h[�&��[Ya�ae>���\{��a
��Xvoܲ[ �n{Ӛ��qp��h@�B5�<Q�G�y������l�5�i����S����3>��y��v����gfzt�s=(�W��t�F�N@��C�t/^�(��߁��-'�8��_�ɬ�`���[j�����~�<l:�?ɵ�M_��M��΍��RḁD�/�KJ����\�v�:�`9��}ށ�s�4�VV�"�����
���Z��E� �vܢm��X!� U2��b��5�X��v�<��xM������� ��h�"^��i5��Vg������;>����{���{�k[�Nm��qh�
������%�:����q��Y)�P�
��d��Z���)��J�Dq�u����E`	,A SP����'�}��x�����M=�ݯ����v���p�D�T� � �0t~i_W�	3 ����O-[�Mi�N�4�� A �����r��a�3 XaW@B�K0�n��x`(~�Y\\�[�osR��  "�qZ���= ���%eG|v��l�'Oʕ+W��w�a= �=��c+1��w�B@��~#'�f�&�����[n���|D@~��!px�6\�xQN�<Av3��G�drjR����J�����S�o����` ���Pr��0uXй�B�r��]W�i�k=�k>l���b��fgU�k�xp�|��	9p`L�={&����Iy��,�����3��ӧ3�f�"�2 �u~a�עD��Dh�~���y1��}�?�]?Bw�ַn}/��?�8;{�,�v�~abxx������S��{���=i@L�Ĳ
�����\�d(��5H i��U�1�R�|�4-4�I i���ܺkz����)�в���4/>g�y��.J�m{�ٞ������S�1�[OFd` a��M�������TSg �/dueU5:S-fXs��3'q8jOe���?������@�[!��,�,+X��DS���IKǻ�	�9{�9e՚�d`y�dV���������8��K���˹:�-ӉF��:���}�Ή9,�/\�K�.��g�u"nm?cc�Q��τ+��������\.������Z�^��Y�xvM2o`�`-Μ��!E6�K��
��#��X���J;L�F6pmּn���M6��p.�9J���s3�^[*�p-բX�]�Fuh,5�1u�B��/zcE䠕SD�C�gD`�΃45����8]������5�y4�e|헬��͘�Me�z�T��7b;=;ܣ{e<�)}�L�Jfo��h����������l-"����~a�o�*�kJ�Z\���@I�C�lhQ��/�l��JES�1��J����}�h�������F�TJ5�$뜱�sk��o}���\�"�� Tz=)>���un���5|ӌYo��FEiKץ�:-�Uh����� M{��L۞�5^�� U�~�7 ���ۗ�@�r�w��/p���R_�&'�ƍ��ѣGʠu����s)�f`T��������Aj��(JK��6h��!�Q�J)��6o2�� �����\�����a���<yB��ť%��t�������Sr��1���5�,��)H\����f ��W��\�h1�~B����q~��sǀְ�4X�����J�5�$1�g����ݜJ7Q�E۲Q�d�2��{@������F���N������������9�Ι8�)'Ng1`خ�',������x��="��N|�&��gϞ��ǏefvV�?&o�uI>��c_pZO G�!`��$���3��vG?�o�D�y��f�@��16pa�di��ՈU\.�2�k��l�Ԃ��t�r+�]���m����v��V��u�@�~o:�_!(�,+�����N��D�,��Ò��Le8�H9҉��	k^�O����v3G���� +H�������{Y���|z�xFDU�gZ��P��o��w�.X����x	|�Jn�Կ�Tw�q��~,���� ��\�@.^�DM<�c�#?��B��`C�h�]:}.'�X��3\��[�3`�� QA�p�|+XD�nj`iFmT8m�\u��5��MH�3mf���A��ƒV3��|�X������3�r�� �sg�҉B����9��4���@CS�Z3:� ���K����ƔW�
��4w��)+�w|Bm�Ջ�` �/Ph�S/o�F�x*#+ߴ'1�R ݉��$��SQH�|���N�j�V��wTP^3#��˟x���|��v����������Z�@[�C��S�\��X沛z �Qk� x�nX� ����P�i!���0W��k]:�/�5e���98YǗ�w��[_X���c}�|MR��b����b�l;p[��8����zg����Hb���A�k�M_9�-�=�]��kBp�R@�K�(�T�6:2&�ϝ�{w��׋r��U���H(����q�P�����o���?����j����L�+�d��#n��	lU<�RI]�"JY|�̬������C�wU�sM���k�s�퓣G���R����ݻ<�> �b���/�+9w�,���}������	���f�ϋ�lb~�~�Fz���~����~��]#�ck�|f��f�`��C@N���MBc��g�Ar̫Ʀڋк^u�Z�k������24��<4 _|�+���,-�ޘ�ťYX|��7�����p�ꑻ��ՠ��M~�X�53;M)�kW>x_>��#���NpW�y�@=���)�7z�O�}JO]�FX_�6sR�I,��4�Ų u���0�9��' o����~ak��_�B?�m�׌I�oܗ`��a��n��['[}_�Q`�ן����v��[ss�H�m���ߺ��j�҄���_�$@*S�&"�~�Y%��m{��%Z��<�1�[�(K��k�w �Y��n�i��)LO #���M��YƬ�����Mt>NӀ�Ш������r��q���;�\���+��`����¢2�r�#��[��u���0XG��Y"�0l�ݳl���= � �D��r�T�X���9x_mە����:YO� ����2�xc�9n33�L#�رcr��	V��w�|�٧�;����=�gA����I�_X�����G���ެ���CV�r�q��>����Z�MQcF3�Գ%ӂ����G,�Fv>���V{{���V�/����כ�|0��Қ��y��J����x�E�q���L?ZI���!�@�d��1֮�OdyeE�=��S�����_j�{�V�ҿ�]�Km}��1�Ҷ�R'P�b��-�@æ������<�����k1�ettD�n��"5��K� �0�b���=��-�i�_R���+	����4Mwck���Ң��3~21�v/d�a�Q`���+�A0`�����[e�Zھ>���`��x�� ��� �B6bs�!cc� �=�ﭬ����0Q�bֈbwϞ>c����6p"k�s�v�k�I�)�u�~�����;r��Eu����=�W�x�eA�n��<�rܓ��߹}q�]�Q���u�Ʒ��W_��;w(��s���}������#��B�����ޏ,,[w�߯��0@b�RC�a�����(u�1簟bZqH����E&�Q&!�����P
�����㆗��X��+�]}��o��w7���r���壏>���ߒ��c�����s�:t�kǃ�Cv��1H=08�֓~y��/GIZ8������;�_��]9w���fa�~Џ�O�&0�B��4������o�iH����9F�Z���� ߕ�Z��2^c�F���N랾��q惾=��##{d�ǽA�^���*sR ةp���yK��ۺ���
 Ͱ��{X�e0���˥ f�����_K+o|p`� | S��3��f�~o
�=ߩ���n�W�
'�##�d�3*��(��
̹���ORC4˳6c� �X�&��\��ܶ·��
�۵vV�F��[z/ԧ��#�/\�@me�������ݵ$������i�g��Yjc��m5�#��Xz�ל�tG0�h؋:�`Ƞ�{���S�XW�V� �Ɂs2=���>�L$�<@a_�q���8�`�1�S��676����2�x�5紃��goNS�F�5�y_��j!>eBٵ#�����|8&�/P�qd���g3�����27;KF3i�����^�I�Gc�i��{����^8�Z�(E%%�=��eRL%�IpU�"�͖�;Y�z| �Q���:B�D���dz�z�bF�m?{s6l���
 ̳�y�����bMY�)���}��-�R���㡢�3.�s߇�y�m��/ċc��X"�&a�ࣘ�`�B�및��Ύ����jC�� ���}F
\lw�*�����lӬH�.�{Q�侂b����o������`�L�)�R����2-tW��ݑ$E n�)�~Kw,Ÿ��X)ޱU:����?Id; ���N6Ч���yXR����`|E���$1$.ګ�J��,��.�w@�qinQ?yJ��gӳ���&��/~��z`-�8/��gΜ&�vrjJV�WJ�H��Z��L��0�� �{�=�:��}4�%Ld��m��m�&�ik���C��_ȓǏ(����`Z��1�<x�p�ҹ�g崳c0nߺM0���<D�YfY���d��$��C���P����:����%�*>@[��U�VjJ�W����^�U4t@�*��`�.-.�ջ�­�%�|�o�}рu�R\�o���ւ��A9z�����Wr�а�k���{�Ξ�]���Y��*�x؟ T笴�a�q�>o�-�`f7�p��Q��w���A_�^��v�����X��ÆS`��~!{�� r(D���`WT�1�az��X�ҴD�H��w�!��Z�U��Q�?���f�&ە������E1ʐ-�u_��5�=e)��F��U���5kFlʄk���\��&It�,�o�L��E�.��ZZ��� �l�_Pk����"I�$��1wۏ��L��n��2,�F��j��ka�KE�B)%�;�.�9<#93��_Cn�B�u�����C��f�;�S����g�5�i^h?��@�R�T9'���3tǜ��"��G��E���aQ������4�5�0��5��_���<�T��7��A�i�9&�|�>8l�MҴ�v�L7ő�`�a���s��SS�i����s����+�hm�A X���L���!e�y�����
��9� ���+r"p�l\��#�ܾ>VN�qD蜵��ȋ�ѪsD[���^k��TE�6[<߀s
O�>K�����w���w�7��+�ߜ��w�+��5����A9t𐌌����#vu:u5�d�Xq�5�7��E�;'uh� ����3�wdb�{�WL��g�7[��C��H]4-���`C����:����^�0�0�\��I�)�f#���cyc�X���P�<g�����	�+��ﰞȻ坤��[[j�[+9��XFgo2�I$h�3�|s���ٳi���R���vu�m�d�wpG���&���,a�:b���ߚ�x*ksvv�}�5B�TU��P?=*©lxP���;���z�bR/=�{���_�H��������m^�}7����?�⟄,�1��Aܽ{��V��++kn?[���9w��|������l������\�ggg�������Wu5�\aM��hn6�����������A��k�VTn�}n�������vM�#����S�v�k�����r��52����[��O�<Ɏ�>�=�����/����ddd,Ƽ�qv�Ø+�;hC�FG����X��������o������}�bL���`���X\[]��w�ON;.Gat��|���E��	��+;��*d9z�8�[�[r��[r��C��o>��������Ag��?�#��?�ܻw�]��[;�����gF�OJ�r�q���#�
���������1�E���,�K�R���Uw�a��ÏT+>K������Z�L����i��O+!� ����6��PDN���zak�(1�PPѭ��;B����V��������ʐS�l�L�]�V1���~�8�@��,G���٦4�&7��k��eu[���6��a+'m>��<&�آ�V��^�(��[�$���4��R4K�.�ԭ,�Ɔ�,�@�juU���Z��2	vrr�n�,�n{�������3]�4��%P�e2����
���þ�t k�F�(�5�N\Zi3N��[ (���S�?>d�͂��� �w`� ٺ���u��IA����V
����_�e��47~-��S�j1hFp�����0��Z�	�,D��5���߈�k46�'��N'�BBfO�?e��(�ς��΁kj����W��q�����5�YH���w���{(@��l�,z�dOA���S70~�o�-���g݃b> vW�d�]So_/�R�> e|,r8��?\��Ky-�nݢl
�>s� ��w�<�Ł����Ç�X�БF�/�S�Xt	R �+Hp�q}J0�Px� �ؐA?�9�~����Q���4��Z������:v��� Go��Q��Q˪���V-��,�iN���dY���W�vIw��[q�h}�p�8���(���q7��0�ڳ=�a�"l!=Zb�ٿ}o�f J�=����(�/�������j����<��c%k��;-_�`��}mw}��;�ݪ������)v�s�A�60������h�p��޸5��/À9���\�ɓ'�Ï>�˗/�o&'�'�=u�LO��Q!H��5i5a}�����˵��K�匽����3p�={G�o)T��g���I����w��"���>���{��]�{����o]�Ko]��4>���8=@e������x��Q��ű��	�wj%��I�YU��K�����;����T�}��a�r��o�OeHc�]�P�-s|����ǎ�����
��m�`�R�,ᬚ�:�cg/|��u����������46���W_�{���ђǏ��^���#�1�;A����]̋x�$�M+i�=�����u)
��_ ���5�-������>J���a�pO���fFif��곽BƟ_?��ѽ�����h6�O�*o��$�t�ֵ{/��g!y��K��"�h/'�c`��<X�џȎ�}�u{�%��ۺ�C�y���n�xB��/U���M��$dB~Y��t�,��m�]���X"xp��h��&;/��'jgd�v�K|v_^t����i,�0pBY�-�h��H�.K�s�b{V�,�c}���Vv�1���P6����z���c//�C�n"ʼ�fKu�䙹̳�X��d��a9w�AJ���>6���[��U� �vO	�N�Є�G@���$-��bʧ2`աXr�"�p���)�8v% �`��.>��:y��o���'�M�H��W�1��|�|�?2�3�7�N1�s�_��>5�8@_�3��Q��WH�Toj���&>t�0�����rpl�������;.���tT R�i��^��٩��x	�C_2W�[�n���j�H���~dd��2���sNb˃��Ԏ�s�C�uyy����s�5^��tܚ���s��y��>7e���H�[�$b�f�9ҙ9��Q����G
൘_���c��y�r(a��wh���:�;1��!Ƶ�S�7	*CWAo��s�Z�&'To�������3��<�oc�J�+,���9<L��i�����nl�������w�G����S[�Vg`x�{��_R8K`��,{�c��:��Ë|)�gD�a�(ڍɦ��>M�\k~��ɂ�6�=��~
f�>�D�|xEΞ�,���re��*{��V�,�Br��\ M�҃�� ��#����'n޼�-nL9v\��i��� d���cwd�F ڼ7n����j��^�{���s�_� r��ٳg����2<4,O�>���v@�{�b��W@y\�9JP�)��6�B�"�w!�  ����S��J��`������,���Lh�[�vP; �&D.�������A-�A\ʛ�����4sN�?�'���������>��=��9;dUff�ߋ2;�$�s+�[����M�۸�z�_�N�0���H�8/���.@p�`#Ui;TB0E	!Q����~��7��@FX�Z�6�	r\��2|�L�5�/��x�����籱�E��W@~CAcXS:M�8��@�r�����}�eYĭ���c����`�����}�ge�8��
����Hn���[�|�?6�h�����ӏ�<7 ��Zk���8kl�:�� O�Ü��u����N���~�[q7�(]x_����HA�N�nۛ��"�.&�]e� ��Ā!�ێ�kJ���L�:�y <�e22 A@-�� ��ڛ�b���a�Zh��b�Z6Y`n�,Ӡ��O������ɓ'	V�I5��e�Լ$ӣ�`��9O�����ߓ���S�8���s@r�i�FP��/e*/��Y\Zt���W�ςx|Hh\��8_�阘�$�P��^�݃����z=<S2�-�@�R����:��1FȌk6�6�hn~�E��$����F�Z�����?tp�}��[���� ��V�d����1��^s0�3;��И��g������?�[/�c�� 6��-�~��l2d�,ҡ6�*��@���lK�\���� �~�5�?�YIptq��x&_~�%��I�S/�Q�:��^��0@8t�G�gV�����#	({y�-��j9b��Q0�K_�{ʲ��j��m��tD�V̑]e@�����]�#��ť%�!",��y)������V��X,�m�s�(��}�a�(��"�#�����| ��`���@��q���@��Bl��m��~�k��N��;�h��|ۿm��i�|�5�i��<�=�����{���4�;�����`��81����_~�?$�;<��m>��Ԭ���PB �2�[v{�G����kZ쯱IV��|�v���}�`D��W�b!��>�L�y+n���H�5ח�\ć�ȣ}�xA����gO�8F�=̝�ǏY��^�ʂ� B�������L����k~��T&>��N��|���<��㰇�={��U��}	���j��	@��v�`�b�K`i��aOA���%���#�LP|��ߗ���?�
0 ��Ld��;(ͬ�>p	��SS���<v�K�R�����Y����g���!�������rY�g&��W߻}�[299!����>M���iCTBZڎ�N�Q��� }o] O�����#~󉻥���\�ǰ}X�ŋ!��l���5��U�ς�V%�2�`0�'W{O����;g��4z����$pU���#�k�Ăx_�OxO�VxØk��4��kj�e�p�f�\
t��Sԅv_��X�n�^,�%���lޮk��3}�4�b���{�Y�`�|�_�Vɋ���r*o�%}����R�H�G�n��ZX���5�f��=eza3���?h�����{�ũ�����;ayܣ��m���~�g���)Iq"���6,#��6��HٯΩIZ�(�����p�<�U��$����qUS���V��uDR��?q��pN�:E&S�Z�c�E���N�s&�榝�����8���Vx�)����Y����Y�k#X�Y�p�\_��Z�cǏ����{e:�;%+�6����\&�v��,�1W��#d�h��*6\/����ŲL��VY�Y�U:L���7��8��fff��.���:Y=yK�Np=p*��XxBp2ǎs�u�Lc#Z�i�?K<u�k�j�|�>��{jr�L�O~��k_-_}uU?�"�}��ԚL+��V�����-2����[�g:<~Ƚ�D @_�=�#c�Y�	׉�F!�۷�8�~��; 0|?�Nh�J}�"���Ƣg'��e1���5M־ޢ����r/
pEgk���Od]�Y
�6s�����3��ߺ�U�U�4\������I2[!��^��i۰/�����`)�s�����VI�ʃػ�@s�- p�R-�x��q�t$����r���9\����䃼<��m
���݋�wd��vW��til����'�k6�T��=�5��1�^�y�=+���t(QS���B�׾�&_|�9�m ��G��C�3�r������!��sA�����2��w�-�z��v���&�?��]ߠ���;w�� 8Tm`�G#���A'���z����]wϷnߒ��m�]�Dq[�0f�8;��r���#m�Ʌ��S��5(�E�L&��˔��@��K泥��#�!P���аܼy�� �c� WV]��r�� k��m�Fi+��I	`��F��h�A�4 w���k����ݾ|P��o�����[�����0;7ˢ��c������z+�����Y�M�����=�/��ε��=�U���w�m���9�p��_W���~�g��nMW�R�|M3���H��D��� cQh�{�9��Mj��xM��r{����Tǯ��@�Nv?�y��� @d�F{ޮa�~��q�)
����^u{��`���Ev��w����������ͼ�V�����b���,��o���y"z��Z�!zW�|�3���!�!Y ���o�F�w�ݷ��D1s�0�r�JN��z�U�ڎ��V�ê�Gڎ����k:�*
�ǃN�H�EPHD�{^ �d�z�K�6vu���~U�Ɓ3]A�Q�nEewǜN=�K̯(B��h s'= �VI_�{�'0_*>uis3�uTRw���OY��Utt�g<�9���>��q�JM����E:��;k�������NL�g��uUR_(+z �:� 4]��f�(
�!�V�x���� 3��k����� �s���0Z��B,�i��i]\r}2H#ipp�:��}�k��M�+�u
�
�	,�֕��ܵ���s<�I�s\0�|pl����2�78��B�gN�}�`Ԣ �� i�Cu���.��R�P�T����4U��/�;k���Vl Q�^*�,����,�
���{R�m��Ilf�H���i�+��mc?��Z�w�B��_��$\�l��`+o �s�@��2mQ��1�^HM��R�RE�l7��»���ݵMo���5�����eV�|m��_4W�'�p�Mݧd�=̡��X
����X���j*((�Yo�_�~�C��d�J�^��X�xMèe�����"dV�,.d�5-�zM����[ul�O�ȲX�B�2��菏�ɹs'�z�m�� 7k�*��3��A�!����{�嫫_�կ�r �S��"�E�g��CF�嵖��a{����G���"`9�[���������7��V���y��-�{6~0���������}���ߖK�.q����~'�<���5��(���nh,|>��t+����
���C�ڐI"��,2oX#@��k��l	�s�]BY'������8��V��'�P��а��1�=>>�~*�{�7�TLB�� 0�H���� �e�[dr��^���[������E��W��Űܾ}�]�A���g�wܳ���N��10��]�L�Gʠ���׿��oJ�@��Fн���_�7�������m���[�I*�����,��*kV�ޘ�k�K�!8��]�)�J���A���5�r��BQz���D���Lhó~I&���[��w[���-ڸ^���F���E�Q�%�k � J!��;/�X��E�L�5u�+m]`����X�:@0��v�7�AG*|N:���Z�>����`�C���ͮ�G9��q��b�.���["���o�c)�v
�U������l���������-�MV�-���)Tg�s�.Ms�Ŭ�TK�w�3M�n�5'�c&0 D2ۜ��a ��/h�(�u)[Q�F@Hn����" �n�t��my41A'�������T/����2�>��ZHb�U;3�@
 JO���t���18(gΞ�S�N �S���$Y��Ϧy�p��FG��
��ѣr��\�zMn~wSYI�Z����b=��G�ɓ��`�jt�Qpolt�N*$D�Q�c�}W����gdx��gj~�� 9����U�Nn��}b�����Ȉ!ۦ�LM�}j.���w���ߎ��{��}�����˿��o�%>�HҫW��_hSB�qddԝw^6W6�$��gc�+ {OO��3��:�gΜ�w�yW�_���t�Y�h����>�r�
A�?|��|��vrr*��Z�Jƹ�A���S��A����7w���XuϬh��k5��}���ڇ���z��lW�l{���k��~i�+�E%�R0*^���ز���`�2莢}�7�	jnjH���b�N6ƚ��b~���/�I<���_ݚ���~�Q1}���JEu�g@s���@7�oo)��%V��h�`�dC��� �2���㯇�6z8V�ډAe۟��PL���8'
�1{hCǄ��ɢ<o�~�g+^+G� W����h���݋-��Ўφf�@����E��9Y[��~8%�����/�/]f �ĉS�g�������f�R�����"��`�����s2������,̊=��>z:���c��w�o
��k׮�?���'��&	P�:0*����K�WD>y�����7�����N�2�Z`��ֹt�u����q>��(��-�i�C�@d��6���3�D��������0zXw`ԯ;���]��{�64�}��(G ��O��S���믣�_ 1u����V���x'l �Ћ>�������(��a��8�?�����F䣟�gu�\�~��`������K-���޻$����r��iw_��O��s���MY���Y�
sב��h$Cdk-�dS�?�৪�7 頏�`���yJ{:�b�74�fb ��^l�1i��f
��DN�լ�������2�<�mVanZ��}غ��n��[n>�O<Y���b[���ꊷ2�!�j'T�N@�e Y��|�����u�埠iE�5���X�LæҞ�����*�)�)'Q<��Mˣ�{�����u�˶ ���QQ�8�=^����aZ�`�@�u�����H1S�PS;��XNBƘ��j���ͼ���^�9z�d�f�8�ǝ�w��:J�1���M��zK��W�3���$N�?������X N8NpR�V7B���M2����X�cGO�c
֑Ðb8B98��s��c~n�}0ҏbu�,�34�2|���c.�?O�/ع^��jE� 7A8I萀M��gR��"��B�ׄ�a�����w�9�ih$��x&�(˚�!�:���{w�2 �VS�Ԕ��%��}=d=��TZ���{�}��e�p�|�+�H�euh.���Z��d�TR^s��wQ:��s���.9Ǿ�o�$`�\����<�׿gΜ�B���,8���$�E��ބ�V��7
�%-�\|Z�2p�i�h�՝{�Ϥ*�����A�m���A�v�9/���M	���(¥׎k��o'ٵ��#f������&��4U6Z���������]�c�e��$� �6�8 ����TI�()�˝[��#�o�ޟ�������s��a�k�~�bn������)�1`>�-���p��:Z>M=נgK3	�^?kE�1�m�l���=��>D�޶_�>h�b K�B|�-Hx������O����뵇'���Vw�D�~�|�\�N��􊆊�=\{�����YnR��������5�|�G����y���>�"���͊�����"Y��S ����$-���G�ȩS��� �S�om�+�������
���I�u\���$�k�W⾰2��:����,���O>��#�������'���Z\�I���ӧ�������[�{���:�Ѫg�2`S��b���,~{����f�a�rl樅�0K	��[��9DV.�Z�ǚ\�Vn��T�� AOfEi�����E�[-֫�a`����ކ=U%=�߽sW��������Ȑ�?��Ɓ�nO?���~7�h�|}�*���Ȱ����ǟ7&���� ��b��=���&��d�f��1N	2�I=�"n�$�B�D��� �튬�
�h0��B[�px�V�+I `w�bL����Sٚ���G� � �_g`���0�P�ǆL����=�����z'e;O�'�G�Xf���S�2��J�k�MM�n{���Ԗ���^���o+� ������TgJ��Bm�{���1&C�!z���H�����Yo)ZD�2�J޽Z�z��O,W(3ѣZ��������b3�TSJ���6��Ҹ�����ޑNy� e��h0��v��� �� "#-����r����do�ƈ��s����r����>y�@�M?Ӣ*p�
��<59I�8_pD�W���6�����^h"��XR �qe`3a�˜s��&&ʟ>��.�by�5"�w��s��9�,en�\f�������ﾓ���%���2#X���C���E:�S'�҅r����p/
+�f�g��>�~�5�^�=G�ŀ��/�A:-���=`�gp�~�}|��T�S�CZ�!�� �[w�m~~�F4�����;�����c�f��\&@�I�Q�T�#��#,�4;7��D����z�:� `H��p�����>��޸q���J�s���l�q��9�?{�ӆ�8ҁ�'~|�>�ڀR�4��}?8�!��u:Up��Ͼ���Vvr��`�c,f��N��	k�2�vˈ-y���4~����S"Ǐ�"���e�;1�3�K���������;�VN�ߣP�d��X.��΍�J�k;3g|���J]jnߩV+���L�<�ݶ��&�e��뉗�B����oi�Q�G�u����ެK� !2Gl,���@��Թ@B!;0S06�~l����R�;]�ίY�}�<����<�V}��eh�Z����[����{�&�䞛]fVt~��8��^5�lFAY�AFB�T�{���v ��F ,[��;�C���`Ҙ����y`�][Y햌����lp��1&��� ǘ����{�|���p�I���3\�;o�à+��ƺ{����`��nyM��V	�b �L69�W��h�h�0�'�xp�s�J)�>y8�,w�ޑY�繞!����=!�
�s
vo�~���ָ���u�6�I��ƀp���5�l�h���4��~�9rl\�\y������B~���O��ģ	�;�c>~�(��,�WZ
�g���s�64� ��������z
��ܽ��mrc`�s��>�,�����2[���H�pm>��}I4@�p��V���nT����=�$�T-���
�6��gZ�����@�kO؛�(T��mm;���۾#�u[�V`���Q��fvX��O����id��8N�g�\�ݬ>��&�9�n{E�,�hM7,�@Sok~N�9c��S��N��O~� F 6���a�z�N����7*�ԕ�x�����?���j����θL������w
�b��`q�!)�d+�r� m�vPY�(X �� u�a�6-�����ϴI�ˈ��[+�N ��p�"�ZM6P����G�������:���}�=26:�"uO��Q���gt��g)���7���f�99G��?��\v�2d�5Y^��ɩ��)��ٹYq�ښ��M]c���1ιh|��I�.+@U�[ C}���/����3RP#-�9lx�����:~��L�>�h�O��3�hK�s�-��q�̢��p�W!r�$8~X��|��S��0��0����Gt� $#��Z�� `���&�+��mrJ`U���}�;{�9��ܽ��ɓ����α�W�������|�-����'>�$�f� �[�o�ۗ�v��gdR���_�������;�Y:� �N<�}��p�"�_��7���E�`�x�\�� �U{��S���	l���X�X.�j���f�����5��hqꭱ�Lv@�m �<�As���0��3c�����ӌ�,��2З���� $В���/(�	�R���Q��31?���3��u���\�bQ �R�]��D�Աb`A��cn������-E�, �\��Ϊ��%b�$Z��ceu��7��O�y
�4�Fk$�R:f9hj�_d���ת*�d�#�aM�  @?�"�eC��2�l7\�i��j�>?� \�LQ�v'ȗVB�Ud!������p}V���lczYFI�����z�ꎌ�\	&�o0��f��i�v���޺u� ����*�n>�����_ʙӧ�<p`D������5:2,�n�M�Z]�9�?Av��+��^J2`����m�X+�;��	��(��Ɋi��0��6�`���sW�L��¾���43��=vtt��؟?��|�W-�Cf֙S��m��ߪ>��ZlO�#���S�sa�s
@i�Ak2n��^����Y�{f���.�;���V-.,R��1X�62��Z[U;��o���ld�'%ܾ�y�}��ӧ�^���,!%(�3����ѣG��F��ڵk����p�]ۨ��چ|���)#v��yY[Y��U���;�y��L;����,$�L��Çi3n�Y^�Lk�!��9^��k��֤@���--��T|0�?'+�̅D߳T����
�!ޯ�{5p�jr=�T�O���dgL�>���RD���1�!��Z+�`��-��Δ�ۏ,���վ?���{�֕������\�K^���_��Ft�����L6�n��t�SfG���pk���ڤ◘�i8z,��G�u��\��?R��C ��Eg�P�������m�l�#%
�&6�Ϙ��ɱ-k��9�q�����/��D���DP(���&���ŲFPD�1�&5��@ |fӭT�i���qn�L.($�K�>�h*c �y����8����0S�y�*�@�+�Pq�3��{��\�񁁎�2`�ኵ���[������IEu�cǏ��Ezr�<��K�0��W�Ȋ�����τ��uޗ����4Tc��酃 )�ϞNX������Nt�,~�ԝ;{�,�ɩI�{�%+�� �3����r��fJ���Z�Kk4�ď��pO�=�;t�[�0�Y���j��U�=�8w���A:J��l0����9���\5X��;u�q\��__�3�����}����ZTp��!�T��]��Հ�:S�1��P�w�������:����{48������76�Й4�N�C�g�S �V8p���-)�B3��XPƺ$@��+�f%]�
 v�MA����(a�9������Ax�~���i��~���HF�����l+����*[��l�:��2����(���<�U�d���ſ��B�V��d�,��1�{�+��8IS�q�L�ԃ�a=�:��@�(i�3B
6�C����,�>eCfi�~�� @�����b�y���!#�N���\�U�]|���9�@��N p�Qf G��<���k�s�����,gv[���++�����_���~cMC�]�Y�ŸȒ,��*��J����vw�V
:��'�.�@ ''s��n��	�c-�Y�:��VV���&U����B���� �����>�����GF�ŋ�ۗ�����S�� ��=�J��
�E6|�찬���`Cv
� d�i�g*������5�y�]�8e����嫰"X���(&��,�m�W�ԵF��Vj�(hR��f���i�DF͟��rQØ�Uco��h� 8�ϣ�1h� �0�p� ��;�n�z̦��a@�Q�F��L�j��1�Wp�j;i�ǩ�Z�Ad�_��O�8��p^���R���j��[����/]�D����a�8�b�5\�~]�<}"���|�!��m������C�k9t�5�3ľxn���F�6C�V�9���,:�%�[�06���q������~`�
M�\FAR��Y|���@�ӽn�:⟍�� ����x�]w0�['YV�"�1���؟����_����_Md�Yooz��|�RH:�a��ߠ�U�����$X'���h��T<	�H�o����u���� �lб��p���,���E�z' ���`3�1�na|����
�|�.t��C�+����īm��|�(�Z�+��unZ�78�	�ݵ�j�k���7�wz����t`9t��vg��Tf�u0\� ��H(�,�iϜ9���j��2�?��~�{6��N-5�{{DB��&�C�9L��E�˫��:g���1g%w �W�^�۷n˽����	�V��y�;'o�o��~��WL�4b�����prp� ��DP�B<=�A�f��'��v�9��O��>���i���G��?�����`�0M��=���ǎg�ms�	MZ�E���2�Ѧ��S�d���;����ݵ丂�L8�{j@�+�P��K���[�?|*=}����!}�>�@�Css~��i:�س $�<8:F����nȹ3g�sz���q�����?��:��+�_�B]�/���|{�{��r�����L�>q�8�Q`�C����Ċ6p��x_�u*��m�N����U�0#���O6-j�sӊ׵^����7��Q�N�;��X#,�ɟ�������O� �6�V�V�U��!&��{9���[Q��蚌����n?��fiK�?"���H7ec}S����|:�����v�g��R�����c��L�0�Tnn���|�<Q6��5+s���/r�2k��u�
P��d`8�������=��م*��"�:��T@��P\ Q����Yp4�s<~F/f��m�a�`b�%������`��:Ń�O��_�-�%��Ll�,,�yj��1�p� ɏ�:Y[ϋ1
��o��I��w7��D���z�C��@�2
�9b�f>�D�s�Z��?�!�@5�^~�����A^�ٙ͝�k`� ������Z��Ɗ��4;;#���e�YM`��x�rn�k���c����������5���u��À�����<�Y/4wY쭢�j�!�����Q�bv�;48$=c�,�,�a��~���wn��y�L<z��U*��(��/~X|�Z�=����d�?
����\�Y��/e<�wQ�z׸F�J�+TB���#��o߾#�~������k�����?���)`��{��zA6@_"�̹�0�2�l:����1�#�OzT��t_�����֝�ޞ�gX'��X�{iX�	"g��Mk2:6��R�myM�� ȇ ��A�����ѿY�_�$Gp�z�&_�����U��_䞒�y��ݝq�?�\��I:�#������F��E��1�x;��K���Y�����_��fV^]���1�iA���/f`�%v����&ɍ)j8��U�� ܋N�؟�$SS��y��E�w�
�Hq,���W�	�xel����X������C�/�~C�h������O�� <����e��MMg�|��ͦ���UU��E���Q��1��չgӕa�1	`A�z(`F*�6�~��8qR��z�]�5���n�]v�^���Q���<|��,.=p�>-S�ف���wh�B߰�ٔ��YQ>����O��sV�h����:� ��{��W��[�ZtӴ�NܣE[6l:�)x^p�Mf������xC�$am˯/	��33����o��"-���Sdk����w�կ��i��GZ�`FM;g�w�ܑS�N�a爃煺��7��ƀ�#�uft|������[�?�奄��;��'\�d�g��=w�i�pڧ&'���#�޺���Tn����x�hJ���sN%ҩ����2�f�g�>p}��Ϝ�^�#猂�>��r����gfY�	,���yG�zkr��=�tׂN^��V��Ѧ7�(�P�3�X$�kJ*�LЋ���a�� �8��K���]]̆T���Ӿ��HNp�m ��;�d��i��QP6�i��s�]9d%��#�c�e�' @��Oo��ԳX+Rsc���:�vvq}�oשS���	H!����~���?��>gޜ��|<��&��uIr�l3�N�գ`�@jc*C�н/즂�[vhbFp��y�?���XNهu�N  ��h508W=xa���<:���B�A�O�U��,~����{yi�}��Y���#���A�� s�n^� u�\�{ �0n!}��EI>y߱�Wp�b-�����hK�J��Zl���}6V��5ŝ�D���`V��Ҵ�,(dW_�`^���R)�A�k��[��̏]Ba~�/Z�R��i�v�ƈ��>t�\�pQN��
�Q�rӭ7��/��KH6����N����^�������.�n�<
�~����7�����r�Oe��� ���v�����ʕ+�ɯ-Cn���2�%1�]���-ӵR=�f�����L<xH�Y��#�c����k�sMܻ/�g�D!BN��L(�SW�J�����h� /�RV���.04��>��;���xùk�~^?�z���3P���o|sC&M��ܯ�;��Ѕ���Z��^
I����q�@��/�ELt�~����:
���;Y{���
��D��ЁA��>�bM��_}�s�>u��Әg�g��v�G��_ n�����[�Y�$!A������@�^rf ]P�"�|���3>����=���̼U� A�7��$j�e���nw�{�������_��y=3�[zy��lK��o$�}'@ �W�;yNDd�-Ta�"K"R��r���D�8q�G[�m��O���L�*���O�ǲޔ��$1L�٤#kw��T�'ۧ`z���<pN��zq��u �g�T�.���/�OP���Or?~��̇�nN�b݈����I������걶ت�{�������w�d���_c��[��.̿�.�M����Y��䟶� �O���*���x[\xD�VX���[�^������lb8�6�m���&O��~���f?0}���O��������|�d���mu���3��13F���,Q����dzs��VavD�@�)ne��^:�W3~�M ���'�RRrȰ�ِ9�f����:�ևU,�$���:wМ��04��
����E��n���S�xa����&�\UK��ଡ�Ε�W)�@F��Y#�����q� �4./�q���о[aA"0��Np ��Xqހ<+km��h4$[�Uh
��e,�� X���z�p�ܾ�Μ9�"Iǃ�>48L�
0�����.��3K˔Y���ѣG�}=F���
�	}2P�d\5-�^F:�ܻwt��)	� ����Y�h����'�S���@x��=l����{��I���/��!���/]q�a�B
���HSS�y/+�����x��
�u5<׋/�)'��ӧ	@}��Q{wo8���^2�����v1��`��r�EK$U݌��������%��`Q:�=#� `q�oϝ���R`�ޮ�OV�*������5�Gm�� ��X�^e%z�L�<�ƛ��=�-o�u�ܮ�2�e��K�<�kR�n���TL�A�"�ˁ��IOΓj>+�`B�#Z֫����y��劸f���m�Ȁ�-=���Q�4��H?1ci�-���)��@��c�@b)�f���S&`L!��I lP�ͲQrp�W��EA�v�)S�"k#.	� ���1ղ�u�i��3�s8:���*��F�)K�Y��{���d�d�H�������j�xc\�~J��g�P�ɳ[~��A`d�l� �w���l� �v��'��QxV���WVas<��@��\��ھ؈r  *1g�lq}?��4��p��{������I������{��Ȅ΢^�<��0'#�IH5}��a����0g��]��JЃ�xP��'�2���͜k�w`j?��p>̳��f>a�˚�aQ_[q�Y�g񥥰K���� ��/����U �=R�>�$��!�H>l<�&U}M�5K��^�ݰ�g��ott��,�b�� a+�Z̒�t�>v��X�]���e��Yp�����3��0�r�K��a����<�3����;?�	���C������X��`������4kS`�q�� n1��uB	��_[K�}�3e��̏���D2(�]H�1��M���}�./���}�+:�}�|��`O��av����iP��о�`���V��i�}��7��>�~\,!?��c�Z��F�}m�}�mɰ\��f榫2O�R��}m��D?��ͮ9ًV�ÌI!A4\���N:y>�{��;m�mX~� 	v�ۤ��J��t�n��|C�[w�~�����[�̖�x�`<��hȱ}_����<鵝���n¢ӹ\�,eN]�@�������v�D�b587C�{�Ҭ� �6��"����L&#Y�*!'8p(���ad�!�s��A�X�P[ԘJ���p��Շ�}87��ݺy�}�������I]r�c�z�:��wl���ޤ��D����Vk(8L#�� 6)���{Qj�:��R�� ��Ɓ񰼲Dfz��E���Yp
�u������:	0���9��y�)�o�������������{��R��S���@-�s�i�7=�C��=�<�qw��I:� ���7� +.��Z�;\#�������N����8C����J,`�{�lAx��kW�ݽ��;L�����:ח._vs��ٯ8@l�=�qp�q��(�41����(��L3�u��~�;�>��Cw(B? ��@��;y�sű�Y2�����/ �:�9j���9ֹ&���f`�˝g=t�#3y�S��n�B���5rdN�X�v�u�I��Cd�b^�=j�3�P�| _������v��#`9U ������HǍ�z��.�#�
kJ�X)�}a$@�$c0���
[�>�	~�>��Ց�K$�Ld����{T�Z�台��(�����%9�s�r����z͘�؃p��w�QzHƞ��.pt�	�֮�>���K����A�h��"Y�X��*w�tíTN��1��;xLS�_�]�����~by�[_�C:�"^_
L�8�*L���}q�*�������ND�$	�U�F�'���2ΰ� |žy,�\Y	�c �V�/��xJ s�/��2��kW������#����E��?�o���կ~�l}"�+�V/�(��ћ�X����������, UԆ���6��,�^{Hԁlկ�k�-�@����=�\&��5�u'h���������^�\���usH4�E��h~�>s����5a�D�L�����tW�\};e�6"Io��`�	�z�G��k�O��##¹�-/�=�`�رc\g�vֻ��q�;�/���׃ό����N{��f�������[������>r�}�3�~=".�j��s�f�_+K`���d#�Y��*!T�����$�(�J_e��}3��X���K�c�t�҆G!AݗY�ϥ*k��g�5�P�}��g����d�	�	��{�p�Tv�b�xa�뱛�����,��IZ��q������z1���Y���c.^��x?��\2�zD�&�oy�ٔ�\[+7����G�3�W� �O�v��-��1@�ػ�L�YV�F���&��E��A�Mw������g3����?�qc�t��b"��ʵM���A�Fcݵ�å���� ���F�V��֦~�Zp�D~�;ed��>˥��+W���t�W�xiL(a�C�s(ַk�n�j��
�$j���O0G�緶66���\	��}�6�o���nܸ�n\�q+K` ��p}����{��d�����E87v�j4F�LK�)��������{�M��M��1��t� �!��R�EfC�R���𕿑P�݅�y��\�>XƫL9M�$������:-�W_}���3����O�9��8��NY����A�!8#0j^	�:R�������"�Ǯ��De��>�2
�~|bZ�����^5Ȇǘ�MV0���@F������܋gθ_>�����*�f0Np�����q:��F�ϡ`�=x��-�,�3=}o�c�����/�~���I��p���BD����EԲm��_�2z^*v�D�Q��>�ȟ�4 ����EF��\ր�*͵��+�Y��>c;5S�%C���	@0]|d�����Ph�ژ�7яɁ�|�U�4I`%��h�p�x���/9ڮ���� �����0x1G�I�"�m���{��0�{�r���1�ט��1.@�
A9��������9P	 Z��)=�i�X�W�A�5qE�E���E�4u�˔��kN��D۔�O��B�&!����Iڶ(�y����u	H�1�{���3�w�&GH�N��x�|aXe�c�Y@���Q`U��R������^_7���C��HX���v<���h3�4�iO�,|֧N$��LE  �^x�}��R̭�P畽]F=Y�FͦY����X�,c`��g������-�Sa?��>��z�\�V�������~��d-��LS�>�P��۲w`��ı&�#������\��u�unC_I�zI�����=�V��;��@�K����Cw��U[O?>?D����0�Ϯ]��>���pmXk�����]٠��A����m���=?/Rr73�Fe�y	�ep�.?u����)
ؒ@!@�.Q.���p�~�zؗ1.`����=����iN{�~ۇ}z=���ݻ�Z1�l�op����ѩ?�~b�Mؼ��<Ƣg���4?�rn�X��+ٞ*�,>99.��<(�~�u&����Zlf�)ʭ��~�_�d�S���ˈ�`Y�U}�=:����j|V����8`�#�/>�M��A��5���y��O�kcH_�2x{����?J����K���§���烍�V�z��A� ��r�-
l>����Nۤ� �[n�Ae8�d�,<����U��Ԁ����;�=5��k?�����?����P�pIf�ر�0H9������NN3~'6e8�Z`��j�pp�`܊�K��`�;Q��M�����"�,ƫ:�0~ͱp	�$$R���`��3  ^�s&�`۝l�������������~p_
�ܻ� 8-�����oju�Ϝ9��Pguqq5�0�-�c����]�������.�ϱ���87U�`-X��|ঁ
H����Y�)����i]��1�\����5�G�A(f�y ��/]��gr��}��gϾB�0���1�Ɉ粴����;x�`_�-��2��˪]��fӊJ'xF:+�_���$3Mԋ�-�][���@	��7��3���c���7�&�i��]p8  ��6�e,��ma܀�<0��׉v��Q~��i��g��8?N�s�i=z�;|��	`uݛ��-�Bdə�y
'�С�T�X���G_���m�y�[s]�3g�R��
�)�3���k���,�씶����P�W��ew��ް6 T�vH�B�ޛ6.�mcӴ���|��;D�UI�W�o˒��)ca&ӿ���]�_�E��.*����+:N��|b<�5��U��q{l{JAK�y%`0�C;�Hq���R�1ߐƎR�i�3K��('���l�1�1�(��yJ�-�U�m�&Ʈ���I737��e0,�?����c�w��o�c��Ym�<6�h�D���(�/�=��]��OU���g�>������=��?ҡ�`���w c���x����,��3t��{
�a?D�ʒ��t�G��� �b�-c<Pf���^�Y�>���`��N����0^?��CG�pO��̋��l�6�	�f��W����_
���a,|ɱ�)5cb�`+�U�(8;3=�5�]dS H��At�tAF��)d-�o"�Z�Bߴ��Tȍ�E�L�A
�χ�p<�K�{���]�aطGF&f�0b�Gx��7jH|��״%tC��Q�ud�%f�h�`d�5[�}�*2%�cx�`.�.0�+:<� :�����cǃ�5�~{�K��G�:�3�c ��=��������_}-5N�@Vw�i@��;L�EAV�b��֮�Q�Pc�~�̐=O��t�y��6���u	T�6�k��b[��^�L��GБ����֒B%t✬D���"��mDו��'y��ˀ���F*����|ж�u������d���hOr�������u������?S ܯ[s��w��_�[����/b�T��ׂ�)��sR������Qԡw����S;���`�	���.���NMU���ng@~�.��T�w�m؞F�T�x��Ok�v��Y��M.U��Ι2l�(���|���9�aʬq����<��G��y.�����5���1�ZI
\�KHqܻg F"�ӌ�'�$�d�]�z�}��d #��E�H����ؔ{��w�_���{�G�_��A�C��7J:U !GG��]&͑�G���	^<t�?p�<)�a�)g`D_Ԃzxf�8Z��,<uC�N-������u���B�Z� ��l!�J��y�駟0�#��_�%2~�ӟ��������G���=�<6�'����&s�0N�\�3i���`1��U^���=L��ch��?@oȏ���&{M� A��H<)09?��Cw'<��G��3/R�A ���Ԣ��q���A?~�$� 8�H��S@��/��5���o�c��cH���@��|�����ݽ����_��RS��<7�&��;�=�����^��S�so4��=+��Q��j��/��㘝+:̶X
�9ɥ�������\jo��f*��V���
��9�ٻ��݌�v |���̹�c�,5����]�"��6�ۅ`a>"�/%+�����u�u�{ͻ�O93܀�e���t� ���\��3� �^)�45X鄱ɽH��L�����c	���{��j@��h�06�V�m�+��`4��7��c8w��eW�k{me�J	 ]��]�ϯ5��]Q��u�Dܣ�E�6��m��gS��������� �ų�U��4�#t�1N��P�R6��,�f�#xa<"�etd�{
����������)��@����T��0�Q��^�K�_��}s�73=C����5  ?|�0�0�V¾��(�e%�и�]a���3`RX�Q�&ѝn�O>���	>��ON�"���2��?y睰��q���z�c>vµ}������FV�z�5����5�3Ȳ��x��-�w+͸>u��������� ]f#`V�b5Y7c��1�F�g��Y�2������6�4 ���q3� ���/`|_�z��Ľ�wݭ۷(�P�z���ƍ�ԋ�q�jx��i?� ��G�E��b�ri�*��t����|��04a�[��}0���ӽӫ���-j;�W�~���*�4ػ�ʊ��`x�`�����Be�eK���W��>��VTq���u�����#��v�{�=�U��������Ǿ��.����h?�f��LҸ�7[bcb��O3x��c���Ƈvd1�� ��4�``�54E�R�U� %SA,�i  ��IDAT�2pTΏ�f��[rvv���;o����v���Zjn:A�웽[����3`� ��!J�ݻ����Y�3):7��zYe��!��6:�ԏ�l+_J�.�PeL0a����p�Q�@����}c8�RE�G�r��)����w��yw��+�I��½�p����
����总r��x�p�q���fc�����p�k�q��sgϾ�Μy�>z4�S8ހh��𫠆5���ڲbз;k�Jډ`Hk  Y��V�Zk��1��N�U �p�6� R`!}���#�pU��'X���˗	ݽw�,�ѱ���0��h����`6�T�� ��5yWR�1���B�:��	c ,���ݶ�y!?������#��+�����~G���#G��p�w��ᵁ��G�*�|��{��,��	�u����?q���8�s��/���
ؙ(x�	��l8�`p/.x]
2j���LE͊�?�H�.ԹK΁WVφ���'�P�m������!��^w��[*�8#)��ra�Y�����*Z+K,^��R�H�'�w�J�d|<� ���u�h`EM\��VH�ݒ�$���N�:��9�:����M0��̱�'Q!�-����1�z��,� �R���	o�*=W�*jA {���H�4��a�9]ӫڛe)lm��#�8�j|,j���,�(��yӃ�@�l���W΂��ZF��V3l6j�R���2-��,g��"h����
���S���vl@�>��rq�_�jsZ��e`�d<dkC������~��,پ,l���m�^���8�}$��{��'�O�/EC��k�! ��g���[8T�S�*���h���QQ�����R�L���vS���n<�`*c��"�ю�~�e�Z�dq_da/��������ȯP
B�/D�k�W��]d? cA�G��Q>���)~��Nٮ�����5,� �������Y��	>�޽SaL��$��Kt�h�#���0/���^A�t����?t_��4D�\��F*�e�e]� cG��^��@6�ԁ�Z�.� 0~�/q�^]Z�s�s�H��S����������\�c�����2$2����`�4���I�`3����/�e���5�-�2eґ5�x�1P�ݽ�q��aw��9�>
k� ;���7�C�U�����뿾U]$99�PĠoa�0�o/y�Z.��5��v�	aK
����%k\�{z]k�uھRc�y����H��Θ�O���D������|��8�A:�b�F}efs�9	��O,V ����|ڑ��n��7l�ųb[f,�q����<�ŋKRL�����{׼������_�q���,�ҿ�!m�㜉��耙�EMGԁ�7@v+ødP��Ԁ��1���f��ц�4p���`�4`�Z�YA�S����k�R�*F�+��>��`Ӵ�.f��M-ݶRⲛ�2�
..θK�pW._rwnO��Q7:,Lm���vMҡ3��Ͼ$�,�C���� ��h]�{Ϟ��ٳ�/��g���_qã�nyi.�zws%8A��IY&�
��K�l�ڰXQ	�d0���q<8ѫ��X�X0��Je �{�㡃��ɓ/�C���s���pͨ�q���EG��G�·�9r؝>�%2 2��_{�U|@5�```5��Y`�[:r��p:1v�\��1`A�c�����1Ov����"�Q�2.�U�cl����w�.Yֿ��o�>sc�γ����>�� �Ɛ�	y0���.i�=h�
��`e�7�x���(ױ� y*`���4Son���H)�c�+�(�/m�4�V9dAl��)�~�h���f�o�q�uG!�S��k�9�eV�S[�,�A���Iگ�;ݺ�Ab�������5&�R��ׂ}#�JZ���;J��y�t-��^�<	�́RehV� dh����Q�Tm�Kf�!�]4��]N����N�r��ʮۯ;�VR���Gl����>1� خ,���) XIp� �p
�0��*�;/4�+l=D��ꈎlop9P�ZAbu�$m�qm�����(��̻����Z;�=�"ĭ��n���OK:y.{}�E�ћ�]�ٟgπ`���ɉ�E��	��%X��u�q�h(Ym˾�k��u�#�)%��1��Z� b./��
`�O)lx�`�F�"��,%m
	~�nO���{�`d1��̠�\���*�8�)�� 嵰�A�	{ M����;��wZM��\��`[2�P�vzz�s�M�&)` Y?؃�} ��+�F3`2�k1u�tfRfӵk7����U����	�ʘ3���8@���s���{d�rX��O��Ν���3ee���G'�R2�|�k5��b�RT���&&����lH�@��0��t̠�~A�^F�M��9���o��X&��8g[��� ���ۿqG�BȌ:�;d�rP&��K ���l\;�k ���L	���{T��Q�YQt�ϳf��k��ͫ�O�k.����)�k��}��iX�K�_��b�qmM�f9������z6_�~L�ד��O����=��O����5~��s*�Y�/�b7��tBd	��=���;�ZZ���׽5.��8�{�t�mXޤن�lJWA��� $#����oc�쀖��ֽ�� �϶=&a��|_�:
����J@�ĔH�7�B��-��Đ�Sc��@�nX'�Ee|�l�hp�H�hi�uk�����S��Ʈs�ں�B��[pࠌ��h��<Y�tF�_��5�,28�pR���С���o/������ Y�����@`�=��{������gnϞ	��tR���$M}��ڦ:�H�5G`�8e�D�x� ��-�9���I8�x����U;�"�
�A<3��ᳯ��;}�4Sq�y�4��3]���Y��8�c� >���苑���ك�+·{���Gn�:17f��j� �dkWp�Y��V���ϟw{�qQ, &��D��l��2������cH_ܹs��˿�+����N�v�Zx���Z0��MM��<)�{��)�����8�w�`���x�#�=���s���@�� �){�d�n�f�H @�%�,	���2�4֙�n���k�ǀ��C#�@ٖN�-(�3�r06��yE��E��k��������v���9L���_�HT�ty��ed���5ڊ-���b�`a�P�[ٰ)���(s�c戓b+G�`�!��d�L�,���u	� D�W�!�A>���׼�Ce��5��5E��S�xT�,0�� �a���Y��=c`i[�}��p��٣�V
L$�$SP'e|H�@!K{�/Ȋ��y �r~�2���� 3}ʌ��^���G�s�e�Rs���0}t~$����L����2X����k�$�����.I�AF��/�<��^dgVeoT�DR���̂}�>�a΄��Ã]�lX�Nﲕj�;���+���K)(�����0�P�1'�Qvz��� ��%�?���=X�&v�
{K�2U'N�lƷ/�_����⸏����~�Q��`n!�ɫ/þ����G�2>��F�F�0�����}��'��B&�1�m���a�������i�bQ���سܵ�r���#�z�|iQS�%�m�ӕ��+�D}�`
��)�e � �a��}Y�%[�4 \�t����F�xtA'.�2�{���:��A^	�?�v�܅l�5�K��],
����U�:� �G�@[�k�L��|/{2�$	"�b�P��u�����s��A�eE��� �x��J��֋*�+�v�V�G��i�eg;�i�C�59��O���H��,��X�2+J�#[hj�:!��HN�V���Ș���ܹ#�>���Y"���C����py��,o��f綢n�8��L��^6sc��0� ��z��<��[����.Lb�W\}CɌ���)�&�ve6�k,�,������Խ�eboU>��:�;d�u"�v�.^t�"�QP��}MaK7
�aBki�p�\��gl�_H�ã�%w���u�^XK2h�L�M��̲��v1X3�+i��(�T�jGn���7E�䳯�u/�y�88�s%8��d��dI_����v����t� ���~�"7 ȪR@�:x%���؎i���� l �c�0��Y�Y>�|px'vMP�XP��xo�Uw�������g���� �9�o�^�Jw;8�؀�� 0�)�����`3���TFG0�~p��\�~��i��U �hW�bA�=�7 ����ӧ���(��#�XkwܩS/p��� @����"��
���x���
�I8g�vi�ϧn���T�1i~Sd;��T�̟"P	��~l7��͌B�(�f���?�PE9�O#N�k�iiɀ���X;�D��[��]q,�Už�d������leq�Mv!�O�U��,�k�i�1��2��W$f�=����s���ښ��/<Z�6*֓%jǶ�j�
� �LZ��v��=+`(���i8du �O��g��k�7���ut�QI��u��UJ`����Ӣ��o�U�V�Tnh�}fbSu��O��]�+K���˒s4���RKt�1fL3<�o~/�׆��N�^_��ͺ�$0p��j�'��R���)����|�)�B ̅���w��M�����5c���X�;^��!����D�RG�9wt銻y�f|~&�ϡ@33M�+f6�IԬ���r7���w��p��yw�o��a�B
leuY�<1��B��ZB�	k��J�B���Խ�#��歛܏�;�c`�B=�[�� &U�L�����E��T٨	�Ã�3��鰠�͛c��k�o )�nWd�޹s�}��y2�1�К��$}l����q@j�: zB���,,�!�x���q��E��zǀ��D?��6Ԇ�
����!9��D`�f�m"������-� �W_}�:ĺ�k��aچ�I�(d�6��������㌋1T�kc�{~Uimp]�j���O��t��1�+ ]�qSVE*\�t����K��������E�f�-o�x<�ƽ�.�z�7Y�k'��`�A��י���Z`77}��f�w?���&��e�x�p#{>��|�p���u�t��cϱ�������P�C�5��vZj;��--Ψ$F��Gs�a�$0èfj�S���v։�]��,�~.w�j���S{��[��,�>��SIaw�!�Q&b��3è,]t,� S�4n �1��j�%��U4Iɺ��KeM8�,��R7d �:$ A8���(3фn8��m�%�\toe��}��ݾ~�ݹ5CI�<���37?�ng�����LE!���ݔ�`q��Y��NM�w��=�^}�%w��Wݾ���E����\0:�9�K��޽�����������k(8�b~SS�������U0k�3<4\��Z[Y���ֈV�o�Y8��ÇQ+[���Y���o��أ�������A�ᙙi:O`�ʦ��7M�i������_~�R8
��)�>�TUci��$ ��C�&$u,�e)r&r��Xx�2�`dY�3��`�!����k�22¾<xp�{��7Y�� �N>����9J{�A�=�;8���8�pK�e:��0|gj�~^/�e��П`f8x�����=��)w |@>X�Zy��#.�Ӕ��"r��ԩb�9���9[>���-�G��ُ�bL%s����"� ���]	jg���/�u�H���-���1 �	�0-h�����k=F=����O�q� ��T��z��Z�$r R��/$YZ�e�Z����tlYe�2=�a�c������N�mL���٠��t�鸵G�%U�#29N�ft2�)��W@���n��J A!)���g��.Ճ�pU��T�����
(���l��ظ��/-f �~��8<lr1�g�r�^��<�����k/�n���&[��pD=T�g(�4_s�������R�-����I�.�/����!w�ԋ�:�裏ݯ�k�I��P�&wa'���HP�����"��n�va�Z{�	�(p������\yl|��5��˼�b�'0չXp����B�Y�vP�T\��;��X�������w��mJR����}{	nR��;�Ej)c�\mj�?f�,�Q��^�"*~[T}X�.�h?ص�m$�|_�.���ؘ���t����hŬ�vgՍ���)-���gU+zA���1��XKΊ]Z�B�ao�裏�έ[�qdA��@�BH�!���jD�G_c�ؿ�s<;ꅭ78����5�_����k͂��k�vj|L[��V���y�A78�"H���d�g߉k���{G�s��!�y@�	��l	�،`�+�K
F�ucDV\S|m�X�9��{.'�,���M_��ۭ�'@�>7�G+���r��)�7���~�`r�L=��u���g֜ټ���_����tl�ͅv�e-\�$����}V�`|�)�NZ�X���"[�v@��,oؒъ�:@�ٹY���"D�Ӎ��ت�����Σ���M���|���R�Y+��������;:�c�K�u��
�E� �#���rZ�a�Ы���� ���+;�4�����N!* Ql�&��A&���pO:9pzT@��{��[o��N�p�,�/>�,��3����ľa%;���|��7��~��;v�@plF�q-�f����W����ݹoλ����2��[���C����npx��2 aaӇCI��p�`QNu!����
��e��tZ��	@�`TZMx�)�xp��������{F�-�D`耝Ô��4��g��������pm�Ǐ�y�� �p|�+��kƂg�y2��x�`���<q"<WIG/ nϔ�1��E'�8�흷�r7���q� =y�$��pvV��𽹇 ����ay���G(R��`��������;��0ΐf�����|�fm���r�@_�wѐO�'��o[C���s�1�d�(GP�۰�U[�y�JL�+1���l�{����Z��nE��ə��3g���5��2��\��`��6aኮ�i��hU�ʌ���D ��>���H��S6�"6���/�����z_{�Y 22��8�5�5{|[��b��4,�kh#���o'�Ttslp,	���A���<2���5��̾F�MeuD���@0������ֲ��X(.��n݀'�i��)�=7�X��63��,���Z�o:Op�^e/�H6�{��`�O잺 �g�z1��&d�1�>5�z���Q;@=����;�~����{*�"���w�9�Q ��#��u�g�u\�6~w�N�s�q|����:�K8��,"�G`��m��@����75�ڈ�2f�@8�u�U���ފ�Zɰ Ȃ���@�,���+Z��D9���i0C#�j�h� �5����B [X�U�&ɺ* ���,� >��O@��+�$4p�QJ��&�� )	v;�U����,���Y~ i��|�{c�@�8$S���C;�/�k����C �����O>�y���YRo���7���!	�p�AVG��Ң�@�He�u���ɡAX�"��*e #��(����	�Z��!VkSt��	]��T�3�����jE������S�c��m��T��۳�=�w��z�A7�C��^�p] �Y˽^�������z��'��ռǜf�U�[t��IRPGjG�1�����/\�Vy���_��׵��h�%t����tl�d������QK�nfFD�M�Q�x�~��L��4��W{xO��7[���`��d�P�Th��$�*Mi�/�SX��4@���s���B���)����3V}��c�x_�ư|���D�6p2��	� ��(��l4c�����3���V���*�X��v��yw�δ;r����~��)���?tp*G��_PP����Wθ��~ͽ��Knl$+�C>߬P�p��wf�3zU�Ϲ�W�+�2�������ԓ'O�&�sp�:��XP��(�3�d��F���(x�5���l@�:@��Đ�`%NVW����cN�'B�.@c8�p���x��`8l��w�>�>��Q�~%<o���a�,��jj�H�f|iG5�}HO��v��Ѐ�a���6�Rt����9|�0�׵p}H�-�0��$���%I����18\p|q� ��E�q9��+�d���u\��j�մ���6��Re�dL��I��R������T�t��Ud���o�a����\�~�u_�� �^Kt��l-J�������kα�Z���J�e+Z&�b=�,Vg-m�0��rxn �Y�!��u���[�S����G��Ƽ�tm�9���r�� �0?P�s���#����� ��~�u��^g���m�����L��3��ߡ�,;���c_��s�M�|�ֺh_�Q�t��j-��V,�,S?�c��,BI���W�+`��U�?�g8�=��| $���a�.��Hty&�#kϣ�i�ZM���5�.ӿec��ؘv��RڡC	6��`�\�>[�>�P�"��6��~A���1�k�5�m��J��:�N�>�^x��- ];�$`��AK\)@(�{���������y_�=��~�!��أ?��sw��9����T��(P��)k��9� ��0���\r��F6q�O\��]��9����pG��F�O���}��t��ҿI�B�厂ڢ3���R�Ru�9���P`��B��u�k�LA���kRe&S���s䠛>�F)T�Y&��-�����G��Ѐ�� ��~�d#�� |YdYY��sOh�@'@�յ��Hx�l<�1F�`�а�Q�2�p-�U5��2��հ.k�����,����������%���ޫ���*�������P��JE	�J��zcJᣔ��X?��@����Kl,�(v�����_���h���/�H~��*���펲��E�_�3k�|�L���v�E���~���a�l;�� �=ZnAY�y�,���g�tP24(E����;��Ҋ�h
7�2�>�^s�3_��amI߃�͒��N��=��~�M���s��9����}��T��;u*=6�Nd�b�]*��� L�r��tG+�������[���.���d^J������J�X��
*v��C7�ժ/�~�J7�е���"p�Yss�.�/>�"8&������r�_<�v�"+���,�3��p/`�B�]:7���ř3������;x�@��Uw�u���w
�H��;����>������ͮ�g��1��Ǘ.]��������n�}��Ȍ�EC`y@�0��ܾG'l��^�pQX	�{aa���p�`|�>X!��Ba8/�g`�I��N���O��?p�/]!C)Đ� �r)8u�O�"���3/�� k27���5�D�� ����Bj,H���[�?��}( >R~�
������l�(�1?�� �;~4|�����O<�t�;q���z���P�������:)�f� �m���t�5  �4�tǎ�r7�3)�q���:�����1
/?X��4\9�C�S�+J��z�T�U�%C���^k\��D&`��\���b�.w�@��K���q�p�t�rR�Ԃ`,kQ4�	~�kƚ��jY��������A�f��l>9�<�"��ڼH�H���!H���B�1��hDy��Z�9��V�97G�.R�-��
�ʸ�n�$?t�M�H��3�\��W��\�^���{�����?�w��Y�y��΋k X����o衂��QAG �޲eR0k=�%4�Q�ϛ a�Ɓ�� 看{LU�7���o ��,mr��� �P�kҸ�5tں �o!�{f�;�)uɑ�+�oM�����Y��=DMU}�[.4pI�k�K��I[�3���Iޠ��ǳD��dm�"p��/�Z Ȇ�c@{~ ��������x�ݻ7�Y���Y���������ko�W^=�9���-�l=�x�^��_�>��w��m�,h�h5�Z�������8BP?V� {��Bu�m��\hPv,ʋ}��1 � ��Y�iC��1�N�'n<�o����sImo�����.@���a>�e��ZS�E��J^��wɚ�TI H�����("�gr�� �豣�� �93B� �`�����/�m�S0��]� ����_��۳{�Ah���^I6l��`�t����e|tB��3�y���sF?q�?�WHb�L��h���Ŧ�q�����(�#�0��Q�`9����#*m�\��1[�����ѷ�Ml�~�e�;�����}_��_o�l����n�um�@���mE�'��+s*w:�-��ed���f7c?��"�]{<k�$_�Gd9Jy÷v:mX^�����t'8�؀�E$Y�^D�O�|JojpB�E��P�_�H��n�D�ٵ�Bi��;{����z3�:�ڐ����{��+�Q��yo`��2@��f�JL��EP�`���㰷a,���]��(�d)�	�b��+�W���l�:z��Cw@%
X4�Z��[�q_�>������	 ��idt�=|0��������S&� ��VR3=ŷ�~˽���n���޻w<�{��u��=�����kw������<7 ��.�� J |"�����#��y�'���$~�)q2�m5;��԰�:©�c��SH�1�W"��@f����B�D�|&�p\�q�լ�{8Gg��`��@A��j:㼇b�B����������@de(���P���^D�U�ŋ��#��k45�J)N؉��p���po`d�� �"![��"��u붛����o'v��s�)�w��!2����qc8���1m�
��
�D�G�ji��|���J�9��ͦx�T�l��"e��S�q�j`' O��RyY�)!��u�����|�J�d��\XUdP�
��T���c[�����h♈����h+�,"[A���{�o��<1`&�V��܄a�]��3�ϯ ��hT�3;��d���]�w��+��*��<Hj�OϪ�sw�M�so�a��ڳi@ v'X���x^��o r���T�-�5�T�<���}8N�#�2��h�RX�����YH��إRL���lM���-��r��0�:Flޛ�G�ǩ{ҚP��.�lx_��(��:��Đ�N突��SEʢ�+��T�����=.Tf��,p$��- �گ*q�9]v
3�����`�k~��p�._�,ӝ�w��^c32v��c������o�ӼE�Y����߂Ō�	>U�������{`���u׌�M�ײ&�2ek�T�b��ܛv3����a�m��-�سy�	��!\;���1T���G�L����T�����������`-��v� �Y5k�p��3׮^c�ߓ'O��qN�>� ��_�� 1��M����]E&x��hJ�i����ừj���+�GK0������=z��uGd?�O�	6�Ң[�g�Ͼ����`�ti߫|쓚K����!�7��J�U�[��}����t?]�Qm=��w��~�:`A;�7Xh���e�s��R��~��� A�Ϧ=�@Ï�e�$�jݧL��8��sc]0�O�=PV��@&5?��%�T��ry!O�߸���˽FX��0��:�h�Qt0�0�`�ᴣ���&���:q)��NC�*�v�f�����������}��[��G�o��� ������{n*���U�M�<唆��-�*�ϭDZ��c@��U��l'�Ǝ�p��/ڙ��*���=�f �"M`��'���]KG��i������8F������·߸��{�͹�t���Cg�Nep q��I��믹_|18@��,�A���^�/���}��[����@)�a�oIj+��IY[#��`���_�����򒤣*�F��=�I*���	z���(Rb�h(�TEp"��8�m���(c=9|��k�*ߺu�U��3�N����Dk'&�C*,�'�qPA��2zP$��P�)�($�׋�r��]�+�%��-�B���"��� ���(�6��~8�0��Ȇne{��̸O<��a����G�4��Ɉ�}jx"���R�(�	v�O [�X�7�ҲI�+�V�&�́�s���m�y�F?՗d�e���"b/�0��R;>2� w.֦��LKg�H�(�d ˵T.�k4��5J a$a�3}�!�D�wv�F���y�R��7��T���xAqa@�ݙ�`���UJ8�@�I5@������U�}|R�z��x�'�ٷ�M��?86��ʤf2	~�s.cM
4�e�,N���	���C�S���k}r�s�1�����1��D����.X\T�ye@�U�w�>���z�_�k��.�>���e��2g���UDS���d�����;&ȕq���JY%(�Z��l���'�����Q燽.�-l�R���-��x�/X��,X��i��˯��7o�6���qDz)�����h*��h���m�a�!g�A�%��U�ϩ��+�k�
׈٭�a^=vÛ�M�����S��42`	�*��m�f�2���\Aa��/�e����;��1J�F�'jB�8��${�� {�rcm��<<�8*���m�K)m�h��B��+<ǿa�H!���?-�-��`� � [�+а��A�4�	���jj���e����X�+e��m�w/��oź��K�.� �W�c�|�ꗣ���<�\���{Ǻe�߰_��W&=SRj�z�|nI�F���\�J�gt�3C���	1C0��������9�\l��'�0��j�뺸��bŰ����{'[���n[ƕ�@?&<\=�;�ۏ�_�@���y�6g�]�����qf������Bd1Y�Ovkpp`�G�K�0Ni��1����X�G믛�J���>t�<p�s�4��h�a�Tv�sy�M�:�q�ËZQ�&դJ�������w��W$i��46���5����[o=������ �=W��y/�\,�k�TE���U��^v�	�X8϶%	�܂Uܹƾ����Nt��4ܳgS�Y��s%O���:�"���.�p�\���L�d�LM�
�����w����T`���Ȣ� ��:q���/��,g �w��b���S{�.
&$6>��w��MYܨli��@�����y��B���\�������nhp880�V �@���(z)�f(ܸq�ݺu�������޽{ݭ۷�`�;�G8�hH��^!t��?}oI��>���]���#��3�����7=MP�;�[j�=�
����ϐcLe8���I6�ʪ�7 ��_î1Ԡ��s/�,������[��4�c]YY#��
�ɂ��b� {,8��ޛ7o��f��a:�`���ࡃdl�`b#=��SS�����d���B���=:NR�6�` �����%�N�R��n*��X"��T92�|�sP���IԵ����}�3��6�#�ln�c.@_��0ٓ��R�1G�+0�i�*5��
K5U���)��+��.sP�c�v�h���O	H�E޶���d7�WZd�7� :�/�����R �����Y�.Ő���Hm9J��n(� hRlט�[el}�  ��$0*E�PU�S�7�/n��r{�C9��X� .�~��)a�e��(�	8-8W;�VX#�Xa<M��9�,�1*�alb��A#2NJ��E���p�Op9T"N�gf�}�>$��Q$�Ut9�"�@�zp�J�"1�+���̦��Y����{2�@`����T����1}��x������uU����NP�^��w�X�0��M�k��% I���ەm�Lr��Ew��5�1X��R��	`ڔ�8�=�A)��[i�2C����--��$�4��@O�W�?}�Y� �I�6�V��T��B��c�~��,
ZG%�,K�3&�����������=RQk���5�hD-{4��/�A� H�>|���ezf�R@��"�xM
�-/�����n'-M��>��"� �z�f00����'��\�퍵zr��@<�ʔ�������+���;�������x,����<\��S��Pǎ�y�N�J-#�$t����o�rY�<�X����Q1s@��K&`y���l�$�k�ƶ��Y��"PV�噂J��m�>��O�U��a� W�y�����'h�m	\�5������b��f�}ʬ��smL���`�l3�#��e;��{��y-Dl�nUi؂O�{N�s
,�n�DnS�	=��y����������8�h���aQ��U���տ�;��z���߫md��~����1���o�49{����G��g�Fڀ,ͯT��w1�k���H�][�W�Iq(m>�����&��_�<�ۨs� |x����O	�������I����Ν;���u��<Txo4��-lߗ_:�^}��0�s4;��`c�ݺy�]�|!8�Wɤ�<��(��N'@a_����x9R{��ڷ����~�N�>M�YXs�V*�Ja��n�9��"	06>��a��m���\��s��=��'��ad{n>:��O� ��ŗ_�9B���e��;�!��X|8c7�ik�j�(�2�;t$WU��M=�E�%�'�3{�چ#�t��@�1�����O�?���C��#�w����XN���u��f���nab��� �����A0�4�{���޷w���|2�L0$JtHfϗ0�Z9�iP�er�ztߤ�^c�,K��Z�;@��l44u�(���(t_x~�4���|3=gHU�8L!�?(�&�V�γ�����e���\|D�b9I`>�߾v�G�^��i0�D����Q��^ˮ3ʑ��mm��y�����l0�}�haQפ�W�+3X���gXR����,�M��~De���"p��>�Yd���� %۫�J�5b$��J������K�T)D��*?Z�^��Ո|�k�ƌ��פ0�>�t^(�/�����tn���% \f��L�3���*j��\L�al���2Y] �N���	�Oٛ�ޟ<u�-�qp'����#w+��`�0�����	�	ǈ۸��Y�������Q�%-�c�XkΪk�� ��mG�J�)�f���Z��·Re��B���5�Q�) *�]|?��$۫Ǯȏɽ���Qd��0�2omͪT$�'�zbIc���[�3?��e!�����i����k��� sK��a�!��Fp��p��3������g����ڰepod�Sb���#�a#����n;z���ڿ�sN���[Y��-ۏ`��:�FP�
��������l6���z"o�}��LG^?��]��_I�C	NU�;�^��[J%^^�z��>�L��Z���l�	�}���#g�p��'��v��-/��zN����ٸGW�f3�zhCzk8��SԓR�� ^��u]{�e1v�e6r�6[T�}������%}�%�Se�r�����棫=hBɅ����b�Q3��Җ���,�@��<�7n	��*0���nz�^F����~m��^H��K����҆�k��wь)��fR��9[e�O)� ���Fݮݻ���f��[�ͽ���V������(Q�����+:��d�b�}��F;l)���{����xýz��	�d�@MMM����>�#���!;�K��a�]Y��:�Ϣ��c�	[���ϟ�@gqxt�<t����"8��2�� `�gx�7�� ��AwO��cZ�pT���`Y2�Z�~���z�*�S| 1׻w�H��<�گ�%���c%p�p_����ݩS�L����,�Q������-SC��8V�_i����Rȏl�|�561N�g�Zϫ�_�R����a��/����?������I��`�T�����<�39,r$�ll��pZO�>��):��?��ݹ}�M���:��-�V�L�BS��y'�c#:{�����C���՞����O��on��<�JAf�a�RZ{�|��0,k��J]ʅ�BA冦,�v���Z�Xp�ي�d82x&�N<vCdɦI�f]V)��'	�ΫIv��nIӾRF�"Ae�Hi�eNL>C��*v�o��E�7�Y_nڶ8z|������&�  ���2�@!����p��h��^E���FG��ێ����HM�-W���h?F0�sa��(a���� 3d���&u� [e�r��"W�ه�1��<��gך�ֹ���Ϭ����7}��\i����xdz]A_�㞷Ԍ-�1$%><g@9�idޠ������{���g"<��N " hrKԐDp �_�%�ۖ��~��TI>K!p�Y����|�l�[���}�TbLJ�N)J\��B#�[-��"`��@>cm-Ʌy-r�J�Rf�U�k��YVR�ϲ�����4����8.�kdt��`�%��0W���t/�F��?�G���[��S0� �1��X�G�ad�M4��� P+��c���{���2�X�@��.�,��#G�J�>\/�J&-������t��(�����(��j	3{`h0J�Q>�SF06	MdA�<w�|��'���eZ��"Q;N׫6�{��x��w׏���`_������WT�ìT�g38�qז����r����{���e{�>|~p�ޡ��X9��zsb�2� �/{˒(�������g֞#`��yu�.��*�g�CT(�m�Y��E|Y��K�������̰4G����* �lrW�1`��RGo,?��}�m��ܿ�����Y3��E�~y���~�4)Ru���H:5qƓ�\��)�3oz=6�#�C�|3~S�r�Tڅ�1c�t�a��S3[�AZ�z��~~������ٰ�߿�M������M�������x�� �R���5��ӱ䦦v��^{ս����N���G�C�RF!3�k��Ш۳{/� ��V�׆�Ω�!:^~�kv�}��s�ϓ�5�o�;��������2�9��<�C#d�3Etmm%j�¡��g`u��+���7�|8> ���G_|�u?��Oip<xp?8���sTP�ɻ?q�~�;��� �!����������,v��B��,N��jp@5�3��J�AbH����:���pm�Z`P^@���WhO��!M`��#G�Xb�C���Ȑۻg�q���>x8�@�6�Z��^��߸I�7��N��s���p@�p{��#`'�X�E�dP������ĳl���=�D.?�;�3�c�<��u���^�7r`� ��9o��
�V��yq�-@��>�U2�۹��T�V�FL�v��<8�뛰Ç� ��s��z�����vS�k�9Pr0��"�ͮU4I�o�me�staAƵ����h�׽=c�X�R0IX�Į�:;���Zl�>�c��Φ ���i:��E����c������tJU����� ���5]�?4��s3p�$^�� C�9cc�ȞP���묮�1���M��I�&Y@5������5���-#�Rb�Z�k�U�[z��g7&b�I�:�=�ň��̜�l�ݻ]�^u��&�/~�s��`�޼uC�� ��
$1�����X׉7Z���]c���d&�u�֯w1�-s��z��{�$_�X́��xN���ˣ#�|c�>�7��Sg��� 4�*�7���8&v�1����,eHI����W\'��
��v��jrD��8�'.]������������߻�������Cw��Aw��fB�a��>� �Q4ϲ�@�&R#���5c��]~W/�^��{��Mg�)oz�f8�Z��}��Kk���Y�� ���5an��D��b�Q�̤�j?1�������r`8��f��-l��1�C�f��n��'9��.���(\?	���x�}[�E{��~x~��~���w�+o���Ӈ�W�[A�M���ر�-�Y�=ض����䞽��M#aO)���z��9��7�`��X ��	m�s�b�-Ou�5˪r�?_g�M��w�O��ߤ�c��ڷy4l[9S�w��7���mu{��~+~��~�IY$22�}}Iiy��Z��t>Tj���m�1���6(��L$���X��V��m:R`�U�	O�6���?8�ss����?���Q������76:�4��-L�^ ��t`�~�ҙ�@H!.I�5��~��1� �
�\��^�Boma�DP���|�b_je�NGX?4�>" mh-�X��
��� �p_-^ރ� @�7� A{Z�W�^����|���nb|�{����t�W�	�>t��4�,�~�#	y��^$��ĉ�n��)��o`�"gpHy� ^���Q�QsV��b�SA ����i������d7Ag����,�����FM�۷nqyc B��,p�,�� D�b=�h,���X���'x�gY<\# �Gd7yS�� ��k�����zJ�����[�޶�l����a��}ߵ��:���JD�#Ȓ;�])��J4�f��ɛ���߀�B�L�A�V.>}֛�ki]����@��)���9�]�/7�-=��翤�0Y�"�M�!:zm�PV�aP��/⺮�����̵�R�zy�f���r�Ռ
�X��?:&�DUP���V:(.^c���W�}!�G��m)c���4�����^��h,�TE+b<���k�n2-�Vs��d}��Ъ�4|���cVw`���˾������'�B�Ik�eL����ݯ?���]}�w{~N�ms*�`]G$}��j�A(�57@��W^����;���n�-$50� X�����fфqv�,�gr\��FiG
}���c]2��z��,�ޒ��Fd�a��A1%>¿��� ��6��d+[�c)87\A{޳7��1����d8(Eb�RZ���g탑����+���������_���~��ݻ��'X�M��o�~�hۑ��aqq9��5ޏɆE�SX4[��Fmɀ0�p����x�J�����,�kz���++��o3�E[L2֐�$�s�w��#�*��\fLߔem|f{\׃by�k�u�!�<b���L�6 �����9�fl���&�R���q�����K� δ����h����1�����-�<��r������6���*�RGe��m{W�26�ƍ�Q�c����=�������u3�g����1:��Ȃ��x�G�v��M���8���U�Z���c$�nm�>'r�]�t��s��7f�<�S˯M�m\����љ�H��1���}����Z��D���LP�e��X� A�V��%�P��{�R�t�JRZ�_�B`��[nl|�N$'^{��i`���z��.: ��	x��q� �]*~~�ݸy��?��|�M�K~��W��o�Q�Q�_�Ȳ4ǣ+ꎆ�������Ƈӈb|�|������fk@���Rp�ׂS���R��T0����q���|�
��9D8H�/_����믹W����7����GJ`���$��?��s`�w��u^����ܻ��N�|����"��"o,ҷd�?�L��,x���Z�,��,�r�	8���ݙr��\�wͅ2�+��mՆ�>�M���G��2S[�ktr1�x������?u�=��c�1��> ���_��9I��oΝ#��l$���Tz��3HA�O7� ��7�穴�}��x���]���fHM�3�.W�B�@7��O"�QD`&O�/��W�R�7�m���j����z�M�V�����g#�=�)�5PY�F�
ٴ�Q[9g*[���¸B�,W����زݳ�t����2���W�=?�*'6��O���l�G�i�m�/E`}F@�I5k�@�!s��t��8���Xe��׭����= ���g.������>���z�p�q
�������T�����G��<r �S��w�?���NgQٞ�.��'�mHn�lR���͜V�i��8,�Y�׺�~^�?R�na~���С��TGP�wP�O)�)]{��þ~3�KpACV�N2��z��T|q; "�f��#�g��3�o� z��b]���se��q>�i��E�����{"
���k/�]��Pfˤw�xP�dK�$``��rL�oG�5�`a��|�k8�I�ؿ9/��V鱐m �/�ؿ��o	ʢ�/���x�u2�!�17?Kk$�`/S�bdT��d9�|n��Z�8��Jy�>�Sh�cE���2���l�p�kJf颒�Jl�#C.���-�C�0�����}0��H������ͅs�/�[�L9f�Z�ȿu�s&w��gUe�O��%���,�, A�kA�$��6���>���}��e��V~?/�(����0��5#'���˚�g�-e���jWgx��>��r�(����Mz�4Z��9؊���k��:˥DB�:T�s6h�ڢf�� Y�O��h��v��W�sW�[ �{�4���y��I��V��=�{ɓ40$�b�!.�<�F���jۖ��7+sb�vu>Y���π"4�vZ�ڡ�O'�bj&|�~�J��y��F�� F��r���������ǎ����P	��؏?�08=kn|t���r��VpPO�C���A�,�=誒�P2���(k�r�v�"o^V������W�ݧ�=V� 3 �������[oF���'%�	�LH���/�{��� ̒��	Z\[t���!7Y�������nWp�����.�y:^p�'w�r�t������`/?Ϣ`V�{����������kw����7_�Ͽ���3 ��pF�#��q�k�7�:H`���<Dp!����7����˔��`FRq��'vOp<C�� �(?4�>��ݻ���"�[�����	��,�q՞F�!<�C���#�� *~���t�1&2�>f)�,�� 6���J[,��j�Eqn:�p��[��u(��}2�ʥ ��(�ftV���T��%�P)H���[>��Ơ��6�IN�8��V[y��Y�ge@��lk�4 D�� �F�vD�"�᳋ˋ
hh17��ŭB�x��Ф���@'c�e&��މd-u�#b���c��=���m͙���Z���������W�J;�z�K,0=I�w�D��)c;��:&���
ɛG�dD⹋^�J�UVl,1�Enw�Q��kO8/5cU��:a���,�d	�\�n_ �y�D�|0[r�ؾ���.�ًSGd�`Zш�����`OD�z?��>���m?Y��CQ�M�I����Q��k�.�}j����^]$�2�l����WϺw�y˝;w�lw|c��=q�sw���k�V��#y��G���P���t��7�-��Y�eܣ�;��Y��NSz���H���v�|@0����p�Mas��?��fS�"\���� -��}�R-�� X�5���Ȇ*�A�L�e�������xݝ<q��<��w�=�LO�={&9�h�x=�L�5�z���h[���ܢ��c��ϊ�f�}��6��Ҁ���峐^�>kw��M����t��[-֜H��7��&�	�2�`G.�.Q��z��o�b��<�'�q�۰^m���7ܺ��Y�F^~�N�'d٦񌃐;m��o���C�Rv��7�mEBꜳZ������V��yY�[`̚�`ܟ�a�C g&[���c$U)O�T/s���=�GP�;(7��z���ٖG�%�f��o +�2���ʭ*s��_zzΙ��/�~�z���骮\���Ď �}sw3�WDT�<HlA��ዙ����ȕ+WF �������˿^�=j3�N۫hi>���o��X�ZXuz����hx�s�����M1z��L*@ �nL��
S�����E�}�kW�>2�|pd��/o~��򗿺ɉ���~�>��jp"v��X���=���#�)XIN ���)j5���`��8��(�`�X��2W޹�a��Ă��5B��;��.vxa��]d� ������3�/�U��4	Ps.=��P��/n�O?��������@a2�W썹I?�����͛�֭�y.\$�fXW ��|������c&8����n��y�=��(U��l���~�4x)`J�B~;;�k>s�,��=Jj���Rx]�CS��<����H�h=���JI�;Hi�a������w)]r�T���3o ß>y*l��i�`���H�H����tc��� �lp�Z����p�?`�
���O	X5�}�X�Zk��>>���(A�05��>6�8�I2��sp@�d|���c茠��/�cϳH`H�t<n�ɟ��eY�d��",n��p����^��aѺ%i�ؓ`��9����u��O[wr���m籁<b����C�n�u��c�"��'23x�$-_�J �����Ȟ+�e�Vx{�N�񢨵�=G^��A%@C��0%��.li�{Sé-l�&���Q`Xn� ��s|k�M6-�S�%PS���?#��oۉ��`�Rg,Ǣف����=�o�����};�p�A�bs�SJ�a���g?m3�u| ��: ?���?K���°�X�)o���F�E8�%P|���݇�`��-#K"�� �=��`v�������t�D`�\����{��<Y�h_�W�G� :��R<�S��V�]�g�$0^ ���f��YE�Z�sP�	�x�6�h�{`w��-����\�B���6��8Vx֐f�3�O��:`sȵ%��Q೩S�(�[8�t�5�����F�kdPXe8�9i�hTO�18�d8	`�����z��*�'ރ�&v�̞�"���H��r�%�����2�b�*JE<���Sm�����=ȩ�K�d��/*���n�)�O���N��c5���
�cRɮ��yڻb����������=?J`�+P�n��	C
����2�9�F8w|��z���M�$e�|I��>�����Π�Xm�`B�=�Rqz�_[+��o|@y;(� ,��j�
��OCٽ��vc�Nr���S��`ē��jG 6Yh�V���T�u��M�,��F`)���o�q��	"��W�t���/����a]a:��_��}}�+:&SR�}}c�-,�l���;nvf�={���.�T�{�Z��F�<� BF��o�k׮�����F�����F�J������Ԩ��Ma.#8���  6�o�;��1"�Ј3��?�������Y8g-\#��)���d��dР4(
��~��g���������H���`��k�^s�k���ϟc2�`����&�(zc�<�ɝ�MPx��Zd+ �S�{�UC�WԶ�kp�q������w�H���g�#��cQGq��p�p�)2��O�ty����V�qo�#���
�����2���ShEC&���/��.)[ ��`����lC𡪆z�>kq@�P�g��z�	�h4����� ����@����gfG�7����P��nL������V���!�s�_��!uU�F5=�V�}T��=���1�X���@���x?�������4僇pߥ�6^k�ph<�:�����b��K� ��`˚���m)��U��� ^X;X�L������/rc\��4�d���+_i ��$���Y![��m�/Y��`�"�(Y+�����G=)��l�QL)O�A��(�9%�0I�Y�=����Ɋ"�,;��s��MG���ϝ��}��Y[]%�ڧ�P�-]��٦�g܇}�ʿ�q��̍��Z'f�H�|+j�҄�*�L(�� ��x)"�V+�G0��O�ܛ�MwǠ���,��?����/�^�L4��@�zº�Hq�n<�&0�n0�s�!	��~�Z֨>��|
�5��dХ/ϕs�!�	�o����乳g��ź�������`�`���~�T򬕂MP9i �kQ��	����#�	�>�Z-���R�&b��F�^%c�6�ha`�O�3�ނg��	p�}dP�`���@�85RD�����)����.�'�GG���N�}j1��{�
$۴,�#��z��g�&�8������h`���,�\h������>I[����u~Q����8�4xk�X��Qf^����Єܣ�c/joYq,���.Ffl�w_t�.��+^^���[�R|F6��d�u���7i��ґD[.A����<VojY~]����v�DH���?���ñ���1ؒ�8�\��Z�ue��	"��n:�s���%.�[�}>����L�j�@x�LW��u��A����`�9�^��v�4�2���n�$���O�޽��������箼s�mm?��s�l�ncF;�i%Ao��p�+W.s��b�AX_C����~��,r�Z�  �b텾1R��f�Y�F�
I�n��7d�I�q�e���"3�ё¹������������������.�k�������R��Z��}��v  Ǵ���6%��!�� }���&�C(�4��ׯ�Ǐ3�xzfܽ����N��L(��mmn�GK��5�ӱƸ��C2����ޡ�pQ4��I�6|��\��6Y�0p�^���װ�-ĂG���C;���k~a�]��ָn\WE��.u*��6ܝ�w�5=��Ҋ�2��焥<6&�$��{7Ȋ^�,�SSa<S��R5^!��r�-P4n�{�̫|��v�����yF��Vyb�f B���t��qmU�٤AM�o)ڙ`������<�c�d�#dM�&'Ɏ��}R��]*][�";V�Ct�9l��\��Wf��a. z����7Cݴx]3�!���4�.w�ϐ�-�vk�
��$(hoir�>~$�1ؗ��[ߓ�;
(-c_F��}C�|Ϙt6�����NM�n�7E��7	X�J�_Ƥ�qq�p1B4����V��u_�}ɻ��c�v�-h���e2���ڇ���G��H<zg[#��B��>=�ח1�����1X�4��`5ـt�C���[�����C����8���k������$
��kk�h��R�����k��H�  k�G;۔~jj�U�U��y�rs�*��K�R���N��A�Q�Ԥ��m��]����4��a�kkk<ǅ�続��~k[��"��T��T�WΞ=�~�_�K�/1���Y��ل���p�qاφ�z&�eק���\#�X�>7K�)�:�o�	v��ں{��	%� �5Ћ}{.��p����L>�ʺWS/��LN2��^��>��=Jc�sWHH��3�T��`g㻢Yo@s6�
��t�@P�2l���w�.��ә�I숉)ѡր> o�q>�{Ht��>t	�#�@9��ih~�������J�TR§t�_�1*l����/*��9'ůl�S���' �o��+�5X_���dk{�|��x���Q�����}#c!����^v�G��|���#�,��sٞis�eS��������g1���������������ɾ�k؏ o��6�5d��l��i�v�qZ�9)�	,��#*�o!��@jѳgϴ�S#�4v��_#.}�R6��{��E������c^�OB��Bie,\�k�y5 ��9W'�z��U���`d�^����ܙ�Q�p���+RJ���[���F�|MSX��#A�)&f��ٱb�E�^�	,��łc��B�`~nN�º��HKn�U����{��Mw��Wa�|�~���g����>�mVz�gl/�#8�dp<Ju~&	6B�Q�t}�O@^)����5:]�\0��N�/tg�Sr��y�y)m�4L�}C�~1K�)��,^�Օ����p%�X[dc=x@����ٜ�`�'����{��6pn���-����z�t��̡@�N�p(����IJ@|����ڵ����G0{X8z�.]p��WY�oee����8%/�q�ԝ����(���]�q��U(�Vsn0M�p� �k�OOX8oqq@��P8��,�zbRXO`�� Y\Z���&��Ss1�H��l�����_�ł���8��ؠ��L��ϟ:��V"˾%�"��>���c�����s�k���S�`�s-�1�K�u�BwNc�b�*j��bGE�l�E����v��̴i���zA`��̰}W��P�̈������ ���*�n� ��F@(0vl!P�(����o����bj{���6қ�B�C������E��i�]"Μ�P��m0t߀*���'�||�[�v�_+���5 ��9��(�1�l%��c�y	�+>��%{�Qg���yqM���w\�1[G �#�5>��>�$n�D����\��~�%^W��d��M��"G^s0��J�B�)t;6�ʂ�ɇ����*l�"�eG�Np��I�,�F��z�Y��l��d�z�l��x�����]��
�� �)F�1�9G*�M-�'�q���@����������P�&�,�looJ�&���K�*������6 ��v��X��M'�d���QK {�n�i0.�:�#��:���فm8>O�r�s>��c����18��*�) ���D������˂1Ͳ�c��J@H\��eHV�*���:� �dvY�9e� ą<�$�ڱg[q�(���$��v�IR����k(���*;n:<ϰ�p]�Sc,�縖�X�`X�$�`���K�]Wj~��3��]�#��o����-`�Z+C6=��sdv5��R?�g�x������!s�=�vl*R�}<6��|L�����?�[�K����|�C��Py$`�G��6;^�e�6~��1�ߋ]���꜈�݈�(YOK��|���=X�!����aM�^�ʾߡ�'���A ˇ�}Ȇ@M(-B � 8ʒ�ۡ3TZ�q�����Ȟ���F����!5�FXK)R|�N��� �E�5��̝\�XpI���h�qe�G�%@9���G��E/N\+��+Z�:w��h-v�`o��vw	(�]a���Vgk����4N���C�3�������=ZZ�1���i�s綻v��&�߿O�`�tz�a©(���R"S]h��'R_������w��w��/9�/]d��Oq���=C!���
�������͊{�*���j�)uD�:l���� ����;��b79���<8@:^�9K0�ID��RƵ���48�`H�]����ﻅ0�OH������;7����Ǫ�!�fvv���?�#�G��][���E���Rth��BC0` �1�W+��V�H�k��|��}�'���|�)�q����e꼌4�})����q�,�a.��Β�@���t�y�����VV8�pN�I�����>�r����A���1u4O�j�~*�鱝����"��p����1�2{�R��kQ�ɀ郍U;�x��TO�43 )H,Yb[���,Y� �N2��tݳ�� ��d�?�9aްp`%������H�:b�r�&����JKT[��sd�	��m�x�8��/�96���|3�W���P%۸ta�%{��^�t��Z&@`��6T}T��t��Wh@HY�Caȅy^�5Y�Z���h�ϸ�m�59��.}-	05�چ�>?th-(��(�i�!�p���={%��W��z���L�0�X�gU
,]�@�x�Ҿ�B��'���c��gf���3{�~ �����ݾ}�� �ʸK݇���c�H�2G��)�!ؼ�7zZ;sg��S�d:�u�$;rW��υ�i�,��,��7����w�e+Pl	v �;��,{g5�.w�Çi�@v�:�,*��g�X�.�W��K��'������F��f�t�=�Y#e�0) \WI�� 0�g5� ��R>#��8֧�+����E���QjWڛ
�:����0��P �b��1�dt�8�<�s���w4��0�Qk!͒�ö��9�� 8�}dI�#�Q���9.ҟλ���+ޫ�|{����H���𯷽~��Ӗ�+ƕ_�����_R~E�L� �ٵ �`]4I��}�'?�{y�����%o�/�� O�/�ߕh�X��w�ŏ�1?V�kɜ�h~s�Nۛh�����������>�(�t�g��m��ڌX�.12rTZ7�`T�L��-��@��g}i�H_b<J��>*�p.�c�dU�6�c��Tz����va ������~{�����X�u�c�n�٪;wn� 3�	 �$�	��#�L��s���u:l]w����8� k����;A
ǭo\���a(i�������X��:KFZ�: �"2�0>�T�ch��f ZJE��yD���iӱ�nP�Y�t��5��� g � ���w���.�C��g���̘�n��n��[�뽡�	�#�����~��������;��X[_v~eY���#�wEj�Ǣ[2Wj'��]��� *��p.E�t��Ϊ
��XI���x��6�Tp �=9�"{2G�wv���2
��)��'�0@�'��{t���9�f�3t��]hX���G���mΜ_<Oؗ詍KdO�{�� ^	hT�֛�!���YC�v ZQ>�le��EV(��}��g��x�::���p��K�eh�ϟ��~�P�f2ާ>G��+Z����'�q8-�*���+% ��)59��������9|b�F�)�t�&c�.2��1�X��nM`�]8��������*4�OmX�ɭ���g}(ڥR1u����,��9̗����B9�I�Y`�{��7�n�I-Y�/�E̆���º"�{=\-��`�R�R�sG����KI��׽�v���~����<��������3�L�2��?��emB
�B`�"�� ��rO�3
�=}��ݾ}�ݹs�Ei��^cu L#=1������B�}� l<����&L����fk �>Y�����ވy����;�۔���,�;al �!b�!U�eAӇ��'̜�x����W�;�f ����~$��b�E�޵Z`�� � ���"���2���1�m�і��ʨ�P�cQ��A6��c����_�ϱ�9*'T�ֲeH!b�N�x~Q�x���޾�Ez�%�0?P���s��]a�{�,eI[�N\�0� �,����zEe��JP��2Z[K���dD12nϟ����(���`:���2��r������G�߯��.�sڛ�T~��L�C5��Wd-�fcC�u}"�2'��k�,�����\H�58��U^7`���ʧ��-��� Z�ĝ
���[��Q�զ���4�^�l�-�e�mά���և�٘@g�;$vr��dT�9��vmGY�����uzt�4-����'�1 �㢃൲1�L���߿�����0J�'����p�]�r�-=��%w��;M�� �:��F�s�ѷK@���Y�z����:ԅ�������ž��p�����Hxg $ta��8�v^���u0��[�T�}���r]�2elݩU3Q4%]�4�J)
Z�iD��nG��g����
�m�`�ga�:�����>������O��$��-�	�|�^�F�UU=����p�_���]����裟�~����32ʖ�D[�����W�gVq�K��r�0�Pp̴�����C_g�Ϩ�W*�[��ø�).2�E�G��8��.]f��N8�eQY�
0��f�� ;�]:��������U]ʼ��Y��GF)5�#�h����۷���9Ͳ�TX,�*TV�l��a �0z+>�dA�ZzȲ"��=>G{H``�4r�2JU(�B�Y�(#x��}E �g
�Ππ��
�'FuB�
��4q.|g��TS��{�u�}.[@�M�{X���k��v�z>�xo�Vcc�����������I{T�{�� ��R�5  D6
���N��\��,�����5g,����	7�p-�`S�u�`&@X��.�|�/����Z����!f�����ܣZA~ٗ�wҸ<7�l�Z�h����z�����Y���S���k䲉��YC`��Hq�I�OӅ�c��gd6@'�W�/@��+�ʖ�ݓ�5O?&[�$�-�A�x����G\�Jy�F��7(V�-���=�u���3�qvP��9n�z*� ��{���&.x]2p��턑� ����2t�ff�ކu 0g;���=Q
#�d�߽{�m��~c]��a���pݐ̀M��W��΍~�����F��`.�u��S����cp��.��a�@�kz���k*������1e�2q����̘+Ο'0�lE�И��s��x܇��9�Εw�cnYP�PXg#[��q���TWPd[� �<�U�)�B�l�K���Ɨ�,_�ѳ���z�0�K���ا�W���J��̽���a�,���y�Nv�~��k�@�Μ�T�.�]���a�K;
L�}�����Z�}��;*�������Ͽy�vb���>�{ /���暦p�Ь�p�9&q"��RN��i�J;��-����a)��Xhi/~φc6���hL���Y�����nfTG�em�t+�Zh�f-)�>*����ccth�j9q�{��_�t��S���p��+�kt��zII�-�)���}z�NK:dp�VWV��x`� |BѾ^�f_��������\
�'gv6����8�n��tNL]cx(5�p^jJej�op4d�� ��7a1�*�Y��cM�C+�U�41.:�?�%(p��
�Wp&�� ��t�=������-.��y�N���C��ѣ��_�����͛��{�]wW�^u�g��/����`4S��F�0�˴&E�C�.�M��5�3�3��&7�c:�q�݃v��sC�@���Hٓi���|�"I8���A�����M�O���~A���[]D�0�����y�ǉE.\�P��L��*��Jx��(t�39��Pf~�1���o�g/��R zR?B�W�@� 禣�}f$��m}W�BYo5�5�pD�L�f��L2�,x<{�7b�71�xdS��tI*A4���:���qX���v��$�g��-?sY	(���@����`�$p��k$c���@���kt�i�ۺ�w���{q��ֲ�HF�5�����{)�o���;^������9�~�Ώ���~���M���Ɓv���؞Y�-��l���Sv�,�_/�+/��U�$�W#�*�:�?4����a�ۣ$�e��dĀ��u��=-�
]�n��B�7��X��4p����XP��ϼ����,B�sNQJ��t����!e�9���`�@���Ln�uj)�ƶ�{�����	+�i�ޅ�E�a0�q \S�:Ő�b�NW� �ݻO����'�x/�`1 ^�C��%�+�Qd9����3�d�k�>���[��13���\�������#À�M[�L�^2j����ׄ{���̌.��i{?� 0>s��Ew��k�^M�S��J�6�bb�F�2�*�k����!�.��z(�8�C7imu/�儑ѧ5f#�b�����c���(���}{�8l?M`��׽?�v�h!�>p
Y����I�O�����.,R.�{����kц�"��jL辈  |�#�u"��$���Հ��uIU2�W��6��=�i{��G�p���Z���ZL ��_�'	�A�Bey&D��>7��{��dWb�|?M�v૲�8��2��1��Z�ց�	� �ehF��!X)���r_}��{�x�MM΅m78}k���c�ͷ_��g��4���I�s����o���>
6���O���j�� �x�J;����F]ChC"�W	��w�yG��<z�]a�8��^Lݗ���2wm�G�I�@�v=�Bz��^&��'�Ӆv���5���/�}��~�����t��Q6d�ٲ���q?��w���R��"��ÇτA^__���3��Ϟ'\�Ψ#�J�EzbQ-�v�F-�BK���G��@��-?{F�on~��qP�l�0^����Y +<|��>2F*t)ϝ'3}���{&72����o����r�f�TU�踊C=�@���7�uwޮf�t��]�Τ*"�S
%u��U���.=眂��K��� 0+9������j�	�GX��v�?��Gؑ�¢�?Ђ}|�b�u��58��)3EJ�No�~�E�6����t�/3��x)�t�G��z�x�y����N-~�p�	X�z( ߞȞt�ݮsϢ+3`�+0  �~A`/jm��I��f�S�97
��VIe#lfaĎ�� ��(����l s~����ј�X�x��(�4�5�9_q�ּ߳9b�~��_�r�t��Sj�g��9����T�PƿP��h�,0���a''�V@Y�m�7����V��U�C�O��5���P_��`s�����>�{���<��΂)�fw���Z����/Y1�~5�  -+�,�G@�dP���%���Ν�n�[�����ߔ����Ǐ���&�q�! /;;�jx�F���2���<Ǽ{�`w�:�Rv�m��5�|�5Z�ϊ�:'�̷�\/%��B�^2��F�H��,�x�>����@��;��li���ի�ƍ����W�s5��K�?�}�-a��Q�c(`6j,��w	X[�@�����%�i��5<���'>�QW٫F;쯎�;��e��+��]��^���X�D*}v͐|	��"wR����*���]�m?���,�5�m}O����ln�3�
���)��Mش��N�i{#��Q ڑ�֨���/pnL�)�t��-g ��*�����-6��N/y_1p�|��'�˫�2-�,���+l�����#��?�����[dv�u����5,�����}��^p:��GK���V�O�g&8g��s�H�M��0������������%���y�����pv�h�=��.,Rbc�_N�}��3�=u�Eނ��L���ɢ�E��.�����֟����Z)���ή8�{~ l�R
͉̄�j�)rr����-��t�n}�ff����~��{;njz�c��Td�@u�:�("�k�`Ζ^����µ�|4)�7��ZpfMK�������F\�\p�Q�mrb*���l���{%,T8���3�¶f����3�}�����A���`
q�)¨]��1�9\�+�ghO��nS��>٥<�3�0!��Ϟ(�	�����"��X�9h���|��h'>�3�20:�)��{d]I��`��u��t����z����/Iu>��3�5N��xّ����K�qp�E�6���F�aK�Ň��"�-}ʏ|dLq�������~E��H�yF� �Z���g�z�Z��XO�JP� �;j?4hR،Ы/a}{�CI$����dتo1��W�(�DEbpSh���N?�U0�V��rf<Ǽ59�E6�maC�����<ֲn��5���ľ/�O@����n�Ȣp�z�K ̈́�rbr,1���lZ0�!a������?z�*�=e���(��4r��
�V�ua`��DFj@',kh�BR��"�Ȝ!h=�p��I�4aɗj�=딹�{�+��G���V �X� ����1Q��̙�ϧO��6��G�	�cna�Y���sa��BG�m���6��2ڨ��k�ª;�7�>_�x&�`�ٌ,��*�' ���7pM��bm,�KP��
����`\k�	v��<	�����"3�?���������l����U�7�e�G���&6%ˬq��[�h�e4�즙v�?�^A˷p�#(Op�����)!!�=p�N��IvØ�����f ���="�/�E;��-v�$��|;���ډ�G[�T�fU�a�i�̶n'n����z}��������|P���Ҫ�Ta6^�A��Z�*:��ڡ����u�^v
_��|8�N�=���Z���(R�]2�`ė�F�_��W�Q0�tj� ���z�h��Am��G-cup%%���r��V�5 ��s�ڏ�st(��WR�����C
�cG�4���s�q��*
��*_@H�`��f���}��ȰTW�u�ᬔI*z̪�����x�����9�a �d(�8���޽{ԓ�x��կ~�^���E.@   � �q��U��[z��=Y:���{�ڵ0n�{t�wݐѢ�#�7���t����M��4���͹��u:x`�OLLSC�sB���#�.���"<�R!`p��i��Rގ�&-jB"57�/�К��]�#Z+#z�E�<����GF�Iڇ�Q�"c71��7� �/^X��9H�������F��Dh\�[�Hg���I� �Z�-P[�9A�[Z�y2Ǟ� �/e+�ڂ�Uf}���Rbv���ű3�G(��b�u��Ɗ7�O�
5;�d��[��0w�^~4��侥ck[����0�;�k���@��dPz߉�@��V��j�I�7���p�OLʘ)�W�W��ČM1O�oA#��)[r(`2 �\�S6灭��s���Cc ��+^2Kb\�N�rrd�� ����G���?���� � )�б�Xˍ�e��{nii�?k�k�>�P��y���۷�g�}�>��3f�ؚal���Xd~����@����-NG&� u!Ȟ5��KV�d�x�o}�M����Vp�ą\G��#O�.ޛ���m����Hz��@e�		�� ax~��*%/�c�eˎ���)	�STUԁ�3����l�!��X�n�g߫��j�G���"�j����/C��3��]�E�L<�$�,ʨ��S������#{������L3�����qO��v�u!�1�u� v�ܟ^,����YtYT�/;Ï��5O���i�s�]�~�t����.���o�?ǵ�R��J�(R���VTf����8���5�d5Y���I���N4����6���XB����m�n���@�&��_��i;m���/�����9�pt4��@K�pIUOc�����m�ԗ��;�@�'����DgB��Rʩ�gj�r��>�뾾����;��=��"�'lf+:���y��(1�"�1��J�'�C��U=$�׳�� �l`!�>0u��3����yW�Oa�#Ք$���$�N��4>�	I0 x"����1��i�{1mU *��N�	~��쏂`�}ѕ5�;u�5��������>��'nb��U���4] �(���Q)#��X~*��
��.�������
YR�~g.���x,��ާ16�e�M� ���.i� �ഗ%ǔld;���X�΍�J�ӉZ�r�&ojr��Dj>��^��5�,(Vu�8g���$��nrd�o��=���P���2X�7!�g@���X�u#�l��דLy�4�� ��؉�8����ȁ��tE̴(������M#,D̍a=t�;�,�x�.�FYW\���Ϟ��-�y�J؎��4�X\�4+ ���^�R�d� l5J=�o�!���j�w6��q~���"���^����#4�[_!��d��^@i ���zcx��Q`Ųt]�������Z�Z�xFe95�Τ+���.�o�X��PY��7���zv�͟�q��=p���R�]����=מ�8єB�\�����m0� L���Ψ<Ug0���Ruz��}e��Z��	^kUI��" lF�_ Ң��'�EVDX�C��
�6/��D�s�����	�H�mzN
��4GP|~~�v��#� ��GX��Ȕ?c�R�k �Ho��	x�k$Ƶ�$D�� ��OO�����($���)=��8�kf�6�.u�K�QS��+���VjwI}	)�9�)<���ű���P b	.����^ �C �߇.?2�0���(AM�>��-��{#�wm�|�:�spl\J���R�"��c0�����)��u]�}U���A��W��p�����RC��Eu�n���R��Wi�������5V���p� >Uf'�(/�98o0�E�^+�=({��O����D�h�٧� �#�fA�rwg�5
,P��9\��҅R���v�N���^E�Mb�>��˲�4ԛ7k-;����R��ә��?>�� ��ფ� �(������s���;{J0t|~��ײ�#V(P9���8�j'�*���aB���4�!zj0�B�3`�H�h��]:�(����M���8�WG����<��F�h�RG1��
�>iu�
�`M/�Y-@O���nJ	0j 6Nz���8��{�G��4$+�.F�A0~���1CQ�_��W����w��?
׾��I1<����IqD0�����쉓�"�;;[�#��_`CC�peeS�G���ʎz�L��c�ku�a;~u]KЁ������&	������9B����e���9����$�x�"\o�rU�J�XK̉s�g9�`���N��]9�U�F�C�p��)h�3�m����'�K�_*\�
��6����0`b�[��bQ`�A�C��j�B�r�v����5I�B���hj�<F�D�^2�Փ�g(I�@��P(�P�ϝ���Je�J�@��K�S [K�y+�gږH���@R�~�T�����^�/u����b.Uw�Zޫ21f�����G`�0�]��g��U���*���ݯ�kZ`j���� ɷ�c�X�M�Y|��ƥ@��	����^YJ (1���Da�L��\	R���tZd�0}�8� P�1�a)���4�ю�N|X� �T�'��,�]��0!���Щ=0=5�.]�����vMP�g�稩�n��,�;��u��&7�� �!5�����B�
�H@�Z%� ��D�3+���S7�h���&'�&���4m�x�:�e~C�w��Q(<��e��N���d9�]Y������̝���\�����E ������b]���"���gC�H���aW��|�TV�`C��k��E�Es���׹oE��~�5���xn�xY��Lt	�Sk[��F���x���<�R8�W�Ve\/�?��q��NOqa�I��a��~b�l����`�aχͷ���ħa������i?r���@֋5�`���A	ޚv��옊ą�	j���v�����F}�Je#���?`�~(�����
oA�beu�W�S�*�cs����e;I�X��1�@���֚��q�f�xaCԀ�c6�9/�?����fAG@#�/FD�X�������=��A�,MI�l��nGS;���4����y���,"�1;;π�F0T�AV)��������W�N, � (�AK�S��%΍�@��)���ٳ�tR�>y�$VG
3�o���l�JMtT�a������T*K��$�~D�]cC
�;���R���BBbP�#@�kFqB� _��|������~�S��<$P}���P<�g�A�� �pf�����Ndp�_����N�-/?!�ł Đ-��hg�e�h�ص�����Ǣqp&�w��F������u5�j���O8�}�+�x�����h=�b��b���M�`*���cV4,,y/�t1'��:�5?7�V{hz�	j�ji�3��8�XM�#SY�3MQ� kM3ӎeŉ�ʼ��Rdъ�T�m�Ș�?U���jRA`z�l6�������D�u�r*�~�T�ۮ1aS�E�ls�7����}J���g`+�U)�kL#��\N�@ �{��6u�h��������P9�CF �Ό��s����:�G�\��4���SA�v����c+������{�1�1&��q�� XW��ؚ�g�<�σ.f���D���kY/���tp�=�y�[
,���\t�i���,A�nOyNp�1�]-v�@����\��G�Y8ý��� �?<��<N����Tؗ!!Q���P�����x{�+�J�e[ם��2���+�'�{��`��o��FN�],�i�|E���O��Z���Y*�/ �)^���??�,���W�]y�`� �e��Ѿj9��v
�ȸ�~���.r�۲��� {� ��l[��:��J@j{���/[��Su��������10�⊆u�,[��7���ܬ;�x�c���uw��u�~�Y������}����-��/�bfL�-,}5M}�A.�D3�+D,�h��z��=~��u�Ժ�^�����_;N�i{�����)�{��'�֬�BHh�O>�`���0`�G<�4�$I*bc���C`���R�Y(�E���98:���5�@FX�.{-3�[W�6Iz��Z�r��֌?V��)G6��m�j<�B�d��C#?�o�|�Ӊ�}\��oi�16_a�JQ)��ռqn��R�P��Ñ���rO�>f�cG���F����p�9E�z
 �ۭ�p]�Z�=2�X�<�&�^% �s1�)��4_R4g0��	�, �ݽU����hp덍-���M����x:M�x/�2�M��^�V��K!��P+�W1���cX���Ru�a8��:�N�Y2B�uvj���7�������A����Ç��'K�9{fV�S�tnq�H�E�*��7�Bz�&��L�^u��?V�����J����qpd�WZ8	�?���W�1�@�q�s�oXTk��+�XxlU�>�� Oa���HO�0�HNLv��	]ԲcÙ�)��H��#SDbߛ/s_9���F�Q@���Q�����P�</���eLe�I �O�bd�{�;�aK��R�%��@�}#\�,� ����� �|���`��^�׭�d�a�Fʺ敁-lh\Ӫ�A�oNGAn!���(F�dLs,�DͼR�f����2ُh&P(p�8�����հQ4c��9��\Dӷ55�<h����M�U�o������X���㊑n����
qI�G����V��>��+��(b�i�;EV���J�2�[ �06���Q���"����6rϬ?��7�b���N�~:�t	�y��h�k��|�sDY��c u�u��hV���ZA�pfF�h{�.0���`]gvR�����C	,�v2�|.c�1�UXˢy�ղY`O�9���<�tҬ�qW���~>ZZb�{�ȸ���!5�!�1��}0� ��&�`W,P�0��������3�:�<P$�'�0��AydFx�߲o��h�;\g��,,3@��c�Z�K�HR��k��v�\u�r�D�k��X!��ApjO��	~
ⱶb���Y❙��}����?p���|>w��������I�Xp@lF/6��!�$(�w}�'3ۺn��}VLY7��Q��:>�q��,s�b�Z�����k���>�5pu����\��\�w���(�÷(�Mv
0����=[z�[/�&k����Ꞽ�|�kɄlaؚ�+L鸇[����N���>~�4Ys����p�;�dZ�a�B}i��Θ�ڦ���I��m���,��o���1��휤�
���_;TNt�c|�`��6���'v���f�L���K�{s�S��.��s-���N����?L#t
�� +�Sso@@O8�E1^�3�����p��.��O�0'iђ	�
R�4@|���p\!�U�]]�G@tum�M��	<��M�̺مi7��vrr��������8f5u�� Sya��ba��ʾ]�|�Y(0�77���'��qp�:�ht"j�F`��w���N��܌7daW'2���Y*�Cq��Ӹ��j�
�����~�����_�;�\�X?|x�N7�5�N`̛��Y:g``��"��9/���s�Ϭ�k�gE�fg����-)�c�����Ё���	ʑn(��<��j`n+;
��R�P@�3ONMPnc��Sw�A8�%���Y�<�R�S����ٳ�Q�ie�k�SV��xO��<[q��]d@ `H��܀��	ց���X8�Xدs{��V�S��}��/o�����<n;��c?t�D�v�033 �n�+Tv�(Rp;j�Z�{�����6(�[*�Ԕ;(M�!"R�V��%���D�}]d.Y����`8�I_X�<�(�;��wV�3<�r�$LL0�@y��KQ�`�	���@�\"�> �]�l�m�cB]��>+NY����r���b,�J�&��&+��tE��E���٫���/�\�{�q.t�%(([��9]��]��e�E���J�e;F�}�d�7�(����Ѻi"+ߞa��$:l�Lcu��P��:�f�9p��%��Q�����>���޲C׈����F�(�;�4h� @2�V0d��w����j�Z�%���6B��1X��E���΅5ݩ^�f�?e�4����V�Hܐ���ΤOL� ���U��HوN��>99M�����(��N����{O@Q��oMM�P��
� �x񢛘��Z���w�'O��8(ԇ,!f�lp]�>==�~���{����W�-ɸ���-�ԩ:LG���l7����ON�8�@>6&�i�Z������ڸ�F��A��=3�.���3�HQ�Z� �;�v�1������BHxFP���w����������k������U�������sֹ�l>/��[EZ�-k���5K�V����`go�����-u�5�j��J�[���+�`�:��g�=I���F��Z��� m�sY�1?$�ύ�Dg�6\�#�T���c�#ްв���p��O�i{ۚ�����K�4��|��?�hf۱L��\'N��n�:�����8�ka c��3�[7<�p�/�.|)M�i�Kfu.N�':,o���a������'g4��Ϧ_^p��_�!':s0��<A��փ&�����Z���lǙ�������N��C���{a X�5�
� a���
�o���N淋��8yp>� `������%��N�K�u��
c�tM%F�6�+����9�c.��L�=��ty�����g�����ܽK�r|bʍ��Z9�ݸ���ͽЗ5�}s�Ov0؃��ϺμGg����dikƦ�HF��>(�Й,�^O�KEP��W._&�}��E2�� ��L++]k�7Vr�c��g dD�0������!G�e>}��=![�sɄ佳(����j3*��S	k�Y�F����/�t����u�0�V�=ǜ�4�� �b��z�*�ylBFkaa�c`���9��=}��&�r��O��0���.4�O��n�=�I�����㶉����H5bM&���3�bb�,�ہ����yZ���pr��/�
{&��h(�+���t��8EaQ1��#�,;a�f�k]�@X�Z Ȥ�kl���-�Bً�R�X��ZQ-��M*�d���ac*�QV�����V�/���Fb�s>2�qm���5�c$9�y�k��}1�h�N^�5��g�׹��F@��h|Ĵ�\�}�8���i�Ve�
	�Ԣ�����l��w>j�Lc�PS+�6FY�q��u�:��G�ֽ�vЪSD� �!2��I�2H�n��F��1K��1�(;����Q[��b�?������ƺO=�=nU�1P����z(�دY�o�}Ǟ���S��ׯ_gM���u�<pء-l�cp��=�o��ېa�i�\˾y��)�RF�����,�򳧴yl�4[Md+�(�bLX�ԓ���^]-��`�IR�����J���i��fVОH�达��=JG!h-�-�9�z~q��kԳ�p {}��숤Q�����y���w�'�|��_��v�3z��[�Ͽp�=�G��lu�����E�q�u#�c,�������ʱ�qM�}�C����ᛦ������{� �6��K-����\I����*q��e�� Q�XcI֩)��s#�<�R;����A���5����VW��O�i;�����{��}�oAS�8�oK_�\;����7��6��Mn��%�X�L.3����|�@Ki�Go�mՌ8��Yt��k�qbwiz|�=�^k?k��ZN�IhGJe�y�X'�[%�����v��I�ȃ��c�%���Ȕ}O�!ƴ�4�#m�2�8$C-��ĩ��� 6���� XYЭ�'I�HQf��A��y�󒲞�E`X�	1�U��J�q1�q0����d=���g!�e�7��������[Y�`a��z��n�mln��ʲ�u:��'i��e�GN�����������s7���EƄ�T�r;ۻ�Nb���5���?���pfVt�W���x��A��7�*ʆ?1�g��l V�������*i\��x�ǂ����s�ſ��hZv:R���Z�;��hczmm#8�R A��1:NSJ� �х�z�zFZ,�)�	�cfZ��ID0��ٳK����ש��07?NG �=����(��!�(j���,��E�0z]N��=��Ƥ��/���V�ژ\�+-�(�"Œ�=5�L)� P�Ο�F�{�j*�&��m=)�N��Dv�E!�bd�4he,U�+L��������┅�Z�<�E�֘v����Ո�f�j���� z�X,�RE�1?�ؒ�.��&����������EA'�D�ϻ��(`�DqH��I�}���x�F3�8��}YLƢ}��ds����<R ��]9�G�q�Z
�:N:�R0��G���H��������j��>����	�5�$M���i�ͧ!I�6	"x�:_��.8�u�㞌kA?ӡ��a�¾B�3�l�!�S*k�� -�7@[y'��N�.Ƹ��r�m��y���ɀ*X��r@v���ׯ����W�˯nXF��� j���?���~�=�ڵ�2&�d�����L\��s��#0�"9��$���'q�'�iOun�C�Pಎ 9@l�	k4T�AOi���6J7��3�̩9�2"C�2��`��{���Ĥ�_���&p.ӽv�Z�E橣�YVؗQ��u+�gE	Y���%w��w��\��?�/o�$�Y ��;-��؈}-��i�w�R�#�_�(��hW`n���ւ���5���c��Q�n�L�e��gV�k��{�}�Z�j�����}�AO- ���=k���z���u�d�i�����W�c*%b�-��N�����G'a�:m'��׏=�}��Z�fȊu*oњy51���r`Y����Pǆ�U*��C��E�N��E:�7���1����U���=�� �i;m/�e���4͌}S��Z򺲾�)�'̝���"�t��+ڂ>����k$��9��8I%g��`�G_G��np^ֹ���)�q]���ܥ��!��m���(ဎ��w7J1HQ1���/F�:8�LE�t���\�L�A�4�`��/,��i�]/^�@=?�����e�ty��a��B�pumC�Sa�++&��v-�ݽ�-"����,��B����2�ܻ_ԝ�5^�!��`Fc�4aT\���O�~�����G����o錂�{nq� 0�EU'8R
�S���d���!��nhommH&�!�����_�oH=��_>:���V�⻀ �q<�-GB�W��Лqss�t��6V���SY�Dv�4c���mW�	 @�}K'=�?@$*�W �������dY�������0g�v���>��!eob+y�3�N��s��ZРΞe�Xc����{Pk��%g۵��@����W;K�#��0�,U;2}3����`+P�yj ��nř
:�q�*,M�4�2��1$D"���#��vr�v��H||΀`�Z��>��8\d`���=�ݝ"��9uebz�ef�&�a��IC�|�5��ȿaI@2u���d������j��f�2@;�h�����b�C��18`�4�v�"�yk�8ye&r��6���-Z�@�?�}��7}^�E��Eq0/���b�D㘌��w<�W`�^�t����U��X�+�c״�g�����2j!\�;,���4��k�?�9t�)Ar�}�^��/]d�_�O���lЕ+�n� "C���4���Yaî��p/~�𑛟��17�~�ly��#��\Da��G��X�Nh+C�kii�}����Ν���,P��q�L&xؤ��V��f�����"u�;�"�]2�e�ı �Z�G�� 8�={�>yL�`�$��=��!�N=��Xq=�;[�>w�le�w��Ի���Q���3Jl�62�e����u�)~����c����ޞ�̘�pa��ϪVpm�H��+H��� h����;�q���gϖ�hL�B���u����-�Q���@!������F[ӱ������������Ap�L�Vei�u�>,Ć������Ѣ�\��	�������X=��Ⱦw��D�Y���o���Y��u6�S_�L!I�?rDY�[,�-�-���Z���R�Pc��� kM`5�J(���K��`1��9EG^b�"Ylz]������x+6��?m��%7y�_\�"?B|���hhƔ��;)�z$����(��,���@�gW�B��+b�8#\Yt��mѢ����F0��%���&�º�C0U�j4�N�����n�R���1�
��խ� ����'O����}���a+�5YEt" 5���p<	P�͢q:�]���TIq��9>���Jz�p������#� +XP?�����1���i��E
0�Fc&�u�����LrΫH7K����ffg��eJ��J�2�����{�J'/T�է�K�G���A+e����CIU��"���	��Eg���Y�߃ӌ�t��H�l��������\%)���d��v.8��LS�g�ȉi����w��Ś�k��0g �O��Fqʦލ�(�Y�.~g�`�1j�����Y�|��*g�/*���:ۣƼ1�j|�%�O�P�E�WU�Jce_*R���e-��
�����Z/x-��@�����N��p锱��JVZ`�$dWU������PV�I�J�x�.�0��u���,w��l���jE7���[(`ƠA����p�L��|.`���7k��������7λh������v����V�܆�ث����;͞��妼H�]�"�!����O��@�z�|�a�~M���ϖUN�'���.Dʓj2\؄<d(fgf��e T�ɢ�з�0��K���y���F0y1�|�����df՟��glι��?4�q�ϣ�� ��������y`�`D��#�����gϝ��p��ݾC� ��,�9���(�!@��e�8�u�����&y��4�������s ˯\��=���3�ְ�d ��4]l�1��P�&{����	�@@ �<���1Xа]�{
{1���X�5��8��i��?c��7߸'��0 Oو�����_���c����{j��x 1��Y@S�;<ǂ�3�����kx��:/į�&Δ"��˜vj$=ӊ�鰆��ΐ��&���XD��+ǽF��3Pg\e���ኔ!V��g��33�)K�9$;te9�K�i�a�<��~�yHثi�m�E�����g��^��5��Vo�xc�6�,�F�FAec���f1���}��_w�OAcR �R�Ξ9�����R���;���E03@���i;mo�	"�����|%l�d�6��~��/[k
:���L���YT>;ob��]t�;��n *��n�����Dc�
��̘'���Q�)PM֢$�in���� ԭ�3��@�MN�����o8�0ݾy^,�1 01�_}u��ǟ��n���z�p�o��U��͊��p����Q�E��T-Y������t� 39�#J�89@i8� E ͆k�q��?����?���|���<5�ϴSHV ���͕9%����N.Ȕ �l32�T���90Ɩ-��p.��:P��@e�آ����V����b�+Rf��&��*U�� ��o�j�X�mYZ�����zȚt{=-�����P��� �(pf%��{�pf�� Y-���;q�G\�5��&H�F�(JT(H�Ϟ������s�.���sO�8�ΤÂ3��K]�2���=�3���[�G����U˼�̶^LOsY�FF#�J�4�j`G��콄hZ��jF<�:/�Qj��i�1��1�f����ŵ�pn��ʢ� �LR#v�����٧����ۋ��8n���F\�.J�1j�ꅷ�3����٬�]����|����U�]�"�$�2�J���_Y/�,��<6�s������L0��p&�=��>��`�;��2�#��������l�u�ƞ�{���C��ĺk���z�C�<
�"��1G!:gk|�ؐ}Y;�E6XH�]�l����޽{�]�|����p7o�$ ��X��.X���G���>3�Lҁ���n���.�E�6Q_��ss�8ܿ� ���a�c��X���*�m%8_�<��^q� �YO�A[���Y�獶HQI@����������A�u�E�y� /�K����a�F��i����1��?%H����GŘa�X���f�m�>!c���"�sd�a���F�D������C��9>_]j{�la ���g6��:G�wwg��|<|���-f��| �xG�,��<���Τ0
�e�e=H�փ���7�����{�k|0W�0E??���2{Q�\�5��tf����ٖ5}�W���nq)/Z&G���k��՜8���E;�H�s�^�Ө��t��k�HW�/���o`�_S;�����%9�"�/�� �=���{����c�٫��+��|r�N�i����?�E���N0D�tF�쀅�K����9�����ML,c敶Ys�ܷ�aɹ},tcn�O�J�TM0y�v��Kz"�"��;���N�O�	 �cc,tX�ҍ�l��,:�QwX��Z���E�,����@�orr� *�;7;�U���:��5KKO(Kq����|<"��Ԟ[��+�E%��j�SOpn�R^%'�2J���,�/��2��K��[���ʲ{�.����<¡�"�5_���ѹ�����}�_���Y7$��4J/���V6��C �"� ��h�e@�����	G�q��w����{~n���\p��j�qdt����j�~���8�q���Ϟ?ѽ��{��k�#�1���5>��u �"5�qS����/���{�I��E�MX��G?�c��z0t[H��c3�/_u׮^�﬋��:�3�����m�X�rO\�x�=|�D�D��Ev�^�1x�5^���*��@g�B�2�g����˜�d5�ZdO�b9�u\���cP�f��+�׎��Đ�-�ɗ8�����O�b�(�yq-h�EM3�qImĳ�s����_Z2"zO� H45cV�S��.��n�zfc"��P-%���"\�I`��f��6;��s����k,�]a� �a�1;�|"��t��~TC�L�q�q[a�P��6ﷁ��8
\��PXǰv�AF�����Uq�l�$!��$6c����0�C�,����J����2'��d��f�z�,�$n߾�~�ɰ��E�lY�����	����U�R!�3�"0�����Y��Hcp�7d�"X�{�l�z���}�ᘿ��o���*ɨ���Rl�l�+xƂ�߿��%���Gq��6.� �R��dP�}��$[ϰ}`;�������;�Vy�D�Rw�L+��pL)����kN����܇|@{�y��[�XPx�c���s���g�_<W>t�������kG���8�����?����'�p�����6e3VW��=뻱�I��������?��[\\��.{�|) P#�Ұ��28lnV�+�Cz�AA`̵lF�z�$�3 ���l������g	�Q*�L��.K*u$ۂܟ���6&gՁc�#�J�j�t��b�TQ���ɲ0�=,�é�{�ޒ�q��׈����G5٢w�V����6|��W�l��MFhr��
Y��2��x�8���O�e��By7J�4��/t�4R�J�ɲy��FI���G�^Æ�ݟ�|qW�CS-��p�jeW�ᘀ
�������i�ԏF�FS�Zo5��J��jc6��y��1���V�_8#�{OD�M��m��._b!5������Z&[z86����mut͵"����o�7Á�u����A9I'Ǆ�.WL�\H����oݣ�G�޽���{,�H4�|e�7��)��PpZffg�@�y-���E��:�}N�����0�!k���Ro��#c���: �ϐ���_�:8X�u�)�T��
��s}C��B%H���UC����#�A�q?$���Y��H�jb��K�{zrJǥ���p�,.�T(�o� @�aYs>���B�8?��'7Q��8��,Ű,6me)�#,E���	�`7�A5d��\����i�`��q���RѢ���}�������sh��G\;tMgn}#�֍1�8v��~tq���\��XH�g`�:�$bA0��X /�� ��iM��
���Z:*kB��ݝ��Y����lca����RC�~׫��E5l�5`�l>��)�R��{:�4ad���me<3۠ɀ�F�?��s�}��^��O��Ǿ�u��{����Ǯj�ڈ�{�����^��������{<㕲p" ��_	đ��ܜ0���GłV$�����l�A?�����^���v�ۭT&����B	�ed�p.��j���yAɛ=O�����Zz.��nA�2.��g� qQ�S^b[Y������$@���)m���.����&�8��1����9��{��O%s���G�/nrCv2m�WX�;<O�.T�{��؀� ħO���A^B��3<˅�*�^إ<����q̄-b1�00ƽ��C���>jD#��3`�k�e;�;������|!9ҭ��pG$\���u�<l5�E��6�{���|�搵�C��/�$YdJ����`H��7�u|�Q8ς��ܤm���cL����w�s�|����L��L�H� ��,X�A�7�m�|�P���w�vu��z�D���l�J�m:���"%��c6�I)��8��R$�p��)�h=�V�ֻMQ/���+�4���H�`m&%0��_��)�O�i{��"�Yz��"�S~�m�Mx٨^AK�h"��	�?�F���n'X~�m���0��\��}~n��i;m����6DCkE�,��L��CƊעq�>@8o-�׀g�;p`�~/J{�B�������3��!3p��T"� p�O�+�ȡ�
�N��ٮ�z�
k;8`c�}��Z�{cc��c�� �4���4Gs�!Y� !��Z::�)n'g}}�,#�rP�޽��M���G��np��p��_�%%�Wեс���38I� &�:9�/ �@ f	��f@��fp������=ũ�Q HD)�ऎO�˗.SW�����Z�&�c����ﹹ�)�����H�U�R��v&&z��D����yg@��4]+����ʚ�����%�]F`p�E�DkW�l����&��|�P ���0���]�Z��L�{2�f�3��]2���I�>�a���jġ1��3�nem��8�/_R��r�}�)�i�����\/\�+��ς��5I���f0*/]�H�� �&��|�X��9��(�sle+.��E]?[k����uG��b��kqM�����'�,d)��1������.��+]��CT�8a��n_�RD2{}���/��Ҳ ��I&vSƱl"�4���b �wI�!~ƙs&���z�&�}1�#ݣ:g~m���1�в(5[#�LK�`��c���ǘ�?��ǜ���}j�ʃY<G�c��SW���PS�X�����-@H�#����j|&�X�=�a���������,쓷�f�����AZ{� ��G����.$`���sg����4���R�Ng�p��w���\�L[����?~��L�V�`P����q��5���b!;���[���X��[��c��y����yf�v$=��ݸq����c��|��u�øn0h!����+����ODyE�OX� �#�Y�HP��2�Nl��}��#��W<` �?ЂF�sx�Ν8�=<��������*}Nh$�^� 1���4X�_��O���@*׈������?�w��KMx���p�w���+W�~���G?�9��>�����$
�u��T������p���sӫӼo0�	!�D�P'�i�	a)���?[��"I�}���
N#[�	��� ��A���ރ��<�e�/Uÿ,K�^�N�Zr�~����U�j�o�M7`�{�ݟ�Q̼8>���N��
��Sc0�ݸ��h?`�;z�0� � �5�偲�U~�R���V�����������Ёg���]c�=2p�]8���P�
x�8�u,�5�w `N�o*�uYz�;���Q&�9�56������F�OE����H*�8 �ӓnrZ���7ݷ[d����R�}�g|�KP�
���<� �� U��O 3�ᣇdB-穻�������u]I���x� H��h$R��\��2]=�ݫ�S�տp>���zfMuVV�2S�HQ��$@x�̽s���s�}x �HG"��5��c�w��5w��=���eʭ��yyi���Ƥu��J�	���>�$�H�f;kk��hۈ�:���y'�2@��
	3�@a�lUI��=@[i�Y�A ��KE<����3�}�Qc9#k)'�RR�q �s��БO�3��%���"w8��jB9	����!�X��p|��*d���a�X��ְ�è?>1I ��l��'��<
��J1��fS�	R�q��;�D �,z�����ZD���@`0��PN����c�c���XvoyKz�N�vʎ�" � 0엢�t��}�Pp1���Ĕ+J�m�&./��*W�y���� ncK�!-B��@�����Ǖ5��;.��h�8d`����z���� k��Ý��݇�y�k�E �U��z���踥������
2^ϡ�O(���?�p���u�T�<�#n���~��T��h���7��V� �1HY`�%`7)�O/C����-�=Pj#��`WS��~���k�SR��������'�� "$������A-b�Ɓe������>򞫌�/i��)�L�6��ދ�ّ�q��p����|�;���O�{P�������+��Á'N�N��]`E3���V��{[�������`��R���	�"���&{�Z��5��Je͙n.α8��f����O��b��#�����7�ϳ��ı[e���5^g۴or��`7�Ť0�J�Ԋb��n�va�l� �&�w��$��F
1�.��>������3;�/�Z�Gj���a{�|��=w���������:�e�g��/ܯ~�k7���@��-�ݟ��gj:�8/�P�����2sa{+֧xM�α��'-���M�WA�Y����\��V�fB�r���}vb7�j�Z�����PLR���X1���mO ��O�+<==S�m��Q^#0� ��f�M�l�w����cz]�j}y������-��������� 4wR���+q��B/�!�����ƔE����� �_ 
bL�;���78�[Z��������o��mkS���U_�RU�/�e+H�& ���-�2+mán�x6p�����;�ߪ2F���ʂh�@�H
��<W&��wcl4���2>���R�MV
���|�;�w�,���n�.�HD��Cj
�mn�x�P	<ϕE"��1U�"�cm�7|�IA=����Sw�����Rs`0b7�7��L��2uVR`�U��M9�S8%����T�L�6+����l2�*��M�&,k8�R���,��d�X��̕���?�T��%%� ^������:؅�*��Et��[P l��`���h�xߪw1���xM���f�*�dQP%"�����5���iD?"�U
���ɍ�ڴt`4<�~�Uf�#����*��+ ��On,,�x�4�%�y��^�����\��t��� ;�|�WM[�R�*CO���wx��,�K�Ćan+:�l����紂��"������dU�Eʷ��e�u$�Ș�5EA?��4U�� �vR���م�˦Z=��y�H\���|/Z�}b�*���|N���X��{o� ��I|�RJ����)�,W>)?�=6�j]�e[+Awe!1�Tj�3;��gk�|5뼸�kP�8G�:��İu�
JX�4i�,/����M7[�g��Aؤ�=h����������m���-Zw�b������5�2?�#���L��ǵ���A����{:�f�!��r�~Nڥ���;L�Ǐ������ޥ_+�$���ևp� �/���Q����/��C��|��U�k������? q	���2>�V�{�
�=��M�
�Ƭ�ӊ�Պq�~�u��[j��0��������<(���ߛ�8J ���!�xF��Y;
{(��F����,: �v���?b�˳f4��F��pᢻ��g��N}:��}{�{���Q��:��"���6�L""6�BƉ�W���j5[a��ׄ�6���:!6fp+��b��`/U�x�����>�kbai��,�ۗ��	�9���`���xbQ`ɴH�zukJw;c����@� �{oR^��O7��~K�u ���<}��wX�C�Hhgz)��@���Ȁ!��˛��o�m�=sS�v�Jҩ���������M��6���"#�%�ma��@o���I� 0��[����p�Ƃ����겣Fί8�����3�,�̽\����p?L��22�O�<�N=�ǽN��� ���	���ƚw�6]к�׉�-)K�R�U�Y hy��)�3'Ϻ�33���_�����,��8���X��P��_5��궀�Rp�`EAX[sT��%�*�C;7�(/tɚQ9<s� �Xuok���U��K�>�H��[��nme���IK��g�VDW�ު�����e�yVjO:*��L�
!e����,:u��=����r����DAR��p�C�2W�˜8��G��O/\��8�o��������./
/A�� 8���t�)��
��慅��+	P�3�{��{����a3�º�8������cǸ��hG��Ϭ	�����i�i�`�[���B
@�Q{C��$�a�e�*�c�/_��K
��u���S�TEg�a9c�]�k� ";ä�`��qSey@ΕEHq6'I�;w�p	E �Q +*���}�}elb�۸�"��SG̕ȁ�m�Y�؄�D��
T��u�?�])��R�4��;Gn�y��\��m�����x�p6��`�u�/K�����K��v��t{[���������똗����H�p0��"� ��ߊ�B��Ro�����e�'�y���ߔu֯��[�,���ܯ���Y[҂����F��h���)��r��e(��5W���inK�[�v��Y&\�E�c����(�B�V��,Lj��m2�%;`5t��y��߫�E�{d���
W�����Q�P����\�������q�# �M�OL2���	�<� 1ld� #6Š������w�!LfJ��~����.�Z�AAûw�%>>>ƹ����k$cw|ܝ>s�;~��:}�[p��?pW�����/8��t���ٲ,�2-$-Ţ�o���].�o �!������e{��ݻ.�,a=ؾ���s��i��T�8Lh����sAJȦI�|U֌���A'ݓ�z(�4��W�պ�v!��\�m��9� �C�#��`~j#��-����*�'��'�S?no8������Ʋ��o�.�R�9��y�8"Rlb0u��X���=Ϙ-��~�o{h�v�$�������kv�j�fi��0T��嚒iG	 ��z���i07*�޴�`�2g�д[v���=w�ZJ�C��e��8>Qw� ;55P�1R5���q1rL�V-�e�hqQ*2ȼ�?�d���� �����[]���?p�N-�cǾc���u���R ��w��ϕ�o(ː�I*���gyuE�w����B�Y~�ͷ߻7n��juu��`�����
�`GA
��h��L�u�Z{����p0!_���!�(p �)/�+@�'8E��L%�L򚰝�����;�Y��N�w������B���*�1����S^_��;��N���*P��ɒ�#��{�i���ĵ����ua�_ ��k���w�ȵ�>p��hAE�ٺ2�Ἦ�������N�F���٦��Mh8�8R�q]�+0%e�V�e�k8�H/FJ,�H�m�4�Cnn�ck~NAsq�� �ZM�\�-ۮ0~#hϽ��~K�����{�&ncz�׻����Jʃ������5	����GLZ:ŕ2W0��Fy�:����� C}(t�͈�Q����h��ߧ�/<��7h��i±�1���X{$p�9�\`uY��i�b����1�/�^(���=Y]	���X#�'S�d���E�j�(_���������b���d(� 0#�r�#ۜ�=[I�o�H6�־���4��Z3��A אq��	�^$S��`�[_Pj˽X�`&�-�ٝ��5�WVpJ�W�Lk�2_�ř=�+�̶6�\��~h�uC��ȑ#��2 ]���C�sH[�x�����ݰ�]N�J��E[�Lr�L�;�L�$��/:��A�\{3���;��~��ͽ��?rG���+��X��:�HV|r����nC����&�#YA��K�	`�1	�aL�=�g��ˤ_3?x��W����a��.��mD-x����V8k0�a�_3>:Ȣ��k̸B k(�loּ���gRT��1�����,2P���FG��¢v�{�����+[~��Mփ)YW�d���2�����E1������������9�0�)#� ����}x������;q������{��իdq�^!�p`|�MN�H�X�p������dD���ĕXV�
��Lkk�!E"��@�ȷt��-�����J��GM��I�!Ӻ;���Bl�Mߏ��<ȵR$0��>ݎ��E4���x�)%���r�ށ�^6�~�9�b�d�i�R�)8�lY�g�V��i���H�9W�Pa/.�y��x�K~^�f1g:���w��X(�ǔ���%x��绞�����2Z7#�`&��؃����$��I���g���縶][�B��ђwcn���'���1J����w��C�-�C X�1*��ZA6lε\6i|�@��mM#�Զ����<@E��rv�o[ntN;-Ug�4�(��-!35�	b��t���*r�K��I�/��,z�k�M�tf�MOO���'�{����sީZ$� $
�A����8YH�~��ff�N�:�'��`�V��4�r���4�o����}�6�Cp|�h��&lC�-��)�B��8��%��;@�E��&Թ�ݳ`�V#8��&,bj�Z)h"`���He�Jq���_���;~��NWZ�s���(�hD����1��lk�#ӫ%K�*��M�{F! ����3N���?�+k+�Sc�
���JS�c&+��q��TA���ett�l,��b<��!t���f��ʰ���:�(��bm��B�a�>�P�t�T I٩
���B�=~���ni�`\#0���c�(ox�������I0�
M�h��m�5D�|Wˠ���m-2�.�&���I���l��m�f��z���IoG����2Gd�p*u��yZS�\<k�G��S"������Y	�b�O�Za�B_(�F��vE�4�Eydx[�,ǆk�<��ըH,��ybxX��$F~׎w���]'oF_��r���(jЩ�\�Cz97��Lb��K%�4�e��s�F�e�G�9�@�$R𼰷�����b}j��
qE��>c��T$��$. '���W����� �����~:�:%0�u��qY��{<^�ԭ�<25E�������_��n�q�	��Zv�^�ʖ�LI��i ���*D�d����ZF`�@W�;�P`niy��=��L� ��n�<S���?�>� �Ǐ�Vۂ�hU`/�Y��&�����+W����o�w��yާ���լ���0�ۚA�&�1K�u3��uR�_o��P�	����"��,e-�i�b֟�nH<��z��x��ދ�)�	�V|Z�����<���z��}c���ɹ��)<���U��~ �	�`��e��׀�����r�������t�C��斻y���������` j!���q�س��=ƞr �0�`Wy�h���>7?� ' kd��Զ�����5�C����$x���c@v�f�Y�;�5�5%��=>Dɒ~�����<�e���y�_��w������͂����o�@�Y"��D���C�^�3؜9c�a��l��h>Z���g�ж��ϱ�&������h����Є�<�����]�2�ߍ� ��[��\�V��]DPbݘ�E΄+���{R�����nm_
c��1�o��oVl��(^
�(:�dy����n�:V��A�m�:��6���f�:�Y��PR��ҠqK��M���Z�j�Q�1)�9�����L0u66�Rr����w��s+�t���6�J5q��,�t��Q7N0pֿ6���Z��n�~�9G8.���I��Ǧ���ssnvf�`%��`SJ�J`��z"�`,9q"���|���ͳp�  ( ���q,K����8	����b��{
�:��~�-�(�}𡫍�c׎4��})�r�������<M�6j��xR��7�Ȣx���Y�J� @d"<�G�Z
�XM�j��v��.o�r�En�ߝ?ޝ>}Ɲ<q��5���IXC�&�d��Ⴧ�n�
[Z�>�0�Ϧ�:��?y��?y��V@	�*܇�K7�Н:2�16VK�ǽ�[�/��<t�I�0�ь�&����a�b���6@�j��s.6�j�]��쨂�Z,T1�ݭ�8p�(0I�4���K ΅9,�i	 �K�,��s���m�i{u�����K�q	�η���3\�rޡ����;�m��Up;I
�ٺ���T۵�Ryq<��;���o5����O/�dƣ`"9d�5-�I)(�4�G�m�nPJg]�E��y�{�d��x����� gҵ#eϫ�\����,�~��;�:�����-���ᐸPO�L���W���&A0i?��C��7�ݕ�w��Z~��G�K � t7��~�����o��[�O�ŅE�����dtI�O1l�����!A��ѝ;w܈�EΜ9Mg\X�׮]c�?����5�k��%zPR-c�	`��:��3�L�E���|ؗ p�C`<d��SC�k�o�4��a��	;��xCC�̨���q�G���w�{;�"�`n���sb�E�A��x׍�L�"s�u���\�B)쯸g��o&�������/~�FG��H��'�*߽w��-C&cl���C}ꊲ��`�d����K��Qa����ߺu�ݺy��ې��`��\ɺhZt-��V�޶$����ց8 ;��K9�b��S7k<\��dQ��~{G�D#����v,���I�JX)�C�9Em��@�dL��-�[��[|)��F�t����'��_�C�����=]�;�SY����>���ˉ�T�$iN��c_(ic�="w���[o���o�F�e2�踉�I��^f+'��m��y��]a��Z�\أ�At�ި���#��.9SI���C-te�[��@giwF3�^�>'���؀�zp��|ma�h�De1���ۤsY���F�r33O��\u���Ｃ2�6�[�CX�@�e��ɫn��"YM ��@�@�;���J�+i�R�i�p����|}�;�#�Z,.�as%�PX��{\w��뛼a7�nj�TXI�-���$@�8B�\�}�u�S�E�"W�^&RN$&ffg�2��7q�?��ۅ=ji�9b���,���Ў�b�o���D
��ĸ��s,?0��ܡ����^�r�;����l���b��X��N�n����6�p5���:�N�:Egr����g2ȿ!�b��|�T�����6	��H�!�1/����u��$�X�Ke����  ��G��H{��k �ǎM$Y�?"�
[6�̳T���46|{�"O lxy��P<����i۟/-Xjh��hG�N������K�CUS�%���z�6K�x�Fs�$�z�����FTg�d��^��%�`��@�N�T`�eF������{0/dR��X=;�<5��.���~���_�t3 �T�Ď�*� Jp�5P�\( �����e���tJ(*jc��	�(�i��My��j+C�i��#)}�,�Ğ�s�5����q�g^Q+@�Ww"j-;��A��d�f��
������dN�>Mm��3��爠�� 6:W��+���;X�X��"8y��]�as�W���H`��^���1@�7�}Hr���5784����/���3N�g�fߨ�,�}s�j)0����='�=�E�ZR XX�5~ �^ Ȯ�op_m�v5����5}!#�c ��{����*��a���u����{~��@��\(���	�u�{߳��h ��n޺��9�W �>q�������ŋ���d�����#w�ҷ��������?C�	r�z2��Ը^+�I&xbR���Q"E��^�%�m*����^m���_Rrl��Gm	��2��
,���Р8ǀ�eAJ@��Dy#2�����`/`qo����h�_͉����*�$ -�1�w�=�5F|㾐��nW�w�v^{9��~��en';�����v:���񹒎uǙ]!�?�����r�2|����X6�$�Y�C�����>����;��_vXg���ޮѽ`K��E�9;�,�S,%f.�h���۞[	cy�!UN��T�\���Ik�2�.
�!m[�R��X�LX���S ,d��\[��M�O(\BD9!ۘ{�`lk��U5��	�1Du�S�x�tfd��<y���W��N�M7�d�ݾ���%�ޡh�٧�d�IQ80p��4��'E��PQ��s��^T+�c�j��N�RE+�[�\����s���Mװ�E�N
�T#_��a��=
 [0��gԐ¥~Rį�g�!�����k���[���_\� ��~W���9�3�� ���#{�/�5\/�qs�$̙j��7��p0y��YT�\�UhkL[m)O��%`0���~Ѿ�Q��'}
@`dtčO���d�׽3�c=��?ele�B*��mh�tKq�`���=U��b�\;�s��|�[���-�˘�k�u_�iޭ},�C�1���ݻ��P�a�VSY�����@Ϙ]��ۚ���[�AF�e�)�D��&Ma����Y�&�"�X�q8�uǓ�6��ɁՅ �@����'W[Xn�v�=�<��cy��z;"����~�;^�����v��׷��j���(�׷&b�r��5�;�+x�0�}��*BP@���}&bss���~=�Pܕ�7	*��+�S�^p��@����|+��s��(xy��������}�ݱcG�
-}/ ��!)(��-(�"-׹�*W�DY�Jv��bσ�X[2b`���N�r�.]b�ѓ'3�1����@��.��c?X����z����^U�N����Ef�+K${{wC�F�x�t���w˫���瘉��_��=~���.���ʊQ����H�!+���)�Ǳ����j��\1��.@e�\��8FP��<��	�o�� ��O>������l�;8�N��3
��/R�Y%Kt�Yl�{���j�"�E}o�p�<`0�����������O�x�2\Z�����O_��=z�� �3��@�L�D�mJ~all�F�Jt�[��*��;��OX���;nrb���V�����G�h9`���f�xCV�QӇ->�n�����!���,����T�P�E)���9�m��Kq�^�y֖����_,��źXj���N��3آ�e�"�х��K�6E�7YHt�k��]�=���q�X�M
6V�������wQ�ٗ��Tk�p+A J2�����{K[\: 
��Ib4�J���2]݊1�4Lon�)������/��~�ooJ�������Bʎ5)���ƢW�׈jE�� ��6�"n��Ɩ7ĳX�!	k^�D��o��5+(��Zx+/;�f��!�Hd? c�� ��pH�0��w��)���Cw��c�X�W�")�p��4�;�o�qKˢ�Iv�� 8tb�����8<u����0z�`�H_�����Z-�R=qɸ�D�.��l����V��@�H\�Ɵit=��!����nP#�xh`��K�2��(�#�,�˭��V��s��Q��_�����~��;z�����nnXG�A�v���u�m���>�	�����%�E0Mwt�t�j�>��CM����y�Z��vN ��hl�Ui���g�lr�H FU�VSpi����� f?���4]a}��1�E�dڽ������cL��#H7�����(����96i��G�%��eYй�Yh���N�8�M^u}�~�=K�.f��Nu4bb;t��;��2?Fh� �,�W�n7	�G���s���e�'�76�r�<��5̴��d�Ue���/N!����O��I�\t�{�B�3/}��®�~<s^�<���;�D+l���(�����; ग़�J��`�E��p}�P�d�{��ė6�g�uk ��5������V�1��n���8��6hs?��֨ѱ����ħ)u�^��7��p��&�&Ac:���-#�F��C_6�����cd}� /��7o�r}��d���W�UW7��`�3�06�\�9�.\��5��u"3�?2)4��d�k������waG�n ����W@�������Q!�u��-w���Z���t�WW�,�뗀��a��#yQ+�R��@2Wʞ>���f������{�����ܹs��X�l�-�Y�~�����@}y��_�ׯ��פ���XG��`?�J뾿�۷o��:|����w���������t��]7�����1w��e�����}��_���0�a��_\����������s�`�����/�u?�1��%���1 �e~a�=�����~�ڠ4�7l +�h~��n�>́VUm}�/	:Yt�M]��k�8 ht�8ʶV�C{���,�+��>ױ���8���M����Z�-V+8*�=C`-����CP�� ҀX�V�f��圮��@�xխ���5DQ�� ��=��M4�B*dd`[�^>_Dя�r{+�e��,<T�d�a͌?yZ�^Z�6@:�K"�r��J�+�%Z]��:7��mqw�Ε�O��X�)/=r�nO���[���X�*����Z�A�w���"ЕF�F4�k"�Pk0�A�圮%�i�����qJ�]���5�$5'�K�׮8��mRp]�`�)`v��Ҫw>N�s��������� �VV���Fa�U-�0������v�key� #tt&&'���<��$�:S��֦˕�l�2)&r% p���X�z��jUعv�m�lfQ�Y-r �3����i%��`�ݢN�K�g���~�䱻��U;<0>�ZQ��%" N �~dy�|˵�� �l�|���u��2 t��,�V��H��NX�U\{̘IU�MR��d΃=Ʋ�ɶ�em�T�.3 >�8��E�K�&�{�Ѣ��d��L�ElZ�x
�E���r X�:�nX����kI���.6̩�Ǐ�#G���Ȩ��d�KJr~2OӴ��3,oY�-��f/�j�lz���q-����+X��t�:K�4�C*�}����r�rg��d8Y��g�V�R�t��2��<ٳ��,���aW{7�Z|Τ�۝�rx/��`��X��s)�Ujʷ�k#��-I=���>�ڀ=ɂ^dL��Po����[���n�%H
�Tb k
�a� �Ί�}�)h�K�q��:��u���b���j�iy��ij�a�wI�-z7/�y�a��>�[o��f��*���6�f���=�Z��,�����x8���#�6��L#�e�_��L�H騍�]����؁rjg��}:G0߉eH���*
l���F�\���U�4P�QW9%;~�M=���s51� !Lz�XJX  沃4�I�V�����+�oP�~���\���l6 ��'�ugϞu?���*k;����=��z�"l��Y�z���yK��j$�:M���9�V�N�m�Λ�cs����*c�����w��,,Γ����v���"�;S
��zm�S0e1�j`�{�?_d@5�έ� 5� �c�<|H��!5�Ski�:ȹ����䗨+7["��_�W6�~>C	�ul��Z^|,��#/������ί$Q������k{|,y$�Y*6��}I���sh�,Ae�s��!g���"�x�ȑ�A2'`qI��P7�7yE�_����o��0��-f'KfCl�$�@�22�`kٚ{w�[
,��c��C%�T'H.�l���d@D֦���1Ⓟ����N��B{�Q�j�3-�H�cB�*oQ�LE���_��#�nѧ�F��Gy���l�\DaHن�y�`��^]�P��<N�F����J�"`��m�,}H�|�\��Jn�0C�<I�� ��Xt��M�Z �Դ����Ql7�A�L�XO/�cǎ���>r'Nq7o����58V��O���7x\��~KNQ |Z#e|� ϻ��Y���&�f	Y0|j����q��)OG��i�be�7)q0��D�J�)Уʮix�G��	�u�Ovnݿ�zS�#̙�g[V O��SJ6�D��GH?����ndP�)��5�^\�"
��x�`C�3d�$���Ǐ���U�NH!-���� Y>`�ܺy�c��v�+[y��ɂ�܄�a�bXV]^O��8<uȝ:y�@������H�S��꨿�!�e|C�&ڈR�ρlk�܂��1��E��7�R��G�3Z��ɉ�,��1*�(���wt�G���G�l��IwZԂl�cTA�4��yz��yTO�%�&Ho4}sclب��>)���9��	޳3$��:�Av � X�`��Y��k����P�Rt�s��kj$��xEvB��L 6cO�r85F�!�#}��)���H�F�ȹ���ba`���.���=�	c�c�I�j�H��o���#��{�d�X$0b�38�ʤ��4���R9����Ξ9��!���4p��Xq�ޠ���^�P�-&�΢ �S	�V���6�^����u��#�(�rNN�G�r����7��؁Q�vK����X�m������"��A�X��8��G��/�b$j�$�9SG���,S�_�A�*?�B~Ȉ ���?�_��Wnbb�6��~�co5�5��e��´߀�3�ފ0p�0^%hc�D �
������1u��h?��������'�|�����Ò��6�`gZ�W
(6��NH-��X�l�R� "�n(��{E��	�9���-F�c0W
%^����o~�.~�w���W܉�'�_x���\qw���JvU��4؆�>�(���E�l+���Ř1�:�u֪�N�.re�������>b?�OP���f�q!cf�ky��/<oS�#:^ �Ѧ�pM����/��Y������4�'V?a\~�Z�۞�Ė(K��&�˥ݯ�j���j=O?���Q7�t��!�\�� �XF`�t�цW�����h�;&U���1[J���MF=w���?:�r��b}��Z��̍�'�oho%�LG:I�����9��PfT��L
�GxZ�� 7;'�E/v���}�hQ��H��\�/Ͼ >����ϳ�ooLK\QxJ_I��.=ZIIvs�EM�,�� (U�Β�4��L�G���P@Y�of��K�uς����Ѧ���ϨS��"ǲZ�`)�N@��gչa�������+W��U�:Btp���Obs8�SG��~���j�;��1������� �p�P]�ѣQe��d�� #��p  ��IDAT�hN+��Xͭ� �Ԫ�`N�[��B��A�=�8>�L�}���3]j��7��/D�<d08�B�U�\��T	V3qЗW���|�ҷ.��` �WV�"�X_��WS}m�#�$�M��;�Hi�����%�O`'#���͛dz�9����Vc#.+҅��	}��s��tt�;�#t�*�Qe�	x$��UQ��;�HagA@'S]SAkdCfdN�nj`�0E��h������.o�����̢�|י1�֠!Sr��)��K:��5J�7�������Ȭ_ᘩ�'r-\W
"��E�Y��Rsm��]TM���4�=59�,7e�>�L����olm�s'\�c�EP�BK��/�^�Y�2A�N��
�A��,R��>���e����Z������	y������u;W ^2Ѿ��SL�~G� �|bM�>�d��&����LC��  G}���mjQ��Ƀ,L���5�]
�4f���~*�'fI��1����1	�:�ڂ)�{�݊���a=�?y��mnn�k<�`�W����!'���K��Kt+� 0C��/���s��f�0��I �m�`>�LZM4Cf�]�q�?���cV�ÇENcdD���В@r���߯r�J��TS��kd ޝ� �q�VWx�ܙ�����I�cL5�m6���� <�N��@��SnH_еL0�ggfݼ�����_P�[�j�痤�����{�=��g���>��������;~^�����˗�w�.Q�Z�s�4�y��	�駟R�*���s�A+�>I�q��$������^+�~J�մh+H�g� �@�y�⨅�n'��{���go?K�`I!i�mHy�Ǹ�X��2��sl� 9.췷���r� }���p�f~PK�o+j��p+nZQ�q?�	`N:FL���^7;-��;��ȍ��m�V���O��#��Xˉ�Q�=�<^��zߥ���Tg(赱�M�YY؅25T��	>O���q<��{�t�BQ�]͋��g�;'n��{�/���;y�r7 Q0��Hm��8c����u���Ƒ�2՝*�v�� +lxD�}[�6�H+� �̀�b��M�$\D%�� \� L� 1��ۙ���\�p������A�tOVj_��x��sw��-�s��P�§��n���nll̍Q���kLuv��Gpym��A�0uX����A=G�lL�vK�E&���9.��Zpo�R0p����!�మ�.3�)��:�M����$5֜��<Z����@ �������i�������'���AI��F
���
�d<��! �x `+#=unn�Rxf(���:{�A}���<~�
�x���n��@�w�>Z���
�}�嗔%�c�*SK���W�T�Y% �\/�����Y�q�+ �*:����\���Ǩ[���icC���
םJn�vM2���]Ɵ��l� ��˙3g�?�Hva�Ni10�q���;w$���8� ��@c�Y���J�H!M;�+Ia��Op;��R#�s��S8����+�:a��Qgz9�vh�B']�G�3%���}��Z:t��tvo�������mc}�=�2�&��Hg�bJ�t�=���z�#|�k�<q��tnXa�G ul��&3��M)෥��ڡ������Sm|��.�+���1!�, >�N�8���6�՗�������A�ױ�`����iwG~���މg��k�00fŤ�WU����B~w�� �q��/�]��� r�Q�X훪?��C��#�d�M�R�AA�\@������=D
���I��٧���W����XO��D�Bu��nm
���IhcM��f�J��C��Eu-t����K2Y�6���@���a���6��ȹ�U�v�#c=cϬ��0���w����22��Va�,���Y�_��m�{sc���Z�����E��W_1��s-�?�y!�u��}��w����s���m�` �Q��|�z�����u(��ιb<���5��MNLx;b��g�{E���ȕ�~���e�G��ta�=��AC��ʭ�����g�z��-���?�^y����ā�E��z>*FI`=�:���U����a�;���y���}�ƛO�득�_������=��0�M~�t�`�d���k(}��[,�Y
���,��	�B�^>�#"��H��g��S	�d���O1D�	t��Y��@K����跐�o�E��/4r0G�<1�E�D�w�;?��[�^s�a{�E�,Y'�L��h��h	�R��#��D׹�ñ.��I���DZ9bf����q�D_K���^��hm��5�YTVV]��QO�Z=��x���?^s����l8� $����-�~���V`G20���=z��0�Nd�(e ]6���,� 
P��"��f�, k���٥y��}�~��_�O/|J��N�h�J�r������w�����ߒ�s�����_�Y��N^XYa$+������r���90|�{��%�9{�4�[ ИN\�$�e�i�	�eae�,�577���Z�BS�Eyz��[[_�ý���̬����?^��S��Q~$˚�)�B@0�����y:�`��_�t��*�5p�"ڶ`�9�T�;O����2s �� õ�ME'�@M�>,�WȊ�~ky�xyy�2��I�0�{12�v���1����Bg@��Ǧ�Q�dueYYbLy��E:˹j��{}G���UF�)�_����L� J��u��w
��_y�������$� �+S��<ٗ
A#���<UՂ�B�ˉMfz��%�҃��@o8���QWv2`�����=Fj����N���������	k 4�k�[�[O�A@�)�^�SX����hmGz�[���,I4v�d��y��X��x� �`�KAYnyGY:�������[R�%�}&�T���s�>pǏ�"�m)蚆���~�Len;x�/�����U���-n���,W�rJ�φda�� *��!�����_Ϝ9M aa~���?��r`���z��$z�	p;���)�? u��1Jp--λ��$���E&ht���j`�Ϭ!�-�B0����p��|�<z�N?�q���Wa�� �e�cKȒ2-�D�̌���y�v�S�Z�y���-� L1�O�w��nx�w�<����0�I���n}c3����6�P4���>_�`�|��Ҹ>��gt�ش�o��s.~憇F�����`S!����}��wn~a��l6�a�Ꭷ�����'�^�H]� �f�
�$�:fs�Z�G�.�~s���׿�����#GX�2��ffgi�d�Ƹ�3߬q|"�#��3�Hu�A�ɴ��VN��Ny����4�c����;�#ov3�Y�Hz��s2�D�(���"P����*9(EƮ�NH�E�_{� �f&V����4
��mٿr�$1�Y�p�� �զ�sYLQ��]mo��-��K���./��0�3e�a�K�,�6 J	F%�Sue����ؤ��SEޗIcFC1)��J�{W�?sU�O�)�wTH�N����^KJ��?"�1U&'���KZܰ��>T'��ZO��16s1�l]K�����睰��01Uԩ3���z1mJ;o�H�d p�3"�p�� MӾ��
�@���3�wn~��<�:Q5~���2;�bH( |_�������ӧ�`�x����8���<r��#�6>��l�`��^��;/|�?J���533�똦x��{d�l�6����s��
���/_��ݹ}�?�a����>�gQ�H|U��Z-a�;`�x�����W_����ѱ!��%D�J&�s�Dǃ����w��q	 p c��AtC��d����P%V�c�T��sO�����I}��I��� E:��u��ٍ>��(`���'�<�,������1��0����T%;N��˶�)���-E�e�ݾ���ݎ��s��c��L�3~iq!��:�'��J�[�0�{�Cr��@m�F�5k��Ϛ����@F�ն�֕�bep'ld�-c��	�]����^s[~� ��0��q�h����w�;<ӎ��}6��=��f��ͤ)��D+\��c�)�LѮ;�%6F��	���%�s��T��w1�c$g��v����0s�O����~�������g�ƐQ�i3F���)`�E��"G��\�F!���H�(֝V����?�_N@���_E�������*�N��{Ӫ[kuX�F%J���Ȩ����G�2 ��S�1�`�!�~���3��*����V+��.�����U������t��!J4��-$$p�[���u_3C��{�L��,y�en�$K��G�WWs�?6�i��%�L2}Xز�
c'��>٬Lɲ0Wq����_�!K2��HiX ���2�7P�����%�b ��3X�,C���.�%(�liZ�㜟��` ����,���m��n��&9�m�;��o/]�T�Vc���&+�}k=�����o����2@U�'I�d�i<�����X��l���e��_P����2�� 2'�d�tI�Mtc�싦�(�&�f�b�#�Nt�
�����c-ȸ�O��/��8_��n{s���^iK�bߠ��ڌy AYF����<8��y�yQ�/d�������!�.�E��.Py��_��}Z׳(��p0e
BG��c���(��H{;�e�h���04�Rn�^��
�0���̊���M��K7�F�b~�����X��r�ː�S���<�h�*�vb#�	�S�$�aݶ���V�s�ߎ%��.��y��'�_��v���N85`� $A:�"E��9pv.'���O,6V���1o�B/��j9+vc��?2*RJzj.J3��W���o DZ�/�_�Nu���/ݕ�?�K�����W?��T�b0���T=~<��o�J��0cA�_���5"��_��[ns�A �&e46\毩�O@�c�u�]�x�;�� A��?�b0l��::6B�짭-R�6r�'�qF�/�ɻw��%8�)�]q�������Qhx,#8�/��<|����w�ԩ3�OT��# t�8�޴!t����E�A� x�c�?<���7��׮s��y5;;G�'a���ZM�U2��� �ѿ��҆���H'#ɉ��4hTuW�͵�2� �[�@p��$���	��&@����F8�hx~(t����f^Q�m<�߀&���u��3ExT�P3�����F�yM�ŌjV 0@��;wn�`��J���d%C�{��f [�-��T΀Z�p���- ;-`�w"G6�Eϖ��6��r+UI)�8�BV`�+�U̳��%�<Y��?�
�vv_A��YT�?;����r����]:i1��������r�o�D:���V+���p�e��T>ɤ��+������pɘi�1#/ɤXcC�;1��B{Op�tZ1>pM%`Y$��Tfن~M=tx��Jh�c��9��}�p�$����tz�p�W0�17Q۫=a�K��J5�Y���g�����B�*�fc�{���8\>`�Z�J�] E�$8]�D�ߔ �HOT,PՖ=��*�#(�1����Ϟ�cJ�	�ή;� ���=yk��JCUuͲ���~�ߧZMb�0��4�@����Q� ׆�꿷��m������U��?����B���.3+����kpL� �ˬ����ȴ 1��B���&�������/��ߋ���_׎`���i�񝙙'~�x�k!�����o,�LMho�a�"���1��gN�/>��=:-�Y�� �bc>��Z������;�b������ի�����_�^|_���3d[��I���e�hP��=���^l��c�?1.`���G�����8 ���|o�޸�����&&r8?镽3-����"�+ �;lb�S���Ň��9!	:ga���`{x�):y��ܭ�wB�{|��}Ј�^�٧a��?)��ol���&���V �۝$�$}�}��Q0p��H��4��N7�b���-��9�8����ј7��ִD��pB�W�,1*�8��b�����!J�l�ή)"������ǯ�2C}���-��T�*,	*���mk�_���/Dc�RX �UR1D��x�V��E-�Y���vNl�}���� ��#�!״#Y��F��X#h��D�XC����yW�EU�MI/�RE��y'���;�ĉ�d,��?�/d�"m���|k5T�G��q�����,8?u@���ۼ�?<G9 �H��g	:�R�<I�d� M��Ǽ��^�p�}��'��s�ܢwl�޹Cg��w��4������:L�2��͍�PT���!���=u���'����'(nQS	Kõ����d�N,@V����YVkG��Q�'#Y�;��W�
k��9{�|�{�O�S����	�����F'�����bZ���cz*��2����,B�j4�	eEN�:ł=��Y���Ҫ��fb]o��;0`37�t����0��c�?ˌ`�����{�������5?�7�7�\���V�ȏ=��8?�A�}�l7B��Ņ،e�����i���S��ƴ}�Dۛ�OK=fF5>�����w��c��~R]�\�$��B��ة��z{C��$U}sc]	�Ic��y���M���Sv��py�^�١�!* ` 0A�P'��s�Y���a�!� �[�J�n"3���vѿ�=�=��xqwĹ��=��͔�}��J-�[(�z`l�sOd"�~��j&�i$b�+�,ϱ���ze�sU�3
&O6QWZZ�3|�� ��k@YS��[�(ֹS#XH�V�w�ׅ�j��n�udj�}��'@8#��4��o��-`��u�-B�/ŀ�^vD��ߒ=;a��R�ο��e��ɱr��a	��Ma����~�������^!C�������R���Q��#L�$��3lҗ+�V	��X���M���dc�CqWj�jAQ�~c0[J��$���R�E����4�!�q��M�	�(��m���\3�6ʬC��1�J�E�+��s-`2�B_���'d#�>D@���Oo��`qK���!:Yb� K+��Z� �؁����V($��@f�ۅ�%���C��O���9������?�ڏר?mE~a�`O�|���>��3���{���5�;�zm+�hF��?mSi��`2+�A�1)��r�>&aa��1w��G�Þ&2:��Z-��V���z�'�+�]��Z��t�H�v���	*C��N�g�t��B(,[y��w��Ov�;`{������[�>3fU�B�BBB�d*�Z�^��ڦ�����;�n{YϾ�qru�-�K?���I��w=��ĸ��NɎ"�� %I�|���dn���V �q�	�.3	,eP	ë���,�m�j6�\���]Tx+��_�Z�h��stܘ�����I71qD7x|F�����$B�%�9>�nFyn,�����Q������n�u{��I��l��)�6�1'j�>2 �������O�̻��G9]�'s*
jr��8f�w�m	L\���6��s�e��,�������(�+q0x�;66�N�>�Μ9�׈��V�S491��@� �?^t�K������O��ɓǾ�p������V�x�N�ݸ~��^Ga���)�k(jw��aI���=!����&�/�I��-2ki��g���e�t�A��ؓ���`I���������?'��s�:pO�n�X��U�X�w�Ȣ�:@�����ٲd��� ռ����n޺�����$��Ʌ6)�`D�(�U5ܐ������wYf��`P��%�N0� 2;v���tXhKNLN�������RG�@ R�+�b��[;6�XhQu�hΥ`�� cy5j��*�%%@����M�v����g�Z`h����sѧF����ٳg����ט%��\2����1��QRP��R8fa8�s�`�(����T ��u� Wt����"5&���᠋}�q��L �#�c���UU�Ka�g�<n�V�^������l�I�+
� ��O��"D �4��8dE�Nl]c�K��?���d�9e�ٸ�J�g�AfI��xM�b4�a���B�h���n��<�?�q�%��1�I���������6!����g���ݴ-f\0�e�Ə��WĜ�ݖu���kHopY��8S�����?E6%w[�jo3ӄ�E���Ǐ�"w�ϟ#�{���0����;��}�,"�ܳ!��%�E�
�%��,n��IP���z!/�@(�%�6��:�V�q��5�Y�̮���S��s[�#���Ҋ�2�=i���ܢF�dA�E�:���~��{��I��%�-��$J؇ ���B�-Ֆ.
+Wk)��,0��4�S�
�B�2���M�፾�=��U)���#��Ƀ�x\���FԨ�$�G�C�:|�]��w��O�z;���Mb+2a��q��~�+�r��g�F3��ڄ�^X\pS�SWy�?cj��f���Q������øՁG;��眃��RǪ�-�u�7H����݄1��e�p���� �	���>|ݭ�|���7���:I�ϛ;���V���VT9C�{4_�}R��#����2t\~���8�mA*Gx,Xe�G�wm��u�2Z-V�F�1�%I��%�t��Rv�
�E��X<���y9Ii,�n���_{��R�I�&`iqa�=z􄬸�'������l�0���?4��=%M�Mw릅������|dI����6���j�o��o���Z��L$m�����4O��ϧE=�O�̣��m�ƛճ�T�~]j��S�B�pl�����ii�P�]�Ԁ���Gk�˫ZniQ��9r�;�gݹs�۷n0��&#�]�_��_c��j-��0?�"H��5 5����$�=���k��	L��ӧO��.^t�~v���U�q�v���4�.8o�3O��[�$�+8X���ƿ`#�`ʜ:}� )��ݺy�l�%��@��3�74JA�����OJH�XV� A2|>�6	���'''hx�/�@��������k����Ȃ��@�g ��k,��2�@�p�����\)6��|V��{�C��q���:D �ɢVfQ�����Z��2��b�^��,��pl�v<H������k��I��hUYH��
`x�s�NK!56X1vj����.e��/�?�+~���;sر��<y���A
��d���N�E$� x���D��(XBm\��z�`�V5M�
8���3^9N�~H��`���}ū:����� el�'Z��s
k���UX��x�Q� �f��,�l���r�/q�<S�Ɏ�b�M,,z��,������Ր������i���&,d�3�0����&�d!�(�P�
*s���)��8Z\$�%�'�Q(�9�������IVζ[���b���N`fԕ?��p�B���ɓ�>�C�������k�b�w������\�U�$|'�蕄�������Q��=���� �{��)���{�_��_ܕ+�S�pdo�m� t�����L	:�r_�� ���ľu���ff�/	���j4�J� �H���1��ט����h���T�H�	�r�����͌�m��%�?\��"��dj�x��oڄ�X�	6G���7БfpW�+��5���Dֆ�$Q�qN ����p5�4�Kx�c�~�ɟ��g��7�([�Z5ʴjS�x||�]�������(E�k���zɷ��Q�?�B������(i螀 @nH�5T�k�� � ��א�dYS5J���nЪ�A�]fB��3����6	�ȱ�0��hS��G��)��g
�]������VX�_/��sn!�͹�0�C�C����� �g�����՜�K{���9����LJǍ3����V˝���5R�,]
�hl�mM	��hc9 ˺��\��8P�ۀ{�DOP��$��FI���"'Ұ�"J�h���,����ر3�ؑ�><ҧ`M=8tV��
�ĭ\de��zlV��~��4�[(W����۫l�B��A�	4���:�uw��{��w��)��k�N���:���ᖗ����4L'٦��M)�F�JZ:��ީ'`��J�[����Ǽ�����vT����>���wd��������@�M�Ќ�O�ɉ��㝾����qw��薖��5�G�M�;G?�x�)�Ǧh�É ��`�b�؋>�	FR�k�/�N�~[9Af8Y�G��d-=":y�GG�p7�����#����� Z�����������ԑ#L�_X�0Qp�E���)�,h���3�μs����G�����K��}l����cd�������u��?����]?��ϐ�^]�@���?�7:\kk�<����åP(�"H>��4�F�Wxodt؍AG����)�2�g�N[�
]�{�����C�D����nk��Fwy=�9;:�U:�<��zV��eC�30�1�����y"�k�>;�Gq�]o��j�n�#�gȸ����2�=  �_޼y�{5�eG�I�Z��յ��v\1I	8`N
�L��al�y�3 ��]�B��$��5��r���m- �ٵ��	���0-��~Y/
<��8��&07�:ammeY�(+k;w�����m/6_�l ���w܄f��B��0h� ےTy��ȣ�!
�s�0�U�-�
��)M�m��͊2�HvI�������z[3$�J�2�X��h���I]�Ho�� �����Ԡ�;-��&�	@�ȑQ~;y�;u�%�L<����j��y��1���7�l۽����c6�%&6=��L6<s �x��hn�Z.U�{d"a�d�O���t�/_f�����k���1���C�d�fZD8a�Ĩs�n���cE��E`�O�-JbM�RY�\Aea/#�+��$��Y
����-�)�!�f�RQ��&��Q���������:cm���!a��q|�6���_��oj��:8GGE��2P(^����k�t��֘��o�[ �G��g��+\�D�usv�Ѧ�>ux��g���g��o�F݈?�ŅE��L�Y�auu���O��9�g����?���MyD��+x"y$�[�U�W"C.���Ѐ����VX��_>��B�b�8t�;2u�t��>����=��b;dRY}{�����+:����1��L��H�Ȩ'�7MN��r�6f�&�f�?��r��ױ�<�9���c�?��:QVҋ4�����a����;�)������#���Ψr��N�A�!�w[ז�zfo�D�[,0@#���é�li�@� �V&���1
}W0塓t]����݃ ��q��:r�.�/Z��fJVU�b�w�����1���:)\%�X�����m)���D(c�v�f�=z*OK�gG����M��0��2��Y��npR� YT򆓞*0T�����R�n�+��^�f���1d�KÎ���1�Bd�ĩ�WUg9ߵuC���'Ö�}�č���p����w2���s�o�7����{�౛;�/���s_��B�Z��f��㺠�g hF ��˔��L* '!�p,|k-��	�π���ΐ�γ0����0�u2zp�L��= �H�s��{2;ôэͶ�����D��*� � &5�0��r������s�׿�����>�	�����Q��͸��|�-.�xGe�5�2jO{ :�A.]���;��##3�� �W�l�m��;t�>v��Al,<;���u�c8y��$�:V����N8�Um?��ae皮ZT�G
:ꚦ��shRJD���<�����0y��Ä���Mg٘� w�Q�s�����x�BC�Vd�bĥs�s�e^ �`~B�U�z�z]Sۛ�	�.@8�3�K�`[�,3,�Τ(f%���,��(`2�4�0�[[[�����	v]�n~�!�5�!�Ct=��d��o=N����X��} ��c�R�+1��D�h1�:�86
�B?�Ɯ���jtR��<z��Pp+ ��Vď��i�bm�Ԡ�������]� 	�y�]��sl�"�a ��@x\�u~�=���O>��k^]����0���x7s����sU.����\.|�b�-�f{��|��=Y(�`�����㓒�20H�%dݾ}�}w�2���C	�f��cYF��9���Y���ݿ�����s�yF}`Js4D�`vf��6����X����a��ù����X����&x3��C)���XMS�eO�y�"���}1ʽʼ�E�~�*������@�i+�.�~���4�Z������]N��(<<6z��^h'/,.���L��'�=�O95ѫ�#H��! �i0��lɠ����8�~��߹�����.9�l>#�y����60��2	���^L$��E]c?�۫�W�x:{�,�l�
L�=M-�&wV$4P9z���O�f	3$�o�7K0?��iЈ�涿Nȳ�׌{F�GEk���h~��}y�9e�c9��/�/���dWd���iX�׻��X�{������]���l�v#��[,��>���-N�C��l:���H�paS6�m{���8��L�d�/�eʝN���*��wrj}!��8���8�7S)脂\�[�Z��I��ΓK�Z���M��ñ����@����6+^��cg���� ��Gtn�,>cV�x.��(�a�m���rs ��*��`N�` *8;p��7��"�Cex��&�w��9�^�t��v.yG��)w��)�c��o�u���99q�}z��s������N؂���d�R  OdA���'��0U�"�Jpdtt�6���i�x Xӡ���V��Ȧ�@"��ޙy��*`����X5��چ�i ��e0��7� �>�W�ן���6�a_������~�~��/]����%Mq�Ǽ~�oܟ����w���U�l���555�~�~G��յE7�p�k��F�]�����1�l�_aʯi�6��l��;{F4y�*X_+�ˢg�,*�;�`l�
�m�7�_��)������]�c��QHsk�ɱcڑ`l�i��v.>f��(���8���?æ>�J�y4����gӥm�/KA���֭;���ߩ�h-�����D�D k����al:y��㗁�� 3bu�QDs5�s�T��:�-m4�ܙ���2@�,��ӧ�[޶�c*ӹ����h(�Li�fC�i`�[v�C0���=5������EGK����M:����׈�o3��o�  ?HҌ �U��U���q�H6�������%�ߍ �br��c�����,���~���i���t�c�a7����c���Q���w.�T�3���<CV	�L_}�e�6���y��=;�/�� tw��{bm�$�hLZ;���� �U��/2[4M���A�V��͵%S �Iѱ7޼q��'�%d a��YtH"�����V<�c��
��ŷ�>b�2|nqi�ǰL�edd����a���
K���v�^ސ�.^�j��bcP:&O� 5���ё �Q5! ���g����N��}�p��soye��=C�C|_�F�̾�*荾��BÐ��}��b��x�a?i?����^Z�u�="�a�_���2�此��V擬�~�p��O��O�/�T�W�w�n9��cY��a��3tE]�΀�#�kl6 ݘ˨9qx�KQ�B�q�IvAǠ��s�k#l�SQ`)��y1��WE&�k	2�����%kg��״�E����������iU+��Ȉn�u�Z�`�K��j���[�^�\�u��7�� ������.�/�4�5�k'�^L����Dl[Ӣtyaԕ�ؙ��9�4�����wc̈́V@M�[��hֈmZ�k4Z�8�p}�,(��E8�������z�Lq����ڭ�3o���oWtk��s�X#ԹwΏjEX�`P�wgN��N�S����Cf��TV���\�6�d+����)�
�3��! #6�f��re�mm��FԶm��9k�q�i -[_�C�;+�g
�;�>��{����u�6�'3�����ݩ�G�#Zs����]����~�6��Aխ8�����͝9s�?~�;;��PEa  & )�l�)�L\8-�S5}F�FfIɯ�c�Ov�ϼ�x'���N`�Rm��N�e�mn5ݠ��~�Nòw����v�N�puHkx��d�Ӓ
�kk�sh3��������v�;��M 6[�ZZL�]�����s��p?\��F�P)��1��������o~��[��sˏf�fB�bii�E76�DS-S+p#Q�?�"���2*��:�j����J'��(A����1WI�uM)ĕ�)��jl2Muk���ʈ��u?�1�<�}��5�יj'ϴy��^~L67��:��IF:��`FYC=V��˞%h����}U-�l���[�T��K���˘sd�A.���
���	IҒgZ-2�^ D┄u�諂�*�2+Z�ocC 
2�q�h�'�$m��o@m�%��i]DFn�9S���}/���DZh���Sا�Z��@������uY�$�kc��J�Ң;(��v �#��4I:���l�0�r������f�,r��OLp�c���k5��a��&�`�!I��'H/kG����X�$,6���2�F��-Kf��L�D>��a�nvF�\mt���ց�^�*���uX��办{{����Q>^?e��0�w�l�W��<����[��=������`w�
8s��֜�݈�n_}�,�z��מM� 8�N�p��寙� �ӧ���ﯸ~��A˩�#d�Ӯ���2�&��f|���gwW�%���$zOЋ�%�����f��{�y�ff�5�����S���꒪dJ�ޓ 	�{3�#�d�Ž �$R���&�d�1;v�P��#`5<D�ȋ=����Ǫ�n���H�	 P�ǹYl r�6C3J�Y��0���^F@�5�5 `��&����U�����233� d'��[C��Q����}�嗿�%Ar�`; F��Pk��`.eg �1:b�W�1g�tFΝ;�Q�ws��6�e�䔼s��(>�2u̙�Q0 �{�I0`���\��r~��~pϰ��)����/�����?~�?z�t\4iO`mEк�2H�~4^�v�䢤6�=|Dn��)2��2�,1f#��wh� Ѝ`����ksӳ��2��<E�o�i`.�m	m�'O� ��զ��|	�{�m����M@��"�XF��@�Z�ʛ47�M^~U�{��<���2���T�h+�ִ�߬��*�"�U�k̗��k���Υ�c��"^T}�	B��6�.+(�ʤ��֐����h�3���E����L?˙��~����m��)�
"8k�a��Y�S_��#d�,����m�7�
{$)���g��A�;\t���EY��C'�����r���z�A.sN�--.�4ٽ�rO&.���0��g�� _[+���)����:}��Ɠ��<�_d�>�`�L��J'#s�$V9��-�J	�kU5Xw��l�0���J7,���}f�wô�=&��L�g������i A����`%�c��΅�?�3�c|�P0qB�+�|'��6Ҏ��MLʱcS�(��g�i"�68d�T�Б(|��M����r��UYXX�$�k����r���ђ;��������鲁ʙ�Q��drey�]�2�T�ߐ,9s�� �q;`���d�&�I�WDx��*�H�H����ϊ���<8����b�ݎj��r<�m1�4�ь����Y���<��x>Hӭ����~(O���7r����lV�Y��y���CS��eZ,�>ҊD|���a�<��IEbrY	�V�KR5~p� y�N�j�Y!�0_1:��nAf���@�@�FшkY���t1vX}�)%1�citȚ�vL��S8N�Y
`�A�0F;&͡3M�BA��J��ݪ��϶����ۨ+]�۾��C�� ��k?�v*"�� �!eL�U �48d���+�c`4l�8��Y�;X��e:���Z��S�EP9�@A�ϓZ�\';V`qc�a�Mֽ*�4�!#��JmMqR�k���y&�?( ZegjŠ{�@���m3K��HeƄ��l��CS���*�<�gq$H��Ȕ�H�z�p�u�����o���;9�Z]f8Qg8��##C�_1�A���m����� �}L�{%�]ȝP���d��N5m_]W�,�=���:����(�����3�*3Y�Rv�,��c�4S�_��:5tJ��u:��=q�$eBp/P��^������p���8��s���{��Ź���Kg��5���¿{�9ȬF0-|g��<�f��ag=�u�b�7+z��O�L����S,���_|�@4�oe�+��c�Y�q"�-��3'�O��'�r��}�u��|����a3��)��_Jf���E�E����kaR���KY���M��9����YS9Pe��5�lb|�Ũ��'�+`�3k��Fy��������_�w��k��p�:���|~n�{���+��������Oߊ/=�x1m����"?q{k��g6u��M�79�o��[R�${����)B�C�����Uϐ�Mn�^��-p�u��y�����K��&ּkZ>�h�jU�~�)ڼD��}ty���ފf���h�
M��(� 9~�<���7nմO��J��#��y_x���B�I�+�3��p�T�/�l�I���nx�,R�s���t���#�2Xg�sFY!T=���_����o�|M�B�b�2�ϗ˗?����X�k`��	Y�1�J����qNT�G:-��Xw ��l# �h�9D�(9:�����+ ���$����;�C�`Q!��K��~�dȵ��Yd 
ؽH[��FJ8���坋	(���G,��{}-8{",��42o8�������K�9�bܻ4�Ç�����]��+�)��Ld�:������z�
,��4	��y��$k���U�9|��'��7�P�DkR����uV�	��f���;w��o���Eu��844±�c�5�U�@�V��l$���CZ��)����T9Jc8h�l���E��6�%���s�  £G��G�/�P��{w���º V�<'+�X�1��ay��~�e��@��PlYc����(��m�.�H�h���FR�<�l��d(��RB�(I43���38\pM�;��E�Ɨ�ҹ9=�ɮ�Fj3�=+�Z��j*h?[����������N�xO���pf}4y6�X���E� ��� ��+"����BA�B��a�A�SuVu�Ь���6��L�(a&��Y|lP���4��z� �P�A�$���}Q�J܁�]���s�.���k�>.��ڱ�r��a9�|�G���Jnp�mAk|����w��o��偩�*�z?*���^��z#X���ݥ���C������;�șӧ�O_�I�^�.ǎ#c�����C�X�(��{G���?�:$(0&�u{��a�ޱ� �g}iMV�W82�b��!�a1?��4X]0X�I+\�U��Ns��>	��^�bu �}L��5ݻ��@���?x_fϱ��7>�sL�����O'�1��G�	��*e���<��kW���}���� 22� �5��pm]�ލ��l5�Pq{S�G�]���˗?����Ah���Z���֑VJ��Fc(ڋ���Vl5u_)�0�х��З�7o;��T�as���p<����ǚ�z$(B���Y�̎����:�c��DY��lc��cde����{� �r�a�@����c����xx^Ȉ�m�c����on��ms��m��7�1�as5��z�ת�f�m�, W��T:�Xor�׏��׋�Nm���;���m?`�u�TW28�H��[�0��R�׌]�HT Q'�$u�l##e���R�6�k0hm�n�������d�T ���XD_j;���K�o�s�0�	���� ��v{ӛ�>��g�:_��D�FK�����udh��=d�@��`r8�MSr����hJx�`�aS���Bkn��YK�!2�LSY�ɕ�)������"~*'�Vp��I4�s2s����	���tLLZ2`�  ڹs���W��a{��mY\~,��X8"����G9������ ��kW�d�S3:2F�k��)�155%gΜ!p�)�t�V�b��e�,%\�P�j.ͼ�`}С��C�o��Xa|qi�������ŅE9r�(�c����׮]�s�`�2E��ٳg���a/�.�{�s(���:m��G��o���>��4i��jSV�����.���ν�?���?��5<R���4�)->��P�ξKK�#�1�D/:t� ��ϝ#[��i� �'�*W-���mgMSJ8��_�~3�a:8�"O����E�x�\��#9u�S��\������P��/#XՎ��]���z�����j~9y#��6id[m0«ƈ�W%(07.�sA�^�&�s����)
�j`�)MQl/�����r�N�
��.��5de����L���I4��r̝H���+�^Fuݣ� � '��[Jo`-�Vt+�7�;\��g���	x:��c,-���<eo+#�.���UH6~��h`9�e�9��_\�M�_�C ���S�g�����m��f��^��~����E�ӻ"��\:h�L��~�Mni�ɀ��f�:yV��`��#��2���
�BW�&X�؋�. X?�'f���}�u���Ӷ�e,WA�$��.9Ap�r�0W�l�V�ڂg��o��E���.]����?|~~�� ����X[Xx"�u��>E<x����x��#C����r���Y^��
����Z�2+j�z�C�n���+�+a�Ȭ����$�%���E��ﯭ+���fp�1K���={|F?P�nn~�����nݒ��hf�������X=c23�Xfg�,K�>�@�<�GfnṢp.�"\�}��=��WČ���Q���k�@��C�P����-��Rf"��T�Px��PZ$-H��u�H�f���.�;JL�b~�_�z����ܷ� ��>�څ�>��	�R�8;[[�u4P7p:n2O��T��O�wȴi�8e����j>;z��Q+t
��Y�Vd�'��6k��o2��3kq/aPpPB�g��Tx�Ae�%F�L�Գ�t/����7����h��\F|����ح��g}x1`���^���~���XN�#Rq8J#��Xl�3��|Vl��H*��41�Z��Wu���)d�ejh��\�/	N�O=@{�3���k�M\/�(1�"�`��7U��_L��F�^/N�,>h��8޳gB����`u�1���Z:Z9R͞�~3�V#n��U����I0��IKb�h���ܱ�]wJ|C'3L�~Ny�2�(�q�
j/�i�)�Z�t�i0�[r����?�Aπ<��I�ɓ���/~q��[�}�� ���сö�,ˏWx��KD5�5��������kq���5#�����A�@��\���ڌ,�h�,|`C��t��I� O���j� �q/�z>5u���Μ=ÔV�{}�R �4���k����9�󟿕�����!社�>/��Ԑ�{����W���ݿ!��wx�յ\�͆ב֫��8S`Y��qN�,Ƴ�5�K>��}9F���&vcc#�,i�-g���y��W��z�ܻ{�2*O��Gw���{&���Mӏȵw���K�te5����,��X��LLw�J��]W����c�޻��^���<zz8ӹ昅�7��_-.Y��i��<�Hβ�Oa��lŶ�{�e0���X���TuJ�P����d�)%�A#ۭr�
 BA)�- *ӕ�pW�c��E��VF��HU��"��ѾI�X.�آ�З�o��>�s���Ѫ݄�0��'��C�D+��-�L1�?�`��R ɋ������5����迸��q���*� `�.kQ5� P�Ϙ�n[斱�?�yU�����|V�#�-��?.�|��9r����	�5ʽn�"SY_�q�A���5m�/�W���xc.�)o��(b�����͋�k�� ��m�9^�{��]����\��½`�*(���224�9�Z�A�0�Q��ii�tU��;�X�K���|BvQ9YDo��=� q�k[��u��? �
�*�	 Y��T�h���pO�ϰ`_#U9 ����Ps�F���q� 3Y�`l� ���゚Ʈ��V>G_��_��P&���ug�����742�L������?�L���W;V�?�h`R�~����< ��A�U�՟Nis���@Y����һ�X�C�#e3������݃�"�nG7�8�ˀ'=s�3h;=7��`�)+�K�ݡ�Gh� 0N��@���s�4OU	�I	���gx;�䟾�r����5{F�d�8��[^[��|2`w�Z�3j��iս�
*�=T�`04��W+6���g��Zlռ��vϥ���v���gݞA���	��:[R-
�NQ�חY�� �TKK�3�A��u�>VZ�l,���],�b��S�!m�٘ś(l��̖�Ʒ����d�U�s|'�w8X��{�a 4i�wu��ٳ�#7"9��}�j��7a�y��j"+#�U9��WZ�� 97,L2�-n�i�u�t������@Ѻc������e~nV���+i�c��h~���24Ԡ.,�[7��{Ha_[]��	6�8m��=�S�V��!�d��H���������������t��*�qp׈���Jm4�����pC��pmg�] c+�hᜥ���@k�1�Q�����+_~��ܿ���p-zӑ�ѝ����[���{/��/�*��ddlX<|(wo��ի󲲺� �_/R{�=�3��9��xл�D�_��_���=���{��(�W8O��9Uʥ`��I�J�O����ݻtF'w�ٙ�&m1,c�aF� ��4��`9\�u:��&ɼ�pܒ��.��������|!R�~�m+8�gd��&`ן;wN?�az����q����q��IiK�c{D�j�A���U��0��u��n�YW�^n����Z����e�\Q"���M��X[�����ISS�]k����#�g���`��Y�+������E����m��4ϲcJ�Jw�|�ДF���Z�LZeY��o3�I��h��� �==_�O.c�Aj��IXo\׻�_�g��h(cсd����9�����A�"�
2���^$��k��dW�9��/\�>��{�����aH��SR���|���ϫ��n�waY�>H��Cn@?�A�9��+���dleLY�`�:�����0��~��m��7nܤ��={&9�ea?�wyƢ�IxH�(����5<$KK���C��>�[�o�c� e�{}nj����
c5
 q��'�3c(>]xBiD� ����a�E0�##Bv�xhBP��έ.*(�0&	R�E��L�� &	R��U�b@�3��!�s@���(�\c=�l'���2�>�P+����������Oy���_�/���O���%��	��m6Vǲ(ñ��@}�
�U��d�g������|���'�Oɉ���o�~�9��Ȏ�l���yf�U3c��jZ�x�~Ֆ�*���/[�L�vF>��`K!@��e2�N)�ܗlI�ßm��g7�~J\��ƻ~���7-P�����S�m��m(ޛ�Ĺl@�h�g/mUʬ��|RT	���m+�-��eȖ�yR2h�U���_-�_=���������2r�o'�2������X�gD'̮�d|�,�^�� z'~Y���V6��ȟe^�!��ԝ�"I��_'S�g
Z�E�X�7}�����xJ��� �e: �����L��y38;j�[�8�~�,eD�5s"�s�TFeSL*{do`�l
q-<�h*Rb �Z��.��@�3���g��!@���<!�Lv�9[��ܔɉ]d������q���(w��
�ޚ��/���a��{,���g��=p��������/��#�e��t4�L8 ���q;�� Ah �op�V�W	n�oe�(k�tHeP�z�0'N�{)�*���VC٘t��Sy���䓏�<��������2��Eo-�0���+��2��_+33s)h���s�{R'��Ƀ�h��|���z�c(ĵ_���ܿ��`�櫫ta���~3�MHu����F;���_�կ�dp��$���*(�]gA$��\;�1E��vB�˂�(,  -/�t^X\���Aܻ�������.��1$c:)�� |̣��Z8ƒ�B�~��3VA��uf��+�$�~bo���>:���'�����*�y�W0��; ��_�kW��xփ��܈�gj���H����i_p�~�]u<tX_osLy�+��9���jG���E�F�W-g�Ud*�RG�������P����Y���9L��0O�K
�S�E�W�4��َ�s��IT=>ۤ�r�W-T�5��!�A�Q��h��=֔n=Ou��q�To��#�tn[�'���r�F� ��}������·�����#h����sb���*x��g��(�
@�%��UA��I�8�ԿtM���^��U��i�CK���8�����yZ^*$��G����Ǐi�@�c�	�A�w߽l�Y�,��n��+g)m�`'�YCc�Z���s@��y1�0�g�9a'�����l��3N��iҵ�I�t���`|R�������gQfB�lt�#��4#j�,��9q�̳Cl�s����j�^m�v��%R|��Y_�U2���r�{�淹T���2��)��N0��>��#�t�}���\�4�+�'��La��-��!.3Ú"�$#=��,�oQ���������`8�UI���	�ex��c�Ǿ�@"22JVq'���cum���$��V�c�E�Zv���jk�1�,�пÇ�Ā{>�DdbE��^}�A<�qds��U��}��m��l<�`8�����@[Ř�~c�2�d�2�$W�
�P�)yy�M:V�j�h�L�o��%&a˳��;�$�c�;��l�����c[�,Ei�[����z���(r�Ȗ�K��Wo�\7�{�8&˔J���S.��o����������J���b�{E�h�VC����$����Kj^a ZRk���K�hj�%1��x9�>��F�>OO �;`�2,��ڳ����>c��m�&R����0%s`p-U�pp8��y��T0��d���� G�,�ס���gvl�>����?=k��U�F�p����5R��Zبa���֛b�b�����:�f&t޲��W��zc^�M�T�s
&�߿G޹xN����r��CY]y"����e���U�1~�ч����@�F���Y	NkJ2@�!:��cQY���E9v�8S��J^'�$�`%�LB�f�h�����(G��LG԰/�{H�NĊ222F6(��	���ׂӹ";�����H�'+��~���͟��+W�K��z���� ��Lv��%ǎ�[!�}��|���~\�ɉ���ٙB�g;�~�-],��V�X'u�c�b�޽��_�Z~��߆~��G�{H�m�3�}PM�L�Ն���$�1?�f����5jF"vtt��;{�,n ��3�����3�|F�ƕMmN:Y@`�C:�����7϶�/�ޫ�/6in�z�.�f<_�s0�9�c|��>uZ>��'����nd���F��9��T3��L6V�3���$1ǝ1�u�	���
�I�ꝥ�Z 9)׮��_�XVp	`؄
*�X�t��Ƙs�yՋ֥I� �
���<��(|^h�{�lm��m��A��7�ഷJ��$
�c�`��;�sbv��e�5�������^|�EHGǢv�K9�/E�2�W�>��I�H�-u��������&��\ɀ�Uu��)j�doMɘVi#���;'X��叨����[q���M"c�y�����O�
�$ U�X��0�}��U���F:,���=�Mk5���Qu��RK���s�L����d@���7o���I��!D�6������P���{7t�;a�b���9a� �����q������xO��Mu`툙�~`� ����@Ҏ 7Hf:�EM����x������9���{�����vne��܃s/�챖��Y�ib�b#A�7�`��IT@����p��]�O>��A�'Nj�B�!R�# �Qv��ALAD�~���:5�ý�=���޴�5=l�$���2��>�����,�~3N�1\�t��ؚ��q�l9�*��QE]�`���D}
0�a�M���,w��-X�TY�ųb�?qs���/��^\^�/��^}�ɽW����8���0tQ�2+��fKT��z��MpZ�����*���K�ܖX�����8���ճE��(}�Z/�T��I��G���O�G�Ta���~6��g��U���o[t2��op��4=�U��/ri���4�R]������0SK�i�5,R7�u�?r��+�7���u�.Oì�cn�������7Sw�15��Z��Ç�r��j�-u�zH�)E�z�оxm*�u��@�����f����{xT��el48��-��s�Jd;z48��2�t�r !wMLȭ����h�P+�D�	b:�ks��q�	�Q�R@�ڵktH��9�%�Aj8XOR�zx���~-.��i�L_]�����u��5��ZԨpM��99Zm�z{CC2�s��2�z�Jp����ݻ��� W�N���c�Eٵ��-�[\����eٻW�[p��^��4~8�`"�P�2� 2$%p�	}�=������dﾽ&CQ���]K�=���:��5�Pi�T�aݟ}����)����Y{hL���O����nR��E��{�-&��=���F6��ƒ:c�*�����P���C~��]*y�B�҂��;�����w3̱���l�q
ig�q�*x��E����8L�_��cM��Qy�m_��R0�,�E�ywx$�������)ס��";L�J	���Ԁ�(@�0&�v������y�`T^���7��6cb�Y��z�PZ�A�F�>c� ��s^-�k� �{N'`\�I�L�@��K�x����K�sjgyDM�$uMr� �h ρd�4 ���"#E�=�ƀE�ڌo9p�VLJt%�8v����-ǎ�<O�:��Rmpa��Vm�Wij*���{�殯;�F{ـ����06F��+̼�{^F��a�)��]a/:}������c����䝠������	|�΋�����	��R��:�٩��Hm\	{.�f�P,!��fd��C���l1QV��X��:�h�'S��[��m9�p4[�`Maa<L˸��q[f�T��V�N��4ˣ�t�ɅT�ǵ��:�Af�U�a�����VV9�ԪX\^�5��O?����ѣ�t�L����ע,�4i��ϊ!�l�߱��o�f������o~#�Ξ�sV�R3��xv���,� ��΃Bl� ro��e�����מ�����px6��=9�GN�8I�5��/�v�zϯi��Sp�����2'��߮u�/��O�3S�>X�3�p ��9[+�jYV���A���f_$�}%��s{��̣���j����W`�$����xL�+����5�u�$�ݷ�ZH�V�}��g,'qp�{�����{�W���i�����-s�Հ�~��y�V�A�ꄃ� � ,qX��1��krc�w���J+��@�:�0}K?����l���6��.�h1]�*��0@?TI�T�7dqa&�Ctn ,K�P�r��ϧ���Q�l^�q>Hb�����8�>���$fd���j�X�33�B �a�A����eiiE�.��Pk<�'�tBp ���.0�O�:E�
+���8�-+�W�Kᬢ�:t�P}~ǎq~��*�#���u�W!%�L�>�H�vm�������&�L2�e��&׺Ņ��o�A������;c�?�)�P^�i�;Fw���?}�}Z���#��f��|���<�L� �S���5�$Q=щ]��X�!�� ��A����Y�ޮ��E��zw�����x��u�#����+r��a9|��1�w'�!�pR^��`&C��h�1�7,P�U��$m����\~��o�D���8n̎�F��/�/�����/��ye��u�-��eju�|@��5�����v[S��MtPE�^e���4s�������81{D�$t�]��V[+1���M�Ȕ���Z�6���|� {�� V��[��ȗ�Zd����꼃I�hX����v]�ܘ�֥j���*Ofo�� G�-� ��V�L,LK�0�
ˈG�}ƺ���E<ON�uJ�h�����~�nｩ}�̾ɩ�����, �����={x�2��x�
xm����#\�I���C�'���}<��\#H�����-�?�f�,�2����8�g7������M˷�~#��>%�0n O�{�!� ��F�Y֌���]guum����`' T�^���[m����LU��QnŀU�!/@/��ee���i'��Txya�ʜ)F�~f>M�,mLb�v_����YNs��S�|����"�LPCk/`�@�R^'O� kbGu��J�a"�u��&}O���FV�}F����_�.�n��ga/���{�Y��)��'zL�m���F�Q�W���Ңg�n�cL�w1(�ll�F�M�q<��Ç���`�Ö1�e2O
�f��m	���<�Wpyk_x�~'�nog�>�r�Oj�ۚm�g���j�e��.dݺ�O�tȣ|�[�z?]R�[OIQ%M�gJ����O�=�K6zT�줶���������OU����#���� ~�?��7�G���X�ߊ>?"����{��(��f����{d�Ht66��r�$��j��iqO]
�ݎ����8��é|�u��j��K��h�(dIQ�XƈE6���m����,�!j6���{��IV�����v���(.�ܰQچ)nT���l7��߼u�k����`��C���m�Im?�\�4u^��,ަ���'Oeh���4v�err�?q��Q@�Ν����eb�yz��^�'��|��yb�}��|�ݷ�=��p8Lcc#�Q�`���4��VX�P8n������26FP�i����5Y�v̡JU;/0�#�N[%UG�˨y����\��p�?���Գ��>�%�#�3�WV�ӫ)�(~6��6��.��.�'���56�7n���Y����8�,�9�K�p"�s�FMG �{����x@3������iE�||��h�Kp�}��Xt	�����R�n��>ʏ�1�`��k��ı(��t�񬐶����q�kW��Jbi�������Z��[���9^_��gF}���h������g�T^� }����D��)�]c�5#�腻6����4�8�������z��me�1kC������۪�
���w�̽�d��kjr�[0��E���Ȕ��N�6hb$�9��(�5LP�^Sā�j; i�8^+�*�x �e��A{��X(l����!^/�rMK��!�1�^t��]Qub@nbb�ee�Qnř�$�a���>*�:��c1��Y��.e�N�U�����P3��L(�=�0�z��ΉI���Պ}�]��K�HehYUx�ł����9�ӂ���óp���n�# �� �$؜`�.���q2+�)�Ѵ����1|��;��0=�(�i����˯e��,��=YL��8{����a��CK �,P#}��ľ��k�\�X��E��0���تY��ҤY^�Kl������6�~��*�	��H���^�ym-KL�I�@��I�d	�fJa�Z��Yiu���8��l��p`���걷i�5�سO�<){��?�`�ek��2Hر��&'�f���D>/�| ;Y2W�^�����IrF��]��}Z����D�d�{�Cf?�
�ge6E��S%`�w(�X��5�HX�U�i���G!�r��i�����6��-���1e�]37m����6��S��ki�OΧ��:�Nen�@�Ԃ�E�'�fy�Α��,e�Q�1����j[�q��ճ��>�`�}�(�o���]m5 �mXeF������-+�O T�nK�+�:�L`�N���\�2<��3�ߌVFQʈw�&�����_~�/jF��?���:jt4l$�(�'�
��-�3�{j���V��y�R帯悶�v��[ɲp�2M�y `7o�d~���� =����=Y�,F����%XP�G����|N��{u9����@�@[����9*��~ CRF�ݐ�@@�F#�����,8m��8$�?�[7o�m���m�2P��[ ��3'�#t��)�g�ܹM� 8�h�܄�l�y]���c���}������F
�����b��y3Ǐ8h64�%�+0���9�X�<}�Χ1��8�}����9����uX}~ii���SS��Ԁ���f8�����]�5-P_�!Y� �4��:���Bw"*//-�s ���W�4��S�r����������G!��?�M��nk�(�ڙ����,��`��g�$�)�i�uX��`����R#Cm�O�D��,20Fy��m2�6e>;��E[,�����ꗥ>/#����^����-�I�E������9V��W_~����jd�,w�:�c�G�<e@�/��㙒((��)�+��U4���Ǩ\Ct��\�M��`�+��T�r(�C�����)g�-�h��)��'�W�����A3s�H��OE�.��=7�l71�@��j�" ��nS?kE3}LK9���_������Ѱ�(�flM�A�����99��v<�u��BWV����������8p�1�P8��tP��}�jtǸ9|D~��_�T�'М�лlT�M�������x�s���9�Ƞ�"?Y���F�*ٞ�-����1��zˌ��yBV�w���ܻw_���+����/���6������'a=w�,?�x�p<����y0_4�<^aa�e���j{��Fi+��ƍ�,��,-��pP4� daۘ�6W�"�[�ȃ�u��N���qͬ��JP��Q4P�����r]��r»XZ�a�RA[z�u-b���4@S�
������~~��'r�칰�޼�L8bC �P	�hk8��k��u�Sl�XSQ?W�o�b��O>���,����Z��cVfa�� W���$�:���g2���c�F���v��9k�;8:l���������v�'���ʯ�	e���h4 tN6X����P�$M�.�P�/�2��Y�yQ��z�B��:C�^�}��Iu����0��6�c���E��6�щ�1�r�FȨNZ���.C�޴[U���������R�^��Y��?�s��v�_b��+��FG_`��'-ST��^T��R8�T;�˰|K��r��Z�k!�^^��3��Y*�"F�]K/���|c�hz~�m�m��Uv�b��TX��eg Tk�;|D+t� p�鬒a���1Hd�`_Om�,�#���e 0��wӌ� 5 ���Z�pl`ĻFjOծ���[�'�<5jx�� �,m�Ņe�\SS'��?������m���:��}���F�9e�!�0#����"���d)8P]�X��|�q��'V8- ����)����ߩW�L�$jD�w8Ǹ�y�zހW��<��!��6��pKP�,�t�����ٳgh�A^bn.c���'�L���������:���b�$����k,��M� *�S�y�=zT�_xG޽��9r��3Ƒ��P����9S0��a	��� @���YSH+v�#�p[�!9z�˸8]��n�r��d��V7�����5YK}�ΟA�Y���%��X/�tC�):���tS��HO���G�/����}��f��R������eڏ�����	ɘ�(c��:Y�-����Id��ft���~����Ba����bvm-�-��`h���T%ˢ��&z�U��aN)@�@�#�F���f���yn�kÊ6��jR�g�s	kT��9�-�O���B����W���kԋ͔-P٥hl.J�,�����")�R @��]-ު�'����m���Bw���g�z �6a�o�z�k�[��{��Qy����w�a�K�&1��������zN8�y�<��/ܒ���6��R�T�[��&��#|8���q�c�av�����@�v��s��ѣ����`
�eJ7-i�̃�;wq_��z�\����2 �����;��&��G�-�ct�`7�м#�tm^P�'�(z�HM���bZ�i��XMj?�[>��2�c����qN��FFw�<Ui?�޸V|U�k�/�M[[��B�
����;�^�O>���;>�{cĢ��He~��ѥ�6�m�������06�{� �$�7_~��\�r����2��l�jF���b����~����²��"FT�p��-A�HuX00��mNʔe2����Q��~�Y�U	Ǿ�{��q�3��ZQ*���rW|�t��}�������X?aj��e���un5�6�d\K�^u۵T��bk��9�^��KBc!Z�B�m�+jd�x`�Fʹ%��nn��R��7����\�S�!�c�.��D�7�u��?���,[�M���=cǍ"^k�Ռ���%q�WS_���H���I����3K��zv�䩦6�n_V��;%sg�Ԣ�eZY�������փ��5���7cs\��Ij�`l�É���>u��������~x�LhN������Z�����������,��`D��<ӊ�7-+�P^��O��.��*A$�PE�����.߾}ON�:!�ϟ���>*߮^�Ȍ�G5��U��(�"��<ׯݐ������Y���������"�}��|��W4\��
6-��pQ�{�@-��Y��+�� e0y�f�2�e��G(K�cə��"O�(G1������\0uU�T�� UG�PhkxH5RwOLʑ#���&׮���N�|��{�ϣd:߻wO>z$�K2:<B�LE��:t�֍M�N<�	N�c��u��%9t� �٣��������n�Sg�!Y78�/H�K�1��ܓJ�<tP�ݿ'�gf��o�ny睋�&[|bb\��<z�08��dy @1?� � h�p��ge_	Y�	S�7�S�3�+c�-oU��ح�<Pf[��$	���wߥ~$���_-Od|�0�q��U������,
JiEnu8��w��&�F�Z�EѬ���(NSe��PҊ)�]����	un�����XKG7}h8��>NL�Χ���A2�bNa���cL{��u��#�b�|�F}�0X��5j��l�x�ÌsI+��=I�:������sg��q�8>�K�+�g��2L�׾�F���v[A���k1���������Q�X�"/��*c���b}�gm�{�ޓ���wr��a��dk&��LH�w��ϔ���8�/z/�͟��Zg�ˬ/�.��$��N��0� е5kRY7�];'�1�uc�6��1�0��_�E	�;w�q�>tH�ao���/X�AI0�w��-�];8?0_ 
��8�}Ɯ�����O�8�����"r����2�xXa_�۔��-3�p�`�Y��d#(ԔV�"�,2c�W�K��D���6m}2P�Ht��Z�Y�����>f!輸�#��mc#��4s���݂v�Ȉ�S��}����G����b� ��hR��6���3�3�ֲ4�X��k��3�sf�Q:����������>W���|x�U�$�{J��h��T�G�QdW��ڰ^9˼��P��x[�k�Gۏ�ƣ�'�אAx����M+0���Qۣ
�o���c�.Y�]fnE�6�e,��Z��� s�*�5Jy��htt���Z��Kj>5ً8��$���ר�Kl�}�� F�m��x `Gˋ4�ӕs3I\fKb0�����=�I������k��?��J��YڠM����z��on��_U�7��6���Y��v���kp���/-.��1m��BQ��}(�C/�X��.,%\�ӝ	_ 3gy�S�X��v�n/ڢA'�f�X�T��f_�ڸ�O��Gs�t�S"�QC��S�3�,'���r��렑k�����%I0�[���h���e��@�D��*S#%:)�����I�@���,e& o���rp>~ ���A�#H�&�(]����gj2���� �|��TX��L�#��H���^\J��$�HnF�O��*�ԴK �,��]�]���N4v���A ؍�1u`��褀�|��M�w����?��@j5� ��A�E���� Q(k�c 69��`P.//�Z����D�5_`,����ӱ�a�ն@�>{:���R�5P�8���<���;�n��;w)�1��1��C���c�M�� ���OW��Y��U��:�诳��.K+c��:�q�n������EQ#��~k[{u.ov���6>�ѱ�Q���0F��o���׮^#s�@J�G-����[Z�CdP�5+��9� `+`� �k���@UY�	5����[�uGS�NM�1c�@lut4��N�"�&3&��O����Y�H7�Ұ�`�e.4Q�s8"���h��:V�WU���xk��L��uMUFr����:�ͥ�G��-����_� q{?`�1�`H�@��E�v�����e�4��ף^���F!�p	cIm�n�K�;�i߱��d��_T�}�D�
��عk�L��b �oy�x_�Z�����׶8���g����NS9��L��=�mu���q��5MH]k�F�xL�����+�w��h��:����'JH��?�C��.�=�����<W�0�KK �}�C9�e�m�L��u�LN���'N��,��_/��I��Q�p�i{������/]
c�zQ��@��48,��ײgWpq���Cͱ?���l���頧�*M0��1�ˌ��I��t\&M�g�d���$,������T�g��j����Q]3p���%�(�D�ʐm5#�n^�+?� ?����I!����GSu��M	j�Y��zF�v��bC��g�?93�6OX�r�*���T�+Q����~j�9b�����㵴��׼��x�u�Mi�ڊ����952J��rv�E�޾��x���kg9�r�-����ف�/�9[�^n��g8��e�G[��s��Ok�w�0��T_�`n=����������[������D�-�y�-��6��*[% �}?RFy�����^������$S!|Y��UuHD�� *�Z���%�J�!�h�b࠲Y��phZ*��0�:�է��_���no`+�8�-2#��B�4ɍݪ�Q��d���m����g��;�#(h"bi�ԗ���No�Rt����v�vZI�Sy	uL��<�<��������r������,-������q��	y2�$�Α���,��!k�5�Q�ɮ��� ԄV��Bp`��9�h���r}GO�^7 �����9⚘(@T��lͯ=���	�坲`��-�ub;�I]XA<�z�N��w@�>F=e���\ݽ{WV�VȨ	@����t� �!�GVTڴt�uY%`��=���-LK1�= �9��}��+���;�ڶ1����T����\�pp�������;�я���2==C&u ��ل����� ��oP79���)@p��ڨ)L���o	T�<���%���
Z������l~�:cr�M��˛�!�x��W �+~��ܽs�@���?|��!��EX���1��߼^�["
�t�M�l��
19`C�j�@*e}i�_!=pU3%؂�H��K��A�=jڷ���L�&�5+fv�sdi�ī ���d0�)�(G;&W�@��Rf!�Y>�Jup���,E��,�5	c�n ��.�*i�^%=庤 ���<(��L�;�~�x�,g	ΨB�+,N���X݅L]w*���%�|r�X���-]����I�����_����	�u:*��U�ˣ8��SpmK�>�����ߟ�U�ӗ U^�l.�~Jk���	]�\�Z�q��?;;� 13U�Z��s|�,Ȑ�����^�a��:u���ɐ��k�H�ئ�Y`c~a-��	�/@Hn!�9���3��Wݾ}�,Z2�-k@���9�@n6$
�n��e������E�4ӑ�A�|�G�`��,^[���� ��{ 5�#��4� ��'d/���C@}4�����g��
`G #k�޽|�����T�AC}h'��R�QY����v!�����;�u��]�s:˰o�m�1}�b��
���{V�Oк_��.����\3���@UNv;�hH������1�V��v�GE~ͮ㭼��3x��� 3/}f��nS��цr[HJ[Ϗ@�J��hn����(8�f}���9ա�TuQE����)Jk8f�x4���iS�ߣ�!9��w������d�!��=-�/�:�YĽ!I��7�m˯��"����s�_���J37��c�u��9N�i�p�Tp<��kH@H���#�h�U ��B}I��x!�jѕ�iƴ���ގ�`.���J�`>����lЂeA"��OM��
Ghvf��0��v�^i״�<�����d��g�V~7��$q�ЁK%`��B6< ��u9���qZO�~Ya���G,��J7[��YKI�D���_��_���ӡxX���N��?�����pp�Fw�je�B�?#�c��ݕ���B����\Yq�=ץ@�2U�<�I�U�cB/)wm�rxZ�j��j��M���>1�����v�1y��|�͟�Np��<���N�c�d�)Ӷ�l���3�p� @��j�u��^����Xp�q�P�`�dp.�;*'O�d!$8�M+��[
���u���U�ia�<ܣ��y$���l����o�й`�o���	���i�R����� �86
��C  �m5���0��U�O<(���"�z���"����>�c��=[n�v��ˌ��]�έ���f3�Ca�O?���~mr+̛+�Ȝ=�sn��V��"[0�K��2-+��8�:��5V4ƶ2zaV��_�})OSw ��z��Jjv��٢��x��<j��}�T��4�"3Pĝ�7���g5�vr�|����O"�nZ�m%�?���I������c�_�k�c9c�։1J`��)+�@��wQ��q��iy�p�e!�k�1��,C��:&���EQ�:��/b�i����x�  �z�y;-�|�����'�A�*��x����ǔ��
qϻl��.�2?�����0�^s�����Y�U��tj�<� ���O"����ܰ7>|D&���=�����[w��`�8s�=r�>~ �B�
��f��]���&2~ffg�w?}���%�wb��#��k�]���ܓ|-a����@�X��TW���Ç[v��j�#o�������M�Hf+��X۰�b������s�Q�g�^ӃM�t�)Y�N�I�������",j����� �3)�8��%�ߑ.?;3��#�3�o\�/����g`<�!�6ˌI��k� ������ú���3`���+V�Vp�L��Wtl�~��	֥�-Gۉ�Ė������[	���&*���6��v{��s>�6t�3*Ӡ�ʟNm?�� �`;^[�j�
JJ�M*�l�x��]��*߉Ҫ�bXD��<f���X�X�a��,������p����{q=cU���HUn@���R��
Xv�����Y4���h�m�9�r��0]ռ�w��s�4����+f�?��>(X�)uh
� Ю���"Xq��k\��a�ż
���L�iQ7\�\0J��v�nojK�9�s�ӥ�r��ẖEn��0��hĜ�<Y��>8B �4���Z���l����Z ���4q���Ph�Q�K&ښ�c�LD�םXq��~&���Y�������e�5L�l�i>��/�ʕr��u�C�>�h'��M�Z�4� 	��pj��]3�V�_`��� �;8��Ok�;`4A:���2+W�����|� �޽c2�n�a�feu�l �: dH&w�!+ 7Rtq���2~p� �wB�xd4܋U����+�V�k |# �g������mc3f4��C{p���߷���g
����}"����)L��H�>%9�+�Y��zp>x����Neôw���8�=��!(�"^��[��$�F.t�B 	n�n�=+G��������q�j� �|�U�;�s�f*'p��q��㏩;����Ç�5��Y��z/�W����R����s�1����Hw8�])s�d��<vց�}��R1�-±�/�� 2K3�aw������|4j@��@�8��5Z�&70�	�7��6>�U�YzI�����&�(��WT�7q�[ &cV��l�ʺ�ྒྷJ#�@�1鎦��Jh�X{���^���,\>��C^{���Ȏ�o�����߿���_|�@>g��H�>�������U���Y +��[X36��q�>��^��\��r�J	��L���	P8IG	c~b-�1"|p��W��?���C�⋯���T��1��}Eg��[e!2��rϵ���e��(�w�>�O[�}�_���̼A���ӧ��R�K�+�ye�d��h�3n�����{�{\�F0���F�R���_E�"r �ɢ�9.'N����Sr��1���=��1����S��'�dk���<N�6�h�R(b{���L7�Ad�������{F���i�r�*f�n�ڰk�UB�e��1�9��9
�)�-�>d�`�i��k@o�=s��������ؽ[�;&gΞe�c�
�6��\IM�Qq̭df���:�3[2��=�[�ײ�k۠�˴r_�%����_��=�",d|�Bº�����*4<M�@�R������@�#Y�^3P6fL����a��ǌ����&U�0?�zc6	§z�L���EJ6���E�B�PC�us��[�`�\�qUk=_)S�I�u#��JRq:�$���>^?y+�l��L̤��t���R*�a�Z�~�J:�k�w����x+Ҥ����7eO�n��Y���B��k�B#m0��/4���B�� \��f��a�.�������J�G�`��W:5*<}S׌r�+`	2	��Z,��r]z�BFb�4���u�~p2��Ôzx�xV�N����{��O�ۯ�L�)�p��y�X?�I�<�KQ����b>8}78V`�"��l��^�~97p�ƃ�'�p�kH�U}�!��d�tb�x�s��]\|JP�,�	'"��`I!�+KkV�b������^���Se��^�Ht<1&�\�E�6�����}0�@����!��	Fݎ�w8G` �<HôϐS���	�6��XBO�����|p�����w�`2s��:0�{V���*侀��?���l�95 s�����O՜�:��{k1������H���������U0_%-� #@e0��>�΅���ߧ�y.��6��On�Ӯ��Hˠӆ���	y�>�/��zI[�Ldg��8�W�T g;���X�0�1��u�$����r�,��jU��<&k!��\��Z롢�j����9��5�����U�����gpל������cX' &��b׵_�xl��3w��#^�r}�BVu�m����hV�K��9�n �%��`�XH�ƽ���G�CT���X�>��'r��;�\�+8ġ�@R>�US���W�l��� ���g�����Z��/��u���W����8
I+H捎������SQ=���N7�3=q��عSv�}����r��u����F�� ��(���5���k�J����k�WX�p�T4ء��3���|�1k3��ߍ�7e`7�X B�C�h�o�������+�C��=���?�.m�Y� 0�.�ؾ:55E=�˗?�]{& ^}�s��|��,���ˬ�����F���CQwڳ� �Bsvٸ6�}���#212��!��KK��q��]�q�	�� `�0i���=��(*��P�|�MϹbR`ön��1��5݇�=�B������T���]�5k#��N���2����b���Ï݊��϶��[8v��5Rʶ#�sjE��K�*/����ύ�P�~*��ٕ�
��Q��� L���h��u�ֶ65�[*/dk'3ݫ{f�~JJ���F`Y��m#")	�j�&����ف�T���u{3��fA�ˢY�$'��3d�d:���Kio1��řD|���M�x�8��`��*��V����,��n����E��wǜUz��DjNW�[]�+`yF�Q0�ڸ/x�MNTIT�����S��c��(b?X$��1�^hD]A�֡�`��B��T��� ��v��9��MPm��6B�1y�7
�9 &�$轝=��E��D�W���RYo��ևXsVj�p��jfv��b1�D�2M:�a�%�V W�\��V��(K�T¥�Y6�f��Nê\�vKv�k��<KeltV ���/~�L�ܺc2 ]� .�\�F?�#-Ҥ`>�}	$�:��d,<p��6ִ��'�#������83�3��W_Sr�n.]zG�=L�2ؼ(Dt�AB�๹y����U��Ŋv�s �]C��e8b�th ���V�52"E�?�wVtF����xzҦS��6ҥw/�ɓ'�hp�L���\K��p8q�ze%&�zx���W�����*��_���ʭ[d��\�2'w�-ȱ�������i�(��%My�s:���ٴB}�]�&({#�Y5��N���[{��zۘƾ�}y�V�7^�Ӥ�.~{�sU�M���to5`����bz�Xo>��2Ae�' R@�Y�%��w=�{ܸ%0����� 9|�*�܈�Q�����uǗ��}I�BJp95pkTj�ҫ+���Ogiϔ�Ib��T����nW�ܞ7�X�/�/�����VT�X}�_'.�ui��!�� ~%�\qzJ@IⳖ����;h��2�/-���W��]
���1/3�R��4Să�e7 �����5��ߓCa=��P�����*�$%����O��{18[1�܇nfW�xL?��鷸.[��>��	�}N�p6��I�T�:6l���ݷ��&:6�����1y��;�э��~��/�ѣi��O_�bث����5���ֳ��65â���f���Iv��"��1���C,̶k7˻��--�0�;;;'�`��{��T�?d��x֪��Zг���GEe��	�?��X���Zkk:�i�>�^��X�gϜ������a�0���w�z�j��n��p� �/�lŠY|��m�w�ѣ���90lJԵ8}zJ�_� ���`��+�%��W�I���r����^f�f�9��Ax��,��p}���dn� 4u���}g57
��;Wjk[�\d�!� 5�k�Ejk�!��5���q�$�\� j�&����l��ݓ�y��E���1dd���y��1��(�۰�ϩՁW�D�����Z�Jm	�Yf����C�#��I�|ma�M?�1�O��\cP#�B�xW�J&�~F,�b�x�������1�ɪhqO�����=�%�~����%��8۹s�j�@:��Xs^W{��e�ҐvօV��1uŜ���l�.W�_�*���Ǐ��E��Mʃ�^B�����[a���[�VY���\S�4:�(�w=�GDs\C���r�i�U�v��R
�o�����>p��{�����a�1�8oF����0�V�	 M�/�mb�3�eT�;݆U��#���J�n��ϨӔj�:���T��3M��HL���N�^�~kIg�c�� �>�Ӈj�ǎ����������	�G�A�R�թL�@jqMW$�!]:�H��ڄs �ؽg���@��C�����4nx��9��={��B+�ȑ�k�n}��M��|���Y�����#��.���æ7)��P��:�����"}��iq��R(�=�e�
�X�\�i���¸�p ~_|�]�ٻw/��!�SU4S+8��)t��(�3��$8�kk(��23���ᣇr���`��Į�,@x��~jW���	�f8�����Yʖ�ޡ�p�����7T�� a���@�s�_���mW�X3H��0�<���m��PIcm���| �d������\�p޴�3:� !�
���ɰ8{�3��W�ﴠVZj�F|-fb�WB,�~���Ƨ���mV
Θ[Z2*�Q�aϤ���>���7QY-�ctj�ʧk���l�z@��=�~��>�r̶��HK���F��������D��>��Ҍ��U�0lnZ�TOwVC&<��Tf��E0��g���#2ּ�g�ʎ��P�Qaz�雿\Si�=�_߹���*�N(�jW�x��,U�*a�G^q�cx���fg���4ur*��9����w��	{Ҍ~�� 쯣CL?m>U�W��������b,X�=��&�w
W�+�@�X��;�� �	_ ��,�w�6x�̆�f�ڸ%pܳ��/��8E"���X��"�w�5 ��ݓr0�|�OM��Sa�c �����u�6��)b}�Q#��*���yeUeA��dH�e|�����U9쭩SSUVF1�X�M�Q�����B�_}��|�͟Y��z�7k�(*�w��X�"6
�H�7x�3��ۊ�f�|a��>�2���`Ű��]U�WI��y�Ƃ�'O�`�c�S �^�$o����YZ5$����r?�+��׹���H�I�Er�x�#e,�f�i2�-�|�B�,��}�����Em��X`5{V������Z�Lo��H}n��6����;�y3x~��u/�m��߽y�-2Fৢ1����˞?o9�\6��c���X]�lV��3�}�T� �cUY���TK�+VFŉp`6�8��:&I_�5c�xCV�[��4�>�'�f�,�����R��Bfi��h��_���U'ѝ��7���޼� �����R�4U���F�����`��8q�sayq�,Cl�`�)�O����t��@e%��1�LòX���	�:[�ͅn������t \�ށs8�(��"%u��"ٶ`����mpVef�벲q�X@�=�,���!:�pVL���x8`H�`|��I��w� h{$8�pXnݼI� �O?���B,/R��zǮ���ݒ��������X�r��~�i4��e.�� �lD��G�����Z�8o��>�G,F��8=�2\���x���ý���wߕK�.�Ʉk�v���N�������c���O!2==K��ѣ�z��LN�3gN˩�)ٳg7A*���V�כe-����gN����Q:�-K��= �7̱����S1��ײ=Tq��k�g�7��V���eh(5����!eڳnߺ�@֞���󝥂y��ky�\t���z~R�6�H)r���w�
��N���J�([���Yʴ��|�?�Xlx���b�+�r���4��۷*㥇E[AF�d���]�똮ün��]� �o@#J)�����ϱ��,2��Z���9��R e�{v>�r-T����E(��j˯~�K�@�@��w��Ɣ{�_����X}� �]ɞ,�W֒j~����U*��oX<4��Dz1ס�(� �a��=1!|��L욐����>���ۮIF:t@����}�Tã#���`C����h��\��%�2vs�����E��5cﾰ�hP&��Ep4�q_}����˵��d>�G��Vy�ӕQ)Ic����yX�FN�
���c �ǃ�w��a9|�;~���<�������._}�%3�����W�6�̡�LD�07:a!ۍ>]C3s�ܹ+��pE����`? �7��%7Hg�T'#���cMMw_['���/��?��\��3�  �����ך�c B�H�"^]�ʢTk��>���Y��r|#"PB.�gǺ�h����@�Fi_CC{�õg*\;�XS��\��x+�O��4+j �v{�m "e�7�rU_v�s�ι��N�A��&�q�%�>%q�T���k�*��7X�ȬP}�J�5ԗ�e�~n�z{/��Ќx��o�9���s�߭��n]��I�6-��Hz �	L��$����m?`9I�X@?�t�Z��Bu^aɤ��@��0�8"�Њ�£/�����-SM%������g7\O��/���]gy�ȵ���&@ �@Z�ZG+/�E�h5Mϯ%e
|Zh���pc,���`�=�c���:?���n��-m��Y�x�g6�S:Z]Kg�{У�Zд�!�#��7o�s��Fx�֤ʆI�aD��>J��5�t��q�K*�詉_y<��`��%\3]��eobv�1��V�G��$:`�_��L�nuR��"W�\%s`�{�]��Ƚ���\�3�s�.vM�����Q��	ta��8Ea�B?ա�,J�|2>���d�w�U�y�@�ݿ���z��A0�V��	��{���y�߸K ��o7+�ҋ�PgHm]U�Q�OV���cʘJl�Wx��f�E���h^7�|���5�ǣG���c���3����ME����!����S�mH=���=�v���o&�}sW�^�����	�;��T��¸"C<��嵨��j�k��^�>
�7��_��Z	�<��8���EQZ� �)���7p|<3��f�F�(
�g��������������[>���E�a��KS�+����U�^��z}��Q��$��܏��ƘM������^��\#�Z	�³ ��<՟�@�w�<fijE�K����G*��(E��9}o���ἲ����{0�T���?�,n���nc�%���������=�z�k�rQH�H�D����Y� Ё���r��ijޣ�,[E�����?�#�t�T�Z�d	�Er�{�{��>���w���3���ݙiA�$��"K�*P�@�������#4�%��, ��!<<�͞={V������]/� o�Ay���[˿��@���h[\*��`���T�9�� � � 5P���yX���+�bi����]�� �D��C5��ѱJ0u0�q��R����@���Ҡ^R  �b��6�s����;� ��x��!����.�-�o8�kR���½$� 0c��q�#|����P밳w67��߾��ܿ��l��DE= =�f+�зHJ0l��������SS�f�NI�ۭ�����n�>}b~��0���ߔ�� b|��c�<��y���Z�;b d�(+�⋶"
���ٹY��lR0Wd.�ξ�PGk�g\���T��FA�b����0���,&�|.�-հ#/^�DP�)��y�Yx�c��x��2ǾK�}=��T�8T�m���2��J.��u�~ѿ �7 Y�!����cm�2��p0�n!-d������-h�g��$C~^#��U�6:J�dYS�5�~�s�1>����I(��育.`��L7�(��׎�uǕ�hѵݏc��|Еg�><,����������˚�����5����X��/<����?�G[�?�j�Nl�� ��v��Ӄ=���\t��,��	 ��� ��xiIZw���r�T1��;��M\a]t��O+�D��]~�~{��&�{���J�PH��P�fk����k/Q�������}x� }��k]kN����#���S5V���!s��%S	s��:�\��`sjD�R`nP3K$��DT�J�\5�S��O?�u}猐��E������{���ʋ�Ȃ�Ysp �� a��k�V_	В ؖh=>_\ �Qu8|�.41�!���>��1SHq�0���,`��.�6��k6<��}��� m@�c�� �R��j���O'zԝ
V!%������\��4)��[f��^����O�p�+��;;fm}�,<{f���YXXv�l����Y�cZ�c�/_Ƀ��{�'���m�B�N֖Mö~���ioG����<�y�ӷS2 ߈�U�4�q����Ҭ���y�5<?�t�@�7�}8�Օ�(^���d[d��,f��� :�_b���R 4�/��L
�p`��4�%��RTT.51��P첼xqt�`g�����)h��}9|�,G{���u?|7���A�$~��Ӄ$�����S����
�A�R|-�+-��l�� �SS��Q��Ely$����8u��3~���ӏ�����5��H�Y1���"���Z������Ҭ�Ҫ����0�u�'������6�~���/_�bFF��|5K��K�hj����WQF+�.P$'�r���̛��ku��c���&���%s5��X� �a�`�ڝh��F���������k�˳�pݐ��|���k�딽���(Å����Y���nuW��*g�l8�v�R���Ep�D���S'5�<�O?��3�Es�s|w7�X�@:�g�� 3��zi�����*�)�`sy�"����龃�9 �7��H0л+����Tz��>#0�9��͌��N���'�~���e�,�|�>с�����h�Qh���"H��j]�\�)�{�&��':����Ƀ�x&��7���Y �z銒TG]�cb��o�k�Ȝ$I���@�MK����J��"��x�Y�!X����?	��ּ���ե�3Y�����Y��cα�pn诲�"mX�z���?h���y<$��bq$���Ɓ��o��6�7���C��1���`B=�&�gc���cwN
62"���OҼ�D���-I��0���8#0F��|�c˶Lp�=�%�|�+�.i��xR0�\x���EsX��x}ٌ~{��}M�l-IBQ$��M�~�D�j< 1��p�,�Z!�S�TӜoc�ey�@�w�|�l#z}�0g	0aB��V�"�홨p���>γ8����1
-��6H����������g�~*��K������W�k�"�284$2�q���`���[�)m��C���sV��'���?�\*`F������'��*��-9\A�H�O���P�Tc��ǧ~7����ۣ6�.S8��ӳ����w����fΝ;�_�}�C�)�T�g�?�}�MLaQ��R�3Ȑ��������g�����B�}����;�Lꪡ�+b(�� i� o|�pVue]�=gP�}�2Wz�~3L�����7��JC! ��_��,��NS�"x��ܹc.�?��}�ޏfue�����0���H���8a��m����L�����%l�o��c����0��C�"8G�a�@�|VR��a<���K^t{?j6�8���tÑ;ތ�}m﷿�c�����	GM��"`���ڥ,zl��<����ډ<M�\*6���0���z��)�/���ܾ}�2Eµ���ɏ��3�Ŀ�f�O�pjw�h����T��pZq�a�,�׋�\� �X�ZJ��]319e��ϛ�W.�E����E�^=5>2�������d!(<48$��j�>E��|�wVxXK����R��"z�g026F�*�� U[-f���/:c`��A��J�	���!����k #�G�6��	$�|���5342f����_�b���+2�=��\��O�_�9��R
�lK�\�T@�s6�������9��E�2ư=�����Y~��kC��gO��'O����Ej+æHM�T�۰^ ����p���`G|I��͋�\2� IF"Y���������nϻH����@t��ѿ�	[�-w���)����{�k[�*�^�\��,�������b�H���_��9a;a�dЍ2j�����L֤$2�J��$cL
���2�(���U ��RB�^�d+��������s��"�0����q��y��"��k�>YWS%
E;�|�����Nؽ��=���J�n���1��;ci M8_*�Y�+�?�уj��L�S�1j}�$D�l��]d���;Ž��V�������W������6t��Z	Yx@������̔�aK}`sFMt9���%II'	�{S��)��Ǎ��m�ә�.\��ɤ��T�OR4K,JG	���۷?C�u�A�`N�F�-�������A��¯���N�a^�RB�X��^#ӹs�p���S	"�pƼ�=�I�[�����Dh.߸q�<{�@px��k�.�
�.��1�R@͒���9�r���qLbrPØ(�,w>����ݭ�|����)v/�I��I7IB�S�� �!N�0�!!108Li!�*W�^57o�d�r��s���!�����!�$̵I���ͻ\�V��m�l8��s_����^�|��w����n����A���͵���\[[�ùO���ns��� �yw��dIe�5�z~���~�8�3t�| �9��;+����?�W�,�c��|�O���`#��Elr)�(�L)M�4�������������&�� ���&s' +�-ۧ�[`�۶٢:+��c w���3�Q�g���=ǎCl;yGſ
�W�!��G��NI�lێ��>^���m��>�l�d���Q �c+t�[u���6i�>��ր	U&8��/h{�� �d�LMJھ�?�U�Y�h>P����&ڐy/�{M���c5kN�)>�~���I'�o�в��n:
�)���(-$$V�U�;��b��X(�g��G͍���?�`����i�=]0/^,�￿ǵw��㒙���0�#"�722n��C��g�90��b�k��!�s��pIy��]�	�׃���B0���NfE@ڬ!ΰ� ����dGȸy���9�~�}m6~�����q6�S�s!�29c¶��1����[��`7��n���54)��so�Z�e4(�9�q �E����+5��YZz�l-�1�)��%:���c��z#�a��#ή�zШ��s��T�KGJ��)2Y �]�+ n\l]�ph�Y�4捲(�}f��+�?0���8 �+W.�Ϝmu��%��*P�x���go��l3>H^���~���=KJm����ʲ����<���>�	u���C�	���Y��V}�P��T���L>�����S��!�3�l,<���PQ�X���ໆ/���~3j�y��]k :�?C���vls�E�u	���FX�˝���;�W�w�2��7�����K3��@�0�0NSu�l��0<���9�����tK	��>xp��Qm-�|��9��J&�7 fg���4�:�����eX��K�nW �M���<x9�9�H*��%�=d�`��~{'[Pٿ��C@��y�� '>�\R� ��
4
�$<x�PS���3'sH�_E�M�����!/��?��!�UR
�u�qj�)�(�� y+Z���gB�4��aA�R����S?%uq�\�r�z�W��4ݵ��C����&�@X�'e��������N=D8 �y�!B�h_\��h-���ms�fV_�?dB0��d��	��2nH�:h&�����*�pD�ܼu�||�c���QM��3Y���FA��Y"F$�����(A����lŞs�7���:��_./��w��>66a&'�ݹM�X�-�w�����zC4�����F���C��Y� �؆�bֆ{���V����7����'������+4۹&���Iϧ�9�S�&?&"����	��є�HW�^㳊qfX� �<#/�R��[^�v�)���<��0�ߋ<6r��1�c����s/f�u�R=Y%�}�;>� *�\���6�o��+��q̱q���s����N��m�6h�R��3�-H`������,"Ž�J��[8��)��&��9Y�G�k:M\���zx���\>�ٷ�	C���-�	�� -�=��b||����Y�6�3�淿���� Ʌ������P�wd�v��� ��Q<wrr�LL���s��w�A':�LҾ�ZɠDfe�k���Z+ �< RB; (^�����`2� �A��`mj@�V�����-��F�'�������۷n��l����c!e���m�l�Lq�l����j�
�`y��YX\`�P�S�?��s}�9
��g��[,̷��f̓��/4m���s��b㈍`i�X�Y�%ES��מ�/�F`}�=H�I0:� ��#
��>Þ�5*��;T�'!}� �R�
��� -�[��_�N}S/��K`�:��o���[�����ZGw���8�}���^��L�qj�K���*�wc�]��U/4�G���{+�׾�q��Q��wTF{�儑K������%B�ZѨ��B��=!Y��ixS�h��#*�vl��a��Y4 =0Nv�&�9L.0z^�~;I4B�*f������
x)��(n�Y5�ʌ��̩���C�o��~4�2�C���j��$,蔜h*#k 1�Q(�  �\�^|�R	@��"S�*�*jp��p<,h������W�聅�!3Y�5�Χ:k(�Б	A$F�knN��ubi�^;�H��S�9N@t�M����g�~�":����kt� �K:%p� B$�¾���ݻ���̓�ڊ�����O�*�D�\�hײ8�*��H�Lu�q��#�o�`ZxԳ���1����x���oKi��`�Q�	]C^��G���1!�_� SIs���c	�f�8'ʮC���g�_��_)��$�ڵ��J����Q£� X= ����O����ܠ�RM���RK'��x<0��i��,F��)�< ����0f�(�礙5UY$`���S�������2��+d�W+�f��#��rY��2NS�-�y��7<�5@M.+�˘�{ǻ�vmA�[����h�o��BQT�S��Q�<���r_��4�A�G���h�kEǑC ���Gk>Д�R�5̛`)�B�d����qGa3�G5S25����ʌ��jp�0W~�L�C��&~�=�c��!�(�Pn��܂���݃~�	�uld�,��"3��������{�h��ӭ[7�G�.w}͚�KKnL=5�篰Xj 3c�L�ępRQ \|��i�O#���Q�p�k�k��8�j|{g{��-�(2r+�p��/�\-WBQ���a!_�o����Z}E+��v��fp�r�6�<}���<5�{��{	Rx�^�|)�"J�/o������/�m<�a`���P���zpl0��̡O�,�>���e G]�D%���C�u�6TI��KΎ}����g��<q��E�7�"��D�Mj��%�i�"�"�891�b��T��6�_l=8.�T%.�]�~��Z����y�=���N�������og�޻&�8�`&'A�׸a��X�������$O�&��@þ���鼇1=�!��9j�"6[��	��)���U�X�$��uI�����砈w��Z=j�Ѳ�������[����7��r�Y9~E����Ġ��ă�8W ��ϊ��,v�����s�����H~��!�M�L�R�! ��D�Y ����c���o�^�RD���MMA� *@+a�*�lU����z�
@1}z��8F ���K�����=�#��1L�h/��Ch�X�b��1W._2w>��Z�p�^��2�lܕ���õ��2[�z �y�|����a$�S�\Y��"i�`�N�O�)��)�:=;�J�p� �����e5)��A��ǋ�|1؈9-�F�T����i6�h:�k�|��W櫯�5��b_��M�>�P��ի�g���T3�ҡ�#��О�w-a��sd�ל}�U� ��A�w��i�;2:�k��H��c����A2V��y����r,U��
���F�Y_�s�0w�AR�ݳZs�]��Po!����h��̆/w"��ަ<S��L�4���=R���v����O�~���"�=��{��{��[t�롷�z�Y����1l���L��	���9��Y�tu2@Ҫ�(jVҞ��z 0>��^���Y����n�66^}9%ӛw.�(��2���L�t7������������h�9���O>�5�.�7�~����_�f ��o�3=13��,�1U.����k�����z�u�^8���'�À�H����Ҫ��RY�;�"��ъ[f�P�k%�e(���rI��`"��?Y�!r�;���5}��u0�����@S��I�2����ѣ�dS������:П��L��f�=�zuMj& 6���^�!��l��� �#��  +5*�`���4��ꡃ�U�"|$-d�5(ӱƀ@խ58���@�ٴs�ҥ��퀦6X� ��������hl�b}uՙG�FA��fgf�9�v�b_=�d֜����(�o��5�����g=�yk/洆J�淴��&G���#K}��f6>��+N���w[���Ӯ�H�Q��ڣ��"�qZ�J�V���� �A �l�:R��v�R�QY��$b�)���bP�y�(`�K!vbT�'����N�r���g�(�2NwƎ�������9t�Q�")�j8��0�� ��v	�(�W�����I�,B�մ�T�'Up'�q�3, ���ϔ�b?�n�����X�=,%V�k�E�օ�{U��x  nx�[�-~��c��@��&��d�^3,Z�R���RJlH�l6E�p�9�s��̝Ͽ�Ӆ�3K/�Ɉ����^o8�ǂs������ܨ�L�U�@&��a��H�v'�'&	~���6"�+�4el薼�B��Q���%a��/&^�������al�0��Y1�ϟ�?������OL}71c��ԧl����j����N"�1��=�s�>������ס�a)�"��[(wT�O:Z�\�e'���[����g��_�ې�x?��lT���5,�"��@r*��1���>�<:-y�>��c�	<�="�ャM��a͎ �T�J����oM��1��6�Q���5����c��c�o����bk{_��|G��޾��k�DnG!K *�{z��L_��mmE{)���޾u��`j64VQP��3۽Ob�h��[�&�x�ߡvz�7c��^H0dQ���+A(`��F��`���nJ1��Ѫ��jn�b]0z��7�~C0u��K�0�h�_8�W�)��u7��^̐hЖ*��R'�HAd �U�S��l5�)�N��A�5�5�)*B,Ez1 ���PDL��,i-J�5Z�Rn+���n^��>���F��m|�c��9�ց��Ԡx��d��=�ِk�f{y/��E2B����fc��d_|���7.˃�xVq,����vUo��Y` 
�܇d ,�t��k���c L���6���E��y�Z� aFqU�3�L(n}m�ş~���u�&7��6�S�����~mS��>�)�o�'6�Ta�����������g�=�%�!��f5�G�c��,8d�uaV =�3~`)�"o�!���Y��8�9o��:K��kD�"�v G�r�5�	��H�˚~_��|�T���T��s�Ć�3��$0�r��~�Sn�Q�r��m-~��vHO=�O L8�dڤ���{������(c���P  �,�T
%���:1�>�g�4��P�+��I��/M3�L#+��ǖs��R�N��kZ�O�TIW�~�/J�ʊ����*�! �/_ֵ{�EvF����4�0����jȃ��Cq8<�6s���?�ò�#�b����\^~e^-��U�a�����;��L8fA��5�ȓ�����W�����T�T��)�j��Zp*��ʀ�H���?PҦ{��%2Tϑ�r*�(��B ���|k��?��ܻ���v�ܾ}��ƛwB�
��a�\�]�K��o~����Ρ��"�_��c���Ƨo�2{�G �{~,c�3��^��?�/�k-�Q�N��G�8H���GժRX<�.2'33��?������?�t��������h���� �J�$��*��rd�Wc�"��33��j�C���Q�;������n��@��A�a<p~P9�����x�Aa��V�_k��{!�hm����m�we\U������y�/���ܺ}���.�ȂHJG�Y|�z|vvI��_p�p��0�4
Z�D�)a��ݦN�+����TA���)��as��O����w�߾���|�g���#���$��x�ܾ�1�-�2��ϝ;��j.;��!+��\�U8} ���s>��>�,ᑖ�fjR2�u$dm��$�[��Cqf�̡Ps��wͬ�g���i? h�1��^>��.PP��M0a  �_��!؍�v��k��Y]Y!@������B��2d#�zs�J[�/���(E�)
ؑr�|��X�!�"	��܄0a�xmc���z�]�K�������DǫW�fkk��8��p�����x<%,�W7{�H�AB�O>1�|z�����6����k2�ʅ"�]�j��~{�Z�k).n�d�o/�FdqM��g��o�f�`�v}��2*P�xRmHJq�N�C��Z
���L��6����Z���"�����ȶ~�C/w�|�3k�:���P�}�bS0�`h�믨�S�T0�����o�i�%�]����j�Qi˲�'�nʚ������r�!k{��ٞ�f}��ͷ#������
.��\�1����.��п
����:"�I�by���{	7�N� ���x&�7�I��{H��7��CVrW��י�
Yh��b+�c#P��Zlt���h��|���i-�s�eA�9���/�el(���+RQ!���b�x�й�88�#�f�9Np���ܝ���5�0(ڇ_��\FI�Ԕ��ƾ��<4���9^�ڦ��2����}�}�D���\���p���`e�,�D���e�xG.��d�� T��_S����J����AY���g�W���_}c���?̏?>t}3`FF&�܎b?-:�8w�ME�������*��A���͛f~~���yD�
`�io��ԯ�Z�C� ����}� .���y* w]�)��؇���z&�l��o��^��30�x�؂�ɭ[�D�ϭ� 4b`�\Q}�<��(��g�5��j� <kv�1P�������k쎥�{���W�Up����]��#h�� ��9�,��w�����߃@�}���z���;��cN�""@�&|�rNF&���Y��	tݯ]�nn޺I�U�%%*�@Y��.��5ꧬ�#���6��x7Z�i�8שk��fw�\*��F���|�lvw�ftl�Dk1_a�U���cp�K����g��3������y���y���k4����G����m����ư�Hd�Z� +�%�0�`��l'w�6dI9��"��F组El5؛�Ł� 6���.Ac/��`0�@� ��ZvJNTNb���:�����u�x� |��&�Zs�=Xΰ��zM�|��_����*R<��J�ؒ8_�՞HD�������j���A�W�kB�$�kȁ@�m�H�
���Zm6Hh1����v�Z�R��K��\w���/d�AB�ʕ���+�~�O��\�Zs�������.��l�S���5YPG"��=􇵝�m�vVu�:��+ͯ���{B��W�*,�b>+��Ԧ�=��s��=Q���a�������I���+c�����%:�-� 
�3q�nhdv�������l��)n���ܺˑ����<�NgȚ��	@"�II5�$u*�yX���'jsy��RqX�	�r����KZ�M##m𜼄2������e�!�w�=���iY��8�D`����+��v,��>�t;0k���Y �s3��e��R۾���m|6E���Vߓ}���`Qa����36��a��)���C2n}�� �b΢�� )�	B�W.��Z� �T�`��|��|�[V�֨T�\s�-�.��Y�&!�Ka	��p8(���ann��-F��p��NI��s�6i !Ւ Z"�G�i���S��;SSf��R<78!e8l7g�b��)&2e���F��+�gMP1����נH��m��I�ݔ@��k�)��� ��ɓ����/��y���ۭSpxh�9�u�k���

��sd��r�����ӿ��K35=�m�/Q��h�� ��$m>x�V��XNU������g.���y��fa���Ϟ�e_�wj*3�Q44�Zx�K���8�=O5[�'�&�x �,�H�U���l-��uj� �������&�Gk �ϛ�l=�x�5���A���>��u����M���ף8�!dM������Pב��8��� *k*m�3�}�;�5���\���dV}�����8��Fe�=3=���^/t]ecP9LA� 7��]?�D��1�{��Q���0DNj�:�ɼ �K̜YYym��6�$�� �k�5�T1�m�����̕�����3w�|f._�l���a�ݻk����KЅ/��������̴�8�dLxMo�äV��g�l�lI�cY���冒fJ/�v@��\�[�K*���%�m��A�I7�����3 &1�j �y�P ����H���`_����Ō!�����t6���8m%|�������]�E�@&��+319a�ݚ�����y�5ط�J�C��s�����>`c1��Hf����Q<��@mP�n��knlR��@�;>�=g�q��Q����MI�_����wg{���I�@�cnn���|~�̹{��5�Ae���-e�s�^;`n5^>��X���m�eg�7�:���p��>�$�~;I{�r�n?x�W��S�}6E�dn.����(��p�|�m-��1/挾b{�wRV{��?��� ���N���t��
�4�y�ux`=ВENG7:K`ٽ�>ޘ�(�F\�Ex�ӆ4��0U���Z-��G����Ȫy��F�K��]� ܂��σ�Gm@�3�����v�ъɩ���
l�~�_���a��1�Q4,�q. � ���t�N(�<�Q!�u>s��͛����4������3)l�,���v6z6����~C� i�����ح�F�i((�9'��+�����Cz�Ra��M�98J �0�Yü��:S��n��1���\30\P��慁�<9��;8 �	n�I�Acc��T�eಢ5о���i�H�M�i�]{.��Eo�.�rES��IV���+������d'���/?�7K/^2h�� +�z�n/͖���ܘ�\�^����2�q�\�v�N��Z�6W�Aң��m�����܇nm>�=%��|���of����?vJ�\�s�`2%-4k �3
i���;37;g���[j�����Z���	&��D320����T�U�&�1�-ػ�]�-g�xUy��8}��>���r'Y��^�
�y���k
�	�Ӿ�}������j6C9~�jb;d� ���kׯ��>�<kjԸGЃ:�t�^KӾ��H�v�m���L8ּ�'��h̜*�(��bGAX�2(G��Ȉdp1=�߿�����+��c������{���g�޿}�7��O?���s��%j{�D-�� Z'&&��5�χ�R��p�02:J�y��3��{�� �Z5����Mͼ@���eHn��-���HTj�~�{�/�:�-u���Cm��a���y���8v�a����y���[�_P�>a�D8l�ٹY����S�hO͉,q�ɋ־�7����YZ�:��h湻�Rh��F�
��/Xd��+���@��2�@�����c��B���(]���q��?�?j[ܾ�	��Q �/�Y�}W� U��#\�G��|����e~�I�4ͺw󎾅�}=T;_
~�0�����a��ٴ Xno^0IvAE
��
蹁��xFG�*x���/�Ul�D�Â�d�k�e�6�}4�@o��gi�I�y%���Y+L%��{�P C	>"� ��d��X���Hr���~{�Z���z�Y�t���Fu��������p:d� ��& �K/:������~�4����)��܍9�4VM�6Y�ʔy +LG�:g�f]���h�4�p�E��r��i�p����c	gN�K7�@�s��¢fJ�	�<��\�(AK�JU�� p ؀sR$�.sP�_X!�����������Z/�����1��v�|rκf���7���U��s(�=���j����BG��:�H8�B�y�.�*���9�<��?������ ��ņ�e�\����y+bRx������n��A�X��4\� .ﳿ.i��S�t��i�8��F�+>+��L�FC5���|�̀�����33��X�`2�F���������M� ��f;�~G��֕�D��õ������$6���S��zO������{P2�R�f��j���0�`~�j�sJ9)�:�ota�,��)��X>��>¾�v�[{��j1�R�Y����z�·�:�/KQ����-Y��n�t����s��es��]��?�Eg,--�����k��^|`}��$�vw�y�n(f�wl�+�XkD�k'�/f0�a�3�ŉ+(Rd���<��-��ω��~�d�������PԯL���Qp��+wMX���kK�����R��dj��P�,|�o� 4� ��eEZ���\Z�I1Ӧb�j���hA�kT4�,�c����5���������vk��b���L�zv2�}�jX`��v횛OnQWz� ʅLe���-��)��G�n�e�|�&�i̹�?۞R���������P����=n����>��=��~��!<4+Ƴ)��B��3���;|�MM�.�� H�o�|��=0 E�L?,��<ë���qjw�����O���eg m��qjc�w�_BШ��ǥ������z��G�]=��e�V���tDY�TdN�T���Έ��g��a#���ݻ?l�a��^*7�60X�k���NCA���ަ@5ˍ��lYj敥��yö�Z��%�̀�Zaf�n6����\1А���=31>�Tͥ�tH���x��5�6�_�:��BK�ejv�7��ںs0W� �"�p�踦�Q��|��H�E9���)���o��ZQp����2��Tچ�rhx�p������=���_������9�M��/^��FM�x�e����p�Р����s}��������s��/l��H)X�Ji��r�i�c�6Růײ����8�,F�Ϣ�K����?��}��@��P�P90��ɝ���r�p(������O�<�pzz��G>�}&�����r?>PV�k�qvv@L��aܛ�OB�J�Ft
o�J�8�|2)D9��^��0u����gw̧�~�ty�hOCFGq��̾�{�� ;ȿ�y��X�F����l��Z�Z��Fq^�Tpv@�u��g��_���7��,F*Z(��s~v��ݗ�1K/�̿�˿�����橿P"���'O	d"Pvk�&3��"}!�j!��, �Ȑ���.�=�S�+�5����1
�hQxo�R3� @^ �`?à�v�k�M�̡�l���p�767���l�l����
p����g��`D�?�/�N��a�a�(�R��/֪��p>e%�5��%�`g���B�aH�i��+�۰��e��V�<[x��`�@F	�l7H�������*琑�a���0�;{��an|���?���������vI�[�d
�:���}k}X�TZ̗1��dB�M����)}σ�8������[��~�Gn�4L�����f���~*1�L�M?�w��6�4���E�b�Z/�vvv��hm!U��ݻfrb28��(�7ZR1�Mú���X� F�2�N��LF��	�_�������L[���M���S#|�����?���4����^8,�Z�8r�.��gU���k������K���T銤LRs5�B�h��Y�_Ȱ�Γ)+�(9n���U�^�Fi2����UF�(�-8; bvY�������L�_�VZb�Da�����u��X��b��_��r�a�`��~��/����|�ͷ��/���*Y@ ���%U)��H8�$!ӊ,*�hP���G��g�Q{2��Fc��Rnc([?>�*S6y��?�����B�Ў��yJ��}��'m��u�����4o#�~�*��c
�=����;x�-,P"��|zbY�D��5wCX��6��y���P ��A:Fb�zG�ۥ6��{/�E���OjN��~�*J����R��D�V`�B?�ҥ��������K�&��P��ȇ7ݳr�9p
:��E�w�d��]�=��
Y�]��.7����e�vOX�+�+\�0�h0#;s�[ �} D����g���̽$ky}}ÍGK0����Sr�^����JH5��b�с��^���knU���w������!P�l0�Cq;��"e���nH����O�>3O�<!���D�B��X�ݥ����Չ	�!�3I��ݫS�E}�_,�����f���畚�<
z���D�63Y�UJ�ܸ�Qx���Ʊ_���%�5 ����y�j��� �6�B���x�C��o�[.\�`�^�&���q_��T:{��D�-��z�[b>��I2��mtR��~�õ>��A����~o�	&n�������[��(կlV�\��ɽ~  ������Ɵ��9����0`#�ҷ�F�w�F`�������}N�ʊL2����-����QY�~^�tl�<x��N���3g���m6%���+}'|_��un��ao�B!�,f%d��L�-��b��JYSH��B����i�
�B��LsP�)��Q\�u�Bcpv^��6;ۻtT�b��G�`� �)���� ��#�7�4�3�{���Q�H��V$�Au��c��:g�O�
�ý����ڤ����a�-<6�}�7s��}�(�&� �o�\U��>Q��;�/p��'�Λ۷oQ����2�S5�nH��a/p���{"���s4�<�n�|�$p�>{�S�9pN��֣�x�Z�m1;Z��~�z�9���fSy	�� d@~����I����}P���T��xs�%�is����E-Oֲ���dn��Q��eG��9����"��+W%���z���E�1  1P�T5�ݜ3?7g.\�HP�
������%Q03���2�z]CQ!������0���d�g���2�f�ʮ����>���QY?�d���
�ӯS����G��1?cb\�{kU׻z�
5�a����$��f�������!E�D�Y�!P;>>j��\w��9�=�M�Yd-��� ���~�� ��/�m�Ao��(��� ^[7���	��=\�������%��(l:2:�,e����wC�D����I��sd�l�n�\�������-�X+���#8GJb�-�+�j���(�wVWV؇"�1c.:{�O`[CZ�27x�`Z����4��� T�D���ׯ]7�ϟ3��. ر�r�����V����ٛy��ٖ�H���[��<�1�Ć��k��8�B�o�h}`-�x�r�;7:�3���s?�_)|&��>�^��ű�lb�Iu�)N^H����}�=5=���Px�;���o'n������Go6������q����R��o��P8�ee�٣���u�R����������}o>xHg�L�S����8�b���'+{.Q��@,��65��2+~W	6�UW�k�z�w�Kl��(RTEwXH��M)��A3�W�/��(��r�9�(�2I�`a�L��3b�z�xe`�$8�V���{�Rs>Sg,%8��x
`�Z+wDB�J,��( ("�!o��IC���iu���j^�\6O/8'z���+�鋥��p]LQ7Ш4�$uT}w׿��I�Ù�Ys��M�O��O��PCw�D�U��L>L1�}eb�E-y�+�h�I>>h�����	bJƁ/$��A�_2����)����n2e|�=ov<|����MaM� I-����:�j%*m�T�������<�p� �6��,�U�Z#���.��usʗ�%� 0�7	:풹��Y�/fǲg6?�`ԕ�����?� *�+i����w��F��N�^����aS`ݞp�l�7oǠ8H* k���+��p��: � �g�g̅sY�oͭ� �/�\�-�Bwk��c�ϋ�fyaY�FS��}���֭[\k��C�}���u��B��X7�ĕ��a�̷n~ki|��{��zĸ�	HU1P=6.�"ZP�,�?�n�k�`O����$� ����K6r�Y&u�� �Y�r��G�E#��lA����I6����\G��� ��n�`~cm�Z�V7OM͘ёqwk���+�s��d/��	 / O=��97�����b� H��~,3h.���x@�:�)�F�����Z;:SY���|��Cʧ�r��H4�I��ƫ��os0���Z�������?���#�����P������ͦT�'�������A��
�|p�_Y��S.�>�F~+kj��r�l*�p��/{td��3p��q�V��Â��˞��d�]��@0̃�\����H��NS-�R�)�wW�� ���)���fF(�5��|����S��A@��S�~���"ȝ�^��e��@'q�&�����([�Ag�''TR���4�<ͻg�}��F��A�Tk
������g~�w��������U:dCCfp`���k�N	T������f�0�ǵ����w>7�n�b@�%�!8�^C���X�´?:Ga�e��k�!���ܯ���oP<`��h��9��[�6���X�Y�t5�x�cA���K�D�\�p���G�@��ȱe%CB��$���O��{;P��B߮���Z��E�ƃ�gq�FW�>���:��޸q�\�z�ܸy��)���^j�P%|������q��x��yp���h�F���Gg<������i�R`�gjO d��;�P��>}[�d��t6$/0�P�o��A������߾%�:�S�X?|�9�H�5�k��ֶ����9�@�bɆ�Y�VЏY[3���"��ui��E��b��?���]���l��Y���8Ue=P�(� �^�"j)��Y4��Ͷ�  �$�������Ԁ���#�ʘn�� ����8����s�Q*�,�[H���D���̝;��s�Λg�(1����y�:��%[ >����u�+`:_�|����y�e{I���ˊ�T.������K�{&�m��dv=w��B�ǆ���2�ܷN{����v���?��9��,0F ~�Q7P��)���o��@"~Up9����r���� ��LCBp���*��)?8
`������8(t��{�޽YHN�ή0\=h�ٸ*u7S"S#����x%H}��"R��g�.��d:
<��4����p���������S�06H�ĵ��v� Y�U:�`%��6A��R�e�&1c�)2��N+��:�z~@�S�'�1� �R6 �y�[�I�;����8[ �WV��ӧ�̟���o�3�>�5�	D�w��Qp�A�_*�vF�;e!����T�N.����vE{0�f��.�D�v� P[��;U��n�����Wn>8��}?K���Q��L���L��Z[�(��?J|�q�1a+H3o����8/�}<h&�&Y�	�2�x����1_e�cN9�� �P7�m/&���W������eǟ�� ���l(@$E@gf�͗_|I��C1gywIU0�]��S�x̰)yza�L�aT���axx��q�Nz�#��:�P'��+%�*0,FP�
���������667� ��/^����w�}O&�[ܞ��v���JHF h�g�6P�� `�cٍa0�Q���y"�ºM���%eSo�yoRd+TO���//��:�dds��K��n��ZW�U��}� 7�E���6�l��Z�N��~6�����8ǲ��a[ ��k�����d����#C<�����k��Q�Y�'0���F��y�Z~��l�]ʑ����mmo��狮χ�&�-+@\��Uf��1P���ss��# �q��6���%��>/k�3-�����y��ͷ�����-��~{ZV>R�M��3�2�L�B�!�,@K�~_��i�>������㬖+HwBa�V�`Z�����N�e
������!�z�����0K�l�֩ �RD	�0��D*�{6
�%pn:�`�:(r���y��u0a��j��ݢ3�~zެ��1v��v����xmQ��V��.r�@�Yi2M�V�@�1�U�d�<�$�K�@T:wΡ$��7 �8t8����� �0;;-Ł�>h6]�a�)ΰ ��L��a0�D�yD�ݧ�)~]�9N��݆�ME��p��A68��NFF���j.z�RuD�[�)m:�,��e6�V3#��pX������/>'�}�P�f��w�S*(��@#�#Nsp��"��-�L��{9�Y�/f �}!�Qg�]��)�/H���	�c�'=�@�����x�4�Hk~������9��}^*�4=�&����l�i���}����L��4����F+�ASL-�����Zr��Ms��΍�66$���>44(�f�<U�# r�Z�}hw�1���x�w��6K�@Vy/Gc.�K\�P��D���K���c����f�_�p�~��7\+=�l^ �������F�eg�}0�=��@
l��@��L�G�����~��ٽ��ˤ0�*���`*�#4��V$����\u�"��!)����8�l�6�@����kd�ϔ���je~g�(ըF���x&��	RAA�%�~��FF]�mJX@��y��ː�,�4>1F6
&���s��!�v����y�J�]Ο�7|�����ڶ�6)�W�iZ
2��������/�lð�2!{�z��&�q�c����>��㷈�����f��Y��;�o	��߿�v��,�۩7�6;CA��6;��~�Sod\F;�RZ(hw�V��zl�N�~N�'f�*��h�Y�ĐM����#S���q���S�T�63�y\�p.H�v��E慄2`��Z�d�d!��e�q/�VL'@U�e�?���Yi�����7�V
ɀ1��Aa��v���O�p#���׈_�geubP<Ot�EzDX�`5�N��ZS�A�aG}�_�I#�hO*����/� ���3�=6�WV���������5�-� �Q����ys��s�㏩9	�S4��cYz�+�+wa�v��؉��)��_�����|����c;���r��m��Y�����a�HIOT���~�(�M�T�㹹9:�^�XZ"{,8fԛ�G�rT&T!�u������[`��h�٦�+6*�w�v$�lӅ��߁8��	�<h�c��B�5�)(ʇbh�MjaG�d�={��ɳ2b'v�sh�t�WY4Z;�=|�׳wVM���u�w-�p٭�5�"��d0[�����M�"Xy����52p1�/,,J��J%0u0��͓鋹�#� �%�3�����"@�( ���L5�`�;[��� ����v1�����p��iKT��C���od&�5Lɖ��� ��?a+�s|�X���`.t����U�B䊌ʅ���d�����U��!`z���,�gx��B��m��/�̮�������)����93;C �K�2���5�(�z��UJ_@@2��ѝ'��$"x=f! �|��z۸��ړ�=���_q�A�U�o^�E��F6�0�V�^���v�,���� �U�n5�1T�p��lZH7?\�����F�`� �E�4��ca��wu ��4XŻ)F�M�x�<G����y��?���E�1�J����i)f@ݼ�f\����ݧ�㜼C}��h$��B��2dI��ý�r)+��w�ZI����VV؟Q�B8�^�N#�P�(�lñ��`Y�r�`j���Qb��)3�I9���+��HV$�;8nt�Z��`[]}i֝S��-� *���/��O��1W���p��������y��)��]�Tq�۰�}����/�V�^a���E�}oN#�OBA����2{��|l�1ul�
-�ñ�;��'�>�ܩ#���Eg�N?  ��IDAT��SϠ���%�x5~G�9��J�=k�����J& ��x�"_ �?zb~��Yz�D ��dU
9Y��>YD�p�A��qSv��)?����Ѝ�v`:�;>��w�3�z�)�����0oz}���q/�y�&�̨��K�TΫ
ҵ�ن�;?�}�����/~m;����woY�f�_��}q���UI��fK$fzz�A�//_�d��ݻ�X�v`p� '�����$K���֭����ys��y�`���W����xjr��Z����@��t�C�`�N�'���5�I�9���%$��P 2���X�k�3=��g6���:�5pmu����~�[�U �"+k�=����ϗ^����`�!�733� 6����"��t���HF��4����3f��9���`�@���P,s�+dsmlnЮ�i��0�,r$�� ��<N��{�������FVAP���[Z@��r"vK3"��0hÒ`i���*=ǟ{�����L����>�|��3���,y�V��U��}�������h��F�����CM��ʎ����?"��«*�ۯ޺1��պ�zr�8�L���![�u���K�]b5���,h�5�u�(Z�tD�0>z��9+d�x6�Oɝzj:g�c�P#0�d��";i�̠i}�Rt��ġF2�Oj�U%�şl��=���:�#����	����ҍ�u:DpJ�VY����*�_]Yft��ア2�*�ߵ�&�"���R�WV^S^�ʕ����fv�0��y�l`85 ���a�3��RDQ�����e�ʽ��������,/�Hᡬd&�g%�&d"7�Z)�TQ��H�&������OY��ʕ+f�9��p�@�>w�uZ �NM�]�+Π� ���@��m�HG�p'_;�E l�Ȅ�lLxλ��l��Y
 [��]�"�"��RMΔ�>�t����2��9 �uP�%�^HՖt�$d5x}li���������*�]����~9�1{t :�Q���p�(�÷���g�kM�g��>�1���>��>��-@���p;��; M�N���=�}�>���/dQ�P����������ۇ��;z���y 숆��އv�L�S?f��Fw�P�S���h��U���8��CF��q�\�B�2���޻G��ʕ����I��q����'`%C�axx����/��F*�x(847lj���ܺ��l�����L즻���)�}��i��DF��;7��3�%/��Jq�a�/]b�u3`�TX�:
���je�6��;w�~펻��g2�s!p���� ޴�!|�t��A��l*Z8��>G�BO_lOC }_;[楳oD���f�̟�7������$5 ���o�2����)��^���}!�ʛwOSfG��a8�o�n�-��4O�Bo%�&A
h��k������	I���- ����>�|`;��R���: 5�Z���/��og�����d1b��vx��g���M[qTJ���2��41>G4��heb{�0� :�ŀ~೧��` M�u`1'IIY�r�D�TA�,X�������&SԻHl�ʚ����=윽F#1�R#��Kg���m(j�Q������f�-[�VXu�õ ,Fj*%/�v�[Z��D���!32:¹H���ִ�Y{����СF
?+��}c�B����R�x�9xHEM�)0����4�����@>^��Sʳ�Kz�R�<g{���f�0�+d'MOϲP�'�|�T���t�L,PX*���m��2k��96c(f/����Q�����)�	]�� ��u,�s��u�36�� k%̉�ˉI�u�!�`E�f��0� �y���t�ՕU2��L2�TU쳔aʲ����.�kQ��*;�1����N��5�3��Oh�xnp�B�{�׊D*��tr��Y�˅Q9<2JPy~n���3�d,s�^6 ���aN.8��c`��h���� ��ȃz����:�캗��� :o}�9��9d��d5�@�) �j}��T&	C�����h��v��D}�Du�WWW8a�B0/ ��٨`E ���w� �Ұ�4=5e���)���g�	h�$j�i�=�|�4���~�Z�X4��Ɛ�s�������%�wff�v�Lk���rI�N�L�+W�r;��iw8� 2 x �v6�=  Ԝ�2\fa��� A�����)�{��Su׋�Ԧݳ�l����Le/F����/]�d.;��}k�"K��r aN�$�M�XdHd� �Y�ّ�>꾏�굯w���`n˞M˽��h�vpm�u�=!������K��a�~;^���vf��D���~;�_�yǶ�W�����#b����@L��+}k�D+C1�Rn�������˗���y��{�.�"� �P ����� �v?��H�`rH�O}����A�ħރ��&u�N���5Vkrp���舀5���JƩ�Wdi���p�R����v�L��O���p�]��448d��%uL=���~�J��OկTj,F���@��������)�El�Pv/��p�2x���#���Pnnn�9�&���JE�`��bS+���A��]��ߑ�
�����ɧ���kR������ttG�G�1ƺ��=���g����aځ��nR>m@��3���b�Y�jl8%ĵRe����Gݭ3e�X��v��˿��E��B �A
����!-��+f{�n�F�~�þ��~yg'�
���XBߙ�Q�X�9�����#%��lrs��Ȅt��OP���ի��`6Y�E@�i����1Q��Ė���b��K#yظ���;���b����B�J�y}�#Z���6)8) lZ����M7�}�w@,d ZZ$�Halnn���s�e��F�xӭ��k��s��.�+��h���� ����WYm ��A�U���366n����a�����|��?�c�	pW�����أBuS����� ��hH�cR��={ dgf�ݳy��5��0��Ƙ������m�� ˿��ks��=��ͷ�����_>_f������`o$�:��bd+�3�ꁛ���Z�{�Y/v_���U�vH��s�ܼ���덛7\�~De��Rtp��	��ƚJ�If[j�y�$�h�̀��<�g�,�N�*m�{Z;���ZV>nc�־)��AQL���D�[��4ZXk������QSF����@�哮�ݘ�'ܣV2� Y��hs|�$*��+�FJ=s�F0L�D���$؄�̳gd֮�o�	�pr�R�&���(7R9���@r�ec|ں��=���> $e�g>b������fkk۬oT܀M�Z���e�i�>�}+ǐ�I��q��b/����IJ�r/^,����,���:e- ��XHQp�����-w�ʶs*��a៍-��r�9r/Ȕ��E�B�B&��8�rIΛ \fyIiO���y�? �#=�B�? ��9G�� �q�;��Vʧ�t��@�����w/�����`�0lbe.��V�[90�	2�6o�1�:��3@f7�HpD�t��s<' oF�F��K����,-�0˯^qo�lqA&B�����Ir�ԳQ��ODs�#����T�N�w%0V@t�ߺd�u�����ᛨ��pN(L�ټ�O������,��� J���'�tS���g*+��f��� �.����Z༃~��  )��g+'ב�L��� *��v��hg����Z�7A6���A���ǳ-���!�鴛y+s<�s@�σ�ZhxF!�!�	��ϓS��>%@����_����?�Kន-e�b^�]��#��׈u���y��)��l�+W����ސ@��g8ב�qJXx9| @8 o|�̟�! ��-��] �&�� �#x���ߛ�������/�0C��y>z��<p/�`�tbym �Dc^�>�΁� p�@��O?1߸a�=y�9��gn�^2���0�@F�)u�rG�Νg���`x����b6��57�`.�BNB�D	?W���`*�M+�!'|>�w�Y/2����t�ô�=�yv��&�Se�6���}�~ �����r��n�}$O�;�R�ۇ������d1N�l�Z.W� �*�h�2~o�g+̴XJ�� ��R"E� ��"R�s�8Q�[I�2�8~�9S9�<� ��<��^1mك�u�;�00xY�ڬ`� ��,�d0Y���J�%5IS@���f$��m4���T�0 `�j�rIezD�>�zyYe�dh�V'o�9�8O8�Ϟ.�'RM�L����6)�#��9�O�=��S
�H� 8��L��H�B�>�F�x/ a����Dh�3�:ȝw�ŐOs���ou=��i���$\���|a����?7>��}*|� 
��X���0�,Ƿ;�=e����T3T4C�n���͔{���j��jSr&�,���/ �%|�3(p��w@� cӭ�A!}�n��(n�v��ο�Q������?
��3�$}������V+��A�ڈ�`� �䄙��a1W�᛭fJ��d%�Z����iHz�H��r&�=�h�FL�B?�|oY��x[���YZ����w�;��y���b��9����?������~�Sbǭ��&m4$[H�"���/�^���M��q�6U>omn���$�c�,kf�:@b��������9�<߃��l)h'߼y���?��Am,�q��C��7��!K�,��~����s�����>p^�[�Ԑf戛Kq2�EQ-���]0�Ao#��G̡��0��$�� �dY�80�R '`����{�Lq� %�@L�YL�F�p��RgrOe���ƛE'y�z�-e'��~����2����m�̃������C�Hz�d��÷>��o��<�J,�0��ʠ�~{k[9���ZD=�im9�����q �Э�%� ���Aq7v���Ρa�._�z�\yq���'O�Q3p���.aĕ)� �k�RV�-������4�SB@,����21mV`�Fs*�Ǯ3|���6t��U��jKq\/�>#���	 �T��`@������@8w�GN�ȒFA+T������A-���ޕ�Uwlp`�3�@�d�3
m ��.#�m�6I\�I0?qm`�qC�zT��z��SuJ�u���S�3~��:"=e1������=g'mY����_ܺ�E����ԛb.�1 TaC89M�D����]7�1��������A�O8AAQ�=�� Cn}c�s�@��� ��3�cd^�����?`��i+0^Pk\�:�A~=��S����ξ8����^�����X��m�t@�bȻa� � ������>�u�EV�HvGf8���1�
Z=��?��n,u��u�9=*Lh��U�tHzl�Q`7��\��B���	�Lf)"�4��J�g�9˂��^��)�Y��e2VVV�
j ��2���� 3�Y- ϰ{�I�%�aҀQv$��b��ܶ5399�5z�폁6e1�M�y�?c �������w�5�q���?����f{k����y���d���nk{�`�Ҹ.�z�ޏ�' m�u]�r��(���${*I���y]w�ɾ�pE����_������N����ܼ�x����<cN����>'(�r���O+kI�^��D�_S��sHv�'}��?��~ُg�"�Y�25���Y�ϗ�7�����哶3�׎��b�(����7 ,��o�s�$�r��p�,F(hc5���"�5�1�,%!L՚R�c|`3'8F�_4S��Α�h^�xI��µ�kx�p���`�h�,��Fl��,�����<��{�0�!1��� ���"�U��|��j�_[&q*R0 $��m!��Tvr���~ c�;i��u��fg�9sd �4�5S]@a;&�b��	k���IA��g{�{	G��s3��9ѤEz)�hA��q�q)tS)�
�²?x�+0�=E�%���d���?�<�n��RL4ˊ	]�Q,t�f�5f�2 ��A�8A�~�,�&Iݳ10h.]�D�K�.r�A:�ʫW+ �0����j�;� �� N�0y���O� ��y
ߋ5?=0݋�\��[���w�^�����7B 1�ZdW���ݼ159I�~n~��K��� �5^�BY�Z4���KM"��a���9hiÕY[ܮ�NX����k��,��~�7���ܯ������=�y&e0
L|����)s�F�AuHM�LϚ����^�t�2ٿ���!Cx��r� ��nf���@���Q2��P�96��C[��h��ʚ��5dԹx�����@������`6XĐ�BƇ@���y����x�IB%�R��8w��BKR�'�!�}��-3<2B������ nS�H�t��T
���'9{4'qމ�n�fv���9��2΅�T<����y���*gg4erV�ٵ>s��-Hj�Ζ�yޗ`c��]�,����x4?|�mjQ�>+���M�����Q'r��^��Iǿ�%[��3e�e&C���@�0ɋc���/�_��	��K\S:{Ϟ>3K/��5gHd"r�<V��T֡]�" 4��`O0{�L Dx'$/"H�T�KY���UűoMC��V@�$�
�E��7:]d�4�L���;u�ed���-)�%:U^6.j�S���nI��Gm��/E
D���y�������H�M�9�=�D�QJ�+�'d���)��i^���n@��ϴ�v����Z���&�,Z�.Ǆ�.��3�WḾ�_(Z��qϊO��tlc2�'&,c>��}ɬ������|�����Ӏ��>0�]H}J|Ɔ���C^6����s';����Nx��|p-�>���Θ�p-h`c.�"s�s���sff:����כ�� �1���y�b)�/�&���Pף���_)�)wy7�!I�ĸ�[*���Cl��p)>UJ�}��\)Xw��� 0������f}m�RKnށ<�ա���4���p�z�x�p[a;`��t�{�P��,�ad`{j=�J���~����������9F�;����i���.��5����`�[�R���쎦\+�:~GKI(��| ��^a`@2�:�7�x����`�$*w��ʹ�Z!g�عZ���(���~��G;������f����ͷn���������a�_�Y7�Q�2R����o�x���v���!�ԟ���4zi[�}sJ�΢yY�5e�e3/h�DɖVR�	����c���F�YndČ���K�/;Ge�,.,����-��ϗ(� @M���?��s�\�A��jLt�F����L�M�*������c81���
\��3�=0�ZF�,�W�F�:ɥr.?���P�'�i`�C��9�z]�� �=h�dTc���$���*3��������$��g�
�r�MLߔ?R�IJ�w�bݤB|@�0����߳ne����x���#����(7tqȜ;����2���̋K�����o��3�|E7�� Ƀ��J���3����P�+��́�}[������em�\�:�����y}i�!��T�I7g��L��Y�LF�:4�h��tQ�uw��* ���ka�ϳC�����`7b�������ԡ�f��¶m{���eo���j����Q�#/$'�D��������A�$y�Z[���{�.�qd;�@�X3#�2�����޼3RK�4�����|Ҝ#��]][Ve��N��0���o���\A���������嗟���~��˘T����f�(��(F�d6ޙb<`0MZ��D������ے���$�� ֑��.����d9�}]�@�l�p�Sq�!���X���7�n��g
>��?�D�-0*���ô�N�jV)/��3��M]8W:�˪|�[�9Nq�tqI�
�'�����R'D�e���q��g���"�?\�c���t Ձgd�B&��`�zw��:2�ݲ눘�2^��'���4|�����Ji	w��S��a���̶���q�r i8��ˀ� <6(�Yh��q0�\|$b}롻`�������4�������P"E���e�Z���}�!���E��*�:OgxQ���̏�V��8�0��j��\� ��N��� GP_���H��v��HY�y8P{������:��~$���K	e�]\z%'«��w㑞1�ɀ���#RƠ	d�`����ԛc�>�7����4����*�mvz@�[�U(;���\�`�&RD\\�zvi.�^�OST3c��	.T�!Ƀ�2�����&���^�G:����`�:�c;h7}�n�e��&�L 0E��+xy���W����g
��
e	"���onohrJ���(y��1q".t������!՞��Qq'/����e{��!z�I ��Z#&��<�*���/�u�� �+>P`\\M���#�;�I-���p������]��.�Ĝ���������~�nV.VŚ&�q5�����_Q�e�ˋ��S�h�N���Ǝ�%��6�HP/]�SlG1x ��$�����n��/��[jc��@u���]�ɤ�k/�{1�=���[����	����Xvz'B����BM�M|���#���_�R}�\���#�����BA�@Q���m{����,C�h�dw�y5dd4!�}��z����Ĝ�:%X�hIfC��;��z��sB��7#�]�&cw�J+�6�.�8�rpK�n��E`�=	(�Ʒ�����E5g�#�����P���������w
:��Ͽ�n��*V�ہ�zZ�^Q��I��8o�UT������K��(�(gx`���J6�'L+[ ��0��$#�� ���Ɓ�qA��y�\,�k�;���$���O���yܡ�B�r��TϤXZ.� ����	&�Ц�D�� pC�j��e�C`��x���#�����^�"p�S/S[S��>��ML��@�1�����:d�'�����g���A�~F%�/�ҲuܶrD��hK�&�Rl�5��z�<�=ٳ�O�L_3�$�I$��>|C��PI����D$>ĿH&#�,�U�έ^����Sl�
q�n̤��o?��B=�:J�Þ����cn�,�&�AS,4�v�U��'^$��j&����	9GV\�:�C�`�������3�@FE2� �e�U��΂�%�K@�&�@�xds@p�ee2ް��݆d.������ҹѸ���q�	}8_Qp��qP`�;�hU�Ẻ����d��+3�/|v�.���Z�oL8�Y:�]�|�ӗ��6�n����ƽWކ�(�&���S��	�Q�<��l�D���vύe\[�����?�})�NC>�I2����Y�͏\��MB~]�����$$~
��1;�˓�	!Ohy�#�7�,5o�����-��)d�c������h���,���<�r��_ԟh	;*
��@"����+_N=�� �,���=#��g��X����}�}/"�Q9�6ُ3��RU։o|�w�^������?|O��?� ��>��S����L�Q%u��~��w�����W��5/�T(s7�ˢH�=!q�v�\͠�t����2���n����	��s^_����뿒�$���A��OR�I~J�Mz@5�R5��t���U:���lX�	Dp%���}�+2H��ENEM*ɋ%)�QQ(�L�;�6�q��Ǐ�F�Rn���|�~��<���W��]�U�򾠹�H�<���Ld�`�V�-�	Q!��sY%�,n&�˲V��>�ѷ;����ƺZ���� ۫ǧG"���F��~�� ��#.2�M�Ѥ�R���<�aBY "I|�&�0@ ~F�x�|�/�"��jp+ɰ.b���.?0v3e%�JZ|$�V�M�=�!.$d������;���o�,��o�'�c�g�H���Bt���%���!�]�_E�mVX�ŠwW�qo6�3F⼉��8��Sx���#�iz���i�!�z���e��?�ج�㒩յƓ����;�>3���g���<ۅ(�����������v�UX��]�,���-�T�H�\^\���� ���}|~�����┃_�?��$3._�%W���l��3���O1�E���0����ןe{���8۔$�s���.A�?�S��L�]]_�h;����#|��3|��;R���C䏃If"��DKViЦ���.?��V��,��UUaCNt����i9����Q0�r�v(���&����V���k��-UǕ%�|'�
���?*�M�m�$Y=ټmG��E�ض�:���Ox+���`W�O�<���X�K	he��f�sL����ciKK���䍸��$��.��~��Ԅ�"� R�I!�}��*%��5 �&pd����r���}�^&����:�Z��f��#��q�6w<�;�K���]r���e[�:�1�r��#���,�j�Ų��RVU:fUHf�[��R=������L��Wj_��zݶMΝ'�&����*��
퉻�&��.x0�!���%��	n~��ܢ�\[�M��
6�����c��Zw+��:�ږm�[�bj�Gp�=�������&�����v�	������s���L���V>�ۡ[��b�6(­"s�#����d�5����ΛXF�^G��:�u�<����+.��%���t�	k���?p��c�aդ�B7F�^v�Įm;iUǃ V㑟���[�����!K\�B"-pУSQ�
�x�>��$���\8��������O��O?���˗?�73�=������`$�K&ny�vn3�-D��pm ��9+K��w	���簎�����h���@}-^a�t,vsM�1�K�����>����w�#�x����tV�m�n��dӵW1F~���zhY��pC�C+da��{����e��@X�~Bk��sr��%�ͷ3^�5U?�Re(J���1<��d?SiK�pX�x�el�
!�QB��_���x�1�į���"*�q�:<�6�v\��>L7n�k�mPy��BtW��ѯ�~l�H=�Ha�[��A�|�����p�����qB���!���@56���7���ٷ���k�H������}�"��U��m<�ڧ{ݕ�Ȃ�	�kfhn+���VV��R�FR�BF�UMS�AV�����P��^:�=�v�'jgZ�A3ю���͇o������n&t
�ᬼF���AF~�p
�?�,\�Hk?���ی(:}OMܺ;2���a�v��ۯ����$]�}���G��)�'�p_q��Di
�m(��(��նݲ�k��_�Y���匽ALJ��pІ��gUT���A�u����Ts��˻a���NaF���В'��,N�cܹE�mX���^�+�7��B�y�f�U�h��G������������s�@���������^W�L��A�?��N|%28�j�7�0�����|��"��j��������(���Ѷw�m�����
�xQ!�����0#?��c�E� �����Ip��֦����{6̡�h��*�@WNP��:Zk7���k�j���M��Ҧ'�7d8�@�kV�#�
V�F.(�Trn{dy9�'L��讆H��ml�6�]�e���:���q��b�{��е#���/��E�&��3�%��:d+��R=�	6$�
a��c_,F.�Lm�����?DB�C�}L[x��O��͡�����Z�{�ʆ�:̋a=�n��lC���_�OMXYҤ�`�<��)�>N�󰺫�-�ë�Z{��U��z
^
LZ��]�(]�������>Rn��`ϲY>�G:�t����gvn��?K��
�c8i��C��FFFdb9c(E�u*��
�G��.�	�Ac�C�o8<q�y��4����c7���U�9���)��-�<ϱr���M�q�Z��*N�_6���KQ�]��A$M�~q��_����_ݒu������3��:	"nKV�I\lS���]Qsqiᗦ~����W!*���P��!b�����A�!��h�UT>�`U��݋Ik�x�$���6����{�I� A�Pv���?Y	��#�"�HBIbA�ͨ�����e�O"��C�B&X�&�R�u���`�=L��@�"(��ϱR�s��m�����C�s[[T�	m�,#O�:�aI۱\��Y�fiurS���l����t�3�&�I]�8np+�/��ޫMQB�]��I�K4�q*ĝ�P�}��_ӫ�jG�,�n.�:�η��j�����cLT��xu"�KvK���2釓|�"	E�|�-�wH��zy��Ox4�ˠq���zx����G�͐��`�X�x�086� ��/�'��%�\��p�f̄L,gL�a /t����r�PM�c�je+d�&"N�\n�u&�Io?�_M��gbXf��1�p(����_e�â��R
&zy�eP���Y��Z���?���Yq\
΃��K/����KБlF3�N%ۿx-T:��T$��}�V,��P�B\v�����[r�A�2)���
���ry��� Z�ou�K�y���[8��}%_��9&��������LW�wdkǔY�ۡ���&>Q��R�!����} �kW���yV����BR[㞧~m}���^Qx���Ce�ƪ�{����� �d��Of�ء�9�D킴���TV2ȭ��"?�h��ߧB�g�2�,+��'���k�[U�DW9Z�\��p�R�*1��6�֮���s��x�]=�s���$�7�]WPNXz���E��KpE����@�f�2iƖ�1���"�'<��z��D�hgͫ���ߓ[��K�����@��l�1o�X��V�-�rm�PF"����L�v�N�ᾦ�l����/N�-�iH@�2�} eW��eB��<�Dʄ���
#tp��9P��h�|1#��Q��Oj�����_.9��(���&�W8H�㙀&���^g��;,�D[�%����<^zbǫy%䥬F'~��RTʅSA�\��D��>5~h�"��evk���>�ܛ����߭�.��#ZQ�:G���0�l}���:�C;#>�MgrY��\���Z+;ͅI����;�j#�F i�H>2ٓ�a-�Z�΋�I���Uy�l?�:������:V�'��M��ʉ�܁�֝����H�W�H�gz^P�Io���`=Y'dy���'ħ�7�����+N����S|��c[o����d��i`��l�[����_989�w���$��\r�1�X��	��U<���ЬW�"�����S�}�^;u�O�C<3x�D;+g�K��"��B��t˴�坈q�~�_ZX����%����-��� �:��q"�Xt���-U @�ݧ���]���W`Ŝ��K+/gŴ��V���/�q-�I��E7_y��򝪣�W�u�M=Xi�܇�k���3�N�p;PC�e�j���܆����G��m5!� �}���&JM.�ֶ��F� W.u�kZ�ig�����ouB��C���m)��^8�y�w6�R�i�&�F�Ñ�[�Z_��P�S[+��~m�D��/gR�
��1-����b�?A)RM����vmi}L�}?V��q\�O�y�q�f��Ʈ�-���k
��H���ՆD8���}[FFdb9cG�@:��p�2pT��T>�>+�7NA�|����pu2ah�/��8%�q��
b�Lq�����f�y�"��>�:LI��xݽ�eX�A~`h��`+�Y_ �͇(�FХ��B�9$���U
�<Q4�Q�]*��:�$����X��yO��\�o� ϓ���|���(o���r����D]� ��!��;���`t���c�ᐆƔ�(oO�bL^��j�]���6��|8%7c�gK������x�>;O�Ó�#�;�v'��x��u�ŬN8�3#L	���aإ�Ɖph�����!�#QQ��Ov�b$��:ȭ�a����`�+�g���>��m�@��y&�3�����H�F�si����wi��|�JeQ;:X�Nހ;M�"��P6��B��
A	n��d�R�_"\�/!��'ƿ��k�u0�.��a,�%�^���1� ��K���|���6�n�h��i�HkO��OC��.2�*�~�c��ݚ$/C�$�K:U���v���k��D:M�Ƀ�%as�Q�,�MeW~�
�[����N�5��K��!����]v����ۡ&�־�6��n��:�h��'Z����4�o~��4{]����z2+u�6����c���ۛ���:���;�\JQDǗʷ�L,g���Q
�����V�+��re���$���}�9c!�'x�^��1S��{Yc����.Cm��}�����ӥzfZ{o�� ��Ɠ�i�&v#��X��c��w�'�I+�|�v.���`�'����e��w=�K�T�RWR�odU.ۼ��=�k!�*�md ��O�����B܎�v�r5SvW�=u5ɧ�ퟁS�R鄔�'��l<5]�,��m�TY��|���N��ES]�z���N�������"���B~)��ie���[����Γ8B��p����./.a�aWf����gUz�y���̑�����%���ڒ����>���އ�>'|�Fc���bhՌ��Jc׌���\�N�����ҹa6�\)_�|��SۂB1��	7
�m ���ҹ�h{`�y]�̳�A����D?�ʍ�h�~��㛂U:��0�:����fWW����*W�km��t��0��L��8�er������6���F_$';ݮ��l��� Rٟs���,mݙ\>di�8���*�M�<�y��Kc����l~]q ?t�q}���q�
���L,g��hu�J) �zM��Q�|�RYLѨ}�\��z�7�Z��l�Y�|��r_�3}ày`Ê���o��넱M�:��%��M���9�F�0�S�Z�G�	>��\��W����~�����5k��R(y�h�F9N刍&�[Q�+oY�� ��u������T��'���S-6�mAzu�T�N�rO�b���Z�Q��Ʊ{m����g��0���C7v6�1##��C]j�#�rE*7��n3�9��\q~�D]���_ed 2��1
�&1eaaN�����@磧j�hrC/s�7~Sqa���ʖ��a�ϨD� $Fp�	�cf�
��M��K9�`V���t�N��D.0"v��)�z��1L���zݚ��eS&�u�����:E�^*�����܅(M��a"��T�ΡʑU��V�R��unEd��J���z2�H���@����¸�Oj�V=�%���+�|���`�v�V�. #cJ8k��^�.U���PÑz��{��$;�X}��|o;�(q����Ϛ[�^�����m�16���������5\^,�ˡq�ͶPF?db9c'�Ry�&�������hQ-[�՝�X�8����Ƃ��y�r|8j�G���pb���Q+�ϼ������O��q�\��6��S�cY�>�W�WYEʪc���P<r��Ώ3=�����j���_��Ծ��y�q�+����tʃ��3����,SO�Fh<��<�g?k����{mQ#{_~��;��Ԉ'��?�F����8?�6B5�h�x���"#��[����$��C�hҝ~üh;���-�pih&S+u�����啵6,r{��w�]��%{�n] �%^�������\§�W�8�GJ�3+Lf vA&�3����������3<>=n���$	���εɆb?͆4��2���ex�M;�?�	�l�@~�T��x���O��r�d�旺��_��+�LՕBeP�V"�.f�ŬrF�p&����t9�z3���:���H�)��*&R�Р�U�ˈ3ȇsC�����:�5�*��9��I�.���I�'N�[�ʩ�����I�F.� mʾ�ǌ�7�Qe>�o�czܠ�moo�ݵMӀڮ��|�I�VmO%@oB��u�U�p*-ǆ���~[���^��sബ�ݘe��������+<.�����5\,��m��Ȕ�"���; O�m6%�����^�E Rm��g�0m��]2�Ûu�aC���
�mC4�A�����bb�Z�������k`��7���[�k�Ҩ�+ޭ�t�oP4ʽJ(!m�&\sD�1RO���yB.C�9!�ϓ��a��e�"	�&�[F����*�h.{�@�=��edC7�\9�ϱ�cL���{����HlqF�'}{$��̭Ml���#��c�}��B��x�G�S��q��l�����r��?����,��p1n��e����G&�3��r���zOOO���f.�o唄��!��qnn1����Z9u�'�SD�V�ҡ6��a�&O��,Ȱ(���ZZ�"���@�\�=K���7o{nk��f{��+��yv����'�9�E��Q���ߘq?�zS۞�4|$,�P���T[ſ��b��� eSg2}5������y�2ì9]bb���32�	3���;p{��\{���>Y-��w��>�[y�]���'}��鞢ry(�f��?���������L,g��S��I����+��w"[(��?C���eJF_8r�xz�qe��J��FL�+*>3��8_�ZI���]e�������h�]D�v���ʷ�^hx�U�V]T=G�2�bC��ȽO�����s5����$oά��K���V���9R9�RW�^D�����L=V�ޚ4V�Hh�]��ܵb@'c�쥭�d����22�ĴQ���_�꽱4��	���du�ؚ��o�p�YV���V����.������\^@6�2����^�He\.�Z����6��Gm7؝�����Q.�#�GJ�jߕ��9Qiea�[Z���t�)�Y���2����x�1�Ϊ��ɥE�R"~�@�-�$a?��]�L�yC��n���-F
���LO��4�f�|��nt����<�R.kc$��O_(�Ԁ�{F+"�'Sr32� m�s߳�零!����<����X3�=C��o� 7k��g�����~������o���.v��3�2����E��_i���^_^`�Y#�D�r[cst]�.��=Lƹ��  5i��=�C����j"�)%bH��L��^�B:����MZ��X=1&D��SV�ߘ8�7�YH�����J���� �ٟ�-b�wj��V}8��t����@�)��TS�>%��XR��� 5�3G1��Ό�c.�'��zlO!��+�����,`�eÎ��]�e�s�Sm��x煘%��X�ٍ�?��V����g�G�C��%Fl��iL���L,g�k`˒|+?�<���3`+&��o���У@B����e�O�KC�O�*���p�S���D�%���n�R�v����""�]���a@ge�w
�J��ή���/�n1�zS8F����˻�dm������Ʌnز¤m�Ѿ�bd{�72���1%ډ����Ú��<��*�2�󢕅@f�@ĺU]4t)�?��YW����_�ͦ���K����mE� h�F�Q��z����6�zQ�M��[�P"�1f���g��N ������]��rF'����??��oe���JYaJ�������@���/�4!pnVɼh���W}+�6��"�����8���~5�E�S��s�9r̡EI�n24Rk�"�q�1�@�Х�-A|�#jMCue�'+����m�q2�߹2Y����O�[��\�Ș�^��:�q�b��m8������~�~��O���7���\^]�KT\�n�D>�-K(�_[�1�˻b�Dr�ێ�����O�Ǩ��%���%,/�?�{���~�nG2�
���1����N�ʏ�KX�����#���B������&�a%R��%�{���U�����d��u]�}'ǧĝp˵L���w�X��vR'�[)�ohҔ����>iC#"�.���s�iOam�@�b̭�=��H�1W/�M�9V��ە�u1Մ٪/����*?�ඣ��g��"����8.�ß���[ZQ�9#�|F� pvl��hX ,+�m����(�������^���������.��u��L�²�̚R�3�յHu���٠���XH��r�(�T��KG0o�.���b�P��///)_�g@.ù#����}G"���`�m\�W�/��q&� �7�j�32-!�X����R_�	f�v���X�Mu<a�5����᳿M�Ô�!s�G�<�*!J8�����Z���3�U�?�[��!M�e��ڠ�;ʀ�g��Brǁ@*���~��_���qǩ%�M�8���J��R��G�@~$�//ay�D������V��ݻ�!�<���n����DQ�����
��w"��Ǳ	$��A�C��pn,�s n{��Ea�B�\cl�#�|E�p��{ww�����v;���������	�5����ݿ$///D*������ʼ��p�Cv�p�P�9�c�T��C�٥���*�y�ѧz�%Ho^�z�%���^���ݾ����L���4;��Ș��0����5�h��͌=`~�����6]6��z
����9�UY@c��^͢���ùY��1�K�m�\!���D.!��׿���~��~���w���	ۈ@��~��J4��N�����}�D�k��v�����������ö��X^�_��z�$��~�x�x��jO�|yx|���\_]��� �m���˧>g�,NL/9����v�Z_q�W�)������,7��\)_���XR;Pl�������qn��o�SZwu)�R��EM��W%ֶ��~T�����^Ll��s�*�FV��&�L�C��{��Q�H����o�z�h�HU�_���6@�T��4����̀��1燩K�:�ɺ�4d�E+��K�m�
8���]�&9j�l�|I'��vH��~�mr�<0[���1.G�A��YӰڂ���5>�@�H�a�_�U��3�u�F���8�d{p>���<��[�nf���lY�J*��^���\,������)�׫	W��� �q��,;��q���B���Һ�-��C�,K�ٟq�M����n��OX�6���9J[!���b4��7�c�@Iϻ��ȉ������%����|uuM3*����ޖ�[oO�4�	b������鼸Υ���fD�#�~7@b�8a7V�?����D�pyq��w���හ4��݀9�����E��QM�e}�Q.��6���{�Ϩ/����l_��4���Xq[ҵ���nj�yM�j�VWޟC5џ����j�F��NxkoDU����A�.���?�>�}�՜d�R�K�M��O�L�Ȏ�^�`~X�M�މ��'iRۨBӚ�NsvzNED���+���2���1&L�Lg����sA
w��2���+rb4�J�~	A�M�e2�Pw���=�/�P�I�?��ӹ�he�m�(��˅#�KؔkجK�=��7wpq�����'x��'�[���"ry���ެI݋k�0D���--,��|��pHFm\c,����(�B9�Dbi���E�@)s��$���]�A��:^��WaU���~��=�%�2��}��7w�������q���,�e!<N��h��0��pY�_Mǟ����;��E�\���E�Y.��u�?���tN~�;��A|��,بc�SӶ���1����C��1�ǳ�A�hzG�gD:vEgju�;���s�a�k��n��x����4�E"l��6��Q34��6�5�Ӥ'V� @.§k�*�~/nl�9�n7c�}w�8�$�,��D\��BSK�q�����x�}*�3��_yI���\^^i���D�ׯ_a�Y��a��쀂DR�����m���ɠ����"Z�����~�KR1��Y\]8X)���/�[��n5����0����VFx2w?���aKX�^�����5�+������$�%B�Ǟ�rWV�Ys�Y����~"ņf��jV�/�F�O��������"b��Q�����8J�T�e!]��������J�oT�Yc�'6�\}ן�J"�O>m�d&��ȚA픜3��9f���IJ��D�1B'o�<W�@��3�&�W��{��C��儊��l�����T+�a�:2�����;�S��]������8��U�i��sL*�ֵ������S*JC`{2�K��!��p��<{hJ9���[� &v���n">|� ��+x|z��}�c///�w+�ͨ`��,h�^�19+��a@�n14&�&�K"��ru�e������)��E+YEA�8�$��:Y�LBՊk�(�=��ܐ���j����r�B�v�n?�9ؙ�I,#l<�0w��Ɂi���T!�M=#1.�r�3��/x��~��;|��٨�v��ͯ//pyuA>w�7���������i�fz�ۊ�N&!)Ie΍��i�#c ۢ�����Ν�+�'օE��Z&��XN��0��s�O5��OD��S���r8�~9�����ړ��t�Wn��'T�:�C�&&�3��QJ��N��so�/�ށpCei��aT�(�������+�������\_������W��=��yA�Q|��� y��$�&x�X�
�.m
ﻙ��t^2ӆ�f`�υ_ק}c�g>;��_+��.5��9̇��gxy~�ۛ+�J7!�8!�-��S9�D�����7��쓿Uߣ��0�opj.�>�����g�+��a�̱����=p����~��gjL��ݑ�|.�Z'�+0C������W4��U���&�ġg++���R#�g$���N�K=A�Y��g���S"�7�L�_�
	{E�U҇58㘭���F�w޵)2�YV��̇ʻ9�ܴ�Q���~m7>�q�9���bl0��$G�h\	�ϻ\~D��C�J�<��^����=��{��W=���G6�I�=Ң�~'p|�So�w�Dan�O>��3�~���� ��WR�r��꒹,t_a7�]�u�2��x\ʭ��a������@�D6rmʕ����\�⨦ OUrd���8Pɾz�Y�-�AT��QU��j�K2*���M�%��60��+q�G��0�\%��m���\�8j$ͬ�e4������1�g9$w$�+�����#Z�sfN!0����c�������tͷ'��L�m:���ş�A>cn�����+��r�[�:'��&>M�� ẳ/��L�����(WaW��z������m}�J��&��z��5%S��`�4,\����=زG��a/'�a�-&������3���K���l�kSu�5#k�V�5�2aH����]�?w������!�v���>����Ϋ�)cg�����ֺ������K��D�sL`Eu^��@�L��gu�b��k�m�:��~d�Ć�9�+x�:~^.����o����'��z��n��c�}Z; ���#����*^�%��#�UF��=!]p
����Jv!�h�j+��F��|�P��Ɂ����j"�W&�����8KbQ���"�5Y�3(����/����8��7�w��������
����q߭U�&ڧ�IH<#Q�Q.�,.� �ϗ��^^,i�h�`8����r��I��
C!�d��yn���/�����o������ׯ�����+F����,�b_5��T�lm���C>��{�&u&�T�{ �{���i�?������kC�"���z�i��M�L0��m����|����G�hA���A*��j�}�>�b�`Үٖ}-�����&]�S4�&^[x�4��	̀�u�c��i�{��>��Y�H�!�&ɷ7׻=�R�Ӈv��ըo�yP�R����db&&�x��m/��$�d�w�5a�����(����qT�^.ז�4�}���ȍ���Z��S�ȃY��l,��>��jƸ��f�_��,�t�֑̅��ٝ�|�mr�e睘?v�-��b����r�?�IYQ!k5�H�B.�!����zbY�Wm���e������\E�*�3FH��EP/�|ED3n[�}�МH����-G��Xn+�)�/���������� 7�����SX��Y���A�o�^~�=�Gj�|d|W�(W̵m�'��0]۪Ā�S���v��HV��}�wu�&̺�h�c����cw'�L�7�]0������2��M�n��������&z3{�)cVh��I����F�n�?�buV�N����e�}b
�r���ӵa��L/�Xɒ�$�m\e��9�@�3�;��.K�����UO�����}vk���]ⶣv�r&R>G�)���*±��a`�]�?�l���Mx��Bae��I|�w�`q�`�����~��/h||z"��ˋ�����~!���J}?t���6�s��FV�WӇu�_ iL�U�\F�E�7+�3�Q�d��l=�T˕[�D�K�Գ�Y�l�e,H#���-�H���J��`$]Z-&.'xF��mG�"1�ql.���OP,K@<M�̄4��XQA���0ޭ-# �|]|>Rc�m~�Ħ%7�7Do�������ͷ����������/����?��Ǐ��w���T)9���q:��b� z�rkw���z��+9���Fjֵ�(� ����F���N���H��}��Ie!�=��G#���-�[q߼���A�X��)�ob�f�I[�2�E�9��ܖ8�7q�P����3M�������zl(Qc[����;��C&
lrS��e��QY6���f��
c�����rH��E�vo;.Ϗ	3���
C����� 	f���.�w=�6c��ϴ�i(�GP'���1H�= nj��1�*Ì���m-���D��?�L<��㧟��_����Hh$�9`P��1����е�Ϝy��0y��|92Z8i|��Rb�m9[X_y�r�%�6@8f��I��75���n;�;�ΊX&Y�S֢B����?X�_^^a�^�j�����u��Λ��D>���;���֪��0V�蠐.����b����C~���j,^1V�J����c�s���ww���O��ӧ����o���t��'�j�V�Iu������`9uC3#c
$	i3]}�tD���_��o�<�u��/�uv�a�fH��(�"����]$�t��_�R!�u����~�'$�I��)����i�5���=w}Nm��6��/�P}Ӌ\����`��]��I�������I��<��3�7y���w�1I4�v�j�J�T��W�ט���������@0f&��?���T�
G���X_o���l�DX?��;;�e��>��k,0�U���1=�Ef�����5�����KY�P����W���_H���O5����r�,(h��g;R�td��\P�����J�L�5�q�nU2��0��2��Es��.���ͼ��w6Ĳ&h�deb����חW��t�r�Us�.��7vja��l�,��Pc��o��V����)�����"�7�����-UP������;������Re��pG�޿������\]��������܎T�)a�\���1�u�M�Z�Z���U�+fSCs������Y1N+i�����2`mR#�����H��tpS�L�_�ך�^a� �<������A��Ƹ?��sDY��6��7oS�ȹ�	��k{+��Ve�`m�P-L_�r��[�Im��82�ۊ��wȭ��he�܄`S{�ڗ�L�Ї�A$G��x �K���2T&���;;w/�f��0��4����hB�D���?���k;�b�i���v��O_Є,�R����M�@����$mP��(5�2f �.\�/㶕�~��7�|��o������u��C!2�5֗m!xi\�|��Bl���%Ƒ�V�a��Õ�M ��<e���܏��fMl%�g{;8b!&;Θ���H�Jb�(^�j*Ɠ��oZ髒�U�g�G�c��W�0�d�U�zFZ*�岮��ځ;��@��/�/��/��������o���9�6�����`�]]]���/a,qgLS2?8J��M��0s؃����[�X$|	�K�ʼ�����j{�ܮZ����+���n�c�2��ᾪ�`�
<������6-��O��4��dFy8v!�kh�W�
�U���vk_�l���겉�׼��Ի3sEX��He�@�ˏ��و�eR٥�5��N.;�<�&�\��^[W�]#����r������>y>LY?fd��/� l���˕��,���T���W�ʚ-߼f��偭�HI�5۫�P[��}�d���h�ۀ&b�X:�OG�G�ed4#L�:;ɲ;�\c ���`�O�~�o>|��~�	~��7���~��䢾�J��_E�����u�ė|��dscP�"��6���>��q�7[�Wޯ��^ıl	A�L����7�� �5A���DJ���{�O�xX�؍w��PK��b������\��B����N�`�{9�\�/�j��GG G�B��l�̖l	�Ϗ��8��^i��^o��陖(���G����?����2جְެ���,�K��6
�Pf`��O~qe�h�˂*$ܬ�pJH��3�A�����F���'*M�q�B�b�{[��� �5U2h>��Ҕ3����}���*,m�n%m��~ŉ󙏁g7%��Œ}�c{�.����
�_�9�j�~I`��������[{���̰��e?��=�]� ��Q��4��C��I���b��U��jO�MD�>x���C-O�'�D	Ur������h�zS�ҷT����τ�@Xh�UJ�mVR�����Ӛx*�;^� by��d�͕��ghR��0,(`�V7����VX�ׄ7dRu��&��!�<&���>&48b>@�����Gw�dqO֧�wYۯ~�Zy�eQr�$����t��.�_�s�ki|'�~��_b״k�,�c�o����������=<>>�w<y!��
���]g;�Y�d.EØ%�9*��
G�+
<֩�IIDt�-��땐 �9�ȯ�~r/T��L��M2;�;�?�x�����}"��`9bY �잟ɍ*����!�)6:/�T�7K��_��w�b!�Kp/��������B2�m�6�#
�p?��|w�%��))���%m+��o����on��>�w�?ûw�x�i�"?8X�TaO���v|~�0�I�rлBw"nLP��N���<Q���隫��>f|^i�1�jP;���;ꑾ��Цj��p��W�`�-`o�s��[*ԟ�|h����jK���@��/A)����>��"���Mb���������&E����d4�j���I�g�Sɢ1�n���y�t�L8;+.��^IV�(����+�!ߜ���6����Fm���T�Uik �z�_�{JĚ�I]�(�Q�4)�$M
�ڽ�C}��)?��bk?6Aڵ޿��'$���]��`��/���IV��I��ߍ&ԅC�c�L�%�;�Ǝ}�t�b�ρ�&njE�5n0�W�sUzfw_��*Q�)��仞��/�V-83���&$;'*��d(��6e������Q�MW�U�l��d� ����C�A$f���p�4�u�\��s�6��h׆�5�no�������?.��P̸Z�����֋)me�X�;�OI'���)$��@<f5�r�wז'��Ow�e�7����V�-n���Bw�iח5�=燳!�%�݆T^���Iy7RP��zW��]�\�}��R��B�V��$q �c�6�y��p�����7�.7�82��&c�}�����[�VP,������/��������m��h��%D4V~"�'�U��&ЋŒf����D3����/���4f̏F��Ր5=���F�(��m:T��3P=�1�J#�5�M���M�J���1'���F�;Ze�*>1�W�E�i'J�n��kl�%��H0Xi�7��Nb�TP~ސC�����~�&�Oڸ��"���B����P��� ˤʞ"���b���}%��0���
�zH,�	�D�_���	�B`y�����K:��ç�V4\:;�?������fB��(�����H2:5���ܰ�0�]M�0�/���G�����@�m:"G�(2f`3�����(���4Ix��d?�v��u��{�b_�%�] �Ha�l)&7�ꉫ$���M&)���]�[.�^�B�l�r؜LI����<"(���]�x{��W�0[�g��r�#��O����P?M�^U-��u��"Z�<uo��O����$������ˋ�W0�*�����_~�/_~��
���;�`B��?(�D�3�X���<���-����\�i��U�5��ǅ5��v$4W��+yf��rj$��gŜ	1�?~��;���2��oD�D亵�~�S ����R٬|a�cR���ޯС�G0��a�x�b����LV=�YJ�qKGX �b�l.�����֔?X���zQX��ꂺj��/���ޫ(V�D+?T����Ўv���5@��k�_虷���#RGG�DNW�Mܧ�P?#qdO����>Q{����������Ք[�OzpD�Վ��MĲ_.�;��-��Y��k�������2��*d\B�\B�P�H� ��㎧6t�`d&2����w�'9��h	�4͕ �
��?��c�[Ü>;�Yˋ���+7�� R�z�L����8�R��!Y��d� ����c:q��QV������4?��e>r�;7F�W?}$L�SÑ��(����T�U7v�W����U�(��wN�#�B�>��L]������KE0�?�e�8F����&��j!�x��;��4�Dp�Ӂ~ņĲL���H��f������=5��F��~�	_��=�pbyf�Ǔ7���+�������� �}`C�r�E�j���NX���ooo������ �]c�^W���"�	-l̆)
��Zp��U��P��s�W��2�?�lI�\�@��w<ݭ@��.���C�67v��f���gC,Kø%/n�AOE�����$��,q�8W�%�S)����TJe�V�%��T�6>�fQ�]Y����~k�,�"�S��\�L��l��oN��r����~�l�bc�´#1�����D���koj¨t.:0��Z�0pX8��I�ilT�ۛNޠ��i#���M=$cr&6p��H5�"V�U��-�#$�=U���T�z��.T�ۃ�(�"�54�d�͚T��BӠ�O�IK��k�T�e?�Խ�_t;)i漤�aa���-W�/�ӬQ7�u}��{�c�K�Ե�&u��q�{.�.�:������(�OWV�߬�o����m�R���>��R��u��w2�}����N{���ky�H�/6"a�CaP�L��]3�=��omo��/��s���`׃���%K}��������k$-�J}8�J�ܒIl��%_��r�h䏬l�KS �Ԥ|m<54�t�����z�'/�E�*���~��1��'NH糅��u������q�W���Il	�*@m�����"�M@�57�*�z�f�KjsX�����T-�+V�~���|�c����Hc��\�n}P}�\Rp\��HF�ϣ�Ng��2sq�un0�fH�b��Yt��&1�߂��m���Qo~ΟTF��,K��~��\K7�a[Ykge��+�K�?Y��8��U�9,u�:�F�}�0	HcA-��L��>�䐼��󞞞��`%���>�>�����3�	e؇d�@U����W���)��;\�Æ����7E��[�˴F�9���,|�G\�:���qY�]=���1�b5�M�0L���똬E2}�Wb�/�m��;bS�t��w)�*�t[���DB��B9�E,�d���F)c1jT{�`�ߘ3��/xzu�����8�����^���A�lK?L�Ng��g�U���r����$�y���Ch����N=}�15�S9��H���j$)z���˄|k�Fm�����e�n�����r��$�y��>ۧy^��mخ���w:���ީ{�ӒU!?���:�f�(宕6����C�}~M�y��t(˯1�8ʘĻ�X	�i#j����}�@�O�]��i?��Np("Y���c4������P'��܇�Gx$�{s�������
NY���~w<�ph�a�=k���ł��!�m+���p�zuu��)�1�ׯ��_~����ʢh�/3�
�%�����"��m���g���.H%mQH	1χ��D�`dt����#t�0D��`��?V�����/U�.�`�OԊ0�ǯ좂}Yzb٫�˄[�J�>�i?�-��;��X��\pw*�@�˵ei ~�@���n�{�>~�>����z�2>ӒH�*�:]�"6*K�
nY�jk��{^���zd�	��g��Q��Q𦐐o�M��G��y�a���;ڢ�n�]Q�b�;EjX�Gڙ��x8=�M@��Qk�Q�80:��D,��#P�������R�$mI%3�V��F��K�h�� ��m�I��9���n��I� 5�D������j�.�����	�4�_!z$Γ׵��ts��4v"�|��W�כ��l|&M ��Ilu�c���_��[W�%^r���0���c�f���D�@��� ׎�@Eʓ�	�3V�q���u+`��J�mԒ����İ�(�2m�o������tĲ"��u=�Lġ�?H��?a���/�l��-A�/,LY���yn";�'��x��˴�x/�>L=I�q�[�z39}vT0�`�.�P0�Jf9^_]Ӫzv�������-6�uI�]׀��y0��-����=�"���8x�����Qy�����&���pj���l�e�,��IǬ���?.EY�	/�}R.oD�\z��\VKM*׭�m�3� ���\6lk�o�Z9�5<�"i�j�ק5������_��>�77�4�^���R����q5���Je�u�k֖�����b�l!�#\�0����5�G�L����h�	ms��_�������R�w�~l(@���5��)��feIB�<k#�,�&Ԣ�Gj�L62���nS�`�� a�9<�A���:��	���/{zX3c��+�K������2�!oKRW��z��_O+�j7K�w��i�o��X���6�懼�V>�ڬ��"�zjqb���|���0�i�Q����_��Da�q�	ڐ�������Z�۱YX5W0ݍC8N)�����v9b�Apy[@:!&�P�V���{����7��X�ϓ׵r���a��e�9���i��g5��±��8�G ��'l�+�wJ@P03�6��)m�����H�&�n�����K��j�����+��x	�|� ����?�����_��酄�k�{Qp��+2 ��Ƒ��ʨ �����'��6���c���D�t����D[�,N���/ΆX.��]J�E��*��{A	]% �;R3���d��	jj��9�rYz��������~���+ج7��\f�~(Y��vA�W��p��~��{���f�^�_`y�3BW�Of��	S�n�$���
$F�B��c��ƾ��v�\C:�,Q���=7�!h���HGj���a��춨9��n!��%-�L\�~E��H��Od2�,_�טq� Ř�U�S��;!�dT��EXn�ơ�zcNb�畃o��T%�=i��Ӑ�:O�
�䘏Ə�T�ú��ہԵ�uDV'u�q�&�����[$�v��43�}�yO?:O훧/���p�h�tH̼����7�vN��x�!��\��)Y��0S}��F��b;>Z,���q��k(]�n�pZ�߶�ҍ��FO1�i}��1��G[?R�)]��Nv-��4�Z�Eq�}32B�Q�ƈMj�����Ve����-0���������?���������xzx��xEת�5�Ԩ\&w�q�˹}/
��q�+��`�N�m�B���¥�������?:�6eB��\�Ӵ|2��K�d�x��BxrY��S'��Ґ��g��My���'�_&�(6��X^�O�w�������w�mK�#oT��)zz��4�&�Ⱦ�4Ѭ�Ϲ^�8-&���G{c(���,���Y�܇�视��}��~Ou��۔6��)�iC����f�cx�-&6�(������C<�7<������`�.�O���f���r�z�Q�r�tm�T�+ZOb�j�Qu5�3��^Q��HE�&M��׮��I��x�\*��tU!��ݻ���}�>7�n�N4����ԍ~hV�����
���A}�A��f��e������}Y�}�"~��В��i�[Bnǫm�L�5��JI�'��>��R�Y��v��u��ݪ����.�0��j�w���+H�Y�D$�N&�8X%
��[�W�Z3c�Ќ�6�X[B�@���Qv�d-��r[7fE�-���///�`������������?���<<<���<��
c�/sA�9�p��d�qr��1'W�J_`y%���o�#$�Ae�_�7�q3���4]g��N߯�ٚ���,���ղ�#�X��\x���q��˒ˈd�E�"��eE)��Jg�hr��jt�H�`��vk�`���ͷ����Ç��T1qf�c��VPT,#d[�7�1Y;@���t�9x_���D$���SH����1�jw�嶑XV����dZb���Y�9+K�*&�&���ж7}�Sx@���������r��O��?|컄2��:h���|3��r.�z.���>�B{�[�� ��5D����!ӓ���cZ]\/_}���ÎlOk���:y&����U%�&��c���W/�n�H���]��Q+t2j��n�n���'2Ah���Q�W�8x�>����6�_�e��Yx�2�uQ������U�ŒT��:@&Y2����I�;*���1�Ml�7W$�-+�K��W����!��x!���ׯ��_�����xBdͫ�T��,��:�؎�p%J���(��  �<�
����-f�MgA�2߸ 
3Ќ����q��]	�;l�^=cb��,���#އP.�w�l$��8
$�&�|q�eQ;�I�v�����6�c���3rJV6��X!�#���X�������kbE��%\��4.�\�Ἰ����L�<��&gd¿��U�W��&�WM���9"C4�)�Ý���P��i#��Bx�Ѓ��j�Jtg[�'��F?=Ɛ�ǠcPe�$u(&����+Ȃ�;�,v��B�5�^�7K���p���N;�]aX�W��#,K�r�4�LDw����Y>�s��Ҵ��
@���m�4��E�O��V��!�C[����W�rff���'��!#�-A�f=&��-�>k���Wn�g��F���`}�&����~w��7�hܵ�c�VG��ݝ��E=�d�Q�Y��HE�(	�B�S�������@�	���ez��'2z��&Ye��W�ʂ&80�*��@s]__������xzz��<o���L��d^��t3�IF*|�����2PѼ7�(SVH���ҍ���lC��7<�B�ϰ��M�[göU��'�^������U�6��f�dF��+��'n*�q▢t~[�X��J9&����w����)�=qmɽ����_cCB�t}q��ݶ���w�}G3;L.XO����r �BN�xm��t��#�����r�$E�xŊ��>S�4)�|3�bo	�Ɏ!���.4���n;�<�Y��f�D4�G����U;z�SQ0+ڃ�Pɡ����n9�������*����$(���֧^��Ԛ�|��o����6=oK�ׯЪ�-��o�tVr�K��N_v�c�s�P���R�ZHo����aB����i�Hol �®Y03�_R_農O��1��#ΨD<��W4���Foi��֠�m�=�k�	����v�m�E+A����u�ݻw�J��ח�n��1��b3���r���*�k���9����}�L���_�m��O�i]��\.��D%�5�nn���^^_�X^�^�e[n_^�d��c�.���iV�5�x\�)6"ՍP`?��gV��PZŅ����▰��9D��5�W7΂XF��Z:����!�)HlQP!��N���R.��Ӹt3{a�TěR�JV���_ �K���Hk>�ؽ�۾��X��T�V�3��ѵŷ�}��/���':WT�WW��E��Օl6n�w��F´� ���0���b� ��=.ʨ�1�w#��3jzl�z����c���)���iM]<�-�����k�e�~w�>�i>?Ajt���C]g.��4�=	��R�o�ԦS�o��������J�mȜ��[Hn��y�ņ\]+Pe21V������Z��I�*I�<�Q[�&�����^/�E�{;eW^Y� � �RVپ[M�g�T�ݤk��O�e��=�=wj�}���:gH�m���C�EX��&z��'��犩 j��"��� �Vv��UD#~ߚ(#����_��a��+x���Xc�-�7vldZ7�J�^m.t�͇�͌�	����9$��[�j��W[./���NFN���fMj|!��C���xT;K:Е,ƫ)��2�,�_#�'U.����E�p1m�3���V���g�4p��rq����e�Af�x��X�c���,J���#@��wj@��'|�_�&��ۋX�������j�W�M��ѹe�Еk��E`2�K�е���>��8|�ϟ?���w���=|��7ps{K���W�E֯���8��F'���8�%b%��X.ɉ<��/�Y.Hԫ���~�*��a>�`%�>��B=��پ�4�;v���[|��[������3���j�,���U=��?lO�i?�ݘ���G4:ǍF5Y/A�b"��Oj�r��ǉ6�3��N0s֜�]놙�v����[�¾9ԑ"�
H��4UFcK�ilS���+ӣ:�����I4��,��c�gj6�iꜛ�b>)qB�2�9r��~O�����i�#Gu�a][:P�����;X.D��6r���/��Z����r�6o6&w�'���r#L�m��]*�(�%3�h��5����B�2�3Cq&*�`���>w�B�ǅ���&e���4��v+G����qKJrv��'Nδ�3�Np�u�l��uxS�c	��Ez����$�����"8b�IS���)N+���8�CV��EEl�ȶ�#Y�ǎT��uJ箂o ��U��fC��\�D�%��Ն$�8{��.��������}wK/�p�($��R��θ�2�7�0iR5��;t�����A&$�� � ~�֟S�LU��53-����5]'���C0�����(���f���l}a�������}�#��gY�������N�С���А>}���/�Rq����;|~�9�1��{{�9������q^�K2g��C�^�;ߓ���xDd���v@Ӧ	�9���U�j{�A�|r]��CB�k"��}'I��P��v��+@��8��+Cd��`���ʡ��3��1�u`��
��Ĳ#�nП�
�ZH�"$O��v���2va+��4�_��W�b�QZX���@��k[RC�A1�X.0$>ڨs��%���M�7� O�{y�}�+�A���gK,W����Z����Jdw�M��b��&����P�͎l�w�2.���rx���T�>�e�_W U�J���I��X.�ݻ����G������;�g].�.}�L&�7��f��H�����4P������ˀ኏?�߽,� �'!:nH�Z$o�}%�T0Q�X��׬%jYA�Ӏ��T�7)����y�sM���Ub�J�3m��pH�O�-�Z��ʹdkn/��7�6o(�#���`ԇ��������KP�oe�!�	�>rH*qP4�9d,����·��'�my�u�b�l't�%#R՚�s�t��&�E=oW��qƂ@�'F�+=O�'���uS���g�8�����Į&�:�D�Xsx�PX����W�U/������f�sKL77�p{���b��`�I�� ��Ճ�����d�`+vu��Sv�o�'�l�딢pVn4D��\j�z�f��p?pi`������r����[�w�����n�A/`��ܿ�T�P�«s�2@����Tg<�ϰ����"�c�G�f�������ۿ�  ###�az��m���j��E���S�Q�f0D�Z�wN�2D3Շh�n�D[�H�5@ɽ�����F���0��R�Gz��%�Ɖ�2`�z��I6=���s�9<�$M�:���sj��-#�O:ON�q��6�t}�������c`~vy�b�%�����,m!-헉�Y2�
{ǀ�<��O�m`BӺ���NdjKeQqm��ADA�e��������'����$������VO��g������k^��Ѭs�����'�A//P��L>�Yˑ�`���9,)\��J�XwKf9D�L�%עZ��Ш��osT�AT�۟uP>K�ImM_��x��SKc�Ktu�/��W���G������U��%���g���euf%� M'O{��>�/K짢���p	���3ȡ����!��W{V��[j�d�.s����R�~O��������2��/���3��6F�~+EB5b���'��.�s� �E�Z���t����q�+9�ռ�ň�����0�#��^�ִb��\R 4]!(� q"�����������}BzI�B@��2JRx��5q]K�8W�UhN��y�@?�������=<�����*��G=6�3��z�/�W.����pB�j���'��O���g�*�d��Bc+��8�Z�]X�_�����Ȍ�*x�<�~ZJq�������V���[�h�n�I~�
����}&[K�sR��l���I�\V����kO�[�ƑL�����e
5B�+/%���\�OHh�������3�����	��1�4�'�e�+~Z��k���`ip��>��9.4��>�)��C DQ���.0�f9T*"w!���^&>b&H���Vb��у'�9p���f��Xd�BL�Z��.�d���@�:S��"�Nq��ȶ���5qq|z���j�2���~F����Wǉ���-:}bbŲ�XT7+��Q�,��	`�HF�K�<ʒ�K��iR\`xų���&��B.G�;N���{��)��������(�w�Ԑ__ݐ#~"��A�rA3�R�8z�(���ΐ��}-�j\��7�Z8B>����Yr��F92222N���m}j����pw�*T3N�I�Ҏ6�L �de�����[��8���<*�T���k�me�qê������i4���*��y��������)�j��9N+�=��VBTceiR�V�G����0_X�ʢ��֢�������D��v��&�h��V�ib�� W����W/�����ť�Ex����#�(���z����y����vb�\ԉe�ϓԥ#��p��L���W#�K�jv� p���ꚤ����������˫+��X�"9�ΐYB$�1����?
+�������̌j+Nl f�)�Y�J�%K�_WkX����\"xJ�G�!�����~I&�W����f�����3j�KU�W�M����JSA�C����h	����`� �����^t:���ƫ���G^C]�S�`���ړ��k�q1
UU�l鲁<�l�84*˪�ӣݑU��w��]�6�nCj?�C<�F�,�<�m��W����Έ@�Z���e����2����%���byuP���Ui�>�4bc]`��Bni�)�EeN���]$�1cć2+��ZyS�X�nƢ�c6�Z�r����L��5T��L���^,�w2��@RU�i��4k����^�2$D�be��C��r�g#����>�~\�>�u����t띹��³"H܋��W	�:�0���vÐ�;��N��2����w���6��d�H��j׊'��FP.O�&��y�6����cf�r_��T���50�+n]���d+ڌ�k�\a �\,`S0�A�`��	���z�p�c �J.���>-�J(�\��sg���I�[u�Q'�C�8��Z0'�􎬮ܼ���A�\�Ab�q����uḙ��a鮤rS�(��`UcD8[��D.+�1��=!����EF �5�,A������ x�.+�,�����~��pssW�W�Z^./���Nq�!���1w�2��!�E�c��E$����攸*;�Pv3����'�/�r�ܩ�+Ó��e�-���,���9�h�۪k��
2���RE��<�8�pD{Lr���JM��i#cv1I���q*�E�5ѥ�F�M2�q�ٚ��T?7��Z��h�DX�u Aq��\v��uL���z�<��_�:�����ŏjU�*۪+|�gR�qf�V�f�ON���j$�mD,�+�m+eD(a��J����P�R٭^jl���P�2�j,+{O���S��`~ю�,�\����������=��7J�l����jh��R#�P�|y���'����iDrs��DJd"��H^��ٓʊ9/�o�t�y���]A�ΓB�Ke���j�eA������SB�5�~��#y��kr�ׄV�i&�ۖ1���=�!����o�}EN�,����#���A��1�������3�)W3�S���A�����WMo0>�;�O�����O�u��I�nc��a{�i�r�*[b#���2�RmG\G���ʬ��!�,���Ěٕ�*����r<I,��f�x�`Y�S�&�ӥX����)��>"%���o�|Id�!����a�}�^��	
c���몢Zfwt7qY\l��p��l4�Y8�KG�.�4f7�m�"�sgQ�odyi����RǠ�Y^����*;TMuK� }*���C8��_f���!%:�����V;Xu�;Fv�edd�+��_��a>�9-6��R6[�rbc�I�ЁD��7�A3ê�c�7;��!��;���U9#/(Q>�R�CAۭ���������ï��9)�	"��XA�l��������+��E�aď�K� X��iK�8�	��0�ڐ:/�	∌3���^"yM��	�+�t�d�LZ���|�M|��ikؕ�')����,�8��p.�_��[G*]
���{�m�8R9����fu�ҩ�7��+�,6����Mh�Sz� Jd5<4A�����Ђ��C{T"�K�j#H岠B��5ڬ\f�9�3�OI�X���fm0���=���sO�j�HQ}�A#N>�ki4����u��p����&##��V,���ɗ�����L3Ь=GX5
�݌��-+��Ƽ�(gW��2�
%�l��yPq���F�򨠖��n@��;9*Lj+����;�3�'B�&�젓y��Ty�M夶j{:���BŲkT�T�QF���j&�Mnp	z�s~H}Pbˆ��l=�nCG��)CG*GK�@]PH妫R9(���!Q�S;�����ځ������+*xQ�����///���e���Vm1ܽ�zc��l�Rv
d���s�p^;�Қ�"��$rK���UD�& �zƢZ���ή9M��Cf�8��@Q%3��_`����N7M�Ys�˞ߘ��BXݸv[�'$�'���1	��dr琑��FX���r����@5N��['n�lmN�%��0�Ԟ���n��YjPؼJ�'@T[a�ƺȨ
����AEn�fx���K.7UN<���*�����s2���~����`�dZ��;'P�M�PϜ�0'��ڶ�N�w���g�^b�������a��\� ��HԮV�����������eĊ���]2��$�(��3<��r}O���zտ�x�����8CR/
"���X\!��8(R5Q�G9��"� �/E!�E�Ldp!�2D��X�e}��o���F�^Qz�!
�v8��:%���$>�}�C�/����/Fm��7�'dddt�ϕK\�f���ˤğ�:��V�+�M��*���1Z��-�Hotp�~�I��W�qq��ѕ�Q]�Q%�|1�m�J.k�u�D��k4[ҤT5�,����ż('�;(�$`�&e��en":���zxl�Т�z�j;�����	�2����CVN�ь�g���Ҵwf|_r\m�Q<J3�mڙ����X�v�������Ȥj��լ�ge���S��=�៥ld��+<>>����
���ʇN�j���nK�[�K��#m{pwL��m �k�0�#�	Dqw1B�s_!�c	 '��*��4��,�c�^��P4��� �2�7�ώ�Z��n)���>��)##��a+�r
Y�V/�%~X5c�q�mSf2}�Ji�u���}�Ǉ����wl��g�h�В�Ȼ�>Ƥ����ޑ��}�=����j#�L3�s"�L��^�VOU���Fͷ�P�1�Z7�|�Vޣ�,���4c�q������)F�_O�%`;,�D���C�LsWy�4���# ,�� ���A�n+��`r���ֵ!�Oz�7Ԟ���}>�l]���Nn����&"��mN�!e���3^��-�àq?U���8ȕAoPS�(��{2�&̖u]\G3��G���/�	�,�?����	}��aԵ�r�����E���ݛ)��V�=;���|9b�/n����Gᘉ���gdd| ��Z�K=)(1^KV���l�n�L����+A���<���?>�_%�(�@69�k!ZI��Xq��s�3�<);h�Ⱦ�^�ˊ:�M�}�-�V���M;\�4�5?���^�>s(~���BmԻ���1�T�2�<"v�8)U�G6�a���[�
eO[ɍ��Z}5�?{���ddy[*sεo�Ykz��͛�����SF%S�i���L2�\�T�sTJe2I� �رcM|���Q&u����w��
z�/�2����締�>���b}��V�w��6�] \ƗQ����&�;$��ú�2�\����v-�b�&���L�(�rke�5�S��w�Ռ�ł�T�.��t"��^�}�H��O�6�t�C�]��q�H�3y&5��?�(���*)��Zk��V��05o�
�e��Ia�i����p`F��FpW3)RsȀ��q��`d�?�b�����:/�E��veg�h������ �2Bg������n1M����l�9�_���mo�~kOn��Cٺ_˘~f^��t��~o6N�3ƩEI\^����-ޓ�8�ε��!����Ƅ rJ��@�������Ԣ�eB��-P�iqR]O�ɩyi�K:B/7f7E/�O�Z2H��2*W�LV��𶾽�A,�!�������H�lj4w�$Y2�-p9���#l��Ҭ�������2��/ X�N��@r�vx1�h=j�p ��������&�r���j���ټX^`v^�}�OMi{WR��{�}%�>��]Z=��`���ǦT,ߌ�2�,Ιpl=��Zk��\�f��^㦎}l�y)Q]B������ޘ��s������������%��&g4��ܛ��3�s*8���i�}���A?�>˩�@掔I͌%G��٥JHxH�X��[-`�8��m^�u�ǃ˫[tY�캁�._�e�Z����3aM�yomI��4V���w({R�:��(fa{�����'�,�l%���Y��\�����q��{���R啥���խ��Cs�4�s�?~�%`�b��V����ßջ��=v�@Y2��%؄Qڶ�q��ƳL�R���)xkQ嗳t>���nfN��S���ɋ�ٙ�qyA����Y�l6�Шl����<@Q�daS�v��ybA@~Å�����Xڔa�N7�{3};�ޚN������4��l��@V.��Zk�� ����l\�?V�0��x���ksyqiá�����G����(&��t��,2�4[H�8���^d��~�77��~��gs�_o�Ϻ��I�JA���8 ��IpX��=ͪ!@��l�^MZr�]���<�(py��ڙ��z���sX�h޹9�=�g����|=�h]����:�6������, &�I?w�hn6�E	??��G �<�?�ɸ���f�
���P��w������a:ޗ�{Y.�sG�R+������L�'3��^�zu-M�bk����2NY�I�
fn�~��QJ�۬�_�ax���8�{�1jZ�@����J�O�^~�Kܧr���3�, ����A9H� ެ�Q�x+�ǿl�.�q�Ȗ^ԡty_��k����-]���2�i6=�o�m�oj"/�|y�򦵇�/ =0����Zkm�J�se.4�E7������'�Y04�w�����\^^���s3��|;� �d	9
���4��^���}��vD�"KE�BB�c:������͍_D2�Pygg������;.�]��0&�˲W�4M�i;�ssK:�-�����s#����f���hW��]y���ϼ od��~�Xt�=�����b��=	��.H�<������}���;�ƣ1�o���9��V�,�g:�\(�3+9'�f*�Z�O��ɴ��i�ޗ�_ 0ykg�|�l⵫����Ȫ��<�-{⽾Q��u�N�:4"��~Yp,���ʣ���j�]	�J��Z�\�$Ε]%+P}eWqk�΅LK���9h��0ǅq���S�+����R�"���S��Å�}̴���-%pE8V	dM���4��#�>(M��_�G��M���͏����BFoz۲�w����R�&Ӑ^�hg��׻��Z�5�H�a.q��̖0�D�Dg�4��ޘo_O���wZ0B�b0��E�0�{~��2�D�w�G�aQ���'6RG4�Sâ�ϻ�[�����-����Y�B�����yg������.-*C�54K�磠8km��tJ�I�^�~YP�����a�/�y-Cw�]�ެ��jm���c����=C/��w�R�~�C�@���9��0g�g�����ʐ� ���:r�o�o�d�ɚ��y�f9�{�c�y?`2�pL>����X�|����|81�GǼ/��.Y��j���yk?�l�il�( �%��&���ј��Z�{�F�j5'�_�fɑ��ׅ�lÿf���4˘���
�\,�$f'>\����h���c���]ђժN|G�.�-b�oj�h�61���?e(������kK�����;�35�̓�܋]>����<��`��O�C�u8��]1U���i=e�!d(���\L�� ��Ti���Z�3-�t��+���NOO������F�� ~�"��a�@�bmo3kh��*{��t՜�)��^ooo���	-�#N�E@b=]]���+z��;-�5p�������2�?q��9_��\��E���[{l��˵��]<��Ҵ�,2�rl&I���=5����L ����7z�1���|������L& ���rA���nwC�-�?�������[(�����3���������� �	1����~��Ks�J������ߦdI�O`CF�>G���#�5.�Y��~��_�^�}�{&�CF�E4M-�@�y�ԃ	�����'r��Y/������S��Ռ��´�(���L�|
9�P�+��՛���V��J4(kヌ�d�R�K���,-(m�Ub��c
Ci�I�7�������E��o�9�:�6������6���s� Y�vk��s:�����MA�p[^~�+u�"2���eHa7���k�c���]pIN��&H���O!�g��l�/_>���锵��B�2�[��@�6;;�fc�5������L��G��I`5� ��:���3�s����E%���f�������=��۠L���n�)��	sYe1�������'�5��x��������[C��VQ��-�~y�,�{�{ۮm��\�͆.��ܳY����&DF����ws��髫+3�N<�P��F�G��7@��:�}���4����h8"�f ː�Opu}m��,�#y��1�������욽�=�	���Ќ]]��L%k�!l�ד=�<�]C[�.��I���hz�Rɍ�[�<g"3�1��?��-Qb֕��N�9��HObq����~���nn?��Έ���mnp��ߘM�$0>s���,����nޟ)��!;N����p�e����Z|Z;�,T�GIv�򕣄��V�:�R�f���{�.��o��|\�>�Yi,&�8C����A�c㗞v����<-�B�8}��L���$\D�rl>$_�F�j����k����B�l��5�G��f���w���*���dܛL�$S������[���7��-�
IO�s8����k��-�2�F` ��Py%�؆�*څ�`2�ϵ_L����s�̗�zc������Ǐ�����T��J!������
��H�}qsk���=?��^Pǲ��Ju�i@y �`�6����c1`^$-cu׊��}e�W?rU�ZV)�ga���Q\�rN���K�YA�r}�U��uiײ�Age��o������_���aO��e}��������fwwǿ�!61���2k����~�G 1�X���뫫����x?���w�A�����͟����Q�0@k�5�����]���e�����u�Z=چ�s���S?T������q�f��FE�
$�Y ������D�e0�D3#��<ǜ[�m�F���5|��w�EF��I��0k"'"ӂ�˫?u���0����zI
�!�.�,K�JD����2��X��Ҕ?fpW��|�����p+���p�n��^����`��U�ӡ���褭"�Q�FcV�B����=��\Yĸ�n���QiuT�:@���F�����3ыdkwX��`�B[��:gܣ�tk��.{��V�����\쓜!�P�h���������w�����4�-�����iqF���$�+���1r�ɜc)�G����a�F4�{�����~#63�o��������1(ն��pNV%����_�淶�=�:��V��{���Y��<({��9˂�M��9�Y������E�	O����Z\��n��I}e�M��a!'�	 ���Oͅ���{H�[������ �bF&�`wIK�cj��)� 5 ȇȘ$�i�]?�$���a��������1����&�1Ȳ�Lƻw�T��6j.�,y^'fR��W�t�[.�h�@��_��d+��5m���s�յ'm�aJ	����w�S �ˀ/�o9� ~�`��t�#�����e���?s� 9DȦ������+����M�#�w����Əu]
�a�r�Y(꧶�c�t]���nM��[�Y�b�c��]�W$�hm�u���4�@�ʗXf����?����hS9v	gnb�`����̭~��c�����}����aL�|�_�e��d�a%M�&�D�����Ny�Nbvf�e/q��E����� �[k��7g�[a�)g��љ�V2͙�i�������P��A�����w�p���"}�cU��q+��0��O�}�3R9~��G{{��x�"�_܂��& q������{���Ŭ
,$�P��=d�k���u��2a����od4��W��6cU�� ͯ�JY�
� �/_���0�ф@��9`22��s鋽�]���Ѽ[PF�{E�;���# [���m�H��|�-�Y�� ����-s�}N�K��� ������B�0��Ff���N��68�ԦmOZc{XkK/��(x$Ɠ���#Z?�L`� ��%��j�ɟ$,J��s���^,���-1�.�FȞ�a-�u�2Z���-Y�g� �6����Dh���G'\��(�ajP_"%+�V_0T�{@ԭ�;�4��3���.EQd�/�5�\�^
=>�(1RUn�2��&?�ތ���串 | 5������'w9��\�~���+]/�_�l����]Ry�E�lZ���jd�JqJ�Zk��V��]pF��b!c���!�_��|���`e��y��ļ;~g�����./��mI}%��N�'��*�L^D.L��L%~ ��?��XJ ���8"M�;������ܚ?���,�̸��օ`����"���a*���K,4K a����n���9W��o�H����|���k
:������i
#�����o�Q���� ������Kk����a}\7�� +g����Euxx@2^�c�~\QV�|6��'����(茬'\;:���h��Zf��i�b��E�YZV�/�Xr�@D�G��OȷM�_w$�`��.��F�k�̳f�,�����a����G"��k�5��ףk
�+�%��Z[��2�j�:�ķ���Hp���k`�@ٖ�N�E���o�@m2�6t.�G��rg�>O�+�z�6�hI^e	�\���y'3m����<�y!�)�k��*X�x�,�b�ԕ���gD��0�X���V'��3eY�5��m��H+,_��1�9O��Zk/o.�?�}3�D�}�|�J -#,�z�mx�bX4����&*Uu��06�p�~����Eh?��ͭMbOC��//.̵_�Bw��X�B���i<v���J��>8I���e��Yz��R\.���D��J�ִ��Z����׽;�d�C���V�� X���A�(����u{f��GG����'�?1�^�A0�i��~
�T�~-I�̮+�׎T �d�S�!�����֖��qf�ξ���[J�‐� -Ԟϝ�B��r����ul���^�sgzb+uJ�p_�������6�F����ngC���8�r?mt	�״�C����20ސtO�Kr>x]��NgZ���X �5��.�$������w�iK����ꛮ�Ve-��R��9h�o5巾ˤ�5�/ y��7�5W�B,��Q�B��yP��*�V$E�hs>Xv�JN�@.Hp2X*���.s8x�:F����,��E[$(=���,��	`Τ�Zk��-s�/�����/�?�����syqN�"Tm�C	��?��wst|BZ�$�1���h̕�!��ǀ���)�hi�V����f[�)���Y�t�.΃v�O����H�l��IOcGq��h(�R5�-Q�v$n�.^&�Y�?��M�b�F���c����E[k�M�#����`L_��ک�2R8��_�����T{������ M�����fooW|��)HW�6[n]�C�k|/�����4}|��}g <g��$�]hl����-���4-����s��֖3��\{�R߹��'�r�}�,d�5�K��n�M�w��ap�ރd��Sx�%�v����C`��p���l��l� ���D��ՈJ��G	�V�ڄif��e�y�6�� T������I:4���O`+��W�ƚ��
���:Ʋ�2*��xY����j:����)W�����]Q$�1>w�)2�)�)
٣���G���@�v���8�7��[k��Wn�EMa^0�͋�O,�����|���`@Em̔�O�>Q����1- ���S�Տ�f ��	.��0nǭ���N�<� ��E�~�"#���ߩJ=X��ݥBBp��8[a-��K��g�yqЦ�l�s!�V۱��-a���BS�WS담�Uk���U�6`���L�2�����k���W��B_ #Lz�ɜ��34��v��#
a4:YG�d��\��;%�h۔H��?��!��$`��q�ߧl+��?���߾�s����)�O޿��4��Qy��/.��Km^�M����3��?��rԔe��#pA,c��gl�=!�(��(}
S���!$v��� �3����\�֖�2cY�Gev�E�U����d�cw=0�x�h&�j7�;��r�jn�u2O&�R�*ͳ5o��%�;���ׄ���vf�Z+����Ep���Z��e�:Ț>Ai�.���	k@�1��]��p)t_\f�H�*;�|�,0�*�U<��Xӳ���Zk����]�:�����|�����Mƴ$%�����'�V�����D�~:���8�0#,b)�c�M_���R1H)�����aa����zss����lmm ���'_��c�3�&���;R��W�������G��!
2kc�W���Z{n��k�GW�Cf��:���������R�����޿OzƐ�@�`�T���L�b�h�,hN̶��s)AG�@i?������`5�}߾~3�w����A������8U]��3^_��2���F������^����E���)�8_�a��	�a��)n䔥�w��<T�fR$g�=z��4&�8��x�X(x�#3�[{9+3��5E2�9�	�	��"m��c���=�8�Q�v�����JfM���B� �ʊG*�L�U���1眅Mw5��d>�,����7���۔Xa������L�!ʔ�00i
��PtJ@��0�-����0��L\�YZ�r��jD��)�&�͵h��֌.���X����3��>ܳ#��',��׿�b����v�N�"�T�C�,[�R�a��d-;
�#30���<�cӐ�Q����Bi���_lF)�1W�ީ�}�767������aʉ<�M
��sئ�i���Ps���.f<�d�h���Zk�h)�p�j/�~;5��_�#�)�I����~������%����%$d����%�H�Z:�����9�f�� �W �Q#E�)�ߟ2��� ������1'�R}	��BFѯ.��k[���R����[)��e�+��Y*]����3�JO�j�$(x�7S.�>��uHwBk�<ɂP��A����1�ȭ
��$�%AA�q�l��U�QSH���
	��"sz��F��W�vn۴�^Q�A��(*��Hv(��L��h6� P_���V���hR6��m�J���
�%����g�H[M���[���,�\�y�& Vڬ��k�~���P#�KXs��J` 3@
Q��M���Zk�1W�8��BA�������j�~	]�O�~#�2��c�������c		��xM���[b/h��/��Z�,�2�"�F0X������������N��ki��a�2����1��6dt<�A~DAl�=k���=DQ�c*�y f?��k�?b%�
�hsk���Z2ӆEBٰ�����_����(���{��=Id��-+��F�8c�T�eO>��r2�Bқ	�Hޣ�)� ��kH^����.<;;#��h'��`b���5��.�ɜ�V�)�-�[w�N�*+�k�sf�?%I�ry�@�#���<���E~��[@P��k���q��L����5���밚{��R���B$�tK_��ehBd�?��(�f��.�Z۬Ʋ1!5G?�q�45���ΐLª���K:@�E���KaW�<H8��\�����~K��V7-�VfS�bJ�-��������;��`�Cs:��t����T)��)�@�|-d�
�5��Y��5�O?C[5��T.�\�����>�a��~o� � XgQ+'�+�M������g#�㺥�=W�S��p<��%kk�����4�cN�p0$��k3i�E�+�� T���"���n�k�8�j5[�HR��7�	KA�1�q��/�/W���<�[���{���70� �py0��?�#d1��9bA�j�\�P��I��N2�	���K'E��s����@�5mZ���G ��,������K3��_XĭBvBaM�Iz��̘�����bk���R�Js��÷�����ՏA�o4��L�o��4o��9������ڦ¾
&k�]]�Z�����e�K���c�J��qj��Yюn�e1 ��}8ǻ���Ǽ��cv��ע`Q&ߞ�'C\B X��4��=J��N�ɪZ�.ŉj�AmZz$���\�jǜ�ED����9�J�p�D�L�=��j��i�}V�PM߬	
��y-��Kp1W~n�^��vū����l�V�3��Q�9׳�1�"4l�Iv����P�x�0Py�JYd.)�1�Z$`qF#k8�f�`l�o���r������)�G��� p�O�[p(z4 x @qw�J�3!�;��	X��T�	m'eg{k����<�S�,�idT�"��̓#����=H��J�|-lr<��9@Kh2�5c�����o�������nL�cp�P,��Yy�
�e��xϗ�1�۪^�I���Z[/+��k`�`A�������ڡ����1�͓�X*[v��KgC4���vKqQ�X�����Tc�:���>��h+��{wrBc6�I�\���+�Ģ����.��)�T^�[j�2�tѝ%]�p] +������X�WV��r,�	����5�D���
��Ї��`�(�+�߰��Zk���ڭ�:ʊ B�l��&��n�FomU��
˟1���/_��o@M��K���>��?��2�yY���"}YX�*�G��M}�g�w���~���9M����$�f6ָ������N���YW�1�{��e�g�����CW�yc̅��#β"��%��Y�2/�ݖbۇ��K��e0��2�:�>1f�u�:*�e\O�l��)V�ګ0��ZZ8�y��R,`�1t�$u&0��0A�_ڹ�Ҷ
N�e:�n�><)���@eA1��m3�X[���QL�Z8����}��6��#|N�Hz�F���-�O �S)&�
��YCt8H��c�Dm:�֦���M}��áh^N�S��V~|m���6gg�s5���+��c�i���B��������
ߟ�Hy�����=zcww�t�{���lm}0�_{&�k=���t/2j�72�RNq�tp��*����K��mYx�W
�Tc�����۴:?E�B��4��9��e
�u{����/?�E׎Ӻ���>)��N˕�I�U�}U�D��Z�1����K��<����m�s���o��$����w�#��FRL/�9�t��g-ן���Z{���2 �f�&LP���/��nM⧖�c�Ų%'�[�D���͜������=����z�d��c<�U{���=��v�zݖ jN"�H���|/\�������'�Ȓm�R�F�Taf����|�X2ZX��J�`�ڔ������X�
��|��'-��`H ���.�{�.3�Mdk� h���{�_�hW�3�b�U	cNq�g4����X&hj=�:�����.ȤV��Y��L�\ʖy�|��������G�ǘ!�EA��t�X��WS�n����i�X�HAWR_�b@
a~W�F/T�W��0lSLY�A�K<�p�u=Y̦Ʈ,Vy�U)���B62�S���)H4����O� c�J�H*iK�8�dJ# �߆�_0i�M����^+�:qN��`bŏ���F��S�e������"I���C�'��v�����!=I��˿ooo��o����i���`�i����<�N�ӵP=�D��-�$�
N��p к�vީ���gZ2�	X���T�~�B�����|����sgz[�vz��5�N�ma�H��A�H�9<�ꪌg���Ė��k�����꒦��[k�M[2>�2c���r��Ҹ>����;{�`���\;yWG�2CJ�b�2�5`�"P��:�弁L���^��&g���Sg�wUڈ�����9:<��=���/��NK�O�=�丁i%�I�ɵ��Ӹ�K17Z��V�L��
@Yw;�~-;,Q\nYѭ:�ߡ�.�|,묍G1Ӈ$شr�z �y�c���|\��cɲ�X	s�xk��:z��^�:�+�V�I�w4��Ż��G��{����*�j ���`ٝ�ҙV�ĬV�X�6�}S�o�b}(������f�뛛[:Ob6gE$��PY���||ܓ��}�Q��V��F�!"����	�R"�L����d������d�Y����>?�p��4����\��P����hZ$(Q	\v�_%���y�֙}˚�h*nln0��~"�N��0�H�ׇ�k�V�cf��JWг[����Az�~��'~/=�I�x?%P��ʓ)1�þ3��B��i��0�"�! ,��x$��$0v�̉|�̅���������z�Z��A�8'�'�R~}'��[������O���w�B�RUm�
���)3ͧ�z'�S�sU���z^��m�O��Td| ::���\"IX�(��7�����w�ĂעQ�����'��cM�Zєg���T��N<�k��Z{��*��0�8��+�x�"
�c��?�7[XD�$����A�Θ:�6:���gF:�v��+}Y3���f�/�w�yCWz|5"����5/D1�i*V]�{EiZ[OK�ԛY�9g�%�ˋ�j�C>@�f��������W�T T���,2�[N�[�"��$Ó}��WCY��B,�7ۑ�,e�?��ۻkxWg<��9�G"��������}���;ZS����p��il0�K@�S����دMwv�ͧ�h�0~ѥ���3�M���*�O�F�y��r�rzL��p�9+e�L�Η=g޾y��[va�[ơ���Y.<7���4H+���/7�?��ga��+�\�]O�ԽI��e�(��@(�k��o	U�X��PhG��$� �ʌU��>�y�t�B��%�e|��꒽n�d�.��	��i�8*2����I���<��Vbc��"����쿓9Ћb,�k�>(@ϚY��iD�//����M*��m�����qJ�&&���_��.>U�52(C�c*2r	q�� ��Ώ�5�y(aU�K�c� ����{���GR#f�Cn���k3&���G7�֚��~�@�����jR&*/� �_0[^ˁ@W��4:�Zk��fK���=��� ޏ��pD pcc���X`qT=�)Du���F\u���CγcdqLt$C�+l�/α��_s�@�s{k��%�_����s���;ʬ�=H���ެ0@� ��X�����mg?�<���*3�I������4�aM(�	6��x��aM^?�<䠫}o��\!<�t8^Dz�.=JL)���~˾֕�:� ME��=.���R��~0��H����!�v	K�)����V��r����'W։M^�Bt�OI�����\A��~�:>�OG��~��D-��e5����W�b���W����W=�&L�^6g���"���4wѳ4g�WD�q;������c���o�IH�>ո�wy�R��|_�x�+Z���7@*ؿ}C�% �(�FL^0��	���WK����3� �N��A.C+6T�*J,�11(Ȓw���lHI���h�pH��N7��2&FZ�.�"�`B�8�^�lm�rc)�G�R�D��1�>e�����ن�� Lx|���\_���;8�7;;��d�8?g���� ��S�V�}.�����R�A;-Z(Bt��Yv� Z�L���2f�8�L���8AD�mH�^@b��>��njD��L
H�0POl��e4�<��
2UT@+��E��Sm︀��r
4����[k���b4��x=27�7���ʏշ4��;�;����f:0��VdvL�ٶ��J��G5��*��!Vu�h+�a,�\���-�7h�CP������n��n�_��T6TN����{ ��g��T*&�f�6Z�P�QԉA-�S@��ħa6��E�f6\��g�og�\gi%��d^_[q���J�ɥ���A�ͭM���k�v�K93/dah�b�/�&�b�2��� �s͉1�-X>?;3���ϰir��z�AF�CĲ`��`*�ڂq꧛�sX��b��Z�)��c�Y/|�0e=5!}ι��V�mr#;��.��akh!fQ�K߂�ίb�E�S�cR��b�ATb�*��$�2V�P���4�%��p� �'tr�I�ײnw&O�%vل~��И$#���m���h�p4�m�J�G4I�<��E��H_i�����Xl�ӠW�m4I��d9�K�:�c���}C�2�|�?õT���by��T
���.~�P�K���k���h�`Y�>���lʀ���
�|<b����Zxp��R��u��
N�c����YƔ�x����h���~IS?���~��k�0����M���͕г,�P5����=��L���ì�+ז~4�U'�Ze]��ԏ{���ꮹ��P  :�?��(;�XJR; ��t�����·�Y�3��������]X����w^=V��t�z&��[���*�,Rd���p��6dP�(0J�%�/�	K,�e��8
+����R=s@Ś� �45�V�ϼ���֚,<)1RLv}}E�*g���Nל�{g���� ��4�߱^�����<�e6~�՘fB0����kV.�{}=!����3"H ��un��Y&j��
�?d����/�쭍%�\��	�nɜXz;y�*�;��F��pڏ�4�<:��f8j�X��ޞ�ޥ�P ��xp}Ѩ�Li�	�t0�E�&��� p�}^e.G𕺺�`5I�u�X�\Hi`����FY�;h��ޙ���	И�Jd/T3���I��r�D���Ȓ	)P�w|�!��ؔ'p�-Z�!�O8��X�8������Q}c�M�� ���0Y�'�26x;jg�j�У)Y
D-k�Q�#ۨa�{q|Bfj����� ����)�䮧��s6yVª��M���L��X��-5����v�k��_�x�
�
9�]a���LE^�t. �s�u2W�,D�a���3}0_�ԐkP�U�7��GVh����H�Z�������V$���j�r�W ���u�����i��N��k6�o��$K*�s(��`4.�aA7�Go���N�MXo)xSC��X��H}"?�8�/���<�D���IA�jnA�1�3��H&�ea.�Wrk��p+uNXz͑�?���J�)Y#��S_�)�+�Y�*�k"SZ��,��r�b�c�,�m�@kK>��;ٸH���@!�p�Mk�U�l������r�ʺV�٧���:��/}B�y��FK��g�f��l"J�t}����16~���n3�������`����k0�`<�u���r�z��6�~,��:��o�Y\���ŏ�jĭ�;x��k�>�����Y�"��s�>���&��=�����.E~�	�4��j�������<N.��Ƙ�Sw�k��k�۟i��2@��3��rf�����!��
���f���@wX@O��bMA�-C�b�.<��o��H�
E��|�b��ϨRm����u�T{�AQ���8�9�����,iE(��;����"�j��vwwon�n|{�*}i�n.��������Sa�<�&E�r�n�
 ��O����6�'���ʢ&j@���̂�HaDu�V�ŢK��f��Q�
�,��ܿ�f8 x=��gD$�cFAC��(��+%�����sS3N���H�i���,�~U4��pQ�ܴ�Zk����C���X�(�q�T�7� ���X�?i��@)�}�����,��_#�	����&�O�]h�onn������k�`&Z��?[pfaA�e� ���sam��"$���F1W����\_�B�]�Uɡ9�ko�R���`���I�r��$�R}��h�~f?�ޯfg[E�>-��j���,�r%8�e�j�$�%y�6��l�F�cf�!�ZP�9b|��c�TSi�U`V�8�"������U��S��?.������I�.�Z#��R�B����T�قi݉����2�vƔ�-��8����\Z7$D�ft~�/-�亥Ss)Ԧ{��
����:!w����(����5�`�g]�J0v1��rz��ÖB�,�Kb֐�9�{ɏ�:��V����2+E�Fa�� 
Ç,�)I9v��H�m�O�F�9$3-d/�Gm}�9�ˀ��o��_o�52�:����.�����#��h%���F�]W��՝�Z@��>w&���ń̇��2L���W��IHn&�C���3������P�fNG�g�_�����p$7�,�x�E�0)Ǵ��R.��D[��A��[�&^�S���*�b�.&��0�+�!�X��^NM�u��"u+D��\�Ք����OthlK��?>��]��ˠ���b���%����/��j��\�o�x G�!���Q��	�9D��x�ḋ���P��E��}�¸�Ngڦ��i�g)��1�Xڦ��qs��R�ccǼ G��<o����/kc!�1�ykJa76���I�E�eX�������*���&�Ef�^Sbo�9�����4�l�"?X�����R ��1N�`�f�,2kbpM��ggg����|?7>����#��V�?���,�a<'p��ֻ�[�`iq�_��Tt��'��L+�]�bR�ј V�9�%c.|��
��]\¸S����pQ�X�8���Q�}�4S��"92b+r�>L>e'��]��p���;�)��&}���!��yiq����5"��Yj���r��<�����Jx6m���h(_~$\'�F�OZ�..�W\�:�L��Y��Pǥ�rvE |����i�&�p`���#@���򯡗;I�~�G �7!_�I�[*Y����������R]���l���ֈ�o�f�f�⾃��3���BH;j�:�^3���~s}��y|��L�;�_�������Q�	7SW$�/��~��hq0�Kc��AY	W\���[����HP2.�ς���F��_�.{���L9+w��l �P��V0��0��]Yf�K�I k�M�=�^��.�O&�~�����hf$��ڟ��lBMNu�1�n�^�벹E��,��3
��	�d�3���^c��yhM��K���t9S*��'7Lb;��T��X����/��ys=$'?V��� �a"����< �`_)�ܓE���;q�I�L���p {ݍ�ޜjJ�"M��>��QM�v�zJ��r�0������X8ݹcv]�LI�c�}a�L&�^+b�T����D-gv�]72m��y��ax�h��h�<�i�����q��*�,,��E��~�)[{��LH��m8�1s�	-��H�y.���.L��Kuy�3�� D`{h/~���|?�N��5=��51d�Ck ���� ��,w�"E�PDO�XL*�2�ʠI ��祉���������<��W
4�28�]��o��F��Z{FK�U�� �p&�N�}H3Ǭ �]
�l�%j���w��{�����`[���������ɨ���
�载]�I�A�lw{�rh�/�6}�����6@�����w����2��TDm
��a`YX6�{���	 ���2ԟ�?.�V�I{��LK#���2�gc�qj<�'��ݝ]�渇8���m
`��+�~qH�]�1� ����_#�,0p�X�H�{eH�Yؐ����<ԏ�����}@X(�e);j+� 1��� 3�Ie�1r_&�p״�rsp�tg�̶.�:Y#��y�砲��SH_ٯ7�\ԑ}��� ��g��3I����&2�� 6�E�⺐�ʬ�g$#͢�1M{� M��0�%N�/�������Pgϰ��:����D ����m�R?���1A����� O���<9��3��3�I�Il7��f��!�s�?ku�5�o��o�, 0��<孱2W���S�򓜶���xz[��JmH\�2���`����}i�! os�GT6��/@Z�@'���w��9�i�"�/���a�옕��-&�C���߼#zc>������e���Q$��Ή�CR����t3��tr��0� nqal���$�!>8�#-�9X�D�Nx�s2e�޻����<��B?��˩��N��֦2x㆘Xp8a^�Cґ�U\�6 ��b̘��f"B�_�0�u����R��|�CC�/�᜞�}��O�����!�'���&������tH����ނI@l����_(a<T��f��$?-�@�2d�P��Y����Q+�@�`�`3���0���Pyg����������Q	�^h<�d�b�7�����w��cj2U$��N4���~�Ks.��A�	�о�q2�rZ{+�r`���rg߿'�}P��r���g~��ѱy���Y�����x�/.���Ս�׀��>�r�����}���	lA�??;���_���#}����չ���� �F�tV�_����!Y��c�����g�����'�/ ����j�O��G�U7���\q���>���9��:�~F�-�m��I`D}l\���C����8���V&?�r���t�!���۩���y����/dn�������ߟFc���G���x�Q`؏� ��~�������ڋmq��~3?. c#ڠrx�������_{�u���gz��V���߅������x���SM�������K1��+su�A�WXӐ̞|W}w�(�5����F�\�>����R���.��;����"Sf&���AE�|��?�`�vx��fe@(�h9C������k�c���+�]6!����b`L֋87+]��x�c�-41��������������|��oK����#CB	H�XG�@;�����;�3>od(�?`m�ɺ�5�S2d���Q��kc��&)˲J�/����u�S�'����k�-��hw�l���b3�6%�$@S
.=6ck�Gm�$�q4������aM�s		�Z׼oȬ����"n�{6	ڿ�ߤ�L�Ǝ�)���E������0&�3��E{�zf���'z�X��*}��3ePed�6���'I�ߦB�!��KF�������Dm���9�R�	I��:i�!���w���踞+�9��� +�\H:��%
�P�9�jH�
���W��;^�G�4���[�(*{��e���pu�0B\~��}k�6�Ԛ�0Y����~���f�i�K���l�5��!���� f# ࠷Y*�Z.D�&k��^�rR���|u�M� 0#I~
@�H�Әa��7��R�����\�m���+EK](���eA�dd9��0*�0�oi�le1kn񧕅��?$��3 ��uB*�ו���5�ep��U�Lٟ3ޠ?�DF��
��3�{�!X� hOޟ0`	���3ߨH��5���0���fp?��׾��f,#0��X�}rOpBf 4�q�`c�������o�7"�Ja XF��M �P �vyAׇ��\[/$^�C��;?~\���� H��[��}b8^^� �U��NtƘ���8�m�˗� ��2' �;��;��s�����qMA����\1��6죛@ʘȿ���� 7�ma_�Ѝ�QN����b2	���(��c�fD�"�W-�c	B�� �����FXO���a�����E��E2��$��͈�D�=� (c�k�� �Y�'/�S�����]����G��pk�y�#�a^����"����U��~��;]f�_�И��c�j/�:��n��|��v�����o �im%�ˈ�W9�>_��I�U��ߏ� K���.�������p����ȿv�UQ�t�׬���L� ��:��晦�q׽�Y�	��X]G�E�v�t�8j��3+Y��w�[2㽵������j�`�vX{�7�s�zs~��Y��-}R����!��.8RLUL�����.�!?i5������%p7t�,���S)�`P�p�?I�?x_� TC-��H#C��&,fT��E�Y4�E��@�TR�C�Aa+{Qr�bQ��+���JA)�$[�nB�b���R2kq���ae�ᙉ@���!�e:wD�ҁ'a�Sh�sA�O>r�"����Ė��T�[����_j�\�3~z�uT϶ff��5d-�Wk^�������lBc[�s�c�Lx�1�i��͜�~#����1�5�D��5CF�\)ŀ ���n�<S���{JϾ��A�F, �`q� �f��Ϋ��й��a�����4R�����<Hk�c��m�M���ԁ �\��i�=�=����Y8�ҋL�tje+�`
���0� ��L��Y����7�~��S�����$ Y�坝M
�`?��~A 6dk�����aaB�icG"�Ƭ��|�k��|NT��6C*��&����Տk�'��R�����L8��x$�`���1�Y��	���Ί����X�sQ�dw�t��(6�g�?�^��g%�,������#���N@'�G�N ��[���<;��'r?�a�����W�Q(&� Ӹ�ְ�@cήc?\��Y�`�.2�_��:���NS���V��q��ш��޳Fua�����N?�7ڈ�ʃ�*~�(�-]Ah�;�(� c7&Yf"Mc��b,:�~J@0�%��P����J��j�&����#i�e� ��`�����$���}*]��9��C�A��X���H��jAt�,ڵNOP��Ag�a{�"�����b�,"�E���5�h�wM��;�G���1�־\���˲y1'��KdZf1�`�@8�����+�X,5���Ȓ���� <�X���7`Kk�
7}>�ƨ�ǯ�$�[��T�6�����&9ׄ<P{���r���Z�m-ǌ7ev��`Y�����̬f�J(����PFP9���NȘp�k��L�3h2y��V��N���;t��11�(�T��,::�<#�<�? ˥#�]=~�@1� @-��5]��#K̆a`�XK��/��bH���iqG��_�wdqD���)��Eʵ5Ҟ�>������T�}�s�̊ �@U{�@�8��۠�8"}B>D�{��0PN-����Q�<��x*U~�ט�������;2�d�^��f}gqjG�� _�Q�{�fPhW�ϋ�}��Qd�=�?�����f�9GK�R�f.8�Iwl���M�Q�kT�SDy���,��J=>�� �����~�������cZ���wQv#�ʊ3gd��
#��q����f��;v�O��5���͝����T��ݤ��dЄ�~~��"�x&Ѯ����n�w�����S�|S�V2���pq�B���:�It\��)m��U���4>�xVHqq�"��w��K����j� G��0v2lh�/�A��)0��7�~=���o 4pط!�B�O���H!�/_����Ss 8O|�@Af,�BU�Hk�tv���C�h7��Ǯ�> ���͠�̾�!@��;;!��sd=�.�T\f*�P��]���	���܈��wb ߱N�� ���_ۭ���]��l2&-�(�.O�H���x`p`��	?�,@0 ��-�w;;f����T�L��<ݾ�6�gg�����Z���ofO�F@��a�[�ֹ�R| `A�0?�tbZ~G� �6���✮����Ç�����a,��x.�Nl�&|��ɜ�l���W�r������	� W�fH��V�l���i���X��������F���]�볛2��f��0e�P!�X��l�8�}��x�S����kAh�A�9�����[��v��H�	?~\s�}Z�8Hfg���S?�r�2	>3��T��L�����?{�3{0�����I֊��f�'��R�����"��nP���z�rǚ��vs��M ϥ-��ER`8����ॼW�:!wy�@{K����`�3W�ʶ�ZW~]��`�����U$��(^�)����]�_�'<�ن�,���\���$ٺ�/4ݨ�ݤ`�������k�4�%U�.,Q8�S��q�%L����rW4��?�ml�i'I�s:�+���y ��I���b}$�I��S:��QH";�B��<�"k�z1�j㝌�:2�;/��NJ����9_�7Ұ(5
�?.���60u�X�P|��98�iJ�8�pBp�Y�� 5&��P�Z��4�[��R���2��f�dW���wlx��H`��`n�Ǟ]��ȸkK��o]DOb-��ֱM���ׯ(Xv(�4g~$2��+��aN�`tO�<�	GX)�ɖ'\V����|֦Ϟ�x�k�5�D�TÛ���ITxŃ�jDs�2��]-ȩ���Ocx�^�W�U�an֢!��	�JF3 u��9���y��ӽ���nA���GM�b���g�%X7wow�$ �L$�
D����q�|@6�?��o�[ Do��>����|,*@�LS�8�?�	��6����NjY����%���w��l�2cm�J !��;91�(l%�CQ�~o��'��3[� -&����DQ-�x�?�?�����P�"�`Jv:�"�0	��&���By�N������Q�!���{ ��g��������P6�J^haD-nH�C�H�D� _ջ������Ucyܗ�U�
���������t=I�[��@yp�^�a��s��@��ݴ���6�a8/1�"{:� �蹒�(�ٕ�sZ[#[���X��%G4�;"t������9��E?�|�%٪,�Ӕ�G�L��
��t�c�Wג��0T K�M*�c�W�=��qOY���j��ݰ�+rWt�/�"3;��,k�'g�2_���P��5]�0�̃it��z��z��su��p!R �f���z�p=&�0=N�E��u����wI����*A��w.3�D�f�^snB��6]�RO*7�œ�s
�a��$٭�\�p=����W��Y~�R��>f�>��f�c��'����lV/W@I����Ӆ���0R^�O)��1oX(���Ȧ
����ӊ4>*�7a`��^`be�� S�����W|��&7Z��W�4n9%M�dF0�k�hXu�@�hL?��e�!B+gb���R+�k3$=:�� i�>^u���i�`�P`�	������vJ���<��jl��� ��W�z�4�����E]l-�s����i�e�+8`��گ7~��k�ٻ������E�!0�!�D'~.���^�Nhd�X?��2B�X�����1�sG�8Q�V��)q����9�#�P����<A2�}�3�� ��=X��D�#�Y��P�'6W�{�����=e�� ��(p�������� f�������p� 1�FF��5�t��ټ����O?�>P�}� �= ]��W�x�9!F�D���H��,��V0F��_�D��O �T`����4�{�$� @��Ʒe/��Ի�c��������h/Æ"� &$|3\��G��!�OO�� f������_���=r&�|�&"����dI+���A�x*�p3��m�8����AK�"-��dL`�ޞ領�t��i�z��S�������ʃLƬ�l>_��O&���1��zroI�YdY�|[�D��̒8�!�������I@��A�i"��g^�$G�4�*�}��7nc%�5B�@�'}��N-�I���P��@����p��alE�3�����65��H���$�5/?����l�8R$e=�^�6��+NP=��)F��ُJ�9W
����a׺y������ ��I�¨f�ؿ�����}����ߋY�&�h�MF���r��R�a��R�M&[��A$��|KzϚ�mkoښn�����
][~1iIufݨ��d�w��I�2Sup8�~b�����Xȍ͹�>�����{f;�,�}!�1G��8f���� +�-�bC;x�͔�%�ΙFxM�n�2�a�D��l��<�a��F,윾��
��O�U�SN{�G�4B�L����%�����E��8�5��H��!XL�;|>�&����e�!������H���,�Rz|��+�4��kk�`��udA@G�尵KF��^���ę�#m���,2�T !���Z�/LY7�Z.6ƺ��ū��A&A�JV0#h����;� �<�c���, iAW�ŧ�R]�>>���q
,��T/�S��!@I�i�Q�^gym���gg-7�����Y[|՚�.�wC��(}{o�
S��3Y3��I��X��\o���=<"6iF��P��F	���;�	;��B�S���-,���(%vm������dz�o0Y�N��Mi�M�;�v��ұ�`� �>�ndv-�&�F�~��6
H��2�,�\����(�����Y���>.Yt��_$�FEA�$�{�$ƝLr �q��/���TgzBc ���sb�c�½��؆��)�w*P&���BC�k">���pM�Lǳ��w�{:�� H����wI
@� q���S�k����l��5��w����k2���	)�b�uk��Wm� �,��d�.:�~��lQ�<�h���|�
�7`V��@����4�b�i]��3�A�D7�h�n��1=��$I�L2�2���-I{��0�gj� ����J'N�����V}f�+2om��S�g��}����% �%+C�Q��*�q�T⸏,��~��_�֖�,}�1B����Aw��O�ٿ3�w6�T�#Kfo	�93��% ��z�Z{{YƲK���Y\��nAX����Τ��GZ;�V�>f?�"zS*�0
f���+��{�A��5/xhQCۢópyH���"'fXfa��ʍ�QK�9�@��z*kD����1� ��B��Y�RD䦢}�9hA-8A���H�kNØR��#�&���,��ɐ�	�q��n��򏴏��tt��+O�Yi(j����`K�^U�+ZtZ{}��s�e��>Y&��j0��En�b��ze�&��c��/������gա����B�8v7ٺ.x�����`p�4�]16C�Y�H��1^u���ρK, �.@L����]맵���h'��&.�,�~�x�_F�VȾ �T��{syyE 2|6}�з ��zp ]�}�CQ����Y��e4��.F}E�U�m���2x֡��>������1Л	� �. M�Oh�H`8�~�E|wo�~�FWO� ��{sSu\;��0`=�~lI�m�64�~��������g ?!�ѧ̅9���hn6�&�9��q͒C�:l1�"� �qiX3"�qG���@7�㚊�	 X��H��y1-��ᑄFR�;��}�F� �-m�Yq,<�`k"���yZ��U����y�3@d�b�B�8��������[�V��*c=k�B��cF���ݥe:?���+W|GNt�FoI�V�����I�:~��9�H�L%`�1��lRe�fR R�c�{�e�Zndu�w,���<�1��"��ʚ���֤rȚ�ą�'LL��p�u�j���|��F9���3Z��^��Nk+�uȀL�y�.��x�8A��a�4Or��f�3�gҿ5�E�$F����O�ك�х$�.Zy�eq[�����	�c.o�e��H΅�u��Q��6�~=���r��(�Z¯�1V��X��p46gM58ޘ��`�sJ��i����0t��~��껹��x�L?L��d�"lM7dQ9���AH~���I�`�R�P�D����v����צE�&�w��;�hp��M��X���G��`��3_�gs�.U&Ǟ�(^�^�	`��ڳ[���-����<�Bd�Ep���K�xkJNb�XR	�MHV��+3'c��L�H��9�h5�'0� ��X�,�.w0d-f�d/���_$��x�s��
�{(8B�ӑQa����Z;g��1��$��H�B�H���� �$Ȇ�7��jJ  v3���N �Ҽ����~�1u��`�t������}��W ��Ⱦ-?.P������N��*�l��^��� ������F�w:�j3|z��|��50���,ݏ�>��0��4�|tW��?�tSx.�68�����S!:�07˷�9I��l�G!�wH��~�'	�%�c���G�A�x4��o���s�E|g8�؄vo�1pww��| � �`�\_3�L��H��������B� �����ha���e��_��g*��z!A�b:!`��F1D��k<#�DW	��-�p��U��f�L���h�]���� +8����֞�f@d��K�^Pp�	��X�i%�R�`�԰A��	�{yO$'�gHBF��HV�f( 0�6��C�
?�9�v����~
ih��sVm�t���ϻ�u/�z��.��u+J�g �C�#eK�@�h��|�s��a�4�t_�X� �*��Uxr�W88�H��(��<����3�bZ	�kv�@��H.aPY~�A�k�;m�����M���c�k����k��q�ŀe���X��,#FG��aP��(xq2��3���t�&(L� ���]k��~1��<��+v��Y�|O��
Ҁ�l�w��R��֛D|��8��ޔ(WRm\?+� �F�49eQ�uM*+aXw0 ���ia)�����u��5���u��䎺��ӎ\d�i���6�n�3��S�C-hQ���g����Ok�o�<�u�߮��T+HVh�P������ h0�BZ6ؓ\��CN�$����U�� �b��ȠKX�t�,��F�'`j�u����Ŋ�c��k�v}����g��_M�UG��|��0�4�ZΙ,���,�\�2�d~�o-6�2��֞�4�n������!Pc��<_�1�������HA6��д����',��R4 �bs�  ��IDATC1<��rQN&�*���@��m��|�1I>܋���X��~CZ���C�{���̏��A�,�]eT� ��t�����?o�[���܆�Q��ڡ�.//h{�SAR� 91�@k����i���i1[��V�/ ���k��ÛThqoO��GAB��3`o�����_˝�mɤ�B����u{sKA60�N�}���gmE �c��5�����H�E�P�ww�k�G�~��Ԑ��8�0����=ei��qL���t]9㄀�N�S���Eh� ���D��G��1�] �t�0}s�n����3Yú��7�w�B��h�E.��AY�E�-�25X���X�y��)Hf�p"H�z�Zs���Z>:l�$��<U�}��c�Ƌ��<�Nf"��v���3���S��D�b�%F�Ϸ���V��W�4 ��_U����q?&2�M�ƬG$�[
�k@��Zc,�v����Hɂ��Y�Fq1 ���Ü��1�=i�M"����k.1���mY$}_�|�*eHGr�z������FQ��G�,P�I�r���� 2�K�%��]}�,����d����D&_^�G�U���uŜ����,	��4�L�H���a�G����a`��&~I�u��;l�F�0]����d�qb=�ۛKZpP���Bp\Y΋���j�|3g�����[k�)-Nn���ղ.޾ł�<�c��©��?��C���O`����9<8 fc.��4'Y.x���� ��tT1��Ju�"+9l�snfX�	���Pg�/��.� v �cq
V'X�`��"�&2��� I+a�.�[9}/+1�b5�*��м�u���n�imM����	da�q��2�n��r�OD �͘�7�
&¿��ا��ɻw�HT zƝn'd�oK �.��h�`@h�R  �h0����g�$ 1�l�-*�L�a0�Yd�.�,)���8�����`�D4@��o���>�~���\T/z� ׭\HMp�OS�� �>9yo>~�H�21S�N�L�=Pz�1��s!�{b�wxmlY�cN�b�����8����ߚU�q��=P�����u �X�>���X�n���?Ҹ���8���`2�gl��Τ�7�*��s��n�i��߂2�T��DȊ@��x������6���,k1T��N�q.a	��z����Px��w,��Q��f�B�E&,d���>�D�*"`LZ�0�<�Ld<��㙤 4����9f)B�A'����@TߗC�"�'�2G�y(�i��/{r��1nT�!>��?�=�z �u�5�CUV��Y�r]ζ�O������p_i�9����s�@�K	�Ș�)L�U���L����g2.��/e��@T�E�)�B�Z��S�T��9� �W���`����j�{ko�^X��'{�,u�X�����2��usrVUO
N.��w��v�'�p��QqOd<����mtq��K����v�O혀�i�L����i�y���Y)\����j�$�n�6Qz�0�����:�V�~��=�ξ�����9�4û-2��<a}.=�Mk���=��گa����1wdC��fi(-5�kO�������^��v�_p�>:"��;b r�7�� I4p��^�G��,I4[pO�LD�� D��2����{�X��7feu��5��{�@�ͦ�W��Y[V+Yc�I5�i�2���vmW^+[	DH%$�ER}z�Tf  n��%m��l���ʌ;��?� \^����hPv�<�i�V&)�xv4�� B���dfV�����'���P0zG>��wČ	���[ƹ��|�� Ƭ��R�>a�<3�*�Lk9�S����1�Yf3��q��f!��-��*O3!0T������͟��'�T���+����� V"�A�j���=l.�GY�����C�X�`��(7�bّ�"�Ƞ@E�O
�lV2��=KV�����C�O*�}O��;�б�`X��|$��Q�G��Q�������0L���Ĥ�~����J@�
hQ67J>z���G齔�����lV
��Jk�Z.ćg�^�30�{�-z��|�L��®�!�ls|rlNޝPaQ�_])���;-�K5v&e@��:����1�a��R���
��!5^��h]��*�s�?�q��sww��w�}��"á�
���i�B"f����;��qs6HL���N(�-���[��,q7K!1먞�¡+�����@�)�8=��02~\�=�8H���L��v�G�ِ��C�anv3s���iV˚գ�yf��ܙ%!�*餵�d/
,��?�����6"`��S�����m���D�y���e[������a��0{���;~2�Θ;��+OP(�P�Q�j�4]`��k�A�<IO]'t�)M�~a5����y�҄�YI,k�6!�r8���p��PY�/���'��8PAط�o�{����ԱC�7ʨk�����s�Bf�j;j�3sZd�@������lM�cf����0K��.�|Rq�8բ9 \gA.�j�% &0��)E���8�d4�l'�/̆��t����'g��q�-��89y���)��T��$8l� /#J�5Ε�P�E��M��yX�F�E�9�Qk��V�>�~I�3�f*���!
 ��S�;TE�S��a,��� S1��+��0N����z��F0@���T�@`�?�j�0��6y�'R�}�d6�����+q���6�3�����h߁��hO,{Å�� _ 7`���,q�au��c���Z(oso��T��g��c���� js]+�����y��,�)н�5��-Ƣݽ]
���>~p�2��`�����ڒԄ��b`�%� NS@˷�����\���;Rdo�ߋm�q�1�C���gA�!Ҙyj���h�a��������6(�9���� �� �����.�T"���̋rl���$�Ҍ�����x�%U}F�
��D�J��������, �����E>��	��M������(S���=:8��u��Ț����������� ��gا�=��D!�K��d��h-��[0��o){cקO����PQT���f��!��q//��=���������s�S�g+F(�1�2��z��d��\$pbv�d"��h6�&j���
S�MY�V|�pNbT[ ���'u�ZL���3�M�L���SX�w��`!z�;�����"H�w�Ƿ\h�df�*<罍��y?�v!��^�3�Ӑ'�XT!Pm��N��ȥ\�ቓ�l0��[;�Qbt9
�Ή�r�Ȋ�0���jp֑J
'̸\"Q�@�;R�
Ec���*�vL����ơj�,�[Ԏ9o��w�'�G3�����Z�,x��Dde`�$\��H?���:k��I'�ȮhaF��'�h��Ei֡ŗV��L��������6{�{t�+������1� M�Cڶ��6� ��t!��*��1{I���~'����3�+�3Ќ6 ��5�� Q�_�� �!�ǘ����&�sВ��J�b� b��j�����̠�l���ߡ"V���1
 ���y��R��t�a���l���B?������q � �H�u�SĮ��������d�ݐ��@&}�Mb����R��� 3_A;���O��j �A+�H�.�e`J����#�����;����?2�Qd<��r��{�# ˎ�4��!� @`;~(��`r����S����4zG�1��Z龹���{ �#��d(8p�	��s�Z��P`���>�h�M-ً�~��0��,�6�����^��I��斮����{9v邑@yo�T[6�Dّ�f4�F{����{��Ξݷ;{ve)�I�7ٮ������Ed��\� ��F�Յ.�M��_�5NMN�D >��2�e��\�M�����l�Dc�l4�)�v���I��XU�����	f/s��.���f��e�~��ݘ��)��a\(�����Ƹ���i[@�?��e,�{!�_G�S��U���9�0w�������h���PBT(OR���AB����#t���[��f�#ֆ{.*�{�O ��>&:a�L)��rN��9cgY��ݞp�4�SVԯ�A�VK��7T"C�J�v��Ⱦ���a��]n�dm�s�X�P����'xq)@��=f�1��&@�����A�9�dMf�� E�ф��-�D1�e �E���TW9�D���~��V��Ҥ5�@XeIX,�^�ݦ�>��������1_����?s�!	���xe+U��f9�p�<��"�S���ޯ���U����eʇ�S|:�7Ϙ}��P��%2�A��8|V��0��`�����}fiA�$b��"���n��ŏ�X��y Y�;?7ǋ��}aS���vT�5kx��,(Mu���-iJ���Z~�L�ùV�4������Trab�̔0��d���)��u�r3�N�Æ*3�R�7e��8@_��`�؀f.>CF�C���YM9��h0�%&����|�U�°�pS���k����}�	��)ߋ��$"�1 ,ed
@�UD�YV��$�%Ƴ�|��(*�z� J��o��a��*�O��m-Z��az ��[���1����)��F�ޚ�����D�ǌ܃
s ���)E�̓�������F������k���t�m�^�z���2���
3���2?;a,kB|���{��,�� �y��0�F!��03L�en#e_x&��{��x`=�-@�]SШ���,f#��خ�#{3L�f��P�;e6��*��e�&d-���Ο�����1ݺu;H�� �`m��8�l�`v/���9`\�� 1�0������&���K���@u�)}C3`�c���ݻ�� ����I�:َIZX��Z��(�����/TV��9��]-�K1�%�y>�Q�dH�g�<��:y�\ 03���U�l��=cY���_hxK� o�i���(�i.�R� s�Ņvk5�{X�"E<�i\�3�^���g��^I)��5y"�n#���X>��.�b:�<�ml�@��4�)ɂ�N�5%�Ԗ�aj��R�]��}������1���T!X2 ��&��ZMҁ��tgD�u�Ε��ҩ��;�=HJ���B.e���;(e(.�T����@�F*�����Z��ʢ	�N��1�\��g�x ����QtM�Dgf���@��)Q+��0�S�Y��P8n<���G�$�����Bы7ur'
��9��?���1���-z�h�z�KF��F��ݜ���:z���8�*��C�Y�C�5��4Eŧz�[ ��:@hjf��fg�;2F[
L4�&�3�����Q�-.����2V���9�;���,�΄U%Z�X$...���iK��Z,H�+R2x��"�Se7D�t��8���6��(��ӄN�k�d~����,G�Ζ1�NS�����TY�rS�\�bk�=���Q����'�����&��HdT=�ugw�efg�P4���ۥ�W�n��ls�"�����k������ñ&J!�yAl�7��|��'�7��� jpn��  �j��9`��M�g���&ʫ��*��8�}�6��� �B�ŗ�S�H�����|�E�p=@Y��6xL+3�&��6,r���"�!�#�6��!��2+;[��K^.D�%�[����,�]�Ku ͧ�*�JY� ��r�����eP��ٝ;���~3���3�5��1��$2�H�Es�I���^�ٰ���+z&,O35��X�8�{t�Lb�4���;�q���&���g Y�G�HƘw�DO�A�}���J����d��OP�A3�4إE�t���Z$$X�v=3=�ׁ���n���=`��j5+l���:���ş}��HPY��Ұ�h�o|�oˆ.܄:P�����Q;	�>a#�ͷ]tٍ�]�>xY���A�+�&�[q)*Y��(`.K���J}Mo$[?���>�>cE������eM"@vV`4>��w}��F�;�� ��A�د���H��P�j<c��4`k�F^>v��c2�j(. �8�1J�e���L\7A��̧>�Wo��ȶ����c��"ʜ�R����!k:����EFbJXbpJqXL��4�r q!�n�G�Q�D��]�o���N5 �=k�d�:jX�����S�<.֗]�D�M�zg� �5\f�jf����pE��9��
L�
5�ܹ9v1���A�(�sFÙ:�Wl.,J�v�㠥0����Ɗ���'�ݱgg��R; �Z��Ð� Hc}&	�h1���1� ���ٙ�)#�6�"��3T��*3Qr��te�fg%hW=�⩦��:���x`�$Ek�BM}R� �Z����X�(J��o�cb��m�uP=s4���`d1xr�p��oo7��k.�����0e��}��%�I4J���w�M��1P�2͆/Ng��.��ו��%'Xw�΅4�g��\_���2p����^�|I��|�������.����S��ۘ�A .�9k�����?|d�/��� t!e��R楐���X�k�rQ?w?�F�Υ aIR�� פ@�JL�� �i�Vxq�K�
�����0���`Z����gm���*w���� �ƽ�2�Q���dHQh��o�"ല�����,���*�����R�e\�ߺ?�8@v�ކ� ��M��x� ��߿ρ;�� H��c{�jA�D��? C_�IVJ�n�7��x-�h�9�a@�8<��p��rq�B[.{;���o����ȹ��iZz8F�٘9pYd��}1kٟ��Y����#=�0q�:m�r[iX�q���a�7�U|�Mٷ?C��*oX�8;���k�V�=���l��� ,��z��S�e��jg	�����Mc/�i]���!ș}���I�����V�v�(z��-��}i��V?�AP	�����f%�a���B�嘜���q�9�&��)dP��k��Z%�즙�~�v�R���}t�֯"3��*L~z�0�m� ��J��H=8����p�t�1�&�E�t2tR��{8����H��Nv�J�{�QgV�ĝC��N�l�nW�6��7�E�Z��Yu(y-)����yv��sMr�g>%�h1o���D��K�Fva��I��|2\K�6��w�%�}��{\�.�_�9��S冴�����. �(��'���h��RY���[��)��D�LZT0���iz���b ����u��N_�SجO�k��Z�g���X$}0���,3׉E(4hy��fl(���G��Y��q��D�QF)� �Q�`�}Y:�D:�䝎x���(�c�Iq�&�l�0�;1�A�c���b�!@��%��u?`ZT�V1
ݩ�gH���-�Y��1�k�>��w@�xvf�؟s}�p���P�/l�ŋTz]bP�_�!���絵��E���	w<N���q(��t������%�cg����AY � ~�t�?�{�c$d=�qg=���n&)�$�N,�?67�D��=;d~�0�sL�\S�,80 Ci~����&*�{	��<����4gI!��n߾Ś�hs OA
�׻����U�������0�E����G���1& �<������1g[T�KdXh5���2���%��͵c�P��0�)��<��su��u�j�C�+����E�c��ϔs|ӈ��s��Ã���O{{��5!� `�����*#;�)W�*��]0&i�
����q����k����J�%u��y������K^�o|����5�	���`Zh��n)t�?wU��#�T�P`9_�B������P�`�&^X+��ʯ=B=@;�����K�3�RF���H��b�����`[��;$%��J�-�3��N�C�
},��>�f�NB��)�e^�LL�����D��[tL����S�UgFG���ڔ�i��]�W�;��Œ�x!C.�-6��lCK
v�|���G��ʹ��$Y�`7ڇ��z���,���wϊ!}����F�1A_T*���>�|D��JS�)��0���C�lI������9Ʋ��Y��n��9���PY�I�ݜ-m�7���qqM�8��;\����`�> ��0�6�2��l���<�D������=�i(h����<���1X+�6
^D߷ٞ� L��`�ܬ��ġ0�+e�� x�Ķ��>�o��K!��C��X����\���-�B�b�Zu��1qJ�ج���qMae�L�}���	F2p!M��̠-�e�8wHf ����}�L�������)� � "omm� ��geXtrQSw�xN(4��yf������sls���MX.�W��s��,3�د�5'>������s"sm�5d��U��'�biZl�p#�QP��R�4+����8�C��3D�ٳ�TVI�2#���t�56�B�i�o�x#�Ϲ� �� �C��`�V�_��j�x���Z��QEM��>κ��B�X5��c��v���3��9k!��2��Nc���ڬ7j��)�1���xi6���lʹ�־�}��n���~���@;�r��w�@(�I22��^���gb`Yk*�t:��r�Ҏ���E���gև`��˹T1�D*��f�X)�0�L��E�dUπ�V��*Տ�}�O-N �͉�/�y���>z�-쭦
)� 	����R�9��9�6�j]&�:�����!�n��o^� �KRhD#D�gs:�[������Z��w�������	:v�<&��u6�v�hi�P�����Z0�������.<�h���E���MJ�H��=�A�Jh��;��g� �bi�iKt_9E>�s
) �3� =�(���k	�^G0��� �B�HƎ��B�:mÞEX�`c���������4�ٹY�*&s�(8`L�ݕ�`)s�lA�:����l��/jt����vpYAn���7R�r�zNG�[�=�^����/��M&���bd�Lk��sŀ&�Ϧ��\�R�Ef��ku�KZ�/�s��y%mx�"j�ѿ�� 	&��Q���ע��|�>3-��-�����}2�� �}��%F�TE�,� ��x�2������~�---/��O+o)C���" �g�1��u����\h�t��̣-�X��f���R^�a��;le�e7Ȟ�)�LI��T��y��a8?�3���;�:�r���fA�p׊{)���R�pf���\�1WC�~�$�X������f����q����
����|ߤ�iDe�R- ���,G�FN�~U+;�R&�id7մ�)�S�AV�~gg�� h�x0��<�|�^�}�i�����t��G׶��l��K�r�ׄ��?�d���*K6�|_3�J��7��^�
\6���,,`.|�g���	�����.t]�O��3X�c�GoC���-�����`,�x���a�
�k
V&)�e��S�f	##��x�t�0`لŧT����@N�Q��T����k㏣�u1/z$�K֢tN,���)�Tqo����6�bqQ�"+��,�[B�"M���D˓��03�a���^H|��74�0� �]�`Zt��I8?�ѩ9��Z3Q��`Hc�R��W�<��e�N�Մ�M`�2>4���K�S3�ڊ�ew��i�l�33G��L�60��ʽ[h�<;("
e
Z�I *�_m���\���$ǡ���1���,K��؍Q(���6)�T���9�.;�zy1Ȁ0��̤CA�b�����+��P��T�k�1jÉ�&�W\��Q�������~5��d1c9��H)�|��T%�5R�lgw�666BJ;���/���������������4��F����"#,�u�6�]�A�"�2;,�$C
�*��؅��Z;����p	���J4p��|�����g`�>|�������,s���^��@��렩�����X�a(�`7 JmD�!.��r8���Қ�	��������Rk����O~�2��@�-{�WcN3���҃����EA�ܧ����p� aa 푞_.I�B�^]]�Ru��`�3�ӽ�����`�0]�z�ڨ-gE: �au�28L�5�Ǿqoq� p�_�g�����0�*k}�iS�������z�e����^�tm�����*#�I����ن��	�Cm��� k��D��'��B�:>~�s~�oz`$�h��`u��V�'ɯ�d�@��|@��L����ͳ�Yo�	��}lB���{O��ak�94#O�{��o�(��b�:�/�lń���(.�<qT>�R���Yݱh�i[���ʹ�g,�}�,��wP��홸CR�"�uK��)wz�������:1gN�_�{u�6�A�m8��Z�vwX����F��G��}�u���a�j�&/�*��NMN;gw�#�p�QPf�ObR��2sz�ip��۹�hѡ�}�Z��UN+���F2��,U|=�ˉc��� �l���춁]Ҿ�f]��
�.og������ �1�˧�z�Qh�
t
v�΅�Yo3��6����ѻ��pC���W��Dk^S����2�� �b>e?��ÃrA�ōe�H@u��9�p�	x��y�M�Qf~��Yh7�������k�,��q��]�eپH�V�X���Xƛ=�	���x ׵���u�M�5]q�`Y���s��7{��#��f"��p�B���#2SҶX�D}�mo��@��V�Q(�Na�j��4�+�A{4���qc��e.�癩��R0���* `l�	�M|@�(Z�}�������Ě�RCC����5�qu4ħ,33Y�����؃�3\ O���>5̈�$�9�����YC���y�$ ��`����¦���K���fV/�{5;�$�6�����[�Z����G�@<p���{B�pnhS z4Yj��f��l�1�0��3�EMEs�|��5L�"��ӌko��}��	��+����]�!�� ���@�J�:h/<�dJ,u:?�Oў��t�\Ne�Yt���	�1�����<�=x��r�}b&f̜>�]5�s�ի���|�������ok��N8����K��A0�؇־���~`�L%W��k�~-�޶ 7'})�!�#�H`���l;�H�fr�q7'N@e�b������}������OE��r�H��L��~�/�+eY� ճz\���C��<���m��ء�WU�~������vn��4%�*�Н�5�s��\��[�K�(�h�n���3uN|�v�v9����o髯��/>��6^��~�����=ZXr��
�����-��T�i����� nl�t:��a[��@L괥*x���i9_���h4�e�q�S����Ee���k��?yN�=��x�b��j��a�d��]��lʥ��u��K ]���e�b�д$����~�9��׹BW�(ʇTk�hk{�����zB�c�"��/���(�:;F;�� n�Y.����%��ekH9����R#A!�FO�&$�t
Tmo�0+���5//-�~-k�F�ʌAH}���^_��^sk���UG��h�( � ���\ �U�⤸��'>S��AHbL�/xc�y#�r�|���b�@�$�C��������~.����²HA��|,[��D��eH��`fh�E��??(��Ɛ31�G���
�EA:-�ڪR��� ��8�}g̴ۿ��l^r�Q�f �8��f��_f-�	��]��F�6��m��*;ѡ�p@��9>G�r�s��p���|.岴!���2­��LN�93����f��<Ơ������ʑ�S��&g�B��R����l�o�¸�w��2O�_ضr�<�$9y>, `�\kZYL�@"ix�xi��giiq9���s:?��߫A�đ��rm�ny�p���xr�I�g���~R3a[�Q/s	}�_Oۍ�!#��B���$�_��:��~�T���)BO�P(#�mQ�T���q+3#ZzǇU��������Z�M;������2(�"��<Ҍg�X;��������֓'���@�`��B-�^����[��xGG���I�}�����+���o8����G�f����8U.��p'HE5R9��4rh2���M�}�	a,�pY���񭩡]vx��O������k����p�k� �¸b�,��k'9�K���9V�Y[pl��]�F� �<C+�L�F90��t�	 ����6?����q)�-�
�J,"��R�!{�S��~�g��٫贌��Q�6�O�h�T��&��1/g1������k/��2+�����|�`)j�x�|F[�t��\��<��f)Sh��	i1L��ߓ���iߑ/ؓ���t��� ct:���uҍ��)1�\����_XO���0��Ż7�v�_�󾳯*�I|.X���8��N�3�K��SLD�YR^�D�o�f�qz=~�T�ml��:�u9�W���tϧ�o/���ѳ5�Wp-��mG�i�=!@����L�T75�nmnq�Eu�UwYWI���F>f���ia�~whrc��P�"�$ֳ��_�L���5֞o��:�U՛[�I�YWHS#���e>���gdn���6���m9��yڐ�0���"O}*~^f�цÌ�:W�.��@�m����t�(|����掔/|v�GH9��L���]�_���b0y�9;���/�ku��f�S2���>��ޢǏ�?����ѣG�ijz� �g�Y6>%�嘄�R�����ߥ�Oߥ��?�;}������u6�J��M�hjr��f�x#Z���)b3G(�9��Oݬ�Zߧߤ΃���{����jx�����z�2@e T�4z���-ڤ�}��z}���{7�"�	i��p��hp�S0�$ٍU�֐>U���QhJ�h����� ���g��_�s����q?��2O�Uw0�X�47��M����NQ6aE��ݵA[׆1�*� M0?�����/���1v�ld]�p�zb�2��2vO,eL��y�	��x� ���q�7���p,�3��əᭋ�0S���sN[�rM��+����Go���1w�x�ͮ�8�>�fOU*E
�e�"���&ِ��N�h4��A��ddEہ����;���V�V���-D���
�b~Y͙^G=��ߠE��~}<d=K"���Ldl���ӑ��h��F�N������}�8�x����1܍Ơ`�>�I�)鐴��y50����_L�a�N��A��y[��kEgv�����59\��܀��]�1�A�ݣ���(��٧�!(�3ݹ�=yX6�o�5&���2c�����[DN��A�e�~�TƆ;[(~�I��h{�A��G��1mn����f�J�|�.�������_�g?�1=~t��禜#2��Dp�z[:���3`�%�r(�Q��M�ڽ������^w�Ν_�D[/k4n��{w��]��I����m��hۜ�x��y���V˭Pa[���7�?���aq����Ϡ��s��<��фkE&�k,����pw'0	�@�{o�}��t�d��prP�^��om�]O�愈�Ë�
X�e� {���j���0)7�D[�N�3x"�H���3	c$`^�zE\�oz����J$���(ڋ���ݗ��c�}����V+ŧi�ɩ[0����&3�0�h4#QP���8��;J\p-)��X��m�MF�a�x/Ժ=�E�����$�c��(��b�?Ek���l����//���^������"qL㌓.�b�<Y/����^f|l��9�� Xg!]`yfz�3NS΂j�w��{F�&��.r�W�<�L\�2Xq��c����f�Ai���Y�íFVlg6�����[��`�N���{��B|R
�?�4��[BI1qAmC:�i�D�xj���eX�Ϳ�洑��]�F�o�M���z��dXo(���ԩ@r���[ܧ��B��j�f�����iI�T�&)�����M�R>��W5�z�M�U��t�u[&c��p������_������y�!--t���|V���)
��x�ɓA���/X
ckk�A���w.�s�n.���-z�h���x��:�eEH|�:��54� s���w\%BR���h�E�{�=v�Mu��>-L��C�W)<xI�)�r���)�j��!`�h�_`�,���ݏs?�x�,bq(���m
^)����;�B:��AX{��k;�3�%�D��6� ���!-�:<�1Z�XD����	Z�w���b,A�u?U�``�u��N����,�(ؗ�q�0.c����u��٦͍M���6ЋD^ZZ��k����}=M#��B��	��7��E����R[�4dp�5���t��-����{V*���q����YX�y��y��ǭ�]KkkK�$#3Ҁ����F�3z��E��^��� ���
�-�H2��g�=����Q�#��ܫ��㤍~K�V�vwwy-��������ٷoߖb�m�GL�!��.�(�|dgd6�=�m��>�>V��K��.�{��4�)�������2�{�7��S9��{Gs+�;��]�]\�>��a�Av1$���VQ�U�-������N=����䨛ùFĺRNX�𫗯Y���^�qq�V+��qDuK4=9M?�я������?�Ǐלc2� ��z��DOd��8>K y�=R��$E:�g�;��w����^2�033G{���2��hnz��n�����M�OJ�< �����H��=�6�.b~�3@�(p*��@�z#����:�B.|�z��FW�[�e֘�n���ٱ��/fRjq6.�3�NM��e�s𞉶)�~/I�#�d��RyP��v}X+(����i�M^�ժ� ��q��,�Fb|��*�UL�^��(((T���H	E�p׍��ˌ[hAW��߷�68U&�n7��Ui�?2CqvfL�/�O7$^W�勗.���{��@;���5�WF��f��և���nf?��k���r�;(w
k�UC.鴽��Җ�>�!:�Zd��߸�c_��E�$��{^O��އ��{�����i��7d8����2�N2���/ƞͭ-���Wi�R�WA���
�Y�X�%A�s��$���k�w�C�jN��)��-=2�重�x��66%�	���Vdpݿw����5���������P�dmEޏ��~�U�D[6y�]¼�A+��|��0�W��vBVq�O+�r����J6���)�c��w��~��������`֋\U�e��'�����⯑�h���lO��@T�ϧ�tu���!��r,e�M��O�5	eӥ&P{ �F�2���4�0�S�S���Tb�\ƦX�Ù X[;6�����6���ئ��^�j�=xD?��G��_����]�zm�vw�T)5hfΉT���J� ORD��7��i|b�������Ky����L��/�՗O���;�ƛq���n,�����>��Sz��ΠLj�hea��wT����gcϞ:}�z����KE�3�ִ�V �?~k��cd!��^��֐�L���cE�F����|;�_�MQ��{l��+4��O ��C�,�U����ا��E��w���,뻕<�W�6I�#u���L{��t�6�4m��H&��Q��(�6z�m -�D�/����Um����R��=�l��n %��^�µ9 Y�xY�6�O��?���*���k7����=N�8mh]���\(����KŶ��l������;�z]��G,ѯ�`�tFh+k����7�L���
3�'&'i�`��|�T��G�7������?���������w�^�8iud�p��xٸ��"�$�����DŽ*�c��_�?��{NVol�La<�s��A���V~y����`�R�`��]?�6�	�B֎�L^7�>~􈥢���{�Z>t� �n���ݵ�\�W�.er���'E�l{�(W�y@�ʿ��6�� r����q�	�f���_�zc���������������*_+־-�ˌ{9qinVc?_�/v��\����uZ��E�E?�T��<7������2t��i8��i����3��
*X���x���Dj�N|��W�>`������\�r�f����v� �a�J~��S�^L�e�T iHo��q��-�W�w��ڈ+~���-�[er������![�J�k���v~�m�3e��:M��� �zP^8ۯ�n�c�T
�-�>3[xo��M�Ǵ�w�NE+��	{�M�K�V����3����/�8?�lO�֩z|较"	����8^�;*Ҏp@�3O(N�A߄�΄52���;��_?�����u@g&�������G41�r�=��)���/��O7��?�=x�D+S�����i�J���ޘ�P�]���6|}?����Ԫ��O�9P�G?	mLf�T�m��S�Q����4
���2 LZ�$�b�C�z�;��g��p+�<�.�6�dz�R�-a��\J�J
<�Mh~@�MB]�ùoyP"�F?����k�T�]����S��8���N�v+�,�Lb$�wѮZ^�b|l�e"8U��`	��67�,Ѣ�|zf60)y��q��W�=C�_G��U���r�<�s���6�Wݢ�ʅ�����F�5��+�˴vo�5��30���"3�is��uvw�[k�����ݨ�qX����	4���A����ډ�ɦm�	�Y;��~�2�b-�����ejF�_�^x9%�{v�Ɣ7��%k�Z��Z4O
�����jm��m���5 �V̵R��B�R�3��'2�9 %8І�0��tF�u��3�b��τ�ֻ1 vt|L;;;�.�9_ۢ��qjz�VVVX
YO%H빝����Ps�cΉ���uY�r��w���]�����Y=���9��Z�9�l�u�����ΐ������C���� �}���$죿s��b�v���l�1]ƪ�5�^砖��3[���o�ܾ�����8�l��m���.T
������1���������↓_���;E����3� �a�����O;�����OGG�\h�\��a���&g�>�������o��~��6? 8�p���C��[���v<Z-�}��o�k�i��V'^ 7>��3�� �1>>A�>�_���7��M��x������菿�Oz����?x���yB�ߙd�a�`���`C�>w���3�E�n��Z{�[N@�1Ӊ���lŮ�a�v5G�˵S8;ڝ�p�o�].�ibf���Пj�*����"�P��u��}jr�&��Xwbb��I�?�,��:P�軍�⢨sb����y� �e������������$�M^ ��`���c����-������1��ޢťEf���k�Za\L��a�T��-} d��j�����}������ gK�1��ÇXƶ6b1	��c0��Ȯ�������\[|��1�
ʚ��g F��LG��F�9���C^	@�D��ldn\��K&�̟Y\\`���&���Η��������r�������������.�ي!蜁�I0�2f[�X�R�jg�5��|ԏ�f)ŗ/_���Q��֭[�3;3#�U���nI2�_w��lÙLg7�^�Yz�d.r��tf�cv�g��&Q�� U⾧k��gTHJy�a3'��!��8INCW.Z��a~L�⼙v�2s�|g3�b;x�1J:P{�!�yr���.�TϠ;
��?����L)�2�hgs���t�ߠ����1�$���I���H�>���a��?��������j�4^)����{o��L�to8"u��[1Ts�Ez伂
%�>�fZ�Ãm��˿�G}H�떦��л�C���/��뜀i*W��w�t��=z0G��_~�>K��Ͽ�gO��a퐦槨�d��I��W�N�<:R�]`:���#2![�c�Q��s������(�#�D��l�W~M��T��)� ��C@�ݝz��KT��C4}�1~�ǥ
$h��H�'W���8����"�D�24:�8�'�_�k�C���+�d�Xuf����BI����/���2�j����� ^��k,��Ϟ1s,�Vj9�m��F�v�����l�������D��0���V�s��ŋWttx��Ly���;1.,��o=���Y7�4 m�vՠ��7{-4.J��M1���B��b9�5��������ZQzg�gz�u{e�q3��=��3�N��h�;�>-d�9�I�j=d�ܻ�������x��ӫW�D
�ͻ�o�b����q��x��&�Z�NB�.�#��}<���W�4륻sz�|�/^8_�}���e������[�G��9/��*�mߓ�*�چe7�ː���+���Y�*��e�;"��5�#���K��=19_����R�8�;Zm.$��6��� S�|(ȝ���%F��.���w��mT�damL~����4���ރ�iLn�Op����=��[�����!��E{�9	Ğ��@�L<�_��W�?�:8أ�Ϟ���<�''E��M�6����yN��K�F���H�.�+��\�5�+�=:<����������/�p��<�Z~�>����?x���Y���h������>X���{���=Z��;}��_hk{�*�c4?1A�z��6��BQ�*��1��G�%��;b&��{O�:M�Zv<�K��\ qZ[�S��>-ZC��U�]{��:)2��������\F;E!5���q��j�t��#z��033KSS�49�i��P0�d�a�`�d.g�;�s�ѫ0��C�5�<�;�wܥM���p��k 
���g h�u��g(�D����n!'L�2;Z�g�,Em�9��t�Œ����5g��)��)��,q�B��G� &��1�F�>���޽�@9����~sz�ô���z}�}0��,�����@{�Ct䴻�>[]��)˨=����9�8>�k��#م��
�ꮤ�:�;��WE��}d�B&M�m}V���\�W�n��2`���_ٴs%Ջ��$,9�������Y�𹷷����EF-�ǝ�w8���-��C��>��R�r��N���՞��l-����4�p�'&�S0�J�����ep��F�}ߵ�F�N��l_���������:�d4ȵ�� �'�&��7ͮ������������}������6e�Z�{�a��,�\�Ei85�'?�)����;������_���W�Z�i�XyvXm��̋zvP�&��I"c�bh�f��ܠ��������?���������;�Џ�c���b��lrD�G|@3ӷ�Cs�u�}��������t��m��p���� �qp��}x�AR:[}�ģ+cv4<n���mڻb����sl�6�������&k*�����Ǐߒ�;��S\��.�.�x����ָ���oiue��?�Okkk�ߕ��[I�2��~aե�����mg`�_�us�:Ƞ1����(ve��,n;\����1,�q��4V�%*����1MMN�ӧOiύ��G[�9���=ZX�g6�4�� �K���Y:j\.�����ٔ�j,d�cm��1V����,)'17t��E�[Oޢ'O�v��抣��Y,.�h`���5�z�ǼئV�u�ݜcxG��{�����)2�F6��4�Ƀ)X�q�vy�>��3z���ǘw��ߋ�K,��)d�B�X5��1�ige(i��h��#�,Zp%�dNMOr`^ �!s��?cjr��"�	��]�7����|q���/�&�*j�J��(3�1��Bw;� �NJ|��TF�
�2F�u����Z&#$I^k=y�AЃ&�q}�܅�9��qf'a��)o�]=`��u6E����B�	u����y�N����0҆�����5j6'(�mb�V�n����ivf�v��i~n�~�ӟұ����F�&����l�+!��JK-n5'�0-�c�0���[����O�+}��3����2��翤���=����$
������C���stR�r�����k��[O��	�u�z�w���;-��#�X� ��G��m vV�³�1V�(����.�1�]�Q.8�W�\z������uq���|0�Y�>���pj���)moo1��;w�pq0(�z��E!�XC3�A�:3;�L�Cf?X��}±[�|wn�&9�#�ɳ�č������F��@�>M��zk��`�S�IZ'�X懷H��	ؚp@K4s), H�{��B��jԤ��L�3^5�c�ʔ��$'������d�mھV��~~�۝���X�Lð�>�Y����W��jGGǴ��`�^�����L�p���v㹀�Ȁ+�ÁL��Q�F��hsh��M����%�Θc�.؄<Ӽ;���P�ݦi�I�A��h�q���[X��%&�����%ݸ�`��6�\ѭk�1#�`d#����İ���� ���o;����xnF�ޡ�}[>��6�ۦ����^�!�.�Qu�>�ɴ��kE㥀Q&�ʰ��s>7$��vE�>�!�"�׊h1����c�}k��W|��`��|`מ2���k���.�z��@�g�(1������XL�J�{Pֲ�Se&4"���8��c���+1�a|aZ�:ۥ0��t�|��f�X�]�(bM��lBt�)	�$�8�"�qxx���S5K�bq~����-�/;�I�m��ݻ��x��g����.�%�|c� �5IiHE�z��k�R���]z��)����_�w���vhfz���<�����s֜�2�NU�2 @G��
�W��#���w���i~����S�Yc=-�B�Q��p��T��s��ć@�@�P.J8`Fc��5��`o��l��i���}�kaV����'��D�M�o5��P��w�q��'H���2�i.�=�\Fݷ�N��`Y�2��STZ������g�؁�>pw�G��ڽ������� ���^�k�����v�#͢ћE�l��H#}\�$��r��z���w<p�iH�2� �����D)� ��W�o3����}]`���&%�}�EK���e�r�~��W���@v�F�,Ĥ������B���#�>��.s;���snlwۺ�}A�1�6(r u���~���&��Z���/.(�s�g�Z̖�Q ��߿��K\�_@S�S�EsMƱ�u�¡���΅��GC����b��Z3�j2u�/��P]W#��cL�31�O���P��g�QC�����R�?�w�W�y�76>�U���ɮ}�z�=q�iZ<�X]U�q� ������
b#;�R�C��������(Pt;�ɍ���������a�Ȕ��d^�����.B���d�[D�.UIGʊx�:7{�$2�2�z�[w~���Ks Sֱ���(h�fڵ �c�V�6����{�V]T�A�¯�H8U�����ٹ9��/���7�6����t`0���	�&{�Xa"�� �F4�@��U�����Ͽd	�J2��n�<���5�BʿD��$@��O>�j����\��Lٽ�ˑ���^�xA�n�f�]�r��p��4h,w,V���8g�dg�?b��Ѧ���{�Y�ȳ<{�����+z��9�߇�ӽ�����s�k��=�7�h~���&m0|쏇��o��?{���7 �~���ݵ�ܧ2@
;J����p�`�p��v�isc��( [�{�
�n��{ʌR�+C?*�0-��@8�%�'��K�� ���P�?�}�4'��J�mX0�~CSxfv�)�畨Z�y�y���<of����`�㞠����_���e����=N��Tҡ�r�\��"?s�sF#�V�h3(Ȭ���Y�r����;���}W=g�-x^hߢ�/��8/0��I=;����!�8rG�i�X�,�Mǋ�o����ow�E#�ZV4�i�8��{	sY�Wa��ihue���}���,�	7��a�R��U��j�/��T433��V)k6����v���uz�'p~���|L|9�v2. kQH!b�y���d�:Q��|o��� ��,��Z���w߈F#b�&P� k���eNGAK���h}�r���Y��:�%�����4*�Nm�� �����[���J͊���Y ٛh�XV�g�xm�*�ƞ{[	���^~!�(Q�2���)v��3���3�f�����RҤ�믨^�����A�8�A�����0���$ ���)!��ky������������C���ޢ��e�s)�+�T�T�ݽM�����	�4����33S\�Q��ir��X�s|}����yp�bPÎ
q���~���sjSH[
e_���sx�t��jc
���1gTY�ZtS�����������7�p���=z��p������������
�F�PW��K��W�C ���j�Q�|L(��f[���͆��8��g�-�A0{�w����f�[��{�J�H�^ ��:�d3��X�ltn&5T)�2a�뿗)��;.��;�JMw�&�#�eH�ةu>�ޣ��������U�(ơ];+W2���؆|���G�,ł�8 ��lQ����*Hy�:��2���,�sI��<�>�����4S`*I[�"tlb��(v	�Ņ%>/��7���zv��׌!M#Y����a�i�Äv� �v&���c�7��\��������|���8+I. KI���X�����|��]h�.֑ ����V��ց*+��P�	�[p��g�Y�^j�l'À1@b��k\���~^W�LV��O@ �%��Q%�PX~��Lrq�r���K5�˴���L��|��"�n�)x?�B$��ߙ\����!$p�V }a�u��ԙ�hÚφB�2>�kk�ת�>L{�#^''>["^����F���m���E�y򦼦�����I���e xZ�Tc�k�NGA �ӓ�4=5�U9��cvf'8=wg�*o?a6��+�D�����t�J%qNXM.���H������}��K�WW�hn�ݹ}�VW�hr
i�����t�[p����Ii{{G�3�3�q�ݥ��q7�ݨ`Y����y�$0��I�#.�&$��pL@�:�{��b�owX�zvv��z	fL^�?�,0CE�&?{���_��ݿ��<y� 0�g7����	C�ԓ��-�5�]�������1p|�W��y�`��5j|{�րZ�����p�-8�h�N0�V��4 ��b� ���EI��J�� ہi*�����2߇��]���.��E��x��BJd�As����ܦ>�,�d��"87�:��0�t� ���,idg.w�'�5Z�]A�]�}3����I �2X�I��?�Q�o1]b=��y�z��+�c�z]�+�=���q@`5���~ .㽖/�V<�] +�̋U>�2��c�����9����:2��N�n�6���cƠ����h;7o����%���둍�,�W�	
y2L�$�{)�T�� ����Y�l.��W�X2��� ��p;�`��o!���et���kk�רr��#R/]ߺT�\(�����9�	,e�\o�$/��Լ�Qldٰ��U�i���PW3�:�:[�Zw^
���R�E�,�_k�ED�8&Kzf��Z����,��_��z)2[
u�x}����T���]�]M`�/H:��6 L�dϨ�� ��E�FW1�_K�XS�&9��@1����97yO��x�D�!{��b��Y����꾃�N�Gޣ������ɧ��_>�t)D����X�siy��,3HV\j��..����ߥ�O�rdr++��^c�;n�4��A��'�W+�6$��$m^%A����VEﵽط���@ˇ#�x�Ym��I�v(
R�ܢO?�����{�������o���	 �P6�..)�8y-��ޯ:�¤ }��G4����?�sPy �o+�?e���Կv�m��V��U�C�S��X&��A�L��5n�H��L�p6!���iy�j����.@D!��%�UmB��-sR��*K.fɶ`Ƹ�띞���Q���,Y����wl��y_t��3�s'�v
61����Af7F��4���G�lfȈ`8��bi_HW}>e��|é��4��̘����i�ch%�����1��"q&7ad#�7!>�V�^v%�m3� �i�~�51u_�8h��d�չ���u!�\��S������z���"�k��X�NtƜ.Z���^�Λ-��RX��ډ1!+	|��`N/.,rMdU)y!e�,�S���h�q�	�C����=�������J��t���C��_�g $%_���uwq��z=�b�fU��r&�q>�f2���]���� �{�L�&X�p�m���ݩn���<`��Ä�p ��� �&J8Ҧ$�l�VG0M�VƧ<ِ��h68��Jb�V�?R�M�����n��E?42��h�Nk��tr8 � ���ɩ1w�}��'��?��>��g�d@OLE�r��-҂s0P��n���I����J�R���(�}-�9�0��2�0A�k������Wtke�o�8���ã���"�� !��h{�-�=߶;}�
��G+��v�O��S�ٵ�g20�&��b&���Y�z�#rI[�`�COyks�'�����ڥ�����)w�b~p1)Nl��.�����@a? rp���&�E_V���H'����lW�N�R�'t�6_���K�6�jF�Pb����+��B��"�X��#�$�"I��kX�>=�+wc!]g8�V��P�
?�ăԞ����i@��|�(
�H]���������<�U�������O���plO`*g�el궡m�s͞?��F.���h�bZb�����7�z���!���%�>�>�x(�7^���2�$c�	>��PN�␉/$���$Py����e#;W˯�:�ɾ��hRg����i��K��aV�f��F6��o��8�ή�뛀�b̞0��g�������<���63$��y��9H_��Dd�Q��浾n|���e����rc0������� �w^w��LTo�Z�Y���2@v�F��<!S���L��i<��ew�F��ʟ�Ke�6��h��jߐy�r��9���gJLG�L6L���ڢN��j�BF���h��WV��n�]"cYAeCJ�o��=/�5��≬r���<�i$�tB�aH6����8�H
%4��LY}lLR��:��	5�nR/����� �3��R�e�Lt2��%U�����G�����o7Y��@h:OO-���-����hk{�_?xp��{�}�<���K����ą� 7 Ʋ�Q)�qO�Ȕ&haq����ңǏh��kq�-̳܇�g"�0��r����e����c�Y-
�]$�l�ˁ��o{�Β
�_M�� �H
�<��	/^<s�Ʃ���.;�,C>��ܭQ؞�h���a'���N�����7$	�������\�/��f݄��q��r��n�M�5����� ���+�2�Lv�rQO��Q1Z��u���9(-ݔFֿ����FNO��
�?e���0&���DB��Gu����S�7�����ͦgN�|BV,�!��H��o����\K��M[P'���B���|�ky������h�i�!�5�d����$�1ٛ2��Aw��K �>�� xƸ︟<�5��3�_K�����:?�4����MB7yJ$^��:���y��П�E��dI�Jp���ٻ�*&3��u��.e�wWodp�_قON�)�e\o�B|d#Ywӥ������)�q&���KB0����9��F�|��=�Z�,�>��`��3�+9b1�Ǆ����D�o�`6
��\(���'MO6��@�H�Qq�W�.��M�o�Gַ&�x�ҜO�k~�6翑�A�@Ne��#i�\m�F�b-ҭ��������
z�*�hCP�He#�>ܿ�V�2�w㹋�Q���v5�0�,(l�T�� BE/��rŋN:�U�5��)ǗN����Ѩҝ�K��0�@�����6^�N3R��z�PXX�ͭ���O�H���Xw����>b}�δ��Xp X�7��� x���B[[��_?v�;��������c������Ӷ�ŵ��PH�����w.����v"$0��1�n���A��̉Lg)��mz��΅ˠ�z���+�����ga�V�N�I��OLML��8�!�[�����f9�3������;D'?y��F�>"=��V`$'�\�,�b+4r�]or�
 0
��������?,Z����ge�c<(ymꦗ����f��/حH����
G����ޯ�U�g �q\�� ���Y36�3�������k.0.�%�ܹhA��E�:�/vph&8;�gݷ�d��+�28[�)�qgS�Ԫ�1_]^���+��8�� ��.���E#����'�]��_���4���N7k F����	�mx�͜쾪6J��U��vp��3�NO)�Ɖ���v�q�����%�Q���'�?��g�b_��>��&_��W��0�aI8����3��\k��l�����)��k���Ne�9C�Ǽ\����28ʓ���2��d`q0�m���(���7.�wٕ�k,˒ڴ��eK����a�@��0��=:K�w%)�18fD�b�y���=��ڣ��-�#%	N�~��;��y�>����5��˯跿��6_C�9���	:::�V��&9�`�����u-�� @�Ͽ��vww8��w�a���$�^6[RrNIZ4ku��r���A�b˶�0�i)���{�9(�h�!�fT��N����f�W�u�p�l��#77���v�3��8�͉Fo�@���3K����5��2K�5~������*����;�{�� �R �v���c]�s�rC*��f+�#��#�F�����:�`,�X�RWL(��s��,p_���~��gY��jk��R)�0,g)7�%�F�` gHj@�Z���֔��B�{��R"���:�n6X�fOO�s����)���Y����G�>�\�ڮ�P�� 칀h��D� �D��s܈£*]��*�<���泞{�@Z�-F6��[�dro��(��Z*x����-m�A\�d���A��j�F6��`'�#��v����x�|e�qV\��W���E��Z�"b]��Od��R$+c,�T��qx9��e��sY��O7 ��u�u��օ�~M?_�q�j�\O̧�b����+����7�?;��W���q`I�h��>��}�v�m={/���Ӯ���� ˝6�ß�LdR��#���O<�!Dk#Ff��x�`c޽{�����66����&���t�ݢ��Y�Ђ�R�n�^ap	����4�O4ܶ����'����/�0�@c	Q�Vw�Ja&����_�~�f&/,��'���~�����~�3z睷YW��q���Ւ��2�^�/�) �Rg��}6�����K~
��1�%��I��ې�'c��2�M^]3�
��5$y�4T .*	 l���%.	 -M#��h�4���08���Ɠ+4��ޠ�j�&�&i������W_}�緹�E�����E�vH�=X��G�����x���m���܅��R�W`q���ݵ�������?��^�|�`���>���
��i5�1f���������$����#����o��n,z�Β7+�+4��	m�W/_���k�B�}ye��ff�Un-�g")�Ƌ獅 i�}q|\#4dW�2H˶x!��]a8#p9F�I�pj?}���ӁS�(p��2���震:N��k0�s4�57�ݲ�B���Y���	�˄s���tA��*��w&�F6�b��3
(�.�G�:��v�	 珟�Ɂp�p�.��g�~{c\���w��~F��ȼ���m�Z�����/x4�q@_�f���à�������>� w{��dWXn�zn��R3��b�B�z�Ӈ��<aS�kiN�3���c�$�d�&R�PD��++�,U�����Ï�ч~H���g:f���ߧ[��iy��_{{��ܻ��E >�Ӈ��O��.=|�P
�mo�X�HT^H���:W�����ZX�hp�a:�X��i��eg��3�o�֐˜�����w`P̋�k,�n���ڪչ����"y G����"�k��������3�(X}`ⶌ4@ ����W�M�ű�09��ǤȀ�(�f����.�� ��S<��q�S>���V��Bw�Rp�� �TkW�'j0��;`��b��#�����ik{�nra6H�xv������N @�1;,�![�,��[.��ޞ�wx_���)K`��1f��-���fr� ����b����/z���=� �3�OQ��l��>z�ma��7�PB���ӳ�`[тN����},4VX�]6��{#�odb��&`%��輦�^f"���c�p;KM�k�����-�;7�"X*oKO���O�w;��]ף&ڞ[���ٶ/�ܗ�T_�ζ�@eCݖ�=�Í�6������I���6��f���S1��:[ԏn��;�fa���2�)+&�Q�D�V#?���M��#�]9`�\�"f'����^A>��ۢ��$u=��gS*���.s�<,���
Х<S�mP���Ac�)�̖裿|C���w��=���iu��X X`���C�s��o�����x�?ff���6}������`��,Ʃ	No�����K��T��ѵ�f��4K�7��O��rt?,E�t�}os:A��C��2�˩Ƥ6��t�]��Ne�H~�'�̷�镵��(>��0����"K,@����r�g���n����ŌZ�`3�hD���]\?���ai��&�P����z���� k��?8�}7[��O,�#zxf	cG��98H.��SM\)��bI�Z����|�@/>�����m��'��|�g|^�62���U�V�]jd y���cw���\@Q'|�� �5���r�Ƅ;��>�2&xÍ_�;�,u�n	��5�?��#qR���l����Έݘ�ǉu�3�Rt^I�#�ld7�
���1b����@�fc]i�2�Ł���ldy;�A��)��RN�	ݶce�1[�v�t��n�P����E`�����96Ьb�&��ӹJ�{�����#�i{}�Z���m��x��`S��`t�� ���&�$:���~F62ؕ�����🝠�0����|�5� d%U$5���R�7m�ij
�-�xy��v�X`���充%�����������/��~�-��l�/����7��u��?E_|�-ݽ{�&'&�o����ez��}���6�����>�{�����-�fkk���S3m�F�LC[#�{��Cj��hS?N�H���������vOt
����n��[֞��tX�ȣ�,�4��ɣ�Iy�M��fQ|<�z�N�{���!�r��-f+3c844"�IW���͂����I/_�����]0�|���܌ ���bP�O'F�L��Ɍ��2�9���*V\�6~x� 	_O����� �gփت� t�ɟ�D�\�����Y�q�;�;4�;��������2�l��a5�3(���ְvzjEB���>ߣ1�uny�j��)fW�u���v��qcͪ �%����2�]e0���[�
��uQƛ`��c�k�b~S�����b��j�����6��ldWײP���������}�\C���1�b�hU��go�7��6��7C�k���I�z�f
����m&hI���J�w�88��k�įi��g�'����=���������/�l8�P`ٜ�@ԣ�Z�9�EZm�����AK��F`	Bڢ�S�p�ãCf���E�JS�U�� wee�=�G����w��?�I�W:<��{�����~M��/�Ⱥ��K߹]����>�pa��o=�{kk�z�5���1	��{k|>"P������� �0����vB�1 �!]g����,��q��4
.�$��T)�v�.��j�c(��d���vLS�@Ь�g�{�"zM���s�E�Y��wA7# b֏�,�v	i���W��_A��]w,�m��M�~C�gO��]-�0c��� y��OWΎ=_#�>��빹y����	�� ˺��{o�Z0�a�G y�aٜVS��j��cO��4�"	�v�霱�)>w0��>���yi6��p梊�kC����]�,'�� ��C2ǅ�>K9����:<<��"�-�Y.�������ro��7hl�h\�������gπ��Fv
3�����᥎#>R��k/��}�U@I��{Ҭ�N�\1���L�������0?yLס����W����l��5��J��$�u��{ʿ��8�w8��$�%^c{�9h)G��\r5QV<�R�'�ld#��b���ꋶ���W���!�w� � ���Ϙ��D$:<8`�
���V�ٖ�z�����ݿ�~���R������W����I_}}@����O��k�����>`�Ș
���g�~ʠ�?�!=���g��hD�<x@O�<a� Q�����Qe*'MN� �� �s����z��@�"V�De�<��kM��K�`�O����ӱ�5�\�yC����t�C�$���/��oh��pAۛt}f|l<0v{�,	Q�@
�W�'���`.	+Z��z�:䀍K�1���X ��$L�`�N�\E�Z[��p�X��J��|���huu�ϹV�1���q����\�`�,�p�%��@�Z�`/��<�ش"Z�>Xy��J�T���ub��o�0�qop<u>��!;:<�|�8>���TF���ߣ:����8�i5:�gR��$E�G6��k&�a���׀�h��9��
 ���#�$;Я�>�ϸ˿��1OX�䛈�,ʘz(������?��-&���ڣW<���$�,�YY��ˬZφS�E�d]�p����~y@Y��~���Z��
��R�� �e>�|4����.X
�R'4�����#��)����]�)��I819A��T�Ԩd���� ��ф~rʀ��76�9jPzv�BT�Q�yH�}�����/_�mW��[o��~�Z�����ãc��ۥ��=ZX��B}��_���>}J���3�P~����wߡF�I��|c6�4�����A��)Z\�f�
��m�l���i�¦����^u<:�7�D�D7��b��A��z�u�Fv�X��w�t!��i:X�c_�/�Z� b��/A������1�������������h���ߩ�[������I:��2����H��u�a7e	� ����pw�����9f6C/`4����r��-���޴gcA�H���N������,�?8`I���L�b�zi���x�Ǳ#_|{:p����K�paD�L��gr���T� {c�3 �p�s�,��A3t}�:���Fv
3��k`�[��`�1�]�;Z܎�ڰ����ʓl�_GvfഒJ�z�����3��M������dm�۔il=��ļM%�I��~M�	�Ŵ��fk�V�D5����mx�x^��?�����a�]�v���}��&:}�˕2��c���e�"���W�^�3 ��z�Ͽ�����U�Y�>������I��ݟ��J�-���C�?���Y���������ѣ�tku���� �ܻw�d����G��< "�W � ��p
�M�s.%��j[֝�+z��9m��p�3 H-���ןc-����*X[��)Ĭ���7{��'��
*�b�d�����3n��e��-)"�A��@�k��� �9�C���Zks�@�f1YN��
@�����N���貞���U��RГپ�HF�Ϝ@��!���P��8`�2$v Xc{H�`b�f+׃��E�Xӹ��q  �J��U���\TP���`���a=�N�g/#�_�c�qP00�,�����c��N��g��M6�\�]�E�H�bdo�e�*��ǝ~��A��I#<yd7چ]o�����{�^�=o0R�pNx�*��EVD���=���5.5{��I�3�mL_:�s��|˵@}7)
�a<��$)�Ҍ��4�9�h�B&0̩��ܤ'��N&��A�썲�w2�3��J�.�S�n���ŝɃ2(�7V��ץ�Z�[h���ӫ���7a�$9�=�� n��MJ5\Q2펍���1�͌I$�(J"5"���ꪮ@�����{xD�;�����n�������}������n���"=�4�yB��o����_�����^����O�B?��+Z[[�Z�B�~��a0�?��3��/x �������^���<��{�ӟ�D���bds�s�loOX��_W�MH�  �ڴ''���w���K���u �~��k�W�����7�E�&U������u���?^�q���	�B_�����&|�ߺYjY��b��~0�v��a�{b�֦������E ��ĩ�u�֢��\��IuH���Rh��X��W���a_ qq��AuWh����ra��}f#�!ame�H�v*e��$ 8�n��D��#cX�:֥�ʅ���qM�v��4-�U�kժ��	�}�ReuX ����c�:�?��Jq |��3�*c��+_���|��=u�.�?�������v�9����Ӽ�_Y1�v^{����l�=�H_�t�o�ߞ�8�u�˞�0};����I����ֹ3��s�q��D��fM�'{�<a��Ds��l����3Q��MEπH+��V��A��ܭ��N��`r��K�YAm�C������s�J���=�6�z��nVc9��*����b뻙�^�!Ϻ56^/,W 
�N��f�v�� �^�
��R�,i��'���7���_ңG�R	r�>����?�ӟ��g��/E�;���~F_}�c��������۟Rs��@�#�c~�X�\��1�y�~��g�֥�ez��%�a d����F}����౻���kz��)������և����H���No��}��v�̀�\�CD��]K"� ѹ~����%
�r�p� 48:�^:<���t}�W5t��%{��g�	:-2|'2� �ajY��c��,�hlB(؊�^�Է�/��8Lk�>������&k��ԤP�S�R��������=�\Ӭ���D�0��m���V
�f?�.+!S�H\��=7;ˠ3�LH��3~�Y�`�v:�-�����>�d��`�dcC���y�N?;�l�����L��K��n+s2���^�x�ߐ�8�7�i����}��瞬����������Y>>d�Q���lf�M�w~���12.�:�q���]��"���N-t��xba��i����Wo��R�^
;�]8F���M��g�9���������j]���s[��0��>ߊ�v#�+lG�Ʃ7&BQ�x��ǲ�*�(��Z���/Gx�̣K�')�'Y�2�d?
,�ܗ5�]!@&E1����T�Iq�#���ʱ' ��ޑ���y��U���<�Ɵ�3���-���}��r�;��ɡ���Nz�{^�_菉G���2����e�_ ����C[�t��䈾�����W?.���e��~G߿|M�7����|�}~E��z����o~�������_�Q���6k��90��󟿡7o�P����`f2���2#����Y��99�aFd�T��e(����1m･���t�:����ٱj|� �S��o���&�a�( '�V)���D���+�����<W�:W��E�7ȏDr��6�����b�s"#r1 CU��Ls�2ش @g���13��:c?e�Z�$+\�oii)�,���{F1����<���g��۷qA}�V*$#������,k���N��?�V�7��fC�=u�a>'"^�؎�(���v���ȞXX���}����]�<q� �n�� �X�6�0�nu��߸\�qc����`����65�1ơF�A�ހ�̸��o�Ά�];2�;-�ˇ�N������Sp�7T���hN]{t��C*�O�"���\Ra�=P���$�L3��g�A���y���v���|���~kN�*x��ͰO{�1ﰍ��O^w���M3F'N�����?g��)�B{p5�\�]�:\�Y����Q�2�4>�65��\I��sȾ�:<Id粭`=�fΖA���L/�ܔD:2�Y�g�X�b�r�r�;�����=ӦF�'�Iѳ;w�;f7,{��w|u�3L;.:�L�.)����f����o����Ǵ��=}�͟�G_=�_��#z����7�L�������'��'����/���G43;��`)���sg>:>��^�`�fHf@�@���!������Ћ￧/>��Y�`+Bw��P�����^;��*;'0x=y���O���A�sh�~�_�3umt����M�K}R����
���_����/҇j��20!2*��A̠c��/Þ�|�n� +^f��z��a���p:�X����-..���5�un*(�wZ���l[HF�mB�A%b.c��'�f\$6������}��E�Y>X߬�-��KK���la|��f�qQ�.k�p���>2�V����ԁ���� �K.UC:��8 d�fWԟa��p��z�v���䲻_�ƌ�� �Ӏ���M,{h�/����c9��Q�H�=��}�Q�����VXa�EV�d�VXa�0-
wB�',}$�p$ozy0��}
��W�9�U�c1�/�'���'�aD(aoa��[ �J������$Á���@�X��'N.C�f*����� ˅��3���v�m�q�x��;:E*C�\���z�uJn����m����!�d7�����hf	���}��?PpH���E��|M�ء� l�y����h�	=~�J��ٲr��#z���}�Qc�F�G;�J~��-��թV[�^o��������$�:�`I���E��u�я~Bo7����.��~��Q����6�x�-���'��;����I��1��;�͑W���n"�eӫ@�ɲ`X������-��'G�����������2��,�۳����&+����K����h�)�������X
����|�(�7&ˬ�3o$�P���C��5�^�0 �8����o����k�Ɠ�����.s�G"`�~y�h�?W�/)J ��j$�83ٸQ������Y�`,CV����&��&�T�֕L	$! �5}�QcIg�f��㢡(��U���`|��f�*�z�F-�s-$�u�i����>�/� r�#f@���|Ҧ�
+��)�K^VXaw�>E@�iGT��i���8~1H���7b�=���Gٺ6­.k�U��SK������wQy2�X�03����W�.ײ$�QVs�}Yk�T� 8[*a?%W��ͷ�,̅��cC>^�Q`9n`���Ʃ���/p��t��C�s#��:���9��稼ݥ��2�ԫ�B���n�������Jvn ���<�js4ל�'O�ғ��4�0K�A�Z������`�JeK߿zA[����O�?f�n��K�H�13��$�F �!�S��Rj���xDG{ttr� ZRJ�s���/���������4���\s�
fT�zQz�ƥ9�������H�f �q"�FM5^�@��X�Ic&�U'%V�L�G�g��@T��d����ZN��Ġ���������Ԝ��`�2�D�ݛ�z�+ �N����J���H;�A�d�;e>��ʃ>�����e`�֒*Gyu4�9��--.���k��s�s�f���6��`!#+��W��:�����)���6[�M;;��9� 4� �q?���5�
E(�9�ǽ�8
 �anv�������y�)�zX'����{�6bǙ
�~�ɂ���%�3�3�ʂ�w��| VXa5%��W���
���18/���eѺm.w��av��|��4�#���,G��\���r'{��,7\����� �㞃��C`��bF�Q���~MK~�4M<X-�A���  ��1�����/rr��v`���m7,�3���؟�
�(���zY��;���,��2���%��Ǯ��� m暖VV괷�K''*A�ק�V���>--/���"��Hx���3z��5�5�������9��? ��M��կh�ޠ���'tttD;;{���b�Mm�x?`;��yU��=TH[ �r!;~�C����?���5���_�������S�-����% ^t��n��5���v��8G�V���\Tn�3�'-Fi �I�1� ��k�F@gm���Gؿ]*W*��Bwֺ����8h�5:�H��%��N]_�N�՘�M)�/����f�]�y�Qޕ�ZY]�ŅEw^�/�o�:�ׂ�`������^�����q]>��["!"�u~��?7��Ӵ�}e	T��j�Q�l�1e�v�wD���b&3�XSު|؇�c���l#�?�>e0`\l���
+�>Y*VXa�ݲ�}�f�g:�4��.��qs
�_gv�U�Li��rr�1C)�:��yz��y=d"��[9��UF�;n���,?I6O��t�d��<��@3�p<�0x`�Ha9�a�eKݗ��@�3��\�gyת�J�`1��z\"��"d>pf��:ҏ��;]����<C+�trh�s��:[+[�E�V�zi�q i�&=}�%}�ٗ���Y�+�|s��<yD՚�����������Ǐi��;z��;Z�=�����:88bF#�$h0#bI�z}�ڭW����̬�ۻ��	=~�D͹�Ύ��o~O�������}Z{�F3�s��v�O}'�n@�E��d ̠o�#��Cg=��dQ��`$��\���&�@��L��].�/Q?�>l�C�֠�L=��a6���_�$��t�~=`h�eDn!�� �@��|�5�Iv�e��~:`�:���������f3�=�������L�+0pz��'W�-��ĩ�'��2dq�"f��|d�r:�n��7�m�6��\����~���T���9hO�qM�r	:�3��V�|L9���O�r�4�1U����F�w�=(^Ϯ��#����=f��떵�1]���=�τ̮��U^��n�B�/���iE�*���
�n+F��v~gr��/3�Q&�ԗ��Np>X
�비�H���r�%J�����o��:w�B��uj0���Vʑ-c,��8� 9�G�h�J�ֆɹHe�^r	�K���	Sa2��(����ݤ�h�톥0ƛv�h20���e�>3y�r��3� ��:`r��S��qz�6���z�D+k��m��}tD��q���4��e �Y�zDKKO��O~�m7O�V������-�����l0�����ѻw�������;f�����Ǡ����>`��	
Q�(�����`@�{���^������o�@���w��şiyu�>��S�����.Pe��$;�^#������!�*�;��Ct�m7�w�ͽN��;���Y�5y0�NXS^V�D�Մ)rҢ~����D��;R$Ͻ��u�
𚲎�,ŷ�w���.���{�M����(8�B� �&���o޼���=�+��K,[J�d�������g��6�J����d�1��v{��W8�yX.����-)D�0�1 �`|�Td0�U.�7�\̾��{���L��34��ecI��0l��R2CI�",�Z�ˑ�꾥�몳�
/6D"�XZ����<�;�s���0�,R3���v�>`��wݘr�v}��Ȣ�VXa�]�]6Ϸ05}�/`�i���m�k�,~�vZ�.����O>���w֑ω}_҂�k`%�>��)�%c=�lt]�^��f���M���_�������B6��Q��_e�3{9�V�'���|YS��x�e�^O��Ɍt
��,-.R�m��^�Z�u;�����v�G�{{��7�hff�fg+�����Z�8����'Z^Y����o�`��ʏ�q����~K�l�Ȃ���O'�6��=�T�>0��)�ٹml�c	�S�-Q�{B���_����N�����ӧ���/��'O�2Pi��2)0��+���YwWf���H�����{����KK�Y=�/^ppDٻ�d�h��s�l�0�/j*� ����-z��%��B"fa��RH?\���3�$�ߧe��~��z�̼�~[�c�q���+g�Z����A�#��8 �Y�+����;�����;�*|*.����/�����z��`Cc?��<������Q�%2���+�UǶ�I��7ܳ!�-�=�hG�+��{b�1���+���
+���ƚ�>v?4̇�Dõ'��F��ks��6�F�ڃ��[??�y�=}��J#�JYߧ��}�5C���f�dgJ���)g�c~m�9��G�5`Y`ߠ�a�Y��k�ƕ��l��\Ԡ�u�������x�sژ���g)��(f��4􁭓I�t�>�ׯ��tЧ��?��O>���u����$�>����.�}�A�~�=-.6�ɓǴ�{L������$�>��������q���+�� P�2�E�~�J���?^�?��_������w}���R�R���	�� �#�fL������:0b}�4�{��KC>v�v����><oc�������o�]!�6ty��k�����KP` ͱ��ҏ�$&����x�Ѹ�}>����Y]X�G�q�F�+�Q�s<�����Q�K?'N
C��r�RpO���i@Q�Z�p��u��_���z�Ɵɐ�P�JFC�$ �|5�O�� �+S��EFK�9Yaƾ �c\���a�k��*��}�-����gA��R��.O��D'�"V+�2�
��61[����X��S��@-�e����aߵhbb7���b�P��9w3�̾��8�ƌ���\�5ϓ#�ѱ���ea_[��ؑ��=$'1���//3h�\�L87ϖ֏fD(���-2� �3��垰�8�f���%xMd��r��a�*�֟֩ӛ�~N��(%S�S� ��^�}A�6��N�����{5����d�^�zEo��^���'�������ttt@�jC
�u�.�\4L�\,�NZm��4haq��W��ߠV{���6�~���/��7����gϟ�O�c���/��X��b@{��fr��A�QT1�ۡ(@�E�? ��[��L�vL�rnٸ��rL����S���2~
�f?�j���&R677T���[Y^�GJдB�&zI�E��|'��8�������d� ����5z��	���e0��~�|�!nTG�`}��S Xe0���Ib��`�"�����Y�k4��g��u�@3�t �����Y>���-ׄ�|��#i��p�V�b,��Z����\q 5�P�p9��F1B��Ⱦ����v�E���k�����	��\��ԓ)\��
��6����7���f��SU��{�V�5����Ԝ��p]V��;if̂��\Į��]�k��Qo+�4�~|!�T���g�II4��{cRӸY���98�رxo�6.G4�X �#��8uf�(�hl�	l�+��C)��J��A��
�`�����*�?^�RҤ�i���m��=�zu���h{��667��f�?.1��W��%�|��][����/�~������?�)[/�'O�hy�1�A����L�pye�f��XÖ�BKK���'������;��?�������'�}������2�t�jQ�}"@���� ��[Ƀ���*����/�w� �/���s�iW��C{��~K�(����alxq���c�f�#��ŀ�۷o����(�8`Y&�ƿ ]8��`���� 7�GA�>�` �|��i֯�Y���@X�e������:~�1�4,�\�s��l@����S� �20���c����i�� r��˘iL"������R�ցs��~��9�m!]A�=�R9;~���=�D�s0le�Vx r�7 �8s$�������H�FN0���
禰���v<��7}5�h{#�e0�[a�v�M W��> ��r}���q>j�\�g��2t:?��Dz�8���)�����i�~����x]�9G&�c�Y�ѯ�:��p?;i����?`9�V��Ā���A��h5������8%�1�H�^�R�g�Vo���L��G���J-�����z�z��6������'�gT���qD3�%:88�^�MG�{������P���a ����*��w�>0�����}yHv_�������g���?��\����W?�����-4��뺟yv�_yv��4��P��e��V�x�ׄ����Υ��e)��x��������RN��YkF��Y��$zه#�O��9�\]]����t||�:��6X�ayi�33"�2]���F�?1��X���#���*C�������
����|�s=g�/��@���
��6N<��	٧a=�ԁ��ml��ܺ���};� �M@��ٜ�~f��Ct��R������oR�ݣ�I���j�A�sٽn�����R�Zg�B�����5ǢF�E��ȘȎ���� �K� !�C�u�b���q"ǧ�Z��"'��I{74�Xs׆��
+,2{�w�e-�*���/������y9{c�d@9�,��N�)���>�1T��M4��9F� #��N&��c<���̔��g��Nw&Sz�E�9��;��m��&TN���x���6����,E*���ڑ=����l�G��҉��f��c	� 3�[��
�>�G���ѤӚ���G) >�~Ԭo�Tfݱ�O�(��3�t��d� �\�T�\�ѣ�D�j�*��~}@]�'����]�=�@[���v��ٙ9N��v��_��ie������5���T���_J踵���5C�n�5�y��n�@��	����O~�%}��\��@��ng�z�����@��yl��2	��݆�<�5Պ���a%�/tc˲�ԁkvJ��͞ �fs&K�<C��q���&� X	��y��w�'�KJ�@��L0o���Kf���7�L/_����}��_��f�6���=:�Z'|���.@�r��`5���۷�ݷ���o<����O>�gϞ�= Ќ� �&#�g7T}ys�7��J��&�v�haa����5�"�Y �ݭR�i��2�����J��״���������2Uk%ިRM�&�5�uZZ:��Nvͯ�Vm��j3Sf�^+��r����G�����*�0�-���믿�b����2{�(��6�8ilw䊈��������p7
+��;cî��/?�F΍۸�w�њ`&w��$�r�]�|O�\���9��Y��x��-�J�o�Y_h���s�����Pq>�։������P1�<4�@4ʭr�=�������|}���B�6��jN��ƅ+�ЯclC|p��C2�h���Rz$|;��.�Aڝ�5m���(�4m50�����r���,����π�&X�O�>�z�N[[����6�֖�`����iQ���m��L�:�ml�jR@kkk�^�~��At�N�͠n��f�Z՛�?ܥ��#f3�6����sz��1=z�J��옃�	�a��D-ne%�ң���
�4`��u]�=�����s. �i`���j<�ݴ�C���+�0*f���&r���\�K:Aq42�e�x��f@�ٙY����yB���"���?���=�����A�s�a28�A/m1�?�'o߽c�e*��'|��O�J�<l@Y��o��ˌe�//��@Y�������|�y�\�,LZ�})�' �o��A׋��?�� 
CC /4������Z�D���.U�Y���Z=��>���Ϙ5����:�7��&�u����@�Ǐ׳c�;/��טb{��i��Mǿ)���
;p�N��1c�Mk7�C�X�w݆X��W�^�3u��-|X.$���A_� ά�#�_aw�T�3u�=���b�b̀�5�_���νɁ;�����<�	X��ў%$�S�G�o� kY��SX<)n�%ͳkɃ�7x�Q 9>�ܚx�7i8�$̹�Ld�0��+M�����1l��+��P(Ĺ�Q6G�,E�w�wJ���l �{�v{��	Q�xa���Z�ќ����ht��9=�^`ph��+�K�:O�F�� g��Z4;�O��
�;�zm8�'4H����=8 :���Lc��w��嫊���'
�PP|tt��A?��@�u���>}ʿ�ڎ	)�`rr�;Q~w��K(� +�,�1�CR`��4a �����v�P,pRwLw8�yf����͎�-�r����>� �	�/b��[�鶺Z�pBD�=X�N�6�c��:��}��H:d?���N�8�gO�{�]�;eŎD_mԖH���}gǁ~����Y����-..ї?�=��Y�8X���2��p���.�U�JY�A�����j'�j�d*���Y^^�e ��׌
����2���9�mW)���C�>�<X�� <;ה�f�)�����ѣu��8>:f�ǖ�1nue���G',����L������5����-_(�ݛq7lX]Xa�v�M/4�d�m�3���͘�>�a7��rj�A���K��^�nW*�|�X	Jj����I?߃T�ՙSd<e�'�0"T�&e�u�u�����|�P��Pd��+�e��>vb�<���F�Gz�6>S|�[�</8L4�'���~I�=����f����Yfn	W&�NY5��Ʌ���g���0��_����"sĻ�RV�d�����֞BT������;h���=k��x�17��K?�ڣM4�5sp؎K�����V7z�D�~���@��G4�0O;˻��?G+�M:�;���#::�P�K�n+�=��*ѠB������-G�-�r��׸h؇(���٦��Z"���괨�j3���$��5�m�`�w8%��0���mE˖!tD��8/��Ӏ� r�,�d"��@es����=8E�8(��g�N��)j;�����M���Ib��\j�)�X���iZi�ʹFsi9��
�M��x�>sH*<^L�~�-���ݿ���=}��T�m�C �L"yq�Sz�z�C�^������y���]����g����_��_
h���N��'X՗B�O�:����,5M����9e���9��ؒ(�mݒ�H�4|&����c��l"���D��4�ۯqw����Mf��/,p��2�R�x�	���ߣ� ΑS���v�A%n� ��Of��Ԯ�
+����A�1a�	Ft/�*��Z)
[*3p��6g�u;��t||���jU�tbp�$�F���)��9'!�I&)�+�ɴ@��n~�`�/ZeY�{���.��y�F��M���P�s��Z���
c3�0�8�����q��i%�Bp�*�#�D�'�c@������%^�i�5�hfz2+��V]�,�ԃ�:~�/�x�J���S��Ta�n��|
CP��\��\T6���a4��,D�=C���Ȯ��^�4݊�ٹAyum�S�۫˴��G�G\Ьs<�N�G�V��n�9�*��@e��t�	��37?� 2�Wk��]�zC�ݑ���AjC���IA�(�db��f��0\!1�Je��┥)o���(��Pޑ�����O���M'>����,�jh����g8�7���F^[%S�r6�C?�D@1�H��� ���&u���W?�����`��h%>W�� ;��@X'(xy||���2>��O�<e)
HB@:�g��R*�2�Wp�V���Sf*��*	�+_��w/U[қj��[߰N�t�-%�7�F�T�r���H������U����l��a�s�7�� �}>82t	��Q�VXaצy���X8>-�y �2_���~+��'eY�>��].l��Ï8�:�%.x;��f:��3z 
��v̻��g"���h[���K�ӟI��/��u���/��)�:�Mr���N9c�+s�T$?�Cc��+-�5P*�Sa����0�8o��x\1JDvMb�Y�sWŇ�
D��Zn��Pb4�9�Q�P���'���C(��/�X��!˕�g)���3�M��>%%��0�o��ia7gwJcy����������Ij4��`��5�.|�Ďn��l*�iff�fg����Yj/����i�u,�ؠp��()CW�ˎ4;<q���̩if��c ��K�r��^Gi_�ڞ�]$J"9 BT�"HL"�`�$I*ׄh��$�*Ǝi��]�ٝ$���S���S�ɠ��f<���Y�'��A��Ӛ�ą�.Y#�R����Ԙi0+ZȻ��tp��V @�d�\.��m��~��#�Ap��ˊ60��gϞ�v�JQ����gU��Е�M�p
����~�G�j�](6��4�a����1��
���W�`t��s;<�h9�#ğb��s>3c>VXa�},��ið��7r/���I�M�$��������7�w���ӱN;����� i�N�y�)�6W�W}����U�\=b�r1��G��H��~�n:��ڭ63�;�6�=[PII�<�i��e�D�0	�,�[\9�#��ϹH1`	�\`�� �[��T���K�a��� ˍ�H�1��r?`�k�[���57+�oL^�e���N��[���4�AǼ+0�a9y�	|��Ќ'�i}r�k�L�
��I���f��,#��s�%xT~�ǥ��(�Vؽ��ƈ�P�0 �x��6����h�c�5qЃ�v�L@��/�V����@&�����sNo��vF����I��8�Nz��sA.06�
c��6���E��+ȗ�װ��!"E �*Ñ�L��R���)�&���� 9�����E��o<i�6�eۡ��ŬFb&ޢ(��U��0�i �Y����wsn��������6ml��I��I+�{��=`�
�aB�EV�c��f�����D�����"͂�-�?�z�_`I��6�U��i���`9��g������w$p/�tv��Ra�v_,��) �0�ks�{g�ǜd��r�E}w��i;� ���d�\<�kT*>�  `��'�(j���{:<8̾���jd�v%y�Ӟ���g[����{�m����=:8<�d�v%@�g�r�	3Y{�Uk�>��
��MV�Z[]��VrC�[��8�)�����s����tp�O��{�le\�`NR�C�t���O�c�'K��C�|�W{���^Q33��ܥ���un3�`��{��$Afp�X�c�>"i_"c��u���g��֝�!BE�@�u��!�Q+?l�a�j���0��Ɓ=x�=H�_HA�w
p9t�W���2H��W)ÉNxc.�W�2�X��5
]5%/+ ウH�j�@n�5�Y���V =$L���F��t�� �;ڠj�1��@=X��z�[��}dƲ�Yzk��k�N��8Վ_x��9n����&�&�)��(kC�ڸ��2G�(Cq�i#�raJ� g��%�tI��X�~����/�>�5^�֯+�ì��=�N�����eo����|Z��u�H��Oqd��6/c�����
+��{ew}:�]YK��^�y�8WO#q���rfWp���x�K�:g9�Y��B�>!iTXjnqq�4�~+H{��,����JKK�T�=�1��<�2�,|I "C���$�c_E�"LJu������Vq�m�0�$=���]�L;oM�K�;�g�����2�	~�	��Έ�"f�%��؎0Ē2�8�����L)���L�0�CS��3���;`n8c��XG.��/ԑ򵇢��B.N�i��r:�a��S�����$	@��3�BN4������EŰ��ކ�cP9,9�@��,w=�*��s��0��U�:w�8����=�Ȗ!�.z��D� ���Ȑ���4�wC
�d���Ρ�<u[�kv�
qI����>2�)`�fz�)kx	��=};��]'�h ͻ��?�Y��l��YNq�����)Bs�>��!&~ݮ��Մy/��~����XYYf���V��a�Y�&�ЀC?�	̥rY���;pR����̅��cY�k�r.T�é���hW�*���!VXa�ݸ)��?�@�����Z~�T~��vvv9-�Vy��z�c�O�1�%}�3��2E��ٙ9��ܠ��=�$h=ǾH,��ɴ�O��o"���#b�!�`��XA�.��� ��G4�1���e�B����������r��2>�5��,�����,�}�:㕲����	�+1�׸�t����`��9�]��gc9*M�P 1�n�ؗ��%�̓��up��xj�(r�@
�g�ǵp��R&�,h�;RP�M�A۽�a�ƭ9�����,����i��*�Z��6�Yxu�1 �V�M��4nH \��géL�lt,�;�qo�,�	���F �P%.4��E*�� �F���D�A��Υu�ò{���v�W,���j�G������v��G@���h2���_�F��:Y��}|t�Y�p�gg%��+�B��~�\��G\�m���Z\Xa�VXaWg�CM,c�ȫs��m�ړ�i��8d`���ӧO0�T����6�;m���p�����a�ɲ��4;3K�z��<y�2��`��������G,� �D�O��/mOR�E�E�|��@d�YK~����cB��Ȭi���95�ϲe�̟e��_��n�Nn�X>�%/�~#� �\K���4��q����I��pw�xw�n^�_��x[&���h��|���=QQ��iJr��Q|	�e�D�1�mm�;+֠�q��T�#�N�6�`��VC���#r�E�@#W`&|���C�[�ɉ���O����w\�V���~�C�6R 2"S�v#p�W5>ҮQ�a�շ����[�ՂE�]�y�́����������y`�u�}�%]�M\�0�[�ʵ{m���X/�|j����:tkEL|�e�zIL�>y��~���q>�jr���D���3���Ic|�dB{RpY�K?ZW��1��9Ƅ�Ej�s���r?�lK�/�XhRg�F��Q�)VXa�6l�|e�1��8� ���eăX���@@yii����GG�j�4�i4Xz@
��R[$�V���7@�9]JYW5TVnkk�k6����b�h9�ۀ���<3��6F�nɋC:::f	�~�'�q�.X7:���J���ԆlK�@���$� ��J2��]f(���Ĺ��f��WC��䄺(1T�
K�3��P�Ԥ�#R���ja��[so)?�;e���:����rvx���I�^#XN�e�W���*IT�0�N�u��|E�8 Z�f��T]�LGN�@�R��D�Š(�+����2����*������&j���d�p��3@E
�mmG���������J��	#�ȹ1@k<���i:^���^> Q�d��ZÙ�SD+ب�o�#Z�a=��,P�2��땅�c��ez{=;�����l�|Q�w&8��a���$�rh唆:�m��e�4�Q�0<xF�{����C�ǩ���?=�\��ȱJ<9(�r=��iaw�����p>�PL(���
+�R&�x�>�vAr-d��1��䘁_�9�d����6�=�����̌f,WF�C�,(�ﳿ������cS%\lU�b�}���^0����0Pa��r��S�'���i���7�����^�pL�w�Re u`�����6�%t����W�^�*�K���}C�R��@��� ���[�����% �!!7?7���R��c>'�r���1��J]�R��/�ޛb%Ƅ����J�Rn��e��i����D����H��Z��R���w1�:��'p��8�#����_��F�
,�:R�K�ŘG1�|v��e��MP��!c\F�
t�Ԅg�F'�"��N���Xڡ�E�sK����(R�PM��������(�V��Ǳ�h�h�1��!�R
��'0�3�+��dܾ��>��j�MC�_�i��)�x��a.ݎ�-�� �i�8��1�"n���E{�5��$n`��	
H��9.�㋍$C��ሌ	/	=�YXݰ��y���qOӤZ�����Z�S�Ka7n������Ľ�(H5\��c����}n�U�����?>��>�;o*;g������Ł���u�q���vvw�Q�7����*L�l=�V�,?���M�n��f��r��|+�B� �y����������<�N(�ǵ�]>^��u�.�eIv����b��D���[�$֛���j�ʒ%n[)w��1|�~/�,;�.�!�`�#���@u�F������/s�k_G�	W��D���um�4
�P�Lv]8��#9��K�� H�ԏf��PR��C�​��<h��:�lu��{�C@�Y�A��} Gʉ�ެ�$��1����� 0�'���W����هTI�rd3�*�վ2��!�Ԏu��X�g�M��ˆ5ܫ�X��@j���nf�w���߅��c,�<�v�}����>��:�V���dr[��I祑rsW�%�F3�m�C�ۤ����T�%ςu<С3�l� (1���{C~Ď�����A�D��8+q����5.J%���c���a�Ϊ:����5�9��1�5��=���+�袡!�ex���F��p�D[0qLse������~\֠J`)�C�ϼ��1��ӝ5=�	k{�@
.*���+��<z{�CwL ��e�ܧq�*-D��r׭����]�\��OwV��~ڕ�ڷk��ta�Ht� �NZ<an4fX�V�' �d�!��0�Z)sA?�>�v��2 �3�ϐ	 ���<
�8���r�;�j��d4��|�
�b��:3�`G1����@ h��"O�/�I^ 0����h{ [Y��Jau�C9�<�Bh;�l�`'�j2g�y�@x���Sl�������+h�h�\��1GH��l� {tl�'��E�������_� 9�cʮO�H������?��3��J���-��c�?��Y�h����8£MlD�
��%JIȑΌG�?��Hb���6��ln,��z����j�r�'5���3/��i�=�������\4M�xG}x���k�����v���	�+�n�������2RC:���aPϞ�"���z�ބܹE��� B�� ߗh��Ah�z��$�;�%t�"��W�m��JpN�	Ͷid��1�ă��l"��#���рe�~�qs{́�㟷q���q��;Y��h�+|C��+ɳ�VM4��)<�|�%!r,�h��0V�+m�����;5ѿ��NwȦ����	S�����x��F;��vG\��
�h�ڏ8�Ѡs��`�^q,da�
>���P��BkssMZ���%P�����A�@I���-�������Q���^�9��#n7`TV? s;��\߼~Á<���|�s��:��M)?k2�c�e��S��b��4F!ȹ���sE�<Z[cpl�y�\f�O�t�@m�C�Ŝ��?���&����e���*(��LjU�P�shK#�2`����R.9���+�6\�of�l���&)*p��>*sD>c&x�19�L�����ˊ� .�e["� d'Y���ѥ�0w6�\�u�4��"b�6a#O �a��Y�ݮ	�<���0��s4.�\����*����W�g��iJ��p��l2+n��ƿ����s� ��~����EN�&�4i��6�ʟ�SB`������pt��vYr���Xy�~��S��x��������.���o6�����)Ʌ<��&r �g'α�b&�c4�tv��A?���sv3'���9���P�-�=)g?�h��dK�)<`7��rf8�Y���D/1��fp9eGv��N*XC
�����"Eܽ�Sc���(�)99`���S��8�	���={_�3eۨ� >#M�\���ݗ!��r�:�Fǫ�8���+쮙��6��{�(AfK�xQ�]��2A��k5�{`^bM�kc�?doK9=�ˬ���[���fs�A?���T^��:|�8�l�UZQ$�fL�=���j� %����~�=mo�0�z-kS��r��"����_���c���̰��C�����v4l`,�\}����ξ���� ��hwg�%=�����%W�/�x;@p7�[��}�� ��,_W��c_���+���O\��LC��r~��V�Gmg��7d&ªTv��bn.,�C��?�y>�H6� Ȝ2��ex�2(����I;˧��	�l�2�-��|��[�f,���N�#��O ���cvl�����VA������8L���赧l�
E�r����t�q�M�`4���荈��-�L��&��1�;c�*�`��BAP�xs��$�*E�'���Վ��'� ι��ڡ��8p�
��B�8�ă:���s�u`����O�'@�R}4���~(�(��F�k�b'i�p��i�r��t���A�½0���Na��t���5�"`�$��8	I@`�t��?Y�G���}c/�q��jl"plO������V����y`�`"&�}�q�0dC��~�,�;�{��:^0��ܗ�>N{0:��uiY�[6O'���B����bׯ�Sf>e�UX.�Ú���u~t;U��R���'�>�me����nw|�I���T��f�u �5�L����sO�� �n ����������Gɵ��=��=!{�D�tii��v�l6���KѶ�;��_�3;/�~��H��6����x�A�V����⢛����<V�}����Tifn�Y�,/3�,��
�����R����:�.�ta�����=��q�V�ug�B�Çm��)F��0�&~'�{9{'Zf1SCw.dƎQ�;=ﮰS�N�&nM
#`���e���t�	�&�� ���rʦ�N)�"{x�q��zp؃����iW�,�b�ΌT�q.f
(�v8��o,6����pJ��<�SWR�g�P�:�2�>�aP��53�av��0�O�ics��3��Α��r?�6N-���m��Ш7�	�`mm-�Y���w�փn8��8J�9��Dْh-㥒0�K�4j��
?��|��S��������.�X>������z�_c�x�fq`N��w�'y����Ro,u���E��\�_]�Vص�]�o�g�|g>�!���s:~�`"ְ��,*�ϋ�b`3քu��
ד�*pF�*���f�X��=f]�HЄU�d�V�lV��WWWYC�kqTJ�G꺌�s�>��4Ԏ�.k�^H�M��7M=z��5�����" �2�������ϭv���m��޳g�h-k/h7,�R*�6�E�r�6f�3����LA�Jf�#x�676y���h�%`���v�d��>�˲�I��+�-�k@���,�/��-��4��{���~>��%��ha��oY�����J���_Y�ˌ˼N�M��SD\��I}R ���M��9��_�=tSwh���lS0%H���i����������"8������cOCE���V���w�.78����ޕr{w�K����Ws����+�2�.�*:LAbcܕP4pE�k�������CDS?�3L�u��>n2
1:�):�Z3��2��x�+�'��eƃ���!�['s�����E�޽͜�}�I��>�!eM*2�g�HJ����I�'@p��ޞ��!���L]��A�3�M�����J��Ȥ�|>M����sd��%�(�1�O��tx�x�����F�W������RL�]�=�"�FV���DG0\������"��JƙnM;%(�@n���w���TXa�]��G����ֿ�G�:a��X��)_�߁d��$���wr��`4����ܞ�	��iEv:]� �i�c;�'�e���LS���O��H��+xP����C9�)�Ǚ_}xx�l���+��%���h���^�g�;�_�.-.���u���H����^q�����?�?��^��*G�G̾F? ���������R1�5pƤ��H}���%'�!r �C�g��w�(������>�猌�
��f�ߜco�{L���Y˼�p�>�ͤ���Z�S��<����qu���	�?�b��(l�v�����'u����������>ݗ��	~6�b03
�ؑ��c�0 ��Z/w���y�j�D{q�j.m!���N�)IK����H�̟��*f<�(����(�VeD�D�ln˫�`���G��@����&�xVط��3q���X��`W�d85���v���￧�/_��֦�GP4d�7�����s�t������V�,����ӧO�v�F�:E�I���@�6�%N)ž�H��p��G9]��v
�A�F�⁮����c�\R�,��$����v]�r�y(o�{&��-�B�UC0��)�]����-�?ξ[�P�Q~�>L���&�6�革o]��l���s�d�,F�L��y��������xN,`�bɮ<H<���_�L͆�K�ny��:���D>���2�����C�@4&�!0/󴸸���C�5+�Wb��ӳ�]�tO�]��ҁ ��g #GGG�X��8��r�,��m�����o�	����i(Kp"'A�ކ�wb�ה�s�؊�7�z2� I�MG��r�Ʌ��qM\焤`O���� ��V��y�j�@>ƺ�&)�=4�T�^g��9�YڅV�MYLR�)qO�1�W�`d�{=	�Z��R�Y76���f*��G�)\@��"�e�'��ˎ,.�#��-�7��֓("����Ԟ~�Svm�,��@�FhHқx5���wj�$"��	���4�{P�J����>]j���sU���K$�^:*D���0� ~��z�t �.����{���S��k��~�ks�1���LRT����re��7o��7�|M��[��{���m��[��l�-�c&st��u�?�o��3����>�O�?�G돨V)��X>x����+�kS�e3ՠ�/����W���,}%bZ��H����uQ�h_�/f��
�@�����73����o��=��L�]��j����:�g<d��y �C�-Z�G��R^#�g���v�̎|��ݷ�z��,���q5��;S��,=� ��䡸B��:��;�!KI��K@"�	0.N&['�1p�_\X-��Ȑ�/����s���3��x���g!7�
�]��\侵��hXI�/���usc�vww�9H-���[���`�p��ӧOhee�5���\?d�	h���G^��%~�i܊��_�c����9C�Z��5����o�ǆ�8�gH�a�g�������Ƶ�X΁�z=c��B�E�.���3�x��`5�y4Kݭ?��'乿�d���r�0�^����d�O~L"����	����1��[`,O׼,5n��1��#�*��g^��>�@��첁9�;I�s�.�Ѷ�F!�4:� 薜�0�=�3g�2����4���9��T-v62�zv�A3\���9��l���	�{�:��c�R��)����>�8��:� &�8�&�YpK8�;���tϊ���9����i��B�\bPw�����{��������l���siX��܄�ډ����k�8rO�\�\�FK�.k0Cg����� ����e���^dS�7�bq_�A������\�ۻgv�>9m�1��J�	��mU1� �̂����l︴�k"N3��}�s�P0�0A�~���$��@�
�V�͙������0�1��պ�j�6���ݿ�euK2�L��{^b��>	��4ݎ��2䲓\`�\�1X������$Ad\,�|K����
�J3�J�x�h�&�3���232Q���4�3�p��� 6�_�o
v* �q٦�B���-|������	�����&@�yz:��;޻h[�_~��	�BwX��ޓys���:�\T�XAk�MJ@"�d��,��q�:����q��fi�X���N#�Xf��Q���DI$��TXa��	��]#}�L�����_d`V-f�JNBv���0ŏ�#X�����yD�7Y�80;�~�q3��؀���_�5m~����\a7j[D��Rv�'�h���0�v ,�IФ̿-������),싷� u��?w#�i�kH_�t���s�NNڜ&,
9H�}�u���PFU_g@1�Ǚ��E�4ӜgG��إ{e��O{®�T�4 ޣ�σ��]3����#����{���$Ѕ�|.�"�ʺ.9kNK����@����Љ+�We�t����;��o��6�m�}X����;�^?-�p�㉳;lW�7hv�N��&��AE����M�?�g����������M�s��B��6i �1s��{1�uZCgM��~��v5����@�`vL���9瀆Aė(E`�%���o��1�3�D�N<>:�wﲱ��'��c!�c���{E�cl�S֑|��9%á�6�Н�{�
{�潄\P���G��]bt�X�>%����_I\�<�3!11H=;XY�"3X�� ��[�b=��$�� HG� g�� �3tb��Y���+b5�X�}������ڴi�`1X�'�'
�Y�X�P��c1�}Q3ŀz��+���`��2�X0tQ��%SzR�Q	X�4��������B}�Y�Zq�:G���訣o�֘��p���|M��5�"��w�W���3�a,?y��V�뇖2��.�]%���˓=���WV�Gm&̝|?5y?#`�&7���f�}A�Y�e͘���#5h�j\&�1J6���?P����i=L�Q�9�\�4�GZ��ݦ�8��i)�|0T��αڰ�D�f�a���q����v��8j�N6��fw��Ef�hKn�y� N����������Q� S뤕9>=�t����p�k�G֑��[ep�>l������K���B����t�:�B�D��z4M�2������8Riԥ�%��Lw�|u�SP３iY���
z�o߾���������9�������&8�����	���I� �1NO&Lֱ���E��7
��w��I�_����Y�����(�.%�'�vJG�t?tԟ|�\��;����S)��7V��E������		�2��SW�PA�ā(�=2$�h�~��z�y��2���T��E��:~�Q��{M�h#��f�|��zS7	��X���{��zO�߿g�5]1��D��b����2M�I���f�>��9�N�]F�������|Ϻ�(�	Rn

�|��Dd� f>�ʪ�rvM8>�Q�g�A�	�}�?��`p��Ͳ�nkw�vwvx�����?'c9�T.���*��z��� �u��g?��g���WF�Hb����m��r}����"���@�0�Mn|���̵?t��`V#��k�C�|��õ��T^]]���d(f�$��|C)7�1�b,��
+��L� ͰP\%&�(c�������f0�����2��k��e?#[�� �⸥(��I�c�0��C�f,@7HV�(��Y-��fT�M��{��τCE������`
"Ze��e�~rԵ�
T�g֮s/t�ja�^��������O{����>isԹ��f�=:3�"��F^Xl���r�8,��J��.�%D�Kٺ�n|L;{��@� �}�'-:�ݧյǴ��B��T� T ����`i�P2t�S8�)����~X?�H�̬Y=K���Sp�-���' �.�3��=W���8�����/�	� �_��Kv������c+���6�$1�Z5���D�����&yMZ[{���hG�gf	�R���Hx�L�)��ϸ�����er�����D��=��i�9ʨ��Y�9ʢ�G���ө�x�M�xR����n�����l�d��~"9`Y��)),K�Lc����N�Th��?������K��bILk��ʹ�m;X<��ädo�~\z̜�#v���o��<����-�<��(��P}�ݝ]��ݡ��I6����Ġ'$ �j#e)[�q�	b�mb��o
�KYĒ%E^kV}�����7�(=�i�h�Y�����}Z\X�bCX��#������Y f.7�K%@�sD���7��.��0��.@��y�
*\M�N���{��9������8��8�]�]o�貟�B}���3�x>{�e�*K^}k?�=`���0���]V��1���O!ザ����2� �1��v���<���U��;�,i�2�=���������sa����C�w}�}L�t��f-
�����8]�!��{�:��2��,�+��,�8kiBFt1�<���
c�&�����׎����5��Ul@�(��c�ݓuog���%k�a.������Zm�^rO��n���~>��.���6�H�5��4x���&�s}��W���S��_��>�|��e��u-5Thuhg�;��zK�^�����o�|�����Oϟe���2��#=��2��p''�������L�]K'\{�g�l1��Q.c�;)iP ���=L����&<xLH��h������.�I�ec���� *���o���ճ�	l�6��&����(����0
�<��Is�@JE������J�����ۊ��h5�]!�����1�v:y։Y]�kA)z��{8��N��~��qo�{�5^���޹m�?��Cǎ�AlfX�z���p�Rp��D�M~Y?����u�g�S�)���R�OSY�[-뷐�@Jo��/���1H"�(C����c����5���U��z���sKǍ�6���v_c�l�&#W���y�9_��]LJ�L��Ǥ�]6�[N��]�f]��u�KʀR��倲��	h§�����n����큾,뵦��M��*Jo8| \�����s�j]�|��4��ff�I}yOL`]gɚ�-��>.����o���>�`=�c�����𐥃���əa5f�"ض�]��x��]��aPY
�ui/�v.��h(�&cf���-dR*�Z�H�V�,s<gd��-�3��xw�0i���m�'��k�s�߁�\*�!رK�6��?Ō�2�2��ls-D���T��\�7�ƣ�q�?��皳ܖ�xo�I�5�wA'�M�%Y�Ԣ��_S���
�3�Xξ|�?��\�!���\������=Ds��c���e,;d�^����PV�eR�<��5�� d�m�����c�,� �2�%��tČ�J����9�`��ō)m�$~��5mn|`��#{�β0�k����G?��˟��~�WE��Ohye���Viq��9*fS��d�/�ٯ�¬�ե%.FP�xtx�������7��W?]���Y�$ل#�����0�DH���޳B���b���t����R���pд!�����A��͛7���̬A
�����&�xJ0Cۘ	�ʭ��t��7���X"��$�+;'�:�1ECnss�b"&�eP\�3����|r�A_ϙ�	� �z�E�vk������|b�&��w�?��܌p<�cN_��f'/�~>��U���e\_���2��q��?�ϺI]�,L���Z��z-D����}�z�N�b���4�R���k6�)�uZ����Oi��m��<tn&��E�v'�?"|p�T��}/�\��HY��5���N���>S���H�@q�˚�vv�O����
8w���>8hl�Fz��]��U.K`)Tu��R��N9��rɥ���3Åi�a�K@d�����`�6���0��qN�c��qʈӭ�t�_^^������K� ^_�lSdv4�\Bʲd<ZK���� ~�"h�����ٶ�V�>s?�����nѼ��s��� �  �������%,7`6s�!Y��";���&%?I6�^�%�7'.���j�KaJ�&�w����I��%&����{���w�]kb���/Z����
�!����h����5W煌�~���c����at�e����>�m��R3c���2�I��	����3仸E`�Z�P�M=0%g��y
.s� �̜�� sd*F��N���j���@�_m�ގD���*UJ34�9;��l�$/�F������������/�� �Z��r�Q�R�#�����I�ќ�ٹUkef�>ZyM�[ٶUj�N�W/��'Mz�l�����C�I'�(}R&�FX$>�mr�t,7@�����
T߻;<��f���Ba�Xf   '�`���{N+e=@�
v��ІT�;�vs��D�zD���AfR�d~ O��4cF�V�~��5O� ,KEu��K�O�d��?L�4+�Toԕ�9P�O2���a�=�� Zy6�d��S����w�Y���~��u�'�a����xh��S>��$��f(�7���BM�<ͮ
 ����<xڜ�-�d*u������{��OI�7 .�&6��fG�=��F2��n̊�_l��η�@�Ŏ:q�Pf9�_�QίQ$��S'���e,���s�ʻ�9y�S�W�9Q��Mu��J�=f�^��I%��I�+|�e��o�t�w�K-%g>'q�gtB�~�5��,�	`c�w�Hؐ�+��|H�q�v]��I%#L~Y���XǙo�k�1�)���]�oT�@u�t��Y �[��e�9��'���H�-�3�c��g|^s�}����9!8��t�����V��:��m�v��`��&�<�'�nS(��i+sA�im4ei�k�o>賤��͔0F[gB�@�<s6d�,~a�/$ӝ��rc�����}�v�m���beԌLF�g$Wt*c���P���Q�N��?Ay��|����bo����tnXV����wj
&O�6�Fj'��4<Σ"߱�4�i����� �>�K�fg��T>><��w{\(ekc���@K�J�#0Hh~n�?~B_��K���_�W_��>��9�?^#�g����|���8�`0�Qop `�Miy���Z�'�߽�mZ]x�9�}�sne�9>hg�}�~��_�������h���sW��N"8}!�S�L" ������/�A0=Ìia���Y�%/�D�!���̸�Rќ�
��z��޽{�Mhfر��,�2"Z��r\��̜<����1�I��1�` � zÑ�����s�&7&`�i��ı���acN�G0w����q�2ߵ�y��C�#��z�����[1��� ݄�1qW81����`�X�®�t=`��~��wc��)��8���;柜~:��:���l�����z���e�~T�%zG�*L~a(6\����7��	sq� �0��X�2Đf���˷1��L�9�tcV�m܊4Ը��`����해��/z�6A�bL�!lAW{2����>u�;tf?��W{c�A~V���\��8j������ 6K���mȿu�;�\��e���nϲv�ߋ���F�lY�ޠ��%Z^^�Z�F}�'i�7*�sؗ�Mc��221�����o3?�Z�10�\es?U�� !u�&(R���������D�C �P?���sC��]�q�5�=S�=�N.9�d�bb�e�9[�V����u����Oů�*GA�mw���.�v$A�E>.��:��_(�e��C�*�K4���(����4�da�v�&R9��kr�=0nm..���]��cs���o���DN�yJ�p>�~�5�����b��9�7�XV昙��0&n���nV^�B�ఽ���P�(��O%8�,g���7���޳K�+�4�P�EUe�Dh���N��Y�����qw�eϒ<g9Cɖh�tj����kfϟGF�
UY�x݉����f׮]���L������~���{��s,����V�޼���O�/�����R�~��<x���5
���o��^O�Nd<�"p+K���漎��]9<ؓ�2����K���grrt�Eˡ($���_����em���/frs��x`����A�)����IW�_@`���p�+3�>����*N�z,y�h<���ۗW�^�9;���2�9��JO��ݤ��_�8@A��6-�^� T�c ��\I����~�������9wx�y��x��3������J&AewȇL�;c����XhhD�97f�W�'�*8��y��������ߎ9,�f���[�|8[�b/��@���x��&{�͎{��ks����L�����k#�ٞ0���0�5���:]~�4��t��J��/z�>h�:�)�X����Y}���j�d�5�o��랉b�.e1��~DR���s\7O���\]|=r7 ��"f6�4`8������,���܎�z�ͱД>����f188y/?>C�ҫ���=<�w�.��1���k�����`���Ll���k^ǻ�P��*�������K[�C��Q��&�Z�h]�˯?��GF���|Xˠ�\�����
�uɪs��J�=`�0C�հ=$�d]#%�+𱇣V�tOON��p��"�z��8���380�; 5 e0�a�:.T!�=�aʙ{"�n�]�&̃�wM���1��D�����;�e���v��U�G�I�]�/�?⁅�2F�i%�=�q8�A�׊�1�Į���	�,t�I�!�죹��\23m[7�gm�f�C�Qp������/X>��sk��5��]�����˵v��	˥y ��e�En�	K�E�r�/ݼ��rg��mӤ�F��Oݹ.V ](���fG޼ޖ��C9>�#hI���]\�/��R~����7��y��1��@��y-gg'��8/w�k�s4ҡ���"f^�I���>������<��<{�*�k(��#��.H��ݑ�9������3y�d]��NO�J6��(�6�H��J^p�l����� }����E�mm�i��*������J��y�E��<��(�o԰�d�d̻S8�w� .�w�9�R��D�^������;9=!���o��ْ�6/��N6�M���zNq*�<+�i����cy��5�X ��Ɇ�S���|������� ��焀	�Q\��R�D��R`��w�-7}}{��^g�8Y��������d�&LA�W�v�hPv=X��R�v�9��۹��%��V���<�,�Pv	���l���5E����ѵ�y��o�W��Z�7a�L8���Bk����l�3��G�<�R��*>3�֩���I���z��3,$��s�0�3A��{�p�!��|Z��������-a�F`/|=�	sY_OBb��CỎ���
��ŉ���-(8�c ��ވ��Ck�}���4[-m��I+f�\�۩��4��na�@��� ��ҳ��ʦ
�A�< ����%X��K$b������hQ���i��w�8��y� p�ޙ�u9�pL0�UZk/�)���;�������e-9�<�������d+�E�{B�o��jC�����|Eѻ|� .�g�U%U.��UC3?��^���	�K-�[�� ��,��i�j�A=�.���M['����lY�ton�������t��Y�����:vF�Ϭ��n�X��Nv�9n�G梳z�<�m��ك"(BC��Ω�u�"o^�ʛ�����XÑdż�wW���#���������>�\676e�Gk ee0@�89:��y?�֡� �iR�����dy�#��H'����ӑ<{v(��y[>x*<�����'�АBT�?���(�?����������=��W_��ښ,/���VІ1�^�ƾ����M/���w�+�30��,����(�V�Zb*��v�	l0��ãC���&�@u��� ,	 �i��ี�(]���E 9���� r6z�c��w�VM�� ��v��:�/�ȓ'��ݻc�-�4`�Lr8Wo�T��;�Q���7��{{ԇ~��Ţ=0~����:�
(��\���>8ЏLY� �x�)�pp7Ü�s��,Z�1���N������{i��˖����$3\�n�6~/���X��gE�A�Qi�Um�]`K&s�a�ڃ}��#��>���u�����A���,����� \F�Sz��O���3��A̋`s��u)�����/�km�ќ�W�f���&��j��*����0�2�)O履'���u_(x��I;��1R��H'������y��͛�{�ʾ+��� ez���j����8�� �H�x�~�e��Af�ˆF�z�yo�g0qL/�Y���
Q�"�`�0�	�%,�.F�f�fơ�pA0@R��$X<�ێsR�2q��A$[;2#o��o}�����`1�6�~�5M6�`� ����ء�1�a2z��� 1���IX��������-L/���й�50쇝0כ��#�������Re�:>�Ъ����jP��;���N0/�9�!��؂�1��{������dj�Aܟ�c${���m��b�@f��b����a.�����a���. �s�������&פ�e�剭y6/fm�nS�LZ�cܩ{��5Õg�]���X�	cñ��r����c4|	�ŝ淘U���Y!���V�1%[��~\�4~�jKv���p��F?��n{QVV���~!���#P�F����*`�`�N������kN'���c��+���^���~x/�/��F���ky��<|����:�^��?�����K��dyi9���X��'�n속rF2N�{'qR�h
a�X9;ʍ��q�~S���/��[�T���Yh��nC�� C�6�DA��PuC��a�x2�%�� c6�рFZ��Y�n�BCi���>:<
�|��J�jtn�G���6u��o ���ra�����������9^]Y� ��
�L�#k�K�UAz}v.�=FJ��G
-XN�i��<�;��fTU$d���@�\춷vN�`�ݤ���kOe��z�ɪ�~7���×��W�s�Wz�Z
A��l�Q��������.@�/&�p�c01в�ȹ�u�.��_N��^A��
:ڂ NA&��NV��N�rW߻k�z�22(���kdK&A��������kYV��J{M��2ai�LӴw�>�r[[\Y��iѰ܊��u����,���)��8α���&d����ٽL)����h�z�Gch�}j�����pOX�h+XU�8UMR��bo��z�I�������������\��D �U3��?�_)�^�,��b��1���?E�U$����}��g�i��t���)5��8��>�Z~�fk��b�$���`��F����m��4s�m �XT�%������Ae��$�2f��x>�B�6��?��e.6���Q���?%���V����DF����%�1 {R�<��t��7%p�/G��c0[��K���/�kE���?i�G�ZD��P�={�����zL7d�쟟TF+� ����B���}퀏)�0�i�׹���Xž���~(�6Yϗ���~����Y���l�Q��g�lJ�s/�R�y�4��h�Uc����ə���Ic�����m'�%M�=r��6pL����<�\���[���'���a�nё�{����k������������tzY\���t�st��Ɂ���������5�Fg�w�\���;����,��/�"�ǧd?��?�����~+��o�bm����X���|8ߙl�����)�����=�w��B���+�[����)Ig���/��mv��R���ɨ�mi7�&M�+�|r��5p�}���_d�89Y2��-&��KFjF��ɑ5�X�����q��Ψ�sQY�)dY�6�e��񳸴�JhʐE�=�C�$c�g�`7�aȢ_�����N^<N	��w��Ç���?g�8�`'Ù�ָ3U4%8��{��h@_@���o�L���Ϟ�<�A�Y�3�j\�	�h�������K_�9�7�2G��wv�W�\�?w�9R�{���m��S?q0`�+�G�A��r��8bU�bz�ʲ���a�%�W�#-���@J����`__�����t����C��ce�$�s����@/���� �2:�	P^i�2��؛RD�e*��\����I���2�I0�Y�U��vD�Ba,6��0����^���p�k`Y���$ȅ{I��%z�0VTG�>�؄�h��g�`��<7md�fZ��  ��IDAT��
����E��n4-{\;V2e_�vW���c�"�3�����{{�j��fq��Ui�=���zP�� � ��d����q}�К,�V�{�@;��p/��y�@�w<�c-�;�]�q&̨�l:��x_m���\�{�ϛ��5��C�׋1;�k;�U�~`Y8��WK�)<��#s8����nɕ5�3����s�\A��~q��Y����
���8���3��Ƭ˫t�8��lk�$��x�i�;k\~��1�v��_����_a�k�m�,y�&���,��UR�9�g�gB�6>~�K=���vά'�
��ia����Y�����~<���C��1�&Y(.Y�D�Aچu@k�f�m��-�g�礡7��
OaT\ժ俗&aMTՅ�S�-3�t�V�$�&8��a��:����qe2<_�^{����]��o����C�+;;{�����R/��	�z�|��j��k���0����꒬��NԜ���?�_��߅�����N����'�ꋯ��Ցݽ�`�t���l��_���{ON�ǲ�+����-<����rz0��BG����,��E�H4c�Ϡ�D�[֜��]�Z�C�p��u>��F D�`�%+�Q���-M�4'Sq�<��߬��Qb����1��	�g
�>]��a��k8	���G���-ϼ���t҄� �/·�*���
·kz��������W쳧�>�_|�9S��	Σ������˺���mlڊ-+��g�����`u�J�����>��{�p������yӖO����$��C�?�$bu��?�V�+Z����놲M�-�ƣ� �E�՚����ZO]^�P ����� S;� W�{5y� ����S�� �F�A�x�@�8�Jj�uc61΃��8<����q.�D�� ��B��!ra88S�u�K��26{T�q���4 ��H�O����ռ��=y
=�d�������_^^"،��DA\�`^��H���F��أ�9Y�R���
�߰UÙF׾x���ߕݒq� �Df���
��uR�Ȃ�ҧ��g�3�q/y�Ǧ&�p��G RQ[��ŭ�U3�*���K�����~\�	����W�3XY]��0����c+Fv,~�5��|D�O������$/"��Y�h�A49�l�Y�UbC�q.Թ@�	Q��<x��9�����ﭮ�q^����؀{+�}}��a�ųdfZ����sq���3E�	�@�{k��Xw"ɸ�1���Q(�k���Ċ��&�Qω	p����e<$!5س�������T����֐pz'�����S*�N#�8x��kJ�;LO��lZ�ٯguɃ�2k�6k?�)��wLK30��V��
`E�b�t1�r]�2X�{�F .��M�sr� �Y��=3��r uKR��g�l�M����v8�Nk��?���X� �u2G�2h�S�S ��ξ��^-��w���!O�~&���o�s0����sLG%�z��:d�=V�Ruf�x[z��.咵�2?7&S՛�m������^K��*_|�k����r������lj8��,-�ȣ�mY�_���,8�rw����8Z�?,�)#g����̚�>#]lDD�X0Wn���Q������^��.X��F\��,�ں64BS?#������j�r4�4Ao�s��I��VV�Ν�ߚm�I?8� {��Ů�9�}��D��Y�#���k���g���K2��޹��Cy��	��U�����{�,��$�T�i-:��;]h�-8��٥.���9vս{���$:�@���*�	�W���J�����ׁI>~��~X�.=��s�w�]q�oq����ot
���l�c�-_U����n �m�s�� ���סaM�A�����钱	���J�Yˋ����`
&��;
��C��L����Q�mtSfaf�r��^�:�J�3����P��� d��e~a4�;�N�}(NI�! �ԋ�\պ���B���������ȀԵ�2s(���*Y�f��CL��ߵ�5��k�������ed�C}6Ԇw)8M�*��g�ݙ4
�z>e7�9<q&����P�ZA�q� C���>�Rc� ;*�>8<<"@��q`�/�i5�����*a��=dq��ϵ�:E������:��ݜ�S�3��~0�.��Ч�> g?��ʢ���:�;
}@��}��`�Kun39eR���qi�,�YJ�q)>
6 ?�ۨTft�~�/���ݻ+w��p���AKA�b<N� �๠���O ���s#��9f, �1��>�f��ͩ�b��ϐ遾q�ؗSw�Lm�:�
��9��]dS�yj�|��Z5e�]>n�+̟f �}�(d��z��?�_e"@���y��h\�3�GZO����gm�~L{'@��^ģ&>�Xmo�"Zc�7�/�?��!d�nUK�/���]���~~ܬ���A�0.��> Z@�^G%)A�uc��<�,5�H����'��[*Ђ��(s��� 8���i�l��^�����!5]��/�W��2����,/-���qل9ew@�88�]h�c�A�C���(��ϑ}�?�����?�o���W�,������|#�g�ӃNrI0͋��e�1������L���_�V�N�������������T��ɶ����R=A3ڽx�#&5l��ͮ}��yZ�%�/55vdU�Gt�X�</��&J��q�Z-8��A��"�aN	�3͠�G�2p���:y&p�[Y��&*��j;Y�t��'�:����/p�O����?��U�Ѿ����'�+0�Ga�ÁOu�]J��TuN[��َ$���!���kS"ceuE^�|%�+̟/ �q�T]�N�5��:�D�mS��v�t�:���@�ث��O}.�g�oU��x�B~�||�rU�u��f"��Rԇ� u�nl�k7O �1f3��w�WK(U�q���H��v�ve��k����C�&p���ʾu�ԃ2�b:�R���MekT��
���=ڑW�
ٽ�'��^���#YYAA͋k a�]�_����_P���6�gU���=����=�:c㒗��P���"�k�� ܳ���c>���e��i@��"~�e�� �?��þ�B��p&W��'脶L{3]���;C���`^��T*Y1664�\(���A ���A| �ҡ��~�2���J{���>+}>�,V��&[�`I@J��W�vn�m�G^�_�>��F���vR!K��g���ꚮ�)8#:?q��^��^�>@p6���۴�\ۿ�4�Z/Z�n�qne	�ςwf?:����5Jΰ���;����d�>�������`{@քr;���֯Y�:r���z.��V����h��`\ܿ��m��+Ejo��0m�C��eg�#`ߴȳ�{�R������;<䬽�VM(��D�-��&���~��y��Rq�*:�Y������׿%�<Q{�j?��*)��lb�eX��Y�e�fm�n_�{U��x�Al��W^�� d��jzZ0��gU�B\MGғ�ų���n�Ʋx$��ŊݓFC����K��m��W:;�T��"P�1g@�2`+��%�󮜞�d�5/�μ̭,ȗ_�F���o��d8���W���n�"�������&���b�=9h!���\^�nӉ���{�/����sg���/����/��Jp��pz����Ȱ��1�8�xz(�o~���,-����K9|<
���￐N�ݹV�z�����Z+3̪�ǻ��O  W$k�7׫�Y]X���M>��ZI#�Þ��3�3������J]8��P�B�qg���ӚlE�95�D�HY��|$;ί<�U����[��cȱr��Ro, �ųz�0��χ�58��Ŭ��l���>�i��>���i�sk��|��w���Gv���}y���_<#�V�
�&��2/��1o3- ���x%��>h������o~)����	>���?���?�{��o?.��x!z@�p4D��>���ѝ;��\^��yd-�u��ܼ��,���Ҹ�Ã#������4o�{/P�U;�����R�ҽ�C�<�Oᙷ3�Q������ ��g55�6q��FIs�6<9��xz����R;Y_�+���ϯ�`��kH�Vي�.6�9*nך�a,T"`xN����3Os�=�zːI�B<k|ϓ��d���E�d�;���#� � y�<��u� <@�n�hTFp|��( �.er�_�g+�~=���aܺDnmg{��&j�&���� ���8��:�CHh�V�,j%WuvF�k���^�N����i�D,�皴6���}�R+ +�viq��L]�X���hBRd����|U�lmQk�c|}
6���^�N׳R�1k�q=���C�h��J"�.�p��������S<��vfkfp;��x�^l`8d�����?��Ԟ��	K��Z��%�/�4xα��H�y��[�=5�1�d�)��,���#H~>��p]	�2HO�<� oYh�9���ṭ���-����S�h3�o�i���t�����X�u:���,<�Xi�13[}"�|���SJ�`��sC���'����L���ς� �0��/[k�����7����BY�ss�ܯc���fcٖ U�L��ObyQ0�o�W�_7`_d�G�p�>Ɩ2s�fg0���l-��ls�x|�Ɔ5�X���
��� ��������^6��-ŸT��p,k�����qv��3k�6kޮ���K�����ݙ.���K$��:��Hv������(��~��rM(�����"�~U�`PY�f6[,>�6����<��,7���Jh2�3Q��K`�qmD^u�i�A���Z�|��S#����Pv�Τ���n����]X�;+�/~)�|�98�Sp��9���J��;����c��dk�5r�y�i�*�q||�����՟��\^�ܑO�~"�����׿�G��Io>8!p޲.���ʊAc���S��ۖã��ւS���������@�ώdo�
�C�$ᐐ$Ψ4��p���2������������5�iW�d����Pz���]BjM��xc�"[�5/Q��;���6>���Vu��W^e�5���al���.�Z$��D�}i�Fе���~�`3BC�`x��l(7}�}������Q1���X^�x)/_� �&�_��Le\��f�aL֡��O�LW�
�L_o�i^����*~��%�zU5��9���������d.lF����F�p�Nu>�_V�� l��ޑ�_�#�a�~lD�����B`�x��
F)��[p�w�����e1�ϡz>��� ��j �FS|�>hS6�AN<�T,fo�:���8��g���>v��뗲�{�{.��%���/�q؎�DI�ccݵ R�*_vUt�2��&��׽�{eX��K��Vf,&F$YE����j�,x����tgw/̱WZ`��
�aj{�z�R��8�L ��~� ��@��feV��:�y�Q�<�]�u<T�����+ �
Pm�E�:\CҹS}|t$g'��}}m���h �Uz��pf!z1_]
�lf�|]��SKʖJT���?g��=���:�ι����� �����Νu�,�)?`}���[����s��poZ��G�l��)ѣf0�ֲ�H�x1���5���$�/*�N�L�u�X�c �㘙�Z �@��,�]�*1��A0�H�]�*���)��{���Ս���� <�Y�,د�����O{d`�)��S[�v�ϵ�{t�Y�0�-���\�^�ϫ�ǧ�]|?���������z����&|�y./�������+��e �۵U鄅�x��tn�W�9��~����]Y_]g�?̝b<�Wq�����pM(҅1�%`u��o}꺌�t&E�*ث*�Qg9��3�� �"+/��S��4H�,y�]���䕜`.���	~Lg����u�Y��r���j�����[�H�Q*5U�1�рXS*�-13��ya^��bf�T"VĔk�������-mY�N{;�=��^V���n��߶o395�}�8{l�x�[��J���erJ�A,|��'�md��sF�H����E�銏���q|~p`�N}�*:��U�*�����68X`��+Me$J�_~�<y��l�׿{�l�p�������1�N6�_������|*O����k��/�����Zp������O���	��҂i��c �M8gpf��#��5g�m ������M�N�:R6\�E���ᡟi��*a>�h�4l03\T��a�ܩ!��h|�S���řE� !�\L���(j/WIį��f��be/2�� �+�������\�g\�8�&,����Z��W�4�?�	0�ɿ��;y��{��>y�I�:~�V�75���}xt$[��n��'PQ�����W_��T}^I@�\����'��e�o��o���+^����Y�����c>�Z'�!"h�$��oomY���R1V�9�s�ڹ�09����a@j���T8��&��q�GC�u�(`hl=0 ���_���-�Gs>w�©G��NC���5u"�QWOe�y0"e���؄Cә޴���ֶ��2��lw	�m��VW�Yc�������yȝTCc�G*�	��(�qP��i���M�@��y�Bx�{{����+`�������
�L8��<2�[m���������VWecsS666Y0��x�ج�2m�.M�tM4/��A�����{ k
�z{{���.�3�6�0{D��jL\�f��[F��	�
�a�0�E�:�_�Q��>2`�b������Uq�F�,յ0�0���clk��*������`�gЗ����{	�+��%�6�v�_�p��a/g���%�������Vn��I@��\�ꎎ��(� ��<�>*�6�I0�َ�M��gϟ3�������"P� D���22��r�n �x���G��f�21��ޡ߶w�9� �?x�U��p�B���I��l��'�5d�>��]`�s�Q����\~���x|ߧc�����,[��-�f%�58U"Kx��{�x��"Q�7�������v$����&��A���i�i<g>-pTϿ���~�;٥5�\�y/��u_ْ���W�Y{��f���Q�cMf�_��(�R�8�jj�v8��\�Y_��A�WqN��-�D�xO��=������Z�D���Ժ�,�Y����VMY�n�T�������R.�Ti�zM0��l��	�9�����ńDO������d��Ь�|��S0�����W#��a�G�(̅`�eCZ�?~(�h�<4�]�Ϝ�ҍ�!�!p������9^^Y����\z�-�����\1�:���D�,�}񳼴,����\���ښ<���|W^�z�8F��ɣGO�������$5Z�0�U�˪.p4"ë�����R8W2	dtj��*��&R�GG�j�4:?��eB��ʀ�����Ia��ZJ�8�嵁�FY�f�"M�S��z�u�����9�ms��p@9��5�k);:^�RG�>q!�V%�*K^�CgI�o+��?���h�BB���-�����H`Ԟ�k���e
t��Յ���X�t�v� \�D���L[wq���pFe�:� O`���s��9�i0��?`ځ�����h������(\G�Z��օɠD����0
@d$ L�l��/A?ޣ�q�k{uuMb�:a�P��H�~���@��3 Ȍ��μ��Tߛ�S����-UxފөA���1�qޢ�s�?#������8�3;9��g
p�r���������]����x���
F;��E�U�1�w̟<��[&��� W"��hmh"v���@����=	��`�"�f4𙰙��I\g1�oi���1�Ã����ݻܗ���\)+����X�=P$�lX�:J�������1l�A��o^���ρ�[�Zx *��)�ُ��M�x�� ������Ǐ��`}I
�7�s
lc̍�B�`^BR��QO?|6J1���k^�����7<�@�]51��'X��-��Bv�/��bد	�v{Q{ytx?f��� '�;�+@ǢP��"\�=�K� �
T��}x��b�a�%h/� _��HV���-	F��=(��ǽ?y�rA��+�ed��c��J�yf끭�'gYG*�P0X��E�+5h���`��Ӷ��2�xc��(��j!#X��4<�V�s���(T�9�٘��bz��Y/�n��e�[��J�&<�3�YM78gS^FA,�oj�ϩ���.�P/���w�v����E�=�rb�ʢ���[�h�7�!�3�mu�u�3f�"cY������X1��$�"Dd,w;$
0x{~�{x�))�wm������.n{�g�]�Jv�6�J��L�$��s��ڬ}|������6>5��Ԭ���X]$�4��J	S�E, �A��za�&��O��K_Ʋ�(���nk��
�g,_l�����w�K��G����2ƣ.�H0����YD|���Hu������'�<�����^p.��"\Y�����|������c���t�a,�	Z^^��Sѐ8<:�B!��K���rg���ϭ����-�B��5*�y�ea^��V_��|8��R���Ca,>$�8TW��%+D��P}��G��,?�RV����[1M)uNmU���ZK��RXh=�G��B�:S�Hb� �Y�@���k��s�I6<Y/藰R@�߉�~��m(`l�HR�zT��ؤ�Jز�Һ&dUx�� �-��|O�e����ӌ��5�7���� ^�����G���ky��5Ǒ��ø�d�F�F����0E�	��ґrlZ����Z��>< �X ��e��(�Ȓ�� ��p ����bCz4�����s�@q�n/��\WN�d�9��mtܜ�W�l�������Q2�kq�5Es�_JKs��Gt���0�E�?�2Dq/����6V� �3�j���#��i|��N5��qG�X_�}cib��<`R��ħ����Y�C� |-*���vww������N�����s��ϋ:E?a}���k؈y@w}y=̅�����?���wɐ��1�q_X�?�˨��<[���j����� ,ׂ����=
{)^ ��p��6F����Z��ހ�P����\; ȣd�����v�w\D�����%�
1��0<h����ٕ��}^�/���&>\z\�P��}���CY�ųa�9����*Jwx�@��f+�����#��nl�E\�ڀ5`�][[[�:��X�ч\;D�HU�����prv�i*�sL|E�������A,���9%��X����39@����rK+o��B0���N�Xg�7��[��@�Nq'�C�>zsm �`��B1W`��y�e�"�o�*����>�k�˵��,'8�~vvʵ���7�3NPP*g@��uX�0*��퇬�WX�o}��n�Κ��o�9.b�wl<��_QD���A�e�a�b���<��vܴ����X�O�2��p?-i+]�p����z�@SX{��>�,��~�8��lh�.{#e}� �ڬ���*�d�n�������b�ț���N�:� �ؿ�����)�0�U�l��f׾a�/FI�����Y���Ŭ��v��w��	�^�����Q�<N�dd�Wx/�x,1�NM;Ϭ�M��G�0Ny0n��酊���q��u����.',��Ayy�%���[���(�G'��8�t[D���	��n����)�Cy�B#V�?�>�|RvO��x�0b �(+��v����y[;���}��$cW��9�g^��m�?��hE0`�m��"H(L����fz�ݸv8�̡������@1��ȑ�yV���O�h�Qc�����w��{ ���P���X���d&���T�N[��M�K8�c2=3�1�� Se@	��HL��� ��������ɉ�y�����Y�0�6y2G�D�� @��ޢ�5
�g�f��g������Xz��ܻw� !�'\ O� ����. �����W�Ν{���#�ͣ�T�����(�+��?� �0*��6'Ϯq�"�9�;pf�SYY����-�_"[q0 `A��m`@��p�X�>���=
n*�7����d���)Y���!Ӿu�L�		$�m< pƾ�?�g-�^�A<�;�d w�>}J�Ϊ��1�Q>#�ap~�m��M��Nއ�K�`����^��W���� ` 4 ���@�^�n���L�(U@�A_\��;�m��a���)Yl���O!��֢1�+�2���s�dw9_
�����X�����:�I�%��c����-+<x��z�M��2]��m��!;���<�i1?�pز"���jr�e-�L|/��2^��\
e}m�����׌\�� #@�1�2���9R`�f^�3��p��u�w�X���T�/��e����+���f���D��k�	pW�=&+X�:�+�����Pu�M�z@�i�2�)��󼥅�U�b�k\��7�y[x��y=.lN'��8F9%�	�W�]�k�*�E�2�6k�i�T��Z��➛Y6Ʈf�H���"׽I��C���~���=-1�?G���6g,ޚ�N���ezɢ��:Z`Z��Y��Y{��ȴ��}����v%Y�4}d�����XEZ����-���Ҹ�$�י��<;�
t�x�/>��Ь�|ۇ����j�;��ɗE�ԃ��t�$��0���R
=�Gڡ�S5\���)C����Vp�����4��j�����LNN�m\)#X(��@���g�?��O��٫�����Ɔln>����y0�e��Gf�8s�K%U`�E嬢����ע�6��y���s��h������ij�moq���׌�kF+hY�z�4�4%�����(~δUG4%��,��j�c�EG�wC&���x��*�c:��p����:����@<	��a�A���<"JV��1y�o8�EI�T�ۖ2^Y���������L�)���H���%�rg�:��,[տm'cI���g@��+��Pr�g�)�vy�C~o8����LҖ��Ű.o)M�?�Y^�q� Ч`b75@��	 C�;;_(3Q*;�6T��(��d`a'�L#w@�c<V�}	fL��J��Y�=��Ѵ�r�`�ÁNd@��q,ӍE��H3:F�JA�JY�����1G�B���US^�&^hk
���uSp��L�F1����0#�����{{���2��E�Fy�Jl���F�܂c8@��"��%@V��	ַ;�
l��^�<e���������}��Y"�l@M��Q�:�����do�`���؋!�Af/�"53#�5s�Ab�+�^V�-�e32�F�A�X��]� /�cX�qN���-�Rm�W [��s���� 1u�3/@XE3����D��z��{����B��s�?Qmv��,c��8֏(b�*��^�%�g�����MJF�<�Q�X��x�y���S�Y-'���LC �l���:�k6�:���`3�nY��x����O�����,e���V�"�������`N��M�w�38��A9�4a�$د�<�H�5�U���1��l*���%E���`�J�@�d,��mi
��H�	�l(��.}&�5����`{"[Ԏ2��@�u;ڭ<���h>7�,_����E����]N�*��r�RLޢD�-�gm�>�vs���5[O����5�� k�	jX�~���c��f�󰏪����NK��Ӯ�v�����ڇ�	"k
d���of���%S&i� �?�q���*�<�m���Y_NNϨ�\ GZt0����ÇШ\�㓭��˃��K�3�bo��>���k�j��V0�	�u�,�����?�ի����+y��ap 7舟 ��t͂Z�m�G\ �]�D�QL�i�MGv]I������q�����ot��N�M����0I	�kz��?y�f_���e�ˊ���-�M�) �yfl�󚥗���	VN���@�"ުj�`��Ht��hA��#m��-鷆��<�wc��9�U���K��}y_M9Φ3w)8�����'�{9l0����{TV���{l�U?��\��YF#[Ag����E��P��B}���2�i��3ӏRF����sƊ�I��f�y��Rv	 ���C-b6 S�R��s{]�#o]���� � ���kBa+ >���N�h���Rڵ@��|@���s�� 8t�&%�,��'Vh
��Xӭ|�i��_�T@��k ���p� ����� +��m:O�.�ʰ�5�F ��X����sF�3J�uf���,��VW5i�����Ma�{�n?��ۊha>��������k��x��30���Ǧ����vK�)���Z�2�s~fyy���D�'�:&�����	V{�3��z�� -"�z�%ei|.v�oĀi�	�OiF�B���d/D
�:�P�if�k�M���ƹL�k]U�lJS��e�� �1�4����^�A�E;�l]��\�s	���Hy^_�S��KP(3����c�����7�+�&�1����;������&}iE����ȯ�$���� d`0fQ��ჇԄVF�n�1���a+�V��,MR�3;��L�	$&^AR__�l3T��b���3���!���+�>K�A���4��u}�� c�:Qw�<����Y	s�mL#2���\�/�#9W�����a�g���>̭3K��]�%�[���sa/�˳v��>�>�Y �|��G�X��} [v���>�Q�w^�z�[��\�pO����C�
��Y!��C�R�k0��pʌ_oQ�9S���^cV����yo�{�f�]�i \��_���	*�?e��.C����O��*���`?2�U���W���d��#m�g-�q�V;Is ����;�b�����<z�ҽ�y��2t��o��ܽ3�Օ;�	A�|$�VN@�'
~��N�ǀ��������ޗ�pL���Q0�N�ö�ؓ��՗,�����-D(T��7� ���	QQ�@ǋ�� s�d<	Ԡ�M��uZ�Ԩ��_[���W�)���hA�zy18�A��ُDu��I�)����@�"#r&������YhI����g���dYt��\B��)9�[���n�0�Y )@)﮺��8��oe+���=��TF��:�Ɨp��������`��*\�q���| 4 m��1�7���u�߶��ڊl\8�ٵ�k0��G���NIt�mޜ�_�-
��7�tӴn|���N���g�4jK#H� �e�:��
�@@O� H���*c;���sO8&X>,:~p�����q�����G&uX���x`�2p��T��98ؗݽ}yֻ�%��2ռ�;�{��6�{�n�m���E���5��uT���V0]h9�*��:���'Zd}�-k������F�����"ثNh�i����s4��,���a_Z!;�k�ʱ �R`�L]��?��e�^�jIo�t��e-�v���9h]����L_ut-Ѣcs�,�|�dh�x�!����6�,S0�XKhA럝s�ƚ�9Np|��.֦�b#\�P~6 ��^�_V&7�[����5-l �����u�� Ύ�F=���l�N�B�D���� �@�� �B�	�����#2��� �	��^�wbW$ϲy[��VU,Hy����@T�&�͙�t����{+
����Ε*>#�Ł `���fVb��2��4ä�2J��8�0�|.#�qʡ�k�IT ��g?o1��~
<�z�n�~f�����%b��;�uo"٣ý��jX`<onl�ܹ �W5I�����8��v��,��M�,c�#(�rg{��e�EC���]�ܦ\��̳6k�vkZ��r�	a�8%��W*��r�$���s�ߚ)<�8� �L�J3�Ų�l���Gn��v���}���r5-�\կŷ����nְ&�e��dd�����M�j�Pʚ�9���Ah]v�uy^��#Ҿ�
������B
;
	����t ����T-YY^��+��H�t��h�H{L]�= x�/�ap
OȎ�#��Gp˧��v�ho��;��h�W�@��$F\M�[�y��	�=`U3f����_�Lg���wK�L�3BS0Y�� �۝�-���f1� ����x���&��ز��c/�5��?��@��1�΅CY�E���c,`<���"�Ԟd6���������R��\�u��6 � ����i�(&�g �	�o���5(^�	`�:Ӓձa|����N�B�)��:|ƈ����^��Q�Y!�ب7bjk������$�s0p��ed�X$�wj��������9ې���?7V�^��T�Wp�2=+g��	㡴{� � Hx}Xhq1-���g���_��bm��1Y�^׾p���+�`z��'kk+}*2q���Ȟ+��t���p �g
0���G���<۪^_����b��g��}�0�G,\!�*���Sb���qI�.Y���ӓS>�$�$:�
�uM�<xQ�X�$����-�=LwowčB5)1+�6����r�۳x�5e57����JӚ�Qj@$�O���6}XJCI}��t��ieCf4�"d`�R�W�}�b�0�Ep[Y�mӣu�u�4�a�k�t
&�9g�:�99"�\Y���Оv<�a� P���e+x�"�g���@_7��m��g���訖R�h���-c�>4��1FF&��L0zUO�>��)@������=�
�b-����T����[��O��	؟����{��S3���`V�ǲ��8��u�
�fqߍ߮���V4�NU�����_�-ڶ�w5��=@�y�m��XK��0��V{�*�in���ʃ��y+ڗjC;��u��3m���k�c~!j�\���-������z4y�(-�vas��<2���0�Sz�V��,#A�.^��܂�(��$�UJ��lZ唉Wf����G�.�Z	�&�;�r3�'�q���3˼��Ge�uܯ�3����������˟��E�}���u�x���%qf3�b��|���:����ɘ5'��4쩏z��Zg��޶���G�粶��b@�[{��ّ/�Z ����}��>N� ���ٳ�­tY���Y\߱<��0�N0:�	j9[�88q���%3�3�b<�m��y[q�Jʊg�R����k[�$�����x�7�(��҅/��t���T�� (~���,��]���@��.��Q�l�����#��0�K5m͡-#q��u����6+I+��|+�Бu60��:�q�*��Ʋ�2��?�Es5S��3�<�{t����p/̗9:>![�L\7�/ FTc��Y��@��`Wv�J{V��	�@�J�V�X����Eu�y�w��\�c�n�T;O�w�y����b�`� ��	�� �����ʮ�C�H�j��|w�?��J�v{��D�_�O#w�^����i�8P^�����9Y����Rn���9��z���,�UX�Z�3:R6L�� ƼW#��x��5�+db��F4@̦cs.-!06$ �YX� ��j�G�궷zJ$Iދ��r�I+�~���iA��,��8T��-��w ��(C�`���
�ǰT�����H�
�*��@��q*�te���~D`c_�i@�C�������R	�7JO����ãC-�$U,P�Z�b�Ǆ�l��#e��Iw��ϰ��$����rhi�P���Q�ʮ5�4d0�N9�}l�N8��k�N�d�L��p���&E�����)�����Ж�O06�8��� ���P��q�bX�,�2�ɤ/,@7�:||�=�j#0�}	{W�$�D�qf�r�_��zsʜ���R�pc�d;�`Uz�A��7�Sm|��V�2�`��t�]�ie��@[�Sx/�����uS�E{�)r�V�T[9ϧ��W�$�6=���$.3+4�cU�����p�zA�*=�5�Bu�޲<��X��Y{�C>���loo1h�E4�;b}�y�+�{{����F��min7c��~?v�����̒k�1�_�zE�N��v�5,�漳�=k�v���UǬ�9`�h	~�v}S
���Y�n���2�|�O����|���l�*��ZfC�%3��*�z�>�v����e~�X��)N I@�کc����Us������Ύ��W����k)�zF�c2g��"����ӓc�j.,̑�v���ecsC�ml�PE ~�r�^#*�� �Qv`~���� ��b�1�J_D#��X������Bq��8�:.��|��ydM�����\t����m����tp]��L��D�q�4�[�*�5)K*^�ԛG�@�:����̊h-�y�����LQ[.�&��;z6t^�s̃0�+���ӑ�*�s,c���9�]ӒР
]�yު���p`�l��R��&����WK=k��4�}��!`��_Hf�
��h�<e� D�D����E� -L� 3S��˻�R �������2U �y������ka1�-�o����z�Pg1������I�Be���W�J�kN�������Xii�p\�b����
 O���Z �p~��.�|:��3���{`�u��2!�`Bj�"վ({r]3(7	~�VM��(��i� x< ����Յ�1�^P;:ݢ�&#�L&fH�\�b��/SZHQ켾FZ�1���?`HE&����+uZ�n��Ȋ�Tc��ƨ���Z�.�.721�0�P���P�o�ϋ��d�N�lX&�Ӈ�}6�p�5�;@�15�;��#\/�Uq����!�xd�`oǝ�����
^W-�Y�W�>}apƲ��(��g,z�ޤ���kc����B�g���3ֽ������0Wu�Ll��Ƕ�"\���Z�Y��3�b�ޥzb��p~Ge.�J���1������8�J��x/�m��:�ı�P�{ƴIm��i[����D@B��d����Li�ݥ~���Z�)�4}8U�����S�X�x��䅁����d�BQ �[�ڸ)��^/aG��Ӏ�����O�(��mo�ŴWVWd�`?fH�,�al��ӻ��2 �:�o�5�ܴ;�}�����������e�V�!s�9� hV����LlZ�:p��]���z�W�63���f Ь�ڭh\\kI*�6�g0�!�ܙ�V4���n�!$m#��˒d�&6e*QcHYĹ��~���[,��v���\�if�봢+��p�ѩ��^�'dx�߃10:aa/MuZ�M����[e������8BKrg���A��莥�3%L�J]��4J�>�#���Q\��`cU���%��@F����	@�.Hd�6�J���b�8����Ǹ�-sE�jZ�Y�`lx	�nmm��A�j8ob����E:x�8�d�)|�M@W�H9c*�����V�`ˊ������̾�$Z� @.Q��M��F7��̋]�u��ن�O�5W�ڔ�;�E�'����JS�s��r\�P�"���XX�3��4�z�2����4` ���z�����P���p�k!��@ءm�
��v=����s_0�V,O���a�뱔��`�'!�U�_��5��S��H��<��pM��y+�4K� -|}������9�f���S�2	�ɕ,����6
5-/s���G&�aR��L!][['K�C�3��`K��*���3�5p`z��d�b�`��:�����\�g���<lt�D��Z�����|/�r�J"�\uiձ�����R�@]g2�bC&�S��x�&�ص"=���$[�8�܁�J��%gZqM�5�q�]0�q�Oǫ�ٻ��FP��bAI�L���݁�z�E,ćWN�/���q�A`���3�c�ӂ�쓢0E�.��y�Q:Ă/�o٧E����蟟q�tv�uZv��<r� ���T�O�@��8.y���9��Z4�U�_� �(e�N-��d���[/$[��Pk�qm.�q�d�$5��
�^��S55;����N��9�E�\�k��v��b|aMAP�2&H���c �Y0�e��m�N�ߣf	��յ5�_�l|��������YF"S��J��Ҙ�$�ŹעVα^��%�c�W�S-�%�`�ns�(�h�s�����絀�����y�њu�J�+�M<I�`ɫ�R%^��3Ѵ �i�_UH�G���n�����ݤ����zE�(�h�<ؗ�����b���#=˘�~?���V��L߮��(m}�5���RZ��[�U2g�����`O� n��}����*/�^�0���U��xMr3���~Z�:I����U6�gm�nC���D�revxm��&O��W���-�ܦ���	��Ѱ[�y泓J�$M�I�|�3k?���e�o��V����Sp���'�� y�>Y=W� +���Jq���`b������N8��T�9>���2�'�J�t���R�Ey��+��O�/�(���e{�%o8Jm�*p	�c8�� OA�CS�O9�{�E��w`Η:�(����+98<&����bd�13�2i���&���*�nks֕�V�hϪM�G`yn�����$�XX*7��A_�o[��>,	 +�q�K���v(Y�5H�)p�E���M�d4He�@ {j9��O?�;wւ��B?���df��U�z��7	 (;��Rɓ<yMAnH��p�EKN��ig@ٵ�! 1VXqq�� �0ݰ�a�L Pˢư�0B Z�=27���A����D��[_��9� ���jVg��g�W�����F^�z�^���)��Y���VV`���7:����7���E�6�QV٦v
 	hyhq��x���ʪh��3
�EI��AnF�T��?.�"ƹs���	�
r;xESg}0|���X���[�O>yJ�4��0���2�6N�0�����=�Uw��:��%k:ջ�{�α��>��s�B��&�t*G-0��?,ρ�_ظǏ�+t�=tqeX�hT��E ߁N/���O֭��;^ �	������`�{4�0���� +-�i�|l���:G!$T��#���W���y��$�Ȩ3����vL���.�(6��_�&��kU���Y��n�fP�i@,��p��Wc���f�^�KW*ktzv��׼�A�D�4��g ]����L�����TAtw(��>.nϳ`��<�3�.�I�yϬ�&����lEg�otm�F��N��ɩ����d��=צ�u�����}0���Q�p��A��[c%��z@���Rg8��ݽ{�{5�$�{�I0�r��(��<�[�&��Hcc�3@�cc���nXRh݃ʎZ���3ccY�d-/�g�)�O��#pSi`�5o�5:���s�QP��s�	����|n齻	��!K[��� m�V��ƨG�:(�v�F�s%�g!��[�&���7�E��޽{�`��{�+�K��8��Ú�`cz{{�Y`�˞>}*�=b�E�![c�U��X�9�l^���E���I��3`=`;|D�[؛ u�b��+�}�k*`]���"ˇGJ�0�4�L���q�X����*Ӡ�l�ڬ}��P��(��d��z���)���k����`�)�N�ڃI�^Fٕ��4!��>D�~��Y6 i���o������.y5���d�`���33::�g�h49�"C�J��Jqe�Kd8;p�vw�){�ɬL�R^�|��Uy������#�|�)�6�ȸ���	F�qL��4��E���`���1��>�awg�i� ����DP.��2����X��xNP�S��Ҝ�2�H&��jHa��`�����]H���4�΀�}'���M:w���z� �%t�#Ӕ�c��Z8�2�Z��cj�`�R��h��
̑�Jf�^ �~��J0J�A-�U����kR��Dg�U����:�jfA�L˒jn)��|�B$99.��
�a~��Q�n@mߪQ@H�]���J����@����5��>hq/��~�8����ѯ�&@�A�H�̭J�gq_e9�3�Biy�w��߲t|+���p������յ��q����༑~��E�.�����0N�E� `� z�L�"nd-�*��ld8X]�U������#�p�����|A;>9�7[ -�Z�q�R@|�V�����/Kݞ��\>,�K��E+
��#�Ũ�Y��z�dV8M��f_<�GsZ�9 �� ��<�c��IU���Yu���DZ�k<v�M?�=��`�� <'�[���1*&lu�yO��9�
H1�px��!�_d��^���u��)^b_�G�{��e���}+�[>�>�1�Y}���q=`"Ñ�7��ô��hc�t��K�)d[��7��x^%��E�Ef� �) �=����S��O��d�/�d=�a(g�ڍq9/�G=�m��3���r��]�����	�1��	����R^ }Hd�-��-�]�/������r�]Y����{*�:��[
�!�'����0�F�}߳:Hv�����L��EY9#~�k�k�Nj<����Eg�/�W�ʝD]+��-�^�=���5~���5������*݆K�M�y��:Pr�X�5F���眵��&ٴ�����d�L���/ɷ�l����]�*�@���;�w����|�<e�^*�U>�ƵVE1?|k������'���jsD��9��Z��C�^�[5�b����D�sdQ+��NfY�\��D3^�y�Ӿ<|�0؋�a=kݨ�{����8EU�{��	+30K��d��Y�p��r�=ߗ�ߝ0-[��LFY�
�1-e�M�.��0�gQ:)`�z����k���Յ�S�y������P
c���hu�g/�d��I�,N/��TM��8ע,0���q��e>��$�v>�Cf o��ޗ��E:��c:T��/��������NV֖��Q'��O,B׎Կ��)hl��
&t��B5��88< s4�ZNw�x�)�A�ܾ�x�80� �xM쓤#.�3�����`�8� כG�8�EdYms���6�m�I
` Z�EjZ����`C1'��D�(��@r� ���<��h;�F�9�ے�&I�  e�{mmM<�/��sZك�bz_f�X!�]�I66#2٥p�G��'�L � ����Sp�E�@k�7�і����O�5���Z8��%g-����+#�N; �b�}t��Jd��1518 yK?)+,��������窷K��5���5Ң�1�t�yE�������x$y}}�ϕ���:����Ĉ0�OAd��kI���L$�V�3m��6�A��E�	���	X�{{�V8���A!?8t�� ��3`��)G
�H�~.�5�x��4�f�W�bl,Ֆ�\�E�hڔW�T��^^(��fX[�6�Y�a�S�
M�,NuQJ8���9o���|�h5m9'��
��)r����_`���y_%�.��aV#X�w0�0�10��onR_�g��'���vjƄ�����Z�w�m��`<u(c���='\s
��h�{h|gj$#3�1�y�Ĭqo��oLSo�����	�݈3�xc�9 �8�Q�ȵ�UEß�sY�L��o�2$u(�����h�"���1�E�>�@�G���-��&�|q]��"������7J-����� '���u�֨�t��&��ߩ�Z��3�Z��*�-�ç ���y�|މaR�d ��CU��r�S�R 1ԋFP%f��C�0o\�w��h�i%�$�k�~4���?���>!�e����~�����<����
�;S�p�̙�x�q��
� 5pFp���c�L�fr�Yfm�~D�x���ė�꽌r�t�uγz�g-	��an @�������~��'r����b�<0���!qB�_XuѵL�#�T���oQ�~�b��c~-.-�����vأT�˵�k}��~��D��^���_Ei�����I��s��L���l�ڬ}�V9Fa��:����O��YMx��#��m�����)�X���KPVy�{_�S�Db+7�_���o�Ȁew^/g-�f���Ӏ�*��"zq�1�Hl4�� Y.U<� l�g��3㬕��
�e�}���PN�Q~vz���>��+������L���/����o���#ÙNH8����wiHP{)�Gt� ���7��!b������ q�1�$�S�epR��\ɔ�7[/���g���+H]X�����]��x���o
�_!�4#+��H������:�H0Z\j��Ǐ9�={�j� ������E��L��u}'�>�]�]�0M��E�5
gV�A�U9\����EJ<x�`�=:9���Ԍ�B�<O���\N�ζ2�B?d�0#N�Y�[=c��+���em�,�C�N ��n���U���&5@����vz4�Yl�N{�HM�{�2�>d|E��Zm8"�R2�I�(�O�� E�2�%R���'#�h"%rN���aη�;F�	�j�m�`^��n)wB?̣�鳾y�����/�+Kd�!� �h�붂�2�<p��@U�23�(K����{���$P�A��ſx��}ِ�Pp���� UVW��i�UGۙ�ɟ�B
��;�8���8M�ߢ�5qY jqO����Oc�: ��  �R�0^+H�M
�ҙ�`�����@�%ӀY�	�w��e�(� W��lQ8�,J��1�w8R���`u�l�9���9+���X$��'����k]�|pt�m	�:�H?F�Z������ygځ8��`��A��
�����20pLl��J>�4����n�&#S�q�1��1ڑYP���	����;\�wǔ�2&vf̏�4%�"k���,�<J����b�����z�B�U�u�L]+���L�� 񑡄 9������q�W���
:�����cZ�	�Q^���y��N��}��x�8�񫗯dk{����@�V�	��jVrfA��̴����<����2e*��h�P5�]{\�������9%y��ƴFPq�
dQk�� [�(�4�:���]D�Q���m�����He{C�cц׆} c{��X_d�@��,͖���,&�K7w�4pd�����/�2*�o�& PYei��۳���mnqmO )b�bøĺ�$�����l2�ɋV����1�/l��`�`?¼�������d$W %a��,�����W�e9dS�F,���qS����p\ ��=�]��{5�:�jh
��dX�@v���ŋ�$�����!�[�`t��dm�5=�[\6���6k��9�s��
/��,�T�~!�e�_d�Fh��0�K-��/`.�ئ���U�˸�q	q�YӒx��n��[�>B`���n�J�Ip�jG�J�U^������"� _w0&���p��N���P`��^0t�����4j���p����?�;��/�޽UMu4�����%��ӧt4���E�Z�`�skk[<x�k�sz
 �������y�,k��[V'�ŋg����(��xd��$^�=t]�."1S�c�����X����.�p\��(�)
�#�@���x�4
e0ʄ}�q3���R� �V5S�Z�<�&�h7�	T���駔��k�x�זU��Ù%����m�O $@�h�c�1�k[.0p�I]�ʌ[|G>U4��4ÿ�e���<��+k����K�{�LJ �!F�W�j���jg�C��9�j�̳<�b^#>[\��#ŧ���?%�me�������*qa���rF�g�A�Q�t0	���������KY|"&#��A p"uZ6Ǝ�)/ڧ�n��Z��Y׹�BߴM������CI�$�Ts��䙕ū����p@n�'����������08� ��=�==͊W%�� n�O����KUڒ]�A��Q{��i�l",ICe��V;�_\h�[�\tt]��G�f�G�%����&[T��7j\j��v���ź �����4�<a(���ϡ�a����<���-i�(cV�NI�g���F��Y�SpMgN$�%��S-��(�j�*6�&݄1 �:2f���e�b��@A ~VTm!���Q�V�ye�R�'l}�^���w�i0�����ds��xoH �V4���4��qΫ�o�\�=g�nG
���M 4\`ڗ��2� �0�m�e�'�r>;~e6h����3z��%3n��6���-��A���U�<2��gYb$���y�ڵ��DkdP ��z�k-\�e��a-��ݔ�/@�3�!wS�Ck���&s�����u��yj6���Tk�sw�9�h�+Ⱥ^4������罞��8��͗��	[֋����AdU���i�BoBJ�J��� ���5��"{�;�a�J��*?��>���`�I|�hY�)Xy���a�T�i��9�9HY�ӛү�<0��m�l�<'�pJt�%��W�.�� �7�kp%g9�-&W�߳�\��|T��v�2���Q�Z�q��j��r�ڽ� �e2iA6"�[�}�Y���W���<΄(�۷��!��<_��ș\���<��erT��?�?Ĝ 탱�`��ᤥm����l��ى����S�"�4��.��\�U�O>�$�|���(�.�Q��y� �TN�9=_�{eﲽc��,���:Dظy?>b���+s �UX���~xrF�B���sz]n�?���}�ˏ���	�*7��GoX�(^����������>yr�2�|���c����&d���/^��bпܿ�G;�g��9<�T�7�#���g�'�y�oE�R@��\��i+p������p�Ӷ�Đ���ޭm�EC�O_�M\�YD��w���^`�y#�!E����	Y-h(i'ZQ7�Q	{��}� 3O;� Ć�C����aX�����gx�"!������|�����*�V��r���|�IWHA.a�<v67������h4`����_0�Q�i������7�=��r�/���S��3pU��	؍�M�<�p���N�gc�P�3���6 V�hg�a�->��GnV �ߚg
��B���^�@���^�f`��?��"XxX����w����g�`n�Uyh�"b � ����I�a,HU7�ŕ� ���5�{�s��-�/�/p��Tx��i�I!LM����	��2.���T�bi@�*S�*�:��T#�b5����@��}h�n�l󆯯E������fG�&��"�A
�U�m⚒iѿ�J��J�E�2�fa?�8+}�-q]x��
n���j冾����kpF��B�~H�T���[�����,gi/EG̼r �X�$���peB�0P��\ D;�
��5z���Lǽ1;&bo>��t$u�9]�%�)˶ó�\�{x���~Bo4�y���t���efȵ3�1��>oy�`�|5�#�5 )EE��6����n�p`z�\�ىq9�� '�C����}b��P>Ñ�f�7
}���6^�5 �l9(X�=,�BQna�7�눦�0��- �`�aNbL5��<�K�8(&y��]^����:-��h���@���ڮ4co���H_���M,�����h{��&+�� ��`���^
sl��#�:�͸���L�k�����Sa��'��K4�(j�D+���e�1��P�}�l ���]aз&QaK+[٥��v�H��~�9�^9�r�g�ׂ��s�Jɀx��6������r��+؛�H2�=�� |9	�G��z�v)>�d8J�f#09CH�#�� "�C�G����ۦc���,����W\t��-!b@&H�{����]m�k`�j4�le7i{����#��p��,%��;Ftb�7����+�BV�1��˙L"{�\���v�ӺX�%fjٵ���s["`9#����l��{�x��~����fv�?Jظ2`�ǂ�0*�����V��FN��r�rR:%�t���^�:�G?���=��ݽ{�A����/��=}��W��O~E����}�ѽ���o���]:P2�GHi,d0���H}����Q�Lf0�~����޻�E�z�>�yuD��*7Y�9u�o�OJGj���P&՛�I�����~��9=|��t46X�y�l'8� Ja!��;���кH�S�m�ls/c����Q���؂������6O��x��'��&}�ixp�L��6�ҦYн5�_i#����$�D5��U�fɓ��� C㋟|�A�Y׵���c�YF�q��ň��;��� lon���	��_�����5�uµ�4�gTn��u�U�N���84M9qz[�����kKZO�W�^{�D4�=��8
�)��[�&�0�h�,��ys$��V�S �����:0Ǚi�E����������3�f :��z�h�?f��Z��B�8fG+����)�vwO�sJ?(�6� �\�H�gl�z�t�a���Ԇ�qQ���d7�Y��k�G���cCt��]a1��-?_.���6eF3�t���9���U�m-��dJ�� �1S�D����E�u�Y�O�K ��)��16����
�g'�5 ��`�8���� �����T�Ap,0{��Q_��Q�M>T�?k�&e����J��ߵ4&��ز*`� �2�z[��q]}-�&lc0!%#� ���d�������T~���f
�c�o�8���I7 lR\c���Ϣ(B�NZ0�(�/DA|`( ��\η���ۿ�ϙ(����k����>}(�b�� $�v;h�q�Fc�:����I���Vf]�,>cM�wn�^��&��9+"���Wy�;wn�|γgϙ�|�ϳv�Xh){Ϟ��n);�tsh�N�����ym,��<sa��0V��������
M-瞏�<�T�{����Ղ��A0� t�E
F�)�M�i�U�$�B�T��
A>fU�<�eǂ< �܀c����pY�D��~P�I����H�=���t�q�<�4c-��Y`@/���<X梽�Y3诣�|�8���EfD�x)Xc?���{J���K���ﴲ���t�7�%oK���)�l�m{{��Q��A�W�y�����[m͜��ɇ�c�'���(��%4V���`4�/�5d	BJJ2?λ��7ks=̊~cn{��z��Y�_�Q�� �����dp�aMet$����ף�\�5�LrN@�g�y��4�6��"鱲��l̮iCb��꩓�C�χPyʜP�ٲ�}BH��0#t�Z1+�{��ׇ������}�l8M� �Q*�j?4K�����%�a�]x���	��M�5 4��K�d�rU�?�S�����J�~�N�D���2K���t���ȏx� ��ϟ����_3��_�����[��jw���"�(� /�~p��g:���*
��ʌ���9����E,N�p�M��l����辥/��}��oX+���Q^Ú��j���$᳝��	� iO��F��-��&H;�L�Y�$$36���uf�ޕ�M$�TT����&o�\��R�uaX�,Kz��o���\���Ç����g�}�)�����e�~�h���=���_~;2@����j�^��"R�lq���# }i��%������2�őA�g�8Gt��Ia�rLR0J�'����.3�R�2�$�8צ�j���@Ӆ�����&��۷��0�hL��lM)@P L6�k��C�����
�q� h)�y�͂e�<X�w��=�ޞ�2�Tm�#Lҗ�k����)����p"���3~m!E�:03]ؗ/_���F�ǩ�'���Эd#�.�V\�aS ���8�a���t�Kg�z�iQ/�Y$#�.�\@]~~D���r¶<<8d��(�bϬt�(sM`F'�Y�:�:++��C)M�-��A �>c�h��` N����`L��}֬�w��z��.$_�������O����Y!ˌ�s p��	����ں���H��=IA<�I�����������A���G�C�UJA2�6����t���N)������4HE.Ey�Ѡ���$�Lf�r�(� ��E'�~��s3��퇱�碱�-�W����T-ko�'$��S�2/_��\$n}=�c7f&i0��E�@�3��2YL���xN#f�F�� ~��G7� ��/��.����Z�ޛ,��u$�$��rH��l���׌5\Vp�	(��������� �s���}Rd63���d�,︯������q�Rw��ўXC���,��C�/Z�a�_��끁�D��X�f�o`>G�sp$i�(�aOjѕ�l1��vfN�s�3��e�ǝ�~��D6�9")#��H�;���}&s`�U��$����K�lԹн�v�����nжV�A��|n��q�βY0��/a�n�/p������𯭡2'���-p��$��wr�oġ��leMW��_�R�*�f�Cܧ9窟u��0tS��z��oS�H3�G�)�ٲ�R����_��7���5�-r�h;-�|1��|�����M�9��[.�'�����[��wFO��HO�>�ׯ?.����d)�?�g�~��_�����N?��OT��7�e�]D�_�zC�_�b����z����r�i��ǀ���'�������O�� I�|���O��?1 ���b�T%��&����8�3�^�^v�m�E]�B�Κ�|p��F.F��{�`�Q�D[l��ؼ�'��}��Z�B�'����i$��S�޾}�>��s��/~N�<y�ڙ�ݩ��1h��Ls�o�&/Y�䎶����&�9G�G�~��D��9�����8�ʸ͔e�R�^Z/�,�c3d�>�;㬂�������e�+W03FWESr��m~ XmugP�my8�`C�8�t���G�k��\���O� v�L��~���{h�;*��5�<����`�����M����'�"= ������7TiJ3 K|v��s @����X�� �빬o�&r�Y��X6Fm��~ؠ��Ep�s�h�s o�dl�XX[69�7�6�?��"�ߒ(�S%R�r.�� �a���Ϡ%�ȸm�%�� �wY� �hsA�v�6�ʻ�Jd���7��T�*4�$��-�-�Y,	@� �8��V�7Rm<��c �Tc��8x�kk´;���)��v�5T�X��P@�[���3l���r���$���/7��Wr�w�7��>˕���o��v:��c@�� +���˰4A����<�� LwZ���Ep!�	�]Y3�:���ǐE��0H 6���z�4�ը���yVrO䨻;d`T��ו�
�$\��H{(>���ͣG���0��GG���`�5�9�b�=��џ��a�g(��Ж�#A%k��abA���3P}U*P�Z�О63�f�e�Q&��Q�5Q��y-�"�k��a`�@u���Ǌ6���b�JJ�^$_�2�;�/��dB����f�Dֺ�(�g׸Mp�3$
i��S,�=n`���� V-��G��4�7���Ⴧ����D�5f��`re�[��.�ؿಾV��̽����20�&!0ɤ̉��B��P���P �]���^��?=�,+�1^׊s�ʤY9z_T����B`�vk�Iϟ>�W�_q�S��X�z������x�D[�qhk	���OO�(!�%�/s��wa���ݬ])��F���؁7"������"켯��>d��FވApH�A�����\��}����.�萰��&
Q�w���Y&��$_m���/˜�m
o� ]6 dC":X[;�&z�����p{���nә.�/_�������`tB/^}YnH����K?|����O����w7)o�	�舋b������w���|��;87��z����·Bd���/� ���q�0�ѝ�w||��N����P�i#�k���O���(_٤���ٙ2\��%L�0e,����.�yw,n��*$E���@�̰!��"� ��v�ӧ\��L�Bc"6��,��EET�uhU� �Y���av�������O��n��"=f��t�����h(y��[\hn�R�g�f����ͥ��hk�Unz;�w��Lz `�~�iy?1���!�F~�bO���Xm��i�wWS�=��Er�8��~�����={��� ��}EG���߸�$-����M.�W�0�F�6�xL��3�s�� +����sa)v�%]��O����'�K��!��{�}C�t]�b  \|��^�xV~g�<_�z�A/��lX���,��Oh4����:C���C�&o:��J���@c��^ �M���Y�����o����S�{�~G���@�u4U�U�K��8L�5r������q/϶[)>F��n�襍M�O�!����:g&{`��Q�iM�A��2��a��C+��е��Y #�_)�elׁ{��(7�w��ʕ}��Ⱥ����Q����u���+�5��rLfor�G���I98��HX��Ɂ��5��;,�P^�f�䚹1t`�iѸ^��9}��H�XU�b-&�ǐ�Z6����=��ڴnvq��q��"�y �s��r� ��,e�|oF_���Y�ԑ�l���c��wֵ�"@b��`_yMD�cŀq�o��DV�����c�*@x�d�'C!�$V'w�_������9�\�x���F�O��b\Įl�M.B%�����\�_�\���["���>\S���oh�B�o<Cc+��ʲG�oc.d`W(�5	xcK��{?d��F�#u:��W�u	d^M�F���ys������!{c�sy����tN�tLA�A����]�6!�/���|���]���q�ŀ[��lP�𕷷7K?�5˅�-}6�XP�ӑ�
[I�+k�$П�EBt���Å3:��}�/W<�eܑ�##n��@����`�r��b����Z�]M�	I�-̵����&E�1��9�(FA�ze+[��������4��יǊ!�c$_f�Y|U��,�y4)��(˹�jG��&��l_��Շl�w/]Y�,���<oX�dǔ#7�tԄ�`v�U����o q���;�k��U^@�a�v:���?|Wn&�ǧ�U~�Y�^F=�Sn���y�\.��T@�"j�8� �ׯ���~���P���ζ0�:�5�s�1k+����~�>��~���h{�g_*�3p��������-}��S���{ě�SM���R3#�5	�57��O,fAIC.�5Ou.p\��*�i��>�"h(c�` ����y�V�6'�*�,
P#��D!�p$��`�a�-��?����!k����hi+ؤ�@1��i
���� �M�s?�j�(��}2T�qPc�]^�:ݾ�Co_3����������BҟX��wfGBr����Ϊi�p���~������+(re�u�7�ʹd	�3��V��r� 6�7�2;M���!�b+lБ�U�R#%1/7? ��{����%E1�M�h~
S���_�|QH��)��sk��5f������ � ��ϜH�Dp�=e��*���L�ׅ��re�x`e`(X�`�՟���E����o��\�Q�!�1����L���J%��!���n�����D�-���|\(��~�c�`���\ic@Z���_Λ^���j�e�l��6� *en�	���Ђ������h(�8<NI�W?����`Mr��i�+#Ij𡐟B��)�w1���1��*R5��QHg�1�:��A[�-1c��C��(���@6��9�����F��	��:<�0[�y���&���;���_0ָ���t�}d�Z�HA[ �`���e,�@K�4\@�� V���yAs�"�vK@�["���9�|!�rڭ��"sA��8$2��B�&d����Vds�&�:��M��p?4������l�\�
�@�{wÊ�<�����"���ܒ�8�HE7)${����})�s��E! �cR(�����0�e��|Yd`+���u#��>'�V�����B z�s�Aԁ��X���K�kk�Cf�^���N����V��T�����neeO�<�+�|�/�2�/�,h�X��B֖��V�V��x�l���8�e��_i'Yn���nd��Ah@N )����}������4�Ι}m��+4D�S"�#Y�r����g���+[�ʮ�R�h����D ��B_3K5#[�1��o�qb\N��]"թ{!d!�U�
�Y���'�`QaJ+�����#k~�7,׀�Y�D9�gx��s�K�ԁ��uZ�D�8KSR&(3Y�HW���3^؝+�@V��?{ޥW�{���^n~o���?g}C9UF.�a]�0��B���o8���'�>��~6���%�8�޿S~r��D������o>�Ǐ�ѭ}L 
��sa�o�������?跿��'{��>�m�Ys�,��ƪ���h��߭	�
��4�$
�
��˦���� ;���>��lϞ?�B"oK'���40����_�����HG~\>#�v\��&�����H1 lMR4p���t{Ǡ �Ђ^Wa&���[:/��gO�.��9�*`�����c�%K�tꎤ1'ś ^��n��=-�9�;Cq͗�0�T+ˣ~'0� ��ͅ�PY虋,..DW�Ǥx�Z�roq<���� ����\'"�Ɯi@�GP}�3Q ˉv)��9՟ګ���p��/�4�!�c`��V��\dU(TI�>�J��EV���u:W3��s�s��8=)�L8*�}?�ܰ�pT����g0+Ù���{^�?c�2�u{����E��t�[�"3}k�]�7����;���>��enG�aR��+��X� %;�V,R�{��2-iѴ3�h ����p���g���V�M
]���P0Ċ�ZA�L�]���v@���sf��g�9m�~(�u�~d����%|y�U	V(3��������ƕ�S[,a�S~�ǖ2[��<��>������oEaCp�n%  �](�%�g?��"�)0�,Sy��@ x)$#�����y<�"���d��t����B��F]��r!D-p'�G-�E��A~ex\��8��q<'&c�3=l[/�~5[��d�|y ��n���E�9[es+�B��`�B����}�Y��2�A���m��F���!��B���Mnd�yem��xV�d|Ⱥ��(9홓00�#E%帱>Cڕ��_�L+�aS��� IN�`.8[�Q[��$8���+���J_��o�����R�Jq���y^-笵�e{��&�k2	����L\�m���n�+�L=��HP�{�k����|�����{z��9�	�	�_�r�
Hmk��$���n�̗(�3ۯ^��Vv��df�2����Ϋ������a�r%<ϙ2ee	�H����01�H�p"$�@�<�x̜K-ݯ�����k���T�Q�<��5FU68|�B��u��D�E<��F�9�o��-�[�u^��ڼi�����6�|C�@��Cu�<ߦ��}�ݽ�@փ�<�\XG� ��~�� ѷ��~���>�����G��{�c�eh.Cf�/���ܰ���m��-R�O�o�c�'��Tn,�����w�������N�G�=�;�8�8����Uؙ������W5�v%zn�sRu�"�>��N$��.b�?I�7_�ɴ���[���]#�a#�  ����� =�6�#-�f��L7��0nms�+lr����U�P'S�R"��2�-`ᵂu�ٞ��֝�b�"��O�d����xk�=lӫ�������?~�o����&��2��������?���Q���Z�;��ht&���C���+�`�?<���_�s����@����b��)i�L�$՘+�	�P�(X^�WۦԲP`�*A*H��u0�q}��8l�U#cm��p�n��v�78�G'
��g��l�0'@��a9����p�E�'���++�	����6�[�7!-����L -؈ X2��Ep�-ֻ�V��
�d��-�\�ט�F=I����e��������;�jqH%7��y��f[,Ǡ㴪�Z�A���2c�X;��B�ePva@3>�m�eQ��:�I�t����$ `m� k!��F�
��[9�ۚV��s��6m��'�`��m�Z��y 7�o'��I��s��X�*���=�\@�Eoq��V��Ha���ef�ؗ��1�#[�B���6.ߨ n ������������<)e�4ب��� ���$7����x5}ɏ�F�
�Bt�9H�Z��/�źfR+i���v�=�p�����ڒ>I
��y+�qD@\���X��Y�4KЗk-��3^��b���,����P�N�W@�Y�-)�81�������(^U�դ,pK3�>���g������Me`��!�=q�+0�CR���Sc=�����Y��`����n���w�Z���ڮ�3?N2~-�Y�7�w���X������q(E�O���$���vG2(��W.Z��P3�~7A/xc�)�w��>���];�CNk�d��O '@^�
S���ߓ��O���͵b���z�D���G*���]�<�����P?����SS��ʙ��x�t.K7�	A��͇���J�q՝AJn"k�))�eZTS����d9߼��5k�e	.��">e�r�fz�d�CJ#웽���t�Ʈ{�i���͖@*V�W>�GI���l�V_�i�핈��5 �U ʀ�*�W��G/!=��AK���SG��]ں��S����{�'tz�MS�)� ���r���%�S:);,  E%0�bo!o��k��t~�������谠{wB_|�9�$�� _�xE'��}���48[���6�Ν��'t�=�t]G}������_~C�������g������O���-���!�ߩ�V&/u`(���χ7�
x.`��6
m�~Rv[T�d&<���]�X�;�:?�w�������ԑ��g
�8.��j9���#�+�;$2lcɚʬ��D��Tm(9�|(,PӰ t-M.e8�8تE}:&Skz��`�U=N\[}2�1������-z�����{����w������d�ڦj�^�ȏր�-P���"Y��)������s:88b�"�E .K�{] ��b1�����zWi<[���ə�ߢG)��ϋF�s
f���>0@���Vl3�	�leF���!��{�n��e>��SH����{�N9g�� ��wk����\g��,�ޅ��BY[H�o��*�����;�̸�T�����ww��m%(R�e�����0�Y���z���`�e��Z��6V4",&��/���)}���30lϡ����F���9'H!E�~�q�L�V��n�և`��B�|�f^��W똴Lm�6��~V�#�]d��hE��7������p�x��� ~��a��kǺ�Mj�D���U;g�`��e>t�hIAg�������&�2�Qqɉ���M<^K��>HF�wH��?��\�tKH��T�A{)^�|�Γm8=�ͼ��z��*�@�e4��Yu�H�����%���&O�Q���U���j�ë�^ y�̰�7�͝2�j٭��dz��ծ�^QLr>o��T�g�h�T�o���Nw2�=|�]@ź&�%F`�l��G�΅|�˾>׽����8�@=t���f��?(Bf���\�aThUɞ3"_E�?P�ጽ˳�^�{��:8�huЈ��m&t~���#_���|T�:Wa�
{S�!��vB}���r �4�H �GJ���YN����U�-�b�/<�]@����Ķ���R�<��[fKa)�x��1��yX���]�	���ݜM ��+7"�1�&����.?�'��8���Hǎ
4���=fHEm�~xtF�'���:x����� ����V~�c�x�by`���u_�xI�~�]��&�/�0��R8��Q�$<��	k7��m�X�a��\��}u�������?����?�#�z��{�ѓ�,�NR�,�Zd*D�l����"�0�(�����u��)�ve��2q�8,�.>�N}�e��:�� ��?2K-I�M���ј1�8h��,ed��&� '�0�GЧ�q|T��_�����}f����~��o� C�*�0cı֯�=u:�<��~��%={���16~���].���x��1��L������N���6����jכ:v������'�s0J�ʓY�U�k�$-L��69`�Q��z`a��W�s{����=��7�k��`.0lI%t��@_h�B� `��f87� �i�<Hl�F@3�Q$b<Ȑ�ώ$�
bi17)����/�pg��%r�r�3���H�w j�Nj
���'���\�ߖ���N�T[�b��C.���>�h��1��1�)�O[�R�}:���ԨP'2n�5�0���ea6��<k�b�J��c�����h���Q�nj����T�e���H6a�±ǟQ}�*�)'�}� �/jW�R-�Zx]f��� '6���'��.�ː	?gT�Nw���gy��;��S��@&]�l w �m�<���dٙu2���	����t�)1���fy�H��*/�Yq���$��>�Ik�X���X}ke��n�2e�uMK�ń�v+�%��^���,KPꖈ޺d-j& i��nn_&WL���r�8?�5���w�&ly�Xvi�UG��?�����6�8n�ɸ�E��K�0�e8�[t����R�	;��^��z}T"2��;;�ã״�'�_��W�j��a� ��޼=v_���FA���%�t�[�7h�\�ր}���[n�O>y@��>����ҏ���)��w��o��?���������ߓ��/>��?��?k����b�KAB"�٠��*|YK���KR�5XCZX�/%�T��
gY�&���p���b��ǋ����k�Ƣݠ0Id� @���?�|� �7��t޻���G�S+l|���B�{9�x����X6  �� ����~��Gz��5��8�惇�4k���jT5�_ö+ �^�1���S��9���p� `,30;w�z.vV�hh_'o S��>��{�:�6�s\���E���9fU�}c�dKk��F�A�|���ؘ��g\2��V.���|��{���O��+�م"y��Ãs�kݹ,)vWM�7]�e^I|�@�:{��	�%_�� �y�:��w.�B���͵��օ[4�#3��s�M�gu�l̰�N�"W�f6�N@�9/#\��RFO�ۓ�Y��e9J�qQo�~}��躱���c�6��qnkH�(�U�=��x�~����-�=��rLO4_s�le��N����U���c\���F_�v�:ڢa�L�aQ��`3�hg{;�3����F)d9c��>{��n���M ź[B.��QvD�[��y��m)�*���&I�<If2%��	J(XY��[f�����J0?]�� ݛ;?u]3��&�ʽIp1��"��*�&�����K��n 9�X�G4)N!�Y=�ΛulIK�3*g�寽g��w�ǯ�ځe���Ҝ>�ܘi���qa1P:����.3lM��^�D��z��>�ކN���R�aa?���c�v����-��RѮM��=)�Vy�����!�v���M;�(�ӣ�Ͽ��~7,���Ϙ���?E�^�)�uz��]��/�(��]�ӟ������,������_��5m�o������%ݽ=Pt]s4EBk��R
�V�-����Kf}S$E��O��,:���f��E���,H��׿fVė_��~��{:>9dP��?.���M) �t�^�����-�������<t���}��}�駴���V�ԋ p��lg��Б�8(�3s0��tt�A�/9v���: �;���8<EԚ
?����͎�ؤ`���ot\ �$�%ښ>h�Fɍj?Fq����vU*z�ɚF���^�7]o�cڧX������(�`�5���ɂN�2Y��k������W����$�ᒯU�{��ڌko������_�T���?� �����ѽ$�����7u�چk��_�����ʦ�M��Z���ֵ�5�qO���c���4���k�ؖ�@�ڦw.�ł�=��m}��Gv�����Yt���1O\�ԵLsq�2�Ws9y�#k
�_[�Dj*�� x(tY�����p �������~��B�Z��t�9cF|���{5����fGZpw��هi�W��e��ǝ��9�\��7x����T�1	����'��K�C7�_�dX&ߵ}t��wq�8�>���5��YB��~3S���[?�Z]��v�
�pu��c[�)܄5_�Ha,�����n�w�P�؇�|���X}��X
v�igmʆ�73��*�h0(XK���қ�o諯��LCD��m����������~N����h�B��'�0����|J�"��2�ai�9����������_�~Eo�t�֭}����O~�yy�w�[��ɱ������%r��&`��nciRM��l���+D)M1a�����81��W�^��~�;z��=xp�<��EH68Ő4q�tZ~���f��$c w���[z��%�~�t�e\��|��mV�8I���g+��\�L�ͅ9�^#����3�:�ME�mb�7ݼ4;)1��b��d����:=%�׽��t�#J����O���U�M4��W��=#튫�5����+�l��\�fZf��T��9ZX��0g>y��\3���,"1���D���Kwa���/,i��</nk��U[�9K}�	���K�)J���E����i�-(�� *�٫6��0Ȩ�*����OgT]��:�>��˽�;���-�2z����K^4���h ���2��������c��5�Ljb��L.AwK��ה��:/pE��r�𞱓3e(��V���>X������A,`�A'Eύ��a��*9�{����d�(����SK�u���J�{|*����8[��A��-K�/jl��^t?x�D��V`�8$��K�t�[��tKN�.�7# jǰ-�5-���
2N�^��*_)���F&C�v�����`H���C:��ӧH��S�{D��YHk����}�l�紵�����3:<8a�,��kmnm��K_��?,���_���W�������!׷�裏>���I��������i�T����@cp�g5�,y���5:(��j�>?�:�mX�N����m��	�D)OZ�U�D�L�0�ي��i`�[qɿn�G�+�[����6�KG�.�t�������k1��5R��j�{��J�>qx�X�Hf�`d$P����:ro���rS޾�π�Ç�, �(�+R����b���Xa{�zV��r>0�&<J1���:�+1�R$,"���B�[g@��`��`M�1W��CzW�P��T܇�lA��ϼ��� �����{H�f�f���}�Y�5��.\8Ϭ����-/W�v�s�k|��!��l��=/Șz�a�Q���h��5�8[xJs���ޕN}���خ���w���i�w�7ncc�\��i���נw���t]K�BYd���X��\���|��IVj��#�Tm;�����L}K���fЉՊxm
&Q�|vm�5V�W�	i����T+[ٵ�ql���c�}�]�H���<e+|!�����K���0�cf�9�W�a��:圙��%Ɋ�k����9	{h9a�@����wήX��J;u�B�ϥ�ч�ߙ��cOM;eu�]��ί�a�U4]�w66��;�ot�����ߖ��_;�V{��'�κ����N������tttJá�bX�)<����~�m�����wv�E����jww��67�￢������������[��<��o~F���c�կMw��Pg����k�|�`��ZyF1�w���p�9F]�VR��)*��E�,s	�{��.�Q��U>D��M<m�P�1�A��L�k��mC��c7kO�1J*i���>G\`<���X.��_p�G�З_~IϞ?+��w����Z�R�r����!��`�[�X �~��%�� ؂�s`�c,�(�G��O���{�h{g�+yC7�����0�p��(���5ko�V�%a\:ݰT��xx?��C|�te�L�<VR����W�%���j�/}�2�N�_������Oz��ܱ�������
���������p��u�˾�E�w��#Ki�8�	���sY�i�B��eٮ۫O1aQ�+��$Mh��
|��|�}���P�k�+@*Z�	/����-�$��	k��q,&>�xVU���g�*��.kPxa/�� o����H\ ����nz�3�ϕ����d_n���E�fZ��j��8T�c,�薂��:@�����9e- ,��0��X OI^>�x���T�lL;y�=ƹxe�݀�2Y��~{��+��7����W����*N�t ��5mgw��r��gmz��E/������zC��i8Xg0�͛�\4+s9�-�������C�����ݢ��BR�������9;;ӈ;
N�-�{�����}��t����'у'��9����^\��e��_Zj����itL�E!ڮ��ځmR�Ai�y��}���Xٔ8���"��ߩ��O�v�|�\`���ASC�Kf�.�&��+ �D0}�j�����R6��[�怒���{�s�6���=~���?.����e���>�E�ڒ�X� A�7����*[��?�hss��f���>i��b1��~��9x��a馅��0��f�1d'�Y�SY����j�p~Wy�4v��sr�´�zO����^"�⌖f��+�9�v�
��w6�S7���Q���\ق@Z�'�p�Ztt�/���#B���)߼���yZ����'Yo������yG�����1��/
yy�jnS�	���i
�6��uߩ�w�}`h�%v�&���c��)�f��j�X�{baގ}]n���6r�76mL�g]�y��yʒ+t����/�aT�z:�9eQ&Q������h.;#-����W%��{8.*�d(���d2B���*ȿ�w�nDcم!1��뺼�X��د׶ʀLV�����D��:k��w���6�������|qL'G]�z�uO���wˁ�a��l0�ç���IU����P׊Edk�ʷyb3����D2�����\ι��G�?��>���<�G����E��/�Q���)�On�9�",Cਨy���#�vS������.:~%DG4��S���}�kHA�\��/��1��1�w��@�9�r��˳���jϖc��Vw_nrD�����@���� �����k�(����nٷOT>>�~�j�g(���Ӱݖ"n�N�����Qp?���["����� 5�;����2
�F [']ur?��CGp���4岚~9�K��=7Mg
:X�!_�3���R�#|�i��ܯJ@����|Q	��̆<��r8�S�����Io̶�h��hf�L�m�-]���s�d�)alcL�ݨ��/�k{ݨ�y�rއyv-��j`��&���iI��U?��73���rw�Ԛ�Թ��3 �˰��-a�K�媬��A�9��&�8�����:����$s��g�ɋ�k+[ٲX}��&�8ٓM��[�k��)����:iە2Y�,ş���t�Y�����X��?��Sqg� ;�p�;^ �-�Ͽ��v��r
�-���������!��P6�%��.LL j�*�vO���s����imw���ߦ����勗���:zSP�r�Z��Yo@����O��;����#Gǧ��C�Ҝ:�ufC }Tx��}Kؙ�wh{g�v�v�ރ�t�<�ݻw���*�أ�;����#7,�u�ײ+�����rx�̥��/ ܲ��klc�JxT{���W?	H�T�64�[�k�63��L����M�Q+'�U�ho�u�n���Y�#H\���w�TD�U�!�@��W�dȏ����9��f�1��Sl�z`C��n��w |!�ﮯ��g�}�@0��|f��Ϙ���
ڡ�ns;���6wh}c#0�������	�Ȇ��p��\.�|�k2����0�k��M��~"�8�(E�<Mڑ���λ��A��2$}��DG,�I:u|��Y������rm��l�,���dr�11�Z���ׯ\�0+�X�m�.׽��-W���Z�2����k��7j.i��L.kl�Zv�c��'yS�m�CD�}�l^�M��/�Ipm�H�/��c�l5��샳����*2��nM:yM��di���:�J4�,HA*H�=?�9���"��KQf92�[LH%r�s���}�Аa�ev,k���VS�ĭ��w�n��Y��m��^���5[���u�����z����c�fܘ�i���yL��ͭ-z����lѽ�w�͋�9a��w:�~R7�����8���X*#�Z<p۝mll2Cs�<ޭ�[�{k�vw����Sg���7
���� 96a�mI�+���|�Zt��5�V�r���k�k������I��
�KdnDg�3>>���P'�0��D��I}�`4&~ �g�>�4��k�(
�$���fF.�֮�0����m�[�����`����]����C�>����ܤv�G�ʄ?/)Y�iq��Rm�R�q�giQ>Y�:kj��� ����P�,�`%�Z����TA���{��A�x޻H@!/ �&w^?o-$��W|�s�m�{�`�K`@G����O���y�"�iZx�~���&�	��}:����`�dO8���W~���f������'�X8ץ^���N��dL�e��f�\�t��֛�O�?W�n��M�렭!UWjA�����4��,�@�u�˼�[�B�>�
j3w�𦦪Y��u=���p��K��&��fcҁ�uf:��\����,���&����3��H`3Vr�<N>����|(�%<&��e�-f�g�4I�A�؆�{=�c֔�Z����e@�Ȟkǘ���*l�u�
3OS|u��Tu�
�D�;�0� �M�����swT����}sR�����z�R��A�yH������5��`[BKvs{�n��3����F��wh{{�%7Ά=��J=힖ΐ�9�$%"�I��~:x6����\�U���e��n����?�8���~m���]t���!Q�x�Bq�^�޼}K�G����3�K>FQ0�;�M�r�-_�I��O�����m��isc��ݿ�Z���u���_p �ǻ��e�W�M�ϻ�/ SQ��֭[|͸�ׯ^���q�i?|�}��A�4m��hX��(��G��3�:����uR�$kg���ɯ��,��Y�2.���[I� ��E?�xѦA�t\�r�sw����P�=%�|�d_�!s�ԽH��ɨ0d��tՉ�\�*��Mh[~/�o�g=|M��.[�aQ���2��3�^����2�����I�TȜ��˵�8���0�\�í0V�s=�6o�\�x�����Ma��ms+����IV�}]}�@��G���<�����v�b��ZJ��]��jϛ$\4�ᚼ���Լ�喇%�O��V԰lΙq��p�˨8����v���B氛 ^���XyGM1�z]�%﯆�H�>��0��z5�%��a��,(d��g��UT�X�-V�l�ʅ�1�|��ͺ�L��Ht��[��Mu�b6߰-��7 ����|�,�pH����`aMM2G] j
y&��@r�*��4��rѵ)��ߠ��5z�x�g}����!1;`b�| `����:����?��Z�M`���NDD��5�U+q������#��� }������oohj���<dz�=@�Y�&횺�E�^��_ä�w>�$���2I���r��kC�ߗ/�r!F|a��7��G�8�|���t����'����i+��#�}{@�����w�ˌ󝝝�g�%O�ҋ�/Y�_~���h{k�N�����tr|�����.��ḡ~��uy�������5J�e���c@r��	��2��Ç.��۹r�>�`�ĲG��I�S��8�~�~��YؿlܫD��48A"!Ac����k�>ߜ�ą7��2�+�����=����;���9&��Y�ߘӮ�lu(�ys[�1���Y�9,�`�*d.X�單�8,�me)|�מ�L��a�
�c�z��p3�+ z��ʓ�W2����3��S|��}aY�e�+�{��'�b!#(�0�չ�t㻓���Ë����EfY�-���h]1�.��-�/�K�@�y�t<��i�ǍT1-�����^��V�.�����z���T����T�S�$��3��:[�{x�5�F��5��D2'Q���fa$2-%����������&=��"�W�)�7Wg_��u32.�ӹɯ�AlQ��#�flf���  �B&�V9��mG������	˹��h);v� G����Lt̖e�P}�,W���A'��ć�R��)o���7�j�7?,fk���up�&mԯdί�꧎�f�SFa9�� �=�b�1p�������-?3Ȟ�~���_|���B�#|����).�h*�X�Y��-NON��蘎���yC;)��>�ޡQ��LSi ���9M���X�3�>93���?�	���1����*�{ڹ��?��������}vk�C��Ip�b�u��gH�9��9�c%{�q]q<;�g�������6�r?h��R$�\�����)�!|
��Wd��!ĳ����A`q����������.0eѽD���&�]e���^�7�g���=?�<��䬂ɵ^vI��	�~�7�ٴ���7��7�i�+�5�������¼*TC���K����P�����Mj1�`�Opcõ)��~�a���{ޗ�-�K2�Wv�aqGQ1��p�͈Oɞ,�g��
���"dV����Te?k ����'����
%(��ܶ[��7���b7#�1q杵�M��9m��9u�Fpa�D������0hā"'�&)�qq�H�kǶ�"�0,�4�gA�w��5�hx��D�Z[���G���X�MP �^e����S�"ad�3`@�IQ:������wv�e�p�g�ׯ_�3�����?��NG���t �Q|o02c��tq�u�Ѯ��� ����1x� �86��!�1������a��&���.�˕�Ȣ��R�v3~aH��_����.M/j��s�Mr�&��ů h�gÎ�y>�&�u�ωV��L&���l��M��M2Oɀ]R[����n����u�9�	3ȓ�Kr��v��֛��Z�G��a?��fW�Z���0��lok��&рI@�U���KV�Uؒ���,O��J����H�4���
-�����bә��+�ߌ01���]�-��>�4?�-�*�lY̛��_�A�ĝH�����o�%���L��ʮJ"����8)� ��B��y�!}9�Q,P�4���k �k��M�ѽ�3lj�)����3���\nte�ٜW�c������h�����寽@ʖt�"0�$�:y�v����2q�mT'�.�Q�,F�ݫ����eD�-�dY�Z7��4���G�v��A����3@Q�Ng�A�Ã��������p�����D�(���^2
�1X|xD���,_��tU?��=r�Fh�~�NN��Ɍ,,��	�z��׏�D�e5D��͟��6Rkn+m��">������Y����^�倇K���-�nT�jQ[���O��:[p�E���9Ɩ/��p��>i�B$�U��A�W��>eƔ/���.�k�I��: y�'�,�B6o����k]�����c��I]�) {;e�RU��������L_��&Wh��⇥̔�#�>���e�rL�{�%qS�_���6�����IKp��ɝ��N"�\7�{�([>��w�����W.�f��qe����m���~쵕��"fx�6��Ь��Ĭu����M�5�w��a!��JCE��I��8U)��w�ٷ����HaD���Nf0%�̱y�K���|���'9���ox���x�݆���	��,By��,d���"O�m\ �Γ1�&~�6�M�K��o������/�#��ו<���n��H���IV��Q Q9�p��t�!�&�f/�x���c�z�Y�\�og{��hNm/'l����h� ������Ψ�笝�f�ِ`f
���S�\��@�l��y���fS��0�q��"�"[����=�UM�k��.��Ǌ�ʫ�3}��R"a3/2��(*�}J ��M�SN"�'��3��0��Z����st��ܵ[@c�����m�u�C�N�^��Ú����;�`7�n̘�]��� ,��:�̑j�:ݍ��L�z�-z�S�O�~vޱ�x�j�����a�_��$��;,7�q��~��� &a�/A��k����ɶ�����	�b���vP?���{�B~R���)����Il>�-CqM5���=f�~_@d�r1��iƋI�Z�aϿ�e��X�������������K\����r��O	;QAI_$���0���p�c�f��w�|�X�����si�B���<��a�� p�ۥ�ɀ��}�F7Pت������}��`��3������ᡶ�g��W�T����'��|ppHk�|���S>�v�n��O]Z[[�͍�����Ǳ�,{�.Bi��j1GՈ�L�x�BV�Ȧ��*�c�eY���d6g�râ����~1k�"�3b����5��1��r���kge��Q����?b��O�p"�2���Wg�O(�	�q�[� ��8�U�t��Ϝ�*�|��v��m�3�G�b�Q��L���an�����[Mc�C��0�� -O��H��;3���������z+ׇ�w�5�?�����`��le�M����q7�����e1���)��1��Xf��Θ�h��xE�����&���"�j�5y+�h�)�v3�D��z\\@\ ^$�s�%�:�qp��*��4��s��!�x�
�S�0�.$�Ss�F����D���{Q��k+��� u�"�.���ߎUgE�pU���)��n^�X�JHKӻn<�#��v��og|W�v'����A����/������@��.6�gggZ�l��R��l �4���3X\�<��Z�/�Aj�0�1c�@��D:����N�������;EPݐ��j��e��a��s�����6�!�k�W~_��/�O�������3�������N��h�9�z�J���(�2Q��<K�tt�{e�����y��� Z�f沣 ��;�������l���5��#�����>�d�Ns.�/�_�����Z�j*�4ϱ]��+Z"�C���9�Rb, z�:P3g�iĻ�?�J�Η����������*����Y�-�)C*ʶpY���u����K@���d_sM n��k�&��\Pme����͟^��NQ��K@����
mZ�;n�yw͒|N���0�<:�-ҺO&�Q�����'�yo���@T�\�[�/�l	��d;Q$���{���+{��υ�a,+
���` �N���V��ƒƲ���)�V��6�`��	
c�@5���ζ?���1H��Xp08�AV~�s�+4"=�L/��eSݹ�ym�<v^�l�Muò�7��]���F�Ca>֦��� ���n�V9�ooo�ޭ[��u�̞-�F����0��,1
v��\�+��Z4.�^[_Z� �#�4�c���e0���>/���^\�=�Yh;�y60�<���L��M˴ ���<��1���1��3������Y���?i�'H6����k+;4 � ��*���
4ËQ`���Qo��H�b�a��b���E@*H%����߯К ���ܔ��6��	�,~$u��o7�����_�y�n����4?���"��v:�M�&b�)E�|����!�|��4M�N}���uq�8A.\��q���\}aޯ���\�M�g�"�V�/�?��6��Q�)�<�Ǻ9������\�H��7�S�
\^ٻn�L����1(,�A��Xt=ӌS�0�N�u�I�+#qG�Xr��%����gs�K����}m5��wsɿ��X��?�ǁ�g.����]c��\^̢���)�[�ӧn���s�q#c�u��c����W�!� �yX0^ 3��O�F2~,�1�58�lEN[[[�{�o�Ӄ��������_���)���h�E�b�dti0;<�G�gy�nWؚ�v��`~�o�s �!y�� ���CU�D�Z�`T���"�p�䃺GdN�Y񷔱��I~*
BV���"L�thV��{i�bZ�O�੟O����/����IQ	{&(���M��5�b)$H�׭Є�w���D�|Qv�-�.��֎����k�y6���|-c'�pr���;Y~�/�?X���8���E��U����	,�Of�"(�땰�e� ���h�׬���}�����[�e]��w^�G
�O� n�J�\�}��ɪ\�	 �X0J�S+�o!�<���u�JDZ����s�������D=��3��i�LMq^s�?vW�a/�`g�U\�o�I\z�HL���ˣ� PFv��\�u-�t�/�ɧ�k\��+�/�q ��v3�e�Z� ���E��U"�I�v�oDlS�F1�eH��q���Ts"���@�ks*O¦Pf�ݾ;�n������\q�Ɛ��o��,�����b4Pޖ@�V ����&m������j�j���<�d�Z��^�`�{_�zY~G��GǇtpp�R1�>,�nݢ��:���i�ouZ��9��B{`ޠ_^[���s��<d9p�! ��<7����B.�m�hX���w�x���ɚVٴ��80]���8X��H�c��\7�̒���n��bi�9��5)7���e:'Z0h�s�Ġ8%6�+zعL��)��M
�g/ϲ��2���Ց0��f2:Ϩ�jصck�׉4Ӌ��Q�t/I&��ӛ�U�?��K�٤��l���k�%f�����=M��7%�8}����d�T��I �O|��̚���<ca���\�4��'m����L���yO᲼��f�|�^w���j�^M `��n��TOs�<�w�j٧�qW�K����NT�~S����X�\h�ّv�4c*�wcE�g�.��3Hǯ!�����V�n����:��PÒ��U��rZi��VR��8.�:��ژ��<�d���,�~>�ą���sm`n#Z��ĮX�ڝ�<c`m�%���;;�/@"���bEY�eT����3�	�<���6���� �D�"]�ݽD��+���?�3������dv>������l��y8�����I���C{{w����y���1!`��}}}��g=n �o߼��Z�����ċ/��� ��F��g{]f*�xU�1��������|=�Ng�|m��w}m-�e,|���E�e��0���4`y��Vb�}2v�3�l^��x�"�1
p�R���U,�&��<�q��p�y�[� ȃ�_��H�����<&�y#%3c2��|���n��Pu#��?��9��,��������F�4�|`Ӈ�C?��d<\x��m�+*�Iםn�m$7�0�{�;��N/s60���BS�����ϥ��@]x��d�c6�E�����6��_	�p3�v`����ű��s�n����m=�_���f�r�)�����^߮ҟ���n,�i�G p���ת r�3��/�w#����շ:��2MH��i�~�~���LF��� ��Y�p��o��E��|�����j!E@��eZ�;j7�3���{BBNu԰?��?ܴ��`b���1v�!�;�e���>?�5u<�md���edef�,�JG��a(t�	Pv������U	 :+F&:�t� �Y#,��.2W�L0�w�vG��XЋ'�"ա�IvT0���u��lc���5'腾�_M�GW��V�-���6KVt:mf%�\� z��w��H
����[:==�~�67����Z1،K����I�=����.��^�K�� D�V��6����:��$�1��0[ד��x�bǺ[(� �\�-�Fzrυ2��Ƽ�1�2��ދ��y�C&���ݣ_�e����l%��%�^�QO��d��Tn1K~I��[��_/}ڑf ��s[�y�����:�qL�?9�v_e_�߰⒳��繺�4d�_5�t���M�\ܔ�)��>����-MN1@�RqeWm�j�X���51h"O����Q�lާs���o�kp��@M�ki��ͅ[_�Y߫�NUK��ԩ��~����׷���Ӥ�n���L��67������)4, =-C�J���}����z��aY6py��H2S��؏�9�uÅ��&��xO[e-�9�y�T� C�!��D��0����ח��@\�=M�g�1eZ�+[�e��v�,e�����E�! �H��\e/Zq�j:<��}��$+�0���E��~��w`	.�-ń}��>���}i�3��M��^�K�-�1R�W�K?�{�22y�~�ǉH��1g͇�'l>+�K�=js�Itq�d�8�Hth8�C��3�����~�x�ig8�O ^�2=f}����gX�XsUba��&��s"�ar�m�9�6�\�s^�-L�M�ڑ9����?P��6����p��2�f�wwo��t����!���R�bP�`Ft�@4���w�p���ޭ]˅�O'''���E��{�����F���:*�}|t��� �̋��缞.�p��O�Pګ�]/|YՁ���.�ɫ	�,�BWa���u."�dI/k��^�㓛�<��x��p�me��%�%u�D��]��m�>٢wó�5Z2	���p� ~����H���qI���,�2�w1;9��8%�+.�8%E�7]�9�U��9QNq/�M���X�ۦU�N�<G�^<�C�!j�};iF#�|�)l�y��8�l����h���ē�.i�����t�h�ٸ�f�����d�ئ�9�( ~$>����;�cB;��_���o[m~��-�q��c�UhQ��E(ZcT	��U��9Uf���XCV��,���HY���'��4a��ΘG^�R������ɹx3�c<k{��t�"�!�M�g��A;I��'����1�O���sj�;�!�A`�r�N���� �l)d_��3�'��Յ���/	L:Յ�TT�w�� ��m�9Y�V��ƴ	����]��񜉀��Ѱ6��@�3��v���a����.���o������AC;���>br2��~RF/6zxA��Xz(��kk�+����}�|�qp||R��}+���Ϛ����=أK�V��Zn��Ie�������c��~S��a ޣdwX����2���x�X���.x���k�2~?��[b�z��6����y|g�� a�C^8�
D���V-�3��9�� �=?g��r�*��%M�R�3y@���We1He���^[ �8V�Ob�U��g]��|�(�ӻHZ4��l�%,f���I>���Ѱg[��g�[��W��4�I5]R�r$��X����_��&������Y2zǮI�6�"���o8�O�V�D�Ac΃��#,7L����&��a`�E�N���(dC>x�r#����u��u`cW.�Y�P�2��"����P�����E����	��8i� ?�ukKiъ����~��j@$��g-

s�?��Xc�ߔg)B��=3�u��ne,s[(�,R��<&���Y� �rH����ac~���{��+vw��p��[���V>�v˟Sޘ߹}�͙�� �~[��{�cPy��F��9M�h?��f��Ac5��� L�Vs��!�q�]�]`}K�$��]���c�η%\Pts���W�� g�K��r7�YT��2�������'�~�e!3�ƛ�QXW�`=,�ֲ����6� �i�2�s�-z2׊�.
�h<�a�Ǧ���7�\K}gm}��\+$�r�s��\j|	��귓��~+�s[�:==Qg�s{A6���L٬RX�5n��bskz���� -�
$�����S6�\k�x�?$A�f��G�L�l�a�V����	h�{�������q�G�,H� �^�~��q�[<{�+ �c��Y"jMS,�V�É������㓓r=�뽘�����E&R��>m^�%�.>V*��U�3$�TG�#�� �����W�!��0�9(��Z n�� ��{7�W��2�d�q����v���N���zy���B6�0���~7�x�(@�@u���V�?�qs���6�6+`�o�1���z�����0N߾}��`�^~8u��m����N�O����7��e�����bh�%�t�OӀ���,�8v�(�Is�E7�š��hI|�c�Q� ғ�k_dꇓ ���c�F�
٭��K�e�u �Ϟ>/��1�]w:w��Юc�p���sz��9�s� �����|j���0en����JDYs��p���ߣ��X ��#d�:�7�_�?�P�yz<�� y[C6��ֵV�Y���X�SΓ���	{�Yn����w��{m��{�� ��H���?3m>ڇ����$\����I�qN i������N���>&�j 5d	���@1ɜa�a�G��c~���Bh�X_S��b�3X���Pyvwc�2��Ӯn6k�5��uCŀhAՑ_� t��g�K�LU��3����#�;M��dMX[���׎��l�ʟ�/�C]��k�!��ǃ]mG[����E�;뼨�=_\���Ѐ� �K$�6��� �c�lW�N�*@3ɦ`i���4� ���t�OZ�'.����b}[�;�I6,al�JȢ�{{�����n��z����{��8�$K��=.�7	�ɬsze�t�����۷e�{�kgGV�++�x� qG"����SUs�@�"�$��B��s;T�>}Z�5$Nl�$6Zd�C�)-m���M&�Ç�׼���1�9�(��G������0N .�1�H�\�g^��0�[�0w���ۍ����Ǜ[_S����H�R��፳��{��5�0�l"����E�kE-W��M '��Pb}ú��ڃ��Ȱ �=P�?�3�`������^�5,H�F��q��0�Nj2T�s>0�c8и�4�p������5�j��K��(���7�'�'�ݻ����6|`�8�����H�q���/e
\��}8poy���,ľ���S��>���&cQ�ma@����0�| �׸.�K��z��.����������qk����0���ﹷo�Ҏ�T`�@W��n�{��ʲ[�qss���Q����5+.u^����W�˃>/�os߭�էٍ86A��?������fx�;���<VI���3����7 dQ�;�h��#] h�	 fq~
�3�݁�#d)�[ab��x�rK�#�7�����C��ȴ3��;��)v��	����p\[�W$އ������a\ ��<<�G�q�p])���|���]���7m)�6~�-Yf]����J�����ȴ=5SD�0����a_Vs��l���!�@����E�d�X/�ޫ>u�0i����a!�:�s	�th���k�Xw�� s��т���T7��qد�f!8w!�y�-�E�Z�������nsA@�YX?��̢p������am����k�}΃{8>>a}��,�L�V�	����d6k6��`�`��iY������5�f��:��"ag޾�vݓ�����uj`��{-�Y)�k��}�_z4��0Kf��
� 8�~�[��9&�!Ǟ�j����2����=r�����W����N׵�m��"2��_D�>[�q,,V��rmh�t.��&�����	"�4�!� ��X$��7�����*n�tj����Z�N��^7lڭ�ho���`����1��uZ�	�,p���u�)N���{7Sc+ަ~���z��bÔ'�6�J�����j>�3�i��~�#2Qh�(�L@�}�����"��
���0�� �3�� �����Զ�oT�c�e�Ͳ�A8�8�9?"C�	� �3�
�-��3w����(�����r'����W�I߱�.�Z�!2%RƨI���M ?p��:�6�;]�lGٝ�jN�΍lR�o � ���<���.�Up�j���:�`O���&�����$Q��K`ɾ��_��Y~ xù��ߗ5�*#X�{XYYf��ROԘ��F3V6��p��< h/��ҝ�g-{G���lK��J�����4'6@��L�����x~x���@S�ۉ��~V�JWT2�} |>�)�Tf+ӢtE�'�m u �.��𞱇���s5x�>��oa�3��"��Mq�RE�d_cl//T�&��5��*e�*@��d,n�C�-�t���F@\���]�O��tf�s`����ږo�4�-�!آ�2�������b���Jf%%1�I��R��sƳx~ogG�Z�"3�c��/��
�s8�a�K>| `��,)�i�P��kQj0r�"Xv�z4�p� X�#�����q���>fO����P��40q]�Df%�e�,q>4c�C����	3�Q�ŵA�����6ѿ����k�����M�Xv�ָ�x��1i��d>	SP�{���,C�_�}��_a/����8��eon�dX6}dm�
�G��������	M��֑�8W&Qr�'�Q��I)��GX�����\z��,��i�NX���[��_�H�)�:���~��2٩M᣼�� L�a��9=Q��1��o�]�}v�����Q�Zl�V 3s�֗��+IF�����+֝�%+�0�̶���i��ƾ���:7w����ŀ��wC���aV5�d�uW�_x�F�P��j�C!��R  �[��mN��Ó�Q�i�b�>
�>��$�<<u#�hZ1�Y��X�vy�斻�cW6���]���̭mT�����޻��[]_w�[[�98�&�R���h\ �OL/%v��^�)���X�5Y�e�L��6�~�V�	&�H�M��}ף3{Ѻ��!�kΘ� 0SK�����T6�(j♮"�Uo��*�R@eL{9`<�)�/��P��f��OM;�5��틵�����w�$���ӌf�
��ȭ(� gl��1�L�Om��֎�LY���d�fm�'�MP^<X�6��@io��?''���'���'O�:/}"�B�7�z�')���Vfz��!T ��7!Ł`�I �Mťh�0�u�?_K�l"�%2
�a�J�"װ#$�0��{�_,�d�1�Y� 4�)(��l�둏/��t�_�u�>>������������=4\���?�OH(P	i������=��y�<�9o�A������=��W8�]�͊#��uB[�5��0�����H�4q�sh�}8�X3mS�~�s����T]�Jk�gD�^�Ӂ|߼Ʉ�kL| �/߽}�?A������N�I#Vd1!�V���n��?��Op�RH%%��^c]�%~k��Wa��ؘ���{�7<O�\ɞ���7c��,���|��~��0�,�<`lc��}�1��v��������ފ����k����*��N��q���޻͍M����wnT�)!��6G�+icθ�}�-� �լ����Ay��S�EC��:���b�x�	&m�u��޽e��X�0?�1�O��e�f��5��L����9�Lv2�[�������o�FM&�����M�-aD
�}�5�V�l s�dFr��C$�x��dv�ӹ Ҕ�	�[to$
�Tgݲ<���|�!� ټ}7��;^��hu!b������c������0�8'ܗj���|:|W��X�T����֚�3c�4��asl��Q���ɧ��{�� ��ퟑ�0�)Cy�9����Ȳiab�F
0XSp
pN���?<s���?<
Fv�ﻝ��ܿ�뿺�^��}����Uǧ`��������dѰX���,�I����vgͧ�����v
�hd~���wMF]�b�����Kg�\l�D}�2~=--s1�y���j4��d�N���m޾�v�0Ԍ'�<8}0B��N )�c�4�.����ݓ3�R���>�%8�i�0@[0�.ޣ� ���Gh��A��勗������]/N�_p<8� �q���`�	镑y@,2�(�G��`v��[�%��́μ���7�=�M�jI�:��qtǙJ����g>����R5�G�xeDE���-��������V��1�~v59��� +�J�����߼!�f�e���M�� ���	�������ܕ��`�h�Շ�g����/w��pe�X�趍SLJ�B�D�7��\�h4伌Ϫ�L*5�%G��Y*.H��������E���ʺ����qg���I|v"��y���{���+�xh�v�x�k���9�c�y���<ǣ���3� ��i�v��.��ǚI-��A�޸v���9WmWd�=x�K�~]CBt`���MS�	#{��|���#Y�Yiz��7օ͍w��?>9�T ��Z�^�Nu�J��#�w���7��$q0_�^�y���8�ӌ�O8/�;ZE�u[�J��3ݛ�k�cLc�ZD��_~vK{KXN�S�t
����Y#�f�5���*�W���1��4��[}�
��eyi�YuV��&�8�����>F\��.�Uָ��2��$'w+P���=׹V;�5�rG�V@-/v�>s��w�,���s;�e��,1�-d�tvq�6�]��f_�!���l5g���b޾��ŀe�<ݖ*��k �M��2/���]��2-��TA���MQ���~0��f{�޿=tG�'d#�<�P�PNa�-���(�f;Z $WI�ng18�m����=��_���;����|�ح�.���o��ퟸw�=�΃����E\�.��dE�r,F�3����Ӽ��+�Z[,a�}�v�ѻiPbK�>��5���Rf�b5u�t�'�%�W�lm�y˫�PsO�'3+�O_ܯ��(j���b�w_�J*k��[V�c^�ƺL���Y�`.���v[�|�~�-:pW0�Y0l��:��꽲Dm�����ݭ�,[z�����8��Q���N*Y�5M�T��9�P�(Sp�^@N�3�ݫW��|�`�Z�P�^u�y�&-`��8��\�>�� u֗���؃��J};?����f�i]��,�#;_3Wi/�Yri��M_i�ހ��5C�G���9�����l2<Jf��[p����2��x5��h�9�´� N��@�l�<��-�� @7��uM�R�BnQ��f/�u1K��;	C6�;ᇇ;;��"Z��M��������{�I$ h�f��
�Z��*���2�8�sL��0��1 ���>�}iY�}����TMv�j�hQA7�?��~��ԥ��[Z\;���� F'�'n�=W����^�g����V�$/�m-]!��w�[��X���>uU�_|�� ��9��.���7;�z���Y��p���C�;.���g��h�`KR �G� ȃ��� 5b��,��M��_k���W~�_�݄S	�>b_�|�~|i�b�y+��*�˳�%ل�T�����u�iqlN���kb��
V9�!+P�d�ՀyjA�xʆ���1vm�1r�'d�X����xZ_����sy!G0q����Ŭɲ55-�ޝdv
��ւ�VP�t/���r��ҿ���7$ � ���m	;�˅��d���2o_IKkR}̷���^}�vD9M/� �%��.��,K�Y�^H|{*���\�7ƩI�5�����ټC@����{���{������X��Qؤ|˭,�@Ѻ���&�C�E�}�H)�_�a�N��ὰ�U�n{��[[�p�V/\F��¿˽%�����Y<rgG�����;�0t��������`ܯ3��lp�CR�*&l��ް�#X*Ϩ"�VU� T�F��Tcv�:��E����L��k� ���2Ƭ�����{������'c�]dCY�$#��koh}Y����&^qd���r97@Y��5�j4G#�z�`�9qx'ʬ@Eh+:�@v.a�:���ɵ�[E�����u��kn7}�_��|r��������h�3*�����y���h��N�K-�q3��u�R����#���]^^a��k�:<�Z߭���E�:�BJd��t<��:�`�Z�a �P��p\����5���ϸ��Q@�~�Au�E��ý�=�V�&�X�I �K�s;<׮,��޸�V�R�Ȥ��D�Z2�gx!����\rj{	��cY���`��`1${�͛7,	F/���o߹�ṁm
)����Q
�; H�tx��X�6�ht�	 /W�&f�x�Y�+ �z��b��=�/�C�Ab8�<6�[�g�禖��2�A���Խ}��66��5�������i0ޙ.=��_R�	cV�uW�?hDk��޸�E�m�6���\��pm3����5��y������W�WbAj�0������>x���||���kwZ�7��>�L��0/Q8� ɰcq-/_����*ط;;dp>�s0Oҩ*[h��c���^����=�<Za��	���p쓢�3Ʀ5���m�ɵ�U^��)��,ӮR�����w�.�}Emt�3�
�b|`��g���R��5~ᖲ�^�Q�1���tmm� ��<�Ҭ��!]��+i�P�&�sn
�^5�A��0&1߱6b^c/�8�\E&��N�ܭ��Á���v;�v�&�x uSi�&��Ka>�Z�K��]�+E���3)�'`m���Y%��/���7qː�@ �
��{��,�H>q��r��X$=P��9�
��7;���֋���ݷ�G��\,�Y8�gjY]g��ۼ�������f�r-�;!�&�((�~o߽{�޽~���Cwzr�|ava�^ꭆ�z������LD�.�S�Q����W��e:
���T�J �[j������s��ߗ�^�w����������-II��9�F42�]Q��c_Ǹv,��l�=MQD5
�x��$�pѿi0�3y�� g�ef�&�W���F<R���lUZU�kj��b�ۿzdsh1�`'|���C ( ��>%[�Cc�/cN�ql�0�]-�0:j��2~�P}s��SG;�@�����V�3O��L�j�1���L�7 `�`YX�����p��}w��.T]a2e�AE ����T �����/z�oW�K
���HX��egL$q�%`�k�� ���a�jF ��[ͦuq�(o��Fc�4�9�8�k.�S��E[L�2P�`��  �J
�>�<���mJK`}f 0��� N 3X���p�����>�ڎ�d.�a�\��c�AVekk+�c)�t����}��:g,5 0��@�\�rpP39�����c΅��� ���C�9�@Ҳo�p/��huX�9q��8 _؄o��k>��)�	�.�9 x��뇽�UF>��r�5? ����h'��	������j�Av0�wü�B~���H� {�����;����/j���ʘ��0��}�`l[ Ox����2�'$v���Ŭ��h��c\](���<Ƣh2�d���
2�Y�:�~�"h]I����&���;�[�/.�(��TK���|��+L[�GPgM�a=��,�<�i	���>>E9`�L����+Z1�f㜲QaMB��vsX�1��F`���RaMx�(}��vu�V3=�5mLJ��~�ʅ��m��-#� h�����b����g����(���Eʑ�9��Ŵ��uA�ͱ/�H�`-��f{C���|dW�������c�qk��X����%-�!�쯴��� ڳϛ���۾`��3���C�*n��:H`7|�?q�^�r�^�u����T�yHSt�Bw���n������nyi�ZM`ʐ�j�ب{p�2:`��2hi-Rk��B��o���D;Qe��p�����	8;��Yp*�\��!�,�X������5��[���5ed45��Egݥ���v��[N�����{y:��\景~�]۴���d������/^�)F��q �S�M��8����6���y:��+kd����N+�aM�Nљo���Ѧ==~.���0��1��%nmd�N=;��0�W�q�QV���.| ������48��N��2@ ��[[�ɓ'���{d2w�2��
�I���k ��S2�Εu�"; �������1�X�i�a>*D�z���gu1��J����<�"~�<7�M KUe�1�kn���U)۸`���vy��ĕN~���k
�
���,�T� &�?,x���>��G��#8�k=[<S C2���W��4�66�0n�)�nzϕyb  �mmR��5�c/̨� R\#� qM�v�C��@# k�d6392���� C�n�}���.�g & ����^"_Ѹg����1k�i����$���={F`{:� ,�a�9	�5�X��k�3�����D���dL�mmo�3cB���܅65�Y�������X�!��I����t�aP)��v�L����aB�x=�[*��*@���!��γ����'Y�!�НF�blb, �ПH�ʀ�9���i)[�	�T�~ﰞP�(����w��fRz�5
�b`��'u�����&�D5y���}ۿp(f@Zj�
���͕��@m�1��*_�mJ�0{vA��eb�Lk�V��=��]���O��]U��R�i��ϠPY�<Rpـ�|$���1��E~r�����)�Ը������v��f�љ�y��M�1&+S˖@"D���|[���9��'��61���HN������
�O^���CtV���?L��ِ��^=�^�|��޿����p6����m�lҙ sd{k�QV8��G4����(1d5Z��`�R]_��L��ۆ�rǕa�
zQn����_��7�o����������'�
������?�����������b�l0ҫIW�i�]�5��e�93����&1�n/�fѻIO\���H�У1/���Z
*�L^�3E���^����/���n��,0����_T��Rt�q).2d�G�����=�)#�ѣG���.�p�pR�����n�\v|�潋�jV���U��w.�}����N����M>Zi�s2�X��K��Ja8� v����� �0?G�A,�n��>y�?~��%�ӥT�� ��a�0�{��F*a0�9utt����U�q�^��y~`} �6 ��Kf��b*���"_m�v\� v����k�w�wѮ+�r&U����n��ty���6�C;��2��Yb���~F���#���e9����#�~�U�J�	<B�����_��i� �t�t;��nvj6x|_�i ]�Ľ#P	�c�Y0g7*�3],R��r���+2V���,��x1;)�s��N�`��\���6$�.o!�?�Y�魭M����q�
��	"��{ ӑ-�>��g8x�u��[a���³C� �ٛ��c2��_c��(�I�'(��A�p:���`� W���T�,lf�%'Dz���l��EYF����~4�x"��O7������t��=��<��a��vs���%���5��y�Il�9N/�B�ZƦ[�a��D0�dw$�AִF����s�	s,��5�s��V��D�Y�"���@4�s��͜��$@ 	s�͛�|��x�B�����Ѹ�"��y��:�*�NV��\�������RF��k�g�>��u�(�^׺�R�
������g�"�!�|���5x��5y�/��`Mk��KׇJ�m��W=���7�b��P��>M��;-Ή_���XD���g���J�)�V+�*S<���<��_��Om�_�"�~��
2,�ɴ�n�l*nl�h��8t��{��1#�>^�d:��S��	aі�܌��c��:H#b����9	׀�Ľ{������\:��:���?3����=�e���K@嫘X�l@�K�R��f�i���-�UՅO4E���>�RH���`j+3��6��(�+����gJ���o�����R4C��Zp`P�-�V���yB�X"x&�F��S�(��TZ F�g�=$���ɻh�LH��˟�hy�-���N������׋w�j�ɷ�Ңn�6�Za�NZ%���#��� �� ���hLUcrb?�Bdz=���ZM��q��-xBGV����|��޼�n�}��scm@0{�X�����A���	�܂�l�� ��C`ڹ�_���C3���@�qW�֩.�BL��,�̶�E�F
�����5L0��k3P���'�����i�b��s��Lf�OX1i?��Pe]�M�(�� 6��W���C��6uؓ �$i՞�� ����,��r�9p� ����I6-.,��r`5���Y���H0ŗS��F��'� &�\ <�x�i���_�0`rVI�׵��N��q���v��6�ح��(��~ZYYr��2��33a9�{���wuN�i���em����
��(��s���>����^|.��ԡֽ����A��87l� W�뮲FA�������2 �fk�`�6�m޾�v]����`���7�i�PZ�NX�ua]���Z���
��B#�#�[��D�)kW�B�g�10�>!X[)(����=de4y��n�kGV
2���{�z�a��e�9j)�w�����?>:"�+A:�;b_-(�@/�E kթf��5�󖳵����B�X�����{���|�|`|��9!���	�@��z�����h�Sw�����y|��_�[R\���L��ZЗ��I�f8۟�5kx|�ğ�5����
Ҩ�4������N���o�( w��Co����僃#n�e���\��e���S���S����X]�I�k3ZkF0�t\S��R~`�w{H_�k+*q�O��7�1��?��}9Ы<wO��VW�t��O�3�>����Ա^oٌӠ���si��c���P��/���*��d����ͯDFRݪ�݋'��K٭���_#��}�3$Z�N�Sj�\�H�߼v����L1����?1m 1S���\ʹ?K6`���/��~��;�<�z+L�:M�����oڼk�7{����![��fhK��[��7lq��)XS;�z!�h.��4
��:�����q~ō�8��K�6}d��{k5@x�0���:u����(�t���&��p�?�u��D���,��"���# �q�Y�R�=)>���76�/`]�����5�Sݟ��,E����:>9�sk�p< �;� � ��8�5�t��(�S��b��Y���h��cAכ]`FU�o��x<)�'� �9 0AI�b�~�w��h�ڱ��w���0�s��
���o��vL[ ��a��bR�^��� a�����Վ�m3��^\����B���Sr�Z3�D�|L��D�KP��b�����>m<)���ج4b������
���+��(��l�2G�>Z�@�g�,� 3�$C�݋�o2` ��)�Y@���v%���z,	Vc.����)���&8�31��`0܏T�F����Շԏ�w�67)�����d¨��]�_�<��NL���D��b~Ť�~�j�X �0&u�Nw)�h?��7�*��\�26�k�� 艵k�?�1���*$"���⟘s��A&��,�bY���ŋ59/d���e0�I�d�!# � юA0���k��\�A���w��O2G���0g-��︊�|[c#�X��M|�@#��؊���=-�vK�2�Y��IH���Ϧ�O!1QB+�Q8>4���!�!Y$���1z�����V;@� ����Zz]ӳ:��������������I�ڄ'��7M�_0��̞�\�djj?T��|��2�d�y������R|�q�lPG�tƛO�L�!��2"�d��!wv2tg��������4�LE6ʱ����=|��=}�C�xs���DP318)`��ѭ�����Bp�qc�a�t�^�Sk��&�n+k���U��?����/^�_~z��ߎ������������W�?�%��/�:3  ��IDAT�nr^Б��Xc��`8�Ac}�% X]���5�ZF�Z
�0��OJ��H��R�"����*_�R~��_{�~�e�5V�x~U�c�g��Y0��/���a�=~�8̑G��?�3V�ߧ����A.Ƥ8��xԁ���v �	e��(�
�0����1�'�lJ�e�m
 ��@$]>�3g�	�X_���v����ub��qM�؉���M��f���� 
��IQu��͑�W v���y=b�b_��0V(ӂ6�S���=n�2��錏G1-��s��.�n��L��nW�3�`W�/��Rt.yN��uwKr2�+G��"�M`���K�`�B���Y k�8��
b��EJ`+��A���0Ga��ZJR���Z�d� ,~uWS��>t�i�`�ұ��/ ����=},ں�µ{��{\�غn��PQ%,V+�d X�
�]s]�v�`0�kµ4�ü���87�vv��`pV%����0J�Jd�gr� D�ֶ�$�3aT��e10�/��V���5�d��SD-+�lV�b���G�<v�b_*71���r�Z�X���EJ:��&x-)2 ¦s�?ɺ7$#y,�b�`��$�([�ֵ���vʄ@������g�{0�t��O0�{����˄�y w��B�s�
�bOFf����y�X#$��NA����߼���E8=���U�%@1۫�-`�ˈc���hqߞ.˽#�c�[���y��2	�q�˼J uu*(:o���5�$���]0n 
c�A�@����UF��]���:����R ��@6�
k��O��h~��'��d|�.X^�b��"`4:��I��Xo c�5:|���&Ju�$s�% �fEm�X�#rc���^.��E���u�m]�:�ϵ�
�;+.�>�z"� �\/,��=1�ZּM�"�[��P�V��bY`{��`��h������N#J�
��ۗk7�qӧf���#�DS8�������f��eG�cA%o{`��e�nf�8�Y1#��e������.[������G��x�뷝A�o�QP�Z$U7�K2RN���p����IߍG ðq�I�A�{�[y����n�aM#3v��,�+Zd�G� �g���S]��*�X2ͥ_�����Ng1����Н��ʵ��{��Y0T�c|��몜��`D��w�21I��~g��n��]_/�tH���{�}[�2��K����qw�zL��u���<~���c���w�����?���>(�U���*��Ĉsh��z|�	�O,W`��<��^X��O?���m��a�
�L�?��)#KZ]q��H��
�B����E	6�1���׍,jR:Gp�G�\���L`����Xu܋6���i�q����TXq�q�H1�(RE���9�(�_�Ϡc��1|���q�V^˜�d����Ƕ�M�Hݟj ���J�R���;�,���c�+�O˰-.r|��&t^���Tr.�s��rͬ�PbPa�{�o����X���F�ѱ��צ�a|0����"�}v&`1^����4���\ ����\�ptN��)Hh��F �c��k5���y��\��~���u�J�e�{����+���X lv�ʘi3�dy�Lt3}L!��e�����E�~h�v�������5=Sa���X#�dX�~}���V~�Aᜂ	M�|�J0q�h���l׃}�j���ؖF/���$cLb�%���x+�.��-0��k�ǲ�4j�z�2��3`�#�"z��Y,HX ��n���sa�P'{<"����*6�q)����� ،[��2R������HV�c��x@c��``?����Z۔>ѬK� ���Yˠ1�S���;�xL�g���Y%� �Y�}���=w6��7�. Su�U2 ڔ44	D4���9ӟ0�[aލs΁Rk$F���u6X�d�͜2�i�r��r��;�L⑂�8�d���/����O�g`[[Q?�w'\#2�{-�k����-�f��m������u�f1b�o(	���. ��xm"���]�)A��\�0�+�:[E/�)p��S��L�y�[�?v�\�ͯ�ߝ���j4lz����VS$g��˒I�����͢-�Σ�ؕ��$rZ���@��χ�����h,�=��~�H7C�i���f���?v��݇��`hѩ�05�U�Ca���{no�����P�0X��t���a�����O��9q����*2s���^���f0G��հ�/�a�7�����n{��/��?���g�W֔9p�\��v4��2�"�'��T���h#�7uf�=��:�728������������~����_���#�) 5Tu��9�#lk#���B����&'��"?]�9�{����_��={��k���p������z��w�3��T�PF}����|yӸ����;��א��x�� b�i;��攱�km�ҹD���'c�PXI���[Y^����;Z��i��s��  ��V��S pΪ��_u!X�(�((�� �ּ�|�<H�	�k����fl�5���9�!��\��2Դ����;%0µ@ˑ���0L8���1/ř����ƛt \��ma��Nm뢬Ǡ��|�p�{�-tN&��6a��\�
��r��e	���@m\;
�Bv����@�t��~�|�9�"�P"�������܂1iN�9�x����j�\�+(F�է�c��p}M�Q�xA��m�S F�Y!U���CkAva��2/i30 ��!u�1�౎���,���&��3�XkL�h#ZϨv.حE���I!/�ak*���!���Z�VLM�@����46̸�T���a�%Mv����{�M��{�T�p����Z�M�dXFu�`0!A�@��!��ÃC�U�w�9��0|�K��G1����7a�c^b��~�M�$��
���׫v,Z(
c�$�H�s��[�;�Tǵ�o�]�Yӕ��-�󷙥7ow�R�����F Q�`�,H@w�d@43il��EJJ�)�[x�#��.�8�H�����#��!�=��v�̆*r6���V��a+��^�#G@��RI��E�z<Qie&�O��E�PW��#6�����c�
ȗ��P�>��1n��G�Ԧ�5ߕ=��8���yS$�Ƙo>����MJZ:��6��G�eA]�r&�V�;�g��f����u�M'�8�ZRݼ���g,'�ԡ�d�#͑)hS��i�b����0�����ِ���Yߙ��`�P%���h�?tgAE�qp���W.��G5�E����W�'�l?x�;��Ţ&�`��U�fii���5
`v%��+4�3g�~�����n���������C8�b0̇�_޸V�r��������tO�r���7^�ףW���S�w���ȅ��k�:X>�|�]u��ݼ}����2�� ��Ͽ��|8`��gϞg�Q0@�i���"��k�$:�a��EЙc!KXlq����*���Ίꔚ��bg��ӳSj8���_h���lE����:WM
��V��"�{��DxK� ��9�-l)ք�<��ۋԱ�5�R���}!i�^�t����b}�ݽO�I�\�\�I��8�h�Zc���ÃS���;�˃��zp����'�'����\#$0��Ϣ'	C��S<b��2:����ϿH`���gL�v�w��n�|@
���D��w~}�r�0��0�\��¼�D~`cfYK/muk'�Ь�R�����Q�[gX1���&�1N��� �b4��+r�R`I�D��~0�q�M�3@v|�
����@f�\\/�	c���̾��xӐk-u3o�4xe�⚍%6��d霶V�b��Y���������t,�h��������{�.��=/�A[\^"C�*�K}�u ­��'�4�S�n��O#�:�BXggC��B�ؕ���ǎg2�T�\�����u8�}b�_�}d�n�s��Px�8���Y����GZ-�+W��H�Lj2c%�j����^5�$�~����k�c�1$ pUZ����	��N"p���9�D�9^?�zwإ-��q<{��a,����������j�%����`WK���M�	�=�N3���t/ƺS�.
�w�t�W�{@�6��i_�E' �A���)��M�k��y�<�G;y�)˲��E.��x2�.����V�1�{�f����V�c�Xl@��wFc���ȷ���y��2�"�y)'E2e-��B�rW%A�J�u�E�:�� 7;:�MNX���\��m�E_CH�-�^�E@=�b��˚l�~��_P�A���1o����E�6! �e�WZT�|��ɷE"�R�B|�"9����j�TiM��~�������2�����k~��l��.�`Z}@b��l���PE��zPY$0d2�)N6�A��!iD_�~�\�q����3�J�F��z{�:'<(OKMG���\��5C}��%M��HF�۷�	��xg�Ѕ3g��-,��b��7����r����u<v�b䞿��T�Τ0AZ��b_��4�U|��3���E������7ތ	��?^<N�@�~@!�m�d���[�BRث s	����I1l�͍��QV�D2ʲ����`"�������@cmu��x��!��Bb�°F�W�^Q��)�lKo������3��ҌQ[���g���ڃ�t�����!Ka�F7�N��Ъ��C`�{�6��[f9�Hn���
k@�>�f�&)�Rj�9
:qpLh�|�E�"������>1 �v�MZ���5�ؒ��5K�;?����� �p2��D
|?�C.Z��-�j=�E���n�GpלX2�;]�`qujy����{�dLi�V����K.U�%[>�ݡ�;\�;�P в���>�L�O Z��kYg�{>�Í��Js���]n{18�\d�ƿ*{�}���/X�yv3�n
����Y���8ܲ�Z�C�^�I7Tvd�JQ;I�k:x�u�P�a��k��� �[_[g_Kƻ�WΉ�!K�������
�����b�a,c,��gK�tk�eL7�`!��D;r.&�"L���"z9�K���+ښ���d8K}�d����Ne�e���O�����'����^ez�b�[@�_߳���ᜰ)�6�x]�?2[mf�����^�7�O�/`K���2/�3��N��E�QZ��BkF���E�m·JX�n��|���|a*���q��n�O�R�P$5X'%|niy��ZX��̳9�<oS͂9q-����b�qǳ�e�l-���W��G�h�k	�C�s���Y.�8���VBG
dZ6Q��	@�����ZV�5S��ą��VC �H��}���N/i2_��`N�v\%��5yk�.rY�-�GP�/�e����@�T�|)�ڥ��붪I�L�S��WZ�+��^��4 s,��9_&���8��y���1ɍ*��ܼ}��2��g4��l��]����M�E�d#Ӣb Z����.�}qc^ �~�������_4M�Ӱ�9'�e$��U��/a(���csvB�K��S'omm٭�`�����۱{�FR	a�������簹/��vW��s�O������?�N/s/^�$=R�ǋ,�����E���rI���@�u$nV!C�,����z�]��f@�dF6~�R,�_�"c������D]e8w 0���9{�+
�8���g�58�p�0߬XN���C*�2���uHW��/qϟ� �^��|7yL��Iv  9��r�:���_!?gs���]Տ&UL!������h$�a��?1 ��;
�am2m9���Hg�_�xֈ�F� `���\3�P ��,������bdf��s�z���k�¢�*&i�q�tD����c,���37]+��i�I� ���n4�'�GD�`7D��� )�5B�,tT�Ff�AH+��
�,{��P�L��%8�����V\-j5&�r��hLV�T}�W�{7����Ɔ0���8��������q��������-�����¬��j��=���h�Lø��࿚Ae�T�^��w�)��� �4�W��\;f�T�����3�-���}�"� vR��ы @�O�R*	c�@�l�ԅ:�)�h@�G4�e���z��Y�K\���c,��ޝqߢ��ܽ�d��'�[ƤHXo����� s	�,/q��XET������HBs���A���t�n���#�J2����Э���B�*S��	��}B���g�ke���Wd}�2S�>�ۧ�FF;��d����(�bϠ,j9�E����Z�>�t�X�����,��c���&���p�������8f
�$ױ���{j�&��p�|pS��͛�}�p���瘩a,���#���y@��N�ovm�i���c]�%�o1��r�>~��Հd��,um�u�N�Z�9B�����"������`��=�E�Ԥ>�-�$��)����X �fHۚ�k�p4�)��.h/�i	*������y���+_q���4��b���/  T�� ~��h?�T��̪�[#�Tj#z#?���9g��Q�u��kڼ}���Ka��΢1�V��@�j��Nb�Ԋ���������(8 p,V�AE�r���g�'<��`(c&PAJ 7`�ln��q:kQ�cs?:y?�s����56O2*	���`4*�=�v�88/#:(���A�p���ե�����'�Љ�G����g��o��诽T]�!!�hTnN�Wc���0'�wT��c����:�w�-����)�3����^�4�����=�3lZo2uk ��h))ŭ0����jk��@��Y��E���R# ��A ���A��&�s�õ�Q%,��EJX%�x`'��X
���O��B"lJJ_P�C4��%GtRx���lqs�L���,� }�'@����K�d��G�p]�pΡ\q��͝=������Q0:����6�( ��E}"�{3Pd��ƺ`0WI~2�C�D�$ i����m�_�5��jf�.2I�4�$lC8�cM�N����9SR�:�=2q�����7�G����KK\OGԫg���)d�����0�����"�& ޢ�_��zGɛ�J@��7S��?�E�9�1�e ��d���ºb����p	�=\@.��/-��E ���a���]����x5s0�ޑ_��vPN��(%�hlA��
�X���ݤ��0�5�X���l�������qz{K���Fa����s�޿�7'�5+�I_�X�(Ń�N���B��\��b<�U��+-�����1�h�,`�b��l��o���c]����5r�S��>�{5�'S�fala8� �h`��'!�q�a���޻���{��%�G��&Qo{"ڪ���~п�������Uc�X���l�̒:6��9�����W[�
�TGZ��`�c=�|�^�{����C����O�q}��)�u�OV00�ӳ��4[9������X� �������4B��Lj%�����D��M&5�4�mq�U��6@������ɖ�&�j�$��p7<b��l��]k�x�E�a<:����T��Z����� &TXA��k6�ֱFAأ�������5��S0֯S�*����^c)�U"�a�R�}�%�h�����u�~sPN��q	�	[Vv�"�yuM
����O �4����w��E[������5H�7ށ�2���Q��B���ןi	�8��V��H�������վ`(�N7���;8j�)c-F�f,{c��7���e��Qᆃ�;9G`�\t�1A;��yp�=x�zzp0�H�'�Z��v���������
E�!8�����t�L �8l�`a����27dI9��̟2�p؟��Ӿ���Z�={������n0��N�2�bv*n��" M��J�oR�[B�.�������W��f�I�\�8�2����آF!��L��YY./�8R`��Xź�RgGRl�صnY��v. V ����{GY�n{]�Wvd�'C��A�0���`���(ҧ��>_��p�͍u2.�P��9
~B �tW5^o2?��P�f"�^1�1��C�����w��)��(�L1�G㱰Lџа�,ś�o�f1��L�x�Ը�� 7�	��>sOI�4e,�3 ��2"ڢ=�0X�b�Nx���
"UU�������d�NƉ��'65(	�d"V��$��RC�i�ۦhlM[X�L��C����B�����+J��:��v4�/\Z�p�SjA���\MF����)Ƶ�X�f'��&�0)�2aO�q5�X�q 4��i�Z�gz8���'�}l���� !�q��q!)P���
��}E�#�FB��)T��R[@�Ke
p�T�"k~ȘC�u�"�M4�K�~�4� E��0�n�>ȅ���1^���(�
�6Y���@��u,V �-a��_��5����֦�ûJ�3�d�5��c1��`��V@���\.X`f��R��H4@;���)c����V�P���朋X_��.Eg
�N�\\K�3�J���Y�5�[;�����"dL�p^�����?@c��G��0��>���b\	��ӧO���I�m��{���m#�G�XQ@<#��3�_6��9��Z2'��|�
��Z(W
ܪ�WI�g�8����y���}9����X��}��HIT�G�����0�%P���;z�
����z��Q`>�׎�k8X�8'�C���,�� ň���R4�8���X�`/b��udf�3X��c	b�P�>W�7ޅ�Fu�Ԛ�Q1��u���2���(�YY�ژ�;5����=F��!$�a��mV�Qv{��z�^��F3���@�L�Ʊ̹��Iu˧�����!�aτ�c�4o�{�����;�
W�d�M6�*�R��vr��PC` D'�Y���LP8C�v�zU K^=��iF��&
����2�p^{�捻�{�-.��D�z�� �oM��e=�����ƶ��ަv-�> �;�QU*P����i�O���ɳ���뷮<8�<��Y�H�hrݸU]�o��k�yC���wf0*>|ȱ	�N4�+Ь��-�͌dsʫ��YFڌ�,��Ȇ�x	�c�-�/����3��m�/ ����0�Qdhk{K��RXv���� ��{�-+L�p[��xY�z i��9�pȾ ��E�p�i�	 ���XΧ2J�ܿ�?zLiد_�v�^��j��yM&HK��0,�a�k����~�	\�y� ��XF��;K�%��R�
�hn�ߠ�{eg�`K�"#讛� �0> -�%�}_5J�$� ���]>�v;WV�#@.2.�8�1����-�ͭm�{�͠����g3�I��9[�i:�^0�1g��P��u��L���os���1q��|�̋v�'b��i��s��q���д�ct+��@ҏ1e7:�78�2�˲N�f�� ���3�`dכ鯒Y��p`H�թ��p���� ��t|z�?֨{a�ޥ7&z��3A��|���fވϪ)�eAex�mXi
���Y�2�Ѹg�q�*�k�-o��Z$��4~o8�X����߻�v��1{����'��s�u�wg\��6C�	RRLBS_t�{���"0��R*���ÿ\&���vYMZ�[Ӛ@p�\�����`McM���p �b�!��G\;m�0���>F��Zq&���9�Lܷ�x����v���$�g�>�{v�2�-۳��Z�=�}��� +K�̛�y3��7�/l\�W�w%_X@{m�IR$Ok�(�{|?��(��}�4ȳ����Xc.c�i	Y&�_�����L����������),k�o�IX��1/-C�P�1�k�V;�T6��b�c��qO��J4�u?�}M��L�� �_�� d˵gQ�����/��E����<��4�7��ʹ��rM�S���;)���U�w+hL\��%s� {�&��锦M�b�Z3o�g���_�����4.������T���
����r�%����ଜUn���H&`0'�b���6�]���)<��Ǖ`���(������$�)��7��� ��f8��b�.��e�~֣#.���%X�gZ���
_���c����u��5���:�+u�r78�=���u�G�[�F�)Z�0o����P�B�$�ܔq*��?����7�����F)ȥ�e��"��rZX�4��r��5�j��1]Go��q��T��Od�;�e�3��z0�!� �ǥ�AN��q�r��9f5�VG9���� �@;��\%��L���b��<R�I ��Œ�7��3Z�յ���s���P��������>9����N�2
c�	�BU�a�Z^Yp�kKR\��SHk@�H����Vd
@�=ixF�VF���F)�����R�������5H-e�9f훪�خ+���uyupK�Ph������L����;�Q+�E�`K�K��=Y���1��	o��d��Ys'�Td@\�P���F�j_��6��z�9����Kk�xf�B0�|.�C�?�*e�s2�oи�%� �B ^�,2�?u���ֵ nv�e���ʉ�Ul��7g4�I)��ΖT��kv�I;g!'����`@�u�`��.�[G���B����E���-�BfL&���\��X����E�a�{�y �85D��L����V�̂��D��{��m\�<��A� h�``��M���̒k1�4 ``����,�˞���w��_de���T�0�� }5`6KI	 \ ԓˊ������ΤM*�bʹ��$�yT��ї� T-,�`��c!���0 ��f��ɞ��f�rL=w�XM}%�&��u����WY�A�pߙH�`2��ݘ��'ź��
����)m\)<�}�������uk�����Н4�C�|Z�G�t��9��˟��]�(��J�Y�c��2f���Q��=����iv�T �]Q������ qv!�!���o�5��՟����?������	����J�u��pMxN���7^K 	�������]�/�Xv��K���Z59�kݎ��MO�	XK��čϼ�й�h+�6J����pY'wg�>=�`pBwro�=��&ml����<��
wmuŽz���\�#��/s(f�H���i�Ҍw�s�����8�����O����~pT�y�--���Q�ZY0����"����x��j�^n��3�i=:r���l0La4����j��˫dH{-:P�Zjʪi]� �ҌL�k� <��Y���i�Y�,��.��{�B���Ņ)ƕ.	���&27�CdHC��"���Ђ0��.�]L�u
�ӹO�Vtp]M����z� qQ (���Dc�� sK�����?\'�=Hx@������	M�X� ݫp-��"H�X�*Crg�2��y!Z�H��(ߊ���a]=��B_M�W���	�B�>�C���A�������P������w,׎�\�lp"��6X4l�3�;�i � �k#���}	��1s|t��b�X�7 ��@^n�c�R~���ʐ�'�h�KC�̿d�'���PEf�~o��"C��5�m˒�ɵXAjK��c��i �F����"�&nA�L�J0c!� �fݴ����4P���q+
 �I?�p��u,��ѺH�@�;���83��B%��Z�u��t 2_�hg��g˥2��2�kr�8��������w%�1�cc�� ���@��8@�L+�c��X���߿���b���<\D!�G�W��/_��f6�|1�'>p���N���G`�&�iw�t�����N��*��3-ʇ�seP��?�|ng{�����ȯ��:���r!0F�d���Ȗ��Zk��k�T�Tr��S��[����%��;r��N|��6o�j�@=."@j��ڕ�3�YJ�	TG�:	�L/Ӣ�^��4yF�1�ą�1�O�/�'b-����QfD ���ۡ1px���\�>�%�;�j�U�g)����lH-�l���?KVI8.�+Xm�6�$���mɚ����pدp�D�ѓqŤ2�灂�>��n;.�;)�k{D����9W��n�}�y�r�Q�d�]�����}���[W��,��<0��6v����WT���/b�>}�ƣ]5e��q勖��16DlB�`h2E�g�z,L#h6qj��ڴH�1� �76�^���!�~#�m��i���v��E[J�̋n�iUm�c��cc����!�S��tQ�C�l����A����6�kq='�SI�J+�RALw���bП��1o��& �	����MLp$�D�f2X| }�``���e���1��F����P�0a1�&ٸN�Aj]��2��f>� �I� ��5n�m�S#�R�b�yY0 ��T�3�U_�4�݁�EP$F��E��z��uYv��G����XQ�E��c)�`��3?04�ޜu�D'r��Τ ����Z��9�8�m�G�!) �1���v��X�%%�p}V�� "8 � N�Fӌ�K�u-�+����F�1��S��Tr<S��)�ŕ��7iu`6�|�t�Ϙ�&2&0���u�����JPBT��i���f��ۈY@ s��z���)8u}���ؘ��+��ܖ��޿#����<�k�a�O�մ1o(����" f��������k�~}
'��\�v]�B�T̡���	ʙ��M�,/��ёdLM佋�5l��NNV\�k�c�r;�>������na����@pkl��T>4����z?��o��	]N�v�5	�-Ť`��r,�����ַb�I�@�b��Lc�,]Ӵ�dWD�NsNp����qnϘ:�Z�y����/b�,��%�T�Oxnn�H�-�an�:���>p�L����ڑ�)m�~����s��̞e��+����A`K��xm}i��c��`�g@iIF�p��0f儽�8<;칐�ubA]0�W� ��}1O	��}�ԯu5�@$|�/PD�ٳ��4�7"�w���x�3W2_k�qA2pd��S4Vj �ƺ�d�_�)WW[\;``�b��k��σ}͂�*�a%EY�I�vA6��>� �a{b/t�o|��}N�%�ú,�Co��s�u�[Q���1�s]���j
eV���ȋ�������ɴE&fV]�L��Le�\H�W7o�v��6���%{g���.DP��'l�J�j/��e�k��3����E�����`,[%M�:��Z�L��z�i	��#^�#�d^�I���1����``���{����rY%3R�$�n�����pH���X�(;���cq�յI;r���&	9���kuP����sj�bS[\Zp�gy0��x�0J��HwL�boa��L�!�Q��wN����{�V�0
�5{#�s�u��HV���H���B+��z��676�gl��W��,���+H\Q�sUҠ%Z� Ya��l 䄅���u�ƤI'`<�G�a�eZ���ـ�0���
'���c#���	����DY��:\�R�7KM�CJ�D��Ţ��Ν�XK+UðE�2w5E� K�߹�!�?VL�
]hH)_�c�~�Ŗ��(PW�B�Ǳ+uL��7�j��9g�� �[���c��q\+�&HIC^�̳��V�.��&`?�y�n�d����5Z�p��h�䌕�r�wݢZ `�L怒��O(�:td�J���XY��J�C2�j���8�������<�f)�#� KOy^2�!Z E�,�X�4��ÃC?���<�{��!�14�/f�m+���b�<�N�xB 
`�����g	[��2y$�� ���7�!	۹�g�Y��;d��X6'�$��f0����,�\lƢg�9�8윱h��s
J��5^(I�Џ�2 �)pSՁ?�N��A[9��0�jGI�ήI�n����4�E�b��زk�Xha'��/@e���I��5�* ����@H�����(� J����:�`H�����:uߌ�fRz�.!#�������/�s���7� �ؠ�Mg�TO��L_��mܣ�s����iF�u��{ ���j��J��dMC�#���g!XRo {02�`��0nE%9��4N�ێ�y�Q��սP��9*�u�����d
^�L��:��K|�M���u9��׵齫�L�wE�E;k�}���I�ކ=�d%/`��s��h����Z�{@`��2�}nk�\�h+u]a�`����#�/X���F�Mm�C�f3��B5��z����|\22���s1�p���B�)�,�1[�2�+�.����B.լ�oиk�eVHjF�a�����"�_��J�p̒���6���N�ˍ����s͊4�������P���.�W]�Lp����iO�4t"XW�d��߱�z]I���j�U<���U��F��c��'�d`co�^p:>��>�u�h��)�`l�jӸ �F���q84�Ta�����)Lqn�����](����N����h���l���=ѣs0l��"���h��p�V׃���:������N�އS��g�%��B���!rU?+���-̖�Ƣ�Y3D�cs>�͚���ݗ�J�,�ʼ}�VI�0? �@Vl�ℋa����|P�RRa�(��jCJ�jNV|^�J1����Ct��(B_r��������'S��Z�9_��p`1ߡ�:VƭU,�"�^��ŵRRe8`�J�$q�ѷA
G_tZ3�W�N1*�g��|��V��q��3z]Ic�3c�:�L����k
@�Lj5������l ������J�/^��	_��e�ʝn;��� 蓰��Zh�벍�"��ȇ�/@��e`ڔn�n���]3��(I1���5���Ֆ��
܈��h,gdd��1����nu�����-�����⣰/��zr���P���.�wo��}��-���n�3i`�Ir��e�9�ѐ
���Y?c�A/d�,k�w\�X��cÉy'�k��Y,i�c�������}�������4�-2ʵ�D�(\3�-=M79aCԮ{ `�R�3��}Y3F�1�`�e:ح�j��k�.[C]&�2�I�G� � ����b���끄�x�~�Y������ Rrc����h�g8B��
֩`1pa 8���XEu��N�,�9��_��K�iH�Q��iG���0nOO��Z^��W��Sp���ۯ�Ud���}j��d#Ҿ�,� �! �.�:���W�R3:�d�#_�gͧ�ӌ�,Ǝ=�2	T��/1�,�J3.4�@���M��F�#2�����͂�,���0>{��%�~�K���U_��}�ͻ�5�ʤ��&	֐MQҒd�IP�(HDX���al��5�� :/��t�	 Zjle!�3KF�@�!Z���"_� ���%��8nW���O�"]�	�K���+"n�W��Q�k�k�'��,ǚY�d-��L^�,Uk<lJT� ���
K��=�� �$إ���t:�`�f���<3��qqY���)���|���]��r?�ȟم��[�8m�!k{2~��noA�l��.�)�c%F�Յ��<v�vҼ}+m�\�xO_���r2譥�i�|�����$%|Y�������f�?�sS��Dwsa*����N��a�E*|oa�u�Z���L�pD_�ܓ'����{�����
$��d�ߊ��*Ts�ƉL��5r�&+�'Et��j�L$��-Uz��HIZC#�*հ@��h"�l*�
6�.��g7!��z�_�M9��ӛ�/w��^ݿ0V����,,�L��h�f�}dL2/��W��F{F����`A|88����aR@����V��m�㊀��0�I����8Z���r�
�<W�!\VѸ&���M�u=��u2qݒ�ףf��)T�vˆ��u�*p�\�P_�r*�7N���&[�%������ `Q���T��-.@�:yc�Ӡ7m)��38J�h��Un�>{���l�r
fZah����ҕQ?��>ث0.��9e.D�ĔY�K�:�.."-�l@����֦�8�N-
�ekkt�W�U��	��j�opLU�<b���5��-� )LT�Z���dY
	�=�i߄f�3�XM��w�l\'Ӂ{R{=dd=ʹ�@��
���Ч�PY�s"op�ӕ@P���&�� ��|4P9u$#`��}Kv���:�)��	�vվ�r��q�q�qx��}��&�`,ܫlO��i�BTezݖbċ���_]i��c� �%��L��>,�|����4��X�S����#´F�j#���y'��S���f��T����ʺ`OSG��A� w����� ��g��y+�X�<P�q��{��S�[ �����<�u�,�(���d(.-.r�}��ܿ�|�f�H����>x3rl�ɲt-p�-PW��1n!����e)�&��lU]�R�%+��"��C�~2��D]�W�Ǆ�Qr�G[YG�*�ez1����l�ʕq�YJ:��ؓ�T�?p- ��=���ڌ�ɣK���1r	3@*�S�=Ґ���~��4� lїе�Y��&��By&�B�P��<�`r���<<3o������(-�" ��'�Բ�����qT��O2��M�ۙ�5r�&���4������y���DcY��f*z��p�R{{�ȭ���3W�7��k�-�r�������Cї�s��Zܰ����it�)	����'�7D V{�{��D�Mcs}����߱R6�n0m�yG�1C���Z����	0�YA:���.�hF�FM-8�H��,My Ub�{}���b�=҇�������6|��=ln�%�U�}���Ə�����MG���ںq)��\dOzu�EʢPc��HӇM#�E����iE�\a�l����j�9�9��c�S�R��k�<��Ci�Y��Xo؞���A��aZ�V|�j,dz�^��9��_]�i�c�'e����z�Q� �7�.�5X�wq�[1�ۜkq��H��*Z���l0�����<�F�ZW��`�;��zӅK��Rd�j�Y8��fUB-��dL��`VM_5�?�}�5K76��0ż�8�V<�4�'�Jt���hҊ�w���`Hgk�[`
# �},]�`?��1����(g�A|��sU��<�B�m�N4@C0}A 1�͘� �.$��	�
P(��u������7�,�Դ�3]�-m�JQ��z�9u�Gk��Ӌ���ٮ�[
*���B��b$x�dk0��:��� 3	b��w�<�t�C~�č���W�.��	0W|���]my'�cjF������+�k��1�򚾚j��#�˥Ra�Fٙ�5|مX��L���e&9��p���~����¡�Ҍ:�̖s�)��6������>�| �}��
	 F���2]X���:�_K�f����5���+&2�`o�o��yF1�U���E��(ݓgI`�u8$��ck��|ƚ`{X�{MJ��Ǳg�ȴ0��`�ßS�E��f��"󘯐|9<��a�Z���[���]	�7�S	T��@��M�_���w���;�̈��e�q�&�\�FY�4;+~?�1�yL��,�S�^�+f8
��?o��ɭ�k_i�ص R�����b�,�2���޴9�$�Ts�7� �Ϊ�j6ٻ;��~��2��v���GP�=3����fw��������֞f�q $2YV�J wsw;T�>}����	:�u;׹����OkK|��y��rb�8�?�_��/:�����B�O��k��z8�a�M'�0�$*�xM��w��2�W�O-�s���H�2lj�Bt�667�����#����/��������'O��n���"�˰��`,��y�ؙ0`yqa)l�I��0�Ώ�9}	����6�g��B8��`C?������$Ոݖ��SG�):3�l��yz���d�y��F�<�{������LF�DZ��>&�e+��;�Ü�����;�ø^XD2�ù�CI�������0�Y��{Y�����ͬJd0K����i��=a?T�i&I���S��l�/�Y��x��,��:#���b��B�.���%�,�Y�@��a*b��ff�:jG��i�0����C���[�4���i���Kp<��?o��4������1�����}� ����ra@Ȣ<y���=�:��X���� ��'hU�ۂ���,��V�V�6X�A8{\$��6��}��u.1ZHh�͒Aj��H�� P�L�W"�����ſ�9GA�S���l�7��{a�"8l��;;�'�Al[�`��Yb��b��!���8��[�R.�0��K=�i}30]���ux�"ӥ {X���;r�ܢ��{�f�\8v8vN��:U���������\�<eA
/�'�fTq��Y��2f0��}0�>�E�Ptr�u_ּ�̬w��/��.~�✛֜N��;I�g�H����Ͽ���)���[oz�R� ���Mȵ�8�ۑ��� p�����Xr�Z�a�Zx�~>� a��DFM�A)�W�/(o.2�1_�f��j}�O��l�d����pf�]��X����6u��xXo�� ��#X7~|�����uK�5||"}/��T,�g��!K��ǽ� �����m��1S�s�;���.H�F
c�t�����a�s.>�,���iWg�L9!�6o��%���&�k>t.iLEa�Z�}����ȧQ�QR�F�e9�>(���X�֤�ʼ�|۝`,_�>�`���f��ݘs���D�&���K��"�.��N��ى�Xf��A"- cO+���� ;�{zƓ��@X���6�BYM0��갹�����pE���)@�٘�R��NW���ikK�:����L��o�4l�p�F�Q;��t�YZ\B5_4}m���z5�r�Ƥt�y���H4"�q[��ͧi�(�$��*u��0V���8�N��Ȥ��+�撎�`KU�I�; �06Q0�R��K*�+l�˝����l��*W��/s"�N��l�Z੒t�΂HϠ@�$k��t���!]lhkr�=F�5�27���~� 2�B�b.j˿eK��M��@������ڹ�/��8�����0@���\p�!��J�"��n.=2�g��5�Ǵ��r�̷����YD0��eN9}��]0�Y�B��$-���=�dVQ�����k�&9�͇!9�?y�
}�r�V> `da^a� ,������̰���f�טO���#Y���yůi*4��!�1?��������)�i�����m�2~���ȳ��L����%J�:���1���+����9�,��l��@��d ���乷L x�W�Ǻ�d�k�f� �;i�JQ��I�?��2��[;
 �AX�1F�E�i��]��nps͌��^�^Ƭ�-[儹+��ĭ� �C�i��3B�鴏�
��s"Y�8��sq�8���i�˥e��K���_�A�v,e;��B`�MZ㸰�j��e^@�����Wh:w�Ae�HDn|ߤ	� �h�U|E���cߍ���;/%�a�p����ُ�n3���5+*i�}&]!Ep#;�!�����l_Vj�-jARd�a>c��4y�]¸����*H�a���fV3�d%��P��6e���VI�ds�M����A��|K�ܫ�k|m[ଥ�(я'���3IC2�L2ӹ![$��7~l1B���6��k�.g��,
Ϥ����y�i��4�~�j�7R���A���Q`F�g6s�
�}�8mć<�3o�f��˟t��߯��9RI��"���콖V�Ş+�A aV|����3�?l��.Gw�,Oa^D��Y(��SF'
,b���XFAJ�p��
��?'��fU� h{�I'ʜt�?���
�9�����_8eI5U��M1}�i�o�;<�������=�<�#y��r��Zb]�X_�]��7�_w�cƏs�WX�S����qey��M$�oTj6p�~|�)��k�ߏ�J f±�u��P�&���$'K��<'<�\��$��}�B���\��*L��LZ�Z�1��Aѯ�s�k�`o��������l���)������9�Uϛ�?
s&H�(hd:�2�E�c�`Bb}I��+'����
�����g�/������.[.�~�k���v�i�6`4C������%6�-4[�<eG�;�ؓ��A�Ek��:�BxE�#�N��M�K.R1/�� �"�#�WՒ�I�R��5*��Ʊ ,h���f_ �dUǽp���(cC�^��������1�[[��������h�|�m��ɍss�$=�5.&���А��,�`��x-\����d}�3���Qd?���۷�8���`�ҧ�A�wt��S���'YD�@���6���6
L���l��=C�W.;N:��K���	������B��q�
�غ�. �/���c˞!{�1�m�=�k3O���(�*��>A��v;�~.iAת��{��>�4	�j�U�Q
c��SZ����Cu�Y6�����{�wɞ �.��o��j�I��1�D���{.����xo�~��w��@ּݠ�� �a�a��btaa��GRTz8� ���l�ӈ���'2>?к#�j�Y�����l��ؓ^�x)���Z\�z�Oۭ����,���&]w�/)��	�����Y ���E�J�Sl�V�_,�Xy�{2���z,N��2�l�����린�k.�����~/�#�a_���~n�)�����{�j�P��Qc-������������yY�������<X��+œ�Tq��ǔ�.�9\��M:F����d6i>���Ǽ������O6
3S��Mi������k��c�TJ*;�:�����]�D�mpr��~'lLH
dp��Ώ�a  X��L�(��ju8�t�w=���hF�=��Y�, ӫr��Q�p��N��mqF��XD��"��G���3���>�~���?6��b�Z��i�^���:u^��V�(#�-�3h)�I_ 2�h��E؍,�W�������н�ah�|��L��g�Ȝ��;� �<>�`8�N�0�͊�o( '�s�� �B}}6xa`C�]5s��qV�~���3��3/�a�C��rp��iV�� +#�E��P�j��f�K�`��a�i�<5��d�ƹB��Ẵ�D�j������H N#J�i �j�i*��rc!� <��
�Ha�~*Ȏ� �Y�ś��Ph�v,҃X�����$MJ�������s $ b��Jk����� �y�-�l]���n��X��}||������z�X��e���D�8[� n�{R2*�ؤ#5��`������f���c��(��Y�a=��1����=�Z�q>?�꼮&�3�ՍW����̆�4��a�;���Ī�Ɍ=s�]d:�4����kA��s�\���i�����է`ֶ>�z}���LY������>?kHx�$��ׯ�nI�3]�s�W�-#�k����L���,A�s���sK��<H[��H�|����7k�j��<`k�
���'O�VƤ 0��Hp�� ��W��*�����o`�ו썰%q\�¸���v!�S���ɸ#�j|�X�@���!��loo3�bY=���������Z�2j��-����&k����%��Yy�*@$�r��0�ɴ��`!"pLG�<@������#����n1���m�
䥓3���t���%	b��� 6��6�k�����H�I �61tӽ�pS�h��L7ѝ4���/��;a�w;�N6Me�/�O���~��̓��1xs�J��o�+؝�-P����w!�}KTΩ̅E�jo�����3��%#���5��F�d�`]7�ϖ@��)�22�ǈ�ɩ���b�b~�Zm�K�s��	#�7o�v�mҨʃHN%H��|�s��'G����v;�����X�R:v��yo�]
�������_�O5@�"���c���_Ɖ3y��)���&G�
�rJ�B7�s�C��k�tKZ߸�ZlǇ��X�V�#ا'�Z���U���Q�8z�l}m���uT�/)��$�����C�M�o ?��+�΅��Ͽ~�������i+8\����#C�����BS�	s�޵�S:]zv�a��}��l�p�2FCr��n�|Fo��K�O��ւ8�]u�v�c\���ʨ�a~f�E�iy��!��4><	N�%y��n��ܢ5�M?�����u�� ���jʌXgc�ˠ�0�hHw�%VWʦ�M���f W_-X�a"a,�V��KL�e?{L��b� � b�a�FD�[&�.U��ZvD㶬1���x��ڴ̮�ر� T��� Jl8=�*~?1FU� ����x�a�h�x^��9K\��� )�Z㼖bc3�O���5u�^���|߸�A� �?K˒V�w}dW��}g�{�{ѻw�����2!���b�Qm��"@2���{&O�W�������A��Y�� ����=���m[��Pdw��K�V��Ʋ��=����yqn�OXs�A%Ҍ��ع-�Z8���L;���6#���:S��oNi�N�?�=TXF�/f<�o��k������`�c�E�~�:/�H����j)�[���}N�Ϯ��]2��4��O�^���7�k�qX�����iް�0OVi6��Q��i�@= \� L%-d̷U�l!�����*�� ���|p����,𬷯����tOýGQL�*��E8�1CxmM��6�n��.F.�ĲC5�1Pp����|�s�a�K�4I�<��n��A7����#d�p��<1�pϱ�uY�vQ23���]s����p�v�f{�?G��Ib~J1jc�N����ج+����k2��d�]�d�rq:�b)��۬�u�A`�@ *�{�"{�@j��K2O��Ű���IShQA���U�k�k�z�o�E΅�E����9��N%�}U�3��2C[ly!3!p��̏�	[\�g㎊��.3{yz��5G�-�:g���,����E�g2����c�����֒�H%ܼ�l;�tjƽa�^2I��ҕ$>�Ê����H�)�ټ�|�g�eO&�������M75Z8�Z� ��&�vZ/G�P�{EJ!2��2o�DW���.�󯮮���*�����nw�O`�+�WuC�΄�+�p��r7�s�$v�J��A���&]�=���9����2 � ��ދl�_����ݽ��36��P���^o"��"Db��i������T�7Y���l�	p���Y1[�������n#]��߾���'�"�?c�!�h�S�.�.`�S��C�*D�p4��~0�P�f�l#�1���}Z��-�����C�|�Y/��ZY��gg<��$\��$���:�K�v��������,�Čo����✸nMLOV�m0o���8��Oc�٤��q&�8�\�E����P�Tk�ܟd4�L58�	Xv���p��p��+���c 2��uq���B�I9�c�g�y����8K�����5�jEfgδ���Q<>:c�a0&��k`�ecj���W�a�*�cI��3f������aRQm�0��� �*�K
�a`��g���ʲ��D����-q#`>�raN/p��E1��2Ntpt� �Ӎ�j 2��?��1�Ԉ1'�_���y��o'��\�|J�Áf������#��8��@��L^��va���F��@d���e@��{��t%n���	d6e/�ۓ�sżhkQT<w	�W8ž��`�����㕔�k�;��xY:9�@"��r��8o3c��þ	@	 >s||�?kk�Q��ǀ�Hh�y��f2m��r~��" �b���UM�ruzs�4��N����ˎ�אyb{���H:��Uv%�U��TP	���2֒�����5��v</����/�꾕ֶ��û�lH������sY�L�	�iӒ<�Pá*b��c��"� ��Ҝ��$�2�5��4S��queE��p����Iҁ�(v˲��C�OY�e�c
-z):ƒU�5eA�~X�x�h�tÎ�����#���p�5��������Ͻ��%k@C��1�&��j���@�$�������{ѝ�(o\��y�n�lR��L�"�u�o�4y{��.ɟ*��^e�X�~/��:�M��eK�ۼ}V`�ãb�gZ��bv\��L�͌P��t�Qj���:H�Pl��&6��e�z(�p\��.
�մ��N{�����?u���tZ��#E�U�[G� ����)z�<��Dw!�EU|Hi�ӿ����/����o�����cCgw�N�N�a��cB��*8ypB�0���%��&��YgQӛ���=!��Z��B�2%�+�5����KG�|>f�ӈ����~����;IG�y���k"���@��Nst놏�q�u����D�=	sN5k��l1d�=(Sq���
�4� �F�<�d946��qީ;I�B��V,r)i�p�q��/db��ү�k�%R�F�*8�H�Ǣ��kI﹧�4R\��_��4�g@�=�Taզ9��Csq!NM,rGV}r^[�.�J0�S5�L:=;���8 z�+��$B �H?���8E��6�Z��Հ���w�f^��D�y����	V����Gl�:�y���.��>��k<h� dpyy�5DB@�U<����7� \�X�!aNhD�s�=::{�{���C ������}�w tV�2p~À����+\sEuW�x���u9���y�[�P8�'�2X'`�B,�ɯ�9�RVY^^k/�l��p,⮵�;I����D;�y.���tJ^�ݽ]����t}\��`o�^���Ԝ ����~_4�a���W�������c����l8����3�,�s ��Ǆ]�\��C�Yp�1�뀜�-�7p}�߼��B��4miP�����S~��n�K�7�].�ʶhK��-��Z�>�ӂ�]M�$�.�������� ��<����y�Y����5=��G�cS�]�3���d�&2��?�8�e������-^;޽��{o���M���$��/��XWp-��V�|�P�s�$�Q��w9o_vKk�x���6ہ��<�`PY�?�X�M�6��vW�2-$��E4�U�L�:$Y͓��t�`����{g�n�}Q�fm��4;u_�@_��BV1�f�.ֵ��S�G�k�`}����R�%�8@�����������`�T#�a����- �>�s�Έ��O��R�O��\�&iƚ��5Uu3��"i�Nc�s}����h�6oҜ�������0a��l2��"�"�������eʖ�W)��Y����;�K,�y�r�>��t�F^��7�d�����.��=e����9����8�^'O�B+d�iY����˗o���uz�}/l���~!�0ǣ��D��NO؉ȋ��uq�����o��0��ِx��3� u�p���Hc?���z��r���ҋ/D�.H
�h��k���@q�V�@dú�K �8h>��R������O��������6�g@��Q���
��~|�_֜�;�K�����}4z�����=J׉񴹹E����C��.A<�����ok���M��}2�K��W� _d(4Px ғ������ �a1�����ʌ拋~8�9�՘?et(�{,�20� � pP�c;b�D�,S�*�)"�K��a����LJ,-���
���)J�P���G&�k,eH�t�S�Q��\a6�"k0�1(R��H,�y 3�ʬ����m&=�vu��m� [�a���,�Am�TY1�8/u��;�w��}� �x��<?�:@d���>�= ��8��n�icL!8���C�1��:���1k��Y[]�~���{��:X����o�,O%Z���dm��e��Ș��'8� ��1��S����f�g�@���q=��������CN8�ĩ&R����Ժ	�������/�Qy�`;�_�{�>a< ���g��f� 0b�U��'�3p���{<�� #�?x�&n�ƛ�+)�W�uH3�8���-r�Z�ҥO~��	�y\�&�E�(����L���Y�����1��=e��bLc�a�A#��򱐞e��� �o�7ˉ�1
�dtl~0�(�������- �u?�D�E�b�j��<��k�l��o9�bnk?�<Tnj�y8#ep}o߼��VTn|O3�jc�jf�Z��B�����9R�
>wTNv��C34]l\��#��ø���>�|oɏi�N��s�A8�ވ�ƚj,dR2A���>c]i��uc0[�`̦S�v����.El˸��t��� �m���� 8%M�B}\���W�7��u�7ؕXm[[s�^.hM)��Y@�p_L�_fs��kN����}G�kyC
�p������s[��յ����S���3��-�"F�%-�Ӽq*�eE �.��Ud�2��4��N�Ϻ}����t��[M��[W�%�أ ��;�V�o=���>�*�1%��ԅ�c��U������Ղ�����6��ac�,c3��eC7 �0�-\DO5�p�S����f��7�R��*"�G�i�9e��~W�Ba���C�l1�b��oԇ����k~miy����1Ř��~�`� ���h�c��m���~���wn�̠��Z�b�g������눫u��U����)��w I|~�|��	�2�N�mM�+�1�M�^3s@���*���vVH��0v�~�菁\��׺y_����(X�A�oE��q��s������'�N�񸣬)�9vܧV4��\aX�^�4���=e,�TMX3`,��tW4ܬ��%wwҸ�ȵ�.���r��C�+gk�b��� <Ko�� \0� p����9)�P�dj|*3��T:n�:$`�j�)c�E�����Z����e�ټMj�.c����0�3�YZ]G�qp�Xp�)�������d'# 
�!���H��Vd�-�����@F�;� �d�$cA�g<������	�����/~��ظ��jhl�su1_��8�,S���@�5�캳���W� s2����k�����b!8� �`[�NI�O�g�u�c�����c7�nN=���sȻ���_��y>��>b���֎�w;��$��;88������'�t�h}�	�gj�Z�������R���O��{R�o�%�O�5[
.Ϙ���h�΍y�������G'�'j�GV�i�b<���>m���	���y|rD�k����	^ ��1$1αC��4��L���=���\�R��݌9�l�5�s�3@~�6�s�&2|�:{�Y& �!���Tudz��<=���}��	��3��X����3\��=��ިu��ڱv@v� /���X���\q��d���Km�4ü��8�^�����U��;��vac�dko�䁔|m5�%��0�����fX���u��C��'������u5��\��BD�YW5�di�H��1!���Iɉ~t� ��ZW1���rH�����$-<%��J�ԁ��d���������Ǐ3�m,�H��g"�pr�S�k����G��m6V�}��j�Lb��ۼ�r�!,L{�3� ���G5P�4Ì}k���r���w�u��i�� ��C'�׬��!4̸���O������X7�2��+g4R���|�J����Gk����`����R/�𦠪ס��}ڹ�M��ѯ~�w�.������]��5miQ"�oѓ���qFo��(8�z詏j�p��v	��W|��r
#�T�, @*�<�{��Y��;�HS=89��~pއ�l4��ś9KO�#޺�sp.1�DR$�Q���g�����j�ƙ�}օھ����©�G�92��#q�";G�2[���{K�5��|Kqt,��1�o0���ZX_�Q������ړ��4a]�6�Y�����E�66im�%�������U0L��P������d�3��d�A�����i���B�ܘ�\��#��@��9<8�7o��w58������o��C�Q��A��>�q�f����
����|h0����޲S� Y%r5�`Q�D��Rf��/�M�oʱϣ�bd�v���M����}fBE�?�19��
��ZX3zt~~�c�wN?>��Sx1�OO���v����x��;�D5%{���k'��R$M���ܯ��)4ӅcT�V<>[k=� UW�9�B7kv��[�f�e]�#N���>�8�0���V�3Ƽ�
�p���.�x� y�<����w��	�'T09�0V/�G�;1�ӳF�ٹD��l��#zeu�>x@O�>a'i�p>�yr|�{OG�g�	𓋾���,��Jhk�H$I�i������Y��z ���@{a�_0��S�M�8���yt���������r�L����0R._�NOȸ�`�te�G�Xi�D��\�?�^�
�@��pA��u�}/iҨ����r�5k��ܵ��@6���q8�����:�AO%�c�fʸ͵'�!7XS��d`��7����y�G�J.$��{�ff���$D �P�R=j~���^�~�ݷ|��0מ<y��,H�"����0w���n�]اVy�`Z �<J!���؃��{{/l`
��83�Y�3�*��j��nq��wЏ)�z�)�m\f�d��\�ӈ��>d�a�@�#:֗Yv>9���`d��~�hɃA6� �,�@[�c4G��ü]�&�]h�f�@֧\^њ�R �5?��E�HEP';���)��)XW��^�Obk�sL:����K<�)��~�m@π�1��H.�QhJ<|�Z����s�u��s?�_�u
��i�c��9&�G�t��b�Yq�Z�l�:8{ \IK�{X��N�Fi�c��ml}v��x��\5�㲞�me/)�~W�X�l�0R
�ۼ�NK�^����g�E&���~��H����]Z��D�Io��)�*k��ϼ�i`9���f�4bu~$B��MP��b�e���.�ͰM�^����c:>8
�9�^8���Ά��zG�ӷ��7����ۿ��{z��%3��
ʒ#A���E�ۅ�N0���:_\�(F��/�܊>�S%/�<�h��v����!u�[�þhT�	�nqL�7rNG�8�4�"n�馎�I������ŵ��Q3�w޹F*��3�苓��ڴQ`��dL���dNl]����c1
s��X5Evl~��Y.2�L���A�Vζ��,������4�)+��׽�.ʤ�(��s-`����z��˴�[����0wi{�>��
]��v?���R�=�mpIug&�	1P�"��1�f$A�n(Z�;��3kcc��B_VV�Y�FܘÙG5���(0�3)E� ��c_�'�`���`����FgOo�%`G�����\p��B7y�,��Hze��@��OO�� ���S�%h�����^�,DvFbq9� ��T�:>i+(�`ZRg �1��A�ER�I8�x�.�j��-��:�`A!9�eK��{}�QLǵbE����F����@���C0�d!$�!�,��EArDR&���}Yf[�}sk{{�A6�ie����c5z�����_��g�YdZ�2��W=��5�Y��6��x�s��}:�,��|�S��(5}C��9)���3�������qY��Ҽ�x����[(2`�R��r(E�J
q�qf,k�# .���|�R
����~�5Zh�
f�~ �kտ�󾷱� K�2]R���F.c���~�V[=��6L�3>��&��hE)rG�}e.#�����3i���:���w�n3��Jr .Q����س�_jH�� �>��蘿�f�x��>�Cf�h��c8�PO%e80��5�oʾ�y����i�@��}~Nx�k�d9͚���.�8���"[����u�:¦�<kC= a�#0������ ���=e�;��w	\vc���L��J��eI�Re/@��ۄ��-�x��
�u����&$�K�k@)'�
t�q�5�8c$����	���I4B&����W�xlB~�� �=�	묖��¾��m�D�a����g��vr��b���KD�zӜF@��������1k^�M�Kl�:֌�m�>,ѡ,�hO�Ą���>I͑>�P�J��^��B7�H��y���	��_���K��c�ӎ��7r�:���1B[U�9"��sN�gwi'�����4�<�n�F_m _g�'��C��:�����C�B�o���-��h�`����������������o��w�Fo߾b����Ga�.�yp��݂�_)�pA�'�"_qq!|$�휙Qg����#0��ȖD��Y#��Z���)�0��~A�sv��nM��YW}��<����݉Q��oܤ	��6�K�/ն���{,�T��N=�a�P��h�PV�J��I�";���f;���ݗ�z08[)�R� *7�3f�5f^���ÝkC/�5�y6��&d��"�]r6
$�,/+jt~>`p����dÁ7`c��'E=����^`���~�7o^s��7�|\bFFJY�Zl�m<6�`p/������T����2�b�A�.�)S����Rp�(����}����6��$]\XVЁa")���\p/��M��kM�L
������p���hΖ��0E]���V��QA*7�t��̐:��w�]��l�w��������ƍ�U�x�cI0�����lb)�h��i��-�x�v����� �+�R���-�=�����_h�>8��Nx��i�y�`��˵@^�LubQ����[EZa�Ǡ9��nd�=g�#ؗqL�{fq�$�)~���R@�Y��Ĝ� ]ZQg��:ߡu�,�����\Ώcu8��tg�Sk�*����?��br��@�����>��=\c��ӧO#�L����a���`���8�	������n�������K{�"%{d^�o�#a ��`���+4
�x�#ؿ�����-�kk-f��^���9K����Q�?j����>a� ���������`�5���{T�x�:�R7 ���87�m�-H�g1�y�`c�vk�����V�}��=
?��d,�{4����/��k )\ .0�q^\+�ݼwo� �U�vkD�d��v�ȩY=!���,�������Z��l�sk�x������b���j����#1~O��&�I�+δ���IJ�m��Z%���`��N�����L�p�n���t}ע{�b�ĜB�VG*}���أ�����q	΍�VJt88\�뀖=�3��֙�Q+��p�Fv�i�kE6�E��on�H����r�}��%�k��`�����f�	p��L��qϰ������AՏ٢C�ɮ��[ӊ�����X;������|�����y��f����}��K�(d_۪��?���Ͳl`cS��i������'����6���" ���E�=w�ak�Ae*��f�&;:�M�"�i9��$L3��//н�5��`���{T��P?c�˛7�����侀�6L����w;���
��*;j�K`\����/������p.�Yd�
�댹��8��#y� ����o��~zr��
���ll�z�y�����К_���O�b���m7/ �А�l�r�qň���^6D�hᏚ<�9d�M��Ô�/2��>g�/�ޏ�����~����.�A*A��8�9�պ����)e�"ՀЁ���ɀ^����e��0�*��@�m�P�+�gS���J�z��"M7l7ٌ�������*����CW�����VVWٸ�ju��L������zp�Z��[�ٴaaBR���ۢ��;+�qrr��������Vp�Ys���ܘ�ڑ�wC��h������	ch�!��wZ���{�2`��W�����p�_���]��Xb&�)�����\h�ͭng��6�X�do����:�)�6�[�Ch|n#zmmCR�Q�ԕ�?�t�J* Zl���b/����5����� ���Y��+n2���-��#�S-Fc<��[ke�k��ܚF.�8@��Y==�$����hii��w";�
���`�oV�]����d�
��qŚ�a<m��,@e�R.R%w�� f*[{8�>㢙H���6��|M� �n1��"���0+a�Jq�xqv���Pf�:�2�|1K�4[�"m�6��4�gʵ��R���R�bXW3��Wf�w$��$J�Μ�m,W)�w�u j���z$�G��4k�3�g}�oY_��eLX1U�@k���e,ˋk`��x$X���+4�~\�(H��B��8�ρ�|0@;�u�4����
�����d�l	l2}}2�7�k�p�����{�A�x�O��C���>�湭��M�`�RnmO��Ϫ�������u�%���l�˟���Dqv�]9�
��X#�il���z�Q���I*�s3F�͛��EkYdpDk��1*]�EF��Ys��&-�%�ט�
�8�����m.mQXVV!�+�22�@L�D0RJ�V�:!VH�I��B�5���,�v���˕�kV<k6�M���N���_���t|t����p�0�����>m���e��V�d٘�f��l�����7��|2ol�����{� 0K�oY�u�Ņ|���
���'OkQW���$� Ѿ^+��c`���l�?�c���5`SX�ׂ��6o����<�"�ns�u�!�������q�ň_�� ي2�<���bɔH��`@��r4r*I��&8���
�����#��)�?=cYA��P����� e�+��a��X�U�y��������Mğ���(\�'̥�E��^���U���#�UT:��8>��?��������o�0{��A�b-L�ZtK���ȫ�W��ӻwo�����rjc��y�<�8am��aS>�?�4|��p�ļ���9�@[�h�a��J��W���uQpb���V�A�bC���s�1Jz'칸&�t��(/ξ�\�_6�����<2�g�B���9�#O���IZ�P�`��J좸"F�a@rq��c�8ꮌNI�k�n=� R��¡�c�iQX��s�͢�=���5(@UX��J�����k5���k|��1T�N����u�_�x��]z�������EY��w-���:�
�H�?�*���<���gv&3�pWJq���������7r@K��g�P�`�=��d�^��сg'�x�0KD�`�>.�V��n#��rd��|��U4��0|�� w'�3]�RӴ��K��s��ŅkX&Ŏ�����ň���������贺N�CI���4�i�ieyI��6{��r����Eq�:<�����K�Xͩ�	��� �o ��ց�乊{��/�1�,��b��I�W�"����e��g�26x=~���eq~K�����T�s0�Q�Vu21���*�<�*ݓ> TF�`7_��.��j��Z�w��>�jХ���� p���e�8�q_�Gd�9le�V�^�o���/,슟;�}�K`Թ��y0�- B�]"��`�}�VZXѤZ0np-3"�#��Z��e�g��\D��Ai�b�T�[41�����=[��^oӌ��`Q��ƺ��I!W0a�a���[{�J�<_<Od�.�S�A�	}i6	����
k��~��yaoX`�P�(+�����s =g�h�I�� �>��}�.��hpNi^�6�7�׷4���o��L� ��g�ey1�蟸����=ǎ��2���
&�bA.4�=�5 ���xV�]���<���`O¶DF��-��� R`���b�jX� P}���ׁZ�:��,�V��g�56��W����"�w ���g4ԢxK��^����}^˥�m��*��W����p���LX��0��^raR}Y���~I{�~��hج����H2ma'��l�b͒9<�k.^���7����ހ�� ��X��&�������X�V� u���S�s���C[w�k񯢈Z�Id�N�<7/p�t]�7�28��bP̜�f1]�Y~�)�$T15�����d>�PNH~߿��mY�|Ry��b� c�Pd�M�m�v�>�,�5�j���fpd����]{OG��ѠHR�޾}K'�����7�zF���������ϴ�����_��	��2������ufE ���fc��.X����iD�Sc�>9=��⌝n�u]fC�ϋ�/�e�����ѳ-�����yx���H�M��
�iA٬��]l~|����x�&�&߫3�C�.����{����{v�A<�tz�d*HR�a���4�2�$��BJ�ӂ;�J��p����gG��)�ӯ-W��9��j7������T������^���N��";
�xI�c�Q%ڙ��[	ci��
�����ݥ���o�3�U���0�~�ْ�J덑�+�o�ň��	��/���N���x�62��B�5�Ƀ����x[u����� �T
 �sѡ0��>	�`��z� ���jLt?���c`��nc����X��R�lbQf���.w��L0��:�v l�0�j{��x�Z ._� �M�v �N����cy'v�O���]�Y��*���� ����`Gj����?����ؖ��+���Bw�<p�dn *�dB�4��i�DD���3�[����+��c �cc�\3�\�Eo�v��boB�8-�\�,��o��Uԩg��%'��|���'���չGƍH܋��`���^��\K +���X
�O�?>�Bp��k���15�zK�Jp����K��L��"�Í�Ҏϩ�+f��6��49�<K��CVK����l/T��2:�ź���J�����`���N�@��a�E?0��eA�⃟��ұ'nlnD�Uku��r�e����4d⼰5���A�2��wT�.������f���ZVp���W�j�bTc�� Q�/�	;�?`���²�G[_#���1�6Qُ�,�=
��Nd�`�g[���L>��k��8=���f�YfE
6�bV�g�N��˒�~��>�:mͲ�Td4����K��JV�\ ��i���Ȇ��Y�G��ζ��^"zԺ�J���;�IqaO���X�������t���oA�y���j��&���YX�SA5��B����,#%!%*f~�p�k�Kb8v� �)�ͤ?�0�tަ�X'l�~˶�:������c���d7�\�f:��ϛ�&����0{ާ�3.�w��T����E�$�:o��/���3��o~C�[���$������xJ�酅e*]�Ӊ[�q@�>�r8���S�[�����&�������a޻����{P�i��m>ڠ�����_�Ƀebk�y�����94�goxo��Q��`�V{㳊� 4`�)��*�y�1������^�b�,X0PX��Ht�3�,��-�x�g���JGeyh�>x �[p]f�����(#��!X80�����=��ub����~�}0O�O�}�'�������e谶�W����k��" ���!���ݻw���.��` ���_��G�iqa)���k�o��B����y� 34ۚ�Zx``R��,�c6_>�9�|WR��ٗE�)�i^J���+��lF.�v)�-eK�`�]+��4�#���-Ĳ6��
�Yj%�e�?��#j�B��m�ɀ{�g�h��H��X&��6��R�0��	T0�Ԃ�q}Ę��E�S�ǎO�	FG���e�V4���u��\�,^��f�Q,��Ç������h3��R!��4gf=�ȧ��|_:���\+K\��0�`rk�އ�^���R�-���[[
�f�PZ���jUtpX���Ri�:>VY��բQ��9%i����p�\~�&S�7ʺ}c�Rp��h��s۹��Č��:'���}N���}��ao�#�!�E�l�9]k��,,���3I�d�<5�7���zQb'۷R�l���ʙ��I�/�3���]nn�U�ۍZ�.z�<��%�eޣ��@�&�&>��b�RR��*�f���� ��}�� %[r�Yg�� ���U�8�#ER���:䲦���2����A/][Ƶ�3(F�zV��#)�f�7x ��qE)��Z㺭~
���Y�''txp��	�z��C�������7ϫ�L>����=�K-���X�ybpD�⋀U��l��+i������ai�.y_+�}��◦5���'ξ/؞G8�"�<X��2�ۗѮk�E�U�twW�\�6�I�]}�܉���2�č�l�*�������f��V}.�u�ծ���cr8@��.=z���A�`��z�a��1�Z I3/cZk�a��BEبա�q�U���V,�� ��w j��{�~�=�~���ܣ����66W��M��T����˽�y2�e8�ed�����!��M��
rQ�Z
�0k\o�>����_П��g���"��+)/�lZ�P��wʆF�\U�j��.��٥�������3T�S���%ũ�}��υ�H+M��[�0!f@�	h��:kt.0����?һ�/�}D��c���_28 �|�e���X�d$�Z��yq�s��~����<W�� x��o~� ��S��n��@�ѿLv�c�2M��������,m�M7#�H����*�-�:fc�c�^�3�$��9��eq���Y�(����&���^�GmΑ�>?-{s�3l�_c�{�2aDj�K�nq�����&4�~srs`�iS��	{�P=�x2�򖆡
�O��N�����'����r���c��e�r�������<Ӛ1��R�E9�$��u��l�Ս�Q�@��f����O�G��-.E���޴}d��|���4���Fn5����o����yz/�`R��ԯ�6;��2�scG��^F:::�������5(]�g��pw�e�	��2ڜ�|k��X��R���Fy�X��/<��weL�"�[AY4�Ɖ��������4�h!�������#p��NNx��9@��zl�[��	��Z�<��F�������b��7o�4ŀ�#��9�sX>?��X;�����zS٤&�?<:�s��ZD�"#(��%L�I\x�?~��\��:p��!����T����/�M�|�y�Y�O��F�Bׅ�Vp�'�-f��*�L>��K�����e�r-3�8Kڍd&��0���~�vٵƃ�Y'x�����Lh�Iws �\F�Y�y���Ε�ۋtvЗ�DGa�_�.k%��5��������;�O��?ӯ�����iw�b�£C��3�k�iڡaB0  p:|(\ �,���<�(R��B���ѫ�/���k:9?��֧Ϟ�/~���RO�ieH��F�$��!��׹�t�����3�&�}�s�&Y�l@.��r %�wd�|N����8��)^��ٖ�Ÿ1H��4�Q�-�9�8h��Ê�ȎOX��`����z��1�|��Bp�������h��/�O����w02��%�����_��2{	���w����	_ �Օ�h�����6��DgM��b*`*�{���/����Ǐ��.��E08!Sa�p�S��4����At��z�g�;��C�8�[�cҊ�}Ug�����Gji8�����P�	���dja)�Uh��4B#K�#͓��,%��-���#�K�z�����ޒ3o'�M7���G���2�y���7����v��P�@�X��~��ɵ�?T��y����1o�k �I>H�i��,�ԗ�D��>�ɓ�\��W9 ��Je�̋���@]��w|,5Z@���"Q#@1Ή�3�>��@b>���2u;�F��׭�X@������ЙZ�����9$�px�q��7
�o9>� Y��Y�� j��XB��9��ߋp���KgA�BX�f�sQ��'�|��U� �SDV/H9������Z}>���s��υb�"�LR�-�i� �Ϣ}�@]��"�,�|�dZ(��HY�7P�x?����e��h˶S�Qm�$6� e�3�1����]�K�m�vIP�� ˓柛�����e�-i���'9Xz�K�}��>�}�aqNU�gy���u��o|}B?|�mп�v��ӳ}��}Og��e�2[袤������ ��b`[�[�+1
���m0���A�.v/h�`�^�yN��-.w闿��>�OE0Z�	[h�^���ܸV\!���F�{��ݱ��Ê��
�Cބ����D����������� ����"i%B����hEbr7���z;>:����Q06(��o~#���2������E��:����=?��R<���y�֟�����/����,�5�����:���^g0���8	�>�2�{��m�
ȡp���Y~	8M �eL��\�r �f�P2	��`n�J&'�:�ۄ^L��� �][K�\�k{��g�C����Z�.�>��T�������y�&�Te��ɰ��s#�e���s9k�}<hp��Q�7��>��>ո�����ް�ʱ�$��>�R�B��ŗ�W�+�~4���5�?���d:"MC$�R��A�l����Y�[�$�r2����DF�H���-��Yv#���p�O��w������!�h�˞�& g���2��W.����{d���Jba��@so��j�DfA&����Kˋ����u=
��,<@W>�\^Z�:����7Xa�Ȫr���T�	��%�����rݒe	�E�?��ni� �$f9��59ك��;ݜ�����?�\��la�O�~�"��U�1���^���;�&�\6�}$� �ҡeR����[���j&x6óq����W>�l!�&`�|LC�����/�W�E��I0(VW[���H_��~��O��y�d�KO���$l|�ݡV١�/^���w��w��%l~R�t�a�]����f��Zo�GDMQ]E9 �Pq:S�zG�I~�K�'�tvzB��oғ��_���=??Uè�A}m�۪�z_5�]��x�[D�0����Y��������?�������i���?v�����ϲi0�Z�^�� ���.T/	����]�ڸ��cm��=}Ƭwh�1#Ze	F������e̩�l��-J��eN�}�����`���ׯ�|��������:���H��!!"_N�3���������D
V����v0������#)(��*<��),�	*�	)���y��v���O�\����������W~���q�7_˛ Ui]�'57�M{v�=�g�rs�C
�͛��A�)L�K�ǫ�B�ot{m��س�.DhB�إ�6��0o_Z��C��l?	�8릮�7�b��ͷ��� �:c ��
��a1�P�'��vjsb�T�iQMo��5]b4|�'K熏���̂�;fמ�I�y��!g�"�����++�Z�N���@eV���?��0�l@���Y��#a���y��1��[R�����j)̺��λ������$��1����99��(T����}�z.l.�@s����G�3Q��( �q�`E��W�!L*e�;�p;@����_l�@�+�� � �E�$�k�dd�a&}e(Mv������	��_����"��طz(I��]m׶&�twH
��7��R�۰i�����-@�NYгgO��n�l�����&�������``����;�+�ܟMD|�W�9��!r#�l�?���NN�ؘ�+��y�G*�`s�`tKN�������(`����C�nrF�n��Ն{Q���	*���|�/D������������sN�K@eƺ�sV.i��fT��"�\([�{�Ն�ջ(hw�=��K��U���_cq��A�-&�s�͆W���-�KS��:cb �Q4�k&9�lX1CR0j9�������\�wAo޼a8�DN�r� ��<}��7�=6�b0��=n:(���]Z�ԅD��ECz�Q�;i��M{	;�C��O~{~�IQ7{z���c�0�$���0���,e����Ww&��>Ϻ�����<������!�<<<]�����\u^��Q�f�>�ᾂ%���K��e� �.j(���;=cb��f�v�by�j�|+��π�F/l\��t�c�y� ���K��\+(�r�h ��f]抬  �k���v�o��3 "�ͮO��������G?V,�|�H���K X>�9��}<C���Ê�{ue�}ah@�sV�Y�-ѷ��^.Ri֦�)���[����@����CH)6k�sp/������O��\��Dm��-'��?+�gE�+^w�/PÆ��~-r�
�&�x=�]m��jwDִs���x��y�cm��c|�>�.�I�׽�qƴk}F�z'�)P��H3G0�u��h��#�m��������۳�i�����z�s0>�{�̖�Vx�\\jk��=㔞Ã/��v��Ы7��?���D#�+z�lأ����huc�6����G�X�:�m�
v�ki�B�ʆd#�T�c�6�E�c�Ȱ���|ԅ�c�������0�^�xA�����2$����֗��+*��%���F�ʹ��7d�O��q�W{)����|�ß��'~�W��8�+���}��lU��bn�"��]��ak�Ѣ�MC]?R)>b�w4���3�Ӣ��XdF���*ml�pEI`$r�J�~Fe�V�Tĵ�u��+���ȟ��U���)�,{���Q�}s0��,��]��O� �q^c*O��F��mn����1��	��j��R��:�����k���Y�K���)��O���8֣;*Og�L���7f?�u�Ys��p�N9�͇t7��'��+b��*��"~ ���ǲ1���p�kr����uIuc���N��$<�}f6��T}����i��+���E*�g�2�l���H@K�����:�Jh������aa�.��; �|�D@�����Z,%׀i1����o�Ȩ9�����'��k`� �qL��\p�d���>���w�j��-��*q���1p<Z�Q*�X�R �E���Xa���v��X����C�	�B&g���c,..D{��~s ���b�=��?\),�|��{���Zp���e.:��Nvמ�t�Z�|&B΄f�����x��{I���X8W��B������hvX��1"U"�e;G�Œt9���@Ei���c}L��>���Ug�;o!����7�������!�8x����%�Fl̑��wXƸ�׉��8�#c��,�,�{t@��O:�R�� .�H-h@�֎���כ����gttxDo߼���������~�;~��Tԫ��i�+�l�/���Kz�f;,�pR�����f�-���?���hM�C` ����ڽ{�կ��W_?c}Y1\�X�X��^�n*g	 ����]�v�EK����t�(����)��|�S𰩛Uq�Y���W����������?�������=^��;9�T|?�~L[�
�C^�k�Vz�U�4�V4*���?03w}]�%����&��+c���Ĳ߲tg�]�;�mRyV�Y\YP��]6{����Kڬ'F R�ls5z �0�ڭm�H=��`̞î�U���Qm�kmm���xS��Ǩn[�v�5f`zά�����1=
�OhSaޜ�|�6*�_O��\�����TWuæL-D��
�Ki׾��[p��Þ�M�?�ک�rw�a������ˬǸ{8c2�`L�ҷIkާ�1?5��S�����~F���=1��Zs3]��7���ǽ_�b�]/���P����M��`��vb�G�*���q�7�r�$�����y���pt5ذ��ʅ�0��0�)�����-\�u�`��_#��?@Ԣ�.�	������w��!�_\0��T�`��U%``������R��XƵA?��}�p�`O���	�=���ƛW �"�x[m���^�+�~���	���O��[۴��E�������2���c�����	O�����c���A��W0L�H���t���9y��Y��V}��!�c�u�g�l-z���/oxGF8��}�~��A�f�$`�;`�"�$�H#��2��E�|�x�������$):[��G7�;b��|s�e�?�3��O�M��M�ic�HRr�K�,2v{,R�g��kb�j��*����^��F;�9{U�6�w����
]W�XS��m)	IK�"����5�6g�����Oh��N� �8J,lL�X�K�u���~����/��P��𔣱�G~��?8⽶�A]ѿ�����W���Κ��봶�"��j�kA�=��Z.ذ��x�n%`���,�&�Y�������H��!���g�������~�i#̊�a��h_,ġ#�y��Z�E1�a*���`�p�����3�?��:�%�\t���P|��-��NG�E$*����Y<�E�~�h�p�i�� U��\d$\#�Lu�_�eb��_�&���/�k��u�xF3p}��S��;>O�Rīa�342�K�/~��`��m޾��;$ً�~�S|����k��_�>�=�)��	E5@߁��
Z $	20z-Ð��$)L�̠�$�@2��-F���.]��!KC��cv�_!d�=�������	��m!ϝ��Ἠ?�0�����.3s�x�qEbb�՚�	��skk�ms ��Ձa�����u��7p%�S��%c��i�߫���qؗ>@��|��s̲�mZb�0d<�|���M����HC�� "$>�i[�_�fb
�baP�LS��� ��z��|Y�20�{e?��4���ƾ�~|�b)��D�H��XW���¥�Qd�K 2O�g���e���l^$�����m���7D�?�|UD���9c��j2J)��3�� �>��6�g}�L��Lו�m��H5Y�D�r,lҿ�ͯ��#�X/�,���
Kc�/�p~|�G'�{a3���.������?��������_x��5m��䂀 ����ે\������u,2b�(�鈒&gI��L���L�z�7Z]��4~�U���yjJ�^f��)�{�����[z��#�&���3�@e�
��qz_"�)�F�j�zl~�=/����'�ݷ�r$�{��A#���q�h왥�z����ɭ��o���49� ߍ����h��ST�u�J���w�մ3^���&`�o�5�����91�N�9�Ӂ��nc�ϱ6�M?�e?�/_
�C�d5T�����&��)�0_P@`&mX7���|r�'��qN9~�[\��<����<�=�}�&rb��m�tv�O�y%5�@���}J���@�dιF����,V|����`�C��\���ct]W���1ѐ��.�� ��Ǐ���.������R��b�􍘵�G�� DX���Hw�~In[��T��2��zBh�Ϲ��o"S/�;� �ܡ�0�UF_�0��E�D��6��{���O��u���>���.��
�Ɏ�㈾s��	>���G	;�q��_�vLbo)�m:�h|u������$�D�j|<��HF��B9���/������>�y���YOl�������"� ���˼��=���諟���3�5�@\�˫�
X(:4H7-,)�*R�L;��W��<�A{�Y�"mq��=��ޠ��m��d����x���!���РwH������
��*����m�E�B҆z����н�{\0n���U*;R(����.K�N�v��'�&}X36!?���M��@�.��; f���sec'�Ã�}��o\F$E�P�1�p��*e�����JA��A"-ȥ>V^��g���/*XkiZ�{��0���y"j�c�b��*����?3�*�y��y��u��+�6��Q�m��Sf�k�n�k2v<~^�q8hӼ�b<���Ŵ6��|�槯,9�g�y>����dy�Od��+_�?^���e��O����@�.���g�Ʉu^W�	��.���ـ�YS���w��"s819��I��Izs_^�S@ݏ���:�~��;�bP�v+������+Rx��+�=Ø���{�v�&`���L�,��Y�&a63�)�����h�<~6�'ų �j� ���g����`�R
�W�,����ZA�B%9�6�X��+ ��p(�C��4�WVniƣ�KN���X�,�߱z:�Wbd��jVm�FOQf0~����,eٶ��uv:�|_p��*�3�0���<�=�A_/Z=�l%d!���2�#�
�Ϊ���Fs��i+��l����r��E�'�&x�������,`%�'��R
麟�C��7��$��ǋ���ϥYf����|6��U�Ze�����:��)]�4�i�Q+�KKK�\M�ps���������"u����hغ�Mk����}:>8���#�b�hp!`f���(3R�P� z�l(�!7�(|����d��˒��(5>��j�g9�:>̐������sכ�8���3�h /Vx��W�^�w�}��}���q����6X�

y!���4 S�a����$�ac�@�A`4➟��X{���f-f��+¥�^vOܴ7��!h��G�Y=�V�j��C~I��J�綏�e�߿"/V�:����R�����HB��B��#Ǟ|�O�{
QZ�z��6�p�y��(�O�*c�|kʧh�#��H���fZ�w��g�=�\������n,'�z�٘�5b�L:����n�ڞ��3��PMe��f�Xk��>z����J3�sq1�#���6_��N��]0!	��&�C��(���AI �(��`��_�Ajϊ�� �w�ho�Ph�u�*B���@�����������=�0n��l�*���l��0:�nw�_��~,����X�	%,w�n3�>�|���R������ Vlo'�����7 �ES���x��7�� �xq��V�Y��%4����ʢ��\��C�$9�� wٽ��}��}rr�ϒ�	}�xu$��Q�y�$�/>���mnƷ]�����6OJŃ
͜m��ξѴ�s���/>��D�'�O��D��o��Ʋ>��2p��T8��j�jg����&6��J,2��Ԛ- ��
H�#HX��]^]�p~q��5 @+� ���F�z�=fM�/4�U,]@�p-����aj^���?�]��]�귈��0`�\�b�M�ӥ��5@���$��V�*�/uBfǘ>Jk�f<Q����h!�߼yM/_�A����`#��v>>�\���{&}�M��h�$�:���4�"�
.��W�yy�yȆ�a����2�6�,��d�t&�0�)�%�Qq^D�Чɖ�Z��V0}" A��j����Q
V�Kʪ��ˡd'��bt����'�ٺ�Fe"�5V�lW`�t��'�c�����:�s5e��Sk&3o�=��!�MK�̀g�[�p#;q"6qud�Z��n�k������Fo��>`8��#瓱7ڇ���O��ͫ=s��e혱����Zͩ�j3~v��/����0���{�}�'�23KM9��nݥ~[�� N������Aa���2Y%����'���}������*���k=;=�:0�>`)�~��x���CYw�|E�*�q }d�[��������ੂ�`X��~��W�ا +Y� ���M�Je�&9��Uz��ds!���ǂ��b{`rW��ߪ4�K���K�_G�|&[�Jх�}8:>b}i��O�zEK��}Ƶ��+���'|(4#RE� ]�S��o_�#4�j8�1��F��\ʲqm	����Kr<��.ԗ�����vK-�I������wX����袪X����'0���\�+���a��x�&l��|hIͩ�V6�^b8����;�1ad���V�k�ԔMl����:���F{z~Y�,; P�ԛ���(���H�o�t�+�~�3ƴ��Nh~6��4[tu�0��%�ʘ�,t�K�����*�m��I�,:gC�@���	�>[|9T�)b��@G-�Oi���!XZq@3����.�^��Fпׯ^�����7T��gQu�i��i���=y�N�����5�]����[��x���Z��@c���J�f� ۑ0BΗY�WY�)�4Oſ��#��r%Py���:9hU��d����أ������U�D;��{�y�wJ�1C�f�瑵��ed�\3�Ai���|�H�Gm�h��D�����漓:�ퟣ5vr����l�HwX�?��7��̘�������c-F�/G�׎y�q��h�m�9�|��ۘ��`h��ƿ��\xZ�k+��������M�,G�XD^U���u?��Cfgi�f�ȟ����ckK���Y��C�kQ]Z^��s�="�-��� �U�)"3=܏?^��X��5�����==9e,� �h���3��v�v$�@�9��ׁ!��b���}�ymHp�\ e �wWWY���F0X�hJ_�) px5ƿ�� #��Q#}ZL_ ǀm�]��5@ǋ�C��~���y�L���as��D~��M����<Ze��a�%�qNԇ��d�4>M@8�?l�����㱮1���=�C����`���۠/���Vdo��	����tϗ1�`#�}xŲ�J�F�Jz�-��x�Z��T���$�V����Y5�,����e��O�_P��,�c�8��}'��]0CU=9K�K�ʀ����\�Kf]7��o�0���3����:��%��DW�Ы����ۺ:��m����<e;�n �dy�!��V�n%)+�!Yn8�:3�:\kE��J�2�6�!۶�[#K]䜇\�̕j���>7���E6�R)��q�x��&��4�\4�k^�5�x�V�z��|�#L�fޜ�i�^�Y�P�9i���>��S���2�8w�5=>ݘ�"�<���Ӿ>�2���ѣa)��%P�����1��f�e��`VR��^�H?�]dL�/v�m3]ۖLٕR&�Z��nK����5�5������}�q�Dҕ>j�������)7�q?���f��Gw��w��N�W�.%1����-��G�N�O{�l�G6m�����;�$ܹ��G������W\cMF�z�� ��^� Sf �`�VZ�h��2�Qi����<|���wxx@0����[��[[�܇i�
ڳ��7����3!U8�}WLV���� �}��E���b���K��l"����$]ݽs�}a��F�66A2ĕ!����IVt��}�{G�ud҆�����\� ����7���>祧�u��)�4��?K_���!���t��,7Mw�ǝ�$bJ�!�0�0=s�pHEE&6�T�`��ay���!�)\���U׻�aA<v{��9��T�4���̨oN#�K�������k�������Y�#YD��Tߜ�%�mG�o�9A��z�YYr��YH�� 3:'S���o��\9 �c������JP�*Yv9�'����h�gH���0��z`�5�$L<�JX�I(?1�Z#�Ƙ�!$����J�����0Q~�T�M�$ ��$46��N`�'R,��f�k^�os&Me
�������ލ��5n�r���v�<�˔�ۄ�\���U�ǖ���V�����:�"�wv���nv9˝��s�N�\],����0��غ�_�i��*�H�]m���=�(�G5�F_���pA��+��3'�޲��3-�#L%ʮ�
����_�%#쓎\�6���V,e�H&�[K`���|��-�ţ���EC{����wd�Nj�ŁTd��s � ��+�Ъ�߿�<xH3@�'�%��Q֭ĉBy{{�=��=::vgg�|�����8�.�N�� C�� �8����v&l�(�a��`wOtK;�e��2ҭ����e���1b��:9މ��ǹ`�|2���1I�k� '��Ei�n2���������O |,1j���:Ax%�H��\\67���[�v�2A�%�{o���N��'WHp����2�u����}8�xW<(k�7����	1|_b��kv�G��f�$P�R
�������-�3g��1��y�&�}���I lF��ej�q�	b�u�l ��vVl �>�v��,�P��n�n�����Ȍ,�Oymhf��O�4�K��N��t�Ҩ��:]���6C=����Q��p�?������y��/6΂����WҴ�Ҧ�1V��s�� o�aLئYG�\Y�}��4�<f:J�ӳ]�#Id�0|{k�u�=�N�������~}bE'F3���>L<砀�j�� ͧ�{����a�a��X�k���t��9 �%?����b�<g:[�6Q2/��s՘��\d�nf?�k�������M�zf�%����뛝�rM� �%2o5 [���"M�ڽ��3�nZ'+R��7����W9�7u܃��bh�I���3Y�u�Vm����WLק��ݮx�_mo����mcӯ��]pc��{㙺����]���/.>	bB��eF P"��_���/�����{|����D���|�(?{���3�s4Ń<�$�g���
��+r҄nB��T>99#��;Z�6�j�`���Ŀ ��,$, =����QS9�������3�ڡ?6n��x����>�/����X�X�b3i�"b4	�vD��� ���>Auc�a����Ȉ�c�;%���2�J0�õ��`�{M�/�/oXuµ>�\"�}��T�ˏG�"���2�M��+��W�(�&����34�ӌm/c��5��?����rI�w�Rn0�e��Q�a�`�2�]�kB�23���v��B�ZS�9�B)e=�=���h����R�]��+o�l���/�Q>�ڗ^��^r;`5pT2ܵ�ޙ��o�[N��[8�Z#����36�p.��2)��)+�hQ岪��p��)k��V���9y��ƒ)�3��zz��%�H����U��r���se¥���6A$9x͵��0c���b��6���}�9X����̜��^hI��Gl�uuưo}��i;�-�����qk[�0�W�6�Om>������1ļ1�B˶C_L����F!��i�WWז��5G����~K,�l�g+_����_3��ڜ|j��}��kpɤ�x�&s�.�e!�W����0��I)�yȼ���һ�c�$��}b�-�F��*J��iխ jG�!}����| 0�GTJ�;�jB ��{{���z��g���\��-]Q�}z�C6�C\@`��R�!�E��M�7�Ï
$��L��`�4���	���DݨV�W��{�Rl#qE�NN�y<"�w�5D.�gj2�_��%�:�s�� t���e�`6�O���W���^ض���c=??�6k�G��'`����m �Mk�7u�Uc��R�&��K��g|��m��S�M���U�SΦ��Yz���k�c�
$��Nfig��!Y�`iσ�kw�h9>Ҙ��?�,�'���!Jʰ���$9c#
 '�ύ�5jSI�&.0���D@*�n�N�o�3���,�X�L�i��[��:٭C#�ht2ca��`9�xT�(��(GS�|&�N�;��E`'ȎEN�t-}���|�\cI��X����y���F㞆���Ę�w�=��ϙA2�����H�I�@��)n ���� m �����~H�S�;H��+��h�:�sk�+"���]��
��FUAJ�ٝ�Y�Z��z�Zb����l�ʲ�`�Q�/��5˺`Z��EZN	Ցj}׀��c_���Iv�L*]5�o�Ӕ���t�S���2 ��qu�Pb��oH6	J7�.�+G;A�!o���h!�l�w���$�̘���K�����Ǎ7^#��`Os�O������G}�����q��)�f��XH�Hx�{��Lw��h�sa6|}��n9���Ą��P���Z&�wO�O`xkk�m��ruh��||r�  �A� �|�޶����.���{|x�ꅏ��/z̈9�]HZ�=d/ -��ߐ� X,�9 :xJ��V���x���P��ո ĩYp%�[7����pxH?q4����c�������'dk�<0_�7���\� p�g����3�w�����o���m�;�4 b��9 ?U�zI@:�������y��.c��2]֯�-Ǘ<T6�Ga�_�Spx�gaw�{��tݸ3)WTR�@��e��^��T�縿����9�����/ǈL���r|�ȇ�ӏ["�1=Bb(f6����40mza>x,b>.�c��.��l�-o��VF���`J��:2?`�ZV�Q�� T�d��o�λ�R*�F�I�k`]��MQr�f�G>��Q�����3 -�Naj!Vt���0^��\\�F�5�N�#h�u��ԫ��uCS���0�y�Z��i��CId�љ�N� !'Π�JK�(Y�����lXp�סs�	?�����;Oı�.�y4z]}b	�en\����Aʶ�ol�J�x�}9�x��nG��`��a�Nz\�[��T�"y�=[<<��;�H�x:���6��uP[�gP �E [>߮<7?�^���F���X��O��?�9����\3#�Eˎ��-/g������8m;�ٱ�q�'r\�nN�8_������C��}n�����G�V"������3�5t��Y��Â��ɡ7ߖO����/��0��R2l7�7>�	�>$� ��ف̾���.�gX�Xr֤{��[W�O��+G�J��}v�}�>���!��w2���K|3P� ��w�K������m�G !�ƶ��޹[3W�q$������$A�L�T"eXBW|n �h�wrz����`�ݹs�ݻO��緷��I_�#�*��w�����zw?n�b8$�`������C��_��J��J�`�����6�q�����O��E%�c��4/�R����+b�&�|�.����okL��4�����1��+l~h=`�z	��I��07�'+�##�`��,�lHO�C-�����l0'y��+��Q��RڣST*#N�|�̤+��
�v9���)��������߬X�U�Y��b�c�u��k��aW����|Z�2!��<�M�B���+�w{||`���pFu���@C�b)6#��|�=���a�v!.Ȥ��pQ�r%�8mc�J��(�nj�-�u�e@S��9��Xn���g4Z�$���7����� jmL��<g02H�x]��&�C��J�7�yc����Mly���4&����)0A��b6�ohK�1������pR��x��B��8��]�v��p6�=�����N oy�;W�cv9( _�X��WCJ�*�U��T��f -�!Y����RR#5~+�G_�
�TS@mh=+U:�y��y!`��ȯ5�T��_,P��Ӎ���5+�I�TN����igc�\��U㦁�"@l��� 5*���J��ڪd��%��%]�6]ɨE��b� h%ʒ�����sUg	2�o�j��W T�{_��8��� q|��߯��x�@����o��.����9�'�S#�#-����gjer��Ɯ����{�1�~��g��'��t�s�6��K+e���Q�%�s"��!�I�ɴ�����~vM�Θ�˼����tS)�}�ۢl[Zt�~j�~�������N׭>�2J�ǀ�Ҷ�`�_	�# h�4�Q�'Ҹ}uM�Y�_ / ���͙c�6 �J��	uU����v@p�����R��p�� �H�Kl�皈e�Φ۾���=8< @L鍋W+�k�숍�%y6�D�ـ,��C��8%� h�s�����v�jW�C�����g)6�2|��p6%�����2y��.�sl�t�1�6E��uO�V�	�?��B��R:҆�S�)ppK��/mX̤��h���������T�f�/�}j�5MY�RR~��z0�&n���v����3�O�,��;
��V�O�XN����S�����	���,�ٽ��VInTfP�Fc�f���6���!n1�4{me-g^�z�q�;�e��	��V.5��<!:chz�d�K�}��sY�7S>�6�j�N�$�{�٭JM1\�'�fg,݂���A����#�{��O$k�k���2��T�̥�a�W��Gw(~�SMKL���ib���d�e�i�5@�t'�o��5�H��x�l7�`��+�y�~�=uH[���98�VB'���o]�ֹ�Ժ4M��}���a�s1X����|O��uX6�!3QJ���x1pt���mu^/����J��(�l`!@W�Ҿ5�d�Nm]gKN��Wi���Z5����˱2���O�4A4�qˋv借Ś�J�M'��o�d��8���@�d�Dѹڐ�2����(lu�������H �B�О��/���_��-�)n^a'�8-~����N�J둰�%�"0�kBh��e�8�3�B\��Ⱥm��6o3y ���m��_��=+��Λ. ���.'����/��
RQ��{M��� |��^��,��r܆юh��e���:��hp���2��@�Bܤ*��W�42����Ɋ���o����{�Y][Q�V�T >C���4�����+�'<.0�K���%��v5�Q�w�/�>��� �(���B���%P�H8��FU0e��#n�����w��u���yHOHe�pX;�J�F@B�����n��v1/��p�n���S��\��ߵ2:1��!�y�ʕ�� ��ؠ��ǸI`sA��d�nk��o7n�l��3�RF<�G�9�2�#�Q�vK��jɓ�ќ�c��6¤��J���r��!�j���F{9��q��0#H�w���>|BZ�p�l�|�h�+��[��� ���+�b ���z�[�k|�X��-�\ d /�Iw�8��>�����|\��b|�3�����-h��fFW���͊�+j�a�a�!Z��o�J+�x��]��d�=�����⬨�G ��X}�l�f6��ւ%+2���@�Rx�l�<���1�����H_��d���̈́�6ך,(���1������e���ߢtߺ�]J�T*�awve��������ܫ��+͑k=^�_�`x�}V>�Ŝ�����X���g�Ǟ����%ۇ��5�t^8B��n- �/�O�9�⾿�y���Q�{o�ni�>� s<�s�\�jg��7p���r,ǜ�H;x��1�\�O�'�6:��f�Wj�Y�+�����wm���І�?�>ץM��RKP�_ikz��)L�:3]�9���d���t�s�WL�&�Kg��RR`��@�y�jg�6�y��j��δWZ�̾�thT�S(ַ�|��I�����+8����[�o�\d��b)��.���?WN"��m�����7�Ukg��4��}�Zet} �$9�a<��yi����]0�w7},>�q{�_Θ;�j�݉n&M��`� qvv�@�g�@�ml�z��d2X�	bˣG�j��lnl���D������{��;>>%��{rr�Ɣ�-e<m`H#�Y[[g2���u�5ϤŐ8�&�1�t|8'�&��"%!�gk+>�� �%�*��l�] ��|he�h4q��F�ޫ�+���&����7nww� 5bb�"���	�'��~ %��ǹ9���?�t��Α��9����o̮�'-�'[C���0>�5��E�-#��Z��%_�Ҥ��h:o+�gti�ۓu��9�ސ�,���(��q?i��bǼ�����s�o�q��#�ٚ�h��K���	�����c-����-��Jt&�+�n�����V�e.=��5qMBz3�H{��E�)X�^�B�ͱe���ھ��n/��׋,�h]�� �mщ7��-����cNQ�ޔ6�\3��b���Ѝ�uL���s�@(����#�3�|)���f�WV�nm}՝_\H������ 2�!Z]Y%�;Qp�ܖ 
�#��:&�Unvd�'a���כ���������_���sp��K�Z҄#`����h�4(���h�c'��.8f�f��5��w��`xv?%�t��A��{�x��y|�{0i�n�'رM����W?���;o�<����߷��9��2����X�i�vq�;�]>-í�l��Io1������S�~��Bm����C=�Y�+0ϖ��**[/(+S4f�I,yM�l;��6�m�_���ړ��:�r�ޔV�%@�^�j�yc:IX&�1H�B˒�L��޶�o�d��Xe�AY�����FA���j���RMЊU7EI]��D!7��/����J.�A@چ�\>Oxq~77r`;�_r�k����:���|%"��<�%<+��X�<�|�m	�t=�c��]+	� ���:9��L�&�ڗ�)(��.���>��>C�2��E{������Q�}�S�p˵ŧ*@���US�������#�/h0y{k�ݹ��*{���|�R�%��jM���,M�Ve�� ���mnn�"K��D���� l=gAjҶR�ý�}��f���@���޹KR���Isp�O����hY(u�7�I���Ij�N�{���{��s���''�.d>h�;b�+����a�������)�,�՛Ԁ��k����0��k�,�/b�"�Z&�]�;]�M��[۹��'�m���T��J2��LO�+x��9�چ?V��k��x�1���EdX���b��D�\��p{RƲd:\I]�Ʒ
V�oO`H��Ӯ;cҩ7kwj�Q0P���R p����t��M�9�hZ���Pi7��]��T�J�J}1�����Θ|��/�.�Ќ�o��ma���m0�|� K�Pdɩ��W]��d�Vp8��`��Ϣ�c�קcFT��b���`24h�
x�W@0��*K�8���R0�_GK�f�5?�t[����ݾks�������t�*��P�{��y%>O���`?�<շ�o)n;���FC�b����E`p�M3v o|�{�]8v��Dy\����h�S�3�n��,ǂ!�Z�r��l��N�N��PyL'�'0��14���Tlz�Q#)�i_��	4!�3.���`�G9������,��~<V��	���$��Zv^CP�}7m�v�MXؓ~#́�?ؙ$t.U�`���0�zr|L�Au�6K�U��fh�Y�`;[�vUJ]�Ϥ�  ����'>�5� �q-4�Y�hU�A�ּJ����?��8J ?���h6����tO����M߿_��
�����dğs-��v�g�Uw�޽����fN�o?Z��� P�rx�'���%9�ׯ���s �F؉Uk=��M�M����}��c��� ���ɍ�2�QRnUs�^V) wtzĹC.�Q���zz��� Kf�r��!�j'ڀ+e�U&PH�u��n����B��i��.��omo�F!g�-����Q<��,��U2��Q&��O���.�9������/�=�|���&�%k�.@�����'���I0��G{ {�xjee���,��`$g�ÓS���O�f@/�,�xN�QO�>q�~�-����'�˘�0��80ڏ�-i|����W���XU��A2�I��*Jq^�?�[wⱜ�颀ˏ��=|�P��*�4'U��?_��(�6]V����}��8�5��0����𸣾@�]�M�2a^��c�����[6���^ǧ��TE�`(���༷o�߉q�h'|pgs���>]�2�3���+X��9���>h�ۭ����>s<&�^������b�ʩ���!��2�*L�8uu0�],���P���P���D~3����~�sW�$�gcmm�m��8���#8�RJ��2��s�;b�M|t|�1E(�\-��9_(�{/c�Ӌkf��\Y�݂�s_G@���v�"�IP���g� ��e�,�>+v/�ܷd��з�i�iM��v���^��%I�\_��� p��/{+_���l����ӑ���׻$e�F~�u �c��]~ߥD|9~�k�m� ��+�2��x��Ᏹ�VW��\�:Ұѽ���؎�AҎ;��4���"����Wԗ�tRS��F��m� ��cǳז��T�щ����;>>rG�'�a߷��D�Q˔���`�
�h������z�%kE<~Р�bA�����������Ç��Ǐ	D`P�������9ˉkc�i�0��y�NI �%Mg̋%����}2ڌ���H�[$V�\�:|4\Z�OD�ޓ!�: � �E�*K-���kcc�W`�9=��s5P�t��6�r��iu�	�3�9�s9S.~���-��C2�l�s�=����
$ՠ��uF#.\s�ˤu�z&t�0�v �}��5�PD�8����LtR�C���N���B�0�-�}��d{Λ袂y�k$������^+��2���׫yy��X�O;�8E�ix��9��YG�e�7$�;x�p�q̨�ޓ.s��=>����}~&~O�[C��m�'II��	��Xm6Fg�(k̗M��C^�{��8;���o�|o��9=9���K��)���>�2�>c�X�h�zT�NF\K��B�k�7��1g���%y|�6>��� �x��7�%��"O�}�&��T��:w�cԒ��sUK�D�R�Bcw��~������K��D#I��\io��}L�S� ����H>�6�}����,~�^v��X���Xv��c�s!�<���0�4~��'��=摾�.� �m,����i撰we�*�~��"�߲�u�ȄF��d�4�,�?���F����p�'R	F���r�%�%�۬Az?S<��qdy	�6s�k��r�.V�/�7H,s� ����{�
�Ch�!g�8:��d'sH5�Ss�����6�f�>��W
Z�h�e|@6s�s<f�vu��5f���s}��	e��ˡ�)r�y.��ך����-�:�ͽ�s�+?��O0P�dX��D�� �|�2����~~������~�~eѡ̏I.��[�ٰ�w���9�/Zw����`B��e�{9�&�뽽]���+�� pd��;����n��}�`՛��[6v������{������]� Ұ.�G��V7�5�;et�4�i�ݾ�? A-�'�JF����o����t��m��߃�$����}~�2�t_	�5'|���_��4J�ќ�ڟ��WO�r�Nz�߼�u�z����v66�Ek2��{�8�>>:f�� �"7�ρ)p�X��;U^O���f8"��S�۝��xl�Yg3�;��U-��]U��g%قRP�� /v޼q�_�f�'0j��n'�r�8}��+w��6�I������>��`]E�)%J��m�N��y��}_j�I�'@f{�mG��:�� �=�q4�J�%�������:~'�O�'Zn�K�	�\�/^��a�b,��F`d�5������7�~+Rs��fϞ7�$0���Q�K*6����>,�\��\��帕�������PK[�եHDY�,<��z��o:=��e7>/�L��l��/	U�:�+ K�\���Q����0� �R���d����dBӚϰL�F����t���␎:�~�xLWz����3xo�C����H�σ�|1nx1b�0��;�lf��n��z�s"�z}�ƹ�����hC�=����x��	��r>d�E�_��x.��XC�m�-Cr��딫+��s�{1�Bpe����|K��ȘiX\;}�׹[�?�X(��r����&'��ǭ�m��ԫ?�،�T���R��x�+Z�Q���*���G@0aV>u����q��u�Y�	��Z�3�H6������e���)��� �s5�O/���xߴ@��P���J���,�b_��^�U�8�y�G��z���&pnlp���!�F ,���hFgPPmN�F�/�Z�z�sL���k#�<_�6�5� 9^����s��lN�P#�7��ӱ�x�|���t�J ���M���ϗg�����%{$�ˮ���؏E���g.y;������G��$��b,jPν~ҹ�:�����wn�,Ǎ��P �}��9A>����D�.$�_�f#����w#���C������֓hC���/!h��ڂN bH�M�f���T����k�I��#԰ɰ�Ϟ=cPNF��H�6T�M��=zt�<x� � 5J�Ǔ���2��d���]$J�������х퀥�y1[΀{x�%�ݴv�6j���������ۦ>2%�$�� �����������l�c����+���� {��N�k񏎢c�e ೱ ��]��Ƕv߼��⼰-^��q���\�����$u}����4�S�Α�d6�W�`�O�7���	���V�|��B��7�¾�к���Z���4��������@"sW��8�1�X�Vp<�����ru�5�(�`L#M�o�db� �p�/�ɶ���3߉M����7�(4�Z];!K]e�,��
�0��:	dƳfw��ԅ��gU$;�R��*�Y�z<�Ë3��O?1������ht�d~����za�`�`�a��� 	�����Y��T.B��gZ$#�)���a?�VX�5b2�F{��X'� ��%^��p�s���y F@�d����M�:3�3�,��N�'���="P�9�4A�KH*�LRux�h�'�����`"W%q��s`Dc���ի�<|�$K?~��s��-���6|��mG2J22EL
kO&��j��[�^M�3��0}�#��>�\B�'���^o�T��a�	��[%3�Gݯܯ�N2�2~��+'��aF���4���7#��脟]���
�����5�6�Mm߸�#`�
���U��U����f��Ұ�@L�����@'��Ē��Kמ��"��^���r�6By��8V��Bv�� 
%�Gd	X'�])][�,�5�۸���x!Yₖ{	0!7oq�:����>:��.ug6D����(���*�\�v����mTi���!3M�E)�{����i�>cߜ�C�F�4���I��x(��ԇ���~����^n�цb{��uw^ /z�|��_�����;�m^��٬���z#��N�_�8.������4\�-�rHi=�T 	*��!���V�v�-���7d~��	U��Л[	�-�v����#6�yg�!H �E�O���e�p<�wv�^(�l��\�� �����V��F����H��ݹs�%����4���4�[+ �a?��s �c l����X�l�� ��;Q�Њ���9cjY�ь�EB�_���(c�1`�|`nM�	8�T�ԋ���K�4�1��@��q$�B�,8����Y.������Zq��Ɓ 9 Xc�����z��ZMM�]]|�������b����d������/�?	 ��@S���A�r_� "�	TU�m9K�-����$[H�(4�q_�J �������loI I�/ TRz�I2/� ��	��Y�[=�[�E( pYY���O� N��N a�2����e�9A�v�7 A�Q�y�@��oW�3��ܡ�k�*ǾGp5tS5_��)N16s0�?p������)�&�C2��gM�*m�Ã���0�/`��>��pm��l��SJU���a��X�p~�1�������%����g)�����Ӎ�ڥ�G��4$9F\+l�w��X�F��&��q���,'��"Ϟ�۝Б�&�=���XT[(J�#���X���V�`탌�2��pU���4�d��<��y�5�:��~ɑ�Qjc\�;A�X}��N�*�*�г�L�b�70��'g.O�O��>�?uG���h~����� ��� �*�B#��Ewc����pw��p1���'n}s�Q\ޕA�Xǀ�.:�rX���37�?��z=g��7h��u�M�<� ��0�o�_�wdfV �����7o��Ύc �!]�W�=����O�u
�A��Z�z��5vv��My4��z<�.�ͮ��}n�A5Y��5 `I�#+ױb6~�{�����&-8�<sæI�i�w��t|V�d���g+\�y�.Yr%_/��Hw�Ԧ�����3H���@����j:g$��6}i\/E��;�|��skRz�N����r�=�˱��YH�z�J��_G����T�E���F�]&�PH���B����y���`U] �����+������#?�X�D�M�X����j�F!9��S;R�S K��Z]���B�M����_��k���*e���0��`�}*z�<�錊 ����9LDIq�S֨��B �b�AF�%<� ��0� �ϛ��Bwxo��u��6'���sl�^GBr86�K�S��S]�#ai�J��ݞ2�8��5�F x�  w�C@Lr�R���V��k�z���]�u���ۣ�Cȕqe?�-��'�Q*��`�4��������[eT��0ч� ��?�S�����x�;��ڤ�`z�X���ܱ�a%��X?�o4Ԣ�̑0W"���2`����r4�S\S�����y�Rt�jŹ��y�r,��8r�VQM��'_?�3�=q �"Ea�i{;��G��|�=���s#��"�g�[؛�V���m".�ݗ���J15�\��l�,`�Õ�1�%��� ��[�����`}�
!i*h=���h�`��F��������ׅ���<. ���m�:��YE�պ6DE���'�}�q#f���-L
G{Xi���o\��w6}��s����N��#�񅏏�%y7T:w�t
�¥j*3��3KG�ז��r\9$y����O�ǭ��x��?��~���S���}Q��LSI�������1�:V�����]�	$zj+"���:�O�>u������4�ُ,4��.N�B|N�����wWX�����ź	��� m,�S���"�V��k3f6�b���p�oӐ�e�ע?���*�X��ڢ&�S2XmpD&	�1W��Ƞ��a�QT�Ї ��t��"aP��Ȱ��M�[J�F��oʿ��_E������ZV��|�%Y��P��3�5�L��@
c��V�`j$,؞�-�f���a�Z *N��&qa��O�V? �dO��w��2p�=o�t����S�3ݦ�����*~���E�[��9��}�G{�1t_}�0��A*q��=@�����4���@_�� ����>n�A�;|��5��vrb��z�c�G�8���p2�h�e�{4w���/fI
6�F������c`v�Q�� !�(/��	 aO�Nk�c[8~|�@	�j�Aqi%,U�ν�o#%�����y���E<�F�54��q���,���G'�����kq�Cf+@4~3����Y -&cP���s���=����,>c������z}/n7�����4 � ����ָ �5�bYw��@�V4پ�"�Țl@����H�R.� �*�nb�� ��&aq��7��	P^�~$���w������{���� lA0����g���+&$ �� ������+�D�_���{��0$e�b�`4&c���h�''�_ȋ5r��~�-�r|~#�$D��B�I�9�y �b����"���m}|��*ʲ�;X� qoͽ���msM`�A���n6�6����޲�'�:'�d�ޙܒiF'��-HS�ϊ�	��BI	����}�j�!�4������Ul�CHLM��^|f��7ڤ��0�����(�s�c�ZY*�r��m��]G�JHXe[O���t����r|�!�%�:$�	`,�+������d�]��}�C)� ��x�ǲ| >�0�n��� �3IB�ߘ��.��bO>���c�/�TR�Ԟ8���tTC��Jqv��3���� �`��l0�}�q��t�߈�3�e8�Ȯ�%���߻��oc��� |n{�{�)?���g����;�8q'Gg\�W�W�ĵ�3�����1S��֜o�A�[��
,Z�0�����Jp�8�+?��L@d���M�wsn����JUp�Hf�������\��lƧ�" kQfr��O�a`�9�t�4.S�f�HٳO@0�������C��'f89'1�# �ch���O �n,����T����_`os4H��-1�C���vD7�����J����I1�l�OM3ڻ�N�2q:�鞒y�Vc
hM���Be�t�gV�̑���t\�|��o�x�69�y;O�����龘���#N�?�v\��(7��Q��s,`?��!i�"��:���(@�'O�*۪J�A�7y��L�6���B���u��ѣ�R�Q_`-�$�U�l	�w6iw��c�|.��]bHZ�����gj�gFË#0���3�� X1@�F"ٰi,Ӑ5r�VX�ܖ�v� p{5�5l4h�J���R=�j�4S���l~�M�1i�O|~v.����Pуy�9ֵ0���-�6�߳� :��Fâ<L�H��s��8wi�Tq������Ǐ�!a��`4Py��;>>�� ��2؍�#0�ш
`'��H�0�P�I��*_Y�x����t V�"9��
~7���䳔�N۷م��'Ղ;܇�B/�&��#�`�$��O�*�OY�ޓ��`9�S���6��b�qn��jlЮ�ٌd7�)�]i`�O#�չܯz�����i}\���ԫv˱�~�'�&9:c!Ko�|{k�]�[�nO��uE�K�Ȑ5J��Y���Ց�z����&�KI�5��7%i���w���~,$�R��A���d:�����L�r>I5�����T�Ͷ睸��Z"ƻ}6�u�&�7W�m�{���҃`
W�JI;Z����k�'�1.FE������g���B6��$,c�:�-W>^Ce2s=�j�($7�5Gui[���m���Y"��D��!�D�Eե�M,
�<��f��^�gu�|����#��q����y�ǡ�G��\9'7�|��Z�0�	.���K_�lO�M�!\�&�I^ 4��ӶB�>�O m���,4�=b��DJH{qZ��n�ͳ}��s���?^�7�7KG��w��{t��{�ࡻ��>J�0cы���ڦ[_�p=��Ώ�׶�c���"�<tO����i�s;?����������w�nu����+6��b�F=���S����M�`�O���<�lܥ���N��aR0�qY����_u[�fn�w��W�z��A~j���S�a��4|\������v�|Ӹ������9_��w�L�{w#:y}:��"`jD�D2
� xjޣ�Y�t��`��'�T�D8(n��z}4mZ���8q{������1�T�YXg]'>m�=>,��^�`�5HT�6ӏ�1L�� ���)J��&��n/0�r���x0�Ѧ���}��Cv
�x�0�?�5��ly�	����ٲF��Գ4���_�F�\��|<7v����A�T�;��0�mH�����rd�?�1=p�����=ك0��[�~\�b�S D�tz�����ƺ�ꫧ��Eb�� �F��Rp�+lȤ&�H��}��~{�����6v`&��G��7�����æ�ɋ��c� �1����o���f�&U�}�ۺ{� �4���2<� \���p� �
�ˆ� ���]�eN|b���L&�Ջ$�` le2��2p��\a� �B"I�ݽ}��z�� e�9T�Hbݪb�H;Md�͌�:kj�m���f�����EJTP�ǈ�d}��5�=h���@�[�� ၵ���c���>:�k�9�>��ς��u=~���94�[��Sd!5_ye�{��	i�%`E�# .��L���1�q��z܆0��J'JqM��@!�圱��
W0D� `T3a>���w�o��*�}R&,��������o�9 ��ObɔnO�����dH��~�'"!V�D�6tyV SX�ٚ��%���Z�m�L�����ftV�BiV�HU*$0ೲ:��TP+C�,宰e�1�����YG�*f���١}2���j�`[���~��YkP��� x��
�DZ=  ��IDAT�ֹ�'0�J܍��O\��?x>��ؼU�p�%���j�{��"���ފ�*#�&?!v�X���B��IP��ٌ��ͨ$���<Y�������c��jx�6�#m܋��f�=�M�����c�LR��"�%��㕰"@����2˱o9\�Ib�?Q��G��
�g�o����!CFG��i�ǈa�#�,������Ĥ����ݓ��b�)qP�������/@���{��}���xi��}�~A6��kk��g��r���S ���MW���_�gϞ����r�;1=��bsM�������ԉ�,:���"HC#>,f/_�t�ovc�������O�6���d@c�&P���mw�~�����-��r�;<ޓr!6��dHa�G fy�Se\*�kas��"Ӟp!�l-)�K�U>�>��b��ۋQy��P��H �XQ+���\�S��qE+���ju:�y��؏͛0nK�O�ƉI`3�V.�Ӌ��_=}J&JS���+	O<�߳��]���P9�Z�ai|u������É�s�6=&��R�Q�u�X��ó�sw��7oR7�թCi9�j́=Q����/ ���Y	�^�?�w�7�����/���:Ik��i���z)p���~S��Jk�G�7����[��\�1���`I#7�X��`'�m��@P������ �h�M���"OE�4����`��i�.���^���Xϫ�sl�s��d@$y���$��y��I�ޫT�}�k��j��D�i8�iL���5��jl,|vӀol+��	� l�nj�X�L>AO�C��wW�A0�+l+^��}�� �0�����6g �\^�,������X�΍6�s��4o�0�߫��h�%ՍFC94|���}��F`]w�?��fS]
C6���N��K���o��:�z$1��+'��} 4��|-^��J�	V�t�QPb���l���o�f��\K��r�\^Ѵn�J�"1�F�I_���1��%=�is��mc�����M�x?(;N0�gzǙ0@��M�Ef�K	/cb{g�3^[�k���`�'�u>��l��*U/�r\{�}(������e�%����d���e p�u��;���A������V�`=BmM[�A���c�/�1>��*���8�Tx`-A�����imr"���A����hM]�a'q&�g���I��N��=h$["Jb����ho�ثF��|UV
�� ����M�
�K� �Mb�C2���	�N��zܠ�v`2l���^TE���k�yيk"^8��g��o�/���B�9&�hF,櫥EZ��3̗�C�����#d��4a�HSC���\��?�{�29�f��#��t�?���8�c�o�>��C���e���}%7��X�x�w��4P�(���g�m#B���V�>���,m�i	&XP�d{���?���ݳ����/�s��bH�E��{��1(�b9-��$ �(p���32�'����e�o�j���;�p���'O����v��7�/��ۺ��v�w�qD�bϝO���Y��F?������|g01gvp9����3���cp����P!���vE^��s��Gb`����3���r�l��U��$,��|\�Ll�Y!��k),�3j�9����ɾBC��Xڭ��gB��ri�2� ���/_�7;oT>$��
ˈW�o
&}�u+��!؉�%p�������CL�`���}Z��\�����a�N��"P6��/����~>���M/Bn<8�	��^׹�4��<J;|/�[�k�ȿͰYPi"�'�K���&�Rr�]Ꙍ���,�SqM|��W�7��Tv��[��8LDjG����1����lmm��.�[��MI V�&�Tc'������(0�B�1�کJ�����G�]V���Ht�E�퐙�ڿ �)1�Հ
���H�v2��+���K��,�=ǄԀr�ʎs�q��  -�h�:�'���50���	�5�`i
�qK�bvH��Z��I�^�<s=����f@�}x!�[��H���H-L=�c8,L�J�k�Au����Q7��h��OƜ�R�� �1��`YX��m����!��FQ�Ӓ}�'��+��]�%���&�ω6�r�v���r�X�^���܌���Y"��\C���P��$��iTB�#`\�l��ғ��-�!��SG�|�N%M��q�$f,	_Q�{���x߮o�%�$�����?Ǒ���SKXe%Ć��/�{؋�2פ���ت]3������k�{{1�0�W�Դ�dZOm1�3����+��+m�KG��Lc]Fr. 9I������4�����:`ūW K���ѣ�c��}�ɸR�Ϫcp&[�U"�%� }�$%�R�Q-�
*eM�~W*��۬������qN?8���Z	+ix�
�̖�4)�=~̘
�s8�:͖c����$=�?�񁗡y�!��f/��ژ�wn�6M���k\�D��Rb��Uq�s��SkBmA�����yy��	�e_���h�H��.5���{�m[�V�r|6�V��^,��� �d�����������������R^�B~�Ζ�Xߤ@P,:�h������v��Nvw�ŉ��6��������q�&��p��P��s��?~χ������������?<p���r�����v����۾�A}gjOՙ���	Jm1�,G��$mZ�6�80z�K"��ţH2�Vޫ���A�%8Qк��?�s���-���>a����K�4RF�9.�p����ʇ ��v�4�&�U��d����+2�����JW�����T1���[�OY���x������y۽���'|N ߉�.�L(�W��A2؀��L��z챑�~�+��/�w�~�-H��	.Y�����a:�2;.����g۽��=	R2@\�c�U>����:�ֿ|���`�2�;������>���޽��x��ڟ� �u,�U&���S�(zd'!�g����``�w�52��Ԛ���8�>~�R=mv�j�:��ԝlj��lZ�2N�a%��v��0m�j��d�������u��QM;&�!� ���]�!#vq��%� v���%�Le����dM� �ʳ�3-��؀H4?D����F���)�O��	J��$U�XF�]���� ��d�QB$��8�1Yb�U��E�@'A��'����ǉc�����>������
N`;+dϭ&�`��6a4�J��q?`���_E��9XBf'̢�$>Ñ�\+س�G��r#��׵U2����AlX g�I+L@v��8ρ6�{L<[ p$.�us��	� �Pمჰ�+�PB��1�<��2;S�O�>�M�rN �pxO��"k? �A�0��Ǎ�	?��VJ�,�r|���L���%=��?�@;61�������n�嵢P�~��Ĭ�ۨ�r�����3��c2Y�s �6<�c}^a�֕U,�ή�E���3*6�#���4���@��PI�5&�A�C��NZ�?�`0�XN�&K&��_�z��cϹ��=$E1,+ T��xM�VZ�S7%�8F���x���L`��__�q��ǹ��la�HSB;j�u�6�$�p�VX���u����W����n�iU.-��g���]��l��h\W��$�T^��+|�A��d.⹷=�J{JaX���]擤��;*�D�q�h��>�y�F�~�0�u��E����O3-\�~��r-��Iڸzt�ß�_����K:�u��q����G9ю���R��ѲCH_���%NR.T�y	��xA�E�m��)&1(;⢍ߣz��-�߬�G�I��������<d�{E��]�?e	f�j�mI�Z2�����Â�������E����J��ϭDHN@ry��/7l\!�� ��e�?��W:!pl���4��2�������̣8����&���ȿ�l8�`#�|������?�@Ƒ�cVZ֊a�*�f�4Re���%i`�	���c�(��C��M�%����}I���P�@j�/_����q.P�g��M�������~W>e�g��ҸΙJ+,��N�+A�b> ]�#U8���قgn�S�ٗ�`��]|o�����S��{�}8�v��N��sV$���C	_9�����;�6l��ݎ5��$��Sf�IVa"�#uJ0v����!�E�㆝��z*)1NL^��}i����EWye�(S���eB�*W��,P؞�͑�N��nt���i�G}N��C�
����$��s�~�i~�j�0ЦQ��[�u��ٌ���X�LVkT8����KG~xp�$+�6�X1����#�� @�����H ���g�{ 0�/��E�$�`�X��(�}�y�܅��
"I,�_����ac��a��1�}�3�{4Lij�y���V�t���*�տ�F�H�0��h=z� ,���}�&�H�������&�X�G	�Pz�dR&�����%��Ƌ<w�l�k'��G�ɚd��ɉtX��5!R��*⦇I�TA��M�и�3��0o��p-�lI�G���a���_�����|�	�e���ɮ�̏��Y�*�1k��$_o�S�a��L�ƻI���7�8K��لM��ˤݪ�`�f��&����G+�4ΰgN$�.�<,�$k�)��Z"�$s�J�ćms� �U%��O�T!ȳoMi�֠6��fL�2�)7����T��\����&� ��FI�,0.�v��.&��F�/l=�9B$�0�{��WX��M�?Hr�:��1�5�ͷZ��?�Ѧ��5�c:��(�j�}7��=?��e�rҬ:{Bh��<�s������	�J|E��Mf��I�%���-1��hh⡅y�����K� X~_�'���6��x]٩3�i���w�vi{� ;~���?�����?Fg����6V[[� �&:���^���.�}Y��ʀ�x�8�T?y�H,�X<pl�D�����:�C�\K(�3d]1�����������MtLN܋%(������H���0(��rnZc��H��7�a�7�u����H�V1߀*�t�-�m��I. ����W����܏?�����f��� H� L�(����Pn꬇4�����<����΢Ӷ���}�=����=TƄ�����RcYl�۾�\�ݘb���������?���b�'O����o)VN�e����-h/[�a��j��w��1�ח/_��������t�㳄���?ķ�F��US��:�Vb4�Y*�ϛGi�yp�:���~Ȓ �Y��ҲG2�}i{�~�2�ss� X>�v.�.����s����?_fR�smM�Rbd�6����7pؖc�0�K:����,�܃��c:�ql'
�C��:݊�a����#�uw��(�kjWu&�$���l5�'G�n7�b�.6���`_�u�=�3TI˺%K��u�
�7�HT�]	�n0�'mdz;����`4`"Xg�Q+ �i�"yg ���K�lIN
�Z�j�>�s�(->>c�U�a��t�aHc�&X2R�t��`]�g�����+a0Ogg�Dp��;z� n B\І�$��(�ZA:���&��x�H7���T�Y	yDF�	��<`��ml 8O��l ����#iHK�/�z{d-K����J����~���N������X*G��D�V?����W�M)��`.�3U���@nBFuS2�����lA��F��$�=b���.(���ư��{v�����S�r��dz��M�\>�q�/�U�Viu���Ϻ��{n����gg)���g|}]�¦�F�4����3�rL�'X�x.(�2��Aٮ����}�F��}������Q>2|���c��Cvnh0p���G��S��I<u|���l�$~�Úpz*@1��6,Eb	6,d��8>>LIKګ�$��D���8�>ǵ�ܓ�b,i���`iwU2C~�l�$��N�F���&��5�>/�x�k3���{�$���?�1��i����M�:�k�s�:&�&�v,�4i���&�,��B���N�-�Xɤ)����c�\�H��ϔ]Z�<���32�,Wn���w�,ˍ���-h���ٲ%�k
F�������?�j/��s��gy�~��Kw�w�&Cd����� ��?��ъ;=��Ra[V^N07���?��������p�����/.T�K�K-{�����Y`!��q�����w������w�?�/������������p��OY���-�n�@�6&��g��[6�u1�T��s�i���D� h�Z���/~���~����z!�� �.�:8b!i	C*;=�����,M�(8r��J�1>	��믿r�����o���l2��W�����钫�/����J�5`�v��������/d�e�s����� �Vs��!3����p��fG�=��َ;@l �p��$��W���oZ�m0-�ːv1,��;��R�me͉�"��3�Z�ܾ6�E&#�u���8Ĥ���R`0'��DY��f<n]�+m�X�1�(V�9���رɱv�n*�����{(BP[>���&=�!I�:i�Nmb��1��-�͇%���׍]�>]?��lgd�O��P@�X��^�J`-���9��~��u{�~Z����@�)k��ή��`m@��lʌ�v�O��>J:j��[�e"S�g�� �?����JS'�N���m|�X�����A��X�:�l��AAB�h��sz=i؆�����C8�#ב�}�dP��A�m�$I�Dh��9��s���4MЄc #��y�E��ٜ+ێͪvhU+�lK��r%��IK��,���Z��d.���������� �$.^�z���L(b�����#X���5����?�͉궶�1Z��K��W����Eb��'@"�#�o+��G�6�$�9嵄u�&M�u]tE�;eYp�l�(q�j-k�{�I��xVh3l�G8>9�u

� ��|S�;��(�.	�����ۼ�/�qZCl���SB�ev�%�FC�Gl��H�rm\=��
�~��޼�u�)��R��I۴/xv�2?�m���M7U��0��[Oc>WAdj��|,�%'HapN�'~,� �*Od��U�Θ}�D�h�aa���]�x��a�Þ*�B�a�I���&�d=W[�;�j��(*<X�AY�J讈����5����~�XV���oO��:&���H�f�i/l&�5$�66M?io�c�0���wI��jޘ�^\XЃL�հ7W��W��`�J-�Cj�g��FD*ϦI��+��c��q�M��v����r�"�� �����L��
b(�a\F�T��-M�:� M&�{���^<���HƷߍ��寿���{��腍gX�*��ņ7�i�#/����<��m�O�s�5h9��E�D�@��XM�y��/v鄿�i�=�+�	:�U��������c	�q
ʃ��f5^t�L�v�lvi*Dv�34���A���\5Q55s֞?{�j������Rb�&8���d�����gk�����=�(c�{�������[��~pO�<fP�F8T��Eɇ)V��;B׸~>.� ��p��|��ܣO�>q���{�?+Ik��Q0���U���Ά4��U���x�,,���ݸOo�k���tL|������J�ke��K�J�W�����W���Xd؞�_P����	�����c�i*�fifW4Dר�ޓ�6\�y.�B��h#��!�� N��t��	���A9�$5f�$�Cf��Y�:\\6{^�T��)�E��Ț�iϑ{��rݧ�QQc�vr�3��A���a30nl�IA7���a��L���k����jT�r>�k	tssl��?�L|Z}ʆAX��s�Ji�5>�u��K���R�Q ɾb�H��5~�ަ%��Ya6H�%9`@bɁ:%��،�M�4��U%P���н�ݥ���ޢm �Pe� �%�(:����1�d��<=�k�����qc����+��5��P�l�}֒��pp�c3@���+]/XnT�K�b�h��jI����ǩ�vo�7��h=�a�6�V����[��u��k��,*�e 2�S ���y4������5�OȊ0��v�I�H�k� u֤��5��PH �x4�hڤvYA��/	�Z��3�)V��O� +q�R�jɇ��#\�T�@��6L{�C��G6r>&���J+��R�bv!��#`s`k`'0�I�� �E�9|N@�s���Z�ϴ�pgc0��D��%3IZx�1��Kc��~1D��犥�U��D&���RYc����1YE	'�-��j�T�\oU��5w�M���E; �<���^0��k'���`�o�y��q�gA�����5�Ś+:ѕ�w�����iP��Y���^.}>�2�h�g=���ch�/غ]%��mZ�:��.c�������RY��HnժϪG'�P)��_��q�#�}��un��ȶ�by3n:,���"�$�����W�t==;�*����`�����TWc�SiL��Y�22�T�>ߍ���������=�,o�E���[p�������?������������O�_���q?=��wn� z��`�tm὎)��bF��g���4��=x��?���Y���'�T��+�=�je�&��!��q
�/�Cjm_(+ac����o~���W�t���� ����gDwx���X�����\�k\F8d+�������4��������{w��}wtx@VVf�V�D ������ec�~��\�����b��G��������K��߉^�&�\nP>0AJ�������G�&V��F5Z���ͮ�*;̀�;w�Pkb�b$'"�������Ҵ��`?n{�  l�<V,3�wO$YȬ�FU�d��O �`	J4q�0��ݢV5��V-����Uj����fg�=�,5���q�{�l�\s������Q�W �%̳ܓ����I�l����}����1����dh�R�]���O'�K��x^^��.��w������c���KGZ$��|�p�筴�RJ�N��LՑ���˫a+�Ds�	� :�
K����A7�U ��gȉŜ�3�p>`kp�w�o (H�c��XEH2�����&(�H�"�����7��C�8����=�$�U�U'��5���jZﴜ�Y����g#��soU�r ��9=;��4J`)�0�=��g@�i����2H�I&�um0�xW�:e	�8O b��!;ﲾT<W+����\�u�1�a,C��x��'q�S��{��?'��dt*Wz|��U	�[TXPu����i2����	���|�܈�^�Y��P�5���p�b��}3�;���z���`���Z�����(|4�� ����7Y�6̪*p?#Aԅ��x@�~D��6Okb'�
�&�Xć�~�@�U!]��dj�5��˼R����.)CW��WRS>�A�/F�08�璊U���{����P���X�i�%�����R{���J%߻	���RՐ5�5Hr0�B�t��6`�U����R3m�2�l��&�#�gk�J؊��O���L*���ي����`%���\�O�lL��y�����[log�wHL���9�.� �+�'�6��V�*�T�t��i��E����X.ť������bqM?]d�Ň��at�z��v^�ý��HNܝ�-w��#��w�v�?��F/ɘٌ��,]�	����x�n��2�����J� %PO��ӧ��#���?�)��!�s�������;�_4��y����UJ��~��������{��Ft�#���f�^�yz���4�&;r����;J'��' �\����q;1�F0��ӹ�C�,�b���,�"��^����!��}��t.��g	7�ra;�zR~�{d"�rs��GH?�y�ٰ���I��vD �Ϟ��C����W���:>>u�ӫ���z�+i�a�p��]���{��n5i�T��%�Nt׾��k��O�c|^�{����4��轝9�����6���t��K�����z���F ��ؕ󋉻���aϭ�bCχ���k�*���ˬ0ʂ�`�ov�0�����w`A�} �J��=�R���R�|�8㊉�����0�G��XxHRu*a��w� A�������>���z�Z�w�r�V N����j�q{����j+�OIb!�>??q�{o� ��*�W��~�����o��& �i�F{�	l�&��Q�B�nG4x0 �{��q\�7��P7��,�BEm~�j�æ�/6_���G�X�H0މ����"gZ�����A�=��f�$�)�1_3=cY����6)�[��=z�� ���:a���H*�����vl����)}��/�,o��h~�WO�l�zvͤ7���}"�e�� �H"�	�t����K<$F�&���C�͍�o�d����ʌ3���f~֬L�2�)�&�H�a?�ǄU�hgP�==?eb�WO��#;N����Z4���X�Թ���"�h�p7W�Hc	������M8&kQ�ָ%D�%j�D�5�� �/Z�� �L
V��`.p/[p��ѧ`�+��� ��	�K���\��d��4|>��b�8�dćcj/�I҄�JkTG��������\� �M�sȚ�W��'�j�QyĎ�4��oZ�*Ơ��
�3�c�8�HB�F�^G�6��5�^��}UUs��t�h��h��c�,%2� �B��;Y�Ht�ENJ�2��5)+z�b_X�ו������Ĺ��Jbg��elU�hd
��i�l����\�����T]l~xi�_�:�z�ҧ]�O2|�_��3u����lR��� �IO�ש2�q�%]e��c��\�?������=2�H^�5<` �{�,R z^� ����<.n�q�� �|��㸨Ay"��ܡ���
y'T�����PR���#�p �=y�(
4@���֫�, +��$HW^8��Cwz6�67�խ��8��h��|��G'�Vv_�S#��i���%c�!�"S@	40~��!K� B�z���켊N�)��zR��U���'�� ʼ6��E�9l�ѣ�񞺟L:g����9d��0�N�B�s��\��ag����g��A�����s� �	 �:�Gñ��g%q��aqdb�Y�J�(�7��g
���"����EC*������45�(�v�h�}����"y��O��܉��8m��͒�Q+r(��0lC�ǐr�|���.� �� *�4�6� M�BM� ���|�{�{^p�X��c�E#���#8�d�����mZzr��kA����q\�ps��}r*�7$]*h��������-}����Fû/�<�y��,����:�{H�Z�xkw��7_��n��2�30�i�N%�HT~f7�3ݰ�V%�u`���r���J�*W��S�x)����*Yo  � ��c±"3U!���4�H{�&}V5��!�����#��deNt;�'
+ iZ�dAw�Y!m�H�P�A���C��o��
`րi�'�+$�X�E�e� i���zdH
�ssI�Ø�ܐ�����ɏ��F4�ɝ��=��F��^�	�� D��&oAP����T�	sC������T:K�߷�7kgk�OٴKl���+�N�����T��\��Z��E���k	��c�GZ�����^]�G֠yD�Ҳ��% rHbf�K��}�sf�O��<|�8��K�@��:e���f���Y���h�N�*E�G��k׮�+ξ-���L��>�3=�}�xӛ���X5��|&n��>z}~�V��ĤEr+L8k�F�GV���P�ق.]��ـ�d�<��u����51��Ա"���hi��J�^�|E&[B
�S�l�����%�0���?؋�a<gEC����v�eׄf �kX/~�,�S
>ᵾe�6M�!���񽬾���G�x���I��'���j�uԻ��2�9�"�XJ���V^���{�g�a�h�ءAbk�2uI,)]�R�}�aRغil�D3A�	k,e�d��ڬݤMZJ�5���D��IY椰����<
j~������*�P*��d�<��غ?k�j�9����"o"�`,P۬�h���m��;�n����u������4�n�H�D��nl�n�{��Uň�Ɔ�N�9S�y����8t�;;��?>�Q���k���>���/�5'w�N�"u͠	L������˝�M��o�Rz��ء?(:6��ݴѡ��)i���,ԇ��/~y�O�B���a�9��:G�a�$�C��3�� bQ,g�s�!��������,��e�&1n�\���z�Υ�#��57/E�`��A��ɽ8o߹���Ê��F�Հ۫)��W]Nic܁c�cx? ���g�+[[���|�gV�Cq�\N��FN�h+l��:�>}&O�<a1��X��G1����g �,��>+r��Ν�8ܸ�ڍ*����<_�']c�R�b+X	��*��XS��Z�Ws�Kg�!��՚�|�a\� [,16j?����*�����am#Ɓ���	���M��rG��@^[�ϩ���6�/e9
�a��>�w��� ��9�w����:��:{�YŐ�5�c�4`?���C��Ra�=|��2 M}`P7��K���W[����a��\YhI>��Bqd�vT����������Pu��s�Zcp Җ�U)��Ct�sK4��9�@��%�:~o+���Q�v����@�붻c�����0	��xñTZB��麩��f�4q�6���^f�e�r8�~��K�i����>�)8Af$��!?�z�:��ѵ�$FX�N�n� 8��U�D f��"�YIh ���!� �g�iz��5�9}�PV+�,<Kۘ����1�U��H�����k��!~�,붃b�t�������'e2y֛j��[Z4��,��wy+B��G�*�kg)R�$�{�kj�f3��]j���x���|�4ٱ6(!`ނr}���W�-��,�F.1��8��N h]6-~�+�+��Y�����kX��b&c���Ag��
���s�0��@��]c�*lj -�}ȟ!���:ȋ}�/�Q�Oً����׋�U�&�"���:&�W��*-_tn��~8Ϊ"��O=H���z)v<�+�}/`��{��X�	j��㹱�scYc/β6�9�^0��πE��kd�:����U���kV۳T��Um�Y��+Z򉫗*q��_��:yJ%7�i��\6"Z���s��m��ʍd�u5H�� ��Y���+,��&��6	�x��U?����q�1Tވ���:�y�d����ӧ���˸��3ՠ��'�[�u�a�D�z���f�$�J�Tc���)�=�AP��׮�Z__az��?�dow��X^��ez�`�[(���3t����O���s�Y @{���ݕ_}�O,V$a {�O�kA�M_x�<�I��!-��E[�EJբ�Q��h:��h���h���F�C�κ�nZo�n�H<4���f��F�Q�z��&a�NR�:���-u0}T�E�� s���Uh����]*c��c�
��q O���k\[۔�w��d�H\� $�E3�Kْ�{Z}S�dt>����2wf�X��Ln�وse/Շd��H�ޛ>o�/�
�c�S�K~ ps��Y���ȍg�`�L���IV��@#i�p�i�J./�_�0���B��;4�!�������n0�1όE�珧;���
�	�[L7�Љl�R5i����%��gЌ��[zO@R#�2�ޓ���w���X=�&:ٞ��ގk䛌���{��$Ȧ�	#�M9���W�{.�[<�j9��w��Bb�<Z2��:�s@0��G*���.�C��@@6C*p�$��FvG|�"Rp�q��j<�z��G2�_A���r먴6h=�3λ<������W�����T�RL?S���2��{�+�؏#�g����,|���uUGyh��d�(�Q��_��$=GΠ%��L�(�1������V��v�SQ#u������lb�6��$�onނnU�+����w�v+M�� X$��o�uIF,�o�Xp�drU��J[ �V�Y�łc#���tG�� �j+kQVj��U�:��s�
���	Q��	��</���'���L�	c�*��{1�o -Cʦ��k��������=�T�bH�}'ۯ�Py�d؅=�؅�ˌ���b�~=��O-{/p���d�<]=1sg���>��s�� 1�W�uF�y�S�Bp��H��!�u	�f��Ou�b݁o�,12�s�� ��<b��N�$,pB��f����be)���"@b�\Y�|�"�^t�e,��3@���7�!a�Y1j�uAB������z\��pM�TFG3( k`3O���z��a��kk@j���Ht���&T�7��`v��i�;KhD����ʲZ�}(����}��{fx����'\7�}�e� 1��Z�-������=�+j*��'y�s���[o�=lҠ�y�e�VN��'Kd�]�5�,��_*;?7������W>��cL�D�)��g�~��3 ������<��Ry�'���&��6�ƿ��F����~�+'�g|�r��dye3n���`����Dl6�0�jf�%v"#T��N't�����G���Ɂs��j������j�+k��I�������Kp8F+��r�;���ei�i���!�t���L>��WJV&����Fk�2z�uPyu�"��i�e���B0G�s�/x5z���|ڙ�29T0b<U�Y�)�(�U��Ek+x�`�:��`l�"�ljL���=��Ց�� ��������s{K51�}��u��^)��;�y*��¨��H�UFǦ��$�k�2�)0���]�_��m* om/�b��� k�
�>>�|�a�te<�R��`�eyA`}�ӿ�X����I<�i�a6����=��]�j��<���A�@/ /Ju��X����״Jgt�j���|wl��Crv�E!9���k(�ˎ;�1Ng�����
P)��YvH}q}��7e�zY��c�����6E.�㿽�vժ�.^��\���9#�R�+�$0��e6<a��[�d��]J�x�IY$��`3!����u�% . �`<#�T��F�u��s�8���u��~�@�Ҁm�[P�5$v�4P+Mg�E��� K���g�c@۞����\�anN��v��)i3�`�P�g(�H�%y�
c��!c`�`_�4�����4��za%g����������IK���,�]$�5��~�sB��\�c.�gV�ϙ�E�G��f>�a�w�y�V�{ ,xc�+3�d�\;���u�Í����`S�1.:���+�����/����s���p�6��V+>S����|�짡��k�?e��쉲�;Z�7W�eO)W�Ԯi���ʬH�-�H׵�G_0nQ��{��N/�u���,��1����� i�6����Ce*������4�2�-�g:M�AD�t*��s��rI2�rh�q<#������K_�Q����> V.lB���Ú��	=�	�����\��R�o���^�]�]32�u�}�!`�,�7����Ќ�$��hSd��Z@i�2P*9˼��n��5n{J�����T��A������!XVM�kN��^�Aڢ*"� ~�a�Y{���kwxj�;�'IYLki��q�u'j�MV�����~wI4��}N\���j��z��]hᒿ.��ΙtϺ���O����PZ�v���&�����䈊..��.��Ӵ�v�A:��{6�4z��ݳ�3y��{�e�(�bEx���]f����r:��"��AA�<���{z%0�p�?��,����;d�ˁ���C�q�wx5I �4���8�Q����zt�cwz,�1rǎ�-㏪n�k��L��Y���[U=v�M�����	ق`Lmn�%� h����ZW�pًQ����j �%��s`.,,�6����#�$pp[�,������vL.Ae �� ��`���.�<�����,+���Ӊ�)�`s�����D���h4����	��j�����-�r�m�}8�+k�$��{���6YԺn�S���vk��W�*�0<=�8iX5�����J�N܁3�@�2��$��Ec�������j��G���mJho�1v[t��������	�+(&�,*���2�>��`B��2I�Ob��(%�l��fq^ ��<��/~![q.B�̰�dUքo0���γ�tY�,�@;�I���@Pg0� /�� ڼ�D���hDS	�Jk ���m{ż�� ^�w ��u�� �1l�ͦ�����Ӷ)g�����xO�E14� �A!�����3 ΝY�{����������U�O�D0�(3e��c�a}��z�E1�td�ѦJt`<����T'ݺ74R�@z�+�lY�G�M���VХ�`���O�_5e�@?�Ш�,�	�$����Bp��7�Q���VC7�)tTF0��Ǹ��� �1F�Q��+�h��.�b�`��w�H�)ZuX��0���{��S-�.��؟qɐ��}�O(��R)ôw�ڬ��1Ϭ2Ϋ.3F�tX;ep�>�� ���T�\�O�^N9�6�LS���y�݉s�Q��ܶ`_S��1�<��9��e�����k��zI�>X��"��=��	>^ �Q�Cy-C�����o(-���kE���}��b���>�5��'g<���ɶ�\Q\�<��u	7������p%\/![x�g��]J.��M����Y���d��v�ɶ�y�J��fT䘑��<έ������3����S'J$n�8KZFפY�x�X�ЮZ��w�Tk�5S���4��37��4��ވ��y�U߰�umC0��ddj;يnn`/�>��������6t��	N�!j[��4Њڦo����[j���(Z�X�W�j��B�>ّ�b��da]#��pr�_*ļβ�µ������m� ���5;Ϗ�cW���: z�Q�$�)���'P?��e(�Sm��^�zY���a�z�K˫Ѱ�4Qc^䩯�[(l�,�F����B��l�ϵ�c�G��L��{{'L�C0ʙ}~ӯP����@1@8�x�-; �ܹs�Le8��sE �`�����t��� �	c �v��A� u�UW���laQ���ݽ]%�8��n�yh�e�y�l|�\o�q>(Ѝ�-X*d*�gk��X�`ķ�}�is���e����+��UOg�k��Ѥ��-W�����v��>���e�u�S>}��:1����� f�@�^%*�@T��lN?S�t}�A��KV�0ˀ2	 EZ>�P�����-
�kV��D�v|��"k$����@����>����*���N�eZ����l�gCJc�6���u�؋@��T��X������=�<y����P��@1j	t�]:� �E
�8�,�^8��ӹi�:+\��@R�_Y�B��=ǵ؁ ����/�;��� �V�^Q��t���83[��RJ��6o�NӞ恂aO�<������%_bF2i~�;�۪S��F������\ه,`���~�%��>2����eY��\���h�b<���y �`��Bp@�n<��l'�}�Rk!�P/���C� ���x��=�N�L�Y���qL���@Ŭ���h���{�B 0Ԣ�n�$_p�( ��C}=H5j�J]k�Y�~z���Ș�π�dY8�l��O*S���b����s���:�$o �&�隷�f{��^-�U�`�b�����ܖ��k@.�D��l	����TPT��ϋ��(�AXp\�֫�]ӄn�n�!2�_ʸ��������_����'�Ѹ~��w��9�O����w�^������gN��=��Yc#u]�M�rGhi���M�e8A+�CU��Ap�ݭ$,�l�����-/�6kC�H���諬��I����)¨�� ��5i5��Ad���)�]2,�?o�`�3��tU=n��
^�тS���sD�.8EH�X���N'Ae��$��i0��2-��"eU���љ�����]YZ��;��B��� Ig\�C�ݘr#K�"���Ң�1'7X�@���E��/���5}rems��W9�䈪GJ:���N*˥E�1B�L���F4ǋ�O�v�m�C�����! k�(��5����%��k��oX�(x]t�a�������|�~iQ��أ7ؐK�L�q�^���ʳ`������S�^�
�
uM��@���s}@��Ω�����i���Ϭ�T���A�,����Q�]ӓ�W�\N��t��=`uo��|=��P3j&�����$2��Y��k}b<�1�{�5���J�w����/�Q��2�ڜ�/^�$��L,��RL̏���C�`2�-�7X� �E�V0	�8�сE��f;~��٤�{�3�*U���C��O9,��tN���2�t�z�E,������SK�C��y�6]�Q��{��5
K��8Ю�����>�nƵz��
��X3vwv��k16MG�u � 4�0v�8���öi\6�]���}M��v�K
~g�>�Cp��c-ıx�3������k��4U;���Zy��eWNN�	�p`݃ƸW?��	U�X��u�;�Ҟ'~��E��~kV�j�Dƞ1\�@h���w�.K����9~���x���_���A��±�N�{r|���΋ ��봓H���z�|��~R�jUbr0%Al���4�J�w���Ǿ8k?S������|�"3����<{��vF����r�ɞy]j�������qM����2�48��Y��i�E2c.00t��a�}^Zv��Km���*�{���M#��!f�*I�.D�o��Z�`��o0���0R,�@./�]ֲi��������	 ���R.j���b;�R�5T�i�k���Gp\�a�;(��b�½±�G@F�%|p���[̾����{C�2kY���gn���q�k��pBHA�4ot�f`�%�\Fc�A����uj��r�8����MFf��l�<u��&�^�+{,����S�٢�I���ӂq�k(�c����Bؐ��h�Ґ��z$���O�����o���<��1��G����`�Me�b�=�NXfN#@h�X �Z�n�@��j�3�]E�ޮ�;����;tH��Oms��S�.XmQ}��O�}���BV��*ou���R]�AI������!��TQ5݊�o�EQ��� 4褭��� p��-�ծǂ�zv~,��W������o���\ük4���`�#p|̢1@Dg�z�eן��$R5b��1���*?H�s]��� TWPDh�+˹�T_7jYT/���(8��"��4�/�Ҁ������A�m�1�Ă��s+��N�<?/�g� �b�Q�N-�����~h�+mTI���?����WV�B���Wo͍�W�v����$�w��1Ǟ?{�TZ�&sQ��o���0�s�5���f�
�g�(!����4��
P��}7�?0%� ��11 ���@���)�X�;��Xǜ_.{0���o��������+�����Ll�X����ߏ׀�e4 ���X�~{�@dӣdQ_'�s�p���·�a��I��W ����<y"O�=M5<[D�qe{�ĵ�u�omޒgϟq�S��#M��"O^dNu|V(.���%>��Ay�y>�o����~�u*G�M��,����B� �3�Tm�̸gx�xn�pj�7��$&^wZ�u�]H����������#jd�ZM]�V��Kcd���[|{���*�ad�h�d�c`$6\�\�L���烝~'�~`�� ��۷n�����|�H��Ҩ����e�c��,���5M�{�D���P����R�#���q�u���)�
�<�.,	�Fy����_��q`��y���O��֍���ζg��\밞a��]&[^���s�2�o��X��� ��kق.�c�2��I�F�
�¿̂��+0޲?q<����Xx�G�5�2�E9������!�W�:2-r������L�	炽��k&�w�_ �Q �-k��&�"Eo}=��T�������ڼ�P%�B�@��\#O)I鈟C0I�n�5�e3�V{g�,���Ih����Oi�4��M�F���Y����4�Pe��R!c���r~֏NR��5�e9$����r���ܺ�7�3��0��y���iDq�޼�%�f��O?}ȟ;[w��73�$f�vv�U'p �A�<Zu<��,��8��FA�����c�4��!��|�p��3K�Gq�EЭ�=�04�O�轹b�T���T$yg�����p	��Ľ/M��*b�#�ib�Vd��ʐ�Q9���j,�S_/���8��.b���W�(�M��0�`,�MS�������$�V�9�l4Z*�=:�щ=���>����9��\�ZhwrR�N������\Y�  ��7yl������| 5\J&\:��4E\�T�$l�Z�k0(���7=O�	VV�Xw("� NH�ü
�A���u`���k��
�ɔ�l�un ���Z�*ݱα���2E��J�{�Ј�8F�<WV�1@ݔ�h)[��:�ƞ��_}y�����)ޤ�?�A}�!\���ӛ�����yq[�o!{ٌ ���i�7�e�¶+�d�¹�K�I���e FT^�ԥ�k�_,��.F�~iI�] ��y�-�c`_u{�ъ�Ќ���Օ�x)�`$��O��E5q+��7�#��"���w�!Kׯ�S}� ��6�Nҹ���x�h��Y�kF��%<��=2���
�*嶨:O��s�Ip�]S��]E���U���u �`g����C~Li�}׾��,	ӣ��
|$ƿ��00��$C�
p|����U0��Պ:��vK
c���u�LOg8Bn���*�	+����CKg���t��__[�ײ�A�T�'�L��5>�3�:v�jg�;�'���g�C ^����8o��|O� �x�wpY�H��Ա�i�~�V~��ۙ����42@S��mr����(��jOԳ�8B�z����,ӺH������IG���@#�n��|��61�c`*�,lM��a/��uj�"��}���s���=�mH���.��u)OD�_r�fS�e��t@0L����D?B,h�+|�2��O�_��,�3|�®���TP1,LBC��^�g�ς��3��χ�|��~�g��G��X��x��O$�X�Ũ:՚3�޺�E0RCӲ
�8�����*ێ�oY�ʡv\�ʅ�����Zgf������2[��5�@elB�\{&�F��P�::oŪ���n�l�t�������ܽwK�������k�!=����Z���?�����G�>���k��7������hԃ!Ҋ��0:eA�����<}���g�!K�P�p�$ڌ�1�3�e�R��_ؘ�!������M�կ���'9������G9��n���t�=�D��t�N�!9˯�t�h=҇����('�:��/,(������ ��!�ۙ��4ĆV�i�x~p�a�L�
F `x-96�����ގ��둪�zo��ӉZGS��b~b�cJ_4�zGً״�{$�`ǰH�W�����iaQ�I�X�`�-�xҴ�	j���`��y?��]���gr E��k@V���&�"���ȺTӏ\P�eT���^�g Tvg��dVܨp�D��9���$��X7�\�ʉHzhh��R] �OŠG�b+�	�P{��q��Gt�+��)�2�E�����P��}����1��6HDm=T�0iP�j��Ql��2	�3�M��ܥ�n
zj.�wCAN�����t
;Y��h�d�/� 6��X{�LY]G�iF�P\����l�q��D���X� S�&����.��`py�9�a�������a��9��Wp/�~�Zb��
8�����;��L�zOP$��õ�/�_�`��X.�'�E�o܋,["��ln�@e] �z�A�������aŶ|MC�~��_2��c{keZ��,F�? �U2�W� Ȃ��ؼ��4j�JJض����s��߀GƵ���qƾ�tt��{���>���ѓ�	�)���O?%� G�c�Y�,�ʽ��dwg�cL��a�"����5���k��H�K�j �,Vj�WV�W���rPM2#�hZ;��Ӭ��#�"�r�hu�^�q�+iÙ�e���mM(-��Վ����H��%���� �`j�M"�Ub���)��vw��	ha�`�z��f����jcM'�%�&�G��fB�u���xtH�%5J��C��^�����)��D��h�����tE�LdPk`�
����k�/5Lnc@���<d<��=��u^|V�J� x��r�O<kg��\���&6�g�y�Y�/��s���sfdԁ?�g5R��9���̘)*��M�O���f��{��Y`������^���,�h�)U�+0{�;P$E+Q��������_�ٳ'��:U�;h�=&��.w��_L'�Af�
@��_n��7_�M�<�J�w���#.�G�����*{�M#�����|a��n6Q��-�L�G*#S|re4��_��N�F~��p�H9�H�MfuH@����!2���@��6u��+H�c
�d�ٽ�(xI��2�w�$C���_pX)���# �q�N,@jj J�q��^���X�!�l�F�0��: 3w�Z�Б|{aul|0|�ڼdX ĝ�fs� D9b�׏4\	ܖ�I�R��F���NO��9\&��U�܈��yVJ]� �`W��O����jQ�r�]gZS��ؓ Rh���xf*4�qƎ*PY�B�pd�/gU����U�/df5 ��Q�+��E>�`@*���.��%Ӭ�ӣLEI�����$�6d*&�w���[��4��s�i�k���ʞ�Ri$��:GmI���r���YX�ɜNV�>wss�������l�\i�I�a��,h!��w�h�|$0�j��E�!�p+{<$A0'*߽{WVVW4�Wd�P)����+֬0������v�D�M]C������^���5 � ���Ap%k��p���z���)��x��g{&�M�A @S��T�
k
(ފ�r�K�Mz��Ҫ��ǻȾܽw�vٴgX�%1n`'x��α6�^��ЌV{lX9C�Ad����<]�ϰ�!֜@<H��Y��tX�n>��qV�3���4�������㝇M���2��zh�5�8�H5G�<�� �[�����ϥV2��K4�	 <R�o�V������뛵��ʱ?�V����(��6�
��q�*���)�W�s/ڼ��%e�k��Xվ��2n���m9�˧��j��?x�;F$�����������w�!#����Ϟ��-��$`�4N�
��}M�"����q��tL'��H⚶��j���G�q�<1{}�/uV��FMu�O�[������|���9d��S�P�h{{��!Qc��Yy��X���
*;�ȋ��?Ҽ��]^8�YJ}�o=� �X�{g�c�c}�1����l�f��;,O�(EP�ɟ��<��U�;���f�V0r�r�o���qρ�q�m5sN��C��o_���� @D������GtL���G�u{�����rz�l��}y��)�b�n,��Y���s�!�Kg�X8�$���޽�<}�p���ad�ޑt{��ؖ�ΐ�h��M�V ruM������.�q)o� %Ѻ.�������{�d����,JNC�a��"����iag2��|S�1LKe�ǂk^���F�4�W���Q�4�:v��73�j�	���q���@V��d�-h�T�ab�U�� EY{65��?6�!i���i��O��:�nX+4y�C�4D/2�����s�C�-r3�+�׊j��޻�W���L�LX0!CF�Vk���}���,��Ց���^��k��1/���A�Pf�y���j=���b[}:P�4>�z6�T����Vm�7�n��/�����Ŵ([���:��A ����Ip`]�R�?��o�m�i��1>5���g�����L����$���sR��n/���-������m�Ƶ`}�v+������u������kLb�8�2VW)�`��b�8�W9p��� ���`�'���#��>���:��L��J�8��+Zd	v�i$�=����f�P�R�ɸF
8t���d#_�8:�-����@��?������tv���� ������g�/��y�o2o��A��O�	�l19�`���Q��R�B��1�]��^|�~pA�f���޿D6r�6*��Q4lI�H	*,�g��VsI?[k	,�c���]K���0������j50�ټ�Y����#ٿTv;e������#�VP�ڨ���������:�{�������E&G�����۾k�Ό�N�

RΦ�����}}l�-��=��`8ÿ-�r$+�֙V�i�$!��	��#�!���Zl�Ȟ�4�VY\fQ��;,�jlrf���w����=�0���k�C��k���3-#w�fJ���T�Գ�fkЬ��V9��=؟�_���M̤���kV=�m�2�'�"�	���gK�Q�`�Y� �$��l���;,ߤYڌm�#�r��cꕰ����4)k�����ٜ�����I��Iz��0�sj��'��ۓ����*���l�n�4�O?��ܹs����䫯����C��<|��)�=�N�|��7��}Hn~��I�b7��jj�Z0�77o���;�]����~��Ĺ�DA ��,�r�T^��9��y����g�:��M|5ñ(���`81E+:���0A�C:�f�h�\0:�^� N�^�yZ�.�_g���DN�lsSS�1>�Vh�$@����X�e��#��h�gt���w����T�g5���y��jvv�e����'���dg*�Y/�4�ܰG�̙��V9[j kU�[�`�u�;x$E9��[ALO�kZz]��ֲ��d4�8�O~��Ͷ]���Z�[���Xд����j�W��JS�~�v�B��"��5�Z׼��-H��Y�HIP@t��30�L�9,\�h�xgQ?h���&��Y{k-�7��w�lLe!�ؘ����&;3� 4jV��4��W�l�G E�8-��o.G�Bm�:sZ�_sr��=���EgAEH+,Z��
 0�Vp�!O�z�!1O�\�'��;w�7 C�V������w���A"�aQ&���o�*�k�����Odr֮3��ydb |/fXV,;<���2��cXs�4>���Aخ	Ei���� ��7�� �=���9-��{}�0���Ǒ��C���ܿ�@`��y@+t<�q�8&���������ҊR�=	�@�V��B;�Uio��Ӂu�,���`�n|.$���^��\3�A�y :.��W�~�_��9����x`.z�Z�)��1�9k�qsP���*RM�K؃���s�N����Jk�GԸ�Q�ع��}��z��V�3�o����3
m��6�d�@%d�����˗/����¿�ڀ/��3e�X�l�ho��[ڒ��l�o��O��d�1㱋b@��l� @�fSח���·�^�}{J�W	���kGF�x;�M�������x��Һ �4k��ƚ�i�ԉX�ǒ�0?�"k�q�Ʊ:�d�!�����
A� &瓥���^'!��&d�f�C�'�KG��6���7��D
R����dQ@3nq~Q�H�`*/P����/���,����B�	P!�^|��������h��ߝ����o�jȈ*6k�޾�E�,�Vt�k���4�������e��-:��T�Z�E����꥚���^}�0��c��m���C��3�9S���z���(���� <�>ctDy�s3�<
�~X+N���c,�2���q��xH�:gA��G ��y2����e5&zf��_���!T?�cl.-��%M�#����]�Z��7,����z1Xv@Y筣�B��o�E�����op� ��&}��x��E��sl0e��
d;@.�u�
���A���Qh,�e�D�'t"1i�HdN0F�V#��ް��Bc'�`Y�K�k���kY� =�y+9SV:�|�ۋ�E(	��bR��#�Qw��HS�,�a��d�`ON�kVO��5�:@S�e&����ֹ�c#�2��s����PJ	� �j~��
����TP���%O��%h�CU|:�m���������@�,[��C�iH�6*U��ځ�z�q��Hq�)�EnLp� J�����ƴ���=VsS![��T3T�Ա���RiӇ������xg�J�����%x�s�m�%�u7h�1֒nK���f��]"I� ������9���*3����9Sp��rR���=���p[DB&�U��_�F��D9G{uٻY��7ٰ��'�^�i+W��c*�Q��u�2�B��#ԁ��YWi�r�γ[�A9������gTt�����I���ɀ*�͋K�&�0��������#����|

���aC�GC�ﶮ"�J���֨@2�E74���M�M�-+~���;��2k��n"Z�7c�H���uH�������ߴ6r���l�~9�c���nЕ2����3��#�9�1#B)A���ͮ����P[�4@�f'������X�#�Oۀetӽ0Y b�v�0iIF�K�g"���S�ݤa+��)�Z�`aaN�ݻ�
� S��v�&{NGK��erQ`owW5 ���n�Mԋ�,-.\γ*���eܴi�d*����A����	4�Y�������O�������ɏԓ�6��{[�j.�E$�F���ޣ�������F.W�P'͜]·�2Uӽp���6A6��OC�GAh8u` H@085�:��2$^d��O� 4J�|m5��P��!�P�OUЁ<s�r�!f:Y^Y��w��]cK�A[}����1vC���v�2c IǔLk���/R7ilCvB�7�*s]�������ZQOѱ��3����#���t���=jkE�@pA&rV^n�'���8�F�L-����i��s�\�Y���zqi�"1��Zi��
c�y�iPU�`095# �o�,K �
V��3��T�	�L�73I��q�v�ʰ�hM��h�|�bkd)Yz^j�����Njg�����hc���qSZ`��F������˃�u-JeD��ꊡ���L����&���:��:��b}mu�cA9K6$�lQ�i��{ڦ�2���21su�-p�}ۜjL7r�4��}�Z�q	�@��-%s\NcR��[��s�4	�] �Ǎ�t3��s�N�[�u�ר�7f`���7�t��ϱ4г��o������+�����,�dՍ_'��}��1�<�ln�;#��R�J����C�L���RRh�jQy/?�$9���4�$�>�jY1a��//�R���3k��[���3�೵�؂-����Yh6^Q�L>�j�j6b��:H]Ir�ڰV��A�?T��� ���$s�5��b�Ff���|Z1|�'8�L[���-ڦ�R�.��A�8��^��������V�R���9P xo��pi�a1LlK%@4R�DdIP��k�X2�����/���\�74�5����ZS�!)RFE]��2��M���I+\��x7Gu�g�&-��`�)�I���~}������d����G��Mm=����pC�Ծ@.�d%�bblo�y��l<�B~�^��0n��Fϻ�~>`9ԴZB
�T�e�?c<����Ѫ��Qc�$X?F;�������-,rSJ]�Y������w�gqb�(����;dH�x��lo?���Si7oI���Ÿ�sYY]���՛*5�����)F�gH�mS�n��نd�r�Y�?�U���/���~G�*@kTg?=?�FÉ�x�L�?{��\������~���]�~y*�}���w$o�R�yo�@~���H{��~�Fd���o�b%1D{��F����*����6�ʱ��9���P����<�G0���\g��ʜ�{�YQ��Xe}(d�c| �kH��G��x�NU1X\��0��2雝�u��x�>�C��;>.\��v���e�qA�-����ϑ1���ܢ,����9���nb��>S׍Nh9^A�W���jXef`����"����{���e��/��\F�����<o��x�`2"-σ 4���y�i���k�;O���B3�Y|fԥF*_P�5�{d�_d��Vi�� ��(���,���؃�y�Ч�3�2���ـkb�_\W��5`.C�F:�F�� �qN΍B)=�v�fA¼a��4�0}̽�+Ŭ��65�e��xK�3/���`(�k�c�Z+��B
������;��뎬I�8TX�i�*�n x<�禌�Bm��t�	g�Q�4LڏK`G٫�Z�:�j⇜�������<�1q�7J�4�Ŵh��z2�{~���V �����x|?��X]��V�V���b%�9R)%���Q�h�A��^ך��+���p����s�aI�2���-?�,d㘓d�.|���!�v�Y{m�}Z��ν��0Wy�/^0����dJ}MI�ƚ��,�����=Pw�o6��0�������m���I�I`��C�6A�����!����o��d�*�Z�K��O�$���>��y�,I�I����r�ҲrfYRϹۗ��;�y�3H��8x<�V/�=t-|ؚ!�A`��A�þ����ǘ�o���B>�f��#k�>[�2/�j��d�𭜳��Z��]x�{
k����$�0�[:ᾇ+_[���ҵ+�a��T6���r%L��$����Ի�Ɛ{�ND!,԰=�_G��Y{��;!�1յ�G1�Й'��ޟ��3�O23e�i
_�@����/4i0@�)<�֜�Z|&k�Fq �6*k1�����8n�HG:;9���EeGS_J����GQr�=����}��|��17M�����6A杝���a, |^[_`�a4 z�ɣOd����=��ׂ>����+�.`���
/H��K�w��nl>�\`Ey�0�ZF h6�T���1�Q@���0i���������b�V��t�S.1dM_��m��77�Z��rM�.����~��&ԶÔFhr^ �imd��A�p�ju%�P������ؐ�<���g��#kEG���|�R犢��8�����K��o�=�>VVV�D���k��`���8	�.���fJ"�l��G��ڱ��xUl�Gc�5���#��}c
�E�S��R��q���.���ǀ�F>���c�թX�~x1&�C���8(���4KNUHA=���Y���޲�n�Fz��K�P}����F\��E�Mq��q& �)%���U�.��P[�+�BY����}
adݜz����/W����;ֹ/(����k��Q�W���	���ʊ	>޲Q�e���I���NX���qR͑�-�/�e�	x��U�4��~4v�ߨ����`b����*&�7��6k��zƘ���?l����Q��r1�q�=X2!��d�=���a��_\J4��L�e��/_���
?�aY�H�Y�LG+i��.C������5d��\�EYZV�����d���j7�K�j��i��w�ɳ*0y#���[AA`���s�
_�,�W��{���B~�����<ȸDɅ���ğay@�0�G=�1�(�����[+��C4�v��n^sh��K�Y��<��^g1SfK<{�����6��	�2��E��� �dW����.�wX��^?�\��[?�L��Ɯ	�I� �n�Zպ�4��D%.���pYL�GEG0[��O�ӑ�ဌc�+΢�@8��XO��m�t���>��Er�!~��7��/���)������'��d����ܐ����<y���ڒ��?~.�E������t�1�`��2S��~�z 4�Ể�t�v�L�TnŘ��/E�D��tO-�RfVL"'C�J��8tC&�>rM�1��¹��8��ޕyj*�I��g[���&?���qi���B46��y�aZ�e��f�!o򞰨\ѷ���7�����U�Dӆ����>A��1E�M;���$@4�A5��	��p"��s^��ZP�jh�Ӌ�b	B�/BZm{H��!Y(pe�5�`�!�mԏ�t����,%���}�"+`ү��ҩPI�R�2L�3l/�1�u���~�CG4ž T�^6�н^a�Ԃ$����u5���Χ�9p�FJ���<k7n7�e+�E��\��t}k�J[�ͦ7ڞFֺpq\g^�D��'�W9����k�����n��k�:�QSP�I�0	 �����ݠ�I�rʽ	�\q��0k�RK���w�3��`���2�䦁���	�8�+&��T�h#�[Q��>Upֿ��P&E� �jq�V* ����80x������K�[��l�KQ��穏��7$݉2j��3s+�w�t��p"L��U��SZ�`u$�]���E�T0�P�5d�]�v�M�1��)ܯe���:� �Y{{�������}�Vٽc���"FQT`2}�R3\�s�����ɦլ}���k��攽�������>�I�y�YQ�V��t�"�v)�9��� e����۲ykCN��Tu��b*�8�����{� si�qS�����,��|t�.���o~�Nޯ��F^�x�j櫫krxp��*0"sKKX^Z�N�#��d޾�!��O�?��'�ⅴ�3�կ���fK��|&���Iv���5A��3�������3\�ޥ��ᳯYo�],���J�e�[fed�����ѠC�\���I���V�b�q90݇E���A���+�Za�8j�˫���>Wl.�̌2���X`1*�(jHy��u�)�zV0NZ���_��^N7F���/Jb�q����R��'(��˿磁�H07����Bt�g�9\?�X/hf:�L)���@㉱�M�Le}.����{���K&0�K;�ǧr��=����5�C�tý�=:8 c�����PC�} �`Oo���(����N�ʠ�����:�}�XĘ�����x�g�����2A�^J�jQ���0S��L�i��Y��Y����~*;{�1߿v��5n����`�%SO흵Y{_[*����YX0���v;���x����K�Ud�2�Θ���Oӱ����*�4O�V��&����{��,-/��8H��`��z%��!�ٱ^Z��HŶ�oE_Ã�5�OHD�5�uQ�?gT�wR*�z
صho[����?2Ja�Vk�Ŗ��wyGg�묽���du9(I�@q�j�xFu= }�~H����ch�.�,�l��3�&�r�K#,L;SJ�>��܈�����T���3׃�@�[�n���<�0��g0<��"6x\VW�г��"�ݕ��E���3�Ha��\X1< J�ˀ����ܚ���,��������ï���>�͍M������o�����|~�������N��7�Z���/�����Z�h[\<�b,^���B]�ڎ��I�N��i-�ܿ���4,̫��3Щ��s|����mz��=�g��:j�VC#�-����,�c��w���rF��qc6����	�Վ7��u� ̄Ǆ����
������\e�bH�O3�Ϊ���
�0=��ubK,���x�I���e�w[--�E�wM���!��Ϧ����)s�9�{0��q.!@pvv�۾,-�h��1)�,� �8>9�gϞŵ�H��
կ�����L�x��x�C: ���$jA����3 ��f�3����uN+��ZA���k�fZ��v�1��g�|`m��ߪ�ע��<�e�k4R�2��_ʂ˿(X�B�f�gV���2Я� zm�Y{��g�H�{�;����W���z)����ڕ�l�����,Lo�F��1�މ�6�̧�HZ�	�~*X8o@c/p���eI',�b�`T��:k�L)�)�����$K�6�3�U�56��Ka�(�B�7�̙��^�@pʣA�.ں 4� %�Z�I��ck�]�P�v���h�y��]�3�j){�
�E�W�P��^��0��}J{�O���D�Ff�^�L\?���2��6�4agm֮�R��؜�#���>���}-�Y��w��4]��zʣ���۳�!�wX~����6�I����M��2q;{r|r��2���ƺ����ų.��^��"d. q���C���T������K�)��DA6�Y���(�UlS� ��ڊ
y��9���_|&��o�&��ߕ����<{�T~��17g�4��+_}�����o��K��'�&��Q`��zЙr�۟nO,TNc��R�_ɡI�n���7_� ��=<W�|��*�=<[���hz��E�d��r;��,���y��. ~ܣn���*夺'4<--EA=�#˳\.�^΂�t��1�O [`�D���ޮ܏�Q������(�'F� �jR&��%;N���,�r~v&����<�}�n��\�e��.iB_��*A���Ѿ�H!��DX�g������B~��G-�qNж)+�����J����*�9Qpy{g��{���΍��y�`{{Gvvv�K�zY��\7�F9�Z��-�"���,8P�Z�.i1G}e�3�[-�"�5q� 2_b��þ2�3���ܵ�eA��O�6#��m�k�^K�� �K��imA��h��k�I�L�s��{�o����v��S��4���$-ƍ��]�L�L�8]^��]Cze����g���z,�z*&�Uc��3��2���ؐ�ֳ�J���h)���<nӊ����S��B�Tغ�Q@2��+zHP�,�:G{��rg��cz�v+���t���wؼM�yĿ�#��
@���E_'�ٰSq<dꝝ�da��z��Ng8�����Ol�^����M�n6�g�ʖ��G�¾���
(�^�|q��M�zew/����oSQ߲�����M��̀e�P�Az����j�*837�[����-K˹����,��ӧϹ CE��e��m��`9n�%%�D�-6���#9;9���FN��euyQ��N�(�1�Cr��-Y^\Jy��C'����i� �>�/�~���������C������/�����޽�rwkK>��3�����_��B��N�m�˝{weye5�T�n���%7��G@�K���1�Q0c*x�0u�5�1��b2Wi&��ԝ�q�� i|(�qX��K�G񌮱�q4��#������l��ŋ��q\d���[S�)�R��`'�Y(�݊F�@���:<oI#ҋZ��&��LkY�?`����S��o�&;;Oe{7��[dqQ��fXB4�K�������g�dc���R1����s�����r�=�y�0�n(	8��<0���a������
�A����u�_�|&gg��W�p����gd6�?@���s�|��#Д��-��pT��~tx��*�L��4����l���0��r>??���f*V� ���v���d�{�Єϴ)w��@'����R,�@8B�`�6'(�j2�K;G��0��r��}SZ��Z���W��K��gm�fm�>�j�)�`��5Urf��Ȁm��!l*ы��U�0ط�����݅/��*}�_j�ei�-��L��d�UǑD ��o�fF-|T<O�___#	�o�$��޽���_���Z�H���w&���`�' �NطȢ��7�����*�Y��Y����"�ف$�aI����2��~�}���N�s�kg��7��������1���=�Ct);��V��z�-���H�D�׌|��{�A!� �P���T����x���h���z��3:�צ ��lF-�V-�ea	��(�5��������W_}����0�tes��򗿒�׿�WG?~LP���6%�6V�=�wO��Rr���a��o�( X�Դ}
�cSFQ���މ������ݷ����|%�}�8n�K��zO666��/���ӟ�$Ϟ?����`���4�N� *��5�:�����ag��&��jV�O-���E<H,G�3�CFλ�p�"}=�:m�ј�EIDؗN�>4|)��GE� ^;�����<��2O�f�U��
��f%����B�_��,l��|��my��G9<ړ�O�<�ű�bL�`�9�LʰL9�x
�/������ĕf0ff�ȅ,�ӧ�h ���1��ċ�l�%inC1b[i灵Aُh��ۧ�,��:��Y|��a���4^��U��/ƚ6	f���
��*A�� ^$'�$+�9�\N_NO�bwn�x��X_P����(໸�u`�c�����{-&9���ׅ����3+�7��a��yq��3���Sh�&�k���K���޾Pc��,�'��
Ȧ������k�+��꿯�M>���4�Kޟ����huc/ԾS3�e�fm�>�V�[��Y�=֛ǩ��f��l��V�Ι����A�n�N�
<����U*"�U7�jZ�/�GT�oJX���mX؆�+ض���b���l`�h�q`���̼H�Iz��-�F�!�D�D3�p.�1�D��E�C�a�CON���`�Y�,�����0&99��ޒ�-����Ϟ0v08e�M/�
�Y����1�>'�6kh� �`q���?UaT�v��V��_O��/�\k#l��a	<���>`m����a� �\ӻe(��� 0��#��q$s���i���IK~�%��7����o�����?�@�Y����v[m b!~^7l 9�f�3v ��`ؼu�)�����!/^��ãCP�6�}�����'_��"n�G���A��'5�����Z<7;�3�ޟE���(��/A�}F�����!��n�Ζ<z��Lד�c������ɓ�j�)�f��J��V��1� P�a� ��v�i2H�bbk_�����ނ�Z���{{�������@`;v���Y�9��M�̍��_ǀ`70a\�P�1-cT��~�R�޻'��ߧ�L�1��ď;}��$��YJ7\[[e������+�z/�\���W#�' �x�XG�y���������#͎��7]�&��q�	��\��86��z��s�O/�Ȋ������_|����u��8_����=�>�L0��p�j�L�}��K�&���Z���
�[�E��}x�Ϣ�5������AL��3 n8��y�3nh�]���,e恼�m�i��Ĕ�.|iT��Y��Y�0[�N'�\yy;��7�t���0e
��/�7�tq�eD�Jhd����)@[d���U6.��v�Z��$!��R���HF0�1��7l��L�z�Ѕe�9� c�  �QS�J��˳~N��p|�n�W�e%��������ׅ���������`���vP���Mʯ���� ;�Y�ǧ<|���u��R�2�{h�,a��)ùb,�ڬ]�5�S�󏯛J9�+>��X�{,;��|�2�:��씋sb��:�藾k$s0n�y֕�Ŧ������'�gYܸ���%�c%�aі������������<��Ã2�0��,��}h>����ȡ]ՠ�M�bMF���777�φܺ}��"�� o ,Il����Ʀ4=����){�?O~|Fy���U���d�β4���Qr��E-��PQ ��Z�n��PY�vߴz�͗�`���͠�Ƣ����)_ݶ�a�.���@mi$?/H!���A2�Mk� ��8Ҵ,��-��
�'�5���gk�t���v�a�����&��n-I�#<?>�]����>�)^@�լ�+���/ʡ|�����?|�O@�+�b&�z�Eg/nne�tY���k6u�ü�����7�o�y]b ���hJp�,��0�\_����u���Ϊ�Ʋ8�<(P�F�;�&Jb2�s�u��ߖ�;whH���&C���1�F�������qy��:���`��������A�$�H����n�ֳG��(JN�-�\���1G�?8	 ��>���ӈ���nc}�2tA�w>����xmȥ�v]�����7����_e�\��Y7�6��� �uf�����
�c����Y��Y�����^dy+��7�|f�)Vx�`�Y�����w�F�(e̝��m�`�`;�Y�RԽp��D�G�`���uL�Ԃ��!�3>}�L�NO�S.��uˊ>��E�Q��3]{y�����o��b�!�ۢ���R�0��G��4 te���[l m�_F�n�C2�I���PuIb���fu�'������ЦFٗ�?���s��h�!����%��r9�^��me�fmj�ʝx_-���J�P�M��7b������i`���KIu Q#�e�S���	 3G�R� ��&�f�4� B!ռl���ۖ��y9X9���fܼ�����4�ʥ�5�`�P��׿��cK�풌>D�{�C��vK�[d>�F��j�ߕF(���k�r����X��揍���'�@q�򻾲"�|��������s���o���C�}q�Ln�[������"��Xh^��u���&����k �x���\Y����~��TTG���׾��n�}�H��/�k?5KK+�ˢ�f!0��4Ԕ��Ӫ�mM;�C@_Y�
H���2���q�9&�@WVW��q��ȍ��&�z��إ�L��O{Z�Љv9���@�vw��ؕ'O��(���z%�䥀�X�.�M��'�� _�/^4��ӧ,������'��C�m0�B��/^}ς����Z.@a�J�N��5��Z���re�t�2(|�+ �Q��c��@֋�=<�~�8�^M�����B������L�;�An2�����Az��+~<�O�/��q=(*v����$�4 �"@K�� #7󉙝��^�\��Z=�vǕ��������F!����w�U�H5|�|_]�Y��7�j�k8�ț�cn?|���P��j.��.��#	��K/x�> �,V��@�����L��8%I�
,��ra�r����0�:��[A���:��%�ڥ, >��gЁ��l?����G�ǲ�@��9�Y�y؜YS���x���/X��`�M ���}�� F�-l�N����X�<�g`��J����"�a�&�������"�+�>�pu���N{���,4][
..�/���m�fwS�I���ӹ\� �5�Xc_{�d�I�%�y�\��ڻ,_įt�R��]�B�kS��4�7s������� �/�4��]	2?wF�eaa(�~N��&8��`���?G����K���15����?�71ޒ۷���ʲ�á��/! �ej�,��,�����Jϟ?O`2�ʪ��M�Ľ���_��_�˯�(�C@oo�Lz���o�����f)�*�RV��׸]����I~%��
mK>��tr�n�7k �W������`�t����E����-��[�[k4~zz��ֺ,
?�)��ԯ�9D�[M��	�˫��6Q�	�U^��t�������|��c�߲ʽ{wT���ޥ�^�b$�1ZW�xOv��w�}'���,҇T��?�<��e���ﭔV\.: �ˁe/����~ݢc���uw����Pg��h�k�H���&_�����D �n�����!��`�sLEC�n<������2��k�dN]�E���"����>�%�)bĆ ��`,o�Gb5~w�@x��C@m-��k��åx��i�9�d}}����-�1�Y���,Yt�
]s^՟�kNy��b)���>0c*���h��'�y,ԝ�ZG�U�����k�^��:I$L=�u��rd���T������X�3`?ҍ@1@O������ 	�B�]��'=�ɜ����Ls7�o �J���	l��>�L�={A?q!�M�-�8�v'
Cf��%���n��V��6l2c������!�A%�����[z-�k���Ȭ�~-�v��.ˁ��$�t�_ �8'��$�K$H��y�c7'�����ECe��8�׭��Jڬ��`oG���} yh�����G8�g�f~�+/���L�d.��5���U�'������Y]Z>��l�n��Y`9Z6�/aJ�eJ���+i��d(�};�p��t�qÊC�(����� W�s?7ų���$)��|�Ց��ō������粶�)���eo� n�O��w����ᡜ��INd�^��{��s�C+�X�ε8�\�W������`��o��߿~�W�˗��|���H/n�s�mټ�&�ݖ�w6S�]n�C�ِ`�ŤZ\F���ݛ��Q֘ΚF4�v�	�pM�g�	UG����{59����+t$*Pa��`���*͹1N�8Q��Y1`/7K���{�p��5�����c�i���O�M\��H�M�nC���߫Z�k6�>��&�5���le�6emuS>�E�A�~�.����O�j�
Y	Z��r eq�A���97Y.�8މǆ۷�}�48�ܗO>���",0X��bM��y%�K�r����E��[�����:�1�=Ԝ���0ba����0}�
,�Ϲ�xKzNx�5��},J{d��C#ڍd�V��+���ZMd^��c-����֊�׊0J�`��%��ȵ "S4c��׻��[\G�B��WVh���[P�(x;�N�����Zb����u3}p62f퍴��9ȋH��i��$"���j�f�'f���c��U�>A�A� �I��*�U���q��%������'��\�g�lp�y��f���j�g�۾]T$?θ#�6UQV5D<���~m8n��	���
�̋�y2^U`h@׽M�g?�V��'�b��vcV�YwAj�H�W���@�ˆ�x7>74Дcz�^��x��1�'c�_�`ha��\Q�!ǲ��X^a>�.Ƹ����^� A����yE������o���$|�����P� 4�ςԦS���KA�
�����]�ڥ�[Т�g8�x�/�pC�k��9���e�ֆ���o �>��]�q����slm�� ��lQ�<���!�8��.	Wն��,~w�ލv��e6��l�Be�q"Ԑ��O�=���\- ZL^�G��߫>�n����wX��L��G��)��cHtp>APct�W��Q�W'�Y��H�A�`�\܈W���U������9:�d�9�{C~x ��3���g��nnޖo�FQ��qc�ƍ�H#T ���NJ��p߰����
)`� �q~�-'g
4�ͫ��i<ߟ����7��M~|������eis^�~zK�>�-++�rtt,�NO�8<˟��_��cNs �۟� ;����%�u�'��a�,\�_H/�����5��V��w�n�Q�j�6��XE>�o,�K/�Aj�?]wJ�	Ҵ����=�|Y��Ѫ"ɒ<C���` ����G#���I��n+-�47F+2�<�vk^���?��ζ|��K-����jT+[[�8%U'��Il���r��<~���
���?��0
��MSP�.�jG�ũ�eI@Y���ѱ~�CD&����s��
�c��vYg�󚭨
����%�\֊aU�m,��\�����������]j�L�v[�)���k@gCN���
Y������R�R�fd��2��Y�[m���'��������v��:)k��u�L쏺�ZJ~�|�e�G�p+��=�6����EmN)���dF�ڟ���^C��?�cX�WF�O�<L&g��u	*쪙��pa��s:pU&@���$g�]���e������}!V���v]��Uf��*�>��U��"?*�[&˺]-2Ů
omѼ�#���7�%�(@�6T��k ���8ee�0+��:��X�h ����e�,f��m��#nn.��� +�q����O ,����,2&�
���̰D�s#( G1j��gH���S�㼲�3f�Y�hq��s�Z�H��a��d�� l}Hx@�mc}�����>;�K����vh|]��$a@��sޓnO5�A���p�+�ں(�M}��~Kk��)���(Y+K�J0��aY��[��D��ô'�nm�Hd̴�[���?{���H�dF$�f�j�ގ�ي����o����<�ys��[�UE��5A c�w��� AMV!�Y�Dfdd��Ǐצ�	�<)yy�����eAw�����fH[2������m�a!/6X�,~S�b,��N�/h�w;=׻l;8q��T����/��_��C���W��?���˿��[Y�Ȇ����~��7�����H@Q� � �$aX����!��ᕅ�)d26�6(px����d(Т{�����G& D�����mK�&g�=�t�⇿wSn��!L�O&�����Ќ��}r��c���
���.9  r�麾��~�����ϧO�ܗ��ݻ��\�x�A	�0!B9�G�C~qq�2�dAon"�j��o޾%[	�k�������Խ���G���̣�{ñ!8�͞�MG�飕�M��yү���$��4��&{���
��n�R���/a@8�M$�F�-%�*��H���&3�=
�F�@�3�g��S!��Z���6�C�ˆ�@�T���+��Ts�+��FC�]�/�$ǝ��Q oe :���lO^���U��Q��D���^���C����0�[�������
L'{�2��dA�
�=����s�3��-�sbq�SZ
�]0)�Kl�����e�c���s����s�3��B�>��d1d�*D�8~���c_	�Fb0��7�Wh#�$A� ��ŐӨ�:��@���c�$J�Wɯu����i�ߠ��9��}0��:/�T�cv��c�쓑�Ċׯ�����%�ݜa۴5�_������3Ή:[)
���=3y8e���4�}#LV�Iy�b�P���"�3*,�K�rШ�l�UM�*���v�h:O�%��su��[Y���&eR���>_����?���?����V<dǹ�1�GY#�W삡ׯy��	xd�_�=3�WV�����%r/.Z�ÍFxY����; ��N�Ņ���?�ӟ	��Lϻ��5���ᶩa�����T;]��5�D��N�F�e�����o����������8�t��0OF�o�/?�����}ύD��K�8r�æ��~�:��Ϟk��a��Y�f	���2�_����C�?nk����P�^�����#�����`TC�=>ş�3�������ٹ��8�~�J����6�$0���m��~�ƺ�&`�ui�� ��h�F#L"a\,�1�� ���r-���2
T��;C�##��h�ӿ��M������2vr^B�o��}�Qm�H������+���L�u��c%Y���h_x��B���D{����8�tzz L�^I`N�*��$�:!� 4�E{�8��=��d2!k{��]��#I�|�l!�R����v�pχ�0$%� �4d�6v1�����s��{K���eɺ|��(9^?~��@4\��`#S�IYƸ�$R��k⿮��+�8\I�����BB��+���f^\���<��������
��Э�-���ZX�m��`�iy6� �����m�x���q����B�,���^�n�@R����̰zv%�F�c	�1	b� _憹�
X�8C�|s���Os\������,r����
�n4��v4 lsa�B���$��b\�L�MzMeq.�o�e��,�,G�S�&dnBb:����+� ���$5�d�a�I��{(U��	�$�Tf�������dQB�(�K��t�F���˰]aN���Ĥ�?|I�Y?aؚ=s#�����ӓ�W��3�+�����i #Y��H6�3���4j=!H5����P{�`�Lqy�b�w��F�vq�}��Y�Zǡ�u��I4$.�e!�m&u�t;��Ʀ�������݋�����}�������?�����u��?��������ȅ����\�H���e����<�w;�;nskC�����B�������?���uo߭��9LP�_�d�q�>�PMbW��~���X~��άը���96�����:�2_ F��~���z��X��Isӳ4����իW���/���'���n�UՔL��F00�� ����c�}�F��H����+�-j�e���ߩ�Ck�����~P�.}FA����?T��<R�z<Lzܤ<f!#P#���m�ڐ�GGbd�5sey�`/��vS��ι����	_��˴�q���*�b&V�"8mw�wܗ/_��* ��q�^][��߶��O�r�޾�:����lj ~܅�x7��c���YQ�:ˈ¦��j0�����|"��z@��������;����%&���?��.A��XD3���6���=�f&
#/;ncs�����e�g~���������\ �>=�N���2��0˳˅ڻfsb��>���~�1Ɯ< gE��NSTZ� P�x���	h����1��萂cewg7��-��_��2t�1�Ñ����� l~'�g e Y���@{�ㇺ�
N�I���F{O��6�^u���Y(8����h@�XB�)���������0O����j��xMg[O�f�K� �ۮ��^0�{
Շg�����U"�qu��݅�'���{�<А9���%��3zI�ۘ\���T���^u��@ɤ34��	Fv���^��7"^��=��0�}�`���I;@|�?���Ɂ�;_���X���%?L�N?z@\�2�����v�I��T�jM��
�0�cs����������&h}c i�����Dc�^�1�.�X�徼�ѽ� c�%�9>9����stHM,�72�Ԫ�nOSc��v?~tsS�$�%�MC��T/�6�T �0�\b[�[��U�;�39ܤ<R1Fzz�!$�_`B�������ïp�k������,���t4��d����:�d��5Qd��zi ��p��.u�5#2T��I��I���%m���D�T��p@�a��P������ <X���m�m|�Jְ9`3���	ɪ ����� k X� ~�}�H؀����۷-���\X�!!@j`��h�:�q��)�� �s�Q��ھ���Z�r_en#�����b ��.*� 
�1�ڑS65��۝��m�m���^�9�A�Ke2_��r��#bj���1A=�U �ag�~:�������&�����DiR�p�R�#�5Jר��)��BHS[xc�X��o
���E��xb&Z���)�Y�u�I\L�'{�=��,���+�Y�H��1%Ur�n#�_�����p�{8��dyj�7��He�4?�����q�߸�iI�n�Q�>|�X#18�u.y��T��y����蓉K����ycY e�y#�҈nf��?��O��4�8)?t�8���K��[�<�%����n���� a
����\-��E+��x*��Ъ͖!T�|�W^,���'ԧ�X���q��tH�J��i�vtݐL�PoNSFg�φ[^]#�zj��k���y�W�Q!�q4z�w�Ʒ�ܗ�Kdr`��h6-QI�!ͰBd�==qg�g��<nB�LiL ����R4����}���[Z�gP���}��b6n�ؼ������}�&�~�*�����������R=�37䘇ڈ<�Nߢ�Kո���� �d��b0�`�"��e��l����5���, ���(� ����!�EJ��pǾ�%���\֙X�?��g�������wD�λ�d|~T�¤L��+�����k7���J�}[��g��x�	� t�7@	E�`I��;k�ׯN�ke[4IaC��	����;�8 � �d}f/ؖ`��D�'�:�$�R<�2A0�PN�z�+���|DC��,�-�Ė�4D�����S����3��wd;�X_^T��1ۡE�j�,�S�Φ�5�b���%�?��h߽}~�3΅��Mx�����;.�_u��	���F1����4�eJ�D�{�v�T}�X0&�(�}>�S2�yq�1o��+�-�]1��d$OM%�q#]XRqq�H�q�Uvi+��5A�{)�<@Y0�/;d%�bc9�< w��'�)�L�рr2�Lg�O�����!�k���A0/ټ 	ӳF�.�Ѹg|���܅9�ǒ	�]�o��F�l�����/k���RLG���VO���t�Hs6�T��A��䄊�9D��)yx*�Z�K+Im}����卤%�0Q��}���X���V�7xD�M������(V޲�R��MA�v�?r�v<�ρA}���E73� �um�n�}䎏:�8�A��..�ٍ�0N0��N������t�F;e��(��KIY��I�_⭚jϺ�E��ݺ���{��f�-.Ϻn8s��;�c���
�9a����D��]1�(k�W�dײ�CC�y=����� Z�~�.O[,�"��M}i �z����5�O@�W2s�YY^��p6�d �q[�F�F�&�W�c;)L2�%RQ��<�w{ Y�������/��� �0y�/��PJ�ZT��t�P�;ܳ����^:��'�!
��r��R�k$(޼y�5�$,��-֨#�I��ɮ����_�H
&1~��&��#�.��X��� zð7�|�JP ����]XXd��]��̵[�s���E1P	�>�ȹ��B���� ��{F�m��o�a H� �$�=p ���X�g�������d����;��&Є��x�ta=ٞ��=�Yv�$��Lp\ ]��S#M�e��}��'{uڵ[�
L�I�}	�ss����:��C�,��=�M
�4�������2��I��Ե�^���KK�=V ��3wxt�f�g����2!G'R���9763��U8� �b,�-컞��"x����l�e읜�Ƀzz�|�`��D�@4��w���D��(c�`�6^��<�+���;�ڞ� �c[���<�n��!��9 ��1�b	�*`��\��(���[J���e�b��t�fR��G��),($g'�b�J�=t��;��ܦEOTQ��P�g��!��n���2ˋ�����V�8o@�������@�:��~�S�{2u��j �׵ӉY\�V���/n>�;[�nss�mmnŅ0~~q){<��N"�ڔ�����Kx�����F�2�UX�nN���Wnqe�!W�����2�jx�mQ��������pH��G�D[=Ǹ��#?�M,��)gD�����@�Y��jd�M�����~6�y�FՉm�18�������ڛ7`Dy?r|o��ZT��Q�UĽ����fsݤLʤL�Sc6�a @-��޿{G0�) -l��n�}8c�&��矹���@S�V�h��@���p	����&�Fb;$���@`ؤ]D�f��0��	#2�� q��5�"�] ៿|���/|��*�`G�9g�\RC��p���5�?#����[B1�ϐ�X\(�������fƪ8�6��㚦M�"��H̭I�1�F�?�o)��(��@_��)e	aL�������%��ƥ��$6�`!۰,�4"4W9��VN	;��^ _!�D�&�\H&v5�o�	�ZtJ}���	`��ʲ[]]�c��h$[:/�g:�v��������È�dfv��B[1:B��1_A������hͮJ�@Gy��:%4y �s	�(�e2��
�y�$��E�� �"�����LF�f��md��	��pe86�F6Y��WS�'�oR&e���/_�28��R|	�b,��F��o�Vm��8o:ה�	�j1{���I��"6����j��Ve�KM��%���g�(`�&A�6������P��p������^���� �<�
|�j�������+����=xv�hd����d�������	�|��I�Y% hO7hHX"���+n��߅�Y7�0�Y����>Ow`�<�y��t��xH{0�)c�L�yz7L7��ӳ��㫥�u��{8�1jq�+H��Eϩ3���j�L�pQ-`,Y8�S�\N#�B��#�Ӡt����i�����}��o;h�e�I�<�/�X��q& �^��<���4��M ?`�X�pFd��`�[)a� ���I���EkX�i�/��ĹD�]vhg�%McHj�\������u�N[�= 0���sI0��n�`Cx�z-��f	.Y�yE:��� ��:F2_���kO�km�u]��]��H�rpxH�����W�Y���\��N�{���$��i���g�fi���Gbs����(����B����aiL��.���S�"3IR�v|}��h��BI�r.`�oN��
Q�5x�q� ~1�,j���t�`k�=��8I��q���ʹ�*�!:���g��f��1>�E�Z��66����	�8$0
�;n6[�KC���|^���i���D�HBj�J�; Ь��7���}f8�a��p�i�����J�W��K��k�~'	�3���p8����s��*[���ѱ�#��M�/�x\~2�'���F�}C��B"�CH�/A )�|�2?�*��U2�iҾ�q�Hu� ��I�����\������Ƽ�jO���܏S^(����7)���C�"H���,�3ث��g��
��2�e O9�V@hR�a៞[�F�[X^r�>�s_ܷ�ono���5����q�.����x�{�K���C��^�h���8�º��@����[Z]�kxr}�࠿�<�F�f���>����uդ���B-�q�׵ޣْ��&��S�]N�~��G-���"�\��.����]ϕقbav�'w�2)�^+��ʓ�l׫I�!
l) " oVVW%D S�5��W����E�ܻ�o	ΐI|)Z�`.��@���M
���@h�V��of�LB�԰A�_Z��s��Do��B ��l��!�U��M��՟�]���M`	R���������N�v��F�� $�j6���@2�w&�"�~�cp�� �����>�5@�`a01	�O'f�3٧�	M̔�T�e��1vဈ}��G��MH�� ��M��� g�����5�U�7 [�n.2y
��e � xU;�{�W�^s�8��^��8cNh��I�Ѩ q�t(��s]2��x]8q�d�V�W}�'�l��+�����Q���G*V&@z Ј�,� ����u��j�{�}v�?"(5빲���=88��Ü[][s?�I#(�������"q)�0��#���ٕ?ĉQ0)X�O_v/��`\�9#dF��(9��������Q�pxX��I[8�����M��S��6�_V�r.��_ƒx�x��[a2�^H���囖06�l��X	)�|9�ǆ�lݮ��X�p�w�߸�&49�?wG��Q=?�CXX�./��Jd��$�Mt��(�I2;MC���L�n0J1h���\ή��Ѿ�G5��ot���#���%�z�b޼�����(���u廳I�Oʳ*��ÏZ�5��A�P�7���4hS�gv���{�uf;i��%!�ү �X)UW�G[π\$�E�۬&�5 � �&3����N�f�9�����ʵ�Ux=C���� `�-j ��_�f�U�����^A�z� kx��6и/j1#4�V���d�i(s�	�b�!������T��]�& �m��ƽ�^da�U��z��Vj� �Y�ϫwO�C�
����H3��)le�4|��bN����FHO���WO ����L�T��S� #f�������2_���>���0?7���xp-�1�j�(��k]�VǏ%'D�yLz��2���\���%�X���
7,W
�nb;�80�S]h�U͆@������CBz4C<oa`��U	N&�$��:�����a�(�MnsΥ�b��0���8H��9&��I���d��[j�Ic�>�~W(��������{N�@kْP�Ę�\yy��j����2ʲP6s��Qf�h{���ﯼi���.�U(u4�27��7�/<��u,���~�pL�^0 �/4�9aD@�)S8N�K-�H�r��''��4�`�E���ˤ�M�e��<� !��c%�����xM ˁ�R��<H!�������;����L�vx��m�c�>F]���'�;Ï2SR�r���]��m	��Gә� �s�w�0�\�Jk}R=<C��;���d���;7��y��I2��q���_~��n�H
c3�G-�u'�5�e��w��*,3����>c�\����՟�h����E¼�Ĝ�<@\��Kv���7���������<����N5�����*[�*�@%\����� �+�̒Glna��ih�b^Lk�C=K�� ���6����\H|`���y��
.m�ѿ��lO	;��b	�o�d[��_Z�_ˇB�*��`k�����фb�d�S���8H7ٳ=�Ap��(��I_���\ù0�2�UQd!����t�	'���d1^�_�
��qnQ~^���Ke�T�ש�$%������լ�����������D֤���BVfj�'���87�� ���NԎ��A�Ζ$�G�Ƣ���M�����$F<���D��Y {������cp]2�c�O�S�#��5n�o�2W�}���a�?�X��W���KR5|�O&R�q�����Xou��GzE�q~�H����"�\q0��Wa�N������1x�k�7I�ی���<� c3,���cǶ%n D_[�s�g�E�;`ٻ��O�*u�囿j��/�gU��}��P#��^А%.��n�5�������ǩ�������	��$���ԁ�"r��l�W$Z|���<�Ĳ�����-m"b�<�bhi�g�Ωy7��c��;ĔS8�}���*/�6�ܬQ��CAkӦJ��n�b_����*��<����F�H�nr?v��0�QW��*7�~l3Zt����&_>�\5���к�왏�����w0<J�=�ǚ8����C�P%��C����esU�XN/,IӰj����~�	�#.o���� _���y�����!#��
\�^½{=O�@�Mڇu����[[]%�b�v�i�0|{[���#�B6F�^�ʖ
�>��c)��V[dڔ	f0��s��==}N�vwo�N���9���),�x����mk�����w��!��*A3$�Bx����~O��=�NNNɲ���p��6@�&���C����2��$,�gn~��SO�}E����.�IS�ɼ����'��c�jl�\1p~������i�O�VlG��wJjVZ���ƴ���x�5ڷ�D�;gB�p�v���\L����矘t�1��\�C�7�z}�-c\4��/�	8���K^�9��2��k �����y��Xwt�h2n�D, ��c�w�OD�N.�p� PF�y����t�nl��T��ֆ&� �+S���~�6���~�h���J��z��=�v4钐�9���8��ф�♙9�)ss��-�Et��'�<8z&Kn`R^T1�V�g8z���!�*C��c��Ad�W��KbI�D�i6S�#/���Չ��ie�I�Kc?_�z	-��]W�����h��T{�7p�.7��}�3�/��95\�d�zZ`9���~+1��/2�\��W-&���p%J�����i��6�����4�:W~��N����.�&wQ4�k����nh�|u� �TrO�'��ma�d��T�\K��Y̓�@j�ۊ�������>��?�j��J̒�7���N8��[GY��66u黖Q�q��r�2�9Юf�o�i~uI�8�f(� ���g0mV�(i*���h��<j����B��9���Z�x=Gk�����K�>�\.<��\��!7�}��μ����;^�w�l��K�%TQ@���U��n���X(��Ⱥ��nt ��]+����6qD���S}J�pӡv]ƞ �㭭o��ݎ[[[w��K|�	ॣ���m�h�������e����>
 �5 ���
 �m���%%2fg�HF}���5�:Ȅ�fg����7Ɩ`��d��)A��]��S��bn�c�r������e���vS��0�}��H���)�Ɉ���\bX�<��fb����N<�2��K� 4?�������<������Ϥ<|��02�H�p7l��qi�tDVB����ʶ����ꌢ?B3������k��?�c�4���G�oL�<�k��pDd-�k��N��z�0�݀�����7
ؖF�j��4�W�sN8�Db�,i�}?C}!Ãq��,�Ϩ��yO�nmu�����b��s�}� �A���lQ0����8G\��� �;����&嗁fQ�2C�פ|'%Q��8:��[1�5�G��i6j:뽞|kd�����IcU���ڰ5�@�s�a)W��qnJ��������2�vs7a1.�m�٢�g4g-?�5�d��u'�*�������_{e�S埧����:���@�s>�0|�� ��Gؽ�`1=�:�Y�Bt��ؐI!.'�A�h(��,�&�~]���Pݗnr�
�������d�p���l�N��u�r��_��Ö;��JH��1Jcc�c�}���mow�}��.��뇜{����VΑR����@s��&�6u�sɆ�8������y�-�7+ۢ\���:��'R�<��^J6eƞ�4�7�Nv�/�� �쩆��w�S�Jo���j���"̿Ҍ�Va�&PC?%:	�1oL��>]6�]�>��+6�c��8�KZ����L�O���V�Q~��V�!�>C�y�1��ՐozD�L�;;�cZZ\Z���A�HQ�X��vvw(��s�i����e��d_^�vo�5���#LB�g�fඥ�hh�"�����XH��qFpi$	-e�,�$���6��p�v$����'Ǽ���M�g`L�<�]���8c�����P\/�!*Iu��F0�ak�ǀ� �f����m�{��G�ծ��~H��G*!��o4)7,֮���	�"�#������!{:�3om�ՉO�l�2H2I'�t�+��ј�?��~��J7��� �T�U˵�`�����0t��D�`a��V�DI�$H��)�E��P ,��7��y��3�h�S[�Y�p^H^�v�s&K�gk���I���e��|(�MU���H���dT��C��J�xř����+O��5�Hײ��~��Űq����Z�"�6�ϑuUy:�r�-�����#�`[�}Z$ ���H w� ���T�8dB�j���� �J�ƨ��}�8�����@y�LF��,���"h9c٦��^��']����V��!��Ň�y}G1����t�7P�1:��n�lI(&��Յ}��K	I������uG���r�+ɨ�L��N�t�A�u�I?>ܢ}2;��� ����<PSgg5�����iC�%��=�%��C�0���j�jV��}��:i?ֆ�ޑ�2��m���}�0�w�?���'3��D��;�s� �o0�+'h�N����[�l}��<]�Xe�d7�$_U�$4��S�3����qQv_�4SW�>��Y63lX;f#�!cD�#(3�]��9O]l��͜[#)\g���~���͝��ʢ9�[��h~����ng{�� �!�33)��@�ϟ?��_�2�������Wdߡ�=w �TU����`#S� �v;nN�y�~�R�c��H|��4?'?F (�1-�1��Ź;>:0<n���v+���N��[�[���%#Z�]��^��o�\�:��w����XW D�G��g):�8`���,�5ʚ��H�6@f�G}es8��m<1��&�W~����LJǒfe�R�4�Ջ��8U��#o�Js2��tb}���:c�1�I����96�ˀ']7��m�{�ip��~���==������I���+a���qF�ĵk8��$P�< ��P��d3�d��`���|hg6rv�Q���W�k�I����u�e�Wk�:B:�X� ��+-sdǎ��C��ֶ����+|��y�k�������8�{^4�r6q����
*��[�.���w���W��}7Q��bz���*AL���_~������@�&Q��x�h�Z����{֢?v�Lٕ�����i�I��"5�M�/��נ}��V���M~�V��������T��ؓ��^�.�*d#��_��5E碇4SC��u��F�'L�9W���� �ւ�e��O��ԀGy��W��}v��`}1%��u1?���R���'V� �e:���Զg�K@0�vF��pS����`�`@n���E9gתֵ��]����=�q�w���a��O;�1J���{C]�f�I㋑se>_���<�&D.��t�k�G�d���א�w|mI��ns+|��=P�=�u�/@O��X^Zf�vS5\���ݡ*ؼxiq�a�	'#���&�C8-�0�K�a��x�����F���� f�; �-q�2 lk�c�	�K�lc���|�$�]�4f �AokB)��`&�^ ��1}N`uX[[K		ٟ��i���Q�3 ɨ�	V2�e�am����bs]���H%$g�6�a~�½�8��Z�<�E&�p����v���jYD�=�t�l~�8��u���Ҩ*� �Ym㞬����6r��<ʠ�v/�4��h4z	�a�['�H\�^��+$3r��\*�;�wW�f㌐q	��_\�v{������g_Y��8���,����������4JF/��@Oz�ɜ*�Cչ�z�7�u=��S�;��la���Z��5ϭ?�q2_z�n;o}^Cϔ歊�ZYW���W�w��+���?zIٯ�d��d�QW�^X����ō���UR+��� ���;m`�]o��]-n"HH�ArL3�ި�o$�T����P?�� �����0v��������ō��'�ŖTN@]��
��e0��j^�mac�$�3�%Q�m��t4#�V�j&bf�<�E�$/�uǊ>c��)!��.�LU/-c&W�S�Y~_��7��j�d4o��%U�!�k�+��G۴	��_��V�>���:P���l���#�vU� �H��o �y��������0}k�G���=������l������4�?�A�IW�x�ʐy�����!پHF�S �F2 �
�/�_�~u߶��{@yeuխ���kh�Մ�9>>��87
���Ņ���d ��f�=�&#	��1|��aR�x~h���LZ7�f�'�����H �1�󟟝s��>qO�� �mT���}�c灦�����-/-������O�Lj����PI n�U�ǣ� ���^5r�3@�j�nR��/�r,d��L�=�M�U�)5w�{�O���~�gka>�?0cR&��(��ſ��R�R(���y�1�qM�ɟ����J�6�������v�}Դ�W��Iy��i���Q|��d�#�٦L�
N����9�0S�2�0������N�0�PI[ةLw��q��Y!5V$��{�W� m��.l��*`�|���6��A��g�6�u�	�3���*|Ψ��{�x/%���19���O'$��C�YA�6'�m�̜� NJ���㸥��c4tfX�&���}.��(տ���X6���+���媱�����8\ݾ6���lH���:�@�aN�~�|���a��,iR^t�1�3P���	@�3�Yf�ڳ��{�*[�y*�0)�!>_�L7���N���~Jz�����6m�$���ِ�����t��䘬W&S	 f�./��s��a��p�7�^�s��s3d�"�@��22d��m���q����恱�nO���U�2/:� �A��$�9JO��GG�lc �����/��t�?'�8E����C�_C^� :����/>s�|ӊ�87;�dR��]��\�d���	���]�m��V&{�^0�{�dTC�& RGwo��!�8���Y-.-񺻱�_�y�)!��>���nZ˄�.m������<��a����7>�K8*
��,���@R<+�����vD���:n��p�������~Ўq����ÃCj |��)�F������R�u��ۧ,�F�B�������s�u/{�[��x��++�,ų��m�v]Xd�1�ڳ�l�i�+�8kx���5"�m�ǫׯ��� Q�捍~6;��>�G'�c�w'�+�R�ᚐɀF3���A{���>�\��s��<�VVW�\��Fi�[��Ka�b,c������X�;�]F�17�SL���l>�s	��z韚���K	����߲L�ҤL��Sl~º	�0J�8�>��KD
�v�L6(�3��<\yiP��Ja�k� ��5vjđ���!}�lM�4�u�8���g ,��<��U�<��Y�s2?��XTu��l�\n���]G�>o_?��TpRu��l��R@No��A�P#���?�[��%��G�ke4y�0���X��mQ'���0��[��a�ԇoV�2��yH�.���rS�uVTyg��2�_io�+��;��k܎����0��f���(�eC+��� �_��ɯ�(_p�Ā��K?�L���K�@!ؘ���d��թ�a��#B������;�� @ʢ�����$�C���o޸w��0Dh��с���38�t�j�D4� ��u���~���%�D UGG�LB&)��n��%�����cq���p��p� ��>��C9O�`z���S�c �� l�]޼~�i��m-������%�F0��g���]���D��u�p踾��v��|��k ������`̂�bs(΅6�\���%�6�@$��}w���pCI@�0�������6��?��J?���~h;�9@��'��E����?�0���`�˗��?sV�gw����0Vl!�3�kt�{z:� n�J~�ZQ���: ����O�웍�; \8%Pg�}?x ��?�y ��k� ��S#��iJ�4j���؟�x}�����K�y<?j9�/������0%�`>ꇛ���eB0 ��g���J��}g(C9�E�]JSĿ�7~��{J����G?A[��6�L��vuu��Q��k�$ZC��q�>�{G�DB@�+����Y�ϒ�wJb\JΣ�ٙ)����e"�q/%�7^Wj6��nRmF#��X����:佔�㔽��>B�p�'届��ޖO>1��IaR�e�O��HU�r����*s9�'E��9�ݤܴ(�2l���h�Gtl?���B<�����$)�v(q�֧���Y��(s����>�bxx��
}2!^�YLX|�i������[�E@���a<#K6�N���ϙQ�h�DE����_�ߘ���*� ��e�	��mC���i(+F�ͱ����+׳@�T��N�6��ݓ<E��/9$�pb,L�]K?��!� ���&�:�|����W t�s�nmu����G7=5C� �?>}RٚlL���' �͛7q�j�e�������od��l����,���p�
F&�䗯_�eGؒkk���� 7^st���>;;'��
�@����+�O �sdUR[�+2HN�qG֥/���	6(�.0f	�D� �0De�B��0�X�pԴ��yp�/I�T{�6D��� H����M�����;;=����{ʀ��5f7�.@�#��:�=$e���!�`�ǽ�|���� P��m2��/_�(k�IPm�d� ���rˆin~�rp.�������e"cb��MV u�{!��vPg�����Ž��`H�m���&<� �¬?�8��t�D�ah��U��	c����ӳS7]�v1�?�թ��k�&��D'k9��d�{��;�"��Ȫ�um-�%��b\��/,.P�B����V͙, ��\�& ��ϤP����|]��f�d;7�I���ׅ�3����d��lS�m��{�yK'�^�O0f*�G�676	�c,�	�U;��`>w.��^)��󹯁!3d�yU�eg�������)u�n��8yJ��ٔ|Y��?Y�h�I�Iy���k0�d/1�:˗իdZa#b��u]��+-fM2<7/��Ї.�`=�}�×^�+~2�-�a9����P�Aj�~��1�RE9��d���
��^�'�S�d�~�5���ϓ���s���-P��g�%�9T�^�ZfO;�]û'5��Ძ�ib��pϠx}w��M�]�=�7|V�[���C��̾��)4�4��<�יc����]p�{�U��g[r�1P��
 ���	��� z 6Dh�l~a�`��`���
�*X��߶	:�<`�tB1p�`��)u���H\2��%A-���� �R�½0S�� h�kMO!�����~t'��\+{d7����Dj`��� ]��A&�C �*���(la�,�#��`��L�J�x
H �ch�&7�9�|���H�c�3�욞J_���� x@�����ų�Xhr ��P8��s�r&x ��&�[���ضh_lrL��||^8?@s ����cR$8?���O��,�g<�3_�$&{�I;�%�hӂ��r���@F �"��L� ���[#P��,���>�i6nf�c��UI�Ef�%6�N�m�%�P�����גZq��5	�0�j8vm��Jy����d\��f�W\�իW|m��B�����\��-*�ģ��x/�����?���a~~�\�D����7niy��F_¸��o��l�_>��{�g8��x��۷�p���)J{�9�,������:l�>�g�@�d�Od1�.���kt�Q���/�����O�d���K��'�E��_�ȼ�BbII�R� �?D��1��Ǥ��NF�-�=/�9=>+`��7���wn>�����*�йz�{��C^����5�����y�"���YS��Ɂ��l��]\�d�QEkr>��Vw����'��)��*��י���Y�),�N���]5��$�פ��p+<��K�B��Z��>�=���v&��Ǘ{+s��Y�v�^g��#��7a������� ��x�;����eRnPBE��W�1�B�U�:c,��T�u�k|N9��O5K��0W�; ����H
����>�qzr�0x�/8C 70ؚ'����M�hAp^z�`M��S� ����\"_�����.��ׯߐu)��Xǽ� LK(�<C�x��5˃�4@���3wt|D\�`�d��.�`�:�* :���� ��6��I:�y�E��p����f�bc'�/̹���  ���;;��nhW�/ ^�� >�
���%�g����9�;v�3����ٳ&{�$o�d�Ŧ�1X��� �ZR7�5΋�&z�M���)s��D?B�Z;C';( �s�R�"%fw|F #Q'����X	�
�H��szr�v�6���%�:^D�	����B6�"�;��`���� �?�L; �%C]C����6]d?�yM��O
k� X��K��D�eiI@g�'��3�m<��ilDs ���K���G�G�襬����fӛF9�N�K�޿{�VWV��~�$� ����8�p_�k�ݞ8/x/K|�`��HG�Ei����Ԟ��2)n ��;������%�a?���`�]{���0;�\����6���	V�K��q�*�r�[ɦ����1ʳ�+���Kh"}=�.��s
҆�F�t[�xo`�w�@u6z�RvPbN�0`�'f�=���e��`�癳el�l�r�]d�j���%rOQRhF��|��:�]7/���i���d����]9����#��[]n@���p���5�Ǻ�P���a�/aȫI�H& t 	$���u��*�`	� d�2YZ� " R�?d�<�/��<�GL(��s2a)Y���9�4��'ե=w_>%�F4Ž.�B �`�]� s�4k/�skkn-��׏y]&�ݏ��фh]���L��"{=�����`(�����8���J2���u6�7l��D�V\>;W���v� S�����XF�rz�#�
,�4�.aG�N������=���z5��?<< ���^��1�9�!�-ع]mC�e>%�9�}����w����&2��@N ��|f�y �%@
ٔX_��E�)��`��yye���g		 ���g�I�|M ;~���6�3@�6UB�V7	��"���@Y�_\�35��uQGO����	��� ߛ^\���`�R�#���MOǱ��F�Ӣ6�\�� �c����D����t����f����t����sB�9%�{E��QjAe1�� �L'�Ӹ�'(<3'a�`��Մ�&7��T�9� ��[�E{*Ց���>L]M�'�;������B�u:[�}��&��M�s(Y��2��C�}��G��l�\Tx��{˺<�E����q*�U��1�3F��9�F�!�v�:wZݿ�E�~'clR�>^YBr�\�R�.���<`9�k֓$�`+nݎSƂ��ػ�����,��,��m1�L�Ebi�a�����Pߋ3n���F���f�7�Z��I��}�u�O� �>�:��ׁ�t{v����29�P}�݂�Grc��Ļ�$ԫX�!1]&2fc���3�iu�ӹk/�kY���9��%d��n��S�[��2����{��c�y�.��Ɂ���~��M���u�1�?�D�=fq.�f��x���w�zʳ	(�N�@o�����B��r��H�6�&c`� �{
cŹ 3sum�@(��D@�^Y���%�-�{� 7�4	 d��lV�� Π��#�#�hG��յI���y��yl��hD&��'��px ��עm�;?>V}�%�J��]c��,�D�tw��le��[�ڛ�P�7�����9zd�v����7�[�U��@�^�Z�4y�9���7�y��������
$V�72���QozV�?�➓��qg���;��+Z���PG�M�w��,�i��2Ǡϙ��ii�\���6��%�W�ӝs�����.��`������v�:Ǿa�zI�'���=�I��<����	l&��K2F���~k�3�^K�Yp��՞xȀ$�S��ֱ�����q��y���- 2-��-�lӈ�9@e3�u|N�g����@4)����������M�������g.�[��� #�X��(MFߑ�}t��#��'������\��<�c���g����PO݋����(��*�E���	3X�ꞝK�T�"|�g�� �w�^��ev����l�|�r2�j/��D��#@g��܆������sH���7�j~�15)�_2[yp�Q��4k���^� E�]E���LD�,_�d`����y	���i]��C70]��bI�~@�w�59742c�&C����ʹ	�>�g-�6�����'q�7�FD�eW�ԙ`��#]m�D6rpe �QT�oj_�����{�ck���_�9�g��qJ���a�>�T��|����X�7�B��8AnV*�5H�����]T�
�:�1����.`uy���=�~����F;�y����)�oW^R+� %�gf������P� ��o]2?!wAY��M�gL��,
J8�����iJȖ˶.
,�C  ��mO��%��s�/X� �mo�J� Ωx�T{Jէ'�FR0&lk�	����(�L2��Ϲy�(��f��2���{BH�Ԙ��\ ����	V��P�v���X�#�7p���<�$w!�pL�/�g��i�.�(�YK�g��{jӘ�{)��9��LPH�&����"��h���!ӱ���>����g ��v:�=\��~��H�h���]��M�>�������s��{ɤ� #L�
�x�����%0� xh����A=)}qr̾P�i@�Q�r///���5�D:lnYRt�Rٌ��z#�@@#�\�j����������s���fb�O�"�vM��ٓ��������;Z��o���Z��9:P�@���T�i�>�k������z�׷b��N�� NO햌͇.Iùk�@|��*YzgH��ܯ�]�8�D38F��v�N�H@T{�He�#�������t!�Ǖ	X.<u�GV�L�qYr�Y9m��]�F>�c�r4��Q�����T��00���;�>Ʒ��f����ET$�jL
�^n)�xꈮ rk?a^��FH2����e�-��3Nʤ�K�q���>��IF�	&fX�}/�\y��M����q�alc2���q�Iy����2���k� ���`���a`�md��D����VO���̠�n���l��n�P�A@�o\Q��ٱh���,,�1�p
�u�Y֝I����p�L��
v�Z���a�����Շ׶Kn4�R��e��s�"���?�%]����<�V�Tws�ƺi[� ��v���}�5�E�6l$1/��#��Bܮ�^�uI ����{��e��?�ga�Ǽ�skG�~��ta����H5�]�z@{gbJ�Y��H��R�����`@3��X�N/ ? `�B� ���<źyp������'�+
٩�+�+n}m�-..1�@���7�5 �������"uv*�<3���&e@�a��c����B �8'�!Q���#h�ĺ�>`'�5��۸8�3���� ���dn!^�`����k�E��<�z ��sJ̃ "�]Zʞ��ޥR��3�w	<�L����k����@�˙Qe�������s��]�,�o3^o�(ؾ ���4Yʍh�t��EC4s �h�g �<?SϹ8#
a�>�$~�t>;���
��m�}�
΅E$ыmV���1�eUb��}��^~��-�y��o߾%�M-�%ѳ2~��(؍0�� P���gqo�^��_�~�>���}C�km�O��x�'�?�m���n���ݵ��o�=g �{�b Wn�ݸ}�
ѱ��A����j-Ԓ�B�e��kQ+7����hL!����6��H�]mrhO3�̀U��	zYG�$�Ut��v]��D�`��w1�A:H ���-��1�^�W�cP��&�4��Q,�*�I�x}]� ܐ�˶�c}]�"�d�=�9����֫��O�{��=X'-�¹:븶py�-T6���6�c���o0
�˵B��tTMʤ<r������	��b:�����J���w�d�#�g,���^�u���d�:9x�sF<N��)\�o�e ��;���(����~�p�h��!����Q2-Hl�/�*)l�����=wV��K]r3�EU��f����L�ΐE�Ss�M�O�M�0��ٝ���䨋��ώ�9��zWN
�WN�rH;U�_7�j-<�7�R��r��̀�0�[nDݞGɓ	��D�f�j=j��\Mz�!�3aC�������h�%���n�mdF��-��Ureds�>���~˘���6>�zb5O��C6У��w뫾���嚾�h�İ^��d<�(c$u���M�0�O;�����F�i��+Z�`܊�m� �܀�R�}�� &`���� A��舟�b���E�1����&G�����g�	�.x��I <���V�R�%�)z� �>��2����aҸxo=�_h/\.P��8�#�--.�Y��������x���]^lܠ@l	���L�M|�C�m��I�M-��hc�m�=%,p$��!�jz��ݪ9�R�26X�"��x��� �q�X%> �3��A�#���U�ߥ�J�4��0��$��zX��:����@�]���gи.�.����ИU�p� @ �!}1�8��R-���}�<g�����C� 5��� �%������ͨ79F�ɷ�*��������	.[��D�J��#�%ߍ�<�c8}0�1j$��S�I�FU"=���9�08w�PO�L2ch󆭉D�K61Y�8o��.TR�7�45b���1y	� ���̔9�l-i4���w���.|���}��oQ�������t��.�p������Zl���%��E�P�䚖�^������eFh�gg�C�41���d�,��Td���7)�]��D�Hv�׹%�F҆��o?^�BW�����_���?��I�q��ϋ���k{[������U����`^S�l(��@F���g���;#���'7A�#�E=����T)�",ԗg�=#�go���k���]��Ja݈�����&�dN����{��r���r�����=������>��`��;�iFdio��%��`K���7(����a�����/F&r�YcLʝ�Gz�X
dj��;$6�9��4�eK�#Şa�@c� m�m�m��KQ,�!ߵ���<�7d�yi�_�A�V��6�V����V�'-7�/�x�f�Jb`�׸n�}<�r���=5��VW)S�� К��zN0���3��1`+����]�s`�nmm���}��<���3�s�1�� !Q��(���b�64��
2`��0��I {ee٭���%e@�!�����7!l�3
� [\�m�  ��w�ɞ�\��Cw�j��А� ���ꖺ~�NEw:��e��;��=�j�u�!�|���,v��F.--H��ؾ�#��.�s�L#qRW�֥﬏�+`��[|��1/�p���	l�>��{��о�� `�ԮQKvO��-�M���e
O���j�N�_��L�`M�5�pb���ϼw���9W�>l#yh� ï���?c�]i�`�7���NfU�a2�팣���i�a��6z��o�3��g���*��U��+y?6n�\:�G�N8:�|�ʦ��~��=�U�)�sp~��[�����k��{����
s�G ����h"RaC#y%��W⼁y������?߶�1�G��d����+�*�Җ ��q\�}ێ?[�;�إX��I*�*Zi-�Ze8��[\e��G�ߘ�&��[yG�(��Ȕ�Ņ�H���E��j/^{c\�9�������إ�:L�� �N����G[#!�oEO=�����<8W�<�@�&��Bm�Iy����4�0'��
�У�ڔ"�Tj4�l�rY�a��������S'�E���Z�3l�'������r�`��<���0����@]���ݴԌG��:O�Ǔ�Ӹ����cwȟCwv���=eY]�좪������o|��0t7����q_��[{��>|��l�0|�p���`�6��PcW���|�2�o������5�2-�aP�]ީy�j���Dc\
� �ϩa�V3��~��B�ɮ��ɕ LX�yS��4���I3L@��o4�� l�f�0�oV�����I�}���e��S��7�2���ÿ~�c�t��'s�6�����<�ߋ.��3 [��@@�1gK����������*'ύ���;MR&���̂�6�'0�7��Y'-�!�cS��`�&wo_dD���iB���j�cn~�����2�il�o�۬36�3���$lC.,���@�~68�7�U[u��	��� ��� Gq��Rp���Ҏ 	�r�jl���W�����2��8��M����sA��s!�1�Q� ;�F[7%����CK�2~ a�k��u�m�:��}?8��$�u{��� h13;�{�� ��n8 ��l s���
�̳����L��@{< =���d&�굌5�� ��=̡`�W5��L�!��!��^w�Z�ѐg��IL�!���}����u�ڱe����9&W_���s0o[�D^�m<dI.W�dҎ����F�@7��p:q2�<�������:�_~�ïn}m���R;��͍M���W����h	a����Z�>��޼~�9s�(�gk�AR�Ҩ/�8�PǕ�U�.��kq.kǹ�������܌��`�0�`���k���ݛ�o���F�F�|���~��7�d�*[Y�N���|t?�����kb�����￳^���o�#�N6���>����'I���<�(������q������^�kϼ�H6�3$��b;;���q�F�w�ע�71  ��IDAT�5�߿�@G'l�'eR���s]��\:-�l?9�PTr�A�$��*)����Nۺs�ݤ<|IZ�9�`Hۋ�����g��E�<�K#���_�W���d��*�W��_�=��d��̍�����<t�;\��O�]3*���Ԥ��Tkڵ�\��rؤ Q��g"�2n������^\ȱ!:=p��z��[��g�	7��h19�m�dn2]���|��l�����G�����B�����Q^uJv�+��_��S�Q<n/�] ��)�w��CP��&q���� 6���۩�' ex0��=�a�U�0|$� 
@ G l�TV�٫��Bس�]��}}l��m�WJ�'\���4�@_1O����������-{�a��A6�w��&�Ոb^w7��������E��jqͳtSS�����p���#�F�� o!nB��|&a���b�t���qʊKD�����ل3n�͉%I���.EV��Ț����W4�ϔ9��z�\�1WaΓ�D�$�P%o*k�DYSdz�
zhR#�m�p�h�q,�Rl�������tn�����D>�W��CC�\	�NNx�2��f(�奰�����<M=�6�
�3 �,g�AJ�%�:��2$ֺ%2y��j?7	���fI�h i�4T��B��;�<c2=cǣ>\[��D����h  ֟��ϖ�K7�y	��`H�n+��}@���������H�~��Q�,e[�ls�A�@�F�����O�f(�?����\5��{o�sښ�tåj��<L�3�m騈Ǧdy�c=\4Z5ao�L��ڏ�����ɢJP�DV�`H��u;�J׋���́R�hl���$o���"K��ux#X<�2�Ÿ���2B���b,������e��&�Zf��g_1\{*�u & S�k��̍X'pسG������<1_��Cǹ!�:"b):��a~��9�$���Lh�}��xs���C��nks��I�E�p�W�̋��{�� }�C�'Do���8����A�vx�N\�uZ��f����{�Ǎ����6x���50/���%����rY�}m�ŚJy]���yђ��T�l\��-e\��ãC��߶�&�4)�2�<���k���`\��&���D����˵,�e2l}���|��^w�7Ga&�&%��>a��6��t�#o�x���ҫ��eS��ҍ���Ap.�\��J�������C���#w�sL�,t�����E@y�57I�P���������7�o�Ƃ����>�㺳��Sn iD\�x�������z��������Odg5�4
����04D��R7)��O��B.����$��Z:��̧�� 5d>����<�nC�G���4���,�ذc� j�c��ϟ��/����h$��F*؊��6�`x�[/m�c̱�����_�=�M>C��)9��FS���%�=�������{��؇_���:]�� ���������_��i<�����nR^b��%���g�+t/l���5
�w�߹�o�r��K\�~;M�<�:/�~l���MX�sq�|�kKdzF�Jn�yθ�n������d#�\Xk������>���7�y=���,�(aHAB,X�)�8��-.��#�������d���� � �������e2�qs���ψV��w�I�� �v�R�	��!�_�-���4���{�6"-yS���j"A��S�3��_~������@\|��zF�!\;�_RȳH�����]v��`�ӑ��f�Qa��LM�>��p�\{�����==3�NN�i��e�/l���%�ay��d�6B��xÜ��v�%�H :g����C�<�`P�?��=[2G��"�U�� �ds�c��-�{.E�N���_�߀���Ka
Rv��&�`��ڷM�Ԣ|�n���d^-����Z� �G��R5��Q���@��Sѧm�=s��aQ�@W��-�1Mb�GS��iU7��5?�
�Fx�hH�YT"X�SS�:� �T���H�������&�%c�(�)����ǗU&���*��v(�p�q/rn����a������mI�Pɿ��od��H��s0>�cvnE�����8����ܷaŸ�����F�?�9�U�W��>��X]]�����ycs��g�=�~Fލ�H�q�������]�̘� ��~p|a�õ�w��և��uέ�;�d2c^��M�ħ�}a6��5eV��x��Xg�P����Z���v��WWW�v�`N���7����$[����8G`^E�p}���m��pm���w⽠�^�Z��k0�\k���o|�3��teb�>����Q S�L�W��%��?:A�F&��h9�/�W�FE����'a.���g
,__*�m��p��zC����D��"c���K��ʻ{\��m캃���쨓B���y[b2	�����>~��g�˫qћ��Y��0����?��<.ܻ{�Ln/���N4|�����gjz�������gft'���{�eD_�Ɩn0ݳ���hW�O�]����\]��({kl�Io����'|��k�����0�ʃ��ّ`��k��dsk��!mk^�q�����чq����h������.6�0�g�:?'Ơ���3�Nl&��Ʒd�2X0�.��_�@���!(�p;a�I/��_�K�s�[�A�kn��N�k�g��FmJ�l�Y�u� �[�.��iPl��l��W}��+M
K_���\~�5,�.J�M/6�8��䘛U0� ւ������Y��%�Ӎ>>��]H唚dM��؄`ӴD�X\�� ���
���q�ĆHo������17�bW�W�&�ˤMk���2a�:Ջ7f����ƪ�k�4��B�8	2 t �{DA{P��r����!nɏPO�!�ؐ$sy�'ck�'J��mJj`��6�V]LcĚ62@��T�||��d�O�#Ls��N / �R�
�Lc��djO��	�Q)0�`S����g�m �;�ڋ65�[j��	�%Ѐ��Oގ�Y�@+�TOY�� ˜�ܤ?.�>{�7��������^/�s���rG>@Wؙ�����;��[�=����W�؋hC��� c�E{����V՝�J�2���Oo�x<6�Xs��}���go޼Q֠0��2,�W02і� up�fK�G@��X�_
�P6"�97?K��}�z|�F��ywX7�	�r�>@?c�����}��5��+JJ@�ϐz�
�k���Z�p`���J��^x��<Ø'El����j$"#B+pǘ��g��S4����ɿ���@��=���J�Ӂj�G��ok�oq\�1-~��H�S:�$I֚�y��YY]�ǘZ�ct���-�mM抨<�C�7�y= �p���� �E{X�����lvfF�M� x �Ę1��C�� �y�8֛j�[�<�V���d}h˃}~�1� �//-s\�h{�5�ޱ?�yZ��ښ��k�4Aaej���#���I���CX�uc���&�鎃8gro���i�Ć�KEĺ�8�Sz#j�/eT {C)DI&���~���.t�< >��Ȑ�`�jR~��Bl�������}FS��vm�~t*�1���4 �ͭhTl��h��BC�����5&���U|-���?����/�!p�(lp�G�I�������g�'n{g�!R0���6���6��_�6���~��3C`pb�!�ə�hx�� 4�+˴5���'+^�����%�n
���ސ瞸�P#~쳿���)�\�Y�:��2Usp��~Ն6�٘�sI��*ll�'����9���ƍB�a��P�`a�y�il<ͅya�c��f4j�!w�L8���
y2�侘��:P��{P�Ҩ��^�?a<��n�1�cE�s��S>��G?��<ZqRXF=����<����بc�Y���3���2'8'�	 iɺ��V Q$L�Qd1 :bNP'.�rKĜ	�fu�~���!�	��o���+hD1��i	+�i��Vfo᪜c�z�܍�R�A��l	$`;�F��������.�Uxq���@��P�R��%���'���V=��&m[Fԅ����/̑1�8�Kh؍߇��! �O;�
@c�H����)�׃N���1�c�����ьƳ%�<c��=<Xcȶֶ#��d�����;�)�KMf��&�r���KM %��(l=� 8'@�Y���q�INѵ��t����X988t[[�|��\4�h.q\`|ĎFpcF0-O�p���c�.�m���� �s���JV ��d�lG�/�!B�1�О_�9$���k ��6X�p
 ��@*�7J��s@0���cp6`�I����|����k�}���`�"2
  ,�s��u�7Ɍx�G=��2���y��08"sm��b�L\ý�2��VJ�\��1ׂ�Y���>/� � ������뉍	��p.-	H|@��a�uW�
�Y�V�*5�c8�ph���DKT�~.B����I��lsJM�+I�B��@����5�DNvp��ъ�
���s���T��07@�$�m2BsXɘ'�'%�`<b�� �;"9��2z���SqX���iZ� ����3�q*��"{t�"�]���wp쓦Ց�S���FjP�	�*�؜�u���Ω;��������V�J����ȼn嵫�O�*D�COY�o3L�J�2;R�g�N(l�Z�bX.�G�4M�wR^�l��Q���`g�����]2��f�Zp�"��8c�$��ح���ř��v�w�Ɨ�h������@����u���_�������o����/qk+�n>n�`|LMō�tS��Fy'�s7.��g�/�XZ�y���Y{&n���).�q3��rG����-���z���������I=������޹?} ���.}$<��~	U�+u{T�.����x�z<�7���8�$��Yr�����[��-J�)W����:���F%�H���?��M1Cd�W#0���q�
�̉6�B�D�駟�_��W^�������_?��?�s�]��8�ݧ:��𢡄"��/{�R=�����^���<����G�8&�I��m�ѿ c&�+ *cS	f��m�!�C
WHF�����!�9��ls�ż�j7	�q�Dr����w X�t� Ӳ2;!�#�����M4��e'i�ѐ�@T@l�q,6�mM4j�T�`d[���e��E��L�jH�Y��PS:n�T�s��D�%�@U������� ��	� %�sN 6�Q�T$"��j�P+6���"��c;t{�>��	<F[@���o�n�F�~É�8�=�� �q�ťe  k�������:<y������ՎM#���*Vc76f��f��وю6���j�f��&�lS�]<๛��1y�><�PU���$��g�ɛ��|�;��F�y���Y˙^Պ�C�N�������ufk�s� -��d�m'��b��Z�����5��@<� H7Ǹ�d�k����@:,b�w(� �<w9��T�+jo���� *?U�Tc�� m��	� �7�6�EȠr� z �:�� ؍>�����`����Y����<7�o#��كG��� � �w�/��  �зv;F>H�ae�Q7���'�~�t���������;"��	�8j6 �jp�X �j2�8׋��b��o�/ȎB�>$Bb>�Y��	�.d�<�hC��m�1 z�f��l�� ����\(�5��3�)�|X�DF	�1=^W���s�U�ُ�pqS���u�L��1�5��b��ox����0t�e"�y.! e1r]-�V�2�!�5Nf�|G��둀�]>�L����z5ʹ�xm0�6�`/X�`�v~W��I�g����eЇ�Տv������o�أ�
�$����Y�(C]�cB��c�[�X��)aM��q��Xk���ِ8��"� ���yӕ6����x����I�l�=����FϘ�̢�g=y��se�y?n��݆�Ůg^���_\��l���S�9�E���޲R�yڦ�vŁej�mw�o��������O`CKb��sz���A�Ã`�v�SU����2ݺ�>}��O蓟����{�f�(K��=���m��N���a��R����KbD�'�*(D���ϛ��l��痃ѿA�oݡ?��~��/���d�ǯx���'��C�E�*���R����S�v���-�2��9���2�i��Z����wy�2��K�f���r�HN��8��Q���oy��gLz8��,�žo,_q,G�=�/+x+��"̨~"^��ܣ���e�k Í�)��W�LA�^7�6ݷE�4��c����_*�����:�kR�PG�9��F���F �i�(�W��;_�8��B#49�`�\����U��?������6�a,
+s�EpN���n��|���mf%)c��)�߆uF�&+�8��u�`��kj-�`�54�{%h�~g�ӂ,���۰�,g���k�ofP�z�� ��4p9޳1�Y_S���0-_.FZ�M�+D&�Va`k]��<[�
�. � ��� ! <�!��_�	"_p-8���!����ЋRI�_Y��JE�����{'�1��n�
ɮ�_f�q�(�	��
N�5�@��)�L5��&��Ic,���ɾ0�0�`6�	3�1�L��x��	��m6En��Q4��rf��я� D���g1ƞ=}�,r��s����3��4#F�'��	�9n�EW3��zW����T6cue2⳰]�,��Tu���[qcv�����|Vd3*tal�����	���X��	�c���,3Q\�������ni�&���s��������}��l7	�?X�Њk���r[ >�e�y�:>�{ǳD_�� ��\�&��}T�&<��HBB��w��,>�H���ǵk��Ŧ��˱�`h�*
K�,y+�������+0�S�}{�U�5����������+l�p��a����nq�{{̞�f{k!���
�XĚ����Y��*g�du��],Y4�a��� �AE�jZ�T��y\+��󚹀#`�Y�5�#��w�ˇ�b��~�\�)��A��q;8�u_���e�����3�r��b����������s�U)"���ŅH5C���s�K�}<d��y=}�"#p�ކ���/g��fp�QB�H�d'�� ��s\[���Z̽7yF#F����k	z�{���ε+,�uP����_,�#�q�$������V�w����v/L�:5j`5iee�7@8�33�+TqR�ga�Wѥ`��0��)��Z4H��rp�\�샓3�\
���#���Z^]&�O�������Z
���:;�Z��L�����|iUI�������au�G<x({�܏����T��?�}��[��i@��-���g�#
v�Pߣ�L ��>d�T ��㨩�
�f��D�Z�W7�c��CbC � 8p<���gG�1����鱥���
���űj�(����=E)�� s�@�}gT*U4b��B��R������t^�'"������5Jjc%�gv���g��kE�`�u*GJ�����Tb�\f�h/8�����L��6�00��ŵ����yvfþ���Ό`�#��0��#�����;�����Y�y�x�q��pf��~dW���d��(~f/����e-�>��3��u��T�����c0J斱����3s
j�T���Z�+]��%��0G�e�Lm�~.S�u�m��u�<YX�E�q�p�����')��I]Ʊ��z�
h�5ǀ��r.Ӊ�l,0Q�h��8��uDL����"�y hF��Tб����lg�O `!��T΢��g_��3.�x�\������+�ȁ� $��[�k�h ���J`�:��Y�� reu���V�͘���s�n�K�(+�[`c�3�p]`w�Y!�"̿c�E���`��?�5�9�vH���{`2����u�����.2�q��8���5 C`-���/20m������L����  ���yh2$8���[���:p ����ޣŭ����lGc�C	:�Hsǵ���W���厦��YXa�
K��9��,;�ِ�^�(�	oA� 7��E�����1�-U�n���%�XkK4�1�11�x\�� {U_��0�X��eS��
����1Ck�iz^ ��K��$�@z��7n2@��2�����A+H����@�5��w�G��}�O�lwU���f
K �2_8��/�:�A s{$�^	�	8[mV�Z��&Ӆ�T��*Ã�����L%�:ݎjN;^�p� �>�j�6���5k~��x.�W�}�3�*� �,ːl(�g�}@>'�B��y�=�´�q��󬙣�#\��ӱ�����ky���K������{�DN�i�7]�̤�I"�.���OۻѮ��Jl��b�;��c��1�=m�_�Tn`G�"�}�r)s���oҳ';���=v��`��V�z9��Wk�i=�������Xu2�X�C���� ��6�=����Z���~��lƿ����s'�Z�F�Dz��O1V2ľ]��o���߰����
=x�#�������±W�������>9��Q+AGQB$/�D~�?��NM��=�v� h�J��!?v�uq�"ճ=%r��͏����c�n��lD!đ��I���G_��T�������xd���s��������p
�駜:#�㏙ �hZ.�Ia��V�@����(ɢ88�+�-�
����0+����{��c��㏴"�����v�m�3l@������nW 8�pf�m�zF�̕x>'N����#c
�p�i؏��6f��*R�S�=1 � ��K�+,.6�X��{����akE�`�0�c0�u+��,.�S"]4`�Om�w�9Rǵ(��L^N�]X���c��0��I]�C�c��:�8�`���ݕs����N$��1��:m���'��������25Z	��:��`����,�  :�X���b���i��p���������^��8��&�`�znf�����cI*1�(�>.Τl2�U���:]�@q�*��p=$�tw�te�2< *�,�ĸW�8X�0��4pa�1E�x�)��N�p�ӎu�
�2(��k{��������7���� ���(��0�jRt�'Z��?���q�� ����F��I�1��=��:�y>����Pp�YZ��5�e�����¶]��
����/�. �G8'�C1f ܯ�+Jt�kq���K�����/�â���h� �}���V]QR��ȸt#��
Ab.��B�,�\E7��Z��0G�Q��IqG�w,����)���j:dAW�1��|{���6B5|�Y��%H����b��8��|��А��l+T�i������fԶ�=�5�@����eWk�=ں!��"�r�^ k�Jn�1�f*j�����A �P���/`�ڷ��P����,�RL����>#���nY�\�i0
�n�6��,�5�<O�8F@ 1�i�'�cǚV.@�G�3�C���o�|±$�����I�Xf���>G�u�$�Z�}㞋k�9�@��m��<nspF�4�ϱ�p�R��F�V�G�O�j�/hO�}B'����W��Ep~��ތ�0{<��V�k13α<'�&���a?�u��x|_���c�:�l(�Б�s����F��locK����� �%l���4��r��F�A���w2��p��M1�v�;lv�E\��G�]����%�h}��w��V`�GP���>w�qb��hg|�#0�ԋipV1�<0Ezb�xqB�@pwnT���U�
�4+��@�`��pU���C�{��U|�=��YES����c&��Q�%�V���+�%��b(^^Y]�����˛����m>}���;7X�Ft�rM3��> 3����xDߥ�fD����	Z��1�� ����^Q�|�oN4?�ѮZ��1�%���Sdo%G�Ez�:�C�����{U���`
1�}N�"�m,��Kov/�t��\����X���a(cl_߸Iw��a'F23���43�|�짃�#5��T���Ȍ����<;�8��[�n�T�}�g�X���ޜ�7.��c��: ~���������8E:� p��U�Cx�S�a�[������w"�s�F>� �իƢa{�EP ��,:I9쫳^��l��L�#�B�2kZn��%@  v�*Du��%}w)�d%A_�y?u.�"��G@s�U�ڦK"5�4ƒ<ߞj)�a��X�6��a�a,#��'�3�Y���ٹ(_`��U�=���0�g��XK���T���q�ZMX�8��=^�5� 4�=�����1l�������\L�̚�� �P����\�y)�0����C�@j��^_���� �"�DYmR@�� ��?��%{��L�0��_2?r�~׽@�QZL�LS��Y� ��,
�Z��{ �4�R<[���G�7��\ss���v�n�����:f�5��M¥�5���Q���܍Z�g��8R����+�#Ǉ��&��0΄�.�?4Ⱦ�]�`i��.+��EmUvDƖ��[Z<�t�"��{"��A ;�Y���˵`������x��J��+��	����87
��2�6��q�; X&�l�� ���E�2�'�L'�b�m���� ��D���5[���X�3�b���6(���#�Hr����+�Nq�,����5��}r�A4˪`-s2@�Ip����^��ˇʆ�&��6X��cYB؈���^���߰VA"D��9�EΕ��A�`�Y�j)LY�5��- Z�F�戝�)� }^�[8�vb�{$g0�X���sk��a��Ś�:��bb�Y��^f).�Z��$˞�Z,k(�kY��l�b\�0ϣt�e�~�g{��o��dA�8��ښ%�B�V�B��Uv'��U~�X� i%+�E�v쀣i{˛+�u6��M:}ƤOO�����jsYOE�V���$���������g��]
O��{������b{��I�ډ槰N˟�m�l�Oz1a
�3؀[G6P�H�1������cGfeu�>��v����**FA�6�\�t�y��nm�2X���))�N5��t3����c��_��5�(Aa�~0fnݽ�Nz%l�;(��G��<Fܽ�(�a`Z��U�3^���f����8�@�jT.��eK����2	v��,�A�����v��@�}yÉ�F�*�=um�|q!tj���'�3�N�N�_ � ���1c��+�}zSz����KP-�>抱 ��00�� ���N&b;8�h0*a��Gv����w�}����Z��
��,�,ۋ4N��8t��=����ﲡ*�hb��{�u�L���ע�zں�P�֋���rADG�0�Dl�Ot�q��@؄`��)x��)�3��\ ��B��k��08 p�O[���������9P,�A�e���"
t�9<�o�0�.�M���6f1�D�F� ̳3M�n�ȅ�֍��,���cʁ���)yc�
�66μnÿ`+����q������a�#��7^?,`g�{܋�? ���6s�Ҿ�S`���R�3�c@?�;W�Td� �P�Ǔ��U��3���;`��R�\���U�IA�P�Nc[e�[ _H��,,�l�,Qq-��"f]�ZD��q%�lo9���v��_����h��ˁ �	p�e��$�����> @3�5݃�������+ [���C��	ϼ�6��qm���΅c�9��!�(�����֙7L�� 
�a���y�5�WWVs�D�<bV�0%T������E���IK�	�����򊲟D������ߙ�_�=���h@ߝ���j6Y�acbN����=A������.���GK�]d�a���j�1P�]3�������G"���1=|���D ��nH�����o��v�����i`��5��PȤ� �jթ�-�/,�H:�p�k�É�F՛�~`�eFs�9Y��Eؕ�laMF�w�;üe2���cp>�)�5�<���F�5Y1M����� 3�@��mk��n|n��&��s@��Ǚ6�.�)�ܔ��a���xk|\+�ū(��Rk"�c�j�60Zނ�Ѵ����;'~��L7�������Ŝ�Y�|62D�C�]��7moz{���57��j��S1�Xs&Ff4O��':p<��#p��*_��ttpBG�0D�`�8��a������׿�;�������>���`�Ԩu|@���s���*G�����a6���	={�ͩXM��J*�+�СkLCK�ǯ�J5i�6C��|�q�B%�������76�V���G]/�I\Ŵ�	t|c�g��yUj;���i��/$N|u�>*�c�4��A\��~_㜮<S�,1�:��;�BMH�#l:�Cf��ð#K* h���j�=�c�3���dܺ�%E]@��&	�w����h��
=�`>�zN���η�ڢH�s�"��� ��6,R)�.�0X��B�A���}��[�Hd���
� 3}�N/�,mP�N�
��	�] ����t#<���g��D�)�K�fC�2C'�mz�/�9�h��,Ƅ�.z�]>.@��l�����j��",4 )p��k��i�3��R`Y��x�VVd�H�{� -ړ Q.�O��۬J���g�8���H]6c�?��}ɲ1f)ß*{����m���$��!�$�i�'96_K�k������4��^���0�˿�?x����!���Q�I�}r��<Ԉ�ܨl��h���-�Y��EO�mr:<2�m\��L���~<��X��j;@N��MM&E��#�H*�F�9���
{�F`g�Ƶh/�݊Ty�K��� 6 ˏ�<=���u����<V��bye<�/8c�Ve��g;M A�I M���H�T�~�\ѢlXW,�c �)�ha`���L�5�q����������c��Ͷ��B�w�eX�LY3���`��<b�R(�9� R#��qk㧯�y�onJq��Ά!�c�x��!ۂς�tm}�}F|Yj����ż�u�=4����Β6��X`�!�����A��4�����ﱦ3�:�!��)LN�	`0�	 ��ϖ�ğ��)@��67�v�;;;[|,��Ț���kk���� 2
o�3@�~��a]y��I�,%����5Uj
2<��+��;Ȥ��8��ڪ��l!���n3�i��w�}��{Y�K�֠�y�H����6��u�϶����Dm�����>������kB���f�NC��J�2�2�ك�l~����:fΫY l�j:qX��UV0Ev��XڢutB'�O���Yڸv�~���@���������rq��?K��1=z�c����A����>�w9"�NtA���&z�Xf$���3����a�.����O�=�o�KϞ>e#`v~���
R��t�?K v�Q
c2�b&��w�w���}_�}�x���F�d�I��i�����}�n�oe/r��-���*��m_� �����IU�inn����`�̲d�� S| 
�2Gc$G\o�~�~�l�'�r��HZ��S'�~�p��'l6�v��s8�pV�ol0�*��^t/x;_��I��X��^�3W� �TӍL��ܦKj�"�`}p��`p��j�B�}i�Mܔ=�:>df~�ـ@3^�&�3�fR��u}~��:u:�i�@R�EN�n��UZĊD	�L0}H8� �q�Xop20��X�1>O�c�O\���I�����5͒�a�^e�̈́�޼V�SB�>}*����$���?����K��s�c��Ͼ(�L�d��mq��EڧY,������@�̀���~�|Z�<��Me�"��u-9��VD��{W>�ϸ �#����4=�rZj鿶gq�);��+2EV�Q��)��5�_˕q�u�K�%Ғ"_)K�3�X��سR�+�10�a�0��W�8 �����c��qO�<:�^2���)аUIm$�\�	U#�# kɶ�Yz��2@�@�#�K�c���])c���6�!���b}�e�1�Ž���nb.��W-�cf�®�x����7؊��/Æ�g ��-� ��w�wd_r啎�+��X��;�w�Q�6��M� 1��tR��ey
�`��h��zr|�R5=���H� �����vk{��_Ӭ��V0
�߼q�	�'\$7��3�vw�s�����1x>ߥ��� 6� 
� �d�6��4 \\3�6Y%|&�'|`��I"��@h<��VK�mb�x�|���
�Z!��U���F�tx���3��|��q��_T�g������\e�w�F�ӥ�����<"����#�}]v��/�sI%��4{��(���6\Bv JLۻ��,k����&OL?���-5�m<�V&������ٳMff���6�FM�������ӯ���G}6�}fk���?������2#�if�A��ݣ�['���o5�)7�R@�
f>2�-���Ά��� ��� &�_��_R�����>'����>\pΟ�����@-Et̢�� � iN��48�^��f�?����:��"M��o�e�,�%>{��He� �	u;Ѐ���*�������[����O�>ݾ{M��G �%������*Fqa��ZL�z�旞ɥ#ѫ<�ݿ�O4�F'���K��m�B�z�̘}�g��T�דkb���F��D5i5~a�h�|�Q���ę����|#���o6���p�
�ꡪ7�b��J0|�;d��ӄ!=���q��XKY���?��N@E	;Y��p~ְc��p�!K�th֨��BKR��<UT`"ϣcG�}[_f` �np�~�����j1���7���dQc�f8�KG��k�/�_� ɧ�t�;�1���D����ܨ�ql��و����/䤸3\��V
�isZ��������Km�e�\i_�Z9Y=��U����?�v������k3Ђ�<	sx�f���P .�>�tq�*��7D���Y��l��~κ�aeP� �(
����~��KA�,�w�0M[�	0lQ�y2{�H� �9��&,�\Y˒����� 2�e0��y �r��,�E"�kD�V�� к]+�%���9�ߎM=�u��ۙ�0�7�Ǳ�SMs���<g|]�~#�s�L�]n�O�Yb�Q��&��T� �!K|�c99/��9ݼyC�(�gr��\T3�i ��:`�JW
i0E��aqd�=|����@�������\���gQ3�}߰�"+⩲��4� �F�@|��LW4��>x虅�~a)
/�`0�ѯ �Ye���i�~�ؐ����c߾}��kW���B�z��I8ǃh��G@���{�.�� =�08��f���,;�t���k��������Q
 O5/���?�����R�';����#�MiŹ�%�7n�W��#$�`s ��3^�
e��l�i{{�+��ܘ�'o�\��~Bh��z/�q�&����x�E��j�(�ႚԬ�y�>��'	����Ej�<}x��4�xD�7�q�x��&5j�q�.U\���X}��T�z0hV92]�*�Op�U&rr����˨�q}�I��m���<���trT���l0J���K!�Kq�x��<���#`��o�������W�J�Q�%]IӅ݊ṁ����߇���o�a`F+�/�����0���(��Т��Z8b&n��{�}z��=����w��39��G�:�/�Cf����3�����4��O0 V"�bS` ��:a��������ݕ>M�_��@Vf���,�02�Ӏ��ݎ��y#�4�<��vhȡ���R��Y�	��:��9�OBC��9ظFh�����T٩0�q�_}v��zI7�p���4Ht�Q�zx��6ǻQ�u�|���s�/�r��\�e��݅�e{*1`i�`��3��	_#��+myLA��"÷�#Yo��Nx�;���]'���&��d�~}q����wb'(� 7��o�4����µ��S8}�~~�~�� � � �5@�mf"J=��ѱH>hp����:���l5�j��|�f�SűG;��g��Z'!E�s㳜��y0[��ZW��#���eo�z�1ìͣ�#�p^�q���$A��v�`-�5 T�'��0{"�?R�R$�0F ;�	��"��@!�r��:{\��Ŕ��P�u���J��MA�7�9b��*�!�!�@O<R�Ã?f�e��a������¢���U7A �jE\-�l6��;w�r0�R/���9�����2���Xr����Rh�a;M�b. ������+0��Y������}#�� �bh�[����K�"#_��iPhN�Ö��ʣ�<�g�i#)�� .�"����.�����9��]w�ú�vz��}Ṹ/��1_Q�S�|kkv�ϳ��,_5��-���~%��Ȑ��*��Z�>7�Ʌ�d2LN!/D��mV4y�6����79I��"�O����+�n�Y[��E'YN�Z�c��R�\{���9 }2�˴�X�j�����u9}��̹�1�9)T ��a0~[G��8��a#[�kk�ys춻t�'�`�C�j�
�WN���t|Ԣ���~H�z-l�k��TD��gg����ж�w���`+;�:�ﵬF���X�I��_�4���p����}�c�T%�R��V��C/���+4��e�ۑԱtWh��CȮ�p��hT�8 U����~O������h�f3��pj�̀�~f2o��0k�°��3��O7�3x�~�O闿�kf�߽��Z���1_�Z�z]�o6��T��3���	�$�
.���p8}0���Ü�k��p�u�q<�)�L6a-c3T�pQe�#�c����wVq�A�^��{�碂��l��f�\�{mu�3���@�`�80�������ޠ_��FB��+�0��HQ�0���A����4]$7��p��~k�0n���T��g���]G���,�N�!g�R�qo옳���X�$[�����E�)�a��iK�E0�Wק0��~f�a{O�Ɖ	�ll�$?㚮BӽA�\��X&�/�G�4����&�A�RjǼGXj8 �U�]�:�ȼ�>���k�t�
jQ\��_V�^��y��k>
q�pܢݝ]ⰧZ-8��[>}Z\����R8Ɖ����<�{��9H-R-�� /�ӝ�ﱸ7�CSkc�>p�\E��Q���MC�_ �� �	��i,����Mkf7f
|.��cAy<{a!�<f���0�6��y��o�V�I��U�3RhSt~��)��d�!_۸NKm�2`�?3�c�؂Kt.�<�1>���t#~ϵ�� �AJ�*Ksy��k�J -v� �9Z�����6�(�sI4��5�| n�
�$�s#�a��j �\K��c�>����O2Ǫ--�\c@��/�q�[px�����y���pm�a�������	dp,�9��9~�O����\�(^��N��4`4���"�d�w1~KD{!~O�g���,��J�D�󜂥M��ٮl���>���ǃ=�,L_�c�f�5
3�0�9d��J��5@?/�~���X����f���7nr��a�ʘx($�(��o��W��ΫlH ���O7�?�9���;(�5ÿ� �`W�M�4.�Dꗰy��O����a���сM9c�o�cQ���@���Z\����P$
gR5�	����_��~��п��2)V`*�o���!{�*i�vp� �0]��r�W����!}����?|M_��[�����?�10nب;�F 6�"���F�X�I?�<�3.���\��/��X��͐c��<���\���a�Aa1 A���F� N��#H���q�k��kU��������Mf�7Yϭ8��7����Pt���/�/�Q��ރAv�W�>Ҕ�,�N�9M����Կ��΃��4@���v�E)�',f `]�m�i���pp�8Xf����jP3˽:B��Ӫ{s������pL ޓ͏�fo���2m��&6�i��w�W�����eN����/�q��E�_d��������Xo�
���+*������hZg�
�z�/"�eR���̢6ۦG�7���=��1�3@�������^�{@�/@� h3�ګ��ɣXU� t��$8��P��Y�
�"��g�VC@ 3�k8�����B�R'�=�;*��*z��Q�hs�7�wb_�_�WV��CFKUM���-Mܖb<�T���lG.Ь��Q�`�V/��>K��ٟb�
�)o)c[��$!tr��į�8 6T,V�4�PzO^��2Ar��+
������1�ȁ)��p(+d�c[H,����mú��2�tҕ`���% ?"}e�B� �lEW�G Ü�Y�,u��_�}!]�g�i\ز���^�dv�q�L۴������=?&�~^�8�a���d`G����y�f�Ŭ;o���뤩k�ζ�,{��cd]��J?��T��D�v<#���4M\*����I)�� X � eѤ��Н���p����L�c`yo�V��8E�?�kz�h����h��>����}޿)��:�f<��#�	XY���g�}��
�jan�>��}�շ�桁���k_�.��i���o|+�/0X����������N����<�T:�����N�A�&i�� k 3�M�J���)�='�>����Np���o��?����_���,ժu��9��1���QY>N��;��}�7�[gtA:bA�rXUu�	�uVӎ��@�}�bvS�'�p�!'�3��c�c?m` @ǹZy��R\^�9ǌ0 �0�a\k"�Љk�� X�=Ƌ-�ۦ�[n�Y0$OR��½Cs�p�"@��		HaΘq��UxS����"�=���Ձv���e��9%�ӕ���\ڑ�*�D�#�����ǁ��O�3�r���V>��l�LRp��F�B@�ӻq���xLɃ��M۴M�[��VI�K�8�� �*/�<��W�lKJ�DX{!��=�0����������Bumt�oZ����_����8�(���e�h�@]Q�)Gp�;��z��`�dU��9�.����;DvB4��x`܉5��`���p�>�kiq�k�QH��h�����\�c�J�;)ܧ�f\;��{���9�[�ϗ=mW�Ev��v��Y^2b��O�yB�p��)��5Cԧ>���
ڎb��9*�M�=�)�Y�鱶��w��h� x�8��6��p.ʂ`�e�Y%�2�J��*R������N�.ι�ދ�a㮋";<m��~� [$�L
*��6m��J�� ��ӌ}y��N��(�d�p�Q��c|{�w.~ޚ��f�i��h���i{��k������m��bP�,'OZ]�|��j��vk��١N�S-�8Ok�7�ڵ�t��V���`��I�EϞ=���U�i,�O>�ex�k���W���?ҳ�F0�������L%l�'l0#�"� ��Ƌ����P������w�͙;���BO�=ei8!�X�HQ�L�vt��}��lF���d����f� ����`(��?������g��cʔAef�l�y"*n�3�UBA�:dx�N#�3*$�>���0fv��_�i+8B�_|D��P��à_/��6S�X#1��,
�e�����n�\p$���"��6�b�f��X�v��=vB�T�6���l��I%v�ۥ����v�}DN��������c  �����7j�/�UJB��j?�g~rc���EX��dp>q�|άʿ3p����sp�V���b#ZX�=M�t�NS�S	cp��]�\ܑ��@���R/���ۚZI���U�HR��BX�2����DAO��`~q�j�w���6c����۴R���WuC�L۴��m(��nY�hୗ�N\�I�۸+3��,�tB�{;�W 0�����.la�YA>�!#�R0�J�����@,�ۇ�Y��@�����kR���~ŅΖ��k���`��K���IѼf*q��^72��7Y���/*���:��{�Z������v��<��+@y���ʁm���T"c&������dFp�l���5�ޖ�e���~4�	��h�u0`���0" *��U�H<n�&��Rҍ���kT�<��CsI�⪖e�G�s�L�a�C���KD�'Kրq���\���Z�L�}�����;*5sl���i{5mTN�3'����I�@�nsd?�5�Cɼ�|��$�|Fw���Sm��7����覍���FA���8���G��\�-�Ġ��+��
��c���8E�+���BQ�2 u���^��zձ��ɓǴ��B}t��;��ѣ',�p�����ll�P�Yc����&����,����A�QQm�
/H���рo ��@Ш�

pP#~�#p�+�����{����f�E͑2���S���g�o�����o�lU,� �`D��iwv�(�C�:`�P��=yM���� ���ir�p<)�؇�DO���>�7��:��������t�vC��u⅚��*?��5Kܳ�H��p/���~�N�s��<�B���}O��f�]���
��Թ�٤Оh��m�Uޡ��V�� �x�+�T_�3K}+kRL�'��f��H�����������kgic����@�}Ic�x���L�������+��Y�^}fh�߱���^o���GQHv��<u� ��ݢ��!�\�q�X�Z�H�eYҸ2�'�s8@}IY��%�֕k�mW�C9m����e�o���Ԯ���Z�FX�!���?H`4����>���S�ظ�6(��>��~�����O�������*}�}����8�<R�?/�G�Q.���cv:}��<�������~����8��of0P\D�*�II��
K�>������|<)�Տ��U��@�Y�����Ϸ�%k�ˢ��YK�-]ֺ0���
�6����aP+{�X��'4ǚ�7��5@TǬ铣�5�MX��ꑰS{ǧ�+8m~�x�w�����/%7Pw�3�p/,���&����d�_����"�YN�G�i���݊�TF+��N�T'��`V���ps�>�� SPYd�*�gY�&�ɰ�$Rr~W����i��i{+�+��]��4�xG��qGЈH�tC����߽M@���F)���'�3ms�����= ��v�::0��6��S�����\���cR�4�!����)���::ܦ��s��4�-��U8���6u�����Ok���2.ߵ�e�|qR@KR��~�����Rg-�j0��\���HTq�X,�@1e�CS���Q�e�=�+ќ�<X�}��f���>����_���F�}w�TnX
�R����
 2���8'~ 8�-�����
�I�v	`�p{{38=_�?�?+��;���o�
'�N�0�g$E��ǿ�/7|�f'�����_^��AD�ЌA"��`=ae�v�m�.ϠeE睤��Z%:�]�sgR+���9PR���8�9�QGc��I�Lӄ�A4�b�n�'�m�7�i|���̶V&��g|=��|}yf�=F�G���)\@Iת���ʚC�u6Ox�s�n�&c,?�v�%��ir{���P�5فn*;K����7��O��J���z��Ǩ
,e��Vt���U�a�K����8X���%��qGތv.�R�L��7��U�P���ꯗ���� ;��>,\*�oܼ�{^����L)���eڸ�A׮��m
� *����a%��㱠����u=ز��?~��{|n � # �kY'U��P�"e�����5�d3���V��R������|��<;�r���-ڗ1`� �ѸI�����V\��� 3�J�,~8��9��y9b ��w�u�{xF������T�9p/�!e���"���K�>#̳K>��|��Gb{��>/�/"�uK}�陰ڍ���Z4�q6���H$����lA{��kg��`	�Yq]��3�w�
�gtZK��+��4mop��Dב�P��*S2e�ke�� �=Y�Oý��X�����f]��Nݳ�)91MM�w��F`9cx�d�~�� Ԧ���?�%{��9���ה1��ԉ)I�z�������w�������x�˻��������ml�
��_��MZ��A?�d�5I�������/��/s1������0��{w��$�a��D Py��~6*v_�6���zZO�˃}���^Q�%�J�Bf�.�:��'�+�A۝��x�b��d��b����=��7�����;���q�Et�1���M+��=�$�SS�r����v�Ep�k�\�08x�;��ֹ���o��R��ݼ�F�?��8v�r�;3�S��n�@e[�F�T]��$ 
cLV��Iɞ�>�3uև�ai��'s�E�k���Yk-c��}���t�k�z�5� ���(�W� .Mur�}dw��8�_�/�d�à6�YHej.��V�X�\S��W`�0ݏED
��bp���\���>櫇u�T���a������1u��O��.ݻ�>�YV	����PeG�����9���j�Mj���hT�蘟n`>�8��Zs��6ʁrc~�5���t�����/*<O��o~{�)�on{��48�|y!�-�W\��A7o��5���?�:����۷�����X5�;Z(���G�.m�Z�� ��2�- �AT��r��]Μy��=�|���ZZ^�;w��Ƶk� �з���S��d� �"�o>��G<S�7�������h����le�K��q���kA_l���׽���Rq������!�L���Q���π����p_m�#Q`wnV@c�ܠ�\���`����eee5�ג���	�Ef���[�����V7qK ��z�+SY�q%��d��a���� mz��4�N����[z������^NK@�R�b�?�+n���ⴽ���2�	��$��hF���π�d&!���͙��!����$��K*�m�l��w�])��^d^�؏LL=��7�k�˲�C��9:=e,{�'��jp�`��.S�=&9�wxR���{���l��N����H�s��ʲ���X�Bc}u>��S��_p�?��N����k��ia��`VdΝ������`(��d�b�d$pr;ߎp�Lh`?|��>��s��ۯiuE�D���5c6
W#g/���0����1�Lc�2#B�kU� �0�F˪��j���G���saȥ�����G�\�*���]>r	k����h/��&��]q��L��#\�h��jd`�1��MS.R�G^�1��9��
� S�2_����$ʽ�(� �>_gV�����:��e�M��"ɱ�F����^���EG�0����5W��#>����ޡ���M6?7G|p��4�  ���g�������
�F	�.
3z� D�`�*�ʃn��^C�uY��1���\;�����E��n����Z��C�����<m���5��]�@�z{l`��(ԊOqa��9&%X�;�w�, ޵`kJ6�$�
�r6�g��X����uv>��/.,0�;�Ee�#;���766xO�9YӸ^���1�,ɫ��݀�ܽs���9�C���ϵ�=n\��{�qq]`:Y`"�iH_����� u��7n�3>���1�/V` ��p�86^ñ���g.Ú�*�tKx��`�& n|�� C�����f����Od� }�<��/��s�i�~ڮB�	D��>���1�ܫS��x��YUy��9cժ��ld�T�y�feͤ���h�X8�Ѭ��m�s��;D�p-�f`l�k������`�l��36^ap#�nq1�������1-�׮�o0೹�C''��uB˽%qj���H'�Uֶ�շ+����q�� �����w�����iaq��c�����z%ل�)� �)������I��؞�}��f��������%w r#X�w��雯�����+z��)�y��b���ʊd�~P��Kf�vSK�Jd�� ���Yb��Ϛ֒+ㇼj"n���/�F�~��ǽ�� �G(rG��o��RV��In��I���&%D��@Z��f���XN�VG�2��s���	-K6Q0y�`C� ��`"鳾0�z*����i�ۜ���3�t,��s�3Baͬ2�]�����1���!~$B-ca��vE7}�O��E��14���ע$�mѸ�����8��8�W�?p��Q�1n`d }�#� �C'a]���qL��vdոQ�Ke�H�Ԕ�(�Qr�.�	x5�����˖��9<_Z�Wo]/���m�.ܮ��NHK�痕� �9�'aHb?������Cέ���Z��$�L��q�:H�Y��Lg�bJm�&�r�����g]y�R���	Z��9�q_ WT�6�KԼ�A'�7�u)�K%`��!�@�)Ă̸��Jt��m_cI����C:}nA߾�
D'���9�޹wg���p�q�I�y��DTdΎ:��o�k���ʝz���̈i�@5ҋ��� ��yR���ߣ,E��U�?�B�N8�y/E��Wl�	�Y$9ŷFvt�>=k2��D��q����ߝ�Z��}++3O
"������b�5&�
1�WT�,�.N�Ȉ02�(�>�{[��F���Ts"��U�����MN��	�����L���c��ʊS�����G��ڻ��`3 �z���g�k�ڡ���b>�'O>���n��@#�S=�l�-߶��JسM�Hu�T�,����e/��^ l����p9��77,��*�����g�}N���<<�[����v��enʚ�V�����/Ե�8�Hׄvrd�[
<	�c����}X���j�e���v�ѣ#��/�Hw�ޣ���O�Qkw�Ep1�_R�~�{^�P�`�WfdZ����P��]�e5����k��}K ���j� �R��YJh����+-Sv��������nG�4 �T�� @_��1�M�wF��آ��$-���#.
HWYS9c�0�/X�b�89|�ꋋ��B�	�,�C�3�R|�p<ַD?�N����t�yX���#.N8�Z�Dq��8R�}̟�u;��aNc�"(����X%����Wr�����
�RY�+Ԯ�3:MK}�[�`�m��I���R�� =��\=�3�\ئ�^�ȧk7��,�c�2o�*f�� m�"����Bl�+�w�xN��@K3�Ќ�MT�����\�k���p(|ͭV���\�:ۙ��lPY�X�ߟ��$/�l��ͿӼQ�S}����a<�p�*��_[�nx�fϴ��`Ë�{��7<Y	�Wqm���}���B�B�݂hBT�'���!����{��>�����v�+�E@Z�"�Y�|�x��Xƴ�����1�sJK��I���"�ϥ2CZ�,�wf'`vYRq�(:� ��,�ɕV�F3pow���|�$��KQ��{��٥�����6�n;j��S�q[�$�˜޷Т/~�}��'aB������w�ңGO蓏�s�#�����ӵkk��2C���TT���f��^X@J��	�~�ӢUM���64�l����u�����
ϸM�K��<��;���c�ȍ��Н�
�\�f�K
��*��1떙����l
m6��-��$�Z�B߇1��_�_��.��8��ʎ����yi���"~P��	ǭUb�����:5f���e_��6K�3�� @sV@�ZԀ��:�} �G��iv1���<4F��x��s}bh��FՋv�������.���p�8s����=z��	k`�DMEa]K���L���
����a '���<{|�����v=�w���_`�w����e��x~ �q.�!�F8
?!e�L'���i{����ݙ4�������m>��7��`�N[��N�);�^+*��T81\��)6�����Z���y�Sn�K��e<gw���eQy#^�������#N7|�/�tod�X���}�m^��m�ގV��/������	ɲ��l�Ru-��^`�. ݗ��bQ�/R�]0���0�d���\�i�ޅ�ڀ�u��v�Eu��+L��-�?NE0'��+�L�e��~�)((�u���3�M��궶�Y6��0K�su�w{��vcz! 4 ��{���E���{UZY�����4?�Hׯ����>|B�3M�=}��A:0a�4\Y]�U�J���{F�;���0�r�1nᆉ�\���H�E�Y�#^s��#y)]=}�M3O-z(E�@b=8<}�����v1�Vk��;�	J�O ����V�ֵ�y>�u�<*�����@KI��������
=~���՟�ٳ����V��u䊀�0r:���ywf���@9@I���z���حs�yj�d<o8�&�EV�!�:
 1�C����]W�ecn�ִ:=�37��$^R\OXJ��eF0������fW�e�}��([G��Y�no�Y5��b1#�Yr����� ���� p��ڃ�lښ8=��$�L�¤�ф��d'a}�Հ%�W���z�Q������h`���u	@��"�!>��D �r?k4M�9����N����|��W��������'fٸ��Ď������ 9��P�z��7��b���<�^�VK
yIV��{�6d7���3�y6R�~ k⴫�����m�y]�%��� ��`�PgvQpy�j�TL�/R���Q��Z�ξ?���m�^SK�*�|d��Q1K( �]�����L�J��P�O�( CJ�*�u1)��H�^~�m�i����5������g ��3��3�N�LR
�H5v�ݑ���W �uf�H�D���7��$kT��s�u�t��O[�����j�oR�A47M���҃�j8�/��C���t��=j�����_��ܡٹ*�bt;�������ݻw�u�G���?M?��cj6Wen��c�?�������F�� c��h�q-�{�	X���}ԧ^�7���i 1��x,��q���~��ݿ���<yD�˟�����Xx�{���9a��X��E�Gv8�h��͢B�JM���AD�Uv�g.��9/�a�Ϻ��ن���M���O��w��_�Ӎ��鸵� !���8�]�I�2��-����G�:�s�����*���hF�*�J?ؽ��^�S�
�a]s���7��v{����R��,�3(l�?
�@Z��+�$�|�{���Zp�D]Kl�G�#.���wJ/�<��-��P`]ђCۊ( �`�b�T�Y@^�2�:a����O�_.� �_��(�����p���!����Xբk�9�biiIV�:�=D���J�Fͱ71����e7M;pڦ��n�[�n|]A�!>��z��I`�>�F��T{H�W��*<���C�&'��Kl�A��!��������c�}������2HŸ��Ǹ���2_� ']�v9 w|��U "���KzLֆ�S��K��Qz=e����10v��㞶i��-����3m�Ľ�H9	�?q�R��yV��'�F]�_�������
�O1�w�]`���o���F)�;:���lf$g�0�\ɮ�-�&x/�<�2���%	�����������,�ys���܂*��^;���b��fhvn���V���������ț�[�n�Ls����9}}�������f8���kT�7��I�
6����~�V���!��D.�6��NY��c*Ƴ�y%��� r}���bI,�`p؝a�C5u!��/l��K
��n��*lv`��1���c�+�ޤosѴV)��;����=z��K�ܼQI��r�:��j��2�o�٠������F;��Y��'� l�ɢ���t��v+*���c;��Zmz�6��1�J��Gtpx�ߝ��smI�ď��1�XV��_��	x�RHp����\�0 �qM�M�s4 7�/c	@8�h�?y�ß�:���֑��Wu>7�!ȎX�Zq�Z��H3�X;9�g5�N��{{�t�:�0��0�C �#�2,�!��8�p_� ��V��'_�Rڕ�W}��/��J���4Mu{�m��i����ko�gc�8��G�\�����+��\N��Xo��\؞�mm�HY��G[Z�b�a�	Cӗ�a0�]����^:�)��]^�>�����^�=�����8�C�So�ﯮ���Ӄ`�I� ���V�P��(���`���L��qƣu1��G��鳼� Ѹv��(��X;�w޶�c�^V\�r'N��-��1�A)���mƃ�P�Y��K�DJ����Jqm�� 9� nڮl{��raH���a�ߙ��?�3�Q2b�hL�w�1�X�Vm:1�����V��V=k��$˽�n����P�^c �������0H�eXw�٠vx$��;</�.ҝ� ��齻�מ�I��ZǇ���h,���v8���/�Kz��}�/i{g������h���K]WO˸���f@
@d �z-�\�Z擾�c�Q\�U_D�d�0�������g�m;~�����ɏO6����L%�
E����2�e��ѪNX�s��)��Rx���� 8G2^�ǉ��h��L����Yw���H9ԕ�=x2F��\�G%A0�p:)n'�o�X�Ԯ�% �Oo�:	�y!�'���#u���\9���T����c���7XK�y�)�{�H1�fS
�zI�>�yQ��H�5�!�[zggÚ�`�ϧ|oV(P��&}�k�D���:4ᥐ_XNg4�u�)z�(��+�7��V��`G6��C�/�,��W��4g�؁�Z���a$@񒝲�W�Ul���F~ʞ���Q�.���V�q����.�7Sխx���i���MQ#�L�8�
��
��[��9RFCb����>(%��O�ogv�8����c���z��=�����?B��4@pZ���7ao��^ꄟ�g��ul���q2%\�8��mc�� 8���G������z�1�,p2�"5�3�V��,�q�lȆ�Z�����E@e��i�-]*l���tgI���)�~v�kg����d� �Wr�~Q7!^��0�2mo@x��X���E�s`��ppe�*��v��WV ��% �S�+e��7�g=)S�eT�W�9XC1n g�6�T ���'Tkӵ�ez����tm�eЪi{:96��Vכ>=}|@+K��3`|:�u��l?���%�Z\X����gL��紼�@3��s��u\����B8p���)�K)�����u�;4?7�@�1K'$}�	�3�&q��pW�xn/ �,鰷�OG�-~A�E+X�)�>�i��]��>��"�\�������H�P��}a�@X�ۢ��4����	���I���.�l�����ło�s�L�$�@C�����
oqp������x�ҵ�f���c@ڿ蟞i;Q������n�~`7(z�m���l3�.��J���6�K�͜IxT�o�
U����ͷΛqvC�A�N��`;� ����B!Aܳh�gZ��젣�z�F���s���� 7\��	�yk�9�X���1��Dv�
,�_� �������0�>��ΊDI|.��䒵�e��ӆv����ii���{��J���j/�?G��5:#?�?�S�P����(A
Z'Kq�w_*�A_1XLZ���n�d���)j�9�A�T���2���r�#7���1�yD���+�9��)d>
�4�o��츲��I[Z����ņw�����22�?ß���v���MИ8aA�1c��G1��}ECb�$�/�.4�>���LrqbPܙ7:q�u���6�����6.ž\�����>p�O�ѴMۻ�^�T�567�	�W�҂x)���Ϙ�Kd��&�*���2� yA#gٌ(��7s��D<���i\����0fb:!Jm�Vbj�3���h�B�"��m�B7,jʚ��W���0a U�~���I�M;��\�j��p �<� �h�hyy�%.���-j�g�i����v�����Uk7���%��~�n޺I�15sM�������� �����,ѭ�7��/���gZY^��Օp��\q��� $:�Z�t��+�\�(&�����a�>�ɀ��(��g���#)0��N��3c�_0�S����s�E��Y�I
I�dT��D?�X���B��4�����9ޫ�5R�����.����I��3.�G��~�l�\ �kk���u@�������L,Wb�fk������iJ�<?�ƌ�c��(�]������,K���� �<�X���9st�r
����ұ�Vq+�����' zn#���y�%0�in^
phfM�J�l<�q�֯��sǀd�W8��|o ��.=�%��nd+�Xb(�����χkS�`��X�*
�W����;^S|��]6<8�k)��7\���u<�:Ǐ��s���ׯl3���1 H\\�.])��8����{/Tje �V>�ν��Ë�=g��w����?��}�S����$ ��@mqu�#�k�a9#	:s!W���.�"�>�:�=�},"k�;lCL�|,�=��N5�S����x�s�vΧ������R��/6��cO���}Ԣd��-��N�����S�Bn6�Ő�E��Q�n��9�w �c�vt���l��ƛ�fpe���"���Ԙ葑k�\��+�bT��a{@�a�6�8�Jk}��KU
�wfb_�K�q��U�פ~g�u�%� ��R��|e�E<�3�,'-��8�6�,�&�\�:N��l� ͈!)Sy��5�'�/�,a ��΃,خ��<)4����Ξ�����qKIv٨n_�}���"SW~��q�I�m�ުv
�rv�v�dߘ��)� ����@sG�ף!��ZQ���W����� �\�bHc��;���kWJcy����s���װ?����H�(gH�R"���m*��
���;;3#)��n�[�J�]`B��_�t�J��)0��V]^^f���ş���*��w���P�9��Ζ�zv���ۋJ߽{��>�?�Ᏼ��E���z��,S{����<O�7�������;���Cֶ]XX �{��4z������:�k`�')���������wցz� ��V���{ ��ȕ�Qo�X{�%�9������݋�(�_�#}�����W�%��{�C�����A�ϪG�z�V��{�{88<�53k���n:"1t�S�޷�c�N0����3�=ݢ��M��_�k�n���J�����t	�,�N�x�`8�iw�� kc�>��!������yq,0�y��@w����?�:��c�Lȋ� � Ԛ�y��@o�5eqq��gp= p�8�``�d ؅t>���@�W��-p@jkk�����T�+��p=�s8��j=���ۆ�����C���Zt�2fK�	�|(���0���"3o��9en{�d��㒚�6�r�ݩ��Չ�=-e즁P~�'�9�=-�Mz��`l
F�.uڔ!6��@%�����y�0JG��_n
��Q���M�֑��s���h
��S�w[���� �U�?�'�`Z���b�Z��
��q��S�|G�̱�R�����Ĕ�)��I��HǸP'�c6�����~͆�+�v����O#��s��]�U��И�����qJ�N�;}�V�}\?G)�\��Bx�����8؊�)�1I�)R�ϊ�\�}?���l��*p6���q�O
g�9�wb���Phr r=YE
���i ��\��9���b����ﰷ��&� �� NjT��c�k T$��6z����Ѩ��3v�<�>�~���>��z,�lN��LԈ�Q��y27�$9{-Υ����N��T������n�J����a�-ؤ�gi���"�y���[�\�G��B?Z�&����@O�����K��g�6�Ǉ����3����2��8^����"t{��a�]��VWVܶ38�G��>�	9f�s"�>�Jl��1j������t�����u`ˁ ����4,�VӠ���4<^�_�s~�|�3Z��[?d���`�ݪ�R!$��v���xM����桿9�4���&�˝���kk���{n��t�nWy|�uM���W��w�}֜%��vC�R�m�rh���ָ�v��^����qS��`iW
X�ps�c-.
1�a��j��*F�,u��0�Ol����z�j��1vx��9��L0����v�K�G{�>^fFe'L�V'��R�q8^�>��v0�`�-��ƍ�>�K��Mz�9CO��0���8G��-��V��oҷ�����n�͛��H:9���߻�������o����yc�0zR��p ������C_~�'��ڦ�8
Ć����g���}Of@���T ��"�e���RcМ�晻�ug�f>DV�lhS$�^t�y�Bs�!cXƯ���t��d�8j����d�h�ǐ8���@��?c�}�&��<�)���\��N5���7�L?�S���J?�Q�}?�
3M��ܽs7\��o���?~���'����<;U�-�<|�oǲ2+++477��Ƚ��#���̅�p�A=M���J5c�a;��O��w�}�}��ǟ�{��e#�)����Z0���52��^g��^��:Tpf�"���񐳓�����E ��a��F���L���1��h��p̬�J���^X?��3��}g���3{��h�ڱ��D��h�T��d]Fr��(��e5 6ܻ�>;��p��\2l��*��R�n�q޴���g�N%�Aa9ɝ�f�2�[Ǫ_}	�\Z�Ņ%��V��؀�"��?�8�=-
��*扁ChpLq.<W 5��s�,������X�5�@)�'8�kkk�>Ec�Ǭ
�0�[���x�f<W��8�8���Rp�����µ`.������Vp�x �F���l���@�B�A�N;�A�sK�ZS���b�� � �9��=���|4&��A��gϞ����E%����!�<G�Y����~���e}��JZ�5�,� ��������{ �4�yZvĸ�kG���pW���k�jzo ��W�e�s�=l7�Qruu\����s�h(�?���J7Y�6���Ŏ�"�S�^��
)G,W�juu5��79 �:��M�p�x�����ғ�OxL2xY��u$�׵����;� �X����DM��a�cO@�	�?h�yK2ΰ_���X��"Ua�.<kd��5Q�����S�}Y�?[̍'O$���������e������>_�a�Χal�:������w�,�߿υ�b�gI�E��EF/y��e���V��x ��`?{��JoD �'{Mf�w��Ez1n�����'(��2[�������{�'�\��g��Q��.�?�d}��r-[��a�x^�� �X���(l�� ��������
@��,#�?Ga����]r����@ṗ�!�W̑[�n	`]�{���ޛ6G�]W��ǂH ����YE��6kR�1Y[k���f�E�f~���1�/�3֚6�L��DREQ,�^�r�D���y��{�?����J��H@���[�=��s� ��>��!�}��_�s��l�������~�˞�����{�)�k�!V#�E���]K��Ǜ۬�H���g߿O_	s��{u�>�=�YP�8װ6�.$�!u3���h�k�	�����L��ób<a;aN̳>�O��ӧO��� ���}�c_���b�+ y��4�}?��Q��ѣ�,����g��%׳���YX~@b�c�_�8��N�;h �3b�s/���l�gQN����נ}{��x�����ڀk���w�לg�X���Jڠ~��s�{S`S�xoNX��E>�'��i���ы����������9g�����Q�����lVt�0�]�^+pVh[��"i��e�{�ڄ���e�VIPp��fy]��>�9�v�����0:��`<����h�����H��v[s}W��� ��snme-.��}��W���ڢ�y�ft�vh��ȼ��u=p���q�q���K�h�䎎*	�ޜ:E5���G��j4Ԟ�_޽��ݻG���K��q���8��Q�ׇ����#���/,=T�,��	�j����������S�ug��*Qb�:�U�y)��\G�!���lׁ�o{p���"�+�y�v�O�?�I��jA-(��ܛI�g�MH@��W6��^S���m�!ɠ���O]#���zj,7?nެ�A��^4�t�qn� �� �餂u�S�50���/�-�5��@n��Eg�~\p&��ty���0��Y�vH�A����f3?8�Ж���$ 	Hp�Xc>�L�� 	�!D�Y�x>��3R�g�s��ַ��1�D8*h���>�?��W�C�����'y�pOu���F�@ȑЙ�ל���x��Xjg�������ce���O��L_��:t�ٹ#)"!8M��<�ߘ��kD9�Ca��1׫  ��C`b|yB�a� �躚����{���\|ֵ�x_�rFXWp�w���wp@�n�E �d������)���T���<������l�YeD��,	 x? �<��鹺�3�s���:Ŕ�j��j�@h�?�N6�+�% � PЎ9?z�L������L���&�ٵ��Vb(�xpR���\m���4`8�Z��0~ c�����,`����g�߁͈��� }���I3)T:r�=f�N � �X���!�@�#�>C��7���S���gb,0�̸P���c�K�"���`��v���>Ăh�˱�1�;Χ��y�}��ώ��➺��h�����m� �Z�I H�S�o:�-o�����9����	(��4g#�ɉ�ɠ^\�dbm"�\X�!���6h�N�H�a�bݒYZ3� VX�7�~pO >2��s�`���7n�Y��3*���-��2[����g�"N܂IN���v\���9�*ڮx��͇�;�QYg��u���~a+x.R�.x���Ob��f �dB�-���b����m���ޥؗ�����Yd�������D���Ek�c�mg��
=S�@A@��5���k�v�Ho�,Hql�������=1�u��sE��c���s��G�c��I#^`5#�-T��9�@�0}�����*t���sϋ�~�2��67x���+��ٱř�W�m�ۇ0���0�O���0���-�+����9~F��Yч���Q��t"R�/�==$k��w�C�u�7~��?@c쏰��z,�^��D�����.�/ p� 5Ʋ��p<ﰏ�:z_�7A���T�C���W1�>�#I���TN��.-���+�_b{I�|�|����.�֧�&�n��g߬�d���u�?�V;~����%r��3�>�KO����̉>A�� �s�pܦ�k�k=��~X�}�L8��y��I����~˧D2����
z�V��Zym*���-x
#b{:WK+�nii�]wx0qO6��Nt�.>u}�KZ^?��?'�������o�����ٟ�������
�-D��{�=:�#�e�����ݝ7�Dc�p��h�L���,j6�4�0Z�q�8:���7��s?�钛�/��,e؋����|�~�Ͽr7n^'�� ��7G�y�m���lB��S*h���J�T���S�iӦ��g�0lڽ�<M��qt*���'����6
����ܭ=�*M�[ZZvW�\qw�܉��wx�Zh pR�C�3?X�(�.���ᩙ��v`�!|�0�~���d���ۼ�7�Ӑ���t�E��B�挩���2�x`~��m�Ip���q�kS�c<���qC���4�ȜU5}��M����ݽ{����K�LU$�` �6�/�!��T����$�; ��w�����:�ا d��h��Ŕ��헙��y�&��.��uh�(�,X? �M ����_�=�)�TȊ�?�,W�'��Z��	p� �p	�@���h�_���y�4Z0�6�#G�#|�2��l�=>�g}I��5
P@X���I<���5�3�Eu��V�� �0����C��1tB�!����M�I�q�_8�p���^|�7�|ý�'̹��v�z�liC.��;e����� T���ꮧڇ,D�n��އti���dwK:l�Z�>����_��?��N?��鮋�O�}���e��� kleq�c	� �>�ӏ�Tv�X�;/,PY�~)�����S2ɬ&�x�R6����3b�`L�����>���<�>'gҀ�G��d�>�d� ��֗8?ښm�T!8��>�B��"[ p�~ Ha��{ �.?y�wds��Y�c�D�M�GSN��@�y#,G��[���>>�`r��l&��_}����}�]� m�r�㜼��!�>@5Yqm,.�=8�J��#�����?���#��-ڐ����X������{ZL�-8��Np~��x����3�����RdL��k �Y�	E��z��e� �ձ�3	�nN�Ii�g�kxn�� ȇ��9:���6�oO�\��&��Я�#���{��n�)�l�/�޻+�!q/�sU����Y�A�I������l�r��G���Q%���yum9�=0��"iOkޖ�YHF�>�l&#h�@8��B9���(�\&�h�)�f�9 B�%o&e���9��ƌNv���fƺ��i�KԣA��#��KP� �U\��<؍��v�?Ԕ�&��øg!ЊL�geIc~����3Z/O�J�G�o왰�HZ��	%�����i��3�ƍ�?����e�6��g�}�{@��(�8f�68�l)B���}�q�z�9�=svo_�0��Kk�>��I�YMq��=��eQ�O8#�)�� �!�y9�KB��Ђ�Y�&'�\���Cm�����>�gu�kx��^8UcA��ټ����DOX��q�笽��� rq/@7Jƹ�J~�4,��˧�K�o�T�����EǮ�X��/�I��UE�!�#�������[]���8��y��]���g�铁�z�[���>vs=��;�����}�ut�?���F<��ODӹ;o�����y���Ed�i.E��}�ƭ���'��=��A��jR�7/ӰpV�}��7�%w�,5غ�?t��O������~��?�u��|�&$����,-*g�����{��%��Aj���`�{P!�������$�&M�3c��I}V@�^�e��8�o�z} M�U����%�|~(��z��Q�LO�I�8/��ܜ_DG�<�Fӎh�ȃ�T���7��z��kub�ĹHv^O��_���DYZ\�̵$�p��6��Z���6v
��`�lƵ��\�zͽ�0�e�'YJ'�>�|���83qi	i�8��W������C�� �,�.���O埤�M���`��!�3�������T����`��sλv ���k@� /��`~�n��s^;.��D����M�*"������x3��Ƙ�	L�86�y����ꫯ��;̂&�(���qh�;^� �)�X0�>�ex�B���6�]���P��!@`7��5����h��CaN
x]D���C*��'@e��k����@5������~��%i��C�j��z���,l	����4y��g��&iەN%���� �4M=u�<kkL �v��ڙ s\��6(&�/r	 �xF_Z�9^0�A�q|�B�p�����^ !X~#���x���y
3�5�i%��\�ޡ�J�7��OK/�6?c=�  ���q__�����S�v�uf�e�T��|�B����]R���d}L[i��Ʃ}�s�رy�-�;��6� �G00�q�g�ֳT�䗌}j�K�&�� �p��=>`*΀��e=� *��� X��7������!�-��`[�π�+�k�ֻ���h<J�I���SNT�s�����C����������" ��C�1��C��� ��+�s�ظz`����e�oJ05�%{\sx���X��I���IۙL�	�
�X�Y���Oں�	@�(��M�~�)`{3�FG|��+d(����HC�_��3��yM��A7�l�zR���X���g���l$�:iN��zW�^��N R��0�R��)����#�%��ReP�D��
�(��g� �y��¹��J����c2_��PZPN@ұf0���n���,���=�X����Mw9�Ǚn&��k��P�fT���ڿyP�e��3a�a=��6t�]죓����3���q�YFBx�-��j��2&�.��:�ε1F��FAj�u(�A_��j[;���}~�7��8���'�#����Z��Aj|.��-�%�3p���~r�L3 �;숄��6c~TvJ�8(;{��\G~$��~ə\=|� a�7w	�V�Z�Ў�lD�{h�t�L������X�o:����B$lQ�lr)�݉�L�JS?�����:�р�N��Ҽ[�XpG�w���U�<��������K���{n�$,4��?s�������!`V�2z���ͯ-Ssiϖ��,�ݕ��]���-I��_��tQD�G���>���lk�����N��ub��?t�~�K�������?%�G�L��Z�k�����"��M֤w��[ �Ц�O�����W�΅�&DTJ[,�j�`�	���Њ�- �t�C�}�ܸ�N���_)F�������z�9��*hA\c#�����mX��N�zzXy����n߾��ǼІ9c��u�
/���)�z�G�q3]Zrp����.����\��nܼ�]�J�ٞ��p�X0� ����p~�P�9L]F�$
{*��<�9��a�[�S;�ƿ/Ŋ ��5S�9[��X��� ��T0D�֝~m�������t���`-(�n�;2B�B��?���K�����
c2�Cً6��<�d�s��K�t2F���b�u*��Ǟ;�XPwq��*^G�3_M6 �g� �l�=����L��&cL稝}X6&'e��{���ޯ���"wA��2�|�\ ������nA��"VX�`]�3�r]�qO�up(2 ���T���U����)+�ΊOZ��n��5ڂZ�V  ��K�_�,��{,��k�r'G�I��a��G�N���J�Ga�Ty�W�W�v_���PGM�1��w���AZs�{�pM���#M5�3ͩ́m-�HxHP�;�ڧ��l�|��K�.i؛L;'����517�2M
��݁��{q�}VZ��f���^_t�g��h��m ��1}��[���#]>>�>Y��ꔵQs� W�~���@]i��^�[q����y�� �I���q]>��`�EMO�)�Vp.�� �����״��2���z:Y6���� �Z�j�ș�h݇�T*�� ��:H�(����u��k��}!��ޛ~u�-vi��{��4̓@��J3�\@à��r� ���Nm��$N����N�7���i�9�cj_�;	��˾�sGNX��֔�3��@�a���n�O�l��]S�����]cn�'5�MA�f��\��!�9�8 m"#
���g��K���)�>�݆�2cu��>Uk�����w[�Ȭ��⋺�8�c�Y�AɊ���H��z�)�P����I23���Q�420'���%���	�Lsc^[�T���+W��ey�#0N:�V� � k_4�{|F�=Á��s�Ʉx���b���%��Un�g�����^��9�9�BI����}�s�Oi,���옓�Y|��Ղ�|���yJ%�3?4��I2'N	�Ud@^�׮u謝ϛ�hmK��)]7�Y�8n���Pi�n�BzE��{�����7V��M��?�<����>���	Y�%'��\N¬/@�ײ%\(��X~�&s��=mʦud��f\T�	y�yRz$-�-  l�x,�8��^��.�����~D���֡���p�bo���������\���)�Vk�x�  H��|p���XuO,(��������/���W����>��o�ǿ������;>'�"��ſ��������>��3jܾ���t� v��hPq�����ܩN����2|���y�'��#e�OY\��VM��R�-����9)uzJ� �s��[O�I'Xt�c�����$���	�|G�T��d�G�U�y�H���{��︟��R
���x�<��tшǚ����'��}�)�%����X!���o���S�^;q��oۨ}]��� A���3Y7�g���9��ej@ ���re�
ѝ��N�0�(�]R��	�����-�\�-S�{�h����y��Ta���Y�V Ԋ�S�,�J��D@j=5��#����T;�&�ic��a��|8�%���`!}�k
{w#��I�O����L{��bw"�1Qf�jg����xN�!�smm��`�	'��`J�-�	h�25  ��#s5:�O�>!(`��l����'�q��]������� �Z>K��)�p�<��A�k[`Y d���dP��gz�3���&�i��� ��h����Y+X`�L��~ !Oc߀mM��#�DG�R\3�(L[�k� J������-|� t{vi^�<I�&{��9 ]�}r�5�����`�!Ʌ����q���=��\R��$��H櫜g�J���\�*@��ż�>���?[2�ϫ��6�5 ��Z���o����}�Dǡd�Ԓi ��q���0��0��z@�~���`� ~�C*��q�;�� ������Gf7��m�G�SE�>ѹ��RS��/��ޫ7;��"�d�=JӀ��l��M��j�j�.;���Y��w�M����Uj�I�ǽ������;���LX�=	¡��س����c? �1�~����a�0�ù�{��7S��<	��1���]��\�W���9(�g�	��}�[�Ь�Ny�v���o0�Y�u��S�f-�H�[�u�/���#�7�Q����lZp�d/D�f�υ�2�p��Z ��8,�8����[��2�F�a�����l0)[GA��0�FJ@qS�װ1�!
{V��1 �b�&܇�(l�5�ev&H�k�$�&�ǰ�c���3v"�Ԑ4!�Z�E�̊��������diPsyD?\�/�ES�}=�P��k��,͞!�R#[�Ã�Č�=��߸Κ� ����}������8�oøb�bNc� 0�3������JP�S���O</5����PFgߧ�Y�R��H����y��N¹3H@m���8�����T��~���t]�1��ư"Œ�cD��o��3)K{=y��}�I�ߣ�O��Xc�o�+��o��Ң����	��6��uN4�����Ἓ�R����h�L��:�g�v���}�}�ɯ�����w��4� ���J�t�^4���i�F��V�Vע!��1�a�h�xc��"� r{k'K�4�.�_r���uj���[� ��|��������*������lRaqy�]�~5:7A�#A� ����7u�L�o>�v������Ӧ�� ��@�i������O7[�
�8�n��
��*�,X�n��z0��Ӝk+*��x�A0|�Tcq��Փݻ�8��rͻ�� ���]�t!�RpYѽ��3nCr2a�h��4�`d��?�3���%��>�1̧���	���pc!��$��Gg=:i7�]��t��u�f���;?C�]�W�ߓ-w,0fk���T����O��+z��f\@�F��eg\���q��+�˙���W��|�˂@���J����Kً{=
G�a� SύAt��B0	E�&c:� �_C�� ��U��  �Q�9@8I�V@_+��y(�@F %8��T�aY)[�
̑A9�4�R�t l���+�����z��,���&�P+�]X|.�<�c�
K
���C�~0�Jp���)�O�Y��}ވE�FI� �4��`��:���k�EJ��01�e�zg��5ɚ�P�R�
�"-�˗S  �Ք��&�N'�U� Y���wG%A#����!T��n��H!��$�#�Ϥ����0-��R���S�v^Aߙ�Ce�+�Z�ݷ�-8`RE�)h�`��E����
&%���׵JnT
�I?� ����G� �y�L����u�=���i��5ݮ��f��%0T%pI�@�g��aL�Q�6Ū���cXW�R����>,���b�8�6.o0 �,�e�P��/`k�@���µ�W�_u��q�B�	���&dR�>m*2�1s��f�7�[ R-. �5Q�}��1�&�-;��[*�~c�[Y]�u�3�v�Ҫ��։��!P&�-���'J:!��M��Bd���l&��(��<�8�u�zV�SX�sq�C�Y/'��{m�^_$���a��Ɨ �lB��3���v���l��N���K���y����c�b��\р��`=cN�oL1�{g��	rx~.�OZٔ�($��l���R"U��Թ�kә�}���!�K��|���N���h�(P��ި!��,6���h�[ �EuǦ�<e�}��������Z�}<���d����fs�T&1�;�� �/e��o��G),�OA@�2n���<����|G��F��ue�Z-�?�u_�`~����$��2۶�vYr�@���ʅ �w��i'��B��W` ��>����.o��,��r;8��IHX>����62O̔x���mi�s��~b7��n���w�'�{�^ek�{���{�f�r�e8�"��Is� �쏝��,Im�;i#��#Մ{naq�V/��խ��z2q�GW��{���}�ٿEC�p��F
��C���*F����h�1���hx����DcN�ha����;��,�re����{�<��ϔ8���knߺI���_��Ѯ�v�J��hk.�{^q�ј�T�yX5VQ،A�6�\�M»��v\6y�9�(�9�ӗ�,�w̉4_ƞ5WݭW{�lrl�p��h��`j���6Ǭ�wZֲM}�LƳ�<�*pͱ�u��>��m�p�NO1��EtF�q����q7���
M��'[v/y߼�=�4�ǵ1��ފs�/�$s���m�00���WFgil�4NA�h�É��~x�Ogȫ|��[�n�3
ME�0�_���Нe��P?Ʈ��iP9��s���ݷ2@(74/>�ab�l��א ��b3i�^��g�e�
�?/xO���Jٷ� p���QD��pޠ/�`��_|N'�@��:�
- G������hœ(R	iŧ�i�����+\3�L�k��
�K�EY&�V�>ދ )@et��b�����!k�/@A�	P O��{ߋ~	0���@+���2p�҇��qJ�s���6����,���0
�`���7��Z?�i���d�WUf����N��A��� ��S�?���wަ������P{���� Ȁ۫��ާOէ4�V�V@5y&)��dwoW�'�8K�������&:��H�/	�n�֦/Y�a�؟�(�}BO-��]�8	x`^\�v���<�g�) ~��=O�3R�Z��=�#e�c=!Ӌ?�9�\ h�U;6����&[�3����}���@�Ӡo����m�I���y���U
���&,l�M�0�<{���3��o8��+P�;���3����@��	Ra�C�e�����jc9؟{
�*��"�g,V��� �4��	���%kj��u%{�e��H��kϕNr%9�FV�h�9�q�6P��R�)4<�P�Jj˫�HUH��ڜ����@�	��VF�BL��5���{/]� ��pS�i�R=ac��Uo��]^�{��+)k���4@+U�?B�ʶ;k	�*��>o2Y������y�Ab<c훤������!��;�1�&�_dVdE�h�`���L�-�O�s8:LR ��B�8�_���Z�-RL(th�\7�lvK���(Z�}Y
����}��&c9��7�x�H�f�Q�X�[_t�ܜ�"��e/�+K-�+�'	�Np�����k�K;��;�6X���"�J[d	���fͿY�Z�s� ӱ?��_���"~��%j����^��-��`���~~�ُ��o'�;���!�$_�N�K�d��>a3e��I}��E�V�r��H�F2j����ه�=#�fn��͚
��ώ�郹i/�	]B�e����@��i�U��Y߻l�;�;k�c��v�5QT����(I��E��T���q��\(�N�1#L��.�E#U*j�S�_��-����o�Ѕ����M�H�'��`{�}��/��̭o,�7W贯������蘭��h07�m>|�m��`jTt���Cw�������6�/�?����������W��������ڪ��������WnP��8/-s�E[|ƨ����3�cˀ�^�2.�Gm�
�&�i�)��;mU��g�tg�dsT<��~��!i��3&N�H˛H������S�ߌs��>�|�%��.�>��l|iRJi�{��I-�ӓ�ɏ?d� �u� (���x��б���V�E���F0p\���xn��i5�sV��|B�E����۷.�߮;�ݹG=(�~VZ�v�c�s�9�)g�uHy���fF��$w�5��o�t� @�"9j˂psA�B!a��[oQk�#m�� p���}s�:� n�2�PDS���5ҽH��6�v�� �����z�BkV⋠��t����������@*8�x��pj��(�g�9������B�C���k��>k�� j��]W0݆�1l >���
)N��-V����: �O�-:I�8�'�M
CZ�P�gH��u��8+nz���C���#Քd��{���yi�[d��A-��x�9�2s������ �"8qxx���\��o�| >������\@`�`�P�n�))B6�醴Np�BsS��B���M]��`�mY���w�8�,|��7�����|�0 �T���5��"���E�󔠳��Ԛ��Js��^h��y���z0y<,X���R]lX�M(�I��D�m��9�l;��׮_#[�[������ͥ�WA�t��x?��y+|f"�O�V]',n�57�=�̡2��{��O�1V �����/X6���^p%E9��"��gP���a�<nam5mƇY�\^<Z�����^}_�ܱ�����VN��l��X�A��>�X�� E��֞wӧ���pL��E��� i�(s,p�� +�S��, @��\��e`�k�oP��@�+p!���E�q�:�K���G3P����Ÿ� �b~��WV��I �Xۍ�kpA��Nǿ�Y��2@0(tO�f�H�^�}s��K�U}&��C���8{(c^b,<m� �2�x ���=KOK͖ ڄ绌��T�������X]|�(� +����RX�����g֐�9YQX)��OۀzϣqO�����/Pj�{։1������Y<�V�%B*�iʹ�ϒ��hX-D��׍mE�B
��r?#��m�X�iB�9I.&D���*2�?v��b�f��v����_���]4��7������7�_s<3H^����`^=���w�p�F5�ɡ�����5>����Q�YW��� AVov��FGHD��Ѝވ��8:��}7iz���c���ꗿp�n�[�n����~�V��t�
T���(�*�MbP�8�?���ʼ�z�{뭱�|��]�I4�Lg��/X��z�����G��}���������.__uK�[��\�>2P9��L�|g��ߋ$�h�|�^���H��`�Ss��{�7���c:�E��]@��`�!�R]s�3]Uw�����*׫*� =O��H�B���t��8��R��c�A�z�]���Q�#~����[ҷ.ҽؚ��f�sp]X��fEzH5 �'�ؕ}�0�w���<���Y��{ %�4b���%2<�w�nE fe���9 �rk �\�e�ʝ�ޝͲom�"��=-W���u�\g���o���{��^d���/�� �]?�P�>���l^�3��z��ܷ����A�֘k, ����3��q9��#�� �UZ�ȴ6鬁5�ɡ�Mɧ\ �!������|�3и�}Ę`��9�∎����W��`��C��%'��h\�kD>bHl8<W��M)�^
Т� @̫f$ �A-���	� (������/=�ivb���'��}�b��y� 1LC��
��v���Н�u�|��h���`$`���fR�s>�>M�ׁ���qX�2�z ����n���ZV���	&Y4/@A�Rd�ا#r�a�y `��Ѻ�JL�F��
�YM ��v,��)K\�@00�ګ�]�)� a0����>�9��b-�FǙ޷iCS�ZP6I{��X��T�9l��+4 ���_&��\Z{f[x_h��>���\�C-�~�D�샴C{ԃ�txy�RY��9k6I.钃=dn��7�{����#8%z�=уN�R��٠�'5��T�e�� ��;� 5�4(D�/��z,H�#�k����4��ѐ�$R�Ԃ� :M�ƀ�B�$���y�>ٰv ���{*���	�%Y�� P{������H�ӆ98��ǽ��Z��.�0Z�B_���0�u�ˢ�p`��i���b���Rxn�Le(�9�\� �c�Ӡo��<ú\������g�@j�$��̊0Nۙ�K	�����O{������u���1�s���܉�M��M��O���v���|d��N��ּ/O3#D�{D&=��܊<���&Zg@��:��7D����͆�ʼ�S�M�#(p#A�W����}��d�s��ϚA�A�}>����Vhڊ;�;Jt��ɓ\�?�fV�L��԰&C~z}W#�|��#�dF�tR�����:����r�G��NQ���N����Ai�E�z��P�8��i8�9���ռ�n�X��!7ʎ���1u1.����r�R'�ʹЄE��=�0������ݸ]���ew4ޏ�iܳh�n=�v�|��{����w���?�Sw��{��;oF�e7�y^Z�s�o���e��s<�K�H�+8�`���Ƶ��=�ŗw��-�������ן�����G�}iѭo,���r��\�p����a4~F�#�����q����YAjU��׮=�~�C��O~��U�>MAή�8/��d�T�Ft� 0J��eq ���U=�����T��haG��A�M��#?���:p�n���{�C��8��A*�_F��>b��g�H�9��9;0�_Jڏ���jem@�_��w�,5�vN���5���(�|�}$����P�L6	F2>Ê�u#'��W�ҡ���n?���/�_��:��ͨ�b��h?���-R�;�~��l ��^�}7�4b�IA6IU'�2���@E8vR�R��5�lR�{�� � �	���Wf��M*����=�/蘛v0�x�����Tt�q����X)���o�t����������z���AH)�h{��R
��t_�	v���stR�6�nOA��i,�(����1@�Y�l�f�a�-,ؾ+ι��>���������r{T� �4"8�=��bN(�� �V����2��� �h�ʳ�,T�c�  �� �������M��-���ю�������&�]�p� w�%_UV�x�惿��-*P��xF��%I ,ż��6���oaa�6
�@4�G����:�xY��`[׎ɷ���w����Lnĥ��J�f	+�Ќ���V7�;���͇��r=�[R����1L�{�,��
�rL�����7���$���u�4ؗ&¬G�1ߛ�k_K�=�p��V�M��O�2�d�A� �&�x~YOEb�X�l�t6׹��60�M�I
�����~b�S�^%}pmcU���q/�>�V7�eô�0�ڇ²5��X�����}x�wı���uoW4��0P� ���MboXx'�+���g mJ~���"��E��Ç��]����b\����1I��^�M綵�=?���x^q��l���� `n�,�C��!��[`�A��ݵf����u�g�,%�!�>������̅��X3WX�|U�@07D��&�5sZX��dn�9�6%p1H�79�rF�c� C��@&��̾(�y ���<�i�ږ>¹�O�D(��:�h�c������ӑ��H����v+���/��L�
���ū�,.�����~M��?����-�AJ�ⱳ�g��a��g	���^`$�;6t[�o�V�KE�V�|/�l���A��C
C�)�a��9k��,U'1N��@����3=�Y�V����ɸ�Q�(�@��R\Y^w���Y|��ӏoB��Ǐܿ|��T8��o_w�n�ДD�/���Ş[F��%,=���J3ҍ���~�����#����G����/��-���j���Y��DrƦ��>I{���4��|��k�Rt��iߣ�a����?s�����w��2c��J� D�H��!`�1c�2z)�:����+�]B�A@�Ƶ������]v�}�����;����LI�gLڅ
���������N�� CB�_`!�r͡"X�K����.1�%���7���&�C�ZT']W�l�,t�}�mW/N4���2��i��k"�:50�@e8��s��R|g�A�e��; 	�`@V�?�f���t�HM�ge�YJ;����a�2�������]�6	;`He��<!q����kPȊ��s���=��RYk�������pp?��:��o�i�����2j�����	0M���1�^��a�v�^��L�ڡ ��gsH�um�}P��I�mu.����T��@�P�u��CX�~���k��h2 Ok� =�c;�2b��E)��x�|��K�:0�1�DcZ@7j��{���7�WL���lE�)G
ε�ڬ5 �e`H
�M�$6���X�>)�% �Rm;�����(;�
D�x��O����ul�cn˝�2v�i�:=G`${��Y%}}6d�A�ck�u]��=�R8ڶ�/�c	mU�5	��^����$ g��ƃ
`�e:g� ��Q
�
�QdW�3$�ȶ�πq����L ��$�]@N�N�!��#!����q��nޚ���cե�mI�{��i�y��E�z��*���4����c�a�+����G��9�R�B�,CqD+�<=WL��$�c���Jٰ^�ĕ���?>�E谮�d~�����PAV�Y�bC��C�L	$5-��y�ԉ�ڎ�Д��=���-��4����Άin�l�Y_�6�EnP�~ӫ��1�K�[���_�၄��h;�0_�L]޻VpݏkC�LB������\�e<d����$@��"3 ���ko����,�l�Sl ��m~���o�� �ҙ�I�H�i9�E�j0�}�>�J�H��`��&Nox�s@&|��԰���ꑘ���VH?����������`���������:����3l̹�*��{EN��t�އ�ה�3^lB�wkV� ~����S��N2��Y���?�b}��_좽��f[�ށ�����������5�RJlh�������n݆y��n�{H�\2`H\^��B4���p�v���{�T�GO�q��1eG�������]�"T0���hX-�k�h��-�K�! IS��M �w��_|�z�oh�Q+2����{�xO���ƚ[ZY�F�[P�u6��O�����Ζ~�>޾^�f�I���� EȾ�#�b,�O������+��?�*���ࣇn|��Z@�%� �#�5���M���$}�{Mw�%C}_Y7U5N)�cT��������u���3���������S^�(������6�XɌ-#낼��~�݌צO�z�[
w�p'�J������s������h?��F@gF��x�����O����缯��ӌk��`��Oz�ӝL���B����wb�� �f}T�{3���Hk,���R�
���h��A�.|�|����9�{�P�  K���Uu�)������, [t"�9�v,ݷP [X�Mb�����J�ؾ:�L�V�M<���,�?����cr]�k-�=�5n��<�m�ڢ����w�)6Fk����tk�|E7D��*� �^����Л\C$%��v+�/�̰�'��F���I ��E��ra���N�9��z�j��Y*-c�$6Ja	b�G�8AKL��pm�V�L$$<u6�*`�J����O���@��^?7Ct�ܪ�ee�i�?��`��E�bq�,|̯P��/ 7�(h������6_ �P�U�o�X@��W��Nӥ%�9/>O 	�`2"��9@_g�J��6 �[U���@�=��-ss3׷�x�o�s�fq��[
�h�鮢 ����^�^d̆)]]�b��6`��9��7��u���E �Q� �5�kc� ��є��Zƚ�[�F��O���
�I�F�	�4�=�G0�6n�{�n��I� 4?�k���Z(y�{�����ٲ~�2Y v��>���A׃x����9�u%R&(@��Ǐ9�&5��V���c/��V^)!J�,-K�VY��0S��y��o�əX&��oiy�c�L&T�9�g 0��=���=�KC�����9��N3i�0p'�z���3X���f0�3y�F��������J��7�P��27L�S���9 ����,ke�n����f����b�Z����3���&�{��5�a
8z���E�D�P�;����V�wV�}g��Z_,��2����%,ź7����"2-�33%�:<df����1 ���"{r{X}2.=�8�M��=\��U@�������յ��H�����h!~��{�oA�t���4�me�n��g��O��n�e�x�ܷK�	^��r�a���Xf��3^�wS��{��~�sjp'�ط/:��"�b�T�<=@_� ��z�[T�j�NuȨ��҂{�����v��=s~P��\40����~v��������|�}��}�n\��^���V����U/��F�p��*c�	�c��+���]�Ͽ�GW�ġ"��0:�u�]�u���`����Pn��/��h;���T�����5��Bg�\�[��vz��I`�?c�pGC��(_Xs?���ܸ���o��=����"V
�{M�1a5������8��s�)�H�l��O��>c?^�l!��n�F�[�_vo����������z�J|�At�T`�4��l-]�
6;��Sw�rk���p�Ν����[@�TmPk����}�����)�y�{�ߟT�HL�O}?�~Z����N����6��^*��)V� ����ľ�����SSC�hm �DWU�T8j�;;,І��]E�+вP�(*¾���Ҭ� �l��9c�1�c:�x=�l�E`�q?�u��M��a�`�y�������3�A�Y%�@����YLYV��,>��d�N0">��v�.�D����Ņ%�"3�$<���{����+��1Ƭ8�>t��ߋ���h���q�.��PV'
�!��Ȕ���Z�<�ҡ���(LV�H�E��12�K�'�67LB�@VJ��,K�2�(M*���Ia�8xσ����([�N�P*~>؄��P�4~p��x��!A)H�p�ݼu3�K�A$ �!0��@��p5n�\�6�H�w_Yy`S>{�%�k8༿~�����:��^3Qp?-0���P}��)eƌ�	�մ}�P�e�����,�uV���kg���H�xͲ�ں�e=��1�<�i����� &�z���C�*ea� Y`�.iaĔѣ�Q(X�f)��f6��sOAZz�h��<�z�tyJ���
^5If���`�������4R��c�]���d$Ⱦ���X���Y���wW���R }-f�g �������!����m{�")���躂L��vl�ɿ#8r�M��|��Z�q�y.EO��B���X��b���>n�z�I����ꊳha����n޼��]��>Y����y�S�d�'˺2��;����ۮ����K�Q�	d�ƹ5 CZ2L���!ӏ΋M7�o,�f`+�\*��uq�Z�r��������%���c�qNIY��֩H)le�캔,R���ä�J]��=�oA�G�������z��Ź��<Vֻ�j��^�;SFN��,
H�ZI>�Z&�?��LTB�����+R1Nm]�J%A�;��J&��}v�k{�IO�+������d���<o��=�<v�ɨgC������b�O��'�v	�w0���������i�\�|��ɺW W�괛��Y�k�#20��Z-5P�:,~^c�d%Ƥ=�I��#Y7`,Mߋe�Y����_�W�^`Y�1��xꯝ�}Ɂޖ�<M���8%*�[�gv��$�[]ր�_�z����{�����v�O�CV��<�/���=z��E��|�Ҡ�p�������ܹ!��a(�c2u������W��~����>���<Ec�ڥU��^ZQ�S+��m��*7��O�����p�'�^	�x�i�X�l
������?�A����O�'?��@^lP,��js3%�T����Jʶ({�Ɋ ��+�/���_��_���|���t`q �kW�j/��Yi�}�+�%.��o�����{e�N�-s�Wp4��pB��-���c�@>#c�V��=�������&��Z�־�O�JR�'��p������g�
XH���`z���*e&�J��2�h�G���]G��aGK�p@c��}���$��ā�<�����Oc>�}���j,[�-�7{���=���T��R�?���)2��y*"c9UWF���Zz��NR�������^�j��F��-�� �����t���lE�ȴD��H/d��it�ub?�`�>��}�y�M,����<�U6- ������p�'�p�M�z������-@?�3 ���<��1g�2a�ſ�Z���n�r�K�,�t��6��q�Y �g
8	�V4E���L-QJ��9:SFe�:����c�>�SV>�
��錓}��J�P{��#�4ұ@�=T:���#�]�^ڻ�6��5[W�c ��1�@��:2����wv���KF?^�c�t���I=�b�XQ8c�b�\<�1����|�M!��5�;ZMDF0hYA�:���@�d<I�~~}�/y�G �M�������[r��b��\+� (@N|�Q8��S@��Y�,�@��:`T� ��{ x���\��#� 4?+^�E!���}G�w*�'A6�e&���b�r�H�W�B9���s;�%�d�po��6�W,ܪ�4%��Ty_J0+g�4g���֔�Ȩ�u�3�u j�DG��$�RTҷ�v[�
�bLUZ
�?����M~�@�OY����tMO<��xOi�JI��}Q4i��ZM=�hN�ن���xփE��&h��[��c��&"���ׄ26"�4��������)�%4m*��G����G���8�RudS.�E�h�mK`~8���WX6k�2e��h�:�����ط}�׺�7�yf˂b�O����e�~����x=���l�b3�}kDt0-�!�������&��}K^����p��n�\+���^tO���nt8�Q�P�mzx��m� ���l�n4�.���f��8�~�Ο��~4�*�>x��ݿ�5�W0��N��n��۸�N���������]D�w��i���5*B���p�Mo�#��G����܄;�v6��I��}6�*�,{`�Dgr��ڄ�o������yڏ�U�=~�Oh�
��6ht	��&[�+cS�rd94R	ӊkԡ�����w��Uw9��_�������gt�8�,c��hu��\��]J�����w߉]�C>��gC��;��O�^���@8�ꓮ��˿��ϛ���G�NC�d0��	P���F�����Ў=�X���g���VEV+�f�	��b!1��/�"@�h;����>{�ųI@ �!F�.�b/2LkP'W
?Q^�E% �U�"|�:w4�Ņ�>�e���d���)%��$��#�=V���d��R���#:� ^!@x��\�X�9����~T���Od��4�&�C�cn ��q�16�P�~0␒��� Y�ҷ�Nn9�VW	���_"3���g=��RJ:���C����iO�e��(L���2��@�g�Ù1��:����*�:�}a��HLk�/�@�G���"MR���S�5p���>��@*�l�u&��G
�{e7:�B���ڴ�c��R�.��>k0y�)��V�Ud��He��wm�މ� ���l?��muq'�M*��plϛѼ�[Efg�E��,�#��	�'nRAO ���PJtl�X�c�}���V�~� ���^b��}�a���aV{�9 ���udrF�a�����}�7�W�՞����{�;d�:�{@� 
����}t��5�Y�:oń�>�!`o�J�@N"H�n��b`o���P������Т�}?���3�aU���|����� ��z���T�K;Т�-8;���^�،Ն  d6=���5����]�+��:�e=������g�XV9�$ב�����y�E�O�C&ぽ�t�Q�
s2[��5]tL�n�2��/�s�(ǽʚi!)�)S_9�"�d0f���:nT+���މ��,ۄ�V�1�%�~�O�TjʤSf��A�&۝2w��F�T0X�`���=ς ����WI���(Bk����s����]p����:9��\�#f��a/�Kom��`��y\[S��86��%���}�:6[޲4�_g�P6�h����f�������:ے����$�F�}�0��i>��h�Jju�k��?�23v����Hب�`, �EZ��+n�҂[�����ٓ�����t�&chcE�}��=�tLi���з�˅ ���K+�d%_�~�-�.��v�`���G#�R#�{M�-)�Q��uz�`��̊�w7��)9	iH|r����fL���~H�崹�`Pv�`/�I�߁y娷��;��*��Z������ޓh�n�e���Tp��`,C}����J;��q�cC���vt�v��Zp�������k�ӟ�� ���:�`3���cY7���;�쁒S��m��]0��HP����x9����Wr�k,}��ՓA����~�N��x����3�fܘ�N
[��$C�0�f�}Ȁߣ�$%��}�7/�_"�5R Z���� $�H�SY8½,.-0�Ŋ���|��}� o���B���
(�H�tW+ţ����b��!+{�h�KW�./�Td{3��Rt^�,�᧦-um��XPy��᠓v���\:hl�
�.�P� G�qP@�P�b+�eŕ����43���q��ڏ��XUC��lm'
ʈ��vП�޾����u0_�h�h�Iz�,�~b!׃}��f�#��`C�tl�R�N�ej���w�I��v�݇g �l���_%F���� �}��=22�@�P@6��]+��_&y֓�dK�xo��]���
��F�0xk��s57�"�qa�%��3�I-�Ċ��(4��(P��	x���d�o���e<_^$�熴m=�����e�xa��$�C=_����h �C��`����H%,r,8�Us]� $�G��F��������� 7i
Z��{9��m��B�GI�F�����b�Q:F�[`���!�"�:�A
c��u��eq=U:gY�R��X
���
��c�����G�*u��^R�Z\�w�y���GO�'�˗���3�_����s}�i�<m5�G���3�N����m_�t�<�(l}�Tǚa�\���W�����3��z����FX���B�X�	5��Fׄ%poM��=��������b��2�uǼ���zΑ��+U�G�B��]a�����d�ق'�( ���+=W&,hy�� B��pQ�S�A��ܫ2	Ӛ�9׃k%E�O�+��
q��t��ӂn+�ҍ���"��D�F�1_�h"�Vx+e����O�\�q�f�%�q�H��z�~`�w��S�Ｄ�>���^�>?޻Ӕ��� R�CА@c{�u�=�qd�V�͋Z���E�Co�>�k,OCǉ�n�v,g���N�s�]���u�,h��3?7pW���	}����z�E�gt�H��Lh<w#�N�)` �)3y��
�	#s0�O�Q�֎�j+���!�h�]3e�:"��h�7"a9���LK3��v�½�"~l½�E��!E�`�ly�;nn�������o�_�E4�����B�0���7�\����|�>�� ��X-Hɼy���?�#���������?���R[j�2D���3���[E\��hv��Ր�h�U�dJ�ʬ�YO>G	`N��B����Ƴ��\��.��o��:��,� x$��4�+��@Q6c�ھ`r��G9��0�w�����Hb���|����j���.G��"w��1�L�-`^�
0��A�e]Ԕ��|�0��EY��B������P�uǉ�G@���9:ͦ���y��c^R �0����v�28�	�1�b.q�Zp�r	���[c��] m�籴o�:�Wm�XIQ2IG�>41q�����i�J��Q�����Bt�S���^�߇:��,4|6��/��I(%	�z���
�hu9m���)SW�+��_�]���ti��2Y�(.�e��g�Y�0DP,rZ�$	��y�ǧ�c�"�����Xf ��5x�$=u|<�~l�X�5��<ú��&�y&i��Ty\�����X_'Xc�5�m��}MS/��߼Na�V�ϧ�E�p~ղ�)��9��{�W���M: ��@��� �}�
�Y0Ċ���*Q� ��h��P�����Ĺ��V|-��ꉦ��?�7 ��_+�9�[��Nvv]��	�d��{��cε�\��`�S[ڹ��̵��Y�Ҽ`���He�ԡ��o,R�D u[gRlTt��a��@�h����}�A�d��Y�HD@�����5~��V����5����i>�]����
o�zi�ս�'�\cY���Ǿk�W��n�W"w^�
�0���i��!�T�������;PjA�J��H��X����/1��
Z�XpB�\�� Z3�c�@��->!�>G-c�!؍L����")Ti��k�1�����{'��|�{�b}��é�I�%amO�{	���tMÞd���7}�3����#���:|��2�EdI@R� \��3�/�/~��|��Kq�/�6�F��)��6Q�H!_�g$h���'I���Z�?Id�U�fN_0�����l�_`9�s�Mۺt��{��8i�3F@��μ�����������H��uO����b��\���hEc|�"3m2���c�E)F�q/KEqI�Ma�=r�'ߧ�T$�Vc�������7t��]�X�u�<E�&���ֱ�~I͟x��MH ,�!%ig���Ժ[^�I4�/�~��ww�nF�}��!r$ ��a�LEY
���{�	ϢL�D? ʡ����}����?t��?��{�w�>{���1uފR�%�w5NMKp�yC��6���߬��07�j��?s1v���{�+�|�ݨ��]����, g{G�m;Xv-��_�g�z9���8�j�~'�6�اw�w���N/���k�r�,O��t!�  �e�������(z��b�W��5o��
�
*�^� �Z P
���A$	���
ӌe��@��w{g�υ{�{cKJ�HA���@�x���yf��-i�y����:w&dsj1T"�!�UZ$����-�ex-�3K5�9x��E���QҌ���'�#:٦WM�o"`6�e���j��ɣP8Cq*? l��sdLq �d%[z��
�x^XA�5������� j�#�s�;+�7Ii���R�.���m�" � �Q8Z�HQ�V�!�J�d	�u��:�@���iC���(�=�nQ��ܦ�)9oL�� ��k��j�� �O�����u�-�gA/Ρ�^�㚽��R�G	"�[���bMYh��2�R#IqX��������<֠�Fe�f��	"�1���N�G�%���DVD�Z1gM�g��YJ�$�H�,�,I�T�:d]�`�m<MR&�8Ƹ'ѓ�l�W������h�0uH��<�z�x$��Y`�\2UFDlf���D���<�B]���'�a+�v��5��$�hrr�w���V��23�%�7��J�͔E��G0]~2L���m�mM�w�ⲕ2p'ZpSdq� ��[�ڔV���ι��F)�����&���;�=�g���X �2D�%�E�uk�Sb&�+$�w1�!>�X3 X��M�sm����Ev�φ��4]+��OV/��~�7��9�ϪT��/ <��c�Y:��]5�Z��d[�4����\��>@����
��#�J��7�f�*e��_d�����/�E�h�]�ޓf Z�i�2e��E��Z�2����i�0�l���)!���!�~0�E{��$�\�2��P��̿8E��Z���3��M����|�w���jh����~m`i�HR����sMz�pm�]�_�ZdF��&�'�&]�*s, c�t}�id� U�%$��)���N\�Ns8�w��h]0Ⱥ�"n}2��-w�l=7`
C}0O��!�?���CA��ܟ��5��[?r��Ϳ�O?�����/���OX%}2�

������,�ez@��0:2`���"�����>�����t
a�?~�)�^�U�C�VVG.Xa��dϛhԙU ����2��t�q���� �o%>	\y9l�f��f��S�;����`6~�o���=�>M�T�΄�8)&���{�Ā�	ù�Í��Ϟ�Y l�}��`X�����W�=`�-ٜ
ec��!%,`�ͷ�7Vy_\�n;>L����T��SPxj�n�^
"�Ա������b�UJM'����� �M�rj�V��G��I��H`/�#:��2�{���'8�7�V��vO�d㎤�ޜ'����Bu&qX��A�@m�e�9��,�
�a��E�'|-�4WB�.�/�q*	��_H�fa��E�G@�a��&E0��8ƕ�� \��4d!�Lc9k�S�=$(���r%��C! �Ç	ꠏpx�d�lk�ޅ��6P�E��Ҟu���Ȑ�>LD�φj ��^��;q~���&-]2�+�6�P4��P�VT� ��ix�蠁N�od�ғ�#+4Vg{��������߽�,ї�$��u-v���g��ƶ�����/��`�{G�������.�&�i�blM��u\ )���.Qvb��� �k5�������ei�C�����q5Qv�Q��(��>�1c�9�f�F��B��P#��U�R�}���~���h����s����٧��3��,E:���$�P+��dك���SH0��Ø�Q}�&��f���>������Z��������G���
���xo��X�2�{��8��<�����M��U#^�j�4�տ�h8�kzq~:ac��gh�yQU�cI�Z����
��"/��b�:�;�x�f��ܘ�&g��M	�vW9�V.B��
�5��\v�kϏ�Ճ�5�	&��F�2-�Hlhp��#fd ����'�F�"�FWۙ��������2V5�]
+J0(Ν�L�
��靋�ϵ�Wp�E��J5ܗ܍�7�EI���U~.���>��g�k�[[O<��&���_���2� �ն�M�h�kI��d�j�G�'ƲI��v;��%i=9[��`A���2fI�X��_�^����ez�~�7������as�Z�ߐ���w�}S͋9c�/θ;'l�� e�����>K��`ٷa)?���ͅa\��Țx�ⷪ�`��f��f�7R-.9icP��x`��96��~�n�g䛞��O&��[�̘u/Wza������ʫ�#�w`��2:5k�wK�޹s#:�߸�w�G������mm����k*O�_KK+b�Rpj~q�`tϠv���z��* '8����`��Y� 5 Foj�%֙<��'t�Xh|
�H�q	��y��i�^�|#�?���s]6�?ȷ�9�?��j/ʢM�a�qW!�l���r��;y����_��7����η0�qX�R��ݷm�{�>gƞii�c��%0 �h77 N  .iZ5�.�z�NA��U/u4��QI��#՟,�G6�&hѽ��"A /K�!�#��3�	q\'Z�j���M�UX)e>X3ƥ�Cf�x�>� X+�����z�u:~�Ȑ p�Z+e_��L�m�5��	IwSd�di�H![ �D3y �|�O�4�^3~�
��R�"�@�ʦe���, � �u�� ���HGk���� ����i��/jb� J�ַAǯ��e)��cgg7	�ox����cb}(����2&�i �	x�=�g ��3O�%��R+=���e�ll��$�@�p�U�� XX��q\w`�];S�|���o�o�0k[$�`7�����(�\,
Y-�f,K�zɱK$�	��s-r"�^������yi�,Οw�{{���t}�9�j��vf;9��XI�I�c�'�w hW��/T'��Ŭ��H<��d`hy�*�G��ƅ́��E@R��������7�C���h�<�{��5 q���V��1[�� �n�J���A`l�T0�h����2�T2���ѨeS�snA�Q���= =3%�ܟ�g�� ������r����V�fHHa�9���9���gc������&����F�!��"��d��(�Pk�W�7�����2�N�ض����'p-��7)�lQ̐g\��J��Ḇ �Sھ��h�< `Ax�_��;D%@�ײ8�׀��6�Ƙ9�o��{��)�1I{���=yV����>�X|g&��Q�5�~��d+��̠�����Q͚�5Y���8֐���y�k�o��8�?ޏ�c��_Z|gL�,Jq�.�E���Wr��ڎV��Ry/��'�L���E���WT,�ϖ}t.���o�[��X�5�Z�x��1ق��^������YL �@ewPlB	�x��i�<�����F���@��T&Ǩtm
�U�D��J������]��$�5�͡����%Nk�n	Y�,�c4�����3�Ͻ]��}̀��6wL`�`����9���E���w�y+p����n��S��Ɏ{����ފ������E��'�L�r�[][I�R�y����E=u�
5@M���T�n#�� (}�-��b�Z�B �y��y��rg.�p�|����ų f7����KN c�]fFp����Y�g�2g���h�K�����������P�;��M�� Da�_Zo�g�����V��:fҦUf̨�PƗHH�H[ �a���QV�>��H ��{��V^$:���>�wn�2���������{K��"eQ�f�"�&�!��b��A�(�K�Z��PÅ��Fh�I,nd�6;���o{ZPIܟhJ�Υ�\��;@��S�-�\�3;�u��kٕ4��o�nP��.������[~5�#`PXؕ�$�!�Z���@uI�2tg=	��6�gG�(�Z��(X��B/������5��~���B^�T����gO݃�x]���~�c��)(����N�R�$�[���e��`�XV0���H�C�.�# Δ��]'ׂ��)��9�\�i@�A�����S�<���K�9j��$�D����"1+y��v�@�I�@���c~/��ނh��TR�Y�&	�5Mw�7�+0>� aPK����A
͑-ଐB� �	H�5.��%9�@i���ZF3OWJI�&�Y��j ���Q
�y���f�;hxn�j��uY�)�7I��؏��)��X_��,	��D��q�'���V˾��m��;��0+���٭"`~4�b~�����<����ݖ�b{K��#v�p�M�[��W�~�	�=y��|�g�<�pݴ6�e��l�>D�З`��̪����$C���bnJ �-�*Q�+gw) 稁�[�[���,xa5���-���`�y���*��f�]�?[nǲ&�]��߰�[�L6�v�ѪF�bk��8?E~C�c��✶.,肾�,@z��:�܌��2��j���{�.�kے��[`��!ٛ�X�?!�_�+������M+���t�Yr� D����Ck�����ZIa����HN��-������ݑ#Y��3��ZDC�����>��?�ٟ�g��~ۙ��3�UY)"3�p[�'�;�NdD�U1�p�������7�L`�`,/�f������h@�G�v4o!���
��ls�%�4ϵ���Ʀq�f�-#Ʊ.���kQ6�-c�Y�C����7�����ǫ���f{������<_��X*��i����&8����n=_��;�<��nSN�����猰h�;&؆^��E���ȱ0eB�|y!�l�t9˫�KI��9ܑ7�(��ճ�E��+���~v��������r�\i��=o�F�sR��k��S�n����u��G?���
|�([�S�յ)�Q�޿�7?��M:��Ր/C�i֢�7�=e;��«D��C��@df粳Iоl���)��6o��n0-I��CӤ�7N�����Kp�%/��!º�F����|i���B�a��_��2�d���$$�` 
`V;��\�m�'��Xy�4��,�W��	�L�C�=��H�4l����p6[Y$�Z ,���Kރ���u����#'�X���a�E�}��W��\ %�^�$�X����M0[��P���jlbK��k��F���h�j�7�1�/�j ���<��Pv�p�2�a���8�q�S@�ؽx���4��X��48*YBF����nZH���hJ�C",0l�e��u�Y���|XB@5p3o��ȏ�5����4 ���j������U�agܙ���e���ؼ�!�f)�y��I�����Ӆ��	�F*�6�����`vwo��Js�u�i��ru2	I���`#P�ݙ�l~-�O0����U9��F�`j� �?K��t���G���IE���U3��3ʑjc��?�$uC�cg����l����k�( z|�̟Ɖ9�������P�*F<�`�����`g�/��_�=,����5j2ca���l���E&����}�[7 ڒ��*�0Q����_֪�d��ø��� D�B�nW������d�PIB�n7��6W`�,W��y��L��&:9�紋3��`��J�l�X
C��_ hQ���Cv��*�yʜ\/�Gh{��,Q���y+~v}˯�g�D�����?�$z��__ߓd�+�����	�6l�����Bt��q��q�S�e�� �-��e��l�v����j�-~�:��-�k �E&��9?kd*�5��� i�47CIn�^��v��-����G�<��JaL�Ç��=a꫈�D�C�S�_�b�d����,>�WP~���.�Z:/������̀"�D@��xj���W677�w&�QT��5�jŨ�lC�ǚh�5�f���sUK  ��IDATo�]����P�%m�nR����u�P���M���]s���f��T�I:���g�>��E!�R�]��ŸO��v7׌�Пd�%��Z���vZ^�-��Z���~w]�݌��eA*_ec}�:� ������(�<}�����\f� ��b����;�+�/��C3�5Uo�4�y3�m��9d�$� �A.!y,l^�N��� C]I� �X��'�0��.z�"�� �\����� ����t^�)xg��!I����O�D}GCm�q�oH5� ���~�gN�Ԓ����x, H�4�ljIH1/�"6�v�7c�������;ϗ����*��${d^Z��hi�}�ֳt��Za�ƲhOB�KM"�)@���l���YV���d�A	'�?-Q0_�P4�f��ӧ���(7ӄg����q��̀�D�� ����S��=a(��ȣ�g+������?'�x�O9G��4ɖ���TxWﵫ��i�Hð���>�ߝ�$Lp�Mi����1l鵿7���@(h/X���tFG����kc��mmm�Z�(�&��R�ڵ�  00d1�RKҥ偑l�b1�4��t��p?��T�q�O�� k�3��yͦ �����2t�(ĩ,�_����NC�
PYj���w�(�����Z�����a��D�]������K�
�ʘk�frO`'E�:C�ǐ��'!������\^�\-�H����ܧ��̙_$��]�cO��-�3�g����P�����y	���a&�&���l{0��{>�I\����,��2�o}m��3��N��d�ki�S�rY��Y�w��߸o�sƆ�Zx>}�ٳ}v�JF�%j�?��|r�.�n٤��HRf�����3�,��i��R:�
���)_�I$�=<8d�מ7�g���)܋����y�9')����9m��$��&0�|��!��b�勇���-���Wj���\]���->)�9�,
!(b^M8�1N�g�>{��"/W�R��&��c�
,��P ��v���/]���N�0�l�-��-����h;��l��.U67=���frO�W*}PY�4�vT�'K�����'�#��gE�
�|��r-�w�	L�]˛�K�b���B?p8��|R�xf;�o\'f3!.��RO����r�Ž �(X6�N<fnԔ��0����E�,4e�%.l�]����Y��W�-4y��՗~-ln�⫻�
)�N��R���~��>k
#��������0�D[YB�ЭoH�oڐPc��36"��́�����D�0y{�0�R+]����j�	���"�"	����x &b��� .��\�|+c�� T�,/��4�x������֥ lG���< ���416�8s�5�c�r4F���7�D�7vk�*�Q�ڄc��+4�HmTH?�=��X6` ����IEXsx1��l	��#����S� �X3��"WL;�< 3�pfz}��YJ"e�f=b�`�q�����"�R�����_)s�LӠo��sqq�m/��}M�%�b Ր�L��)�K1�$l�	�3p��@d] _��F����`M�mc�'�u��S��1���V�;����*��8j$�_�w.6#��Uk�x�y��i6�m��<Q�%ȲU��_�y~<��~�9�2���&��?$��z�=k(+ š��di�uuY��ƒ��bp,�͋&��7���ĸ�X�b-Wc�3��$R���hB�0?s��IQ{�XS"��W�����,��3�WO5�_��l���a�$�.�{��C���LC���:�H�
g���`�[2�q$M Ν�FNH�EVD�g�g��q.�-$9i����혭�_��j��1�	Mx>��	�^���ɐׄ����<p��/$d=hY�r{�ya�Q�:G�ߓ�pxr��cN.�Nּ���Ç�瘽�����&��1&�Q?� e��<CwŎw�+�h7��������yF=������ɓ�071����jE8�A�K}CZ�C�&!u�5����������9p�H��q�H"R�#�cu�`��������RFa�i�xdmq�9k��"���{Ø��)8�d�aNC[#��g2��`-ғD��֨���ʸ����p����Bxe����$�"
��O�&XR&kG�s%�5�9�)�B1|'���W=�#�6���{p)�bD���6k��S�+
��a�)G�ծ�(��³O��||���ns�:r���)���:���Q����ۼ����#g���<�q�]�:+X&#]Ԍ��&a�e!I
�����n�����6���,n� Ж	3L����y��$6����&푷�8�ay�v��S����H�.���t��T���t�����;f�&:�0Sbb������c��n��������;K��8��S<7�[�B�l�"*�y���Y��LF�'�1d�^,/1�S�y�{oq��t΍�jcq�:�H��j6�������׷o M�ge�M��<0�Ɠ�l��0q���k �I�`��M�h�
��6� 2�N����e�k0��j�F�h:{���4UK���5Yg�4��� 1�& s
%NXx -n���� 8����c1;�8�]�'A�G6���pʉ�=뀶S>��])���`V`:M�6Qi&�8T���r¼L��:�M�!@��e�@�6�&k��M�UԌa� FV b6���ҝ�� / ��k`�%���{��ၴA[�� `�>}��L;]�N��,:�c��, dH3~N�ܛ�tD� X����kT�!�2 &�Ɉ$�C9�/h3Hr���3�"l�T����0�L�1��~@6��/�笉3u��زgk&�5Q7h�Jā�Q��J-���"^��1�b��U���@ƺ}��}�F;;�� 4@R: ����8�Vhoo��v Zr��)f�\�D'��^��5`'�/@��dbY���ʇCc�����?"g#��m��8AD"}��&���R��1��H$���l���$�ϟ?��?%�FH 0{m	巄�hG �H�WyJS��+��!9��g�]�n-]��#_�e�H1���`�焿"Cg�Y{��NA��C�6C�*����g�cgBS�0^��cw=�_��~�H�C;��ӏ��qź�������8�\/���n�6o�`��n�ֲ%�4��?��u�7�לw��A�̝�܈g�Ğ8�uM���d�R$s�$�窼]�}��B�b<���@/��C�,޽�]&hd:����{6�Y[x,IM�~��G��aZg�s-�ߚ�ޑ�}�6���;;[|���c���� �ϱ�"2���\`������k���A_r+�I����:�ڐ�Su`�:��u��h����{R��m��=����Ujd�����F@����6#��T�=y݇���9�2#/��8�&�:�j�+�'S�'6�.0���a�������v�+����z3*��ཎ��O���.�EY,��:z�����w����"+I��I���g�H�x6���@6� �A�=V=4{D��<<�a�9��e�\{��)@�P�*�X�y��p4�i}'�0ώ�����&�S�g �����.�@Q�m��p�E����+�O��䯫�)��yu��<r��\���w_����zkw�|K�Cʌ��'7`�$���&�k^���>ۗ��bLʂ�d
��B���sR����M?4oy��:l�77י���R�q�D������B�s�	w��Q�WWe��<W���e2��f` @�&ͳ$���T"� `5�0���LdaЈ��y����3z���v�7� sYS���M=���(��u)`i�z��31=Sf˳d�k���f˒ ��e��D����$Nt��\Ds�A}��j2Bf��+@I�8.6a�]�/ѮE�!�y��3hw�_�D�,
� #LR��4��j�DY=Nh6Q���;����De;�[ۻ��4f�I��Ο��[�.���Ax6`}�>i���䄓m��9V�#���dr��f��bI�f�ܖ��Ø � 3��LS$�t�X̃a-�ec��D� ��$�����6V��p�4$}��J���o�~��&'䄆y=Y>%?���x��ۺ
�bPFA�3s�����ʏaLnnl2x�k`>@�66<�GT��>�XX[��H��$���G@h���sD��$� V99`E" ו��C4Y�%!E����[��nO��}6�����\��䘔��tm��ٍ9��(�/G���u�>8�%}�)�Cpv���s�����&��1��Ø @��_r9���b�omF��LUK��6Ĝ� Ɣ����{�yP�ˉČ$���I�6�Ȋ�p�h�A�1iQ�t���o��H �������!K 0��E?2�EY�=�ip�I��3��2�-bm���ɦ�'�jW�J�BԪ�u�D�%*�jbINܨz��/L*�m��d�I6��<�����E<?�:�×�?���^3��㭦�ˋ6��[	����c�<y�D�'cq������R��p|�9)�� �B�M��D�]y.����e6����6v(���A���14r��KJ@0�W��Ԗ?"	���~�Q�}��35ĸ�b=dֺ���͵-o�����#K�Ae�{x�B|�Ҝ	t����f�Ǡsy����"s��-R���S�]h���(h	� �>��*��gQ�T�!������F!do �裶��������nU��-���*��K�T�gV�_<�vEPk+-h�"p��/�|x%�#�L��!� T�\CH46�#R����=}�4��2(�ML���fV�>"8�PV�0� ,����W$k>,���od��v���R}`�%[
�/�H�06�����d��H����윙O�0D4G�P�,����"Rf�0�޿��}����� 6���$C���j\��/��J>�c^�%����v��B<-���E��>֮�d���NtJG���hmK0t9�����A.!�q Z}�`�%6ù���� ��@�3����jԇ}`�����,�Dٻ8�X��@*������4LE��H�`�@8���ɷ����B}�x@�Gǁ]]jG'N�$�������?.��I�1f7cO,m��D�.<���d�~�H��6д��~ g�ev�(��z�N��1ׅ�����H���+�Ƅ��9�yw�-X s�c�6�.4 �f�\�yy�;;܇0%1c6��T�������}s'@Cr:�(IR�ST�-Q_a���|Ʋ�r�@4����
~o�˗/��߲�X{��=g�7�Ս�,��%rq�����1=C}���*[�9�����\3EY�8�~�lMS��%�$��e���mp�6�g�m�f��X���Џ�XC?��A����[��а��-o�jBƼ�y���Lĳ���R�����"(���8�Xg=/ogw����������D]3���n8x��w$��ꫯ�sD]L��c��}�^���I�X���,_�=�ʑ" S���VH~n'N�<D˿�I�>)�B��!uR�-���c��2�ќ�9� >����޽����M �����׷$�"�֫����<��[�h��m�:b|��Oر:�9hOH��#�Uha�\�>�6�2��S�[k��M�A�Wa� �g��T�f���W_o��VU*����x��^�W�\h��j�����b�����\�4���^�y��P���x zӮ��J�R���sn�#��?�,� �x;:
��z8=�ͻ�ȋ4M�+>���Rh����-G�{�,rSMTg�z҄�r �nYx�}<�k� =�a}���&WW=h�Z^=��ʋ[AS(��_�ݤ;���mO��ˎ�����\��2e�����.6�mO ���b@ ���D��Q��Kr�Sb>�fc�whcs���=�M26���]�F
ܭ0C�����&<''
ֱo#)؄�����5���z��$dbD���9*f١qm0⶷��.&�K(z�.��	!~ &��2XkoI�2�:
�`s,�������,�� f����/�I���	��ə���@�h���B������K�����&��g7��H2,�>�UK�����R�f	�Q8T�? �NC�O*�a��E=L�e)ڢS��V<'I)���¸PjZ҅.���t�'IC�!�,̽�����$&��]������y	�@Q��x!A ���������2cS���)˰� �3����.�k78�c+���"��S��X��Xj�����\t���h��GK���A ��~GB?Mv)KԌ��L �0vp,���l�ѓ�XW�0�K��	;[V��o���F0��ovz��i������̴��<S�1�(��,) V7�QC��g�c����B�B�>����A>/^�5F�??�%�+<�����2�q[1ù"��A�݀�v8��7���F\� ����93SQ�S\����|�ĸ��V���T%�V���&/�q��K����J����A�i�Ac���F9BVA��2��w����܇��d�NS�8����si4��+��u�c1�P�X-�������F��U���	5e�#sט���;P���x�y��z�K�,I�$h�C�	JѤ�PNĪ���#��8sb��� ���y�Եg� ���s������(/`z���3�P�$S6��'��)=��=��Afm��rTć���жƜ/�������ܰ�'! ���[��h4RM��Y����jIX�t���	?��I���X����)�������is���v�3�2p�#j�q���tO��bl�;f�Riq<�D2��d�H����������T�,�]���>����Yvt?��߹���ʝ�UΨ.����PQ�P�O3��?�8�?k\.ʋ�B��36t�U7x�Ib�y�\Ƶ#��mFw[�ʀ���1��僧3]�%�3��*|����9�z�A�k~N������_y�2�^կ�<30ݿ\[��o�Y��e-8b�?ѤQ�lsů�3�@ ��o��ut�2*&!�`]��F�B��3�  ��Z!�XX`2��~^�w��"�i� 2o�/�ʰ!�\- H3����xcIlJ�w|�lq�4�zƩ0��NL�U&��M�S�`56���<�w̖2�.Q`Tn2�9��8�0�}0��r D	x5Vd n���@�["�	N���uaA����ȐD�aӉl���^�E)���
`�@Vl��ct^�˔!��Ɯߟ��3:�_��k�o�ڦ�थ	��H�e��Dߑ�Yc=O����*3� �@����I�r�����;��Q��]��u#0�p�&o�$���x�|a%�ԃ�M�y��|K��z�
\2`���}�?���<K��ܖH�����,�9��Ϝ����t����BK�ט�Nf�C���O����bև��o�3����G:=;�>�RN�P�2�'I���������Lס0:��Mڮ�3ج(��IYyu�˰ȁ�9�d-�C�*��B��X��	[sB�I�ƓqH�h^[/�<�{%��-�sU��ӆ�y2\4a�bQ'�"IҐ�,��4�"&,�b�� �c����5�o��0H��?��� �m�3I~Ȳ�?�D�ü�R�d"�����B��d�c�^�n%��D�	dω�1�bNh61�i}���8��x����p�ل�H�ǠDBhrB���yp�=y�IӲμ$%l��nN>�����^ЋN4
���7I�>���_0���=�`��>A:<7+���yc�
��'N�g�6�\��'������o��r���WRrα���n���rt����`�8a-�&vP̛0�7����GD"ge7�����F������H�+R )��|�Zc,n��e,$�6���Q�������}Cm7�Z�S[��+y�?��\&�d��,R�-L`�,�Y,>���s�Ϣ#.6kD��s欓���x�6�x\f�?�<��)i>�3h�D���>�4�����Y�`�I��g~1s�� 	e��ے.�'ʲ�Kh�m%�-Z��rcVZ��Ԙy��?'k����V��y77/'�R����_7Z�Kg ��3�R��~f&l����k�y]�sm����}_7�|��Ɇ]-n����6l�1B���P��c�!\�͌7b�� Ƅ%1L`;��a��s9�[�ш,�B�1�vW�D��Iذ�/Y" �H�d��Q �`f@�T��˄���)^�j6o���7_M���޿�ɅXے��c�Ǽ�`eg'gr!�ؚ`+c�lɛ8�w  <�A�#��s�'征��+��R ,5a��A�'ɟ�����$ `hC����v4ַ�F���s�~�Yx�s�v�n�Ͳ(x2�ɚE�
�5�������ض�5��T��� ���� x���S'����f�ׄ�+�
�L#�i2���k��'�'Zi
I'�p[�D�nÑ�,H0�ڢ
@����O���r�̀�D�F�J�� c�4N3I��v/X�S���ҤkU'��a��i��+��hnw(�g�g��&m�'���@��g�ς��5�}���%Lt��1n�&ER6� �
����$ �����g봶�΍d [��\�>����C�y]%��$�g�b野�k�A��ָ��"��ܨ�WN�;��X�9�p�0�ߖ9�e8�+��Y�h�DDB����Fɭ���/�U�,B�,���lI��-ܙv�i�©Ⱦ$G�E0�Q��		ǡ;���b�FuN�Tu��ع���5�{Ay�ĀC��������������z�[�9yS�3�u�  wʠ����f`S��~��ߎ��-�S� �H��n��a�sWZ�"`�����\�܂9Դ�)��
�$5]deK[_����;�`�|y��Ы:��k@$� �����K�4�o��8��H�_H��u�MA�Y��IAwv��u���{z�旼m5f&�&m������w Ɯ9�2u5U��R"3��� �T=���q�a�"i���4Yiks;$����>��ko��"a�%b��H���Fτ��8��3���q�u�O���X�5�|�V��Z�\c��K�{Ʀ�̒�e�~��Xa����oK��^e,�I�&���$41�3�뢓&��DI� H�Q��-�v(^����-���\&+M$V�bn�@��&gH�5Ƹn����'��4:������ #/�	{���`x�8Rɤ]�~��:!��\y���O4��߀�V����8�A-�1ߜ��U��c�Xkwp�;2�	K�[c���^�y�[x�0��~�ˀ6r뛚�H6� Z�wCe�v��vf��䢄͸� �y9�(�V�$uӐb�eI�
��zl\9�\KXNH���	�!߇1m�7��T0�Ę�r� ��_��\�[S��H �9�k�B��|&`�X�ƚ�p������Q��I�`�"�*���V����f1�]\�,��F���	����|��E�����&px�^�b���϶2�E�8�S-�c�ϰŀ-��]g0��м����P�ݝ]*K��&�!!c,M$$�����n֯e�h^�V���h�sf�����Z;�'����"�\� ��v��	�X��Q�>�:,K9� %�Ȇ�!U���2����/�u<?���,`ZZ$�	�Y�W�1�����F�@��  �߿ItWWx�`ܠ�ۘ����(�Z$@+R��!��nnl1�.�i�6夡�5^�z�Z̸Ξ��T��3�%�I�fӾ�
P�s.ba�# ��Jb���>yJ[�[|?����$I�����R�����/��Q�%�>��uRf5��3K��O��A_y�ٸIDC��O�͒h7D�t5�@@<3N&����H2��ࢷj�#���RE���Ɨ�NIѾy��
K������u\�oH����7K�4���s�)��X��Q�����5�"9�:��+�mn�F���$�7�ŻF�9�x�С-|T�]��J[��,�i�e;��������]�]MB9�t���u�������j����@��"�P��'��2�mI9�&��M��t)����Q['08���]��w�c�T��N��"09�͎+8x ��i�km��������D�7'�9��}\�Y~��4+�9�Y���-���L|��
g�W
�w�O~6��颟g,��i���Y	�gzΙ�A�yZvT�
o\Q'dl��L��	J�����d�8�,7ɨ�UZs-4�/h�!$:���/s�4f� � ��5��>�+H�Ѱ�3�?����Tʋd�T��U��˙H؆�I��l��赾��'�\�s��\�؞���o� U�+ۋ��S�O}�6�=DW}7�H�4w���P���*, p��1������{r|Tʀ )�� ��v� Ǉ��|���3lַ�\�\>víCNq��-f`��(k&�fv��!h�H�-h8Z�.6�8��~�^�D~Mh�p��,�6� �֌	�P���uAmCp���%�-bdE.�ryŻ]��Uޜ3[,�l�7�f�ښ z���Tՙ�������3I����PF��m	 ��'˛�!뀆p��kr���j�
`�����{�NKb'���K�rE�S�'2,�sDy�+o_�ц��g9�1�b�^�={�ರ�[�d���l$�C;�5
p�ٵ(#IT.�Ì��	!z� $�͈������s<;?������kB7����.��bN�ݸ$��Oq��IJo����յJU߹�w��I:�(B�7���ZY�0{�I���mY�
�k�6 R�������2��	�q���D�6$Kfܐ��!t��B�5�pP-m!Bd��'��`nü-G;Xʑ��Ϟ��s0ߴu't�1�{�vK����tWѼ꣍��Г�ڬw��������A��]�8 �f���M,��<+%+��m�K=	NV�+4�W�$vט̻���|H��<&�'�~�9�g��s[�+�K�*���@q_���jO��-��l��m��������Tf!W����)�@R�ymZ�[������ı ����9�Q������]�!]O�T⨁6�����~���F�xN�Ϣo�v����,�j����M|�I XL&��z3�&���W���n���(+��п͙�W׌�9_?z��b��ԗ���X�]�F�W|���e'�H+�nb�כ��t�w�3p�ϩ[���2a8�0:�h�y��9������g'g̐�$�=�h��.���0��r�g�S>�Jkn�.������.�WT��Y�Ih�}u�;}�Z��x����a�"�M�se��1 �Y_�ơm�D�8Y���mZoT���Bux|MS[dƞ�����7�jL�6O��g��0�(�ne|��ٓ|�Ubn!�*�ƭ>�h����<�pҟ=eA7e~�@`[0#f��/�E�9�0(9!��������9,۩,��)U>�7�ц���{LU�����l6�|� �U`��&��3�i:Y 
��, �t�Β�IM�I�v��~n�F�I���k,���{ ��U�Y$%	�*��{l�a����F	)b¬D���8X� � ��R6 N�u�uR݌�:l޻*����i���do����1d��>�z@G�Aɦh�:2 ,Q���n�fo�q�6�hq`�\��j ����3(�a�9�g?���~��
��iw��u!/�x���`���i���^��ʒ�u��Up٘�R�kYF���d覎ɨ<�>�?K*��j�3�����t`;��8ʮ�;�������1�<�WY���Vy!�ԙ>�b�L1�̮آu���U�S�	�*pe盓:O���~lz���Q��Pr�&�R�MWDT/@��OR��3�8���s�$�;ԡ���X��~�*eA�:����t���S�|�_����]�{��V��̆�IvaֈN���REB<>6�g��O�pS�d�k1�h��o��|%���L����XV��L�-�ʋ� �I3�$>G�ϊ�Y�,��qs�rt�`����l�A�f����������X�H��@6���Pĕ����!ko?�DN���&C�������!zCZ�X���kju��@��e/f1�"ԭ�V�_�a�m�?�� ��3���Ʋ�L��9����/8�-s�C��~�y�O����x�c��f���rr�1m���1�E?ܗ��s��`'�f:9a�#�����~�~�{"�����w��(f����<����������1L7�i7bЅy5�{u��'.��Q,m<����̴>qU��6����h�r��$��I�$ٖa��Ht|�R��4MfTܣ�[k�T�6~�N�q�{x�G�1�H�*��|	�6�j�ٹAz����/��m6��&%'�J$��-�EJX�3��T��e��Yv��� �00W,���`2�7AT��c� ��^Ɠ2óJ���$NF�����ݜ�I�{ԧ�E�@�̕��b��r���\�ڳߺ����zѼuE�����g:ɍ�dC����(�ۚdYKd�}�G�P��G��r��h��]q��&�;*�Y����4�M�$���H���1��Ԇֱ�f��s�?�t}��ǩ7#-j����e�X-�~��E;��')��t=U�4�B�����9�ؙ����׬�`�:h5�')�75vd񢗭��*�^���v�e�x�k��x.\�B�Uƅ+"d�CcM���)n��Ŀj���1��^�� �����i֕3�e���գ��Ә7�N�1�Wk�(`!s@�kޢ�Eֶ~�W4`�~�g.�1��E��m{*��\`��b�{��'R����2��J$������hB���������t��X����6��L$D�D+�[���7�p�����/����^Z�*%�&��/o>p����)�P�W_����5[�?��tLc���0�=	!c�&W������
ݩ؞O<�j�h�N��T ߞ�#F���nԵ��:���_�5������/̉�	�t����	r8~&lD{W0A�0�:]�^e6^�Բ>�Wp��r%Y�ɻ���n��z�@�]�q��[��B}K�L�m2u0��| ��`Dn�]��h2������=�`a-�"��709_�C��<" ��u�~󱈷�D�L�uۆڴ����L��H��=��ge1���o����I��+��B��O����{En���,.�E��j�"f��v��l�(P�jU*����;����J@�5.X?�}N�i��0�1��4\���6" �-�3gz���B�B_�~�U�N"� ֐�sv��?��Y�Ӊ潈_������;U}�d�9˒ \�V��(�l��)��wr)�����'X�D����wƬ�m��f�:/��*+����,\RU�N����m��j&SyF}?��Tq�!J�"�x��+M
��l�����UGޕ�\��Z���j�g�-�~���7	2U��@���;4���|��X�ˀ�ٟ�1���%3rK��p��tVΜ�8y�V�Q�\is:
*+s�\���2�rW�t�a��41���5k1�'g��wzrF�'�ttxL� ��K٧A��,e�~�%��o�q���˿Ћ/x!������?���=�R�g�y�G��h=8����'\���3j��:�$M���x�t�/ک`�ۢ�:�M9�F�����=�c�|�[M��P��:���$XY���}`�l����trr�ڴHltzv&��^�J���L�i���5[��4	�7679�5gsG�mR 	N�΋���/$�Nn&�b/�ǜ�|S�Dk;W�o=f�7l�=��؂�^<K�q2����M"Aps��-obzx�|Tld}�o�:��MW8,�u�,UΠEf��iz]�`���\3@�p���.bN�R�����_U����op27�����Ps��z���c��^Y���]�k����~�Hh��ej+���3�%>L
&��2ב�*�ڜ	w��lӺ�f�n�&�"Ds`�Y6��4������5񼲪c�8NuÞꎀ��	����*�A�eG����{]�>�m��V[mK[��~4����9La�j���s9���p*�OpɊ5{��61^3�>&� K�����∓�����w�m�a��h`T���d �����n��c�oHG���{�״�]OK<M5�X���L��倎O��:xBGǜ�i4�β ��V��V7�鳧���+z��5���Sڀ��3�#!N��b�&g����`D�i��
'��4�����zw�Rצ�}G����V �\�u^ﱧ���ߚ6E&�/�	��QXʚ�)L�]
e��Q4}9k#���zD ɜs�zǋm:f�cj�(�Ƴ#���x����e]N�OX��08���vʿ*Cb`<�,̈þ��������g��pAB$�A�y���FV]���{�J�zgX%�\�B����2�o���c옲�2\Sp�G�ˡ�W��V ZT�0~!����ڢ��j��b����+��-<���$?����Uɓҗ�����A���un�U���a.��nU�;xT>�'��
ڴP�L�vOn1f�j��4�1?�>o_�
�k��S�UD�;���w�d��.s��X��R2=�u^E�b��*��
�<�Zz�=%�f�0?ͼx?v��ǚ�&�``B춌B�Yʗ����5��x�)���r���,��D�=��l��E����vV�W�S}��k��7�W|�cm��j�|L�Ǿ�����JǇ-��Oc���"9:��rJR���˻�֯F���b^
����I�<�,�9��V6�myW����-g��}�r�,��_7@"�~U�δ��P�&�F��%���E��	s�:=���s:�x@���_��a<���X��mq��gO^�W�����;z��k����67�����/�3�����r&��z��'�nv�fB+���N(u�Ǵ���������z�G����/��k�h��J~��q��юC>!Ȝ4�h�y-��&� �����p�B��:�7�\�6�i3P���&������j�,aU�I̺;��ˇ���_~�>��>g��������.�ȶ���]~ar��Gp��_����������|��{B_��?�Z�7	��ˋ�K$�t��zD�k�{��\э��}�f/��
[�� ��/-�	���9�g���2� ������71@�L�Ų�?)5󝆷i?����kVm���z��$"6Ϩ@�Nc�̻;�{Zf��~�_3�FE�#?��U6x���-{��c����b��}�֮��3'�{Z��|2�-�o���+,�4�nz�g��W�e)s���:<������e��\�	����|Րhu��۶��~�������`�k�j�}��Z�Rr^� �^�O�2W_�m����;�Q�em�}&f��,�� �w���� �f$H� ���lrGLrL�z�����[a��o��(��&+g^yIX��G�iί�QYA�X�X
�l���%-�'^6+;e��Er;����L��`��D4\9��-; ̐�@(? ���������<;�d��X7��/^��o���^�xEk��@<;=���-z��y������{������!�������%��ߖl@Z��BH)4M���_���E�V��f�e1N�uW�f�6��t&&N��̛=�MpM�Ie1$y�̶W����l��.C��L����=��=�� �?~���>|��8f &���0�}���<e��B3ҳ�䘋l�W��������ce���ӿ��_�������g,��F�!��T���C�6?��_`�bn�@��w� �yE�ȃ~����-��)���䥢������̼v��k�qN������NL������;Ws��I0��q�W���G./m׼��A!{�lQ)�[�]��+����]��uq��wi�1��r�Фڟo�,W���	yV��e)s�v�����z-�� ��Nrn�QD���];@n{������W���e�[��������j��(��̫�$e�.r��Ԙ#�r, ��2&��=,Iz�h2y_p'�Ў�,��K9�tOj��JIHK�������|�K�[�8�j�o7}?�<��)8L�@�Č�O�����e�z]G�r��ՠҙ�Xh��Ki2�p1L9���8���C �G���~<�㓏��-j�+�i	 ���K���G���7����r�wFH����S���Ǡ��J���`\c}�&��d�:��I�&uV�j7�n:�.����Hۻ-J�>��������(/�ǀ��DQch-��ʸm�����^�9m, 0�Ӓ�p4G8�7lq�S������U�Jxp������
'���g��A��?��o��_�߻df���Oi��3��ۣV�?!1�j��{e-ܓݲ��i6����v4sB�f�E�߿��ل� BRfss�ˆ�8��Jn�!��%ފ-��ag�I1�d6�
;�i(S���LS�s��*�Y��9����3��a��?���Y�re �_��5��C?����i>��孯����9_w���� �R�r鐇)7�����ly���{K�������%������{�=�����Ye�q�qwgW?�꾇x�˷oX�\W���'�g���{�ܦ�ϭEj��˴x���E�Q����Ę��8JL���.@c�o�6�G�^�W����x~2����L���Y�E䍈;�ʊo��y�Y+?�=(c�`�y*�?_�y�G{�&�.�?�g"�N�d2bؿ�ѐ./.�X�����1�?�����)5��4�h}u�~�����_MO�>�f���W�Vi<F"�	��hoo���m�v�Oz�����/���[:88b�e��g� s��B++]�8���Ih#/��H��i����������?џ����?���������5;���� ҌI���٫��G�/��z���t&
|�sK�6��i�V��*s=xl��k��m����<zD�,NCr|�ן~��~�W��矩�Y���^��~�-={�����X��i#�Y+�� �"{$�$d�M!��J�����~��W���?�����~�-G���o��C�"�P�wZ�8�AzKvj�����T�E������g8
 nѢ��=�M�[��y��xvO�y׸���S�ț\�q����-��v���9��Uv��s�����[]�Am�{������9�K���c�n6v���j�c3Ɋ������ύ�� tAFS0��f��33��90���C�/� I+�K��ǈK�v����噟z
`�R��z�Y'�9�'�g^w�@�)���7� 8����, ��H$;�x���./E���v��Y��O�3����_qb�~��Lˬ�$��A���/N����O�����	���?�$}����V�%, �J�Kd�n�h�2�n�Ckk�4^�u:g��V�IF_�-���@>9���zy�I+c��$�PH�2oQl�ހ�=*_���{1h'�g���\�|�IQ���8��Û��_]s�_�k�/տ���svv���������u�^�z��2+++�'�q����`t��З��ш�W6M�٫�����������88<`�2^��h4ҙ5����>�����<&�D���V��I����]�]�<jI\��[�^|�i.Ӗ�HP�>A�>�}�;���ѡ�w0O>�{��9ms��sr�_wW������3���?v{�5�����6���n���Vۃ�a��K\L��4�l��H��BB��z.���� s�&U�y)S�H����}1���|T�f%pmaOJ1����#�A�y4{7`��(�	�&�Q�:��C:;;��c:99���S:==�� P�%)��wT�����/@2���v���������>|xϬ��xH������nu����F
i�65���&��v�$�V�X�����!����9�����O/����/���zF��˻�y�\ �~��^0k!�7nH_L2�a�n6�3�'d: K�����V{0Qz�$&irm\��������wvm��3�<����1M�ǎ�1��?������,}��wH\�]>>����� ��� <��@�	�}�GB?؜�2�������$��D�W2����ˠ��o��>p͠ጱ�p�$�|��k�Xb��>�y�Ep	0�o99a�4�uݵ�l�=c��:�E��@�C����n,p���a\�b�u1�Q/q�&�}�r@s��
�'��V/����������J�
����j��4���BNԩ>I�d|!_��V�\�7E�ۥ!B���1��K2W�9v������D$\�E��5%'��D	��׵}�aQ{8`�d����`f@c׮�\�oӪ����>��`�qiy|xi�PA_�%<��[0!�$��G�Gg����w>�A�h2j2�xc}�����o���v�w����4�j5�Ի��p���Q�wN�;;�`�/闟a��_��=ױ��N�k4���^P�9�0��x���v�DnwZ������z��G�8��͛���M{����O���o~�&���H�F^Θ>i:mÀ�(<��Re���0C�dԂPXդ�9�'S�s6͌|�9��`�3��ҵ�azzxD?��#}�����������?��?�&Q��h5��H�|������e, ����W�dA_`���;�� 萏o6;�d����#�)���o�����_�V^8zPW���dq7y�v��ʱ'��I�EFf���G��� t/{������Hn拃 6L�d�	5[MZ]]�ռ}:�'}��� ��V�� tm��ݓ͙�\}E�1A���G�%=����=�$�Vu8����9��I��jwc��S�^����j{��A�����j��K3!�e�r�,�X��ݒ YQ�-��h�2Έ��� #	�\�#���$����Bj��o<[ۗg�X��-N2įb6��VC`��"��(����"��ձ`-��f���䙭|zv�`��)X˗�h/��qj���:=�ۧW�^�����%�S �p�3�6X�� lQ��Z����i4f�y~���u:mڠ�p:MZ��3��		���g;��d���E��4N��is�E_��]�яo~�l"�yh�4k�X��3���o��k�R��VP�=f�YK����X���*�+���q���E���Dy��U��O蓳F�2^y̱�U�"�����/ˉ�p0��wyѧ&X��ftU�}�x� �������|�����t]__+���B�U�J\��F��?�u�1�} ����5	��6�T�_3x����e�[(��y�_��0�www���e@�!5�q���s̚$HLE2�p�H�&�/�g�+<�q"���v�%a]3�ʚ���~
V�]�����������{������j����j�틵!M��9f 3I(��p��lI������SxX MbY�2r���B��	|a��<u�]�M�u���i<��)~Z{x`Y�;%e���+�	!/�+o��e^]?��L(�Q���� �A>@��������4i0��/^���M&'�;??g`�����6ֻ��tI��w�7���C�|�����q4f��]c`��b�Y]�� �K����p�����H���5�do�ק�u�{4������Ni�����2���5����E����(�^H�gͦ���7��ۢ����p@G�G�׿���da��ݷ���ÀgИ�U���z�Kv����-�p��e���8议�J��sH��)��40�I��yH�y��傥g�i������N�q�U��^PN:��<��K=܇�v��W6�H�����ى�m�Ϋ�cv.�}I<��O ����pD�р6.6�}����2t݇)+4�ê���8����H��zN�k��l�G�[ͦfN�/���d&W��Ů>�MMA�W�w͂C1��>�";Mm��V[m��V[m�Є��Xz���lI�o�\���� �����$U����,���2�@��O\�]�%��UV��ܚ�c��������([�W���X��4fV@�s���6�J��
\��f���Y)WW��������@L̋�>���%�^  x��I�O�9�����Ɨg���f֠T�E������+�;5�ŋ����^ѫ�;��O?1�n�P��B�q��O$>��9cuu�666��x���Z�Mp���Jǧ�����~��~�����5�Г�MZ[ݥ�_���o�����5����	�0{g��S��1�1D�]�ŀZ H��.;��3��@>{[,i�U�?636�+U���>r?���c�2$b�g ����*1 �M�Q�>�n5�)��e
�uD�I//k�q�:1)�E�ȓ11����)���?����N�׷o���+ꮮ��>C�/�ӷ�k�ž
Z�|�EYh��H�PmS�4�I�2~�����I�+M&ó�j�x�B��v�C�k��~[�t�H���yPq�y�� ��� �߻���l4ya�����;�3i��i7�����7�ɑ��˚jy���Y��n��j����j����>�9��y
éXydŉ�S$��d	D��I �Q�BwYc\-���4�q�#⥻�:oe}'f�%�im��b�{l�X�rt#\� \����y}G��#�
�(z�3.4�~pF�ᐙ��G�trrN����P$�J��h���.3��{���[��o����K0Q&���?P�7ʿۤׯ���}�����@�?����I��5��#Ip��l���G�l���.��߾���iON2PN�NO���|D;�)m�m�w�~MGt|rFM�RfG#q ?�8T�Z����~����|1��9qx��?n��f!M��l�:s�����ޢ��1���=<:d��Y�={ʎ�ӳg8$�'Jh���Y^��:�Uҿ��VK@��Ly�s� ���!ӥ����Û����t�����G����"�B�*7��a�C�uH���v{F;��E�豅FfR4�;����\�-^��ݽ�&˸� ���<o\���9���
�yg�) ���Sv����,/�Y�rq�-j� ��`���Oj���Y�����j����j����~[&����Oc�p�y�.ɀ�LW�4�W,�t�X�����̺/fR���9�:3��O+�����l��>����1�<�� ��n���GQ�7��-����kqHB~]$��Ǐ�]���[8��l����sf+L;���A�'O��4�a�$ڥo߾�����V�K��^���mnnQ���B����u�$f1�!�@6�{u���>�/^����/�����j7�i}�)M�8�:�:���џ��o|�N>�%���F��!K`diR賒�ʘa;{�4d�=�����@O����s���t�Y�����	���3^__������qs��5��@�GN�Q�e��HUx�8�P����������^<M�k����&�O�+V���#�U��1���c�..��k?�W��
�`aP�>q��5�1��� ԣ-����������	��>����7>_Y�(Ky��?�|�8�Ü�,gg�[I���{\w$D= &��tY�5�!�ݍ��m^�/@���j����j����j�����!K_�WJ��L${] ��{h,f�Y���c�dr9�ȴ���le�손cBf��۰���X:y`m���|{��ƶS�M�a�2Ï�~/�����8�F��p|�	�NO.h<�'�1��<D�Z��mѓ'{�Czyqκ�8���<� <��tZ�� V6���}x�6�.�v'������O���p������p��18a���?����C���+��Qs{'?7�3���M�JO�3���\�n���uZ::8���j��4TC���YLE�������
��I���J,�yO�E�e��^�]9����G��GSU.�����;'���xُW���6���2��\��={���]��d�x1�9�b��0 S�!�,1��agHޗ ���Cc��I����C��r��F�T��x���0���M'Ǉtx�#V����f��\�)��ǽmT�G�̫S$���gg�tzz�m��=��1�LkK iO�D�m���}�Cf^?y���>y�N+�{��m�6��@dD//����:�h�F3�{'tq�q�B�6U����H#"DGle�O�"��j4�s���ڑ}W6�����b�(-hn�V/y��r�cQU�����qܓ�[�3��>���l����}�g�����(��-���&��1?�/������8b�ވ;��t�y\6#��l��Y`.g!�{��~�E�,����"Ef�gRHg�A�Z��J�P�۴kE:3|�ئ�ߺqW&!���ϣ �Mx|X��;��y�P�e�������&�*�7Y9:-�`�P�D�ɘz�>���S�G㡀� �}��iwY�Le�{zz�:������2��n7���0���4)�F]������=�����1�dY�4E��FM\JϞ>�F��,���m�.�z�{�d\Mz�j���]:<Z�:7�)��y�G_���6Z��١05�m���j5��l,�H0iSD�\G ������A��2j?�̋�.g�o��)Jd����I�T�rD#����O7��-A�uG-��1G,�r|r� (d\v�w`�ހl�x��oؠ?`��h�f��R0���O���|~ΐ��߃A��f�k��#}!7�L��˔��"#�����ȸ<�`��.S/:����38�c�k���$ ����2v��K��V^��P5�Q���
�쬭���E����A� ��M��4����n��$��|3a�8�7c'W�ݦ��s�` �q-��(<�`9�S���r�#qDs�j^�G���IK�Q8+�8���o\�ǵ\�6��I�V[m�Z=r�׾���T��ނ7��Z[m�YA�Qr�c��4�$�Kx�9Ϙ�Gس�a1'A#ӈV&>�Ŝd�d	Ke8�Fb�ζG3&3Q����j��7��?gJn����R���8���ˮ`4V�%�&���g��o��� �qjV���=�-�`E,3򲄑z�����Mɺ5:���U�n�t���=�tf6�nT�d���������;%�(��3��ht�c��`����z�`]�����^2�����hkk#?�����x�>~�H�[\�+�,���t@��6�o��C����~~�Ui�ЦE� �g����)gV؅S�|�vSr_*_���35$���'�?�@S�!Lǉ[	/F�w!%p�����"Eq~q��cOg�8���~�����ӳ��ێvKY�B4��VWy\��,��7`�~���l(L�f���Z�`ى����X�
�$� �;++*m!� ���*;Ðm�I�4Q( x�q���4�f���n�^�x�'��ˆ4��F�|�I� �M�#��Z�������C�ў(ǩ�z���^��j����j����j����3��,Zf�#��4c�� �^r�`�V��sU�6q|�\�>��k{,Gd�����v䈞_tjXgN��]�To^'c���`X:��3A�kF��k��D��p� �x����=K�'��X���M���K��<��R�%�]]���6�c8BR�>KZ�-����th�$� ��p��Vk��������6�Y�ڭ&{��c�	�&�u�[MG�;[45)�4�>;K�پ���  �ˋ�����1�E
C渳� �ۘ�=r��Vu[T~�7_���0X��Z����,�I����	���=��Y&/?DH�O��p>$bX�a0`�- V��T^r?�ƀh0'/��J��?����D"H����,c������vm� \�v9��2��N�b��`�r',m$�{�gp8a\p?�7o�Ԏ��zmu���78�^����YG�d������r�ty�t�;��DWt�,��> �����Ю��h(cY��Z��,��t�K��j����j�����&��
q��߀	E���Ś�9m$9� �G�>����ز�jL������|�����Y�p6��f�c�o��M��s�\FTf��~���
�I�����m�0Ck{8[�5�p��+ K����#޲����1�ـ˙���a9�k(�6_!����|l~T�5��<��X��| 7������{{P3�0 ����W��.Y�}�P��I��8�|8r4>]X ˭�|���`��t��F�������m���IА=99���3�3�� ���?��?��j���(�9ʏH�M�kk\'0{�}fG��ɬV-�G0�����bF���7����G�u��,AeW<o��?羂���1�ّ2��
���������I���h� ���K��D@k(���o2�2[ۛ�dR��M�t�#�Hƙ�c��C�C�f6'��\�9� �N�<o8d���.�B��E�,�^���(�KcvA��������狃;��/��n��f?�Y>/l�j���]���|��`n��m~�Z˓�(�N�? z]f�|�A8���@Ԅ%K�b�v;�4�TC�=�E-����S~�wY,�V[m��V[m�-f� a���TZ��ˮ/�b|{3���=����_�\0� ��g�M��ݔ��Q�wiB�r�h^/���	X̎I� �d��;qr<k1G,fˡ5K�x�0�v��cfW��-j{�)���5���/�$�L�6+����V�M��E|E����8�AgRN�8dR�a)-�<�hi��wZ�+�elʄM	_�Y<���F���2����r�/�ۦ��U��=��R70�q- k ����$���1��/?��?�Q&�L:�I(}��yvzB�(h�������}���Ӛ硊�-PΊ�2��9�/���Φ=]kK��~{�p (��6�N��l}
˳�xLA����З�U�%�ʲ�Ƙ���/I9W���؀��fkp/�����3����}H� �Q	X����'�Dt ꔪ.���)5?BK�2����4J�qvN�⧧gtzy��[�����=9>	����OF�j�XCz�i:��噑�$���h���s8v��<���p���Q	s�Bkk�q?�z�����E���j����j���;2?cAW/��|3�p��Ú؄I�e�d
��ܗ���e:.�-c�b/�g�=!��"G��Q��h|��1�9џ2�%�_�����,���U+�!���Xm��u,����ʝ�)��8v!ٚ��Fg�.\��1�lH]�e[A���ʱ(;$����\���7,��pb�*MF ;���n��<8&���"g���q聋4o|k����!� κ�-�d`���d[��n�P�O�`��y~~I��=�`�VM%������s~���p�|�%:ϐ��_����r�~F7�4qh��gQ9���b3�ޒ'1�<_�{jB�%J�'�7I���$���j+&�⽂�I8։�$)��ߡ��1PZm��^�p��w�ú���hA���}��-���s"C���p]}���<f�P�D$<V�-�����8m<�gt���$
@g	Kl\\\�\��oe���๪�6�Q�l�\�8/�G��9��h!2Bt�!1�y^|�s���:K���p7�W^�qʈ���S����j����j������t?�mmW;�x��0"S0i?�,фs�����=�'1��\�aa˜��d�M��ך��q�|��.%R��E���>:���vb�#�M�˂8�|���6�%�(�e��[�� �7��	c��b����L
����t�s���S����3�wD�*�@����<-�4L>U-�j����qkB�Գ7)e��S0-Q���>�Dd'�����Kz�b�ZmG��:�8���&mo�S��ɘ�x4�~�A���ҿ���Gx̍d�.{`#hB�'�/i����hgw��3M�¦F".e��Pu
M��^;(����KM�o��3Зb�����Ǘ��� x�rpnL�ͯnO��P�[��9#��p��s^�%2ƅE�_:*�nPZt�'��7�	5�%V�3�ˁ���o����F4ȵp���Ua'��D�7`�c4��/�5j�d��4'h�D��"�#p���v���Dj���W��3�`k{'/cU��)�1��_"�1��i0<�^����[y�	�"����o�������;+a�iL��Q
�9t!Vs=�k����j����ngw�����j���E�j��ٳN5"���*
{ٹBz�˶�~~��DG���&6��Hd3d�7	9���M6#������{`Wۣ������|��i��:^�<(Ӏ��\#B�!�1ɲ�wl�N\`'�}:::�AoL������ü��K�n��ˌI?d0�&8n�����������O���c�������h��s	�pB��o�ћ_~�'{��lv$Y^Q����A��s���[��כ|��� �P�Bmb���H�ܑ�����Q[�c ��D�aT<TO��X�`1�������ءD���1x|qq�/������s$I���# @jQ����������@����.�no�ۛ9���tO�.�:Z��?37� ���RT�u�B����g��ddR/%1�f�(N�c	gHPG

f��\*�&���'�5������[�[�^�Z�C_���p��+����l��y���;;��[aV6����)u���'��(�	0~u��5��>�R������G�n��1��x=��k��Xߖ뿐�@���E����q�\���|Y@;Hyt�R^i8�'*����*����*��e\�˦Pf�b���k��Ș�aw]��>�ν0GN� {�9�U��$y�׌�^Z�H�{�F�"L��s���re��9����^����S�>,c�-�#iA�!
�\Ʀ-�ϙ/^%i!*ߑp�	ŷ\�dV� ] v���j�C:���[|��Y	D`0�����vV�H���Wtxt@g�]J�
�u, �h�`�/���#j6:�nKskk���:k)?~��v��9]ޫ	P��s�9c����x����j4�%��o�.Tv� Sh�� k&�̿���g-E�:���D�z�\�����4�y]ȹ �mx)	����ܤ4��Ե�Y�WD{J֚�.R�x�F��I�q���|Y�:��?ǥ��$��U3�e�
+ qq.`Թ�a��6w��G���w��#X��޾�h�Cp
�ec��NXJg�]g�\���
u��uZ��^���n1����^"�a�^���q�,��.�ް�.N�1+~_Z"�h�n�-8�(_Ye�UVYe�� �B^�bi�K��e�� ZqC�a
ۭ�*{�l��1R��pNKeX��&9b.�%9��KPZ��e��,�ߧ�;��տ���6�j�%���Mnϝ˰ ����f� B��7~K#k(���%c��i��&l�D~@e����-����.����5Z�X�z=ᴒY6�H����/�ʲ˭V�>��)��Ώ��?Rxλe��E�L�n�P/^��^?pj����v,���Ч�}D����v��1����p�^�ӓ:88�^��sSd=
�B㙆yO��Zx��0*����`]O&��l=�g:�O?	 �������3|@*�C�@��ԧ񬭮�ޣG����Q�4��,k�
�̬h�͓�����&�PLyY����v)���7��)��nӣG{�BCY�طn}G�]P��XcY��֨�i���&/C����u>?죹Ң &�,3�;�U�����d*LckQ��؝����q��,��Ն,��B}��3��  Tf�~<��#�rh���ό��viOZ�[��^ߪc����*����j�ř#4���� ��|ֲ^�lj�����م��}?SE�+����F6>T3}a4��*�e�r��MVG�2O�L�̢d�F�2�Ǌ�� ����`�-�\]�J�,_%�T?A��-��Z)��hڈ`H���X ��)�&j���4|�>`[������2;p:�� #��-}����Ï�����@���&��v����٤^��h��_����۔���x�ۖt��NNF|,I���Dq1�h���.�iYt�lA��F���^x����]�LH~�(Y�<S�%4�n%
Z�V� "'�x�3�&���1������rf�L�r0�ۮmmll���u{]f�$����X��){m#MZ���k�6�otX?=Mhoo���h{��<�ã#:?ﺶ8t��5��@h�_Y�,%R��+�C9�O.�h�s�m�	kk�tvv�m�r����$�-���;�tpx�@:����B�c�d*�[�\��>ך8��we�A��C��n�ZTVYe�UVYe�ٲ�R��Y:g�MgbQ�E�b�l��*[j��.g��[�W�e��L�N���L�<�X灹tF�3��Ώ��PfA�� <�^��<�y�e�Q�rI
C��U����r7Ne(,��W�.�����ey��T���b�i� a��LY�,K�4�d��k`��Z�Z~9�s��p�g�"0�1������������W4�^��[�^�r� 4�������;:;=�@��Jc��&u��p���]���>��Sw.m^���G�Z��!�4��zfb"2V���i^��6�|PA��cB�ZpEFW��0�/�ff0�g��lWT��g��lH1;�����I�B滶;~��3��00V2@Y�+o�E���5�n�mb�.隗�`�2֟�t���ҧ7�Y�{�mU&����t<��`�5����N;;�,�aU�Ӓf�sѾ�o�I2�g�.�1?�Y
�f���4�/�8ju �M~eS���0�뉾H�|�ڭ6ˉ����*�Z��v����#=��Y�EM��;�������ם���?����U]��u7*����*��~��Ea�{�3�5�v��GxQ!˗ZO��+�L� _.G���+i���[S�	��k�@�r�7���/���um�$ta��ML&{=���U�d���e�z8y������Y�԰���~ �A_�*>�C}P���	{> Ķz c@�M���"ߐ�ߨ$�s<+�h�3�^��&ӄjf�Ύ�����t���,��^]���/0fhs{�66�hg������F:��0u�Uj�Z���������~��G:<|M����T�V3��f�=�/��3��/�?}��W�n�������z��;�mZN�m�����}���=j��rl���>���W-���g� u��v�7�4'�Uz���"8ghLs�D�M:���y�F�GToL�s^��˔�]���P�� 1���q��)�gZ��	\(�'�1��q;0����WMř�h^ �#d�ԭ?y�n���/�	�W�^,,�H-�&�2;��6�{��,�y�\����S��lI��З�DE��g��VK$)�g6w���l��M���V83, ϸ�����-�G4p}WZ�����yEa�ݪ����:��g��H_��,8f���G<֨v�>$�d>ɹeV���(���~�����	��4`��5�m�YX�"���|�+����*���6yc=ӂ�Q`�����ϔ�`��P|�Ÿt���2Y!�%gɁi����ܕ^$�A���|���[���C\S��Bdf��g��g��[�VcY-����L�/��j�:�!�(u�lW���e�D��׺��T�w~�ۛ���� [dT͛FJ���Xp<��L��&29(�)�
(�E�Fy���d�3$h��8�ܘS�'Sag�`�T��Ͽ��h�LJ��C���J���4���ϩ�5�Mn��u֩Y�ӷ�|C�����\�����p||L_����;z��5���Y���!M��}V�2{=�����֞::>��/_�,�Q����l�9�����Α�P�8Z�W��Z~�Q E���W���3:==um�K[[��yy<c)"���X,[H4�{������гf�%e,�
J��S� �BWZ�+���y�����¸��kr �f�d��C�a%Em�T�Y�7uKG�w ���h�=������,hZ�F!>�^���� PZ�x�/�^]���Y��P ���ϩ>�p�T���n�eyV��UF��-��n�-ص]���B�S���,��dA�_��O%G�� ��@[�)o�,����?w�-WDJ�K�&Es�r�U�^Ye�UVYe�1]��s���eH�ts��&eB~8v>�_@����Z\P�;��,�����˯��~u��)�$I���3
�{����VV�C���F�e�Y��Ohw�I��n�w�T�t5����E�N�3�e�`kn��[�K�e�6S�Fj���K"���7�7�+h��AO#�!���S�Z3/���� 0G,�<P�Gv� �Jk��5���2X�yP�{~�)�k��4�aƩ�R��V;k�8�x<�z��14����E=?�җ_�����[�Z� �vw������13.�cv <���_K��z�u{=����CG���?��/Xg��^c�Ul\�4���E�"��_7[��D
�dzS���ah�'	
��s]o<{h��Pt��&��a�@��aq�~.y/�7�ᐁ���*)\�K�x��,h�s}f����7���`)?/|T�d l~���q2qBÌc����k���T�٘-֒�S�v�����'��� �s�m2a`y6�n�)o�F�k�	��~0���@�%�1��8�|ŋ�U�Օ���V�&(n/�t�ʌ���/eŠ �g�`bYd'3�}�l	l�k(�H�I�%	���j,�N=���>/�.�`TVYe�UVYeW0;?�
x+~��uH��'J�"=���2b���z 0A�r�c��~�����H�K|��Hȁ\��b��p�����q��t�pˊ�}�
d��6-<z�����#*3�<�3��rL`2�;��Uh����X �Pd3E*w:�����ħ��q��ɧ;�|iW}ٮuZ����^Ia�A�,��&45�Bφ�1�ːm``����)&��:�����ʁU��`��܀�Rg0)�UCS�
3��	M'3ꝝ�w�G�}��3j����Ni�ywD��}�t0�o���3Y����3����۟�/�������9�z�����8�Ω8��>�����p�LG=o H��9�z}���6�6�5��n��F��Ώ���_���/i8����*3��N��k�£a�F0b�����;fZ�.O�]�o�*�>��/�3���%�y[]�p���9�=���?��mf �Y�?3�Y����g}�¶99H!@����0��죧���E�!0�_�����OXlf��ҳ���ħ6Y��lee� 7&8���5�E��� �lo8��qeY���%�� ���_cMz���V��1�@V�pGC�<4kjwڮ�i0c��iׇ���ղ�i�0����f����@VרV��u$b�[6�x���+Bξ��#p���2�`���?�"L��Ӫ�0��z�����k��p�q�9��$=��\�u|��2ߗ����uPVVYe�UVYeo��~Ad.�e�
������g���{L��eX.�eR�G�	�֘�
8��ưo�5;����S�nw���"�k�`3$ڸ�PZ�I��DD(��-gRe�ݮ������g�~c��l��'�}D���R1vS��l��(��wg +���EC/"���F׿�7������p�CV��������t�gi#*l<l�a�L��1s��X&?�@9o�D��Oޛ��A�G��Zi5i8��x��촞� ���kzz���>yB[���u�ɋ��x/e����^�� �����\Ii�}�����/��0v�|�x�x"��l��b_��&;�Fۭ;aYKp�j�c������Χ���'�>#��ݏ�O��z����
�� ,�h_&�n�L������ �U��"	����k}����&���jȧƲ/�tvv�1$(�b�g�6�ՅQVX�ho`C�o�ܶ�!��\a��f���$�<.F��!���O�^�b��vooO���;f�Im���c��#�bmu���<K}`����Ƴ�f��$�V���k��l���+�B���b8=a �Ś�7aXc@@�h_)(,iY`��^��u}}-8M �1� ���# �,LR޶��n�]�Ei�f���f¿�o��]Xr�O����yebs�"�|ܳ�`�lt�� �|���3�_ x���O��cR�/�c~_��w�g���1Y�Q��	i$�n��%YTYe�UVYe7���V����~8c�d�Pv~X�w�|�s(O��2���l=��8�����:_�z�O��c���}��;�9��;(����;,�X�5B�]`X��\.�M�>VVٻ�+C�C��Y6��7U��l^�#u�#R�����)�9���<����X.8�w`9k9&iF�۩�νp���ʦw&lo�ʡ��U������s�/�]j�a�I|�Q��d��YKc,zQ>PFi�y�:Q���hn�S��b�Bi��{ȃ�JKR���������¾��j�[�Ҕ�z=�0�G>|�#u�k2���@����HG �mB�f]�� ��0x }�Vs���Ɂ̦�Ym���:zǬo �׿yJ�}���=�n���#3�;k����d��j|�<(R� I~-30�]5�|F�p���Rq7��O��v�����}|r���ӧOX�7֒��,4���嵄k��+ �hH���#��8��V�.��{���K׾h{g�vwvi� ��f�sQ��S��̳2X^,`�o��l3�����%��{�k�[ Θ�m�db�k��][p�ߌ���H�D@�2&	k��,q3u�o|
V��uר�e.p��E� z⺮��	
��\��3`�h\�\����}�\�I!�c�V=�v�_ń�{�]�٬7.�/��o������T�j.㙀^>&�x�-��~�ۈ_���*�e���l|����UVYe�UVY�
D�K��^����/�7�y�{������tv��[��o&d2��X��v~�-�M�H�-����7��;���3z�>%��ہ����c�S�43�u�Q�_�-"kD�7��*��.-���� ���iɋ6<?�),)d�G�dD�����M-�C���s���~�}��M�w���d_���=�)��٨���1�ĠX���1�Sl���] �;H5X��+�T���tC�//��Ǔ���Qw��mYSrk��g}�����A�5�ƈ��	�`�~���������A_|�F4[�_����!���׶���ɩ{�������[:8��z]���p
��y�?Z���7�7��������w߾��#����ljh<�R�6��;��Sw,���?�������:k�������:8:���-�����4�#\��V��/���V�[�f��,�%��~�<���u��ݴ�Wr��н'F@�~o��7���~�	������_�mJ�|�)}��/� 2�� <@&�ufM�9�����m8��Y�� ���3-�bX6 EN\������ �<yJ��;n/�a��:~wE�_��f�Vr��n]������~���k�TϽ �o��KG�cf#�4�@�k����8G���dĹ=���Ɇr� 9K��9X�4����ALL2 ��O�5���䏮�&o��W[D �K������:��u���`0��U�.�13>}����:�k7� �M��qm�0(��F�o��y�.~h�{�^������'�A�o)��(_��k+����*���fKi�g�2�^?�uc0 ^��''nNxBggg�'p�k_s4d�6YKXɐ:�{�-�|*����}�)��Ǭ�?�5��~Q��@������68#�I�n	"��uoG����)U�reѼ�U��D�c�E�����o��PL>����y?�}��c�E�9a�/Wm�����m�Y�>�-ֳ�li�pD����F���d�)�����%B)�֚�}������C�ލ��n����)���4�f:��t@v:�QVc=��� ��G����G�7�w����R�O?��eS!Ce��V6��|xp�����p���俹Ң��M�{�G������*��n��Sf=��3�(��4�Ѹ���=��~��_��~���^3������@��Kv��` >3�$�g���@���ε�
d8�.�����f��OW5S�V��o��/3)6�Hik{���GG�trrH�fݵ�MN���p䙰A������	��x�EK��K�1PΚG�<0y_�z��4 �vwwiow��}��H��;��i77�6���4�x��PRfj��c�M�He�)^��2b�3���#z��	h7��"g�k���
F��[L(�>�rmm��������L�x�kf��,�W��0�K�ZxN��%?S@eM7�&u0\kd�`B(�p�7�{�8X�kk�+a�0��>�x"��e7>�m�m��];&3dV8O69��{��X�?O� �3����b+����*�����*�E6�d�e z��
`���:�b�\[A2��ǘ�yZǽ %�L�z${�r&	��P@�����ܺ`3�f�� ;������^���q<�!�):dU��,7�tI�R��Kg��d1*{Xv�9a@m�5Xz���,� �[��/�������*�ξũ�l9׎�g��c��ð;���֚Cˠ
�~Ϯ����ce.g6_�*�α�����A_��S�݂��5{�ONy�?�h�̨>���M�k-zux�c�?������;�������o��h�GG��-�I��0�   ��~F?��3諫-f�$���/���lX:>:���<�w�)MV�������O�����_�W������_��3����_����?�������Ai��ۜ.����s��̎Ba���k����(*�_ˌ�����m�%����X�!�3�J����}��)3ݿ��+���w�O��g����lM.b�ݜ�����P��lB� ƌ��D9/� �z��?�s�%�lC�����k_��&��]�j1���X~^�Bv����cn���'����Q྇n�j���q������Y��~3gGN�k��.������j%����&8��F
��[�P�n��/��GO�cI��I|p�/���/_�׋ ]CaE������r�:�G"e���,��
�t�s�k������@3���!�����	) f�(<���~v��*w?7�x�y�y+��m2LTVYe�UVYe�3�K@Q�~����b��/_�`�Dd�e��A�`�.�ȄLU�d��f 
�'(�y2��qѽi��x�i6_��t�]�5�:(��c�xrzJ�_�f�4�e���7�~um�v�/���:��1��w��[�U( m*���Ǹ]dY񳒩�TW	M|�V�,�y0$H�y���D�2T}�؜�����k�	=����J-��lZ*�6|]�I��@��ae�%���"҄��Ǻ��v�&���{�����_��%M'�C�ѣ��;���ɓO���_��_2�����1���^��3�37��������Dg������`mNK͕:���a�λ���w�����C��m���������I����@G''n�5�$th}c�:�iE��4�l6�4{. e��a~���u!BF6��0���5-,�P����� ��8:d��/����y�j�^�xN'�G���#��/����&��v�)��<����,)�X�r�2����m{����/ <����G1�
@��ؗdO\ے�75�� [� X��FF1�8�+
�)�����ݜ1��o[� �D�� kَ��f<q����J��jy�1�w���8�%6>�����aL� �(�����gg6�H\ l��j�:�v ��"�zAq�z*�v#��IR�4X�:h�z��M�� �p�˦������d�ei66�h��*�ed=�T��+����*���%V�G����i͟�����|���#�R>;�a4�x�l}}�66�y�F��K�b4&�����V
8!K�؜�y:��2�����!xwI�:)��2�y��g�"����3�Pp~��Φ���Z��x����*���y�*Ɗ&r��=�k�;*#0�n^����M�����L#3�0=ԝ�����+���r�r�RSJ�)�����Ue��� dk\P��L9�9����) <���֪�9M�ݢ鈡T7Rgdg);`��~��������}��.���������#z�d��N'�s�N���F�);���i��`G����K_�oƠ�h;�P5)ԟ�)�)}�������?��?ї���Z�G��6�dXi����P��3�Y�.�j�8
_+��&���p��]j&��*�C�t�F)�� ѧɷ������O?eɖnw@GǇ�L7=��ʬͺߎ�Ԇ<w �B@Fa^��	�w<s
���>;Ő����������Tn��eF� i���K���wކ��"}��ƖL  �/�T��� P`�,�0��8f�ѴIގ�a8"�Dr!�9 E�Egv%�R���|�e:����d/0C�`}3���{�H=�Գ�;�b��/�(�ĸ褌'o������� ?	��t��"���q�w����	�9�q �U��Qȭ3ٚ�d5~f��_e�UVYe�]l��d睝x��D�,	�t �Ϝ��z�5�IAb�󁡼�ɾ*d�����'l5)�XeMc��j'�텹+37d���6�D�!1ר79{
���4��A��Ȥ���]p!���7\]�9Y�OU�[����V��ǝ��;�?�3�}��|����N���[�x������g*�[�?����\f��h|��DV!J��p�7�8���Ŝ�EcT��#`i��}��`���v�?35�[�����;�Y������|���9+<�tYw��g��^��??�ӓ.eSÅ�� �L�� p ^�xA��p_�n�ĩJ���<����O��/�B�ӟ���:�5�z��v���G�hu�����^��J�kvN�����O|-"�>��C
V^p1w���P�.׶�{�,W+LWJD�����f�	K�@�muu���0��O��D����=z��	k���o��1pe�N�cM�ј��/~�������BC�W��5}��'���F�@Z��{����Vw
j��������u`�3�Әfm�}�L��J�~�����g�`���~�3\L� *C��̏)Rpo�}-RX�=���c���@^�ҏ+�J�ܙU!_i�MgF�fka�6,�����}���+@i�q��~o��H��G\0vccÍ;�<�b��TVYe�UV�f�ܢ�}�ey�ׯ�\���\7d��n�l�s��G�h{k�	G�;d��yr��C�ђc�/��$Ql��t��`�����������#z���;Y��{�sY��`2ïΥ&��*�`hj��C*\����"r�~����D�0��u��af�"��r�S�rs��``o���T�����&GU�������L���'�( �tc���[���x�%.2_DN�/PP..7��=��R����Ŵ�љ���B�I��	H�:�>��M�لfv@ȴ���������E���V7igg��l'�����CT�NiU}W�o��j6h���nsQ��/_�W_}��3j6�n�� ���k\@��_�+}�׿�7�|M���q�J�&�л;��^�5����6���h��Q��;8$Q���E3/R���f�U��s�,[�y�u��O��i�F4�%M��k@~��0�|tt©��^�dG��HA�N��W.������@$ �}vΡ���X�[���ѳg̪P`<�5(t�^��?�^�t�
('o��_ЃX�@?�OC���`�Y��^�p��J�ǖ���/��,�k|S��,�T��G��>7�:�c�������m��O?A�����Y��:�"}�l��C�d��U��!�v2�]ìc�,d�ڏ���X&"��ci��3+�N�.2~]�[nb�b;�LAC� 82ZN���p�5̸�Y��i������n:���_��6�x?m�����*�Q�.l�s���q����$_��\�ϟ?�#� �9�ƾ�����P�����1�I���ˁِ�$�D
�a�mI�,0*s@sJ>@`��6��'��x���@�{�|"��O����l��4��*{�-���J ��h�<�\=�`f�Y"v~8��1��i��i���`��*��l5��c�u��a�o��O����9�v��(pb���2c9�`!�7�<����(,s�)H
˃��DY���Ld����~bPԳ�|��.�6��e��G�( �X��_@1I�'�p(FÉ���i:��׈l2f��&`2g|sϺ��P�vd0F�&�X�w��ڠ�1#�W�>$�67����r/���&��i���6��6� hq|zH��o�F��=�#�G�9�f����kk���I�@H`�60���齒� �p�56d��d= $�,E(��c�=\� [��H<�4���y �.C�&un[ �T`gg��_�ӊ���G̖���6Dgn��38萆��R]����uյ��-vtQ�L�/ڼof}�I���U�6wr��
,�km?���Bq��N3V���~�����@�D�$F��Xu�[��Y~����R�MB�sGJ_.��\?�|i�N��x��1�䃃}��1���l6�g�df�?y��g,	�X��2K���|����K�����������j��ز>� �V�??�r%x �xvP�z�m�1e�_u�z�'���>,S��v��,=(���}v�#����R`��s� k����8���0��<�3j� k���GL�@>��yӺ�����\t�q���w��`R��c���
�xIa���<�Z��Ln�i��ysp`�Oݯ���mK�S�~ :�)�ҥ�
�4�(ngKZ���X�u�w1��T�[�� �?D��(�9�D9���<�wlqg_ ��¤�siB1v������;�CF�ew*����$xI	-l0��a=�l�(ҁ�ږY`9�>�`���(P��d�9���A��jj�L4L��u+��L@4K��,���G{aP������g} ,��(��T|���S�2.� �J E
�7�ͫ��*; `bB��_��n']j6kIFA���S��뿺mpj6jH�^i�ܱ"ei��gϞrj6
1�NV� E,��^X��F��=��_z㯳h�j$\�{��졙j�]��&���+�� F1?<�H��>,89:f��t�1����2�48G����&9���fl��s!�li�>ܡ�!�X�ۛ2��,�*�݉��Φ�|p_I:�̄�/��\��1J��5XG���YRb�L�{VG(��ݣ�?��676�q�c�N -���c�qƔ�T�Y����
�ƍ�u�c���ā/�Y�	R4`�K���.�����d���*{Xv�.��X��TvL�=�R�����W�_�\�x:���n9���(`͌_7���@�W'��C��J��{��H����,��w~O�<f����C�{�d���O��y	�(�.���\Ye���#�?ܲ���/e���ʾEE�=iiL�?�<�Uws� ��%��x+9i�DdD���*{���<��l4^���D>�X�)8<c���c^Wٳ4Vp����]`UZن�ٜF�q��P��'ۉ���u����� ��k=X s�>M�c1�h	�����v.�t`R��߯Г�GtvrJ�n�s8���!���f"OgC��b=M������1K �{��%G����s��s�N��uf*�=�e'�>���5��L�E��7�o2�R�����g>pP�����i� ��2��\L��!Ή�������q0�x4f:�K�$E���t/�˂�	 ��I�\:��A���q/����^�ȶ����;����:�N�8�X����J�$��������|-z٪~5L5�qpp@g����E?
C�/L�@ $?*Mo␚%K5d�Ae�
yxg3�4�-j4[<��,��K���,��5�r��C���C�*>������ƴ�Of�Y����ӂ�4C*�'��
��>�1���w��{�'���܀X$`l-��]�C56���n��R�#o[�A�ʒ��p�?l>d��l���A���_���Yj�TC巕Uv?m��V���5rdyѼ�L�
҅K�Q��&��I�#)���@�2&̯s�ЗU��ô���vL�՗�C`���(k,�|� ���Lʒ�)�L o��$���˙/���T���Y�E u��1 �,��?xK!��{a��W�X�5j�����X^�����CJ�}�tQ�@��z��`xNGG������G��G}�E����ѿ�˿��_M���%6NO�����sa�p''����+.�pt|@��;.�l�e\�zZ�f�E[ۛ��x�91�����d2��ё�z!�?������)��P��G&i��R�U�P-�L��]���x��|�v6�����mZu�6@���ؔ���m>�e`L <��K.K��﹍�D�����0K��,������9v�"soL����(f M�c��xQX���]��X�z�����o��ZT��ǟ|B�?f�22Kt��o"����od�oL`3q������ѦZ�6=}��&��g��B�X�3`e����$s���P�==�{c���<�>��ػ�n�вb�����Xթ|0A�)�i�^�s��ztt��
�6u�'l�Td۔4��|�Х&��ā�/ϻ��N��cB�r��̭�M�A���s����K���|�_Ȫ�z��*{˶d�.HH�9Q��b�~1-��+�X�'���E@bQ�=�� �f���m���������R���!�;ƲF>|�E�Z_JQ
��F��FX�3�R"ߤ�Y2�o��y��lfX8!��g�%H:([�
[97�3�o&� >c"G������3��9��� �V���p0���ᄎ�O����Vlo����6�`�� ��pސ�8>>���Qgu�Z�7���]ِ̓���)��v�H�n�{�j���S�Ȭ3���gi�I �L����&&���غ�ms���x���W��m1�W��[�L��
�3/�"�X+b�H�$�SU���6����e�qV�k�$���#���Q`]h��wGN��}5R>%�cH`׃�)$��yl�:���R��y���"�b,B �~�� ���O?��W�h4�y�2iЏ��#�����W+��C��讕!�E���*\��ˬ���L:��Z� ����<E��X�A���A\�>
�$�+n��h)�$r3����i�h�Ll��{�����9�9"3����T���*�M�:Yj�d���&g��ϑr������gP(�\q�}ղ~+g�V�>ڝ2�u�R��[X��}F�{}���g���bM��o������]�L�G�=��e$a&�T;X �< $��{�f���H�x�7Ok���֖�C1��:��T�9�"ũ>���)�����kj�:�h6��
��wvv�m�6����g�:CJs�����a��wGĺX��Xiv�A�j�0�6���pz3t��|�pty��欤L-�r&1YR%b�|4�U��Z�2��B���Pu<��4ؠ�o!:JT2,3ۯd��Q�vn�$����ֲ<��4�Zp�#9��Tv�L�G3w�����(bF���.��nF�bA�)aPy�&��[�&��;'>(�j�|���"}�Z�rNZd1w�f^�?I��3�}���k:kqV�S��2��}><<��;ǳ�3.��	0@r��L�pb'�*����d��^V�_fW������3���W?�����eť7fp�t`S�tU_��Zt��g�
_��4��/�����������N�2 ��\��1{���#0���ٳg��>�5Q�C���՟���fs�*{�v_�$���c����O��~�E��y��*J�{���
���T�ڝ�+���!���?�5�����*Ӑ�S�r��㹘&�f�.0c�<H��r�Y�NX��t�"������[���>��5)n�u8�2Ҝ�T�������Wn�n�UO�of,^5q��N�6�����L�5�!a��j{�j��$�'�ބ�6�n�3�-�7��L��F�A�봹�Ŭ筭Mꬶ���s����"�)b�}i�r�2.�%�$ꬂ�������Lq����SI���x3:��[�]o��{��X����|��-<�<�����ゎ�E����ڂԂ�X�[����y�S���1���gˣ��
����#����C�_��9 �����G2�w"^2k�Q�rp�S0�ݶ�v+`C���x�&�;�v�À8�!���)O�Q<g��8"[ �z�{PYe�=,�������Y��ƾ�U�eet\7�r�~����^���Ȕ}۪��PsT�)���e{�'���H,�<��ӧ���C��(��f��e��,4C�*��CH��D���W��%}��
�A������� Y'd�Z�W��M�]�v��K37�K�3�g���1���hvct^�����U�N��`y�I/KI@%/iad��)��/��x�L�/'�a~�w
6��sf�k�=B,i�3n>Y�T�����Ǆ��S�$��.�s�LDz�+kM�e��43�Q���r�_|����|z�J�!�ddY�x:��Kt����d�z�""�c3Y��)���_���t���t�����{mJ��[h{�C�����!5m���t��;��\�0)�VcY��r����d���Iچ#�p)���]���Z\A�X�:͢�Y1����Ж>ϕ�?��1�OQ�{S~�̒_�ח��ʠ)�0z���������e�A�O��ݥ�?����+��x]p����W������|������}ߌ�Ź@�1�4\lȍQ��J¸R��+���s���~B�s�����C�)f��ӠO���r�Y����.mM�E s�ʂc�N�і>T>ieo��$��Y9_>��#��}���YB[[[<��`s�=�߻�;bb�`Db��|Hzl�opf�0��W$��ݝ� �XYe��ܮӆ.j�1Z�:��'�!�q��U�}H_Q{���c��P�6�3`9&��� Y��$*+�X d�g�I�nƒ�b�\v�K/d^w���a���	��zє%�@�P�d��9~�Rl�bc��}�<��XT�űwz}f3�5�MiЇ�ňƣ)3�q��qB���4�k5 Pr  ���p�Q���5�&�r �������@�A�C5?��2�*!��'2u&��Z�,����m.��GU^�5e-k "�"f�2��K��!-'���^�U�C4 $�#�}~^�&-�h]�!�q���l��0}3R<OONX�He`(?~�Y9�W�&���Nx&� �?���y4������m��q�XO�
F6���|rz�i�`,# 9�����YT�P�6��2`�����X�<��-?W�`9�Tf~BYw�G��t�0���[$wt��(w(��]،$�����:��ܯ]$��͞�W����tn��υq��9xއ��+d[++<�N�?�y�\���Jx���6�W�ٍ��[�R�2�L.w������eaU{;�[������?qe+�n��m[�J�1o&0cP�0���ᚿ�Ӗ��[6w�X6��l88.g��W�|JQ��`Py
z1���/�4F�]HZL���O�#�A�#Μ�oUGS@kҋ��ǾP��>�?s�pN'�$]�����h�丐��> \g�)���C�V�6�����K�n�'����u��S�^�;�z4i�=U��$c��B|�(k6(qǅ��յ5��C����XN�&����%=)˦9�쵐in�����ne�da9���//�� ��S���	%�����-s���]ɖ8O������X�h�Z�]���ٕ*���t>�AB7�t{�t�=���x�})�x�?���mb��_�1��������0�)�A��.j��o>W����t�h۝O���}��A��b����i\�M����?�'�J�GQ�T�[7���r���|"�o�2+�i1��7*{F>�5���|����u�i�?˯�+�3�ŷN0����$Y�VLt�ZW���}� �)L���Le����|��{!�	c+���P��+$
��@������I�S��8�b$U��)g:T���2>l�w����*����ta��� c����_ ڔ��$��f�T4?L+!�7���{Ʋ���H*!>ff�e3�:濳�K�"&4�&4�D"�ja�K��a�bb2���m��%D�;�������d�g����xx�MDVBe7�a|��e7��u|a$�w:-�@�r"Z�,�A"��I×"J��CG��wLx��X�y�T6y �|��OH4�����MB�v���Z��(��ߪoy��+V{��T>�Y�3~��x��f�(Yك�9OE�Y'@T����O��K���b�:�s�]��g\,���YG��q,��=y��V;пO����|��3��
����71�����#�=��z�h�����
�
!���]O���6��ή��j����������Y}�:{��5�nҌ�=Q�H��t����>t�3?\����Rt�������S_���5�M����&�\����itr�!�E�	�%�8�0I�A8���e�vp^�f�:�v臥8����g����y���6:��zY�(s1~Q>P����#��^���++|M�D�B���0�G�v�����!�E0 +����v�C��2�?[�γ.�|^h��C9P��/���Y��K/�أׯ_3s�	����w8FYCTuܢ �[����j��;Vs���m	�	�����J�%1�ޢ_cx��J��ŗ@�6��w�L�oYu�v��r�I���g0��)ѣԁL�����b}3�`��\8�c�Z ��3�gS��%Ҙ�|�
+�A�O��_Tuzm�r�l�լ��lHu3�oy�X���	&�(!VP�r�;�p��+ 1����2�&h�QL����n�9�^e� ��+�&����/�D�|�&�!A�����,9blw�轝����j���aU�m��H<�)&}��$ZݴT���E������?#�x�����+���U�R����|��񢔩7>RtF���+�p��G�e%
������V ��O�����}�ץӳs��U��`g�=z��!��C��<��}f9��e�[�8^z6�����W`�@�CЀ�j<�^"�i��.ϙ/ 3+���:}Aؙ���վ� �����3W  D~���`
J6YRh{� yBm�Lo4;"b�4��4���-y\�/�H��u��$/�,��ۂ\8�˾#�����/Ɉ��tdҡx�J��Y (ԩYe��W���'V0M:��M�ɒt�)� �erͰ�^���g��_��D��X�w(��x4��h@����g\RlW�-������k�C��.�HݱG��&����a�|ߌ� |f��ុ@qd%
��y?''I��z���k���k>jx_i��O�ݡ]E��|��V���� 4��x.��7x�%�g.� r�]��˖�,�C��zzU��E��j���W��~� r��2�i6p�w�IP|���z����+�lά�1sak,�5f�{;�䢭��Zԛ)����o�\�A��du_vZ�)�\J�kQe��b8�,�?�j� ,g���C$��??�3��b&�Hcd���F��/ �K9��p$G��vi����ym26���w�u��8bb7��W�Z�b�]��S�oE�Ò���Yu�49@�h�Ei|(TN��RvF3��ı��$5���n� �u�\O'�Ұ��ib�qH�gS�1�#@k��ԁ&�@��5���œ�E ��#�8�={�_�iƚͪ�m�ð�0���gr�Yi?����g�1��q�J�z��0�,��e��Cτ��Y	+H��q��b�p�K�Zd�څ�]�n;y���Z�BP9bw������^�.[��� �u0�Pe}t��ˠ�[c��:R:�tr|��*&G �=��O���y�}���Y�֟O�0��2�.8�˦\�xW�q�ǂI���:��F���s�}��Aك��+�l�)���̷��,K����!9�΄�r� �ɴ�~����i!�g��<0�m ;�:߲�b��H3Q6k F?�$�/E������-��HG�	���� gr�v��������0ePlA�'���h�eop<�Z�پ8��G��x'���<v�rpp@_}�
B��W���C6�g������O�b������˗/}�k!@�;\g���?�|�"0�v�E{�;,5��HǤ��2��y�x���]�tƙ(��1��o�����wv��Ai�%8n
g�1�����7�2��h����⥰P98���<�,�� {w|����g�IևYv��A^dוx��YXZ��_���e��w(�5�.AB��G����0a�Kf���f�K���*y��o���D�� ��cy��3��R;���H��<�^��}f��K��5F��v����<Ms�p-*������V�w2�=s�bPe�oBZf����#�l&=:` #�Q��'���k�Y�����3)�d�@i#�"�1�U#r���6�zP3�~3�.=M��M��}�	cˆ��w��)RC�N�ӒV�dc6�0H�B 0�)��C��(:���
*`v��� ������2� ���MBXt��ϲ� +�9�O�p� 2�����7�������Jz�26�����8��@�@Q���
��kW�����)<�'bp93I!���O�����F�����۰�'�p�>�y�s��^���o\<Sa]�咜!�����µ󀍰Ԓ �����)!��e0
=J��<&�FC�"��Q�C UH�c��X�� �e%���)/�����L�����n��4�Y ���Z�	���hZ\i��T���=@��f#���½K�u��}��l/�!�}��wrBi���kks�B*���3.�Ӕ�0M��].��@<�`�b�h����!:�l�O=�omG��� �h�k.l���?�o���z�눞��3(��2�T]P� ��<	��t��cp�-��%m��	��� v,C'��;fѬ��, x���q��n�˿@���V0��_�H朞��l��	���m<���r�;�@<���	@�Ѩy�J@7-���$V�R�@ 5�}���G�mnom�>�;_�C;kK֟��ޛe���.���<:J�W����k?��{\���<BC�Ǧ�ߋ�h�ƛ��?|mS]���`9 �`Y�=�L��fg� ��sє�"�ףLb�_��7���ݼ	��0}t>��Y>忉��/�s2O�/�>X�k������os�!���2^�m�H
|�*.]�ó@�ȗ�%�i?S�3�w����|�a���sG��(�yłe��#往�߲��!��}�c,�ƻ۷�i�{P�wW�O&�EZ:qg� �r����1p�H�t��,L6$]zҨQo��	���E�@kx�zJ[�D�$n�o;��Pt���$��_�Lp
�ܗ7�E���%�<p˅<L��	x�Z�*(�k�Ye:K��|�����[3�4�����U��S��/1>Ϣ�.��,˙��d*��]�	a��fU���-�x��Nd��,����?eF�- �w�,�T�،}�eS�J]�39\�����-�~�
@�%�U����<3�\�@�1��s˷��aչ[|����x��9��� l��<�ާ�G������������)�JFs�.�N'�E�2��1#I�i	�?���L܋���vx2�6&̽~�6��< Z`�U=��e��ޅ=B�.�	P�֟��YŻ{��_��<���Q'- �~���x >�?`v� �nB�BNf+���1 ���3��E41vAfL�` �>��^�z�����6�`.�|X �A���}N���Ǉ>��@�4hc� Lwwv�m�і�&AX�D+�p-��ã#��`㼸��;���pLD�Ɲ3���:����5+�,�r��8�D�ڥ���� @����uRvb��8G0���`�;0����7�k�A���2�&����e]��a���x�(6�,��N�e?���k��|�O"��7�������!\e�� �olnf���@Dfk2.�r>�����8���E�`����3uݳ� 0����2N2���DEp:�by��pۄ�ޣ��<��6�`n�.�,����H�L��P#캸����r�ӱ$����cƙ����a��}�k (���{�B�+{?L��V��x`���ª�qB}�l.��b)���]�����y������s���a�
ۍ�,n��Gn���n���w,{����_qZ#&�vlY+y��<;o�ȅs-�I	T�$x�&	���pN*��A�l�ӓc�}b�c�����(�܄e��l�P6L)AYӘ�:�s�M�#0��8�^`ڨD*#	Q����T�XO���u|�_���]~ygy$����`t���.8)9/�mY
gg����p,�)0��z�4�*���r���rG�`eo��N}ʯH�BPf9��6���?CE�x>�.��婱oɮ,�bp�p澗~O�r��u.
,]��iH��4d����]�G�{��.�i��b�`����h+^�C:�:>eb�b�����ia5���{�@i�?
��Ǘd���P������_��;��6W8U�@�o�z@H�VEm��ʖ�>�!�Q��6�m�=W N�#�|�Иu�����`�H�@����^����`�����X��QCϔ����X����}����jw�@Y���&�T"Fһ����	�h�6=�0�2���}�oq���1ۥ�M��4 +Y���k���1@��O��Sy��B[����F?��s����AUd!����l��9}�]#�̸�d<8���{�}��@�6�Idnn����m��+Z�s�]3����
�\X�21�;�.?'̀^[��g�-�gld�+��p/Lϝ{��=`;�� �p�-w�D%��Ϩ�>r0-f�ly��8���5�r��S�=G�i�}�t絾�������sG�	�M��9_��}�GC�v���2�чh�O\Wh.CT'�gB ������	Me^��;D��� ��T��ڜ��sJ�
Z�¾3�v�h@%c)I|�A5�7ԟЀ�0|�lE������q]�O"`S=���w6���D?��IئX;�.����c�,��m��i���\b��!%��\cѼT�����p��e��6�nBz\6�Me�b �s˓ L�'"w���,�1�ߍ���hIC����n���b8��盌��;G����j֪г �
�)@�r�Z+�� 75�vUrx�zd|Ǔ�N�  X1���@����V�^vmm�W��Qw�y��K���H�$*}O=�/���ha/6�3&��8Ts�}����b|pP}�5Ln]�� Qf�1�d˓�����&�ы�������^��CP���"`�|iJShS�`����}� �EpY �$�g�q����ߔ#��$[@T� �F�@�O���Ϭ���2�e{��ͨ�������	๰LO|������6��f��1#���:vq�3����O%�W����(B� O�p�����w���%dl�37�՘�	K�:k[���o��e�\p[�b�M��`���0�	�*�� �Q�m��p�C�h���vP\
��fרF0@c�;��a�n�%�P��)�j=���O#�+�W���c�����8U�|� �l��SZ{�~?���h0�_�z� .�������0�����h�����1���$��2n1`�"��ϰ��L��X������I��R̫���)d:೻k�k`�ɓǞ�-}�ͦ�8vǄ�1��	w��� ���8~��%A�A��p, �ܹ(��*�bs_��8F�팱����s0�9g}���S�99���m�빷�+��Z��1 �LNez��>,O{����1v��v�@��� ��i$ٙ~|������,�� t�	f�$�P�3�C<s?�e����W��
�Z�<#��3��c�b��DYO�i��X*�	�Q�'�|���S��Z�}�6��5��x,C%P?&��Ae���΃��d�L��Z?�ޡ/������y�@���*-�M���|pQ�Ha��K���,ܿ��� >_p�UO�f��aA��u��v��y1 ~<FTs,�?O,�*�n��@��� ����g.�r4
���cc:��U��ι5)�Y�7d��d4G���9�f0�NCa���U�30�㌪���S&��#`���S9:��b�O��G�:SqF�-/�e|���Hڒ��2L<���/�sz7ܖР|�����_�����~@�N-��-0�4��=�Q�%V���}�kAWM�(�KKޏ��m0�a���3������I� �~I��5��_A�/��((-��$�����
GOD�K{�;
 ������͍u_�&�S�a������m�#��]L�0�@g@�}ӏ+M7�W`9�j>=���5ѵ��t.Z~\��sh%H3~,Q`1i�?|�E"c�8��-WV[�	��/�Ae�Y$}�4��.���7���6���Y� D�2E;q-�Y|`���O"vP�nw����8�� �~�� ��o"��c�1�R.j��@�{��2�m��A����s��D��� ����
�4f���	����6�����
���,k���~E����O�>�wmDʃ�f:��/�� j�My �?i�Ώ�A}=��5@�Ld
K3a/����(B�g�| ����uק�8p�L(F�2�=��w�v�/��^��ǁk)�+��W,�}�2��ύ)<�1(�2 �g~6E.�VKX6>9k������@�@ ��V��_�#Ӂ�V4c���I��~M�\؜TԂ�|y�l�H�|O�j�	�1�,IF����@����!?��jF/�\,1�Aw�#�KM���f�������EB�bF��Q[H�%	c?L%(5��t�� xT�曯]�������2��n��98�O�z��D*���M@e����2��ķ�0�qA�9�2�����O��U��&�x�J����M���;���qO����*{K���E�q��]N#�3`��d2c`X�[Ӑ9�ف��&HqCj^\n�쩑w~�I<��)�n�t��ġK���J���8�u<�?dVFR����0Rά���%���m��ePJ^�Ǥ8¬ˬg�h$���V4j�]¬ac x\Hȥ�"&]tB$�#w���k#:b�,�8�K�8nD�}��ɴ��D�1�F!=4�̂�%?�]ك2y��������>%��"gg��\胄Y�U��M�,�������/J71IgE
�P4�S�B ,�p��\��|:WpL���l7�a	�Q�OC���^���	�Oм,�]6�36uB�w��a�mum����c�~�?����,�Lk���;tc��s�.�f�1���S�) �(0@��<�`n���@��bu���s[�[���wZ@@J�q��H�H�>�x�^��}M��觟~���C�a L>~���}�Y����z*�{0�����/a /�.���m��.� ��o�s0������	n�	ڵk E�	)��d ��v�W�"-h��W{(x��Z�L�{>>>���S�G &��/�����o��[9��sʃm������}=�[_	d�u�.�MO�� �TgMc�e��>��tlr ��7�3xV���^(ڷ�����H�̼��##%@��N�����~a���
�/*Kd@n2Z�8?-N�q'&v"5$f���w�nu� x�Ɲ���u>Q\�a�oo)(��3	�W���>�V@v��������7������a^���v��'L�ե��8�ky��l:d�x�h�,[�n��!Ϲ	�%n>H����EqK�X�O��Q�V�m�ܕ�<@^�����LǷ@6���۷B��/<���3�]���m�	#T
(�!
A�آ�07�,������,�_ə���E�9;�gk&~���k�}ne���x� ��PF:ܐ����ǚhp�x�:�T ���Y��Eq��>�p����uk/{��g��z�_N��;���[�=���Ӻ,���2�OLI{*��}���x(.8�\�y�c��A���,�@������]�i)p����}���_� @����:�;)D�0i�Ef���d�>3���yD�g�
"/�\��p����,˔ީY�� Z�394א&	�g�h)g����3�o���kn��>d�%-��"hG�?�0��l�e��O� ��H5�b���c�����y��Ae�E8, ��U��΁S3�t��S�����[`I��O�_�n��H	h?���� R/^�����ȮYf�v�0er)c&�瑿.2�є́6�}@V`�]�Q����,���@3�,)�)~X M ��� [�`⹅n�G�6�ME���+��)���fε���
��,���:��jQZ� "�/������]���0z�bM��z��:��:�+��
ޠ�F���LK� ) >r]�����@7�0��2���Vm�"AB��!��e����,݃��� ,sѾ���+@j\���4(��Ǉ  �C߅cKk�&>+W��%��L
�f�����.����@���}8֑���vHc�sMCq�o�־Ț�o*�@�������4��~�>��n
��!n�R]�R�8m>+/L�/�QeW6���CvѼlYW�$NTBA���O����dK�c��Ђ|�0�v)��!�D2L f!FIAQ3�O���P`��,������������Oiދ�3�:Z9_A���i=��e%_7)d[��!����q���3%��9i� K��!}ӽ�$��H�]��2?G[R��Ļ[v��g|g����da)HF��Y�tT���{�k�Y�K�09����Z*n���cw,]�t8ay�r�ه��W�KNǛ�S���٠�̠r&);�#�_,�����]�A]�!�0qvjB�6h(��t�ŋ�?�FP��]� F��ܵY���R[,(���eF~�KH��A@�i^�;������1�\�6p`����T�j6Sƹd�k�W��+���{n��"�!�œ�%�/���J{�����>>&�Wʸ���fӧ��tjtbF����8Eg�g�z�5�z	�V؏ !�8np%�4�2K�������4p��2v0��(R��˩����~�U'->ݹ�7Fg�`�������D3�����o�D��p?9�e4����)kjW�a��p��G������n�όW�{�� ���(��@��� X>>>b0��Ϟ}� * 0��n���<�Z8�EKXdT[`�k� N �l�o0����@�(����=j� ��
����F�ս�V�H����&��	Y!�~��ϲ?=���fs�fw7P&��*�sD+�� }w�y ���7�L±��� nAG�u�M�@.@UXF�<w gY���kQ�x���w�)ZAx!����a�uX� N������%����<����>��mmm3��uq�`Jo�����|�+,��(dDb�-�����֠�_ ���� ��^Ɯ��l,�bi�b����ܽ��L��4�F��A�r��k�izI0_�3�g��>�A;�&�m!L �7[B�Pz��_5\�X�u�Q�-5�d<�����>$��<ڨH�$<��`��OHƸ��R4�����(���w�������}z�)�� ���L��hQA��|;�Bp����S�2K�đh[�AL�� 7�I01*��7T�k��Ɣ���u�L9�������'f����f*{�٘����~��
E�+{���% j����{E(��6�Tc����*����5ް.O��Ϧ^��t���5��8�1���a9Go���ޛ�7n,Y I�RI���{gn�����Է{l�]�RI���ǉ%3)R[iɰU�H;2#N�8���`�,����)l���F�6j�����aw�?���}�$�wc�]��
�z2�T�����"�`=����t 0�!9h-��*��Ț���ߞT��?�gyh��&��!����BLwHH�?�l���VnʀsS���l���1���M�O��-��6a2�+-�[˞��{>���h�!p��� �yq^��e�.3�jn�T38E�D�˺A�,[D�ҋ�Q=���@c � � V��D]�5��r@�����G"v����af'7�K�V�p��I��+Z�mt�I�4� )���Ef"�ٶm܂0�9�������8f�j�{e&��^6P���;\\���h���s�W썢�����Y�)ktbY�H��9�}��FR��{���n}#�f�s�d6�wRB ��<�����9 ����V�8����p�,x����A���Rx6�� �D�F�L��7k=�Q��K�sٔ@�+�7hTC��;J�9��s�%�8�`S#����&�/o|T�0v(�7U��vE�r��!�`�M�)����22���a.�_���n|²`Ic<B� u%���d�����e~M ���s�X����K�����cYȘPR������us'�bz�#Q�e�TƜ�%�#��3g�����8��K��h�%�%��)��mm��Vs�@���p��@	�,�EM0���$��1WF!)���"s���e������ވ�/�ђt����>g�۰�oߎi��*���9.Vk�=$�&���P&RWÍIil�'��Q���u����b�^�e�q����G��`�{��4@~Q"�1���N�-e�V�L�q`��C�^�0��R�ӾN�(��$%�4�$r�"�����Ӷ^N����>x���y`�>8Y�"�h%&�-���!�8��RY��
���i��[�p����T>��$=Hܰ�8~�u����Ռ�L���SpԊ(���XU��j�^-5̤%zgr�St�.�&��Ú?�
&�{��������Y&e<#��Γ�c��8r���j�>�ץ@�.��C���6� �-�' �{蹛�{o��$R
=���jM��~�|���^o��_�q��?�X~�'�T�͸�!�˗��C;J���)�Ug�N�#4Y:�C��Fg<>��1���j0�4��p�������U m,{@��4�.-�D����al�$���j9�X��IkL*
6G$�T���iZ���-�$!Ox�4�PP���Y�,(	�pB��J �6��$�p��ݰ,F���u"�1 ������H�/�喒Djv��=|t�<����+� |4fk�G�D�cc�/�u`Y�a���F�N˽� �}���I�c�ʸɠo�[]��`@0�7���$�F�����&�j��p�A G5��U$�X�~	L��c�8�k�Wb>R©;OM�w
N̘�m�"��X�,}wN���(��3d���8&��8VH]�
������[��#�4�1	]C�Зܼ�4��NƱ2w�`Pc��� ��ۼ�{����0�^���c���뾘ɼ�|�oi�	>C��Avr/j�f��D�ڒ��Hj�e}�MN���X�f�V�E�-��6�e3�:��1�ב����4�7�8���:�����?�gcC�t#ԷPߤiQ��uS�
J��2n[i�]��K0���}.���,?����sp9(>��lffs	d��惱;��q�1�`���Zy�屨�ei��C����6ׇG��� (�i�f{�=Yp=d��^�0��<�͚�F0C�c�X��ԩ��tF��Q�	Q���������2�#�R��NHw�26
�_�ܝ�#@�z
���J���4&�=���g�Z�ϐ�j�i�Ä���}1�Ogm�sz��\)� d�%�,�6�4�F���Yɖ��V�ʊ��xY���dZȺ���3z:�aW�X��f�n��ϱ�Z�������R9$����Z'5���30�?���J��8�5q���������o����#e6*�њ	F%���%���M,;l2 a�x�Yu�767)����9�A?���@$"�$�)�7�;Ϸ�kT;�Z�$�e�x�� ��3���b��<I0pP1� >��!)yb���c��F|�4�7��d}�0�'��M�A�z����Q�4~v �����hbՀ���mnnw��%1�!q�} �w�����KZ/@H���ߛ7�hV����ƥ�t �c��c9�n�M���QM]���C �� R��g�s=�t��2k�r���> 4�^�XTE�'=>�&�@���]j�ź����P9�����*��� #e��82�[v�3H�ɘ*?Xך�[Hr@��@�n�X8::tGo�HR �`�ݶ Xײ������5�a�m#�(I��ˌm q����t+�[k���'��N<s�'�wz������k��}�?�2�V��Hw���:�!i���,ߞ6å9v��*\Š`�|��$��w�o[���M�H��xD>D�g�*�&D�F����l@�f�Ǐ����uW��ꀓJ�� �"��Q�J�Z�^�g��r{)�8�<�mz^[��s(@e��@�Xg{��$��I��쁒��$����S������l�S-�����*&�̡<0�:4�?��\o��p��6M|�@cY�J���1�N(t�[G��g+���jhY
�Qr�xr�F�f�L?;d����d��c�h���3n������f��&��5L�m�n��E� ���`�m��ׅ��aq.I;Jg&vzh{\"�Z�S�_���Be1��Y-ќ�����#'\^����� ���Bd�+3'�Og=&>?3)'��ّ�E��{��>X
�������u�_<W��\��x�J���ltn�)�#�[wzvS�M+k���R'3a����°,�����淓nԧ����VR�����Ŋ���1KP��Q���F�����O
�kcc��Я ���h�+�G�l����dP��JoоU̠����k��&U5Zҍ���:��Thٹ7�x��{�u����:ʦA?���v#���m_�u���
��+؋+̾z�ՠ�p���	I��q�+���q\���
��=N�aŌ��8N�4��=]e�
J�=99힛s�z	o�k��ǡ�u��$g1�J8|��� Ai��N6����$��X[`�`��s	�b����A��xn�A(�[`	�"�M�	�+���!mi��W\��X�|<3���A��_ �CW����6k;W�gQgM�t���,�����qmwgύްQ�f_"�z�����H*
hU¬�}ei=m^�}�q������$��08�[�;Pe��Hi���JZQ��z�����Ȃ,'s)������v��ѻ��C���,������{c��Y�q��+Y���5�C��
ɸF�S�������UjV����C��"O�+�R��TV�qUqyz�}*��d�r����Q���cކ���*�嫔Dd?�9�U&�XO�W_��}W��3��C�8�bk=W3Gs�tc#&���ט��`�s��pʳC+���.�|�]�af1��悻p�xk�ۂ�!���Xn��U:�����q0̳H�#1�>Q	Q�g�n6J�����f����$����$���,�{�a��	�J��CN����FZN'��,��N�@�i������c/�-�ֺ�|Ƴ�3[p��;4y�K�n�`  ��TQ�{6�/#��E�y ��J�Xl'v� x�ui�5h�~�s~���N[F�h�������8�+�M@���aLx���?��W��'�N��>mWv��Qް%f^��0���f�k������洹�ؼ~��\q�K�rna�Տa�m/�z=����Ӕ�_a��O�&Y�D"H�b����Nǳ��ñblp�
����^�#.j�;�?t����F.f�a��?�SF%�C�܊�9�X���Q���v5�\�:�P ���h�5w�3HD=� w�V-�n�݄�a���1��L�	�2�/���9/IO%��յ�3�(��*}�=^��������7s�] ,�¯��2�M��}㪥�q@��ݽ�g�� �ܘ0��r^����P�X�(���#PwB@��O6AN?x��� 4�9X�Ď��S��5�����j!+� �x���J,�Kn�E,�ш@UH.��u#�>H��f�n���}iP(�KO�9Ok]'},�2B�0$�X&���Z�8nH�����h�u8ocg�����1�ى3���9�~�c�U���t�:�]�@61�IZ`=~��x�z��{sx@����j�푰�ܚMZ5nTٹ�A.\˶j\zn�׸/�|�g$����"Q�:��e�5ˣ�����4��l �p;��S�� �r{����$u�+oW_67<30N��$$�½�slJ�r#�	�?�t�*@������XM�z�1��Y�#���ąm��OA��T���4���s�����3�Z����"�D�d_tW�p���{�D�b/���iȟ�ܜusJM�q#r��j�^����T���s���qw5�dq���U�XL)� }���؉�򥄥��]C~ �:�?�$��g�	�f�������m�{�6o�i.	��>	�7`��Ñ��4�_�|u_�~q_����
?x��!gP&K-�Q&0�t��$�ꚁeb+w3��_�Q7��U�5���F�9)��䆁0�`.1��M% ��W�@�ey�GP���D&����srf���Є�: �/S�P,@�	�gq;�8��{)��|���a��?1�auW�1�c ��h�>W��%6�{)�L�>r&�O��g_�x�潀5���TS�r �x�jb�}��JaE㐃J�$Ty��W`J�f%���V�e6��Κ�
�8�ió!F\b��iؐUI�@p � |�ww2�7j�U	DD ��#(���~�.Ξ��󵙝K�ڗ~�g�1�Zh���~(�\K?�>Im����4�$p2`K�D�K���Ȱ�:9�������H@UQ ���������k�t�5�1x�!�F��׬��H��#�2��L��q�������f���8��n���Sf� X�3���]n��\�y���@Ϣ4Tv"8#%"��L[h����,�p©����BU5�	g@%5*�1����X�X�=XGX����5;�3� �cfc��Ч�����}xt�޾="=e�*���=��A�gGє�� ��8Ǳ�W�0�`����b��C�"�ڦ��� ��c塷�,6��?	�Um��l͠e7.��psc)�=Y�����v^�Q�m��>�8�g�U觀���0��02	��ת�L�����j�i�1��C^� �Ʉ���<���V[�� ���x60V���Q�IS�iⱦC�O�Ks�b�۔l�=4�_��AN�iU�20�Tj� ��<��ab@��:7Ei3�C�z.�b3 FBh@���kn�?����{��%t�=T\Œ�bOژ��O{� �Â�{Ui0��)M��?��L��ߴ��*�q�n�5�#�o��Ts&t��AI8|߾�к��FAJ���uB,\�K��T�tڊ���lsx�k[EQvY�e&�n��1|X0��hB@���`�ɼ (��G�/��Tt�d`hӹ	z��]�R�<�e�˸I@�2���@�h{��]5��������j9�E6��2�-�����s����{$��~x�w����j9�������uL�"#�fi`@T̈����e�5��U͠BuFYo�T�4�1i�7���ky�(̩�g5MZ%��3��P⼮�!�ؑt�'�FѢ>�����	ٜ���Տ��������HSh8����$ή�H���:����g(@!�ȋ#��$�N��P�����-p�xvvJT0c�x��@U.[�=L �m*�l�Āe�b��&l$��@ Wa$�6��W4�r���;>=�v'�
f4�5����#���w������1�;e�THÍ���v/�	2�~�؁��ڴ�,�}"� �6Lr �߾}#p�I���;�t��Њ��"��k`�%'�+S�'P�Ъwq-A��F�\8ƙ�T�$�]|���q�8~\ ��*P�L���D^蜎 551��]�%7��}_lE�)��>��l�0t�d�il������5MVS�t�wqYe*c�A@`0��a�bV�'�$Y�uϦL��&��S��P"lq� ��-\�
���*����Q�$i��l��5���Ɲ����s��&\�J��IªR`9I��|P��s5Sq�C�nk�%rH�^p�^�"���qcB�i�fζ2��apgʫ��� �m��ןVFRM?#)��W`��"I~̽4?K�[��Q�5�tŞ�Y�����μ6HYX*��&����D��38�WQ�m&�RAv�G��%@TAI	�1��	�zu��ߙ�����80-�
�H�������̒���^
b������ �m�����nu!%��gbj�C�望>Ӛxp������Je��:��:�YVv��3������Y�F����%g��0N��h�v8�X6��߁C s�b��^jH@�܊�I*�n%a�ɴ�N#� JvVh�Jc�-;ki>$p��0���r�v[3����&R���Y|h+�9(nx�,�%����fh�ģצj\��Z��t�Oq�2��l^�@��㨧���j�v>6A�΋�ٺ��c�߰dK��Q6 ;0�P�Ơ!?/V
#�3�s��v�W=��$��7�VA�c�A��?�lm�g�#(J1��$��g���Gһ���3�&���|I�xӰ^2��_f��(�Hv|��/aqD}�������{��BS9h=z���wlX�-�q� ����H��>������#����Q`�zѝF�C��X?�������q�޽{Ole�c_Z��EF�%..ɷ���#�:�l g���X�GH.d߽{���	��Ew���d������������������|r�͝|?��r��XSo��v�!1E�&�1�G�������`��1.�#Y��h?VV"L�'C������4s��3�&4���Ƌͭ�!��}���>0�>~��>|�@��X�k�� �G"=���D;u_�|���(��Kl��ֵ3ىR2�o�H�i&R�|�b��t��U�����74�:+��Rmh�o���d%I�6���{��I���l�<rF��,u-U�u�>sj����#�<�x@�����}�ERf=2��(*�
�5m��~Hn�gBĤ�$�C�������wR��,�گ&/�D�3N
���R�A
ׂyҖC�뗯_Hw)�R	���P#�Vw��Y<p`�"��?�{¤�t�8܀�������}���&S.��� 4᠒)gk�nB�4��8c���<��dI ���5������ia�G;��{ʶ
��d��]���d�}û|��l��E0� 1�e[�5D:]�=�3z�qn��)� �W��P./���NF:�e@+V�5�6�e��,��i\ױ+Dvs3�U�)��ф
 �l�Y���ߓ�(:�S98� `(a�������f�X	�?�1 ��' �t�ij��	�:�
N7��]������(;�Abk�����*�V������*���ֵ������Y\'�p �9ې����m A����$5p��M"�m��{�M+�NO�_���,���.`a��S��Ć/$w 6-��7�o�A��%�pw�w���?��?��P(�� � �FG&���5�1�(���D��xv�E[���)5���q��!$�R@�r7.�^#�s;p�k\����� �@b��@'HM�X>~��~��W�����  ��W��~F@�97#�y������_~�ƽ��Ƒ�s؍/�B�����1��ٌ�!RA�n�N��D�N���R����� ��}��j��;�sC�Ki�xv���+�ՆF�Iw�����_>QR�a,�|����)*"t��٭��wĤV"J���u^�瘎K}J������qs���D�I[Ľx.:yy�������3&I�ͯ�s��b�/�E��`�+HP	c�[�\=�4�Q}�u�Y?�� �E�|�4�����t4gr��7ݒ��3�1����1�����(�K�#�X<�(ľa�:��G��s7o&����.��̕1�)I�.U-T������I�-�8��M��TB�	)��綱�Yna.��M	����0Y}h��Fb�*¤��f_@]aϊ=��y+ˋx�	0��$������� ���bm�+u�L���� uj�i�R�A�LJkX;N>4�H�b:� CKp�]͚S(q��b�X�	���g19�.v�Mǭ�r��`ҝy�ݲhh�g>M�`l姛��~j`l��0�8��yV*d�����P���˴h`��˹�NA����Ũ��	9�(�~-��53UT_�X>���ǰ0�W(#S�b�ڔ���R�ڲܒ�9e�by(�aϦc��|���	5�:xs�~[�L��t��(.��&�늂1$g�Q#Zjdq-N�4�2Nb�ʥ��?�:�	��ޅ����?�'?���>	:Vˆji������l� �l�^=Y��yڪW���yή�?�{�	-�7k�\|�:"pR+���� .H��X��\�}Š� Ǜ$�0&�2`���  y���;<:��k=�& � t�߾ 0�]��3�����@q�Y�WW���WQ�oW����}~��=cH.9��;��m��p�:<����B���2@�����/��_~����t�(��	��3K{*��*�yCl�?��LaOͷ�?������]Jb!	��	<�[���z��g\O �2��f,Ư����`���2�ONb����2�������-i<��LW�J���,���w`�u�
�:��J�5ҋ�g�PͲ�چ��ܜn8��A���.6���[</zoQ�%�*��H� N�?�'@�Jxp#`nv��*}(��$�(�a��$��1���؃di�Ϧ��L��h��l¼�,Eզ����ma\D��1�N���c�D;%!�sɉ%e&����A�bŞ��i\d]D����&B`�,�n���3��0I
C0���A'c/;74���ju}�bbjN|��(�/�8�W+�kS��s$ w?77x|���oi�1�<ĚC�Gs�n��W����p`ys��H��e-9�����cL����HJ���W�f^���$�3��+)!�5M�TSYR<��HÍ��D:ݓ��pӒ�t��pQ�*>���r�v׬P�\6�;�kc�0�;�ˬn�)o��HK�I2C37�s9�D�p��=�/�IPؽ�� K�-y(+���e�`0��Pt���l?��b���`)��9'0O�nj�q��X�b�~��s4m��g�t�'�>�F{��a��?��ñnlE"���?�� �+�PtM�����8[�us�O��vs��S�o�q�=��t��V�h�;§��z$�Q0��u��I�2��lC���^%0�}UUn��}i]�[�\��ޝ0l����Z����=�<!��*��zf@���ɱ;���3qg�߁	����/���G%���4��7O��gaW:�K��;%f��`�g����ELS���:zs�����w�ߑ�7���� I4�]�f�n��mom�Ā=;�{��ؽ�B����`�� �Gbƪ��}����0c@ubOK3<��2c n�}�VX����t��$?@���+���� 0E�z�y� Y0��u�z۝g��4�%y��Vwm��� ��
~;~ |i��Mc���/>x�ST�M��j��N�I�z�$��  ��IDAT%$d���y0��G�q>���rԱ)�oBdYS���!%'�9!E-�\^����Ʋ��EO�|�v3�4�%��M�1����*�Ӟ	Q`#���������b���� b�w�O��j6W,�J��-����{>1�!�� 3k����kM�05<��A�
���Hv���es��R�Y\U���σ�X�R4U�w�,��ʈ Z�k;Ŋ=QNe��s7\}xHI\$�!w�U4��I�����5�(U-w�9�|�b;2�Y���H!j��؉�N%q��L��N#֖��&����qHz8�qt~�o��qŞ�����^�4��f�����?4�IWf:u�R�m�8�ΦL$�Qi�D����S�8���&'p2���D���pL��}Ѳ�ٴ�.�W��6{	�Ľ-T}��¤��)W��/�jǍEbEw�;1*z͞�M,j	�$���,�T b�Ųld�Wq���/nq�5uzE��!����v�>���_��֌����\E�����0+V�防��s�q��FR�9Kǩ�ZXw�  �}{Hl@4�`��1gPC-)�֚j�p}O� 	��Tlc��\��ԏ.ػ ���n�(�S��h2�X{c/�Db*f��G ˇ�.#��n�uTtI��&+����	ᤡЊ
Y鶖'po�w�`b�2�4�6�>��P���"�2E�>]�$���a� ���%�_6�`��?ʄU � ��%`��͡������{������B`��uq'�ᆻ��V�4��.�>��t��<����ƃ ��FU
�~��M7~�73��	L�w����s{�z����� N:����|��Ǿ$��\�������t�p�� B��p �I�U����@���<����28�(���a���o�k���{�������3�=ɌȰ�[-�{ZA��_���!��5�
��~��ž�^{��Hd�������5�%�$��d�aC���<���m/c1M\vy�G+��Kov>��z�G��!�M��>~��s1�3�s�6��H�}��h|����`�_o+����p~qN~�o]_�f�,ƨ�����D2�d�6@����H<C2ڲ$}�RbX'��6�P����c�3Wړ���Y��;�J�]�G�ğ�+�9�q�a�l5��~5H�<�
.��
*�,똬ã]G-���&�Um?�E��ϯO�1�C��2X<u[X6LXi\�YXf@��J�Pʈ�C��;]�� �w�I�L>T�c��P��Jk@�[��Z���/~�;���s)�e��W�Sb9�LAs�Rӏ���,���H�9J]�x�Z���ʶ���ݺ��8-9�1���r��/�zU����}7�1�s�5�����AB�E-�>ǬC6XE����w�O�6��0�M�,r6���rho��+V��J�a��e+�:p��8%�s{&�! ��n� �5��U��k��S�/�$4�ȃ��k��H+t�Z�.2�8��y׹�4�P�o6ۧy���;>>!��T�?��l��	)(?ʊa`Y��"h��,�w�8Tv�N�O�hS��<�I�1�ݬ�JsE&)��7�����]��],	Տ�/�{ܶ�i/|>��m��F�c$W6X�BQ�` �*(�R
����7��$ _���	��a� ����i#�5�o�P�!���w�0�ƅK��g9�F,ׁR�*G�%]g4뛈�i<3�J��@�A*Sߧ��$�~*llOl"O��"�E�!G��@�	?�ן�2w��o�:T>C{�,2\���=��伲��k�wHi����s�`Z�۩4 ���!$~ ��Ƹ�{��q~=��Mҗݔc��_	X�r i�a��0Ǥ������ �)�8�}��:ty�������@� �n�׍A��)��&�N����.$]�i��L�L�(���`~k���!k�H��� ���^F�yzͲ��]�65Je�%=xn�s��=7>n�d�������̂�����Δ�\�^�i��e�/�{i��3v��3����=]�OO�y�Ún�cJ�$�֦̥�~���a,�ĕ6�LdD���r:�R�}o�|~lX-~�$�}Y��aið�t�[�_�Q�V�XVm	��ݶ��<;��~�BL(8�̄� ���8�iKNgXS�75�l���i�&hIA#��=�����s��E6`2D�$8��4cA�A��h"K�V�utH�t���3i�o��<�Q�B�K�s��C+�de��o٘|1N��o��KL�0[]��jv�͜��˅Cb:�}����>d�b�)�DA7l��:�{���u�\�̡+V�-{�������>��uF�d>��Ekj���Si�G2�l����.pC��۷R6��O[��� K;�3���f.a�1�L�Q�n6&��l����T:��AX���s%MM��:�i�\�8��$f�8�*��$ ��{�?tI���+�ֱH�(���2PlA����� `�������}��_A,���H�|��_�M���X�tnw"�˺����y���0?�bx��06�AU@L�n�����nH6!�",W0�ԡc��R�JCkm
��e����1��m�ʚ�@���]����鞁����h���s���2�.�PH��Dƚ�����w��)�6��,m��2���~
�)hY{���;4�i������^r&t���<��� i���{~��Dk~�ߤ{�����8g�F�U���0A�'H� ܟ m�5?���q��#�I@�m���D�mȖw����a���_wI�"���	b��.ʾT��D�ؼq �1�
d?��8\�_�>��4Q�<=�bņ,��@Y1[�u������O�S�P�O�:\�U���	��$XT@,��&1�t�wLM/���K���PuO~����i����niHwt�a_be�u%?5ds���V��&�W��%4�v���S
@�L�����m�e0�3j�G��-��zV��<�4�P9LjHU�G01�m@�Qed�t�w͎#��
�*X��g����7�0�c�G���F �XЦ+�*�U>!=���4Pûnp�J���fF�=1��B[P"�2�3����-��z_����f��<�����l?��z��{�v���'��l���YDn��	��_�5٣�$K�`�E�0�cp}��P�X� � �nosl#�FjL��10�a�EB�6��'����"���[�A��
���8�\Ӿ�-�zon."�:o鲐�j�4@3�=T=BJ�J��U�qm��s����x·�I܃Q�B�:z�% ��.u=��:�x� S�� <�x&6DMwz��<�����oc��Jز�ؐ$D�k��q��ϳ��0v�/(��8�C�B�� P_RN��;�]��ub���d�6���/�K� xs�1>�
���F�۱dE����	�i
d;7��$�K>#��U��	��zA�[a�s#oeV-����XtlU���˶;�N#"��ۍ_�Ll��w���ۃ��m�y�{��ҽ����~�ǛZ\UKCy{&�F��ŉ�ѻg%6���mv�ku>w^*�9�q�uE��i��!n?�������H��H"2�\��b/��s"�P�H(!'"Q�*|nk �친^c���Lܟ c��Q����_vN��l�����![�{��}���N���o*�x;g��\s�Vo�g�s҉:�p߿����$}�LgKaY�`+��,b>"�L�*`X������5(#?\��e5�0@/Y^�h�p���4��$`ek>Ƞ��&{Z���3,1�]b �ket��|��W)=>�.�Ic�8w(UȌ	[�~3� 39�<[1��%濫�7�fB��i ��D��T�]ڹY��5dT6:��Iw����X0۱(Q����d�B?+�l-{V���v��;��آMLIK0r�[i {�=cj^��:�=���?�U���s��&7`#���uO-�\/�����حL��.@�X�����r�%;�R�m� Z�i��Ѕ�2��a�LY'��uM�K��k�q.�|l�g�E����ƃL��,���<��d�#�'��*�����Eh�r�q������zkh�Ƅ
�R$摬'�sA)(I3�x$���?7��(m�f���G���O�~��V����8�:+:<�'���$#�t����{"!4DdQ36��>X��Je��c���������K���:K�-;��2�<��=�'�?�>XR����$B�yc�8$t�RvF�e�X��+x����^�}��Ox��D�9Z܆�g8.C)�ذ��w�1�g��ph�r*���oą{Q�u~�Ҕ|\ܴs_�e�쟣b���/Q"ߨ;�tȍ���2Ҥ���M
R߈��gfA�~R{�q�6μ�ŧ)���n��E�}�h�S���6r�mvӒ�Cߊx���,���������$��+�*K�_�R7n����C��������
�L*�d4��|C�I�`NZK���\�I���%F���m��@���X4���_f�Vqu�Q� �q�s)����9��ۧ�c���&ܠ�	 �A8e΁���*�٤vK�:�n���:ϧg0Ȋx~#���n��J �أd�u��gnc�^u�������� \�]!C�A�%�s����Ot�Z�4�f��bŞ�e������=�{}�V104�q��o^u�Ք��ѽ}{g�،$EM�j�0�

C�O�����d��cp� �I*Ocؑ��Ie�|���]�I�B� ��:�(N��KPS��1�9�u�0X���Q�X� з�coL�Lܙᣙ�"���m����f�D��ݒ{��`CZF���4�;�}q������|��,��Pj��ɛ��-���k�{<�n�� �U���i_K�4%�zZL��	��Ĭ�*���͑s:�.�u�CI&�jA}F=b!�d�N��@�K��G�>�����DIKך%6*a���L�V#y�#�e��U^���HF��6��#��?k�{N}�e�cD)�F1�sT���S"�$������g�۷o$K���s�\Y����ٱ���,b�����G�
�ei� ��Zv|�L�ɩǚ,�&�3F�o߿ӱA*S�8�C�[UL���]��]�z����F���иЫ�2�~6[)���r��%ǞV�u&�ն�so���Z�#�_*OΏ�w��ױۮk�l27N*�־E�V�~�\��=�Sŗ���(b�jK���Z�����D0������LX��A#!2{巂�
�Rc '�E'<m�'P	�C�?�m6�8��7�#�Ø
އ6j+ǵ*�L�Y���Nn5����^��a�E�X��(����� ��P�\�T��%y��iF��5�����It�q_�P���R��P�,�����B�ͦ~���-wz����Q=�-�8EWU��:�E�<	�����;�;'|�{v��r\|o��[��tܕ�b�U��"��Ϧ��g�Ԝ�����|55��vdy(��<}Vű��L��l����$9���_��RV��V\*O̾��
��캛C*�!suAA���e\MDkv��Z{�{�Z��Wb����ɗ�3� ���>}�C �Ѹ#DP���_��w|�pɷ����Z�x����0�:�J��7`��_*��00c����� d���{����z�o}v��^�!�i4(�۰�?^�1�U��!mA��Uͯyn�����{�X�mwm�\,�Ϋ>*J�������C��8;;�y���HNg���	��xNܥ  ����J.���I���w�8a�;�5я�E�Kem�����}?���ցu�����d<f��g�X�gf�����<Aަ���ޗ��y��X8vf��M�ZȦ6r�}[H{���l��F������h��}�v{���%�ꬿ�JˤM7�k	YH�Qv��ة��.���~$N�A$'H�!��3�`���y���	+���C�SfN~��51�aC�3�.��`L�1Ш��m,Mj]��sp΍��ՅlYl,K�|=�[�A 2�5�1W*}o�Ddn�� �2F�{�bP��3���F�4J_�G��S9�����or����Ti�R]����w�q~w��
:R�س1o}3�l,{�{+pi��g��9���4 xB2���˳�?����(2u0fQW-�nf�iy��^Ы��� ����ŹӬ�%�xK��^~1�<�bf6�K�T�Ѷ̺ ��&\87��JpXl�Y�[}�\ho_�}w?��]��5���|��Gv�q�v�\�^1_��
�-Zf;��Y��y]wXӊϣ%���O6&�?���:��~F	[T����/4{�4�����t>�l_n>�;��>_ �i\	��|�
��|!��J�Ǳ6�_�|�?~P�>$�U[P�v�z����bŞ���-�5�N���D.���E�Ҙ��6n���ַ{2K�+���7��Br_�J����}5,[ 2M�V�3
2���]��
<2PJ���4�D^[{���Ot��P��Ԏ������%�ݾ���D+k��ZΫ2���\о!��7Ǡ��QgEe'ǳ�O��vgkR9���@kX���0�ެ�����������*VE�7kcSqh�Ͷ*)=UM�*����nS4zb�U�1�p�ī �ekk۵��]w��eb8/�TG�c�x_v�m�\I��� Ŋ����P5Q���U	���i�5��"��i������	�ǐ��~P������5�� �� �6���N�GcnB֍{hT��]�0�4���h����\��$j>G4�b�Dx
�B���{ùgg���"�����8z���D��nY����	�)������s�G���7s����&��O�b�`=���UL�y��h�{uy�~;&9�������o���Gi�;�X�`mʍ���ږ�s|f�Q���,�ָ���D^��O����ߤ��AcY�f���q(��ed(���g��YT��Y��]���WR]����}��>��D������`$wC�'u�E�F���o�q/�SH�֋�e�:�͠qCS�Gt��m�����˝b[y��r|�
��@G��)`� WU+���Ĩ2�R,c9P�>��鈂{d�ueI���4X�YX�
����]�l�e�Ƴ����m�Vư��r��]�l�e���=�f��9끚����|[��N��f8R�`��32秢L=r��kp%�*꼰�7g��͛�3��{F��s��f\-��ނy�{�cY4[u`y��h�667�����Wh�����|!�4�h�d4	�U����Ͻh|�\;���Ф��q�U�X~�Yؼ~��i�����V�M+wq9���2�d�
���l��۷�Hh����Y �b/���~��}�9�:��]�b�V��y��a*��$ V������������B����i�6i�+��{�n���p<I�������S���x�~�ꎿ�r`���@c���ߓδ6�+�r�b�m󴓟��;�~�s��{[����<f��K�'�c0�~��l��-�S�2�ZW���JR�G`�n���ܐEC�& [�U[qv�i9�����L]a,W-��*���d ��&PY�(\b��jsP<���>��v7�<�����w!65R��߽\u���/���0p+z�
+X���e�	�~��Y� ��d��2��ե�	Xf���0V醴�R�� W�R�U5�?��S��ԁ�h8P#j�SQ#Hd�ů���#F�O8� ��-g0Zݯ�"��bŬ=w];��>�z�<IF8���K`��	{GH�}�ã�7.p��D�+���RK0U�H���9�&U"I1U��q�%�_Zi2�^9 ��z?�q� I�县~s�OO	T�]-��@���|'��X�bŊ+�7�� �e�R~���@��tY��?|�j |v��֮Y�`7�T$W
sg�œ�}���C�/`P������ǟ�q��:?B{ l�Ư��*����m�bŊ�h
p��g�=��0&[4<�Xa�95����S�6ށ�g��^Ai&���8n�=�|e�`YWcY��R	:΢�~1��(ub�Z�~E`Y���l�N^��y�ԯI��Kl⠭i�2LUZ�e:t/��٬t3�C���r��t�{'�@E�g��HX˙i馕Qt�r��f�8�֘{{m x��]�^����3٧S�R�
,�#�ϫ��0�q����}�愪�eV��ވ"�9{�X�b?�X"Xp��6%"a�����������u ^���������˘?rM��V�����;i��1t���0Wa��i��~��+_0�ͮf��5�P�۹��23���� �O����q����9$<~������̽���*߷/{�V��bŞ�����~C_z�&��*0k&mmn�O?Q ~��}���I\��n�vH&�O�E�c�E-P���3ԫ&�_		
�X�ƁB��8��%?���������杝m�+�e߿=t{{{��x�b�~�=?\����ym w���Z��s��|��?�=��a�;�c�����#��@��c]�[����}F�4����mnlQL�}�T�i5`�+K�AR�Q�����$�Q9gB�:2s3Kl䤭,Ѫ�������곟U
C�
���x�*KY��>���Dܖ����ڸn{X�3 �J��8s[;m�40�/�J��d�ܜ�1�Ԃa���$E�9�� !_�6e��-[i53����F=1�h�Ngz�=�-nf�2�8{Ş�pY�'�t��Q�Z��#�hR�(P��2*a�Mm���f���y
>���*D�Tb���u^1;�m�(���y��}8��L�@Gj��&��5�%�ܛ�m�n�_��mvA17���E�w�{���\�bŞ����,�oZ�G�b��ҮAH6�1�b�$��ƹH@���� �l�܏���d<�&��4xg�e!��pL볘l�z�N���CVZ}�(^��8�>�� ���p��QK���ǰ������-+����8+�,���_>7,H���^[����N�_K>�O��v�cv�@-��I"��dd]}�+&+)��Amc�����Ԝu�r=&Ҩ�J�r
��]%#p�Rn\&�h �04y9'��m�gX��`L`��-`��l��kb[��n����;�� ���+S�=�Pg������A�s�b���ϗ���}7sb�"�����ל2��$������![����Z9�Ş��8rJL�W6�I�u�wss˽=z뮯�]<���:��͏?q#H` x��Us�*h�*k6��<m�� .���j۹��3��������5����{ �鱅��3��~�������ll��\�_{�`��T,	զsbt��+V�X��g7G���W[�]��1�i��~*����\`pϺ�w���}�� f̳`5Ï ��yz*Pܴ�G������(��8�n��A�v2$=�|����J:÷P�����{���4.��Ŋ���g�;����i���=�no}Y���ݪ�L��߹q�>�{���u��X���Uk��jCsm&i�[�j�rM�E�L�G�@mE)��B:0�cs,y�	�T�����n-;�)�5���� ��T9��S}ϧ�Fo�M�m,?v��ME�WYX1[�Ī�N�jcfr���㙓����z~�ޘ�W(e�5[=|u���`2���ܔ�������e��E/���C5��	�W�azH]��'Z뷂u�s�+���e��r2�Ŋݯ��&mMn�V�3�L[�JU."�N�GG�,���Rr@3�;�v�/ݡk.�mҰ�攆�{g�jQ6��!�<f/>'f��+psc��}������;;;�*�;����Ad:��F����bŊ+V���}PP��=�L,وJ_":E��G#�C+	�&omo�O�>Ѽ�
��߿����A�����reg7�|��4�b�Zbܵv0S��-M�O���~d.�/@� 2U4mL蘰OБ���'���j�>B�_��~�r�Wf�Ȇ�],�����>���k�^��cs��p��b��|N�3��`���?{����Ai�W{�U�J��cg���]����q�6��f�#���=�+k,�F��q~ ����r��� }��ۺx���B����DN��e�Z��E�G��Q�Mp������O���znf�׋�(~ �X5�}�Mٰ���`��䛠t� {��-=|�eڲ�Wy�gv|����l�6�n�0�������K��o�������C�	n~+�^��mH��������օ��	��nM�@���~^�/_��sHY\_w��)IX�f��	}���,V�8��i�LJ�h����1iO&\�K���R�y�[iF�휜|w�����?�i�PP����-���;���K :�ZR*[U�X�bŊ=��5޽���'7��^�� �����P�
0�ѷ�舫�*�ۺ�� ?>�WW�s���.ͽؓV�F�U=Z ��3���Y���u̟�'h2�%���qJ	t4tD�'�k�}w�Χ��	!���3~�m�^�Z��=�3~���2I�D��?G�N�d\3�6 \� ����o)~*�m�mXn��
[UO$_�k}�1�6�� �:b��͊�D�7�����ҏ�ǫ7�s��2]ݩ ;�B�9�g��ۑ<�6��D�+@"I-v�2��h���*��_��7 ҉���H��ȏ�d*�d�4����O��|��  ^�U�ܭl�x�Sz}r�s+ܰ��� �w.x�Լ�uK��d@T�dp�!?G�1�}*���2��bŞ��xA��3�5�:'4w`��$�����o���DK�!6�:���{fAFC�`'A���,�+*�0v��i��{��iM���������������w4���٢�
���礏������Ӿ!�����bŊ+V�gٓ��bl*Sx�^���{��\	F;��8I�������h_^]v��w�d���%x��{ ` �cx@�Vc�s^~�8#?�}qp pd����S���[b`��� �{��H��q/�Y�wŇx��T���n+Vl-#�10�&o%���V]e���c/������ek�
�a[�Ի�0��ߠa#e��Y�pp=��S8��"�c�9Đ�Y�iD�65z�ߨ<�������^�:�?��0`F&�_�4�nG���뿉�9�2^"C�Ԩς��= �,��B�  ��qD�?[$��e7X^f�)N��`�ty7�|G��\6���df?$�`�0d^��[f.�^dk��˂{�Jt0�<�K�_�yXz�l���$ ���ً�cX>m&����W9P�\p�k�+�����sq�=e�[�j�9f��%�!{�a����3���̹��___Q�HzTTڲ~$��f'��,Jn�I��<��3?���1�nE����};��N�w_�~q?�~Hy-�)������T֊�4�	NFc��I�����=�=n8���2��9���$�����X�nO��oH�A���-���c��M��q��SIS_| ������cj|~~N� U����jJ,`���:��*`�H�*$�|��[&�7�������_���Kj������
&���MGG*�}��*��f�Щ�gX|��򓸹��iE�BR���q�̰����`����r͟������+�\�}��Lv�|5�lcl�h�D>e�k�9%Iܲ.q�l���
F�{�,�*��7�k g}�|,L�RO��O�]p���C��׼:��r����_� 4�w%���y�6(;6 ,�wk��e�R-�v�-}^�{T��2���8��O���.J:[!�ԁ�k�c���9_�'\�[�L�|0��0s��m�x^��tA�D3���,oR(�^�,����	�b�p�d>���������O/�F�cl�w�j��݀����.�������_>k��<��*��ޓ	ZrU̾��,��1��+��6���:��P����4�vƻ��/�h����{���R0vvzBl�7��now����Z�I�q�#bB�Wf���QPٌ�����:]i�f��;���������P��@o���k��ޞ�׿�EA��� u�:�yI*:��Y,���G�v���.���}�g��:�t��m�:!(���M?�U]\��6�c�|���n^H�̱�{��?�p��;9�F��_������%�?~���J�J��L��������7�b�!	�[ K`2$: ��$<����J��"��~��8 ��&�M��n<���0���ܺ�$��rh�|��u]��ҳ9�꥛.���`Ey|�3�l�o���%؜�ETg`&g�tIb+Mҥx*[�7Ë�QU��J%�o���"�=��)���W��Z�9��_���+��}��������qT�ȪגǦ2�$0Ê��q���:ӰOv"!�v�'g�^���c�#T`&�^c�S���̷Okh�j��H{�y�y�M�u'���a�0��g$�2�F���v��d�n#�s�7�V�����ͿS��k�^%��n˹Ԩ�U韆��A�����N��`����ݝQ����y�q�{(gݠ�|J	��6��tT⨷Q2�yV#a>��Yu^���.HTmD,��&���x��X�� A+�C�V�^�c�'�bŊ����+�9��_?�����{�����@�/_v��|I��w~~A�����n�������re�ϐ �Z��I���@$��4�e<�5䫠�
s<*�T��,<�R�����%pyL ��w�ܛ7�������G�r�����W��'`xc}4#���I%e�a�'�E�b����`& W�U�*1d�g�Zo���1 �+G)i&������ �i��Ϝ�ZCs�ʳ�!z�tc����6�����ܠ��V3V�
y74r�}������̩*��9�����:�l3���6�������f�|�N��gO���I
�촬ț���@��3+��r����!{��Wς�-����}�jM���q(�}��ܲ�As���� n�%�y����o!,xg-+^A�gi�s�jY ;>UV� ��x��t��ڻ��3
��̦��}yy�..) ��7i�"�ܨ���b&*U�!��C�_�=��?״��.=!�g����	�k�%"PD7��Go�X�J��s�3g�Ŋ�`�AyY���|Lo�ui�&���?�c�5�� �0	*��(	�6�^ecn�qΌa�����f��ފ�1���T�-L�`@+8	,�żN���m��{XFZj2�~���{��;:<�����á%�re�������'Zﾵz��.[���j���K>W2T�bKm/3$L?��7x�T��L�uJb(���z�1�Иǯ�wN�Hv��s
~slD�������q�w�x�2�24�5����S��{h�7a�� �7oc5`�O6�}�-?0�����Uvl�	��	\�E�zV>��+�6|'��ʢ�0�X��g�?�=p�\�$�r2u�3�o�8[W=Y����r\Iq����X� �H_��ig�ZL6����>��������?��??���%p�����7���O��]p�@ͻQ��qF*���c}tP����z��>B�/�펿��htyᶷ�i���@��ǏH�ӧ��b�hD�#	a�F��~~�HY��� +V��Zy*^�?�i��4���ę���8����� mQU��o����$_u=����$�{�� *omm0�,��4��8q]�T���%��U5�����P�2 ���gL������!Y���#�/���	س��(O�϶��[��#�M��J��ɍ{���^��X6b�q��[PI�t�1�����LNe��h)UbB��8�y���{�̢�E�xq>���D�vGu^���S2l��j���S!�WUc"$=�^X�:�\Zq��_,c�+��,)KD��ɞǿyU!?]��}�-�j<�e�d��ϰUn���$vu<{m�˫N��e�,���L�p�5zt�tA?�8[E�z����>Ŋ�$S'�QS��Ǝ�dL]ҙ	|���ŝ����3.'E���+w|�M�F۔٦��X�A
5 �q�K;���0���?3��ÉC���G�c���߾w�@�����ۯ�A��>��RцX^��*g̝��K���Þ�+V�X1W��b=K�;���.s e���`��su�dBr`	�|��O��\���5�C)������c3 e�+F5��2����2�4���e�g<�:M:�(�~��mi�u��P�ͺ�c�{N��ų0M֨�[d~js2��yY�J��sP�s�Mq�(ѣ��q9�L�TDV3�q2c���g���lee/�W%	�V�PbI�F��C���eb��G"MT�ʑ��n��<9J+�#2�}0��z��B`9�4;����D݃4�ĝ\ D��z��S���]l��4���,�n ����Zf�w!�^޴������ˬx���0ߜ������_}�,Z=:qb2�	4��Il�g�R9�2��bO{�{N��O���W�4��
0�P>��e�nw��4������Μw?�O/܏�S
� .k��@Ζ���������X�6��R7y��˻`��L���d<�ǂ`���t��b��|NZ�v |l�?7�?^R(3c��ͯ�~��aʯ*ױ�14�Xr(���"Ёx���7���lv>���n���w�X�����8�I�@f�m�����l��y�6�`#�F�F�'p�= �lw�}��=UY!Qκ���Ir4�m�#�ǥ��+��-�����(Q��Vm*���=���X���	SXߍ!V�T���"����@��>�����ym\�z��a	����V��4F��%k�OX�����{�=�@ȏ����ɹt�z;����\����}������4�K(.��Aa�8�f5�>��g�@Y�i����b����m]&!�V�x�ʓ�\�e���nbz���жuhefw"�*��Czh_q쬙&�n�$�.�{*#�0}`�2�Rf>�]�G��$+��-�����Oi�Q���a���.h���7w�������k��@�N�8�Y?��g�r]qf��A�ϸ��t:��.~�S9��o��J7Ow�����R���u��;hc��Fq.e���-��y�b����̛�[l~�w�}۳a�;��6(���2��#�p������Y�S�E��$�QՄ�W�e�z�ф|� � ����6Y�yҽ�����L|��(� �A�tV3���=��]z��<���VV?2V��b������#�؆�%|5�c��$����hUkL)�r��a'g�	��^�y��ݷ:�e�a�vJ���;�"A*����ѭ�n|�t_�\;C��5��;9�
sok�˂�Wra<��v'
7&�`n�赙Y"��`�b>_.�g��zJoι�'�S7G��DY#�`��;P.7��*����ˆ�W������_A �txM�z�浃��t�R>u��e�:-��&��(x�d�nc����}��<ۊ{@3�u�XJ�M�ϡMFt��X�U��9�n� ���[q��N��ɑ���ú ���AD��b��I݈���w���O;�]P9&�Z�Ln,Q[� {)},V��˶2�=)끕�_�u����}����� ��b��Y��x��5���{{nz}+/\��~r���̦��Ũf `��s�6Ig�|��?sHb��jN�`e������bh'Aa)�n��
�%GX�uC+��I���?V;�&1f"u�	3� L�YV�~'޷q[C���݊�OY]G���B,�h,E�)H;��(1G�N�l��N�UF�]��=�������\��.8�rf!������s����~Å�q������S�`�~���y��R���5o%���d�V��
��{o�ZsN\,�A�&P�6�a�����k�o�O�z���*^�C��r%ٳ*^�`��C�LZ`��� ��<)H�D�}�|�,+� �¥��Ԗ�蒚�� u����I<�x�|���]^��/_��L�3���Iނ��N��	Ϥm(��|L��u'ѐՀ���~��G`2JZ8"c�6\�A�j81��Ŋ+�J-���b�aÉ͘�]x)n�F�\�<X��]��y_ܺ�u��)���ߠ����<���� bH{�:6*G��A&[����А����u��'�ţ*O�s2*q!�vQ��%�r�u�{%�A���K��UBBqŊ4V�=�+Ǯ.�d�Z�4S���&���"U���"�����i�b�}"^0π� '�6���U�E���u�b����n	cٻ3����H1�SP��l��f���op���
�%�ف�����"cl�ef�ݯ6���ȫ �y���N����fԍ�}�H~�Bz$��?�dq�4�ϱǇ���>��-O40�O��zɞIf��� �y��:=����C}��e(� ��-�����F��t_"(R��
������޽�7G4��E����sj���L�G�o�my��<(g%�f�:�#�=������z���R�J�ؘ]�!�c�T��bŊ�x��R���P~ݪ��i�_e��Z"���K)lfa�����Y|ޏ�Q�d��i�IyzO;��k�k�%��!g��k���m7�_�\R�ؓ�~�@q\o$$p-�3bc�2������b�,[6�}TUZ1Qec�I�����Tى{�ȫ�ecL��xu_s�1� Ӵ��s���5�	�����%YBy�P%�x;�v�����Rz�C�M�]��z���Jӂ��e	�3�y��.� ��>J����s����K���-ujd�m�ܼ�Y��.o���z�야����'�{$6zF�w��Ŝ߉�s����^�Łͱ��\��k��� �#��!u1x���.\X�N^����/�068d��u�Z���&]�J��}HQ�T*HUt���loo�f25�iMc�^δ���z�T�*�̤�\�X-ڱN�j�=;1�[�X�b��2����^��e.V������;K>7.����o7�U�B�Z�'x~�E�thU�����%P�oZ���91^�gaFޑ-a/ �@�	�e	��-�r^W�Zl���H^�k�TI������[`,S-yՆ�݅s���﬒b0J
���'�y_�&�{�D����N�dm{�C�
�0��#x�AM�X�Uv�y�A�,�5�������K��7O5<�.�,2Ut�Mւ� �������4�ˌ�ʥ����B4����(����rC��-�T��a��qpy���Ĭ7���-��؆8B>��d�� @�˽p:N8W��bkv�\�^��1��jo*����'�J�)8(pH�6���O;��L~ڤ��Dq��� 3w��y;r�MT�X�b���M��cBJ�,x�[j�A��fjm�We�[5q��j��|�s�b�z�Ãm8��/��4IjR��!�n���֖|V,�;�����Ih�,���=Ű��}��e{旾?�oC�oL-
��b`
"sQ����3��� �2hX�ց޷�������an�^��+���olr�> ˼I�鄖�n^�- ������8���+B�S���PX��s!�gt0�9ع��'��G�'+��z@:��O���q�c�J=�N�FG��پG��}��[����|�3Pطx�2v�2*B�jXn�ܧI@�T��	�:�>���wҗ�ʟ���,��=��A���eְ>>#Pϑ2���K�e�|!�h�^�=X�iZ���z��pJG��N�D��@���:=��{Pf����dm�4��:2��&hޮH1*M1i�.&7��yy�+V�9�c�֋����FVr�	Q�W-���V;;x�:��r�a�@ו�'��k��h��-!q.~Ӊ��~�W4-���7�b����Uq
�أ�57p���ϐ�JZwzQ��K6�����VH2�l�/����r��=fBZ���D�����2$N%i�m��P�޴������%����ll�A��&7H��ߡm�6pϛ�WcK5��+<�j���"�����j�S0�V��@�D�l�����$u�JC�V���4�*{10����s"[9�H�)l灍�.����cצ��cv&���Z��I*�zy��zO0�eT<�P����UCM����s1#��ga`�m������d^ڥ+L�b�ea���5[�rӔ�mN�϶��|L�_��+�?�d��{��"��X�bŞ����,q�A�V�|�|Z�Nz
��u����$#�����Ql�XE�P~�Į�S�[���٩�=�={-ɰ��h4��~��#�3P�޻���{U칛_�]�}�Bl�G�����S�C3�%1�k������e�Ǽe{$���e��(�j��]��:�o���鋭�-j���=H��k+Ja,�<��M��&Ma�*#Y38�~+�;���ΩӒ�i[��l���f�{A��G<ݢ�G��O���	և�n�fM֥UƸ�+M>r�²S�k� w��u�'�;��w`,;G��Z��0��|�j_���X��d��3>F��1��T�R��bŊ+��vp#�'����VY���Op{�`M��OkC���b?����Ta���T��F}���4�K�s"�UgU�!(�\��f~��}.icQ�O*�U��/�<��r��!�c,��m8^���3���	{TK����&n��'����+w��g|�,?�-b_͙�XqҌ��/C%�$n�ʰ��t�>�`X�L1Y�;:�u�����>1��#���g>U��"��1�X�5�.�����^Yv^ �p;��37uV��r-e� 4�TD�ewM��]�$���OC�S�r�bOՒ~X���>��/_����χ�sW�,o��̺�[�ޔy�矰p�>W졙sŊ+�X���ǒ�x���V�X0�*��0�L���%l�kߴ��p~���P�(���KOr(��^B����X�$!�̸�#�ľ���3x1�`�\&�2�xd�T����ޚ�C �sL�J.߫T���\e�ҸEɛ�u$ʔ�I�W��R�Ϟ{~�=`�l�q����.�&9�3z3(�8�-L��v�V�Y��Ӈ,�_�;u������F���f�8ȧ�P�Z'	MI3��>d6��A��� �.��>	(B�#M�T�M�S?���  �^��*�cܿ�����xߑ����s��t��;xߜ4�ODA��{�--����?7m�^k��l�7A����^���bŊ�D�cO=Y���o�u������W�5����q�=Ꞗ=�����Ĝz|{j�`uKL�`^�-�/z�Ж�mg*�cv)���*Gf[�{��ͿC�H�'�'_�B��<&<�q��-IR�b:N�ǿ���p�"J^���CO˞����D��K墈��8��&H(�a�.��v
f�g��ߜ�
�W<�s���v��Y�"�QI�?Fgp@"�����aɎ�g�[���Z�}�Bk��v�ۦ��gS7��>�gI�(q�2���n/_b��.����jηwK�Ł��w�R+�� ���c����(���Ŋ+���.��}'&o�^xx�=<tI�-�\��,�-�t�瓡�e ��CxR�O��cV]���d��q�Mx� ��M�e0!�LPG��f�Y�R�yiF�4d�(yQ �1ƘbO���O�q��["�T���t[[��V&�j��8�i?'���K+v��D`yUt�.4�����JcэN�"i�����Sz[ [�U�eL�~�Ii�n#�����9���V~ӽ�h�f�Ĕ���gRV�
S-6�ӹ\� �׽{���5=�`&���{@Ɯ�Snp m�J���@��v����P�K����cz����7ʕ��?�8Y�zl��`��#٭AewW{BN���%�Is�_�{�w����o�&+�s-��Zi�f�&����qhX��:+��W�ܰ�CՆ�t���䘟8��=���(YЯ�z���]��f�����>N*�I�����c�b]�   �!K������4�r��{��#�޼�r��T�������m��<%CLHa�e^��d`�>�[��F�C]�ܨ��hF ��|%���8i���ٵ��ȿ����E����
�yq�XNd2\��P����ǱửE����W9o��)���g｟$9�t1�,պGb��X���G�3{FҌ�����x���nwq��F�U����C�*�]�]U�tUj�n^�Ե�k����1�22���x��G�˸��|^$-�zȭ|�nH��X.�.C�,��@N�t�~U֠)�.��8:�\#}2m�r����ݍ<u*�����E� c�,�\VB�$Y*�6�xـ�U�X��0�������������N�p�L-��RIiy��������u9�����pO�X�@r4.ul.l�mhJ�=_���X��̷�zE-��Krݢ��OU���ѵ�$����m6��]��^?Y>r�VQa��<��(�B��7���HV��Z��p�o��x���E�q�\-\���(lt(#�LB��С�<�8�ˊ�C"���E���ń@⌟�[��#�=�=']�(�2"o�tc5�dG&Y�Գ*�ie����t����.s}I��(���BdY�����_�,F�t���_�[�\�6�:e,'YR��X�	\i���s��E�����T�\^�W�N%�>/v&�W]�%?r)d�*�yJ�Ű����J�J�D
|����%��}��o�lI�S�?�.�n}��ZjEn��z�-}�E5��c�0�w1�������̠r��B��Q��n;��h���g}X�U����]Uq��p�-%�~w�	h�>)�G�"�.�X����*�����	��>�y��wy�H	�_E������G� �kD��jˋ<�RBt~~.e�y΀����=���l�_���v�1^5�bD���L�֫u/�-�3�����T5VOv\Fs�O��{�+�F�Q��K���
�<��g*˭�J��2m���%e,C��n�%�v�c�-��͘5>�1�ʥ�W�����Cْ��8g�X��*��zP�������{����W�x_�I���촲}�씐!1�O����tXVi���tzQFi�?�~��e�xG�[)�E�A��p�b&}���`�P_�����E��Y`9�8ge'EV7�M���=�d���,�S�;���Q�r���r���Qay�:���8Aځ�R���9�e�~��Rg0�)<��\ȌOΙ}1��R�pM�⬤X8�P�Dw >� ˈ��FCʍ2�ڣ���n��D�uV��pa�M�O N�$u,:1ג��(� 4���pcN��!��edT��[���Y���U�TS����et�SV��H���h�7u�gly��'M�ōT�0�z�g�O��� S7pE�r�+�7j?ϩ�q�<���%�,����nd��\bJm��~|/��|���xY��Ҙ�֒�窚�@����T��Z��<�A��-��<� �ʺLe�Ѩo�g���\���][
�i;W2 �ͦHݶ�����g�6��*��*cY��4$���8����^$ZG s�dv�(m#N���ե(z՘v���%��#��J�����^X�W�b��wnA��mǃV ��;:I��Kc掝.�Dy��==y�ݹ�O���c��0SR��U+E]ũ�ìi𯂔�xTVMZk����'g|���Mb`9�&�0�6�UR�Z�fu�!�v��[��	��
n�UxWK���ո��\�M$��J!2� �8j��$�)އ�b~��6�������Wנ����d�&���t�n=jڧ�_���(�k�#ë%L�A��� ���nw��m�9�W��W��s��6l٦�cP0�}֑��4X�t]�rV��
�^)�AI+e���v \�����<�M%\��R��hTF�u�]�ç��\����z�6�Ɉ[q��E{!�ҦHWݜ���FtA �A���/~<?���Doءv��j8]��<�W�W=�9y��Z����)WMt��HZ���sy��f]nW����a����Ő޾}K�~����/i{{ی�<T&�1\X zڛ9��L,׍0*#�W�d�Xy�*�C�DW�W@]���B�e*���VIZ��rRo�S9_=����2�:��e�;\��^oҗj}/�R��40�,�C�����X��6�'�����z�����*`������������4,�BM:���Lw�����e�U�+�c�Ҫ�O���/�n���͞��9<7�Ɣ����b��
f����0�d�[�����[%��{�]Y�)��(/@}!���p=�ځ�Uz�VБ�a�c���S�o�q�K��A1]�p8��p�٨��ȋ��p��r��_ę�0�#��K���2@P)i�g�T�Ԗ��]b�����Y��׮��#�W���*��z�*Q���'��Nv/ny�<h�H�0<+����s6d'd��*�/���q��@�-LUZir"� ��@�VO&��J4��s�v�\�����9g,��Ï��>�^����q�qarKp�M�����B3 �����Ǎg<����f}P��y�YT~z��3+�w����d��H����ʘ�Y'��(���{$Los��Ȭ���;Fec��@�g����,٦{g�-��׺�]�.۔a�t���Lp`G����Z\��i������&�2^O�e�p�@d1f�b߳�s��,�z5��R��t���jTs��� ɭ�ګ�=[̫�y��	��>m6h�����	t����,|_��	�тo��y\��=ƴ�x�-2��+J�7�MM�f3,U�oq�?��4�@�r��L�����ݪ�d �:��9��4����&��iz��K�������y!k�M1�~s����Z�5�k�����E��G���E�3�T�dX��Z�U�-�}>Y�1�&ia�pf9�r��i���4`�ur��0�>��!�������;trz�:2v�&�u�_��5��Y��Ygggt�]���J�L�5*�e�=W��y�a�ޖ��՗*mU<ct�<�g�W'��Ϙ�/j3c�Q�󨦔9<��޽�1�:�����J��&��$�X��{����vZ�&�4:m�D5͞�,�9��N��]
(���5x��0XnH�IT˔�y�KkӍ�j��p���W�$YIi4���h̬z��<V��u9K�[ǲr�'�.Y`���(|G��ijKb� gY'��=��v۫5����z<��k�j��m �h8��2E�8��t @[J�զH�ȅ�2w��VK`^i>j��Y枓._3)ŷ���G�q�f�WH�0�|cɒ}��{�%_]Iy�̜VT�]�K`3�YN���=l�mp5db��B�y�8��,wQ��I�����bx�A�~*c��Ю����}�p�e��ĉ�EZ_p���vV5+3Ψ�t�,� ��}�`gy��<�u���K�ؤ���q�r�dR�]��yk@CJ�`T~oR�_��ql�Jо�v�Xn�2���r�6��D�q(�^�	j�����uQ��+S�2ӰT�6��&���Jgu�2t�ggU4���n9`��	O�dE��'�0FA$9#��^�HT�u�� ����n�z}�W���e��U~�V��oF�X��Щ�gM��0��D�6���Z��O�q������/h��҈.ϱ?��[��$�Yԇ�ËJ�Ȃk+b�M!�G�2(m��k6��|��@�qa�-7��5�M5��ˁ�hu�F�b�e�-ie%v��7S]&pT	�hΊ\�i ��u�禙f,����h�hss�BsY;��1l����~M�S���N�`(}����?S<(Zy��t��3�JN�{�dپ+�]U�����e�#V�ԋ�g�����e<者c��s�R;�?�N�Ӱ��殃>��UY���![��2a�����v�2����SK\��Β���J����Z_�U��͗���P������M>�^��^Vn�<�G�uj����1Bc��qT<�nBQER�,�B3��jQ\V�t�Y�2Y��~�@0,gyws������(�i_�V$\�* �[]}��%j�����@�h��el\n硁J�ɹ���*J3h�2���ܗ�G��6��0a[������.a�Xg�a[cj̼�e#���L��F�<�s[�ҹV�9��+rXBvA��#)=�2}e�\e\�03��ZM��M��W�r�SGcp}r���2�*�SidkO/�Z6��\�y���zs����9��{�W��X)�ܺ}��ol�v�I�2z����h0�ۦ��&i\E�|+d<gS9�3�׭�X/ϝ����_�����Q�He���GB��n@�N��J�Jigp��ڳM� �:��t.�E��2�%k�nR��`��C>�xkpV��������� C�׼�ʅ�Tj�p+F�v�y}�1q�6�B��1A���ʴ��1 ���1�ۏ]�����)��Uq��,Nڪ�|��T��r��2���K�"s	��i;�C�<GCJ��9زO�$c�1�]�6a�_���`hs������^\vS�RQ�$K(�+�I��}غ-������tP����d�,'���^`���*�U��h�T��Q$�������b0�ta3��cy���+�m��E�����ƒ���k��k�Й��֞�4�p��L>���f��UԤ��`���T�K'{�z����~W�&/�t_�}�n�5��,I�׎���3��}�s���$Y:���4�[��wu5M��Zp.�ʲ!Jr��+�Fݸ�����m�',�Tm�m�E-�V���j}��&1�S� ւ�Ľ�06Q���v��F�?������6�&ɪ�����DHf*���1�"�ȼ�oe�
�o�6���,<q�t3��<.�n�����B=�m�dPbd�7��4�0 Mh�ƀ-aD��T�2�[�Υ���Fؕ��ߋ��,���^ދS��*rkOjt2��L���,�i�O�� K��j26Q�fP˒_���j�R-�;x�O-���7�Į�7~�A���T�rs��U��Z߅ʼ57�wF�=��$I�S�CA�5 Î�|�̫�C�>���\�	/In�$`9��u62`Y������{4�JSV��]ٮ�X��Y��*�Us+���9I*�$iI�2f��d�Rũ��[+͍�ښ�����8�qu&�
9f�sQ�XY����e�W�V�p�Ւ?�4K3���D27`y�u�u�P��-�A<(�rK� N�ASc�Z�
ϵn�OB��%�Kv�J���ު?K��\���-*�}S�q�t������4���xH2WI�r�H2P�o��K�d-3�l�fW�,�,�Uf�K� ��_8{Q�\[�le������bJ{$)�ɢZ'���$>!����ݏ͋&��W��h��`�$����o�Z��o�����C!�n������b_��*f]_��4��[|�n�PNv��ZϗR����꠲�teqU�ؑ�����z�?�,��m�
R�&Y�$`9���U�;�? ���9d�x�
�fh93��5Ts�:���s�^���Ÿ\��4�l�L���N���Ix.BV����R�.q�Ti����e}�I�1i�Z/@�]e{Sf���g��$�!Z)Rm�_��4���ėZ���J܈(�_Q�V@.{�K��I����ތ����������{u%g���������u�|!�e�R�J�t�I=%|T��k�p�,��2�Gu���(0���$I��,�TW��� ���F�-7ﳙ��.g0�,Ŭ�8�Y;���]�K唩���e2�'��Y�[$�����0�=T��j�/�$W�g�M:N��q�h�ȼă��}�
�����ԩV��K�b�P� ����W(��e_���jX��T��ʮ�F��q����.��W�o�������h���>�[s��U]P���$�r����+�B��
E=˫�c^�>Sad�&/�	�ģ��)������Bv�'���BF7P`{v��cFA�P�b>a���F��n��"�8qX�,�˳v���7���Qv_�h�%�J�($�%z���>8�����%3Qc�c�9.�6O�M�4]\��(�����>g��5�2@�$Yq�1U����&�
Q�/D�(�>�ý��p5-=I�^����ޒi������b���K��ެِKv�l4S�d+%�E��+��6B���d�J'�D�8�P2�;�.���eJ�d�$`�&���m�J�mP&Pё�]0�\p�sQ���.�-��%�˞\^tF����񼺲 \�gͷͧ[�����kU����(�<�I�z�pkB�I�N&Ts5�:o�A-�9\�.��:�>%�����;\{SOz��f�" $ LT�Jt�Hۼ�5Q���]���v�di�]X�k�Vd 'I2')�B�ꌘ_9�SfA!����t��Ara]�ϻ�;�:H��T���UY���A�(��̟\��Bܻ�:���ɕ��K�>w��C�q}"�:e.���PL@%۠E�30exs5H���uk�nR�Ր���ȯ����2����1�S-�ț���*�6F��0�i���l@���J�6�����W�r�îT}�rk�p�T��6���1�,W�˶Ѻ_�$I�E�e2�dG7d3�P`�,ǃ�ߎI�S���E���%r�
��tqAT +FT(�#_�b��.���҃˥VXT�\^)�Q�u��z��Jی�eg���^YVyMJ���"k�P(G3֝ןM�_I�,�\
\^e�Q�e}��+4���,nA2���Q�jfo9�f�<~ڮm��h0����\��VL�qS#�����{���0e�yk"�9E��J�4m,�J�dU�}|q\�M3e�=��DɂD\y�1�����N���.SaԷ�h��]�['	XN2F��
�btE!��O��Ya�(6�@e4�+���WX%��	\^))�s�+S�SNW,⑿r��MJ>�c�f�EU~��ױ�2�*�IVK�ಓ��BZ�s���f^o�qH���� �{�Mv<2�z���a���2n�LT��`�}���{N�ۑ�`�BE��t}�*�%��^��ȝJR��K4(U���a��2��ŘUD��ep���*L���H��L!�r��0O޵�jh.�y8Ƙ��k�,(R��_�ɢ�VI��#���l4��dr9�|˭�>�mGq�!I�U��)����}����%^M��3�Ӄ;���}����l[�ͤ�7����o�w:z8<�|���J�ҕ���H���Kf��4��8�Y/��e�9��ʎ����N��9I�6I�r��E�E�t��T!�ͧ�U��Zy�植nF-��K ��꙱�[�|Kd�ׯf�5:��ң�e\)Z�IVI���_zỲ��\�϶�M�\���C=�yMܫ�Q=̛�7�j�J� �<u2<M�wL�t�@T��l�&�Ɨ�$�L1��1�n�ݺM�dJQ�?��ޯP�¯l3�Q	`�����}��X���I�K�Icf�TsU�78xtW����Fa�e�2�iʎ;�ۉ�a���$Z�UE�}~{�z�cYٺ��+'Y%i��WE��)�,���J�ę��Sה��ɘt÷e�rm�d�F�/�V�A���8P2��*]�±2M���̤�1��ͭ�9Q���$SJ �pC��<G��@e�3%��T�}��K�%�If��&�5���>`�| (�h�k������zռ�5�D��dQ��4�<5M�������n�զC��m�5�U�5��f��.^�;7^V��T��E�c��β�:'��S?�1�*+#�n����5���I�e6��x߯z�WM'I�8	�#�F�J�=�@g�i0��
�J�]�T�$�H��� �4�`%��·�	F��r���WhDJ�K��N/%��$I�CԥgҪ�a5ײq�b���b)��β�5w��\I�L�rNg}�MȲk��ѵ��\��L�u�C+t>5�p�~]ْ3�GU�5��P�(<R������r�|��^t�3�����l/�T4n�F�����NvM�$�X����Oj��*���&%�9���r+��z&"�����I_����
��Y��@���)��#�$I����7�Y�"E57êď��R�q��:�x%%��Y߸����i�(W�CX��9�[��2�2��j��̇=)��J���'�J4%Z�V��e �Xĝ��g���D��\����R�d5�<UV&I2Oq�+�&��(�:u; �;�o��y��2r{��$s�����ɣ{T�#�"/�#SY���Փ5��#���ZӑU"��
��5��NJ1�b�=c��ɋX�,��vM/*��w�z��I�ր�
�@�V�u����Է�|���BG��.U�W3��K��$��D�a�� N���A�y��epYո�WԇKr���r1�I��(Y��� -2�G̛�t�B:�en�2K���S��F��J˵5&\�Z���9���-)M��x�˗�J�nҚ]������y-�@��e��2+�fm�3.�o�u��3U4��tq�&��,=O���\n��ў�@-L}��ڶ��N�Q�5o�e�6���|	,������T�=ҵ���$��YM����q>�����$�Z�n�r���@7d��^�ǉ��c�C)9(�_�)��d9d��e���F�e�e�Ȕ;o��Bi�t2��O!���r-�
68��_�j�5���Y��Q� �l���Y��!�c.ۭlR�Ӄ����4� M�3��Jr^Zrq%͋�uԧx� �+���2��m�e)_.s�V����<�ӛ4K�\�!�%?�5GG0o�IPy�!U�jhz��̾�x�`E}��3�g�W8~&"�z*W/�r�쩔)�l����C���\l�1r���I��8�!� ������_hd)#9 s*W���/d[���ZF����I�A\�
j�Ae��yn��uƍE;�\O��1���2�����.2n9�����1�r�lI�Lq���iw�U��T��4��~��f�鶷��z�,��:�*��L��,Ӏcd��H�+\�Y��2Y��p��p�^���S��#�=͈�l/ǵ!���@��Q;�6������Y)�iQ�A�cf�a8G�!o>�M�K�%�sd{T�ېi�вC><[=��|`I�$a��4W��m�_��Ӏ��z}ꛏ���Ɲ�$�DI�r�9�D���0%FAy���"�yp`����y�3U�n�V�$�S���ҽ�vf͐Vm�Ԋ�!�S�I}��$^Ք���U�/5�K���C�J�o�4��n�3�v� 6���Y%�nE2a��}_���UE%������X̵US̩ ��m���Y�e���}|O�����][ʹ�����	��ظۆ��m-�~����)YDc�rsi�d�$I2�ͥ��`�Je�#?Y3�l��hD�~����Ǳ��碯��
�N�$V���Aͮ(���N�:F)u�
ݥ�p��()d0��(t>&*�U�$�,��Z��eGoɥ�'m�q�r�Ĝ�y*%��%9Š��~�I�S$YEU2�n/�6�i���
��
Nܬ[m���z�B>.0c�W둨z����I�(m�T!j��X�ߺ��{����9Z�*��\�/�ߧ	
��O�V�T�p^Q����ݳI���� ��]e�%%�$�t�yC���I�p4b`�A?���oA%?�Km���IZ%�I�$�lJ�������s�4���F\����yI�Y���$=B�%S�M�V }���k��f�:��Ѥ�z*��N���w[}�h�%�fI�C��:�}�d�y�S�2�妵��xш��!��X��^7�O�ٜ�Ɓ?I��IspTW�M��;V&��h8���U�hel�
Y��l�6�c�1�,8]j�5~���uա�i�-ȶ%l�l�H���R�s�����D���[�YI���
���9�,�̔��Ø�f3���J�)ӓ$)K���]�1p\t
�;��:�e�e6^�T/Ҧ̒����A�F� �xZc�_Yb� ��M�f
��NK[����fGO��64 9q�!�a)1�g�iR���m�B�{���6^�Y��f�6�=�S�fl>&�1��LW�O=��{���g�ϗ�JU� ����4&��1�r2�����g�c���(nj��Ӱ�X�6��aim�'��D��-�&^n��{�������Rqi[���*��>��͝�<��$�z��T�A$t�����}f��UYT3�$�)	XN2'Aǌب@�GE�(�N�Q��p]H3��R��AgI�z�l;)�$I�I<�S�d�@e��_��Gq	$=��+F[���֟~_�U԰o]��ȵ�U��l��rIVG�φ��.e�P��Xi��"7�,b�=h�4���ˎ���-|o �ƌ/\���w�Y���N	��{����hD��ŉ�n?��kNg穆1�؀�nA��A�`�\N7��7_�P��h�Oc5SCՓ�V8zd��),�M���=��|���m :F��=�O�U^ġ2��y�/���I�$�V�ߕ2��N����lN�d���$s����Y͔�5f

e�g0wئ)��*
I���Ġr	Hn̖���e-��4ˍ��5/�XV����2f���D�*�`�$��.�9 ಽ�!`���r"W�%;7��ٔ5�2�#�~��e�Z�K�-ȺDE��i�>���B�i�CJ��I���<)zO?��/X:Ǚč�� �ꁒi�
�l��J�t]/F+O%� �u{�.R^!��+m����n�^��ĳ��x����t�ee�F����V\�T�a�^�(����B�h��4f�9�� ?�6�$���Xh;l��шA卍M���J6@�+H��,H��3�;6�[.�\�u���/׍&U�$I�DJ��*M�������6����P�ѲA.��e�@�UEv�⫢��� �צ�2�ĠɳU�/7�K�N�C*(��;����xSKs8�2��3��%�^�h�j�$�$�T����1�����	�$���)���/����!�Ļ)�
��k�j@���[�w�l�:܎��V(���v��xv ��lZHI;8Sݶ
��3�����X��#���¼ HG u\I���U��RY�= �ox�h��������޾uH��6H����f%D�# ����	\NrEI�r��5>T�:�.u�a���ꐯ
gpY88�y4j�N,�=����$I�L!U�E��<~�q%��D�T��8T�`e�	&�^���]��X���|
P�ҩ(�4V]�V�(�t���[q�՞8�k���<�Y��I"���a?[E�"�BVb�?!s�]�`�U�E�+�Ϫӣ`Jt-$�9��G�S�GC�>�GI�)V�8L����r�`�D��i*����;f]d�e.���I��x��M��2��FX�|���P������3��(������i�on~�,}8�0˝Y�X�ј�t$9�(̲��0���1Y��6����(��EO��R���z��z�cD�1�i:@�<qsu0��f3�����uFN�8]gFS>ou�&U�*r1	�۝V��,8�T[�[)͠�O�a�e��H�J�#:�by��Cl�l�U&Y�I.#	XN� 	fg$���1c����ed1+[�e+>gX5mo��'I��R��4IT3��)A�Tƈ�C���_@���ց亯o��ȴ�Cj���)$��ks5�2z�u���S��ᛮW�j�c��L�5��M-+o2��<у�E��[�����G�ܷ,|��ᨻ��X�߳�J�g��_m�.t�܋�*�p>v�"�z�﹮}����RrR�)E��T�t�@�B�sټ�=5MU!C�4�ո�\,I�/a�/wJe%`P���LE:Ɂ�F��FgC:������0�N4�h8���9�����鉙�{�GC��pÐ�9�������b� �777��ta�sJ�''�F[�����R�ߣ�`@�[[<mcc`�����c��u{=�4��]Ǿ>���>�gᛩ#(g�e��]6 Ғ�m��KZ΃��E��qV�k�ئl"��lM���=�$�
In��k� 2s���^���9�)��$W�,'Y��і����Dy	i<�i.�,\�dk���� Hr�J� �&���X�F����%.]oj�Ӛ�L�m*΁�L�����x�SV��L7U|ٛ�e
��)�G����<�:�'ݙd��@�]&�)/*k4��J��-��>�1"��]֐W� 	��F������dW"�,���/>�σ��)�9*2��oC@*�\d�u�bL��L����nڸ��*Ku�F��f%��x�ݽC�A�L1X<�߳�S::<�ׯ_Ӌ��������[:;3�ۜY�姿<�e ,?������/�h{{�>xH''�Ԃ��&��t��]����1���`�r��Ç�q�4�w���a��O � �GƟ�pt����������Ӟ�������e�����G�����s�ǁ���� ���5q��UV��q಻I��b��R�1EǔW�i�'I��,.yo��A}�i���/�����$U���,gِ#�,�:x�rv�ĘȬj+l�gu��	m��x�%I��,.���U'�����mX5��9�w�k�g�, .-�^��@ႁ������VUF��#�ڗ�{��K=�vq���u�8���L 8b��L)i����Q��Sxg�)�|f����S��;+I6s9��r�	�\���^��Aɏ��C���,�t�l	^K�d։KĻlg`x9cP@ 9'�gtxxL#�F(Sϥl��0�¥�ϓ
,��ml�~Fy�ݯd;ʴw`�r�2
{�>��].e�R�O˲8���\�Kl(��Eɢ�>��Qi���s
CSTM�@���&%�dARy?��ї؞���k��� ]	�8{#�2���[��������\\��쌞>}A'''ttt@�_��w��1������{����o����1�Ϸ���'�p�RGf[/̶N���3]�������ˍ�"u��'f�Cnl�c;::cp�ި����#4��0ۿO�>zD[�[L��c|��-�|QЩ9n��1nmm�Ǐ>�up��Y{�{t��]ڿs�>�O>`{�cu���mz0�D�(��Q�� �m�'�E���Φіb��K�a�I*��\Ϫ�pm�Sx'I��2��������O"�m�cEhn����s��r��̺�n�^��νYԘy3�:II��d�"
H8�r�������q�0P3e�&�����*2j�o�I{�U�$IT��в�{1O�BU�+@rp�,e���9PH9P�6��M[��0�˲#E�r�!Iy@�$�aXp�N9�F�,�e��0��4��d��SDg^�q��'�����8dA����_L�T�2���9A���k��,^.�V-��ǓV)�̕��.�1�i\� D@��Gi:��/������磔@�hXЅ��t����2��kp�nq�<�s�4 � s����u����[���I��;z�7��
���H�*��e��s�[����Ƃ7�A��.$���A�!dڒ`�U���Me�$�2.=K�1���,[2bP�SV���H	[�>�-Y�2��4��A=� s������7o�������;z��=�|��L{G��<N����8�ӓ��nn�5�C��������:�87���1͔��A�һ�ڬ{JC3�),�Q���c0��m�$05t80��է��m�%'�NO��q��::����������*�QΙ͛�����Ǐ�/>��Ƞ��ߧ��3΀�Z����ձp�2[]���1�;.��3ru����$2O����NZKl e�	�O�1�-��$7!cB�5�4���ݤ�/e��I3�Cu���o�d�qW4�8Y�LW�Pn�޸D�Z޹J2N���Z���Qd���}��d*&#k ��I�$��f����q��)��
(��u��%���8gl�H�P�B�!g��l��*�<d1[ ���e�PrN-�	'o���.�/?��գe]�����zb�9$�B�uee�	� �Qf�������_�B�:5;a�{$��
%YF)W'��-�#%�����1�\��:M�E�3�)xI��O�Ç�$���GG̴��Ç#�LD�*7.-E�6���H�u��q�t��-؆�aΎ>;�y k�M�$��]p�f������D�£��������G;;�f�M�Of��(�4..��zF�|��g=w�.�EЕ�Jw��<*l�B��$I��:�`S�}E�t��J��ΊA�,L���A�kL���kp�*������������~~�3=y��x��>��*�ȹ���ca_@��f��+f�y��U?��#�A?���'O��u|e��`��m��# �������赗/^qP6���󌅡/ ���w�z����)g,?��#�~�_~yJ�?��~�����_��_�>�Y�~�٧�y}���{�σ+9l&����l�/K��a�"{��:d�!���DpY�'jz�&�W}�J�|��5��K1ɲ�${ ��MŕWP��bj�r��U���q-����P�ռ�$5I�r�k���"<rb�IBLf336JT!YH\Ν�W��NزK��I�c� �c^��8�
 Q�H��f�D�s����t�}�ueY�/9�NH�!d����Q���ӑ��������L@8i�:88��<�qv;=�\���8���o�)4�����,ˬ���7��s�K�%k��3�q)��b��X�9�/-���@�@��*w���j�k�2��܀�y91��"�Ѳ|�Q�'���\Gs<����R
���D��#���y>�HY��)r sHx���Ms��
��,��O��Z\���8�Cn3�s�m ��N��o٬p���M��E Lw��Н�w��;̉
���=�3.o���ڵ4B#������C�r���u��?�	�OA�$mg*��C%�Z�R���!8mw��6��-����|..�
Y�iNz���}3VtF�'g���zn�7o���!=y�~~��x��P���@3�h�v ���I����KF�> �ٽ'A��`��^�Ǖ�ׅ���s��k��O���	��`w���v��Uh�Ǯ�9.�Ͽ���:����t��=���z��qx14�b��6���#��=E�p_�Q1������~1�p,'����f�;�F��0O���6�Vݮ�����zEGv��QP^eA�(���>ӹ���v�L���aӥ��n�$�$c��X��]΁����M��T1-W�2�h�:�Q�Ҡ��x;���2]U������e�0v�	dn�,'�6�gq�Na���QMm��⌚$�%�m�E�դ�g�Le�DeM�N�]Wj�dC*��Qq�JXힵqN
���.=7��S:<8bN�w�����wtvv�e�gg'R�N&�tF��Qʉl?d� dz��9�Jj1�����,�P��Rzކq����t����C������nn��7�������li���:���f%\�Nցas�.gQGv
��v�"�=5�q%����jC?;k׌RN�$Ij�`��k�U�BTe�S]Y�2f]	�((8G��� �i֛7�zxxș��4]qƟ�R�HG�.�U������\��&���R6K ���X)��'�W�1R� LOr�;�Lk�m�2���S�l!�<��go�赻���K�?��?��=zD���c�e��k�LN�gI*/X�� �L�`�:ѥ/I�N�#ͥ���P�y-[j��aO"Gy���l��!n<�xE^�V<���Pc���	GG���+����o�+������+z�����|���f�P �b���ޱ4<�wA� p
���#����I�9�Y�|��w��0��Ш>�3�����bdl��9�]����}��Ψot�_|�:���W�����T;/^�d�T���l�W>�h�A2��>��3�B�ͫ��O?0�}R�i짗�~r��^��o~K�|D�{{\u���0[([�(� ��2��y���Z^5�o&W�%=�$�8	Z�UT���}�=&��o��F�<��7���*QI�ɬO�;�sW�S��(�w&�e���)2����1>����W��,z/e�@f�o�^�X����ĕ���3(6d�0 ���DŔ]>.CO�>2o{0)�K����E�fT�g�rn��Fz�v}3�Nזj�����������q�Ыׯ����w�Y�[.Y?>9�ӳ��7������%��1 �����o�NO�>�������XgQ2ztJ���!���舏�W���4�*8z�W[���������;f_�i�l��i��\�LFd�I��P�8�B ��sm����q���d{�d U���g�Bf��Ό���,!�����n)g�i�z��X�Ae�M.������<���>�?}��'��̛,ř��3!��Qt�G�d�W5�A@ū[�
@� ��r[-�dA( P�b���[h��Ît1Ȝs�J��p�>@"��4��������駟2W��wPllrU�:�K�@rF��>�0H�k*��g?:��� J:�v��"����f;L ���MH)� r/�_]:;��{�==��'��o��/O陱^�|F�����N�]��=ʺ�Z�TȻ��\雨���d݄c�`��za'��K5�2�� 0��6g���6988��t8�1�p�@�8���}�1z���}���9&耝�m���A���w�y>��[�[���+�D�px(��}^賓S�߹s�v����㟙"��=���2`C[��Lñ����ߧL���� �p������X~���':$��;��+ā>=n�$I�����?(4`�K�:�w��ؿo����.W�g+1�H���IR�"����`���d��/y*Q1��JAFׇÿ7J/3�U���Bs��シ��t�@�$�I�O��J�)�3�옣�Ҥ�C:C�fƀ���+��˗�i�/����J��]���j簈��AH�@d*��Ho���iM"�;�YB6��(1��8�e�G�ttx��ЫW���;?�8j�D�,�R�^���_�C./�Q�����{c����̲>�<�����8�h��1�C�X'(���G��{:z{L�_��rT��nx��A� ���.���2����{��d ���6���3����ΐ�������̚\���L�Q�a0I�uǋ�x�vԒ�1�� ]^�����qrޒ4��"�x�[�����l
�3����8C���[T0�c�n�uzRF��/���������zyp�7��1���_?��^�?�m�Ӝ�#\��U\�0b����5�Y;,0�q����t|
`k����'C:={gt�+z�B���o>���>6���A��.���?��d��]�-w�ĉ�(Ӑ�Yr��5�Z.���L��5�^Yj���CZE��׏�Tl�*��T������	��	��y���^�8�7��ӳg���?��?OO~��}m ����7�a.s��.
Pke�o�i�sY9�C<B�p'۲���/�msc�1���6B��Y��M|F�զ\%��a>b:�b6߼~�M�w�hg{�+�A.h�f>�$~��pp�@1��wo�r&���R�1�����&��9Rtvڣ#l��S�����Ǐd��g��m��𣏸z���w����.W�������d.����)(׷�/�ς���0'I�$�g�C� 0Ol��ӳS��>2�������aL��glc�/���&���q��c�3-��TV���~K���1��PM��	;X�U^�e����}.��Ir���rG���E.>�ێ9%`9ɵ�S
l<�4::`���@�"xG)d:rgs.7�'L�+��A�dye,>!���VfX�H���bb��d�X�����,���B�S�����鳧"#�~p����o_�損���]� F& ����nw��p����s�\F��:t~ �l��S:9=b'��8F���;w�1���VA{� �5�X/w��p�zFG�1�9=��s?��!�\`\q^��p��`x����Ч�}�Q �hx���}��m������7�*hD`]v��pg��yw���_�X�n�ň�w�9R�
XNN'I��( S]D�9�-�9d>����Zfy��3�g���˗��|�� Cc��=ʿ��
crh�'ɘ ���pl6��N ٍC�w�mr�8 9;���&�K�Qm�j�C?v-�f�d�t&�͎��k0���mm�9���������43���1�y����޾{j��s�?����#[�hggW8Q�Q��K�4����S�Qa9�V�c��񙇀��p�[T���h�\�)K+ފ��Q��W.K��Q�j�TA�z�JI������@�.g�{�����{���o������������nll��^�3�z�>��ާ��}�w,����� ��]�#C���`dp#ь�v����u�B)c]ǣ��'��ۀ`�װ{6Шӂ=��9J���lG�p�h�=��cKABB.z�A�*���.*�p�o�v޾y���Ga>�~�i�޽{A��⣽}�����߿���'�g���3��:;�,�F'}��G@����#���?0�3�::ܟ"�9�ﮗ�L��^�L��ϭ"7��$Ič5��2��	c~���7��
3��O0����AP	1=|�A(�7:��G���?��N�r�.K���4V�O4p��T�vZ��-[�`2j�|u�_7�>'=J0��tB��8�]ֲb`�B��y����C�[ {�3]WI�r��3ֺ6{�n�;+s&Q�rّ�#I�k������f1/��.Ym(��F4��7��f�9}8:�f{\5d��J0���П��'z�
���^�y{� d���/;��l;���%�ơA)�| p���R��P!:g[�1-��C��F�22j��}�7Y�5[�/��VOu����Zْh�#��o�o����[�Е�~�Ox�(�E3.tw�����?0�1\ۢ���L��)�`N�ڢ(��BF�u�'�bPD����$V�K2T!(}�b-߻��c!�=´f|�=d�S�^�~�c�|�AE�vo�7��_�_7���o�z$>�Rjm���*�r��4@����*�v�y��{�������#���C�gf���ޤ��>o�7�qcR�3�(ó�s�GS-��w{�={��iB�0�!�,�{\��y.��0�PB��2���"(I�	��BӬ�K)��}VZT��o̎c�c�E3�ׯ���Ǐ������˾ѧ�l	T��[���|�A������wL�����72~;]-��M��ǁ�c�5�<�O�v���6-lE$�
�0~s ����"��ȵ{����1�R�f,#۰p��NN�G�Uy1Xd��5��������Og�C�`l������{��]�X�v��ۓ�ƂX���R��.�M�9�}c_A� I �o���~����w���淿��>��3�P�I�`\��y�Vyh�т|?	M>�(F�y��!J�*I��8�/��A�A�%�;wP��1�g�;��8�_��g���_���w�0٘
����X���Aj����r����+ԇ܍+`�%��K���y�����VQe|�7P��t��6��i�����f�\O�RB�������$W�˼�]V1"�s�D�5n�W��nO�'�9��v�$I�	��6���ed����A��N2c�_q����K���D�_�p���|��W�׿��8/Ǽ-�x�9��yD��	�|��E�,ec��y� 83�YG���^�.��c�F����p�u
Q�j��:L��{{t�s��86�(۴G2� 8��//;8<5��s>���3�و�R7��������/���ݽ��XW���4��v�P���ϧ��:�Y��f��O���
�ز�4d���=�C)M�g��R5�KA�*�wf��lF��
������=�\ �A9����볩����Q�F�d;J���l��?�C揀�a<8���ؖ�+5Yəp�����)���Y��:	�"<�'94=��8i���;wz^P���]Ɂ]���µEY�����l�}�L�pyk��� �#�hAv�	o4���꽿d�)<
�[?���Tα�zzTv���4�K�e<��q�d<��}:;%:<xGO~~L?��=}��7�˓����sA�<�G��]�٤��ef��0�X	�䶚R�̾#��_���#��t��td�=�3H:�څ=�k�=�앂��tB0ʹ�s�Y �p�n�۳�P��g)s��c	��ײ =� 6@s � �p��  ��،��l�39�_h8�8���Ѡ��f�u�����l�������͛W���z��9}�٧\9��/�V���A<{���#L)寑�q����/�qF%I���	�[�l?�4;�s��ƽ4���>�9���-����iеO�����@@�3�����:�1�zg�f���b\GOa7�W���*�U�o.WeRޯ�-����v������k ��)̨��v`R	XNr��#r��3�z§H�K
�'�u�q��ȲSBI�$��t���9�����z�.��!iTg��o��̙|��3���G6<^�xμ�p��� ���1V��%Y���(=�V�@. 8�Bs�P�� @"���-�Yd<x� +-��:�gCs�p�47�Ӻà;~�q2M��ߜvvߙ}���u5�@ml #HJX����c"Z�f7��Y?��WϘ����_����s��{�����������D�\hD���ͳ ��LM���e2M����7O������-ɭ4���������Ev���ð�ad*on���8p�������=y�3g�`� W9ʰA��2 �(,l�EpbBJ?��i2n�AJ�ˆ� �+�nP�r�Q�]��~p6����b`�}�2i8_��h�me�� \�玫D��e(ñ�Y 	z�UIp����X���A{d=~����\���O?e��#:�T��B�yD�G6S\�/@p������*ɒ��S�[n�2�Le�֕6(�U<(f|�濠����-���g��?�'���N�|�W3;����;|��) V�9^t�Aӓ�o8茱��>���s)���]3��zt��:��:z�.��^O�e KT�`9�������`S�J�,��
p�2`a����t|��{όSp@3�k������>F���)���;f.d �4���vA�~�@�L��k Hϸ)����o�m��=�u����8���b���vv�S���!}��5��?=�����{c�|����y����,c"O�lu���G��L���{W����I�$��⫷H*�X���f�d\�@g$� ����_�͛S�����=���W�䗟9��Ad=�����n�U�S�E��5Y�˅�]E�8P/����xu�%&b����'!�Yt���2� �8\��}4O���o����$W]��L'pt���7t�D��S�l��3
W��-'a����9��,��s�7q��p��,��ً�^wik�Ɏ�k� >d81��`��z���1B^������C���_�x�A��]����oY�	����+��_t�+5�E��5��ئ������m���la���?�����B��)YF=�.��)���`d��1E��=\/D��߿��^�|E��Y�����G�_|��2pMzF_��R]8���Y����78��[`�$Y�.}){��0J�i0�@q��6p&c|C��@����<�d���n�!{Vy��ה-K��.��m�M�k ��6��"W�	�ˊ��$��|��y\9�k���ovD�aw,���,���
���շ|��	ψ�_m�5�{�N�O����8���@�Q��ñ�͜�Fϰ��f�����Zi��Jف�B�~	�=S��I3��L�W�,��˕�e*��b2�+�u�W07�}���������?���F�}�`����|�ٿz�`�L4�u 02�Xz�,��Ǳ s�8V��w�CE� �2�̐3�aOp��|]3��۳v������Qo)�.�1t�	��ܿO��n�E���9�����ϩ����	R�nLʺs�� �`��ނ����q8F� �}sv���
�ݿ�c�8
·9�\P���67�ڂF�2��p�t�1�� (�~`��(�7]8x�$'�-Ǌl�1�Y#��e7~S�+ɲ���imyg��f�v���e�D�
2 ���|s�z4~H���������޽e���3�����A<H�q��F+��Ab`��{��fC|���)�$�!-�m���;�,`Q6����z�t��􄆦�&��e[Y%g��$`y��a�L��7�a�������.F��d �
ʳ ڼ7���-!g�:�.�#�.2̀��B����4 t÷E�G]�5Pѿ�#3�w���LU��P�-M_|S�(4�2�ؠ�=IJd�	�<�?E�=d%�a���2�U0~ �Wr�s3��u��������4S> d�C��
��A���7�{��6���Mݍ�=wr㮳�s`��A$�RV��5���) �Ҁ�O;[;�؇��4����b��:�d����U8��;Jv����@�����sc��p��1@�pF�`��׳�����z��c.�s�og0 �>�N���٨pY����R��5���-;��G�L>
�O��M��k,�U]�s.�ƙaag�k[���s0��qR@��@ � *k�%N�q2�(�;Ɓ�d�����L]�p�|Qu8������O�����9	��my|�K=�C�:P9 5�b��m��)>���hjy�������6r�����n��b����^�AA���L�o��G?�gQ��IV�q�&� u
�)y��8�^~^d7#^`�,�K�'DT�`�3�K����Pq���|���S�/����}��������?џ��7z����	U����`N�������5�&0::J�.َ��V;Ac�x�4�w�]_DTΞ�&Ev�u���������:N_�vD�ٲ�^O�֏)�2�MT�qA�=�u�M:Am10�tB�CS���t���ݣ����dy�MGO(�`s�z����|��;7��4>8�^oDg���9����.��6�<����{���� (��5�0����>��@�������Q\����S5<���9
�'I��2���>��p�:��U+�h���:� ����1�I><�;����]�x��qE �d��9�{��ǻ��U(76q��T)�����hgG��!Y�,����iq��Kz�u8�����"R��OsV�>J��.��TF%����G����n�m>���F� :<5��\��F7�9^/ǿ,��2�V�Wp-N�ȵ�;;�2�U�v��#�m�j�ugŕ@�B ��#�@8F(�D�"�5����ǝտ��kv쐙c�A�	�����P���肝�;$݃��I�\ ���ۣ�?��y��?{Iϟ��g����=z�����P��ҹ:ѱ%aAT8ay^W��� �Q �QTp��� �5F�>�������mHt�G�k�)סMoS���YJG���>�^d�f]�6��|�|�;�px_з�}G�|�_�X�O�|�	��?�+��G�}����əq�mS������	� 8���e���(4+��j��5�RԄ��_�<ޚ��p[pv^���gڟ���ͷ_s×�O��s�e��8FG��
��e�;>I>��	���ǥ�pJ΃	��Y����0��H��w���pnu��d��T?`l�w}H��Vn-�u�Y�\�n9����1L�T:��hJ�j�K�Ct��
�sp4�,�m�~��ʺ7�©��8�/_��_v��G��3�b~�_k�@��tA�1���ZY��8��_7Mx.�V�?c:Ze�ڗ���Q��l����#��b�B���nkkk���f������_�ν~y�،9d���} 1����Ki*���_����S�j'~w3�i�j>�q�J�N/4"�u�E_�g��ƦTK���F�ͪ<�aǡo��W��#���΃��F<�:�L��X��M��1�Y��+���lk��t?0��}ΕOOyJ�����ׯ.t(t���F61�� �ss��n����So߽}��q�8`����4�����R|��ѐY�cnf��(�7v�E��Qg''�Ĝ�W`~���3�d4:�׵}M���7��2 �v�k�ٟK�d�R����T�А���SЬ�ZO��� �Ã�O�*	M�M���_qe��w��o�� 4(��c������UT��)��RCS�L��1�]\@���u6S�fD{�(6Zd~Qߧ��B�Uf�d��CH�Ļkss�ڔ�6f� �e�$`y]��@"�0��yl�j+/Q�.F�$�����Y�a�U)����͠���qI��;�����*��3 ���B�}7e2,�,B�U���7Yw�"`Y'D���M��I�d����b 6��O���~�o����C([G:�,��ˎZ� E�%�0!;wd9����2�����x��2�e�]nH�o���p���y9�|�"�q���+<��X�D�l�����u]�N8P\�5�r�h[��$@K�Q�9!p 	V��{Ұˍt*8
Φ4��]��3��(9��7t�׿������Kt�?;���\Fzp��~��1��7���?���Q���vs6�r�r�`��;�F
�ԝ\�F�q�T�W
��L��g=9wK,j��R�/͋�wo����t�l�XA@
��$����7Gw�tT&�/��|���X��-���^J�Y�KЁ�M��������8P9֝��X�D�Dy}�T����4��_)�&�kBU����fs�g�Z+�.M��`�?�zDY/h:L�e�׍�>E�d,՘ 2FO8"b��ŋ��v;16������l$�@��=��f~.�bG����= 
�
Qt��1��j9V�RW��+�@9O��&�n�'��C���*������.7��`��?����?�������w��o�em�*�c���>o��Z*�dE��P���Ye'�P�ь��=���=X� ����2��J�BzJ���M5�nÍy������kc��֖�.{��;c#nX��az,�W�|���~�^(��F(f�O?>e���#� �#�x�][Ǝ���YzH5�:�Ѳ�(m+1`��y �e�KY���&�ڦ��������g[�lGJ��sc���~���0Sp�����s�����e���c�MU@�L�{
[�A��]��|\�e��̸eǌqT��#�n�����ХN���1D��^L��g�`c��i�hv��d�j|������W��S12e���f��	��$`yiE���-�1�r-휗�޴� *;�(��G6����H:�qP�Y���n���]�aL��������2�����c�Y�d��I���D��4C�$7(q}�!}٭+
�O�y����NM��P'�������?ӟ��':9=c�	e� S0~�T���LyH�9"��m3P#d��  �'g����ѣ��]�򂑲��ŀ.��l
�t�r�I�HӚ��j�`2���'q�@oq��n�".m�:��M.���2S�r��q�2�{�/'	@ya��C��x����+˿��h$xp��Kf/�M�;w9���{O���+>^��}���F��d���K�������-c�IF9�˙���kb�k�%��5*kدsnk���ʶ)C�q�I�H�L��h��n.	���)p�"��!d'?��E1�猃��G�ߪ��t`=�Ѹ�Ggǻ��z�`9��#�7�� �J�ؕ�l%�r��y$#/�`12����b�3� X�Yv�����z�f5
5P�)��;^W
v�͖����s����+?��S��ydp�𐳓޽?��>��}�����A�����1�,M{?�2#M�){/b���I�)M��D�%��aS��m�L�������P�<�Ȣ}��c�ӟ�B���K?��#�.
�������y��F��S�${� z�1�u��T;!@�!������B@b�|on��Yii.[�$�z"���4��͖םy������w`�)f�g����8�P�sꜟ�q�**�j[5��{���K�aO�Dl�C�߽�������^�(�2{f�]ڿ��T#���0�� GC/���A xB*�����:t���Þp ^��2#a���_����������hg{�u�{s `��b~�5�'�%N#�����^J���M����b<E��DG�x��piW.�&����H}�8�x����6&�4����r��2��vkO<ƃ���K�2g*Š�����לITe�3����|e�<�yn5H�uP�i��o���_U&<^���؜�օApvvʆ�@�!)�YG���xh�wXi���xJ�x:lp|�� l�����3���a�bK&M^�N4(�$InR�%}�@���3o�|\!�C��T��]v��

u�],g�ɠ� ���u8pdvw�|3� �5�������,�����|ɜ�kt�	��W-�c�������分3Ȕ~��T:�w�ǂ� �L�s��ň�3��A�H]�?�����r\��6mm���;;wY��b�k(�tr�jsCbѻ�Ga�E�r,��&�u�Wv��!�S����9������ �!�a�,�}x�e��|{H�����w��￤�������{ֱ��ѳ�I9����<4�*�l�2Ǖ�#|Kr�X��~�=`%�3i�U~�O���am��qf��>g����������y�V�2Ld�x�e��fXTT0G�4��Cm�G��P�c ڢc~�<B��A�0J�*�����K����Wʹ��3n@
ԣ��oP���y
��8[��w��L�K3>����,�\Zt"=:���-�yw�ti99M�����f��N��� �ˠ2{��) Q������#n����C{�l6�R�qt(�7&�2���BRU�b]�ZfO��5��$�/����ߪ� �g�QfnT����R���ԥ��=~?����?����?�?��ۯYܿ�#�D�Cva�H,gי瘳���~ ��<��J�I�>K�f� t_��1u�+ lT\��&���ވ�pF���?( ʹsM��uix>�� 9W  X��7g)� �:�U\�L2���X�������=46�����B2�o~��ь��˗��@��٧�Ѓ���T: 7l�������W��Jp�c��۠ͭ�����ad���!g�/c�߶ٕٖ�ŔjxO��?��o�+�ۿ��˿��9�'�X�r~ξ$��Y���qp.9�I�UJ�e?��;�\m�T��ȩ@�����8n<�+�����C3�Wp@�E��>�ȿ�)�+��l��Qm��k�{ɬ�K�&|	�r�p6��Q�f�+�^)co훋|�4u�|�:��\'��ȕU6�#%֣`H�����:��q��l_Wc "6�l$�-_���Ա<`�JFc���l4p7�q@丄3�Ip�N�?�;�q#�L{\��͙�Rn5���U�o����>�2�U@e���`LZ�鐔��ـ%�0�'/c����kz��=~����I���k6걖�~p �d��.����&����-�w�.g��̃~C6�T-l����p<��DaNh��8 SON>��lq`,s��El������Q�"r.��8d*��s�9�m�f����>?8ZȐ��3C.�NN�|G���@Y���]�=�5g"Z0�:7���8�짟~���]���҃�;t�ގ�:�g��{@��W�:|}���;:x�Y�H?��!ݽ��YAx�������$�X�J���]�����&P9e".�8 �~oY�y�*�*92�� uN���˃ $y�3W-�Yn^���J����U�6��2��hx-t����D�l�ą�Y���R Ϣˁ��V��[o�e��+��fȜ��:��|�6;�^u{������XwHR��o�r���c	Q�����_��p�S�g����ۣ�p�wÉ�9�H95z:�R}��UI4B�u:ޡ�s���	L��}��Y��$�&��=kHnZ� �L�H'�>�|\��w����諿������ы�XE@cIS��X	�
W��:}�#
ٲ���~��������	�grYŮ�Ӎd�f]���Y�5��o�#��x�e;��Tg�r`9w�%�Ph�иC�BFy[M.�q�G����T������>N��Ć�ǲa���{��zw9Sc�.��������C��$!te|������I����ٙ�ڥ�D�0۹�����(��n��`���tEu�h�?90yj���>���=��+*ee=��2~�-F٫L>f�喠��u��L�fɢ
&,깓����$��q{�<��-���kӔ�U�:;�K��&�>E���]�t�f�e��W�\���v@q3MF�FH6�?�fYm�&�W�W;P��\G6.�.w��]�g����3�F�BF�� C5�����M�kh8N2	��)�0��H�W��;C���6� ��H82�_�zE�^��;��u�].�V�%���#l��1�@�Ç��J��u9G*����J��$7%���S�8�����*���֩)�-kn,4x���o��#��8s��c��]��5\M��tk�2���34�8��a�ͭM�So����\=��{��#���s�^��wv=����/_��*4��[؂��N�V3����(�竰Y>��4��/�@e�l���� ��Y?g甛��YV�����XR�x���3���qƲ��%�溾{��yhq���m�m�s-wwү~u�����+7��z���������_�������ݽ��YC�k��;:C2��GR�_DF���]Z��`|  ��o��ˆWj��$2	T��z�/SP)�#�Z�L�md����+w?x�Vx��}��v=�HQ��T۪	`	RTP��˘�<��A��*=��cT��)WQP[.a�D\ ��t9�#��� t����ns��s�)���lЯ���<��n��9��,r�����2��X��?�K�8��v�?{o�%�q�	�Gdf�gW��A
 R"����z;CI;;��j��}�0���V�DR�����Y�]Y������Gu5�h4�@ueeFFxx���}f�Y�J6�!��yNLH)�G �wv�\Fvڅ��9�yeeEd�h���=[/<��I`��?��6��z*cY�h�x�����dHT�_��� �<�\f���i���{�ƛo�;��s��ٕ3
�rF��u�Y
������|�)���v��0���n�֭NIu{)��� gx�W���l6��d�dq����DN;�qR��O�W�-�\���Ph�x�'�&�=�����|.��A������{m6,����: lIv z����E~��ܦ���hm}�#�WΜa��c֑"������g�1]Y�m Ï�l�L���{ �]%<�(l\6����H��1N�r�T^#[�7 C��>s�>:�����^~���S.H!�B�vH�͜�|jZ�C2ɇ~l��۷�L-w�דz�e#��$�~�s�.�fܲM7�� x�x��ʒ��Y��;·�%����;�6O߆��2�/��ko�/���α=~�t��w����S����@I��
X��w���U�.��o�Ǡ��cG�u�
�,��\ƽN��R#L�J
^��Y�J���,9�J5 &(�#����)�$�Է�vhmu5l�w9M}�q�Ź�XO2 �H����\l�(�Z��O�&�mH�c�����3
5�RT���p�q�G߾�^�N���C���������A�z���Ƅ)�Q������O>�˟}Ʃ� O���b�<��F�bZԊ�~u�F��/���	��sAf�Y����@��P��ʕH
}M0-GȘ۷�е��9�51-�r {YD�[ ��9��3��sa)6��A�����(	��^���k�6���MM�����{�Ʋi{$|��(�p�Z��s=���\nH����i:��җ_�����-��%Nkm��g���0F���N��}��{��~3<���G��B/��=:w~1�S�,z<����G癲�E͸��@��J��&��h�q�?�vZ��\Ɨ�5:���l�8~�^�F7nܠ��n��.R���ZG
�A����)$�-s^H��+jP1��@)t��\K�}�o@��ˌ'34j���=�����PMN��b��,��ܧ�~�r����@���za����:d(�q�!������}����6��R��W)��M�޹�\�$��Xx���+��
�☶���-�D�,�p�x/�ʯ�f�C��n��e|�D�5{�}m,b������\r�g�l~�u	g�9�Q;s��o����w�gj���Q��0�|W�"�:�-�����]^�d/LѨe�l_K�:D1�TN�~����_��:�ׂAK�)����_ ���)HSS�i��J���>з��(���o�..r�N�,�B�^�Ւ���(��b@��8j��Q��erI
��DA�m5�w��z啗����t���u�6;�Q�Y�O2�$ K�^3��:$�h�Cx=99%�Ï
4d\!�pV����k!m���� � C����n�{>����x��/��:֬���^�2pY%��1�`�ਃ�љ~��c)4n��e�7�Pj��g&X���f}vLT�D�7��
2�X�,s	uʉ��b�r�����i��ȣ� f�*}g���S'��<�Olc`��9�]�*-N(	
��GZ+�r��ݳ�ɳ.�~��:��^��Y7�e�V1%��@N�i��*�H���6Z��A�js���%�?0��!�pnnN����*�(Ƈ�7齃R��~B���<�0�Z04 *sDt�+���#|RY:\I�(y8�$o�����x���Ns�����'�bd���Hei�"D��[Eq>��c�z�
Ƨ>�ƚx� i 
C��p0�A6?;Gg�,���,+���c'Qdgq>�,r(6ʰ���/*!z4Ӛ���k̹�����!�ʒ�D��2�,SR&btb+X���f>Bd��{�t�� 2�W6��bz� NP=��D)	_���Z
�\FE���a���uc�S�$�u"�i��]�A��ާ�W-��DJ}��	����	�鳺z��Vwhw�)L���g���g8*�՜PʒJ�,x}��.(eh���2��הؔ�R���5nOV�ў����S838��)�z���s�>]�r%ȓ{\��	��u,<�i݊W�j[{.�*��rws�q���ݡ~����5U�Q���@�{R���5��K~>���f�,�s����tHTV�0ÕȮ�R�""峂��z��yBk�Y_�~��p��9s����bfK��TBwu��rA��L��
�@����M�;����k��e��jH���=�+��{�6/]�d���	�acc�y��~�-��o�a
,ȏم�Ы� f�#�1�~r���\����$�G���f�fb2Շ:�e�V=��g��D��Z��,��(7�ʦJ��ߊ���Z�~&um='j�f{��	�ƞ�ѓd�xq^G���Ϟګ�t:��﷏�9�B�i&��[��'�
&#� ٱF�4��X���g�#�)9KU��=�<�Bu#���,V���:�%5;�Q���{{L��ӟ��^z�%.l\�G�NL���,i9��ԉ۞��1�i�T�}f����6��6�<�>;*�����πdm�x�Cf�����ɻ]-�J���2Y�8_��Ns����܉�#L}��u�"�W;M��1�<����S4LO�O1?�m;����zxtP[Pm\O����u���M.�A�8%w��P�0h�(7�4OT���tFNa
��]��p5l�?���g��fQ�*w��z��UZYYf�:�A#
��FH��J h1�w�mƠ��p�fE�8�>��9�!u��#B�m�����Q]�DZ���u�X"l��Bt�o�;z��7����i�M�f^-dX���h2�pj�P���T�3���s�|�[[���"}0z�Ͻd�0��\�B�IC�*D�Bv��yow���78�eXa|aI���qTn(���Q�&q�9c�b�y���B���])pS8����0�Z��:N� a�	������dr(�Y4�$��+���Â������A�H����lh��� �/EŀF���E�T/0/��kw���U�F�䓏�.�_��_ҟ���h���0����,�VV������7*2�8���'����ߐJ�\D��(4����vw�/.�g�}�����������k�5#Ƣ�϶���B�=�7�~��4�G\F#������K�N�����9ί�R$�B�I��܉�d���VN�*����j�r��"��LPd����Xt�Z�EI"@�>�{�2\_[�������=G?��O$J@�;�6#��4�[m\��-�ieFi���R~tMM��ߧ�b�c��(~l�d�;�����)�sg�y�����._������H$8~�� �]dE4[�:>�߶i|��Sa�v�xT9�e�J����a��ɉI�&�����m��f��c	 �q���1M�up� ����ɱN����R��j(}�Mi�P��|2�y�hCʰB^�J�P����}^u>��<�v�����@��n`�8�a��Ν[a����evR���Lm�U��5�d���o�͸��������	^�8^��F8�!U��{(]k|���D�75 ɂ0�3�� ߽s�������uX�˿�K���,�`�G��R�M��z�F�`�$,��g�7��mܾ�&sy�-���f�����ˁh�	�as�t��ZZ�b�\�y���*����l��Tj�Y����G��d�[��ծ�e��ۉ�;,��ob�Ka��u|�^��l���
W����[1��
B����}��B�o���Qt��|��ȿ�����"�V#N��`��ܛ��z}}�=�P���r$��7�\�����3�2��1~
�ٚ
�䤦LYz��?^��xHI����N'�l�;�-���)+��ǋ}���p�Ɇ����;Szk�pٵ�n�F���������ʗ_��΅R��SK�0�8rga@���4�A�i��>"�Ϭ�a�x{{�eD�JD�p&㽞 �$OAV@����sJ�L�r4���:_G"���1qST^(TV 5������I�\��`|oo�fg���B�@�I�Y�w�;?D�����PX�B&���s�� X�kMc|��b�w�ʮ���n�X�goS�3dr�9�Q�2�ٜ�(#p9�kNL�i���i6{�m��$����t�ޗ��?�1=����Y���ƞ �B �gd�#��	̫|m��$�"	E0���W8n��E��2��i����.�2�,8'�w����;t��紾��N�V��~R��c�%���e��nTq���^4$n�M�If̘V4d ��T��
<�Ξ#eQ99a��U�)q��1 .�%+7���"��FDA'g�ډ��j����_�Q��q�o)b����r�� �2�+�&�7[%;���<x��?ХK�ҹsg�@�9�8�cR\4٪Y���E���g`3�����q;e�9��ǝB�$%��b�� ��{�Oo��F�;���{���(�¹%����s�s*���BrB�UH�`O��X��ŌL�=u\a�����o��:R�aJ#��~��4�J�Na�����C�5��H9Z����1�l�#�#���S�N�b�#�ms��w�A�Ϡu��Y��!�Bψ��3����P��L�othsk�9����PK�� y�b�f'�iQՎ3T��)�p .0n���e �������Cbq��+p_I�A)�j�0G��+��oݺI���߄���G?�Q�I��2�	6��.u��*n6G7)���2%��<s~Y��B�_�۸}3m��������U/a����2�59�M�{6{K���t]��N�s����~Rd�������a�C����<x��i���w8e�t��;��Ί�����Oݞ"�;,k�qL�կ��5v:�U����fx�%X����(�	0%_RMXd�������҄�}A8��:�9U�h�"6ٙ��3
�'#2`��$�� \ཞ����}�Ξ]TcA���悫#��Ϭ�T�0�z�O�t�1r��͔>��m��	�!9n�6�e���?�;q���To��Q���Gv:�ߦl��0��Wx��-�D���e�j��Ǻm�0�׌�3j*
v�%�! � ��(�	�����a9�"wgW�J��]d1Xv����@�4���A>�&��ǜ���� K�rP�!�Q`���O��f����0�DJ�~KQ�I�*P]ht�QQ���VF ��PCA.�K�K_�t���w�hD�U�M�o��w8����l��|)W���hX�����{����Cߋ`�����ݺyH��᳂��=���5��ߡ��uz��	�~�%c��ڥȕF��8d3�,����R��9I�`_�=���#�aT*dS0�iq��m�r�
��ۇ<��c
sW�V���۴ً���߲�1@���7���g���r�j�ć�=Ї���w�g�t-8���L����rX����`����.{?�SK_���d@A<��8-�(�Ц�V�Ν��ח ߃LE�J�u`�I,s]�����\���������̈�s��j��9��$��E+����(���"ٿ#�r�7��gMT���79Bua~� j�,������Z�>�xǙa��B�����M��b'���>�$������5ؙ�(5[��J��x]��g��mi��F���#�*���S�ق��#%AJ�t��k����8�i]�i�T��ne�3�OUz�y~��cD/w������],�!c.���8�y�''��ت8�Q���`������Ҭ�go:6��\jQO��Y&�JG��\�s�Ԣ�j��u��%έ��k!���RE���O�Ӿ�k��U���q{�ۀԍ�N������d�ѣ���G'�����Mj�)yO���S�����>k�rN%d7���W��]�4Ǜ��}�Q����]Q	�2����_(f:�#kO����S4����O(
t5���������%"���GK<C���--S"��F��*$�E;� 8ҲH��ih<�b0�0sA����lnm�Ұ�|��P��[��y��+�R�>���b�v_�N ˮ�lJ
X
)c�m�{;�7v�!��ߌ'���ۭV�� �C~�����hsc���w�fggx�Yv�ji�FW��a��S.
F�B�	�hyi��+���t�q8;3K��8�� 2	�
���n`x�������(!rR�TwP���5���^LB Z��Q�r� ��1�y:
�������)����9նS�q��!b
�d:��|���\8H#s �3���4��l ���r5�x-�6R#�L�5 '����|� 88�`��A�M23=�����=@�E�<���{W��I��k��F_|	�U�����^����\_
�(�ۙ� `Q���=�u�a��\��T�څ<��!uY���s'J�,@�rk   t�+W��p��<Ag�b�>���t���S�a���?Bū����Wh�9f�G�G��'J�$��f|+:�Ƴ
����*�@�i/��AtYau4���:���<F�������+d�f�\n6<G!.�/�<��ۥ����^ 9j��/1��Z�{:��~G:�j#��m���
��[6�~����F͖'�_�eN���V�T��QB1�|������/�J�������?Gw�8$�4��F�|#֦��R�������O���BAbuBcނ
��LqxȠ*�c)TY��TU/�c�1ȦB�b�2�A��(��8���fBqSdAq�v��r�?��$K�c�9Z����c���R���>�sʢz���FqP��((���[^^dz�j�:�k	�dНf�{���x�߿��Xn5��;����\Z2�v±�\ԯ�q��yg���oʳ@ftJ���s�q�&�����}�?'B@TW�� M��k����2nT̀[���Ph�H?�qy�q�$ʜ\vH&eU[f�Y ����D9V�N=R9�cV��=���:z(j���wr`��>f�%��e�a�>bg{zp�Gޞr`�������7+lN�f��m�K6ϳ�� R�D�uC�-�"	���	C��#����O�6񸹛����<�=)����$G	+\Gi�e@�y���&?Ms������F��(+,#������b�1��Pȥ�z�\���/�Sn�����mܲ憫����x�`�,R/wL����Z��s�@��bX��^@�?�g�~ƀP;�7��y�˺L�X�`8�"U*�����F�>�ʠ� شT(���A��\���A�2"���<� Z��TI ܠ�@�����g���{I,Yetƙ��IңAe��т|p�4.9���������RT��QNU����N/5�#@��VC8��M�m2O$��q�Ai�7���Rf�X��D�A^�q�66���s����کԨ�߇QVQkb�xp`//-��͔G�k���1'���+����������v��D?��ς�8�D�Eh�A��w#ʣ$��q��8?���i�F��)O0�2�%Zq2�1g�f�ݼq�nݾE�nݦ��]N/�5�)��J������r�R�sO� D�<.��YJ�z!��	��Ͼׁ�����*'�.gL�l�@��͈}wZ��S�5�z� W�I0�B]�PK��~k��DQ�ez�"&�jm��SPX��l���*M$����[7o�����l�+f��6�����<��@)���T9����ټHO�(�x�
� ��cY�z������/����i���(cχ ����5����;�^R��u�V�G6�g�f!5b8AH��.P��i�2E#��z	(L��i�-gU9\"�s3�?�=��x���0�ǅւh���?�8Y���CLG�ϡo�h�y�&�j�7�����QkZ��T�Z���1vx-�,x{B�Ƣ� �g�C=6Q.�}V%
G��`�y��qh6� �q�yϰ����˩ɠ��8d��=�(G��<���W=����~<�.Zƹ�#�ݬP�ڊ!CE0���]��?�1���ϳf���+���*���I��� �?�|<��c]ƌ��mܾٖ�Oer]%��x2���5u�@\�Qm�G9"�"��P�L_��Ҥ�ŵr�J��~�g}�Z��cv� _���l�g\�/���Xp63��Kmp�)����S,�e�ln�膊t���)f(T�f)N2��,[�5�9��4>͆�]��{!oL�&��@�kJ
<�����>G����~P�:43u�f�A��i(cإ���hνHfNvu۝�}8�k�O&��Z��S�X��!���F��|7�wD�_K6m-���`���;���M׮^���y��^�B[[[�|�LP̧�ydEI���3�����l���qT�1-�\|gWV�p�=�c#K���*��0>`��ETv�u%j�B�$z���[7or�� �'���>��`��b��������B�'Q�{�;lX"}�+w��C"�K64��`v^�%����&s�69���b��ɠ]Y�Ӯ�<e��hV	�M�dp�8� W��3a,�hnv��;m��B�`$N��%��ל���gV�������1A&�0���~��t��&ݾ�ƻC�g/�ŋ��=�zU}����Z��}��ε�L����b���ӿ.ߧS���5�Tj�n�ˀ ����~��uNQ��lqT�T���N��E���TYj��g���h�tF��.tp��� ��~�j�3�B֕����6����x\�־9�Fp�`3�Ǵ���n�!���=��=�B�sj:��"���ѱOi�ӵ�ꦃ�����K�o�!G@*�E��.���,vX6D�������]�w�>��;{.���zE�K�`��wY�U1� jձ���zÜ"�V�������4l���P�Hy�}8I��;2�Ef�8��2��Q�u��:
�hEf
Ҿ����'�����p6��@+���h\�AQ�.�N�dDZ�XV�Օ�EG{����9|����I (������
-|W��Թ&�Ҍ�c��u�����H@�
�A�b����v*o]�4Z�P�`?���F�#��oq>���1����_�F.cqdKV� ˈ�f�`��.�>�-�F��I�.�# ٰ1~���`�*#Kپ�p"�Y�R]����q H��h�c8бqvٺ���Q�Ψ1z�/���4�y�����8�/��ą���Oq~�]�̕]�j`��zH������ԑ�ɖLjҸ��7�l��3͢�]�q�s��d��'ɞ"�a ��X�Ϲx=��׉ *��6�WeQ���7��~�3�V��i#��k���N�8��F��1+>�,�BR���e,#�t@?�lNnO'V� ��gsM�����0��,������ �|��f^��ɝ8g-rł堰��
�:����٘���gX��G@��TД"J��f��;n���Zf`k]H��C|�OI�[�	6�}M'ź�w�>���o��}Dw��a#�X�x����E�p4����
d d|&�T�"��HX^Zb*��`$���п�� W�9"� �G�3� w6�\,&�]�U"q�̓������"��4*���Qx�骦��j<���$���r��	�j��9��������֛���{�q3��c�:{G�W���T����S �,S��Ё��^'��y������$������>�]�u��~��?�k�V��?�O>������;��o����?&������˼p�*���H�׋ ��	��G�g.����o?��z�����8� K0� a��9u��eZ_[�5�ܜ�n*8󡬧`F���9S�"[��� �v#U��.���
��huPB_/�����b�.��� ���U1z��)i֟�$�|$Df�X�3���ʣ"��;���5�<IA=�Hd�1�ϼ�"��#�����E��Q7	$u��T3B�l0G̗̼����T�����E�
z �/��?�d�����$��ϱ�X����\���HE��q$��#KI����U�ab�I�~�t�6:������Z�iE����A��#��_���;�͑��(��SuK� }`oyTh���p�"�p�	��*"�wSeW諸n�+CZL\ V�1 �x"+ӛCF�� ��lT[�VB,��5�˧�7F ؒZh�Gz���$Nc�lj2(��͠q)�`��k��I��"��L�R�s�<��+-�;����Q���Y�@%E4�_v�p��p�Wܫ�q��X��{�.����Y0���d�}��nx΢�kЂ�V��>�Yܰ���7��gX6w4+̲`G-Ҽ�2��s�y�|��z������?y�E�a��u����bĞ7���6�e�c<! cHy�w ��Y6���'�f!�{�r��(r��P�q}'�g1�$�"_cį��&M&V>Q����C�l�Ǉ}6����jV��yǁ�t&�#X��Ja�{�6i�3�j����}��j��XK�SG� u�Y��`��r/�)i��br�~��sp�":ʹO��X�V݇��KJR��	�H���������tpR�� ̵�Ө��ˎ�}���w�@��Q�� *��Dtx���?�75/|�緶�����\iE�֔�\u�̅��aAm�`^���p��1=3G++g�}�=7Px�H!苁,^�Q�Z����_��(�丫������-�{�>,RLB��$A@�F8Sz"xQק�$E�����O�`8� �� �\���"��l�'lQ����Y��Q������)9����4�W,�꺩E����B�Q1�$�f=o(��d4�W�LH5��EЖ�\\� v�Ν��h�7��o���2������,�P��qDa���{�+M�Q�:�yT�����c�>��"��߯p��2�֥H��j��H7�E�l���۷9b���p1J��o�q�ư���tf��|��^W�!Zp��FǡF�E��S����w.��=�8'Ha�'
���b44U��QP�����M�w�э��o挏�w�s��&��@����H/͞Ӿ���>������RG�z�id@!��9#��E��1��l�,��}�W���C7n\�^x�f���=�
�kGxQ��-�E�\1Ꝃ$Ȫ��]��g�l��r7I��;�V��\?���
C���ӇuP9?�.��L�ܸ}�}��g�ګ���k�������f �x̚2�C�nȐEZ�d�Of�%F9��I&�X�s��S���x�z����Y �M&DQ�����9r:fn
�iAK��0\���z�=.�=�(�\���EY�)��D[��Kv܈�TE9��0����˾d'4d��,�qVn;E�*�j��G�	�ԁ�@=��F���R�<���7d�qC��y����,��0��'�uo�#�[�>�����;�>L��f[�Jo�9�>��_~�%��З^y�e�3�z�_`$��HeB^H�ڃ"�����3i�j����cmiܲ��2~�F͔~�R�^�wrg��ޜ�U���`I�0`{3юU��39�L��{��I��=��>��!�7:�|,R�@ΫB�Ny|���~�a��ȏ��}����6�� C<)�)��m�O�r+�-�ϫ�:
��[ �W����4���>y')b&��n�}��u�x�T���e^d�����5�h��].��,��&�����ɍ�����o}@@���z��v���G���rx���^�B�����7�dC�>x�+/��0|�B9G�0�J��DeT�v|t�T8gV�Хg/�aP�������D(�/����f���˛�D���@to��$=ӗ���E7oަ7o��)؉��oM-S�D�A$1H��R� ���Վ�q���E1��"4� *�S)f53�b�B�����Ҁa�A�XG�6 �ר&�Ͽtq��b�]�z�w�>���1�m.�'�SC�zY��bxF3�z�D9�\�9������R��0g.��[�h{k�����i������w��M�(8�%�S�f���Z�p4���R煯����7�NNԿ�������k�h�$o���)���u�q�]�~��-ҡ��^�s ��[iĊ�<�O}NrP-ݗ�SeS���1`���6�R����v��b�.�1u���ǃ�^R6r���!n@���W� ��������Y˦��yz)���->>F��ivN�ZG6"n��fU������Dڰ�Ȓ	� ��S���E�7� ��&�[�q�<����e~������Y�w��`�Rˍ#H���
��̜�.���}($8pΙ=���0��0���k�C.�y��7�ؾ��.o�V��I�Z��٤�?x�~��_�G~����3�
�{;�u<g)�-���\$#6K/YC� q$�A���eړ"�Z��	�td5 H��?��,;K2t�9�2�S�aк,E�)��W�嘿���Ō�R���Q!�.�����h_�qnPVpa�i-�[��E�!7 1vG ԍv-~�^���P�h�� ���%ь�w�@a�A�����3�p`��Ǭ����Kkk�><Ƹ��
�hbK��=�D�	���v�.�P��H���5>@��чI����>s�"�y�C�A�q���'�ˤSF.'����I��k諵�v4n�Zԫ)�@s�E盾�j�;�^?d�4�l®��f��ΏL�B��(`��d�p_ni����i�1�@�	g������B�c'�CE����qR�"�.�\��\�H��'��?�.~�B��~
��7Y4�6���g���f}�����nqN���
�����=�ő�s���@��[l�!�)Xݮ�f�ToS����[5D(�۸}�-��}��y�)ގ}]Aȁl(�X��t��/闿�w�r�*�4�����1+�l�	��ɧ�W>���)ٞpdbSE������� G�d��wT�W y�5�����ٰX�_ਞ#��=d
��gK��>ݹs�����A�D�������y��J�*sfc�o:�_��N�:�{<"8�p.�Ln������H�3 ���	����a�AfD��(�D$5b��]����Ab),�,��𜗂l�=�Ǣ�d/�bC3^Ok��.�p�n�9�`��<��K/��3I��n�믿�c�C�����/Ly_�~�.�1׫+������ӡ�N��r�����Y�)����iC��QEf�Ԇ��� ����{�]�~�� +ѳV�A�s����"���F�F���ƀ)�P�T�e��~n鉒"�x�pa���	�{ƺhTh*u,Ғ+3������܇X 0��{�ƈ��X���rQ��g--�*\�R<��#�w NX|v%.xV}�Ņ��E��_����w�j(���f���2٬�656a���)�^��+���翡�>��t�s�[^6�L%-𬂸��e�`4��õ��ljr|�J�8 ��4�&����v0����	F�R9��N��7����o�?���_��\�ȌļE=8E�� Y�c�r�%P��]�����łw�B�h�/��0���(�cKR�P˶���L�R�U�:f/�@$�5���4S�,�1�œKI97``lK�Uq�W�Ut �h�oUI���N@�`Gu�ϡ'�0��[k?���zE?�r����������J��Xk4� ؏�h t5.��Z/����>��p�#��8gy@�cu��Y^V ������� �v�H} X����a�_�� >x�KK�A�:�/�������?����<n��c�İ��M$�WF��&�!�]�siWGA��7چ�2&�ǎ�h�$ժ���ˊ���a�4�E!����j_mP�|�h,�"�U*1����e�Go<�1N*�H�]�v/�W�G�*SV�.�%��B���"�B�Q1 m�I��`<����$�,Γğ�͙�H�R���͌<�\������v@/������Z:Q̡� YXX��壣}�:ߦ��|-5����T�۸=I��Xv�����i�v\*;5�WY"S{t��]���O��wߥ�W�1���u$���ͳ�����)�,�|�$�����5�gg9�C�y��n�9�g�H�b��~eSS'8��Ӷ'Zd����" �*�����������wp}�b�$?V�U�#��L��h�Pm��+;N���5>I���),)Uf���-�F4���MOwe<�'���;����hĔ �69�76�:,߻�Ο?�\�bw���cP��i�ɉ9qļχ����Q�f�ή,S���O?�8�W��)����Kg��h�9{���bH[m�8����8��YA��I�bs���=T;��Ac��
52ԁ��V\�lcc�>�� G�ҽ{��SiWi�8;D�:Gf~�����&{��Ź`�\��� -X��$D�A���2X3 ��f� c�1[A�=8�Y�n,h�V���h�h�2 Z�w��4>+��#Oj��GeS�]�~�Ƨj�����8WDx�'�q}�G7v�d��ސ�r��]vRDb����;ʊ!���g�}A&�_]���6�����^z�0�"pZ�J>��Y��ZY�C��狽̭��~���Z0�f�c�M��KL}��t�|�^�����%	���u�lЭ[7���[o�Iw¼��\\�gp(�� Por����w܌4�Zή�cJ��3�ʎ��U��	 �ԗ.y��|����MV�������,J��e����0���go}hJix])]�j
�؀Kh+���31)�6���\kKY��Y���S�DRj/�4�i)�(1֡�������~�	t<8��2{�5PhO�z�.���Uf	���� ^��g�:}��UTZTK �V<�%;�/_��u �[/��ֿ��r���Ki�Q�p����5Y�$�:�M  ��IDATj5À�G���'��A����9�un��zW�����9X�V0���SѺ,-�`�ǲ0,(�-L���r��1}*E������݄�g}s�6�`�x���S>����Aj`���!H�y���a�B�����*C�u�����yu�Os�n˱=���������G.�(r�h�GԽ�k�3
@ ��{��B1����K�U��4-_b�2wo� �j8�ɸ��m�@��*c-0�^�-��9�=������|�u����L��E)�wp��@b�	�$rJ��[XrR|����9:���;Ήc���R\F��0r�����K0~��_�*��F���L7�����1��[;1�-�b%�ʓ�����-�	�2�&;M�X�_�o���)m�vݶp��^��Y��^0r676i!<�!�ApbD|��aIuwœըE�{�t`��}�����̳̊WT���3���q�����.�5"�h����j��۴�d��5�g��q������66������������³D4��˄�| l�?���MNI�9�کK�]��������eX�N�(^煗�@  ������_�Z� _����E�}Օb�P��̝Z0���^������:���~��y�������"Y�1�/�|@���������P�R:��Q)�Z�ʀ�D�{e���S�[wZ�5@B4?�{��y�/�ns�#Pm�U�9��q�m�4s��
�`N��u�((�l��w������R����Qd`>P�c��c �Y�*�\��bj��D�2����CW�]�C̿���g��Y�RD2ȍ�a���E9��'��{�#�]�l���%�#���ތn5��+��t)�p|�������\$s���sA?��(坝�������^�=��tD>qDn#��c���l�U�����aPtZp�w�ӷ2(�I݂�v7�7��~����{��9��V��	 4�8[$c�E�Y"�{�|/���C�{oCe)�co���ڂ��>�uV�8���8kr�?�� M�m�����y�z�=�#"��9,�Фz��x�Q�� d.~ZLk�B�g�KK�Aw��g����A&-.-�����@����m�Dg*���������\�]ɔ@D7 ��5����;+gV��4ƭ��:�Cz"��`��M��ow�=�+ܞ���4�?����լ���$��J��"g<)u�i�i\h�����N���L��:��p�U�y`��)0R�b�d�2�o��})o�r߾�KoN"��T���C����2ˮ���E����q`��i9�ѯ�>���[6_q�&��@�F�a7)�H��\����+�&Z4�2��}���q�'��f�D�K*�I��%;1znݺE_|�%��֛�
�;P�a��h��WO�e�5�u�E���b��ʳQO4�<��zfeY��`�������b3X�]M�Du��d�Na���
�C�u�r8?��a�HJiUc�`�J�N�^S�y���-ϐ�Az:.Y�s*>�.��ič(�K��b;��B��`�"�2$��v�=�ec�!
�ikk���3 ��Rs� �Q��aT���3��" �s/�H����A�����3�|��/��l���>]�~�^{�Uj�_��_ӳ�=ˆ0����J�y#V�΍��e��+U|vq<�2��N�0�7���NDǕEz.�CjK�GO7nޤW�*���t���kh%�F�i�u�=���f�3y�H*��1Z����CQ��|�3 (PT؀v��5G
s�Mu����V)��s
Z����|���e9�H;dh }^�仚�I�X*XVia@�B E��G�n��6/ Y�UR姂~i"F�].t<2@KƤ5�@d)RR|�f{n�x�p��v��䞌2 r,7�XE�!+ح@��O���/hss;�qE/<�-,̇�ԕ���2Q�%��"q^��g��]|sф�ls�?�&r9͛\�y���`�D�	���P�t��d ����o��ަ{w����R,������!���lhEc�Т�k� ��H��R,�#E�O,�4ŻW	��n�J�_=D-s�TW"�E��Q��u�mP��\�R$������I��3�l���=����D�����MNOr��(�R�8�b�=w{g�)��L�<�����j
�Y��p0[v�R�����El��e�x�G���+��5�oq^��g~�fCAu��i4�Q�����sh�5�B�t	�8�\j��çdT�G�Y����
-�q��O~B/���*Ih1*z�� �E�$>i=e����?�a��15��6����7��/[���'���^�hx�eA��z�s�N���Z=�hGQfgE�)	�X�a�s���@6�톬�\�Y^q/;,��\�Zu��'݋鲕Phx�r�q�6����iP��+�{�^���<u?h|����(%�A�"F��
����;c��:�9W�T�t���v����;飁�}���YM�TcǴ ?��S������͛�n��^��<7D�r�^^�Zd�[qZ<��\��sqK�4�Ls̫<�T 3���h�l0���`(n��Ca-#F���F%Ŧ
5F����M�#I����Bkj�l�xύ糡�țɾD� UT~T��k3Hū��&fU�͠��Y��呷��x��B�s�RN�%֕�5g��c�d���B�;�;�x0����v�yN�&��Qh1�S����:43������߹��ܩ��4---���) �W?g�G80.��Oxބ��.@�f�x����|�\��'Af����0�\���4<Ku���_�:�%��0�-h0� ��/�2=�.d��:����u�+�z�0��UL�jj�,���SOp�F���x�k�FY:8��se� *;*��gG��Y��X�1s�ۋ*	Go�}�1`��6�-5&�&8���8�Z�ƅS�2]�QU�h�P�-�ٖ�QPD�׬pa�W����X����Y�����<�#ܳ�)�?����צ>�?�? ~ �������7�g��0FA6N��<�y���B��G�ppvώ�$ͦ�#���Ҁ�%��~�ځu�����@V��˟ћo���I�{g�,��=
N�6S3yj5�ud��J`���8q����`��B�F��Þx�Ja�.����ד���ݸ�,�ώi*��dH��=�^�"�r�4���d����{��d�0��A>�7��)�'�>#�����N�� j���)c8�����R�t
�u.@��o��)"Ms=�3��7|tN��x�N`zj�l�gυU�aI�3���9�@��k�q� ��ׄ��G	�Gע�:���:m]����ɲcWkO#���=I�����*N\NZ̸��ci�> �Ps�w����-��l!��"�Ó�L�~��(<��2q��*���EI��|nȧ>9*�_�f��������F	�8&�
��?��S���ƈ�4��+aL���ˁ1���Z?��د��jt���@1��h4E�3����E8����Ԓ ;a2����Z�?�����.��N���������O?��~����'�~BZ�Ag�*�\��u
��
.�b��
^�J#� �@y�AA��N�>�bsZ0
�x ������%6$z��4���1�c�7� 3��
�@#���b�p~8������C�:Ԓ�Uc���H��p@�H�X5�K)����S/Յ}��fP�p�ai�@c� G��؋J�Z:��1A��G�^�t��#��ܽ�QL�M�4�m>7���.]d@c���dD'�5������Sw�#����5C�����;t��U���z���e�����a��P�8(� |�D�#��uNC��< �L�H ���HqJ�ܸ=��a���c�,�0@�)����a A�����t��}6�A-Q�Yԝ�Jc^�9�qZ��ʠřT~��б�c�Q�h�oy����I��i���*�*��V�3�C�-ؙf��Wr.|Vr�Q)��
����� ��4�8^#k���tP��mDP��!I���3`
rkoye�)��לh��C�����:�l�9�`�AW6�1;�""��!��X���y�G�n�b�O�́�"v��x*þ���n1�N��͛7����ZZ��_���n��AW��]/Ā>a�F��]oi&��O<�Տr
"�&���]�W��}��ʟ���Y91�������7�(����h�g;B}���]��d	��2��}b�r�[���CD �" ZF**s�ps��*fx�oj�.�U�:'���9�}���4m)������ΰ��uwv���%�7@f�<���c]	�2t���Ykp0��S��0��p��DA7��e���cd��@�Q¾.�8�I�v���ݮ8��)�S���RIF�� tk�������1�5�:�S9��w:�P��M��̜����1��[�[AG�4��ۿ���מ���� �&?��M���f.p��<\���fE���҆,/ΒZpRU��f7�u��
��� �� �{l(Eޝ�C�8����(���v�u��\e�3��Fe��>���5�{*��c+ �A�6�㬯
�*#�\��	@.YR4�vI��E�_=����p�l>��jJz�?e�_:��n\�W�hPټW1 �@#��F��r�W���Ӹ��ކ��>�EE�>@e������x������s��'Ζ��#��C���H/���U7��r%2g���ͳa�����1++++Ju!��*�,���D�tϽ]�ad\|�^GR�9JE�9`��`�H�P���*�`�1(��q����@c�Lһ|,�% X��&�u��a���\��Z�J9WK/��8�5�%�V��U�]@��}�%n t�"�Z�O9��`����(G�9�9�sa��[RM��Q��3�733���%ɓS�2?G/��2ݹw��z�nЙ�%~��TՍ�u���ع����/����>�;��qTz3s�}3�#1�E���9:��G��R��mF��MAD���e��
�a.J2�s��_����;�_��T�y���>]�D�Uı�üp�TwP�ZxK��eQ~��Jc@�E�7s�EO{U;Q28�4,ǐ�R7��P�����
Y�iOi}v�w���v~o@ze�^"R�`�_y!9q��� �K� �C�3�A�� ��^.�	��m�P�\0�ً#ܭEYDy��em?�0<<��!�G���ٹ蜳HB�; ���y���X����P�����eZ��J�C�L��B����֞���鸘��C�Lg�,D�����ǿ����^��<O�Ǉlg:�Y.�$ݰ���_Cl=�?�2��}{�N�xe�(�󨖂Xr����>粷L��qo��d��9<���m��魷ަ�?���k��g��'�EvVy%&|V�x�%�����+����н9c�JѩE�v�A��OqT�8^�?c�Gc �Re�d�{8��k��sb1�\�r̂v�T[��)���c�̵Rv2&��"bxg{��[j+�5t3�<��p�2sX�׮]�Z
KA&�	kc	�\���������쵞Fw�3Fw-��(� c��N�q.N�m�p�e��>Wǘ�#��:SS��݁��-�A�^�Q�Я��MӨ_��։d��R������~�);	悬��O��gX�'}���i�̩�ND���]�!|u91�~ƭ�����oy�;����}�}�>�z�s�]jHP�I�^��{7f)&�K4�B��t��}08������'ܐ���Wx̠�qJ��(��b;�(�L1��	��k���ޞB`9� ��Wi�S�9 K���2OI�����t�ΐ�1p��٢��G��&G��j\Jz|}M���~P<��_�eOT-o@���k�z�q����#�C#N�L�F��(��?���z�M�2�qq��J$����G�p1����Xyd؈r��&a���,G%u�g��[\Z�J�pm �H�l�!&[
�3a��>��V�ˢHU�A�Q:>'��X �stt�0���zxYJ���%��
�0cC���?b�p��f��+�kq�I0< ,q��e���?�}��b�ȨT�3����E|�Nﱀ�ö�F�Z38u�"_���q-���@�gc)�{ccS��yI�_F���A=���h3=5���\Hq�Ǌ�x�I�<�3uk{3���kr�SVg�f�u��8���;�\@����}�j��{J�e ݩ���B��	�Ȣ��:{O���|��d�`_�	�y���ͭMvP���[�c�H98&�L�9�N�Y�)ҥJs��E�����d��^�@u�[$P����,�NU�uJ�����nk6���1\�\9�e�7x}p�3����, D-�r��6mm�0�� d�������e�Vk}v�@ӹA[�y����tp�~fy��?������~�4�Pd���ZO�#p�H�ϩ� �� D�w��@��i;�I��� ��*uD�s3�E81 "��8'�+�}� ɰ�8KZ��R��HtL���>�{@���+��������G{̯������Ω�b^u�'R~8uc���~e�~�!�2Z����5A.Q��z���o^��.�Κ�+Kd�民&��҂v��*��d��m��֢��o�<ƅ�Ө���0hJ�;`������l�V*�G�i����/�Ӌ�:�����~�$�x�u�垲����z2�R��i�p��~���s�|�`8���k�mu�A���]I"�����NE��@��z���2�r�V��mz�1+t����� �w�-�ge�ׯ�uD\�)ې}��ޙS(�<Ep��ӄ�KR���=�u\�^a�����̅<�C��g��gռu�dar~�0�K��è-�+|2n��62�*��?�%Ou3[/^��権2�\���R���%ɨ��p_��`�72P���2Q�v�:bo�a�Z���㢣Քd��=�-+�����f�&�}���ID/�RIQh�DvCeP���}���~����=���=����ԢDٶR��5-��׫�s3X�T�y�戮�h��B�j����v�(8Г��Z�PF	<ۢX�UZ������a�2��$��1l/�7ɩG*��yP{z��[��4ꠇ��f�{��z@�6��s��]z�����������iš��Q%�q2�Y��'��'}��<jh�|t�k-ss�l�Y����ǂ_�����p���9F$�T���9#��3��x�s,0& d����nv{ǡ_�k�LO�A��� �ܙ�j���P DR_��A�B8j�--.p�3�S3���ҋ/�t�/��/�d` 3DN���g��@ep��[�|��=6T�5Z$��Pf@���p�e���~��̚UM*����.��9Ҕ�I�T���.mlHtq�+�O��D��Dp/�֎H����K<W<S 9GGmj�������̀s����!ϷK.�Z�[���y���X!"jjr��f�hye����v���-ai�}�Ye�pSؘ�qE:�v�Wl����Uf�2�AxVH�>8ܧ�>������G�n7�� d Ͷ]�m ?�ȮTі�C�d0LMM3���%PYR��=cˢP��	�����m4[#`�}��/`�b�3�c�����x^A^��n����9ʖ�r��@��A{
��Z�����d��!վ��ᬈ&˂����ޡ[��"k����t��y��ڗ� )�ϔ���h�w=��@Ƈ��i����{H���h��P�a�Os���f���Dev��E�p�F�=�q>��s�W9fJ�i��'�6Lg����xB1���i�(��	��֭������yQ�|�����-�8Iazߥ,�����ˎ�ȓ�����Q�j��?u*G�|�"��9�}s2��C�^��Y�����Ν=>�cy�T[��1% rW)TЊ2�P�}�Tz�"�e܏��E��)����!�{��b?\�6�&�A�<�:�����PD��DW�Z���5��i�9� ؒу,(8h��r���!�Gvʔ�~_�� 煮)�8�}/��Z/�d,uXO;��-}�aD�:�Y6頵��}��M���e�|��Y��*-���V�*I]���)ar��u��N,��?o\�#�q�&�]|'�s!��t��ZL�%�2(��"�4ES� ��)�"�%�/��8B�YP��5>�y5忨�2���(��=�mwg��y��p��EZ
r��,�pPL�b {�l3�l��f���)��a�S v��o5Dt�G�r+v�<���Tغ'���_��	$��ف3z����!f�{ʕ�tB��Ma-�7ls��"�}��� y��6�y�AJV���"�c��$���XK��N��h�����*����=��r���Z�2�yVFL���x#��< q��o=_��NT+�S?��U�ya�ӹ7y�̴(�̛A��)�c�}!�P#G�[-=}}��>M��q����e�E�ϲ�g���#{J�q��ڷ ���~�ƏL�pە+W��w�@���:ݿ�����j隮�s�o�Nx�غ3G�D�eA#�*��-��0Xm?�՜�ap'8c����`CׇQ��U9 E��$u`m4 *�E��CD�ݸq��MK�p����D�S)�PS ��v�u%	��`������6�7��Z�P�t�p~\�?GPU੖⃤�"����G�#@fIQ��K
}0����e#R
t���δv<uRTσ���#��P�i�tqu�v�dĽ7��vxtL���gl(+0]f�  ���ߕ�킟s��K0pυq �~���p�#���fP�� �F'a�\ߠ/��"<�)���?������L���X%�Қ��|���U��ĸ��,8/��tO�b�� ���ߦ��z��^��sf��U,�U��/�hL�aj�0�f��wK�H������^�+�)��GV�U�q*:��PW �����+�+�z�j���(e�U ��Z? W��Q��'�-�3�"
s`��������wF������cKZ,�-�·��rk�"���ReT��T�kJb��M�,����c���]&^TQ�GWr���ҫ�sx��!�X�}1ǫd���r�����W ��`<���
I��?����r�k��"9�p�_I|P{�c��{r�̫��ZsCߑ9"�/*،9��-�կ~E��{���ar*̵?/ �Jg��+($����s9�]�PZ�"� ^1E�80�le��������*��j���S	{�FQ�OJc p��W�\��e �ǟH�Z! 2����$5 ́�9����Y	�ʂ����p�8����8�0���}��bn�A)��&Q��^��S�с8=-�d�>~��n��ff%S�Q�
Xw#5N�Ϯ9a����+,R�F�B1��Ԍ-��(���4- ��ɞ�y	�M�U���{d�g?h�2YPWA��V�A��]���ua@����8Cg%�<?�_~F�>{���������{��f���T�qzL���dϸ}7[}�$�d4�ly��I��l:����$b�u ���}plɚ~�J��X�H�Rvɣo���$[�1r:�O��\䐮
�6�u���M��{7]˨ŌFv ��)�R��S,�AP���J�����]%��N`N���B'�}��t������<�.7~"��TTO�`�C���^�fj���}@�<X'�����V<a���ily�{G��������޻��o�G~������B)\�G��Z*�e�8�̨A����0Ǌ6+�U�F���_�$���Ê;D���)�
*#2vrB�� ��1��SJπ�onnq���ь`R���h������lr�0�l���Hs��(k� )�C-��("[Z�n}m�Ο;G�����N��r�lG����0_�CZ��o���lM�5��G���Q>	wZ��HԗTn�`���?�q�((+�nBt �	وϪ�I���p����loIq�0�+g�����U#�����skL�Q�{GT���߸u�v�v9�cpkmm-�wP(��ߥ��cN��A�H���y6�1�8ʲ��.���|o���(��O�?���e� ��K�L�f��p�@� e�W��}���<υ�bB�>:K ��^z0�-�2���.]�H�T,N����@vd14Z�0��ȳ�D���d2�Z%���y�G)��
�g:��߾}�nݾCk�k���v��ݤ��L2g]�
�G��%��
�UY�1`!�����:�	^�x�e2.����Uz��'����� ��Pr�9nE~Nh�̅&G߈N�F�KA�Nm�������
�����2�޽���lN��A�~�4o4��)�j�qD�G�?{��1�y����o�L.?��dB��,��!�u��i�u �޻w���O��ͫt?́3�+�D�s�Nr�,��DK"wy�]����s���F3rsw���hZ���E�K3�7��:׻����z�Pt����"��	���Y�]����U���Ba�'ɬ�9q�(�[*3gFi�S�MLh�>����:�yMb~�a��|���c��/�3��lm��w�O�עP]|�s�oȠ
�AOr,�����v���<�Đ{�ABN��TJ/�$x��s���)b��fsN7��X�w�9�QVG\���e.��X��{���D��v��J�D��S ,v�=j_�G]�~�Lr��9-*؊�d�w5G)Q�.9Q�q6?n��M47(�GM9q��g�~F��cV�1������oț^W�q�]�F1pYְ�2P}��G��s,�hu&���,�-�eq9Ց�Cqb�`!	�q��,�,W'��d���	(��4jpU�
@�~L�\Qqﻖ}']|�b�Mw���V�_"�*?Oxs����yĥ��(�������?�x��oB�۸=�-Nw0L���4���}�A�/���Ӈ%M�E�Gg�aoQ��z�����D�0���2b(bc�9
��lt��J0��r�/�CF.�7/��17;���؄Ɍ�7�+ V�ZLW��:���R*\� La��0Hn߹̀������յ5Vx ���7�A��q7�F���8��&�<�݊�.pY�����~L��ߥ�W���˟Skn"�C�676tQ L.�9��M��
@�SK����� �gՑh_񀋒��<�����^dD���=KI;��|+g�J��S�A!c���K����cE	�"��`�bl������瞻ȼ�GGὝu-���{��]��gh~���)�[�r1�*F��<d��Z}�)�_�TS���6�5�E�p�<GKH�D�y���և~L��/�}��'<�Ϭ,���s*5�D�t>?Q�Z�\>��?���G��.AU�,sR$ʀO�vp&����&V��K�<"T08�{]���N���k�=zp�ϑ�hS3�����5�+��6���ai��ҵ�D�x�L���AvA޻�F�oܢ�_�!=��43�������+���Lu�u5�`o�e�8	ա�
����ш$+���YЄyJ'{O�)h+���x������%�l��C�S��-��'|�r��Z��?�3�������7���S�����f��C|a(� ����	هę ) �����W��5���47�
k{2nD?��䆂�.�P$JR�U1�CC#?�gd<�<�x��*Ȫ��peb�9�A����ݝ=�C��쬠�@0رÇ����X8r �N���z �q���ч�b��SQ���D2s�_�<GG���A/i��n;\�B�V4ڍ��
����\�OWX���p:��I@b�7���"�) �Vb�L]&�P����EQ_K�n* ���R��� 7�a�I.���ňb"�Yr-���)@\��8�3>{���-�\p��ȸ��w ��f�e�Aޫ�y�}�P�A�?�)���󊓏ї6Oc]�ȬPs�S\Mf�۸=�6D�N��@��Z����>D��t}B��؉=3;=���sF�i�(ZI�^e ����%���;��d��}����཰��ɉ���kc� ���t��O�>���k	LN�� ���Ld�m6��=��������"�3���\�C��a����Gr��kQ=Ҹ/��Z�����Ё�b��n����a-����+oܾ[ͥM+��$ڪ�#� �k��F׮_g�}BSαy�tI�_��|4�K�8�h�u��xBT��� ��zc����,K�g+Rp��ys�*"L���ox6� p`��tC�8eQM�2�ф�> �
"l�0��&��>` y{{W�ؓTR(MAf��l�\U�b^\u=�~�h $Z��<���{�\� ���p�6WZ���e Eu�&xڡ/���1�Ԟ- X�h�3��JY�1��?{ݘr����}��v�`�G��N7Rṽ'{b2��Yy&9-:�~p(F6RR��6x�|�p�"�\������v8nS#ͅ�qum��_������9��r4�R�Ռ�BR�z��a��w%�l<�{��@�0� �j��?������m�� ��&�c���j`�1�0u�<�C�$�g{�)���O@+�&�D�H�����p|�D�N�A*R� _@���=b��� )�R���ugYD���j�YM����Ō0�,�O�sI&[�H�N�,����o������e��RR��)����A	�%�`;��찜S�$9�}�A��BV6������/8���;L�4�@]ߨf�-@8N�=�	j�s���&����o�\A����g��l���<3�/r�쉏0�2'l톩~��Z~ߎ�J�d-��5���Z�Dh	�9���O?���}����3Z\X������j���N���^�b���8+d�=��X�ꩣ�����v��X�UG ]�C县�ky� �%)�g�y�U����Ɏ�y�EXS��U"�gA�>����4�.�[�IԴ������j�z���:���1MM�0��:	M�����
��ӓ��H��i��X9��<�Г$����;T�dA�9s��z��r��N;��b��Dc"�x���Ԕ�^�@��B��)f���g�=��H�,A5��H��i(��������鑕����z�������0���)΀�`�yf���T��"22TWWWi%Y���܈�ӧO]�[.��C$����z`a#��
��q��j�x,�I�ޡ|e����
_-u_��� 2�&M;��Ǐ|�����=$ϰ� X��?y#��x\J�9�oI��v��$-�]��m�f�X��kFK�h���~���+`9c�R|�f�9�`�I�ɴ*�7����s�e���`�����J�%�y���I�)�r~�m������j��7��q�rdG��ep���8Q�����e$L&���/#�aG�:��r?�A��+g���6j����H���`<�� ��
���~u�����ii�g�د������|��]j���� 8g;���&QQ�=�NM�gYӲ�C!|t���d��� H�N$"ېb�\��1�0Ye�f�6���8��\#�nU�����to\�PgȊJ�2t`�!S�Sr��i5~U�Ǆ85=%��I/,,��g���K�J��t��314��UQ�a��bu�1�?肕�h�FZ��̔O��޻OЪS�A\&#rrz��'O�����?~b���^����!D kG��Z^WG�[� o���+��0,��d�S������Q�E���Y� �z,���5Prr��@����qy����:��o�[-y�lNM�e�bsss4�._�@>���p��j1} 4A�<8�ڷ}ہ[�{���Mgy� ���I����)�`��N �+�:楎3���B�(���EW0��'O�	�k'	@�܍h9���H {m<`��N�cpk�Xz������L�u�E9k���#���U��{"[�:�Mﴑ7��)�l4����g���OK^*0� ��aٓ}f�X�g��R���n��`l�,��gϜ���1��$���/C�,J�8�N����K�L��~t��~6���'�r��z����?w>���Y	�&٩�ڋ�:�%Yd�"��s1�A6�x� {Pp�����UΟ?��	��ڞ0Q��Zv?�2	���e7k�el�����ɟ�V41w��}���ȷ�����l����>��J��{�$$�v�P�s��{��c32U9�)}`�,󀣨�9�	���Da��Ijg��:����:��,��G��=4��"X�L�m��
��]��T��{&��n�+�H���_��a1M|��o�ȣ���8_�/a�������`�p������a��y�s6�C?_2JI3H���$���<26̀�_ -��0h��Gv�ܦId��X��@���W��!�����>��M�_�͙�K'���j��F@�P�l fm4�`��.	���k���� ��:�S�gp�Ѐ�|.x�h5��O��]����E�KzҾ��"���A_ ��)~��m#`�B��V�6��7�[x���3%�Z(��آ�� ��,+{l���w�>�<|T�cX�& �g��T�5�a��_��
���ڭ�-��K|0��\�rJadf�D�6W����I<�M����W�?�bL�!��,�aPI�~ۀ�����P�F� ��Dj�����s�^�u�\Fו���X�ݟM��jcL_�>[���U@T�����Z��f@��6�=����Ʒ�Y��x�����������9��T&�p���3�jN醘n莕�S�vl��M�x�� :;|-�Ao!��B`9⚙Z������*i�bRCZe:�X#�V��j��i�Z�)+����We��S�Q�Mѱ��tE�j Ej��?�{���Bmc��a�DA�F}$ޯ2k ��4ڂ ��#]��*p9Y�SG�R�K��#Ur� ���<�3�pG��	~AotcdMFGr9n�_׎,-ù�~���3�)�t��?[[�X4�Z�yCP��q��{��f��:�Y�(�@ÿq�N��4�뻻-y�|�����;�jd�qE�t�� :�-�`�9?u�wJw�/..P�djzL�ͣ��w%�D��nz�z�@�`k�9{�`_�ؖ���4���#3�qf�����*�I�����Y��8u՞���:H �ڵk�����3�3&)Pj)3��"���%xF��7<2�B�'O��<B&���}L�>�t�[K&���@
t6lNm��&p��C�k��'W�kÍ������2���dQ�4�a �­%��ةa��+��a�`�瞤�͕U�L-�����2� ��d.C��˯�bz�{�M`����\� O���X��6�����JN�?�v�`j`O�>B{X����Sm�u��~�"���o��2VjW�i��r�)��׎]�{�$�&7p���c����?��0�1x��)�)Z�L]���0dD賶gh'�b��z���*[�%=����V�-W&9S��8�^�7�|�b}�`����7�������@}0e��:�"�Xk1�"wY:1��"q>����C0���ncW3)1V&'&	"��dq[]?4cɏw�5 �k�MГkd6,"e�u��r��	�t�Ae���ޗgO�R��G@�ikC�~O__[7v�^_c#c�@��*^þ�/f�X�	�4���{t�]�sͳ��S�i�w��{�؟��f?!ht��X^C�ҥ%����CZ�W�M��> P��f��8&��xowGu�Sx�ıW0� �`yE����3YҺv�ƪ�h���׵��9�k=|� <�z���f�E`y���7X�����[���W�X	��Y�3����P���/��ao�$3&����G8a|	���?��a���F��6���~ ��&-T���.�[a�T���n���B1�,cFm�sڇ"��}�����=�� T�cٟR���<dU��P������ ��4�F̞�S�r]�A��r�����7X�"��t��δɔ: �ڥ�1���a	��rܐR�:n��ťױ��9Pc9�[���E?�-/\�������;t��H��y��Z��0��a�$8���Wf0����|����g_�&�ZE,D��3��ZHP���D���+|���f����)�>2�� �� �zb�ٸ��L��t��$/ <v����%��\�_�I6D`��M��|'O����UU�&@20��T�O�c�){��V Z�9���E ��(#i��l)����,c�:��GH9m��y\�ѐ����h�P�h���$�� :��ˑc29=(G���Ɩw��eyi�;��U��x�-�,�v�j4rd���g��?g�� ���j�ʶ�s���ܤ3`�@*�d2ǽ#	�c:�H���I�c1��! �3d��@kyb\��G��>B��Ng�_?�B�n���Z ���	]e󔱸��-S�eWV�`�HHo<��@c�GJ9���f?����s��=��|Ƶ���3��1�0G���}��!H�����������b@#�!ʒ��{=� ^��^�ZfA+0�11vɆ�ג[�92�  6L	�Uy���2��[]Y�̊^�T��sI&;X�F:�*{)�u�.��n ����lFx'��������$�5���en�f=x���dtl�:�:'���W�B� @"0�T7$ +h`O�g�\2��U)�U�>1&��:�MaE�DY�fr&�SHo6��ʊ�1��jfҸ��]�>�����/���#Gdz�(�1�����5H�UE!�K&b�z�(��oݐr�}�m?y�������1H��rA��~>�	|���>�驩	:��VS3�l��]�nY�e�_J��l�"���
��@ը�mP�,l\�VO��}pph��Nػ:�+[�(WeS,��
Z!J�lԼ�E9	���Y�;Թu�&����@-��E| s����Yp�;-�{;n�6A�fpp��n�|����}l�r<[1K��f2a�W����� �8�Z	���(�:�����<��������u�S�ڼ[e�v���HQ6#7"Am���.�D�O�~k�c�Yc�?:�hv���V�!H�(��C��T�� ��*6�Ť�q��i����^�=��ɐX�ׅ�������02�W��E����$���=������C&;l��m����R�9a�L�`>�`.�$e6; 	��Ku�Á�x谁�a��*�졃���tx`�%@�=_�l�`��2���2��U�S �(���.�1d� å��oo���[y���#� ��AO9��f�0���]i�ebx�dC�^Lu!e���,�f�mhV�������^Dż�
�9{��[-���9-j6�*-)k�ou�����J�������~C�����f֤�Z� u0_u>f���s ��^'���l�ҀF�>�d�����P��1:�@��S� 'fr��贅��n���:k��w�j$���/Y�����VZ����?��E��ܼy��ܔ��q�b:c�����8p��'t�;pcЍ�?Hup�NT�G���e���3�oV9��	F��5��m���6���ݶ�ϯ�y�Y���)�����%u��i�Gdr�-�o��o�}��N`F}�/��"�v�]�Z�,6����=3M�:Ϊg]��ޠC	P	��Y�f{��$'S� M���a;��D[xVp�<�V�2�w	��ƴ|����H�}�W0�J`��m߷������_��a4N�h��6f�^2����
�Ԟ���.�<�-���d%W�
sp!-�T�Y��cΥF�a2	�^���,�nT���v�]s�whic� ���j��������F���)�t\��s��H��ú���\�n��\�z���@&�zc0��U���4�x�Z,��gb�~���1�0�+�r�s�Բ�ߖ
�t�!��hEa���{G�;&�������Fd�՘��d�r�<��V�tТY!�e/�,��-�����)=q�8%+���H)2,\3����GL����Kg���g��Z۟}�����u���T}����,�0Lo���g�Y�����v���C�ɜrn�7_p�*�֙,΃��`�~��'������ljr��e|�������Y<C��*���`q�S*)�j<���� r�BAJ�`"�~sF�)��`�B��R2tM�X��a,<:�S�o�����U��N�}X[���3iaqQ?�p����ɪY�J�0	]��Lk�,0��=+ �O�rVJ�U|��5aM��-x� �1��ؿ�d	@~��EP端��O�ig�	}..-����o�&և`[ @�5k{۵m/�ͅ�������O0p���\�+�W� �uH�]���5�'� :~���b�3�/\����Gǭ=�l���q��!~��� ����[�(]-w�{�
�e�u�s!�&v��0�.w}��?A+�N>��^8�r����g�zI��fhű�+	�NI�W͒M��@���=�ľ
w�^���\��OV�;
�6iB�4���nP[\3y[V�F�͊p�:�7X�߂k��H5Vr���OL��e)U!I ���Y5���*�����]�v�)ݿ�����j{chg���m��N
��;��c)P��,�0I�^���a;l?��_	�6�:�-�c!9 ���?��oy�l�`#���!"Щ�f�t���+:1(��t� X�6�	�6 t! ��c,ƺE�q�f�&�7��*���Yi��d��$5_4���σ�����=��,щB!��g���.�@�\�z��>�������p��&�
ע.2d1�Ǐ�`U�Q����W\öw:ч���bT_`��0�zY�����=}��;��d+mm�P�bcsQ:�wF��w/��˥���OZ������>�ɉ�rᭋr��uy�pV��eb
:�`	��:yeY���w�J�h ��(�� �)v����|�&o ��j!-��e<���I���<����gp��h���&�C8`+�c�gdiy��ҭ>��s0pt��ݿK�����,� ����=�RF!�cV�
NY�}��^`�^��L*Q�1�Y`�ב��g���۷���K�	�Ǹ�~�)�6v��(�rW~,a����s��1����	J�w�w{(4I@_��@o�{�) C &��F}Ș `*Sv�����r��M���i@��ֱ����-z�I���I�@��^��s����M�v�F�ƢO�j����"���lTC~.�D�B��Xۦ���!?�fׅ�(�F �V���O���52(/^�@�� ���aoEd��,�v;�އ7Xl̯ՐC����r�_�o��o䭷ފ,�`W�Ս�X����I,�#�#��༊��ұl�؞�2.�\GV��U�z�YY�����m�&�?o�6i� �ʰ^�&E��<��Qt�0��複yA�,� �L�v��m|r�� � �Fn;ǵ�U4#ฒ�ӿKvk��Ae*����{��'����)���0��:�  �q�`NSF�VS����lB���X���ɹ�?����i����S@���}�5���S��y?'>���qX�?��֬��{��b���U�@'�ޢ��6�k�KHm��]�2���lֽB3���Ȍ��43A�a�}�����s Λ�[��G�f$�QJ��'V1]/L�ę�R�+�xD`��jQЮ&PV��B����{2;��`t�K������Xh(jc����l�8l?���~��h�=�DIH��*2�	���e�V� =����$��i7ε�H��U��u���»�񭗙k�n�U�$��P�{Y��B�8�?u���]j�:���7X�2Ё]�N*����
H&;��DK9��6l�A�/2~�9\d�\�+�/�hVP)x��ɥ�}ǹ�v\�����4�.QE᝸�dJ�K]v^t��n|�	�׼u1��R�͈�i�s���.>����l}4�H&&�4�\�UQϭ�R2w��u55J�V	��U�QS3��<�#�p����Df�]4�,ڀ�s(|30���!Jk�Թ�(�Z�p0b�n������7�^�Ͽ���0���c#._�P.�>��N0��@drj�)��J�}�1��fKפ��A���us�;�G���@�a���a��}��m�i���7�+"������.t[��)�kgϞ$ �b;++k�vvU�ō����
�ՠ<y��mş�c����ȹs'��|���֦��ހw�u�Y�Qe7��@c-nMise�Щk[���۳��i�/h,"�~,�BW|  �x��
b��X1��%^����p�[=F�ی��e�wey�Z���ݓK�#�ʸ����J(�M+�K���E#B#������}�O'N�K����t#?~,�~�<y�$��hG�K+��,���_��Jr�� ļ�g{�ϧ��a:W%b��v'}��2Z!����.� ��dP�@��}����E����{<���{��`e�V)���V%ݓ\Z�_�}� p�����[�A�3% X���{�ss�>������TPkȿ,��|��#3A��f��}Y��T�lu�.�����[�c!���������k�����8�Ԗ��`(L� Pa�u���ܗ���x<z�:�`v�����D�,�(Wv�3܋K��7���Op���3 #A�"K����D��?�����}�L�~�չ�Sv�{���"p�~g�Si��[�������l~c��^�kbA�vK#�ʯG8�Z019I0�ӍeȖ6W0.���#�j=�:����d�5s}C&���&B����i�=���S-���͘[$� ����bd
�DTv鞬]���JF1�{y'ay�O�\2 ���A�t�O�<md���=4Ԡ4��|w�G]��؈�=L���g���N`:���2��؍a�M�'a$�,.�G.>g4���Y�u(����'��ߒ@�'��)�A7�:ׁ��%-�U�ǁ����\�������(�޽K��\�Q�Z��)�V��K���"?$���0�O`�Oga�5?0S_afœU��d�$��ȓ<�c��b�FM"�%��m��k�!5��=s���e�ʎz�l�p9��;��j��%d!�6j�O6rJ�zڛ,�"�~Fb!�
���E7;���*T+G�X#=)[9�ӴҢ��o�W2h���������'�1�4��k�����(	��F^�7�7$�r��պ@�����Ȅ-T�雐{��Ͻq;'�CLRR�	h����9���E��_�)�4��g�Ã�+��*E$ص*i�����m�4E��kup� b�AЂ��phE���-:?t����Vxr�������|��d�9G��ޓ������_�Fnܸ.����?�3�8HgΜQ�M�akaqA{'k/d<.\8O�3R�����:�4M�Zݤ#���z� ˕g��cI#���8 k�r���oҩ��3X6kǎyG�c}Wȣ�Oe~~I�<y��	�LP�������}��?>#�OL������k*�E`�egkqQ��-�n��N��!�"<��A�Pɭ�G@ �j��!�5�[����8/>�g�����q�������ޔ��e:�0F�ޔw��r�{�Lf:�t@)�Q �g,(HXtht�X���_vR �%��^l��hd I��zP��"�ဏ$�i�����bJ�l��Az�W�\a`sul|� �������}z4c����>}�R
8^+q8�^�`.	L ��k0���I�?��W�|2	d1\�~]�߿Ǿ��u��T۽4P'�xa>u����,GG���g�z>��a��������^Im�,	L���^�T}�v,Ppѯ��* ������`��� A#��>jjxakw?Fk��U!���g����3���S2Q�b�W����U=����9��K X��'r��E9u���;,���r�,�2 �/�Z$���~6�Tt��|��@2����\K��r�:�ؗ�NǸc�:�+�K��3�`�u�������ٺ��⌸}^�;BV����e]L�
vj0 0N�4222�5�Cb��&��5cum�kH�@� ׅ@��#Ӽ7|�/x��#�[	��f0i����s_�jխ�D2&B �M�c>$@f�-���+�w�+�&�������2�6�/�"`c3+���g\#Q���������q�@a�Ǐ�(�Qc�\N?� ��ΰ=��Q.d�`0O��`8Pb�Vۊ�Zq�,�k��u�2^�e��A�fxh� 6�	zѸ~�J[��*W�gX��K�4x3cG� ^��=d-���mʞ�l����&�! ������_,{-2��~+��`s��?�Eఽv�A�����v\۵^L��r)����O�)��`Q��<\��|)��{^�a#��T1��J�t�O��g#:퓰o�$]f��:�z��ͦ2�՛�� `9�"���X�]�H��a!,cܥ�"M*)�b1w�/��3��m"=h��gU?Hl��҅w��{�!���;���*��ޔ�b$0B��)�z�]'�3^��>CX�h�#9���NtƐ��������; ��}��/������$Aϊ��|��W,��U�fY�֠غ���3*��:�����\a���]��0��081d1�A�bYY�b)�߁�$rЂs��P��18���O����{�y�ll�ә���ꝷ�f����T[0��&�v� .�յeYZ^�ba�� ���=�?M<�&�ha�����b��<YyC���5f|u~��ܜA0��!��_�Z�q�!_V��x`��$���ޒ��U���0M�%��)������:-�{���&���|omuS��Ч�qXˬP��L��N{p� w��*`;���`	l.����cp߫�,յT+���8���.�PX�~s3:��<�C��FFJ�� "O���<�/'n���v!�t�61*��bTe�QOvή9�*��Ϯ� �Ӳ�����~c�����ʊ\���\�r���oX���'�BSa�b/�Vd@�`�� ��/ 33�N��@z8;f��m��``ײZԼ�]E��o�ܠ����C5֦��5y�h�̲T�1[9Dz>e.#�%�M �+�/������ｏ*����
����^J�7s�L��A%�K�K�Vcyf�]�\v�g�t��2���Z����F� �"ɂ�B��ho�g�!>h�D{�Y	X/��=w^��US��T��(ݔ��v�q�?� �B��N�j�����o�(
�MkQ3�!�^6w8�2�^�%�;X�%��R@��+(u�?���'_~�l���vԏ�F���>n�b�Щ,����<@����/<�$۳â�-�{�<�)��[��0vɼ�,+�@�~p2�Q��5"�U�7�����!J����Q/t�v(�D0z��߰- 2���:{(8>6a�q�K�־�����F=���{�M���4?�I�c-ڷ��z�r�u5<o�5s�Ԭ"�?�@PH����-y��	ǇL�� �!���� <��X��Ņ%oW)���[[����d�q�8׉�4���� �=�H��P��_1�`��k̨����2>1)CC:�jM�9<e =ŝ�{Z���q��_��.�p�j�+)=�H[��)�P/�Z�u�.�jI\2�� �a�u�N�{.��������e���u>��b&��H�;���@��V�v�0'���%���u��#ν��]�����lj;Y�	ѕ1��$ش�H��2֔<s=��μ~�5�{Ze� �Z)e��f�vJ���	ZL��\�굝NZE�Im&=���WE�*�ٶ# ��lV}PK+��XgŒ6 �w�/�QVђ�۠��L'Ơރ�j�pY&R`9u$4x˹��\
;@GS��� %�@���4]�r-M=ǆ�E�}&bY������}�ni@�]�\ ��q��ؒ���i�6R>��Ϛ��eX�*F2���5=��r��Rm\��;MW.L�z�ީA!���,Ԓӑ�|�	8�=�y?`����1M��EG�V��� 1��������Ê�O�:-��:'G�L3%�?>���(�����o	,�\O�>��w�6��N?v\�y��~��x����4��y�ձlp�Gk�svH��禯����$+���V-��{��o�2\�)O��ZCb�ȤL�Lh%��yYX|杦5�y'�9Ni�ՕYZ\�ON��/���f�c<y��ߤ��z}�{�����JG3P��"��+�H��K��ٱ�����1���m�;xms�]��ת�p��p���EX�q|k}u]A??N o��עSzg6�T����(�5�� 7o��3�V3�.��j�"���2/Yi��`�N�juO���V-�ϝ�%N➪/W�� �mW��Qc�w�5S�����D��T���1(�x��Q�#��a1���su�;�*@5-�2�}{@�M���jCA-�������@1 �������g����c.Wj���c#f�����ˁq�������[:D����$���V��8��E�ު��.وX7.]��{�<+���b&�� ?���fK�|���Op�@Z�v�� a�Y��p"e�e�LM���u��i>ǹ�'���Ŀ�z�Ѐej�W�S���븿�A��2��4��1}��i�/_�؇��Z;���Q�3�o����@�O���*����u��4���; B T�v�����k<��VSY°�C�f�ȸ7��tf{D�	6H�N�氖Q�kD-�:u�Ef���������y���N�>��Z���ua������'��Т�~��?��kOǏ�1�W��8� 	��Ђ�N�� ؀է@�l����8d�����C��평1��p������e�����~=����O�X5硹����(�* ڐV�ը�	���	?/�i���@P	� y<[fpe*3�3��յU�-an�&
��N#)-&/��	�S��ۻ��ϋ���������,�XA�g�C��a W�!㐭�e��(���Z���IV˧��P <��e�|v��c	�gϞ���-�[!7A��9���d�3�VI9l����BP�*f,�/�����L���w�������"/g������� �/g;�#[�����ݛ����
�W�Q�N$������~�Ԃ,��uk�9�ܿQ3�ժ��D��v��i�P�4�Y��^S�rH�����^� �e���۱�ʶ#U�	T�:i�@+���L���.����Q ��U��4�P`B�i��j.N��"ھ_'{!�ѓ�n{�f��	R�Zd'���j�0چ5���39l��'�����T��E�k�ί���=�
볳�thtM�ȋ��y�5�.ݬ+ �L4��3�M�����
�Ѯ���@�U'��2`�L�t�J��n�m=��=� �yn߹#W�~'��QB�)X�gϜa��3gN�7�|K��.�%�����/��}�i��c�?N�֜:-���d%7[���s���*�V�k�_��T�/d��~X��H�n>��b Wdg5��<B�����,,��	lm qX�B�C\�K�5:�hI�mȚ����9w�u���q��/�B�=*�����<�_�@!���hnl������+�0�C����(	 *�b���`�9V �q0^`�s,7��4���U��?~��|yy�.p�����y#=Z�O`)C��=���-jb��l#X�G'v��2��a��_��(y�k?��WN��n.��l�?�$\\Z���a�s �K������9W�h����k�B�<:N-ۣ��M=f��B�gc�����`�H`C�k�q�
fmQ[|��>eS+3�c>��Q��k����	�P(�B��4���x�����-��_h�@P�E6׾��_�=g�θ3��"ʎ;qvN�
���Ż��H��ߧ��7�6�o P@@�J�]�7S.*� �Nbi���)�	h���{��gҎ��\�^=������u����������G�,\��krj2J(P� O6��]ڻ��~N������~��*p墬UY�
2@��O>�z�1�}cF��UZ{
�8�zx
s��Jȸ	>T�$"��D�DD�T��i�@�H�������	׸a�!3���\�.��! ���ޠ�UY�#�Z�޻G�����������yR9�Ad��&6@Z�A�8 f1��' \��.��m���S�W ���"K �>ֺ��v�\����1Jy�Q��.l����x4;�m�'�o9��poSB�R�����V��(���$c�y[�����_#`,.,�Q�� �]3�	�?�}�{�3�:/�c|>�N�N;�GF�*m=	�H�lڡt
�1��zӰ��ͳ +��*+��?2��@��۾-.W����X���v��$L.��h�d���K��&;�>i2���w9l��'��2��XܭI������+r��>�p}��ek8��̴V��	!�oo$�Lv��p�E1E$T�$p�6�r[g��U�3I������-�e`�U.M��4��#���3S��Wi���
�;�YyZ9xMV��{����(6��i�mj/�Q_�~��,���]-�ϱ �Ɔi��Ҫؗ�F*O����7��̴�AMW�b�#���WH`ܺyS���kY��nd6���zf@�L*���j�Y Mb&�"����V9�%�0��kZy�i�����ꡂ]���#���y��!_;2s�l��o�'�
gle�˞<uR��/!gN�b�'.h���#R��(���C@��ihЋ����*��?������X
����#Aϔi�pf��50x��+�7!AR�k!λ��U;;��5��9yb\�ޙZ�z�lm�I�m�Hg�ɣ�y����w�W�Z�/��J�y�wx��c����-Y[۔5�Q� ��w
��NYS�u���4��1 &�i2�%�E͞��*�'�w�q<�~`�OMM���w�Ve�����j~0^N������s���10$����s�4�
�
c�g�B����Nʄ��"��ϩ������4����������e��W_}M���G��Y4�um	�";m��0׎�!ˬ��.�b51��"^�Sژ�V`���=8��PM�nZ��20?�3��M躣�&�A��=	f3��8���������N��m�pz	P�oK��\{��>��=G�.h�0�k�����4280Ǚ�`�0f�_@�v3��5��`��	;tOG콦p-�Er��k���-/-sl����v](�qmGk�M�c� d<p\�iO�8IM٠���03���+53�k�+�jnuC~��c�T1������q]�)�ˢv �v�߿/׮]#��@�K�+~�u�m%�1*)�0��� 
1�u�f���ۭ�2z���$2�K+f�һS�W�]�m�!�>�5��)��2nB�� E|�����օ����N�=}�F�g�/�-����u��Ǵ-K��׫��gvw�g��,[[]��6鞢h�E��dmY�^�y�/������h��`Ȍ(,���9---�cl��M�1k`�ry�23��d����b������2�U{X�z���ǎij�Iv@���nY�,�Wr_RY�FԠ�]��� p��^���JD�D�g���	���uˬ�}lc3vdyeY� �F�����ʀ�Z
;�3��������u�U�ϭ�{[�}��uM�=�X���̋?�5��U�5�]~v�_��Tf#RT�Aٟ��z��s�ci��d/�m��l)�i�r�VF��j
�n�&W��������U�;�E�3��G��N�9�U�.e�EE#�,gb~l�5�\�7+��2;wWn߹���299FCF3l�(�
eƂ��3�Y���8�4E�Z}Z��� q����Rs�N�z�\��@�Q2Ak��W�~KF/_����[�Y�>.�%�gG��/
����i���r﬌P�p�������a��`���	�Ƽ6e$��%�ra� `�---�7_-�|{�lC8�d�;C�2�"h/����K�.ɇ~@���?%����򗿔�Gf�p��;;��꘶�0 0Jp~86�n�� ��IX���s���A`=8�Z�g���ёq�X��o�!�\�dN�8y�@.p8�Ϙ����ږlm��)t\.�Ӓ/���,���
�A�]����21~T���}����{�h��3��l8��ӓ��Fx����l+���YiF�j&�|�ؿ\U��k5dIP�&d7B��Pz��gje2=w��D�Z�K8Z�~}o08���H0ga�8qJοuAN�<.W����|�?��r��[��{����D`R7�"��0�Ka,E3��p���@���F���B�S]���Yu�ś۷n��Н�w��֚�L2�^�+ѩ*���e��:��)��,����� �U��:E���2� �TS�����@�vR��U�  .��#=\-iB{��x����
��m�k�>���{�������Z�y͂����d�u��Y�� ���~:}�L�u#�4���u�LK��c�G�N�ߊi��>״������S�{���"w��Efv<~���	z��mZe��ʸǠ�,]���.��|��wr��E�w\�/R���λ�`�Dbʪ�dO �5n{��s=ˍ�v~cl��>�[~MA��ӧNq�ܾ};�%+4(�C��E���*�����g��� S	b��5�G���X(M�"���]�{	�H�`���A��f4�>F0`)֙ё�\@q>���/����F�����1s��V�� qq� �����C�~�f6A��ߗ���:2NKY��$h���8��d�k�D�$�U�~#;��=�(��gf��(�?���ƾ`0������9�96:� ����уYo?��<�������?~⤟'���2v��B�l�@
��䂰�&�9o�~m)EWP���_Y��jd�媥O���.A]�S���:[�v���P�=9��l2���\�������>���x�k&�,3�Pc�"d.�r�Z�4<�y���sn�Xos�����O���U���]e������Q�1��G��rO�ї��/�B�o��F˱ѷ�H�klª���Ƃ͗��(��,��A��"-cE�ʽ p�8{�A� T7�0��4�R6o���L^�jn�E�+��n��Sਲ਼�ک�&@�&#��~0!���a�.��x�-���ZM��4�H��U�E����u��h�,*����d�)�������պ�����H�o7�N
�}��7��#���azQS)���OZ����ok�2��`��@fa$~��`����"4(LSW�W�W%5��6�C t��ׄӆ]d�ʠ�
��޽��#�}��N�:I��ڡh
�{睷#�(�ip$Co�5Xsx�ue�ۭ� �T�a�\%��V��`�3�n�y�`�h�!���� p��g�|�5��4_��±��2�������}����ȱ��ȲЂ�h��V��ֆ|�������~��Wt� �5�u n	qkk��
�`�Í}� =oF�9��Z@�c @�kC��P�U�	ύLm�E�N�˚\�w����ޡ��4�R6T��;� ��}�j�d�t\H(����/ɷW���~'���&[y�c�ӆ̟ |�J�0q�z=����!������oK�
N����a�vz�ʏ�k:gYx���ZR��2��fS��e 4T�����(�D�l��¦��"UAc�W2=���R��G�Ā�Ύ�a�+��{-�l���]��Y +��b�!]���/��b�,t���r�����}E	E�߹]�/�Ԭ�j�v�x�z�҅��m*�F�ҕ%>��Xa
��Q�8U	�N�j�a|*��-C�!xo_z�?�k�z�n�l��Z�}Tv*�{'�XX	.o�P�w��M�<y��)�.>gR ��ά u�_
�Mia]�XK��WL+�"XK��z��e��4A��y�bQ7��!� �̉ӂ�eK�5�kɠi֖����CmG�k����m;�zB��STs��xM��=��ɓ��z���%�
쏿�կ�7���L�}Lz�IϞ?��.^���Ԏ�[c׈1�P.e�(����r�L�n.��
Ah��|j����{�Q��W�|em��:˰[�X���.�͉� 8~��!en ����2`x��	e��ʊ��,���"mIH^� ��Gf&e��'΁���j@0�Im�̗��AN+��הݨ���f��1c�$���8�$(�+rBث�y- )�� ����yڇ�VQ�_���c�
�Z0�g��R�W�� �TdF������Ϲ�ڕ�g�g����9�c�a�jў��������t�2�2z�
=�� �����u��������H`����B�̖�!�б���6�r��~� �!uT[`�v��*W,
'/,:�2�o�I硳����,��I)�w���R�͘�ް���+�Έ�(#dΰ�C���P���6�I��~E	BՕ��L�@�I�3EQ��cs�ۏ�R�&��0�& �:�p��s��,xG�N�i;\^&��Q�m7�a�PUH7%�zl�
 ,V�>��a�m��֡�!3�	���h��Թ�,n�\h�^:��޹��.���j�ǁ���{�й�:����uxjr�������"3oHu�є��, e��4U�NC^���5�9��i��Ӏ�r��H6��1�i?�����ʢln���d�zxp�N�qM����mS��Ѧ^a�"���:�pD���yGjhh����5��ܠ���裏>"c+8��⎀�����Ύ����S[Mۧ����C�[�����,��00��'P��yPP��	k>���a݁2��B�{���'���~"3�E���昺[�mj�ooo��۷L�<11fE��B�$��t��E�3,�,�ۣ�����l��.���Ta<W�5's�s�)g�Ïɺ��BI�z��P��>kG���{8?l�0Ƣ�l��"~��>碶%A���³�N.
@b܅k�l�} ?O�>e`%3&j�F���:+�Δ������;�d	˦t�Zp�~������^���WJ�:R�u݁cӒ羿��z��Y+$���q} �bWI�% +�,#k1J\�*����L_��Y|F���A��⥋�сn>�wmmA���;YL�zХe�{�j��E�p�}�=�����Ҕ�2"{�Of'�Y����5��p�������1�gu����{��`���/�l���L�h�_'PL8�1����0�f` ׊���V,*��D�6 l��^V�Rz��LQ�`Cn���	��@&��"�rAMb�c'N��~���~�,"0�qO`*c��@�WȞ�dTi��X��^����HS�eP�ny��/��;[�P�1 ��sF �ĉ��8ֵ\����b�# �h����ML��Ō5��� `�I��0��aP�q��_�{c6�?ΰ�/+Ě
[d~�9������v�A� �֍ D�m��m�E뻚!�4ۄ�5��@�o�/U�ki��������^��?�ipX��,�t�i`�'�������, �<1&��*RX���Τ���/�òr������5y�O5��6B�N���㵙-��pYXs;Vw$JL����C)�׾1��;�Li���V�ſ;毴�P��j������~vid����|P����fa��d.�I.jֱXM��^ �_���}�`��uF��4�F�������;R'���ޮi�y&t`*GA/�f�1
�)�.D}Y�݊#�,�i�)w���n	�����d�2�ҡA��-�~��<y�L�nygMS�^��Nvw�nī�, =���ڔL!w���!0|kVH�E�̫+��hi��8����V���A�>��������p�=q�٫ a��%Ȍ"{*G���'�t��U:7���r��^y���i
Th�߻M��M�p�p�*w�=��N%�)��0���m�����Ҕ�Mi9e��1��=�`�����'����LΞ=*�c�������ϼ�{>"o�u�R�3�)�es{�Ny��T�B����^���gt`�9}���K��;�{�|}��m����o��*4����NP$ul|�N�fӴ��C�z:���y޶bG�idTRf�ʝ8>g`bpx�m�o�Lc�����0t襠3֡aFG�Uͯ�`m��X K#��I�w����	�\���Ay��|������������b�Ve;��]�U����9�8�,�a �0^ �B�
����G��g��%�d���4�L�8���!.��{�1�0_��Fܱ#��T#�� �m�7�MY�ȠNz�7j��&���A�pL0�8A�E�J��z���"������5�{)����-=gW�%����
T6֣3� �xJ�?qs`��h ͞c��͢��붫
��9�I�D@�gv��_W�����2�"fFp�Y�G�y��#�]�w92���n'�a�a-� ���РZ�@k�	h:��!p?��k��ꚱ43��߯ݣhm|Q�|G�8A�lm��ﾻ&׾��{@�ZM� w�V'��{"�?]O��/n����z�M� ��|���V7oݖ�~���X�ё!Jlom��sg%3���dΥ��Fi-�A kA֬�#��`i�x-~�kɸ�D<�V��
��vul��@�����.l
�1�VWW��b��V���������!C޶�4��k�)k5>��)E� ?{�����?��!�`h�7�l��m�v�m���Aj�9�s���5yvv�l_�|��F�F 0��04CJP�slm��2�~Y�é��	���A�R8e�6ֹ���׏L���-O�=�׸��{q��Q�O~F��-�	�݀V6m_��cd��Dk���3����H�0�1}>#a����sv<S ����h)�e~���;�1ӈ�ln����>�j'��3�a@�2B��`���g(�d�(˟e��a;l?�֏��#�����7Z�"�x
��~��Ri[���I�E�TƲT)v����~M�	,��#e�P�!7���*�F��Y�:����"f����#�;8j�)�E�r�R�D��"�
�		#�1:�R���67��Nhmj�<
��4h��yl�SG��*?+��Q]Wi,��I�j`ha���e,/Z?r�Q��bK�ܞ�H�� ))�p��׼c- ��7��`v��1�u[7��}�Mq��i��T�.2X&��Rpn�� sc�;:M�� @�r]7]Ƃ�(��8['O�`�*�$ ��7�~|o����_��#׉TI8g��><J����y^pLƼc�c�,5�S-��Zes���1������kP�׎��C�X���ݣ�+p�w�}���_~y���Ϟ/S'��w���w��/��p�yB�ڠl���Κ�J�t`7��
����Z�du����C
�XU ���r� ���T�q0��t
��lCA��!g&J�%;�k�3�;����}Nt����n<s-^��oQ�N`��ϋ�ø���#�=�C�?��,�>��l+W�vs�)�e��d�@����kKG�w�Ū� ]0�1�x���#
��1��lΧTle� E��<�VFq+��x,���/I����+���ܿKF£�>�87�G2��E�X��_Ҽ�V@���u���g����l���0����/����Pv������20|�� f���A���յ5��={�LǍM�� hT*��'M���;h2Gm��8`,���p}�,��x�kLOJ��?����ۗ����'��n?��`�&�ȹQ�����9�( )�A�A�5Tؘ,+����R�o�Eۢ��2x�m�L�ϷgZP���mʖ(x���62��	�e��u,v�� Ǆ�L�.�u"I&�aE"Ë2O~L2SǊ��f�7]; ��˿�݀�c�Vh\�xQ���������c���̤µOMM�;��2�p���bv[�d>�8`�n��.�L�>7� e�����n��:����E�ndd\%� �`{�fh8�����u�v��d��,3�cn3���m�e
���(�f���B� ����u���H^������{r���.#`�@3΅�1��fӲ��]1��T���W ��b�K������F&��ԩ3f�} � �7M�{A���PH���>x�̂Tc���6u��I茕�;���=c����L�������:K���~R�į�:s���{��r�d=�c׹^�<|Ce�v0���˺ռ�G\(�'oL{#�e��<����'Z�Ϫ�����Uʪ�O8uHԨ�,�Q��2I?�m�z7���RK���bF��S�#s�0���\���}��M�Æ��Y�-�h@2�ef�$����±��7� 0��L����絲r���	�����r��=������&&�e�){N��!�pY�k�~��V�ipPu��,��C�	��G���&Y�ΊVCoZ��̀ʐ���������[�������F�*�@�p,p=���"���`.�:}�ɐ��-�G�����(�?,d��,1�^�}�5����&pMp`�d�l�}�2��&�h����B4|��igr�ά|��Y]Q٤V�{K�����ޑK���Y��FA ���`)���i]__aw�)4A���>�X���S��9�kF�*�Jh-�9��֪�_��Y�3O�\Y� k5]w���Eh;�J��ރ��i�uC
;�UǊ�ᙁ!�:�k�)�2h���
��D��]���҉E�����r��1�x�d�h�U$�e�S.�[\Um��R���(��j��e��27;�q�B�:���]I H���*S9�K2Ώ�y�t�!5��փ�,�r��5gTv��A���υ�C����
���ĚP	 $�𔭉�f�Ybפw���$�	]��z�Vү� @��������M�ə\���O���Ul� ����l ��ٹ9�8(�Uob�P�& ��K]� �AR�k@�n������%
vV0�����u�܍:�~-;}�4S�!������rȄ�ܴ�����R�y��o��/��e�j�����[���~)�N��kSC�v-�m�T��벨��<�q ���{�O Hx�q��l��5 ����.��y�i�I%��u� �fma�Lb"�u�*-`����\�1ٲ�*�ᡘ�f3�~����''O�"@�L)����W���kk�� �"��Sh���i�����ŵ1����b��ڏ�8.��.e)��AA��(
��Z��f�]ah��F�}�����ue�/Cᜰ;`�P��7�eg��Z΢��BG+�.l��Ggp���``�(u��SdU�6[ԕ^\���bǡ�<þ�={���s¶�=g�.�9��ؕtI�j�X�Ae/Zme8�,xH�IcR�ÿ��nE]���q�����fݤ(��Z�E��ia,�]���^t���Iu)�Kq-v.J�am	�K؍�>�1����`�ދ�
ޗ�Uغ�^ݛS,���ح�-T�^������3�M'�S4(�~��9N����Kŵǌf�Y�P�'a:w����ϵ����jy��
��)`Et���<�2nf��nJ.GxX^8�\��݆x�y���^~��"�c�j��)�4"�٨�A�Ӫ�)c[xu���jy�tܘ"��qQt����O��|����3ձ��v��m:�AC<0��R��0G��ÿ{NakXY���*�7�d ���A����O�FnE���	�f�
���S��7�O��E� !qNh����y��5���ǻ?��mG�Xu���t��&��P	���yD�'�\ �F(�RP��V�BM�_o���_�
JA��;91EF�J5���Uۇ�;UW�>XҸ�S'O�{�`z(�2�㺶��>Fѝݝ����w�����;�����#��y'yU�^�T�ސ�7�������et���_'��I��rٮm�nm��%g�!�pvvNZ�u�G�����\������"O?��wᭋ����;������D�e4`�fQCc6#��V�	2��1M��:���FР�l��U��Q\��b��yg~�N6�����G���u{{ל0��+�#!@X�q���;w�����˗Y��J���6cc6�RQ%0^����*�Z���|�w�.Zu��)��,��ĕ�YiW�!#���A��ܹ3d+c}A
s�AKƑ��Jy*�>�,�r�<^�x��BM��&CZ���<[7<�-�|���wrc���艶��ˈxZ/�����M�����w��&���l�����-<Cg�}����Lv|�>y�XN�5���S\[&���AR?`Abx!h�e(jձL�-�\L�6cQ=g����h]�af��pyqq� ��SY��=��F���o:Y��M3�t�3����Ϩ5��s�c(vv�A9���I�֏~��볦�!�v7�����u�~ox4�H�߻�̒����f ����X��I ��ڍt�4�3����NF�Q��s�_4u�S
.�4�����N3@�A��ac�28������7�ה�@��+�����{2���r�
�:�(��)O�����q����)j��c��[�G~�˿��t��qJ�`�mm�Swz����������|�����O.Ｃ�Y�3S:Oi��p�"[{>�;�H-
�p�@yI���F��5r]�)/����� м��ʾD�]�x^6��ȃ���=ږE�W,H��o���%,�H�k�B���wc��E�m�h[�{	솎�3m�o���?����;�(sv��օ</$Ep� ���p� 3�N)+�v���B�`j��C��P-|�����-��E	�6�Bw�\s���͒�:l?^$��̉.[�,{�|�����*i��}�o�U�u�ӞVv�����y��y�UT����5'~f� ��s������9e]@��}�H���v�����^Ʋ�ɫ��t}� r�����?x�v���j��dȔa�#�b,c�(f��t���1����T�*�L
�ϒ��QoY\�o����i��:%^$��)Z\��[�o˝���a�$�|!R�wH��{�U�z�>392j�{a�n��]Д�����\D(4���� ���!�� ��q9���?sdF&���^x�<Yd�<D�i�d�*� zh1;0��d��p��u}}C5��t��=� ~'O�='�V�9�������Y�^]��d��}��d\��Y�D�� ��~;����u�;<�5�{�������|�@R ��5����ݽwG���Uϭȹ�����I����>(�6�,�d�C'y��K%��u��`fdaaӺ��=� ��I|���@X�7Ӑ��X*�t����̇qV׎��X�f����w���p���x�,�� �/q}Ԯ�����X�W�����I�R�K+�<��x�b��4�Z�ې.�b���8��:2-�B��px��`j�@���(�,YBM � <�z���Ӕ�Ǿqqo�rp�Մ)��2CL�M6F�B�{�Yg�`,�7��yz-�ӡ�SŐ665�� ����&�������J`���+ۦ/�u�+8��������^��`=}P9���YI�k,����u���=6j� Hb�C|�,��A��A�1��L���^�,0��eV�c�Ŕ��@;�1c�ާ� � ���M�ۤvw�u��1F�ԛ�r�gq/ ?��s9}挌M�������S�)_�ue��+q�T�T�V;�nݺE��� rc��j
B��� �i�� mY����;���4{��L(��j��i�I��;�;|^|�,dQ!��u�{��\��Q���[�R��P�
���-,�Ql,���j�?z��`!�;�7�HV5������<�7o^����Y`p~J��xf�y���D�X�X�t�w�� ��`N �CQb������р�h� �aΣ���fd�����g��[q�,��m0��ڹ����{1��i��l-|9����9jE� m�^Z}������>⚮K'�yQv���j�;��Ǵ+p��l��c�0��t�����k�Ag��(��pӂs�4�5�#�6ޘY��-���j$�A�jj[�ԡ������j�|2��-8��'�B����`O�r��|���W|���2������rR��%��D�&�'ޔ�F �hJU���$�B�  -�D�!Z��U���Q��}����w�����s}+�������,Hu�j�!FX��ֻ��>kFi��RRTp~̰H�e��i����e��,�*�W�� 6���a��a��Z��DGX�0��T;Qv��¢ܸq�Uʑ�)��q�T���T ����O>��	�L{�N�D6��Q ;d��T�Zú6[K�)MKO��� �ܩ�):$86�B`�����_Q�pjrB�=B�L��Ǐ�%�	���Sc��0�@������lI0����"�z���Hu���|�U��g����ѱq:�b�M N�����A+>�֠���`P#��A�jLV��������7nʵ���� �;>1�8�xm�Ln e�����.���/�g/����W���ݼC:&'O�x]�f�ll�'�b8�p�pms�ϩM����pF�b��U�&Ƞ8_o:|�@ e3�u�1��:0���r'����Q�1 �t��٦v3�c!�^,��#��PlŐ��%�A�6����%t�0�t�A�"%�ʕo��?���q^���ZRJ�s�qK�}�0�w_{�u��q��ǹ(��l ���ܽ'��ާ��� �R�=��Yd��{q��? �� P�	@���V; F�.�c�&E��Wiq���3�� �ܑ����I]h0�;�~� ļ���/�l綛�`O�U�}�a�����>�\X�~�孷��}�bz?� �v
�X�i�=3H�@�zmu��*��[ �bt�*#;z�(��}�
�阢s$U���kz�1͑*\\rZd��8�}4+�Z,M�p��8��t��}N�UY��R#��ͬ��e�`=C��?��/��;�)�����\�Z˄�\joB��oҰ�c-�	�,����=kОa������`g�1�g���"2�X�΂�����E��쬲�;=W��]�i��1�ZX\�Flw6�^��'b��,AΠ6�0`,�����w�~�6�SH�`����^����{�0xE����4��I�;Zlx�ckiq�Ņ!��En[khf���r���}�揻���lW>���Ң��ͷ'R��լ����q����i��߶�� c��ڐ�֎&n�K�.�Z0'�92 �Ν�M�#p��$��1o�P��7���N�����Y,�^��e�1d�yM��I���-�3Ep d��� `�N��)a�����
�Z�1�������G8��ƺ��$8�k�%�"����pCfa�� >����lfaL��L	*��e����<ĕ�����:��������}��d ������L����[� �{��U�ս��}A垳�*���o猜c�윖����,�1�r`6��Hn�b`��i�%�q
��KSoJfB�y��$�}��f1��]�Jٵ`��]\@�k���/,
��E�JL��]_s���lA�:�� 5��U#��\��Eb�hs��-�C�k�����k� t�f��̩�=V���W ;�~�L�p �Ϟ=��q��=�,�Dʠ%i�{�)Z�M��0�F�ȾPFi�z`��0��0d8U�p����z0��X��jue���$1��nic}��k����1P��>���|J�z�.��z� c�@�}��13��dmø�#��Rgř����:�/��c'Dْ���/y��8~�� G��deyM������ӧOd����c�nܸIq������Cv(ԃb7 �YN�@�)՟~����w��=0���8���s�����Ȁ�e}m�?��dc��n��h�9ˋ�2�h��p�����3
��{��#�;dԴ�N���2�Ŷ\�z����Ξ��0岍j��]�.*���6�&0�px�+�i��D�ـw|
e�� 4��s���C]`W��t`�
y���3��ܑ���,�������:���аlB��4s\���򏬦:�N�F��ְ��MV��q��z� L��0;Q��a�9l�֗Y+]s�Tu��D/�l9ȼ~������-E�d���z�
R���V��A�3gNT�MT`m)5W���8�~��J���n�$',���k~�@� ���`
 %:��x��x�#�j8�����K�z�NI�Sm��E�@�*y�?�#��s/�T���Z�qR����^�  �<y�}��E�/�8��~܀%��4�fE���T�_oI��%�z$8�qT��I,�lD0Tq����.��g~�� U������Ҡ
k�����  4�����3��ܼuӯ�����2��t##˲͵�����'���h/r���cwK��F� ��|ݸq]VW�9s�$ԍ�V2 K���\B�Y���S(�d�+h�C����D��D\�o4�wS��>
�v,�����p���(֐z�ބ=듏?�ߗ!�t��?���]'�999��c���|��/�S2AT�-1���,-�;��<@ٖJ��$�|��}Ϋ��P%������G��>|�Pn޸Ō���Qo��r�|�"�(:@���v��ZشŤ�,�4V�)���]��'�0�vX��]GffX��)�Ϟ5df��a3Z�Yc`O�~�視p���ZAs�&���'��b@���� }��F�L��7d�a-�5�;2�vw�	��\)!�.w��0����G���Wx|�R�i�R�qx�,V�EY7d�E�v2��a�>��<V ��\��8T���*"E��J�?y���[�g*- �b�ݘQU�V�2�����=�#�t����[$%�޺���wgvz��ߝ�e���v���JU��$�@�č̌c�=3�H$@��(��K �Df~�={��12G��3�� ��x3'�4&VYY���$�P��k���kM��#�R�w�*4_=�zbR�����[~�eW���̵�#b)��li=�������|��sdΞd5�6X�yX�śo����}iu������������D��t�k�r�����5����3�FQ�wWvofz7z���=�'�t����_�-]ҁ5(�����rpf�Y%UvC�U�G�p�k��.�Yc�[�� �a���B�8�މ��T�N�4#�R(������8 ���j�?��x | x������ݻ|+}��9 K.�/]�# ���C�&�@v\;��.�C���L8eH���6���]�w@�&ޏ`؃�y,8P3�����$ ��&��Q�=$W����57	M�p�`jBV�0�<~���_��=~�D��2j�=)�`��>B�N+�@�[+�����[[[�y��:���)� �C}p0�"9��B�19h3^��ipF/1��� l��� �Dy�EքU*�FR8�8>�q&��^Ԓ���`�{�|W5|�J�?̂��Gvy��7���GQ���?���t -Т��4q�	�u�=�C����}�]�J}m�`��	������� �>���tR�a�Ӵ�d��=m�?�o�:�Ff\p��@)��㖂~EaiB5�Dw1h[�=��ZG ��VFV~�l�7@�.[2.�1����*˱�< ���B]*�U���{���g:�1�|��Ҩ�an_�[�bj���_��T��^��W��D����='��zmz 9 τMh�O�]��E��z79�T��CT��qݾ�l��%�4�ˊ�_Z�D61�A��.��QZ�δw�h2��EQ��������#��ͯ$���w�녻*&Q�;���r���ן�\9�ƴ��}�Jʕa��o��3� �S���"�*�% �7Vg�jR-�k�j>�/��DY��<y.��,v��F�#�S3�eLJ���w�O�Z����*��j�)�s?}��?��ɰ�@?7�R����lA�}��6�3->��m����Y��
�ް�/�6(v�,d?M�^��p�X�����{V�c0��8���c��S���!�ZHpxO��# ��N�Lӆ�	�2T%@�j��\��Ң�õ������3�p�$�]��j�&�0ʩ����c���\�X,�sR�j4���ryi�|i5����oRIͶ��خ��}C2�^��o8V�������\�zl�q�n���Ap}��"�֖�I�5�N^���ӵz��$|��8�գ��tgy�6��[�ٚ?�k#�Ǽ^�m��l6����]�3��"�xk�8l?}�Mϟ��W��5�H��H�󌊊�0���d?W��M��
����l��~��FAسˏ\�б�>��B�u��@�׹֋v�~�&���4[&_8<?���[~�*@ɬ��H]0�G>]�l=s����89����R����m�`m��[Ύ�(�1��@J@۰yq\��"�h �`���2�!��٧�Q3��op���v��[���}B�@tz!� �%�?d&MO�./��WV�34ł4�ӳ���:�Z��W8<kk�n/��^��!t�?���x�������\�W�
���ଢO���Kg6 ���p��1�����Z���Aoe*S�
�:��J��0$��
���S�c>~�~��_����WRx�@�Am��$s�R�~J�:Z`����F���C��cS�(��a�Xu^����nܩ��� z2  �U�H��v���m��s���	�q�+���{�:��0ۧ3 ��X�m�0��e�$�RL4����������=?/������V��ʑ�'΍��U������LV���9�(v���S�����-�&�i�:��i���1���|��?
lv�j=��A�`���i|�y!ū����.k8��X9א�J,�Ñ)�B��^h!�F�v�UV֮�o���u�/�T�'�D0� fu�q:p"A�Tc,	8|���l�	�����H}�7{��4��ֽ�W�2���7_�5������H�h���Gy|+ §O��2�2J ��xƸ'`j�]�JƠ*�cD����3�^�,)s�m]��dÒk֓���/1?�iTc�� N�	�
��Z������%pᵈ_�W�,�%>V�����T�k!�#�$�K�GpXK�� �[�w87���>�4|}�n޺�����+�F�kЋ~l��PG����T�}ȐI��*�q�rZ��Р�d�e���j.5L^�b��4����B�{������0�\���- g0_��}�
N�G��!�{e�b��u���e�W�) i�5�=X�K���5���`;����8�`z웜��;6��>$A�EM�:2h	�3*"i��@x���1��m��Q�t�5��snqi�Ǆ\	�+@,M�-���p�3��R�O;�1�m���p�~?w�+nw����^ �O�D���Y;��7��)��7a��<���������s��Wk�ź����v���8r�k��CUǽ���5�Oj���d*�˵Wm4�K�����>��X�C�̂KK%�z:`�%�����؎?�RC��տ�`��+�1��ж�ƀ⥀�����H��k����{�E;�M��ڈ�C8m(�����C�
	Pc�����[*d�Ep�Y4�){�B^�. @,@O/1�	ihp�
e�dy��
���
���Y�?�W�y���o�Y8#�UF��7�0��@D�= DTm���1N�����a��A�(�Q�\��/ �_��+Jn��B�a���d�BR��o���{��Ipp�?���Օuw��-��_�����j�HP����^�<t���s�Qx��;j�����fV�k�2?�����p��x
@�0�f����
����$�+Xy=Ϳ�@��}x���p�)w磏ݽ{�ý�c�C���X �l*HX����v`^�g
c':��6|�`� i��KJ[�����}��]����VV7��P����O>���#�����rN��'^R@��&��N;�����������߿G��ƍ(��R��$3js���8��n�@����3�B� �!)���cj�͏����F��RS��������C`L?ꢦn~f��^�����kBs̼�lG�<ճ�����A�"ӣ��vȩ�e$;�mjvI�|<�w���gYH� ۀ�S��vh�]��$�&uW�%J�Z���L�����ݗ_~���F�ȶ�����Z��;b��XS�ǂr̄	k���FX��s�t;"$@�꾪�eJOEy=R�F=��W�b�\����UO�<k���C�m��=�dQ�ɏ�c� ��g��(-��X�!�,�8��0k�$"$æ��F���A2)�(fJ��j���`���hc���1h8�����I ����ng[�X�{�V����'��{�'}!�D2�"X.��DxHx�潽Qq�ss3�F@�u�X��Vm*����|+[ va�0hS��d�c8����J�t �=�?@�E�r����/qZW����>�&�|�`�>z���1��<%�+ww��a݌��;�`po ��k/��}�`B����A�v_��
�wf��b���dV��l�*m�����u;,�!���ԑ�Z eLh�d˘�s8p�.l�)JZ���|�:����YUQ's�Cm�>l��Ȣ�Z��oEIG�l�*ݻc�\���5�Z��a�������{#�YZ�m`n����'t1h];�����c�r�=�Zu�na���N*��n��I=�g߮�^�^�	UP����75��W�O�t�:��OHGx���X��zNZdN���";��dc3���p�܋vn���bD�v���*��@��@[�X$ecn��.�M�z��|_'�����Cn��i�0�ᔀ�+���R<���2'Y�Ñ�M-ƭ`{�NNe;� ������7�?��)��UF�;�WJ��=2�q�`u �C׆�J��0�/�R�;tt��\��n!|����ߺ��?\> Ci�{LX��1�����-~G
�nb�]�z=8���q~��$]�-��͗[LQKN���4�����dq��Z��ҝ$����B?"���۷��fq"M�miZk�qR�0�¹�l%�:����W���X�q/�W��pdq��E�Y�70�+V8mTI�D�N�lUK��1��r �|���}*�wj��>��3��������_�^5�#��ߤ�{[�3��3�Rs�o�8c����|�m8�\��I^��[K�f���cΊs����#h�M�qW����E@��W#���ڿ�nA#{��b]x��0 ���U&ţWrµW��ѩ�C����ϲ��o3eY��b��8�1�y����l���k~�)4���� C6�̭þ���Z�lH5U�p����J!��g(���ކ����1���[�<(��"�Cu�]o-[��������[��WV���bm�PG��0_ �a��G H�r�iX��O������*�W� e�:�:��0߰�67���������5-�,��?T����Rf�(��뺃���u0-8@׊�Eg�W�8���s?)2�Q�`�H�u$�}2�t�Y�q_`=#�`(������ ��y/E
��*-6�Xߥ�l���A��t5���V�خXn ��1�/�(�7�E�k��4��,,�㱰�Ycyg
z�壟�|u8�ԡh�C{-λ���6�����g����FEh+���)q����U�)SY���>��ɵ�N��G,ը�8��!�5�����E��$��d?em����.4�d~��6��.#������@��%���@�e.hp��w��\Ƨ�l��c	��^�b�_���8.���R��E��Zďm� p}����@Go����&�$*ʐ������ɍ�Z۾A��2��h+��v����+`9nD���\,�p���'��#)�g8�ǳ��q3$Mgg��ݯ��8#�]����H�Zca�-I-�M���IQ�R��RS�*�f|3��:�D��>�^�b��!;�g,#��̽��x�(��)(�Q�*�K ���{����o���ݽ�4�+���1�S��LM���^�J y� �>��\���Y\;��("'��?dZ����O�㟨�F�1�6C�>8p� ��u�>�����o�� ���gk���B:%t����=~���e0Ľ�� �6\3u����` 4��)ٙ����D
)��&��\q���o��N�!�-�OBn]�*B��n����8�������p� �������PSM���N6�@HME_
۸ЂI�+y=L;�u��"8�BL��������CQ-a�-�g�Df��~�w��:SpXo޺��]��N��[tV�ڌ2ʵ���0���O�3ً7o^c�0�Sn�o�	�Rk�
�*V��ew=����ko����sљ������1���#X>��#�� ��;��|�N�|�Q"�H�y���v�,��|�����;1Pi�Q�ԙ�s����#��1��G�*O����<����ѷ�ܶ~����ck��ËN�x�Nq�{̵�ݍ�ꆱ�q��k�6����$�4N��_DҁI�C�0t@�����!�t�������8�h�v�A��=V�a�NV��ߑ5GPegvv��:�=  3'	�ι��	f[��m�o&��%�	�w�z0�1W�| ֤�l
öpR.%�1�VvG��V�P��۲�\	���a�����@I��(L��c��� E���������������f��ξC��;��v�T�|\���|�5V��.�c��T�2��5��Z^�Hi�,5�Yam��$`O�}��}O�i���}�Z����G��y�kQݼV(PS��Q�$ �#���`	K�#J�!�����d ��`
4��,���������gV�C싾�E�? ��8���<:]>s�m��I�D�-��X�EE�h$H�FI��)�,�(c���e�׏���@��7��4���pQ��hm�%[�2�j�騉�N, ��i5��91�o�iY�����?_aG��X�px��{,;5�q�҆�:��8U}$_4�)�Y�Ms6)G1�ҏ�<�R��;�~IPY7l����Z�c��W�(һ4\�s�J��:"�o�l@���ȼ�zI')�σ>�L�W?W��aƪә�;�9|y����H(Qr ں�a�,�$�"��� ¦�`�z�d���T�����&p١����3������H���D�� �`me8~p�~	���2�]T��L�1t�i�s����z������o(� ����R�'����� f׋��x? �~�'�������H�6��M �Q�'W) 8�l��ɖ}Ҕ�D��a���4U8>p�>���w��{j=C��ߥ�3R��Y��ep�$�Ϥ�B��Ip�xPx;@��w�������~���֘2�6�] 뙎��+,���<��.��C��D�R㺠;�Q���?�
�Mt��A1���P3��?w7?���/\fAB0{���~���k����9/�$�J$H�٥8�ʽ�w)�q��[Z���"� N�%��u	JC�N�kCQ
 �g	���{ k	n�f�[����Md�0����۷ns�#��Qۨt��M#���*f,��?�έ�Š������F3�)�:�I���gZOe��+���N��Ar�[�X�עH��#���а��}�C�295M=V4ѽ�ب4��r��8�X�8�!m�kW���c�=~�E �Zʀe3y7�)��e,�l��l�{R��.A��?��k3Pb�?�)��2���zRcVU��>b�d��	� 9�ݻ��'n��%Q�!s�����ۘ�R\�H������=etVE��e$�^�F�g�򹱈��u]m�Z��t�۬#�ss��\��v\�J�-`�����y�v���Z{�	!A�,S�| �.�mѭ��W�F�v`��������K~}��\� 2��5`]붻������5-�g�7h���ߊ���E=�$�T�$�>˚��>�냍[ �f<C����>�m����ǽw�@o�E}?z�u�iHeC_"��ʕ�a^e�^�i����0>�	�aെ��,_(2�חs�o�weP��%VTj2'�׊���u��w�¾���Q4�Z��i�`kP.� ƃ} Y��JfG������0�Z��: �S.�L�fU�Di�S������Or��u'�H�x9�
K8���E�h���~��>pT��iFrE��3�[�����5d�0�lE�ޥU���r|�\m����tTj$5n��l ��79a��s�6.�3���΄�9~��H�*_ݟ���e�!Z��pD Ѧ�)�sp`��H���#�� ��0R��Tx���,M2m5�s�X�ksʣvb*� �R��[W�5��4=a�`�B��޽{�O������	��h�3l����`nk5\ ��:d��_��� �͛7ɂ�9�g��o�!��|B&���h=| ��؅!��B�H������	G�s���N �*h%�	�~ ��LI-�cz���*Re������Yo�8.�������/�W��+L?K�,�%gF���c�1�1��,;t����������oݧ�΅���=|���,+���Z�1
��8�it�D6A�K5ݖ`N�<O8�&��� �(��t0��}�#w�����O��!��ti!<{0�|�Z���x���0.�0��s�`�>sw����:�	!(�orIZ��+ZAP��|�j��T�KCӘ`;+�+���Gi��dK	�}Y�nFIQ���� K33, E�hZ��@�ܸ��~��&�f+�i��x�[�R�ϕV�X�.�T��p/�d������}���ʸ��3'?l9n�`�@�4��O}�������~Xs���>�#�%d�+�2Wp�h���gr�p9�9��߸~��r6��yל+��%������\�K8ǋ���G���g��(��\���Ed����:�^��|���OlnQ��=<p�am���Һ �*���J>C�UAX�ǅ�G�gP$��뚔B�-c4�Ip��.��h�ZQn��:��`�X��$iѾ�~��	٦C������#�ո7�k�}��`8�_]�L`�hn��1 U�O����/d��^" 73=�&�=�W�� �(3�X�NnE�7�3�#>�1� Hc�������`
�/�K�Ym� za?!�H��p�7M߄�#�z�5�sz;ؤ诵�U795�L��́���(`��~��V�(@B�?����zb�lR!qC�d���0��QU��� Χ-�n�l����C�����*\���c��<���-��(RZy��n��9'�-Z̰r���/j��LO	�>���N��Ůu��V �E;���캶k��ؠb����r�얋v�N��q������*�b�=��e5�}n��R�6�#��P<�z!�y�۴=h�D�4�k�ޕ�� ��f���u�dyM��x6�����j#����|�����\Y�[�]뷋�n75ah�L��4b8npdȾb�\��h`�Z�?�����	V�#k�U-S� �+`�s��U�SBѐrC\���n/���:e(�&f �?�Rp~ ��ۿ�����(�C43;+�y�� /h��n*�d `��V�4�M�R�^0�¸��+W���7� m�o�'O�Eg1M�4zϨ�X���y��{�Ч}�=Ad��/8Tp� �#RΪ�7�V!R ��۷DW���m��
p(��w$|�賫W��ܠT
��#���;�x�;�`s� ��QwP����W.�Q0��N���/?w_���GW(��+ri"�j��>�̩U	�v�U�5Ŷ�#,(�����G�P��g��RtQ8�`5M���B�b��e�����S�0$P��
�;�%���y�����v����nݺŴu��	��%x����9�ͺ����v��?�z=j'�$ �˫*�1s�se�Wz�y������D_�x���z�Y�[ �S3D#u��}��@C�[XGp]H�F!-��ѧ|�x�δC}�C��ӱ��w����k}vLQ�u`���g�]��,|�)c�ʴ�9�=b~��z�{��k3�����`?���G�y��8Ο�J;|�ؓ��5�1r��d°���b�w�ޥ�׸��`�e�	���UD[�
������q��K��k�
�3@e�`<{�\���8�N�ڿ���s������)�C@��s����hQz��2��:*�
-�l��\}�a�\�~� �-����E�/>#K����X�w��c�:(Kģ�Dp�� �����K�P���y?O[�� -�� ��'����d�a�ԉ�Y2h�[x1� ����8����߹��O���k`$�Y��bW�\�����O��w,��=�N�1���ż2�
Ah  �=~��}����=N�z������$]YY�| �⼐3���n��:�YU�OҤ90�'�l��dA_���h';�1іRr���T��Ƹw
B�4Ϩ3*��nqi�MNO��x	�>0	`p�ʵ`}���Z1&P�6�-
؋r-<�9+! 6�e�$����f1BZ�x��˽�O�8P�z=��#�`��ֶ8�<v|�ߏ�{��Vu��	j�[���,r����<т?��~l{��Jdňa�5:)�~�O���v3��i���W��yPk��6�# {�{
L��w��颽�mL�ɫ^E^����N�Z��Bo�����p6�� X�^�VRp`uVk�]����^+��CB���C'���p3:�S��#P���3j��L��V�E�&8;+�Et3��w3��Rϓ�	�(.�>�}�6+��q]~��=x���Sfѿʂ-k�0�`���O,�L���5y�R����6��=e
�fa���vܸ��kdQ;eL�yA�c��2�C}��3s�{����>8i���\����!��hx�=H����g�pt��ߢ�ף^q��$�D����u�{�08��&#@�$^%ATjB��yN��VʿA3�s�xR$}G�M���.{/�>L�·�����oH����J��`��罁d��
��`�z�p�[-�AWz��'kk�n~~&�^	R��PnM�5�B��O�G~h�sM��
@�ۂI�����^q�GR�#���:aoa��-���� �(�Z�X�_+k��x<���u[��V�Q�Ժ��=�+)!�3��.��j��n�c��3�!�i9��+��(�9��@�\1� ���)�e#�V�b��+��$��ZH�y�t���Z�\�2�-��O܃��06I�S��`��5N
z�o�-�k Q�>}J`�-���JHy3A�V�����h�d�6�u��������u}�����2�OXO�ǜ��u�h�ȸ-�ݠ��&'\G$�_e{���NŌ��P������
�Y0�Р�i*�u[���ߴdȐy?2�9;7��t�u��창=�ᒥSrܮ�x�"�-->YD���wS�q���k��0�C���ۑ�Evv�Gԑ�� ]`���ve�ڭ��)�P2���I��i�;	����X���ֿ �+���z�]ks�K�pϳ�}�u@fM�`}�,�]y��M�5 ���C�E�[P��)����o�p�_�t��a���� �a��ZxIb�&��K�<��v�m��i��R��X�؏�E`Yf�k��Юo�����O��,0�~���h1�B�O
h/5&�f��X�s�$��dzI} |&MD��b�$i�J�ٰ�s��_��Js��٫�ϋ!s���v�}ߏ��l��t�L��m�y�:�X[��X2
�FѨ�Zj��Y@�H_��i�'o���m�����]�󇁽w��3�+~��"��X^�H*�B�J�q�;P�^y�����8i�3D[���h���T���J{&��<�u�q�`����d?�2$XR"30P�Z������:��#������[*=;+>jU��T�H�Y}��]pM�>�ɱRy��e����H�gZ��˴��a����Z5��-�m^dL���B8c0���\�v�ײ������߿�-�dзTE>� ���Tm'g���dƚ���ţĄ�k =bln�� |���Dƭ[7���R�.U&�I���q �����r|�����-���8�q��.��-$d�� �a�B�
�l{{�
է�Ø���9�U ���<i��i�8`J��*ف�y��sV���É����g��P��2���'�lg��ڲF׌/�V���/X�M�D�SI��Y�|(�,\+�F�mmm�'���g�|�`!�����!u�8*Pٻ�Z��M����p��=�?{ƢOܘ�D�s���R��	B��2>{��ejj"�le�����x���A\iڎ��dƜ��TvH) �&`O[�4����UpZ;A�UeQ�����so��LG��1�q�~�'r&�6�o�<�+O'��Z]"/�F��E��Ә6?��wtmC��ڷ��P�	�Ъ��:�D�ca�Zy���yN+�f
�GY~Gx�`i����HTA����1;�N��u���u�����˫��M�K�FG�9�b�ND'�,��!%��0�g�3hl{���2;yFedJTRcp���z?�� 'w�y��J���^p��f�������Gp;��,�0{	�yx���uq�����B�|���dFk���tE�6�י�7J�d�L�51�^%5
��eV�AY���K��	$�0�E�,e�s����}ꝳh^[�������X[���-�ѝ;����~����w���lnnn����0�676(��ޝ`�@BL~|���.�d6Z���� ��aKRB���i�R���~$ud��1$�YJ��"�|d�!I��-cE�V����s3ڄ=�/��'�!�79�ǽ�ٮ�m��ǀ�Fc$0!Ϗ�H�-6&`k5�e�ˮ)i���/ �v��'�&��v��j�Ⱦ"����ǁϣAs�8o��ǈ�w=n<�:QR�()nNP�'�2�L{yL;�<?� ��,;T�L"�	����X�j5���89=�]m`��XVG���%�r���I��"H��x�.�h9�E���-JF{8��@��92 LYd3��p �<�����f�4�zN���SGI�	�lN����p�ә��Ӣ���p~p�`�����b�N�˗R%L�ɉ)V�G��H��i2�|���`_v��+c���� ���8���ئ���?����<y������P��f�8�y5��i������Cj_����e{���������<=;Mg�Np� ��"�݂�jt79�p�_|���o~�.]���9 �%���}c��7-aye�$YU�׋�9�˃�����d��}�LP8`o�<�3mB�V
>��G*��a_?a�����d bS�1�_8� ��ng2��$S�{dV�(�Q*˹c^�<������=(�[
���>Gp'�
��3�=���?ԟ�dI�� ��H�V��:�A�s�Zj�&5F��%,M�S��:��} )�S]��^2��;������(�.a:p�y�UZ�'���1UpAҳ�|������/l�^ $H�iqe���Y�Ύ_:I���� �<�8/�L��Tт�a��#�3 _�u k����(����9���{�yǠ#�MHfO:dV�C�^�J� [C����%c�{NH]Q�>��7;9���מ<}����5� F�&rU�D#)�,���3�=Na�4�ڂ��?������ǏG�p+m)�Vj,V{���l�,�g]d1d�V�
z�2�_�"��z�<JT��	�U�+������`2� F!!{��v`�t�d9�� {���Jt���CrxH۩ם���F�,����z��e�% `�W��w=�K����mA����F*A���� c�R`��
�..lrJ�ε�u����VW�"�vh�������h[��}�������N�R �c�����%��[�5 'ɋ��������@ �I4��ρ�Ni�"���2|�@�,6�6Q�i��Ohĵ������Rߙ�c����]�F���IM�X�S���p{��LF�d.y�L�,��O��?���ꐁ.�z�<�?�^��T�D��!�ي�::N���h\t�hu�.���ky5t���T�m�3��N��q������ظ�:
&3({7I��{�o{/�e�*U���[�6����q�7t#[j|;>6y�v�w�
Y��*x�(X��q�/������v�~�VV�֏�����$������ש5Zv�NQ� m����t
*�B����뙰~R�D��n)-��=�R�88jr��R�����:� 0�ќ�'?Ufm��J8 R����	�KO���`t�ʼ�ۂ����Q�n�z�����n����Dq( ��}�<��={B�`T瞛��� c�.�gV����}�i�dg"29�v3�Sna~�����d����d �Gg8��������u���E
X��}A8cp[i;\�6��������4����@_Qkz�tT��$�'U.Q���N���Ӑ�����s �����s�,2���N�X�Ca�RCPAs�ښ���(���1ӹ��� 4Y=�S����e�}�����2p���0����&����(�`��i��mO�����Ͽt�n~�x���H?rX�d��-�>��0G��9��w}u������8��9�C:}���#�`Opc6̧˗/q.Z�m6PՍ��8a����m�Ӽ�]�Ň9��dx���2�@�\���YDЮ&q痓�f��O��A[+�We�Y6K��}ƴCI����̮	k%�&a��E�6����.ز�9c��:������v��5���ls�z.~؉`L����\]Yu��	�A0c���R��=�x{{Gd��uc�=j���ϩ��}��/�d_����]� I��MML��r����B� ��� ��� ��t��fø֕e%�S���Mu�c�#d)Ќ D[3 p6�%�N���b���F-j��^��k������/�Nca:?�Zr2H�F�SG3Hd�:����>Adg!�+��H& `��'���i��W�4E��y��	m�X��ݝh+�|��ً[7M��؅`V_�v�]�r��|��ҥK����P"x�����;�2���T{{��s��<��/C?.,.h�L%9�L�v���R�t�ĩ�-�ˢ��"�P��\�]�uw4����Zаb%�S
�8Qn�{��
�� KZ�KXL�T����J��N��z�7���^��shm�X�,�Ù��I���s�.���^*���c�^2��_:�Gm�J*��=r\��ۍki�7��2k�ZVĄ�
uu���es�u(�� �^��י�Z�Q���ʀU�n|=�A�c�AY�d�F��"�?�T�E�ho��H��V�8�/�r��Py�9XS����ء~7 ѩVg�u�m���穫Zu�,�FA��̿��_$E���}W&��4��]<��)�z��	�u���akP�t@f�$VIiǱS�Y����
�ӟ�Lg
�^��Gl��W �H��`љT4�&��9�/�����z�ᖖ�4�i�^�Xaf��ёkwO�A,��ܩT����`/�|]�V�Z�i�������Ђ� �6��G����tpD"���33na~���gϨy����BpܮP�p.���7����y�c5F�v����U6,��X�>D�npBsu�,m�6�څ#���M��j8>���y.Ώ���3#�N����Г��{ �gD�EBCdD�Xt�Ms[/��V�f�Q]bХE�}p(�Jq�0���ߒR�m)hVtQ�8��:�ʳg���}��ZZFf}��ژeTc�& ~�w�J[Vf�Kᐧ蜱 �����ܰg�F��f��A�
,���䟘�b0	:�-J��}����O�#+")��	B�N~�zH��25��TL�iCgC�\UЫ	&�W�_��۟�/���^�UVE��t&�Ve�U,_T�*l�>� �x� �P���4��~���L��x��j�Q��@�Xj�j�N��j�7 e�v��qU �@����l�����~�3]��hF;	��!��gn�����y�5�2 �{��{��rM����~u��Sϟ=�W2���{2�a�Cd�zN�vR��Lve�c��4k��Y���i�L)NX����KM� ��p� �(&�Y�C���2� ;WV^�յU�9�� �� Pݡ.f�c�i��`(2_�y^��oib�Y��{��/��2T ����Z}��_R����-p��Y1�`ϠF��om�c����$.v�]��o��pU����Dӓ�e�g?x��բ݆u8	��t����Oݷ�~K���
��XO��IX���L FC�����K��(��`���"���A �k��D�̚B?�܊|I��и��-��)����e�}ۤRT_��o�?�bD��\އ1��+$ �z^$(��ANA�$Itܵ��k�!��>���酲�M���7�$��9{������@����v,8|��{�Tu\ٟ'j^Ge��Y4<��H�y��H[�(�� ��/�������v\{w������s�*K���DC��V�`�d�Y�BQ:�4i�œ��������|d�D�x���ņ{��G��S ������΢\B؀�����V�V�*�6�-ϙ9vոe�G�_8(�+�JR+*Ц���|B*)$8� F�|�?�~�0j��|sc�ƿ��]a'��$5��	���:�{���\J=�OdSƵ4��f��쌛��r�n�t7o]r����p	4�������#�ۉ�K��*h 'Cu^0�P 4 @{��u��_���z�ݽ{_��y|�=@0�p�`�?L?�R
�?~�Ľ�+t�g��Y���u�3��G
�6��	՛&��'�Iw�P�\n�$�Lʢb�n(�+ଃY%}\�������:tdq`���R�4�\�-�x��t�Je�B���}43ͨ<���� �vs�>j���˽���5��q�q���Ls�3&�n�}��~��|Ԥ�93"�ӱ�^�8�����{c��p�� c:�k�iʒ��cAP�Z۽0Y���KB(0�QΉ��5٪u��Sfx�2������OI@c@�`���{}a�F/c6���j�]��lޜ�JN��I�mk�>њ#�N�R20�,+F��*���mDVBam$�A� w��`2;�o��,���y,�U?���@��L�I���(����sw��u�wq�>7��6���|��[�uZ#�<��^����;}���Xc`�@�\��{��+nnn�{(�|5!�q*� �J�u,˚τkR!�~��uQ��w�@��)c�Z5���BI��
�'�w�Pt��^��e��L� ���>�@'rB�;lÞ}�"t'�nRRss���>w�|�jc���	P��ꄽW�$X�B|����X+�0Y\Ǣ[Р|�{�h)j�D ���=^���!3�2��W_q}��\�կ�._�쪛ny��֖ia�PS:I�¾���yf�����<B߶�W� dkq^�P�.M4@�R���qP�2�(W�i��Q>.P����^U�����I����細����Y��$*=U����V���}�(�-b2��8����CI�7Ʋ��^\����K�]t.ڻ�8^}��ȟ��9�_N��s�����v&�B�_���v���1G��X��rN�{[���TSvz�m���.��{,�dn*�E#%Y
�Ul�Y�?�W��!�<*G�q�(Ox휶�_~Y��,%�b�$/�h�GBl�_��gp�ho�@{������e����U/rYgX���u)U`�g�lիm��`��IU�słb�j�a&������Ȩ(��,Wl�N��FG;U���4���mu�^*8��Ca�Z^RK�E(���ĘK¼.\o�K6%�gfw��Tp�z��y�67v�3�uy�+N�0i
-��>��a�2՗
������_�nvv!|��AQ�1o��V@G�88�A�������s�d��ri����_����A0}P������\���T�<�&:u:c�$?)�V+��Ӯ����dLk���%
��x5��<|e�L�+F+���ŉJ�Bβmw��qۻ�tN����4�M��@YRM[���U���6�S��Hd�I� O�(IT����y}�Ed��o�E�w)�Rx��.5��`	��E�-� �����c11�l����ݵb� ���U�\,�6�(/�"վ:�N�T�Z�Ō X�5�S,G���UF{M�uDF%�8[�)[���"��b)�M��/#3�X�1S@��{���~�+j�hc���4��b� q�.�P���o���a��I;aO�����Mjԯq����j����F�פ�J�ݹi~���D��S���V	{����"�=}�v�z[�idy"0Zj��A�*�%{}QpT0P2U*�w�s���\�x�딭!旱X.e*dO+���i����wˮ���� Pa� ��HM����!���>R�xE^8�U���x]�`�!x�~�r�������_�����Ƹ���g�W&R��6����11�	Z	�1l�o���&���i�l�{�̰��W{�{�yأ'��vԒ�����RG��2��#��C�З cA8@�v����M���'I8�b{*�e�j}��`'���K��R��B�{Yl��=�ݰ*p�\���+�b��X��q{f�Rt%3,d�~1 W�Af7�:��]1 ��rIŔjaG�,Ft����\T�oi�E{K�?�%_7�o���q��ٓu����&��^�mGr?�dv.�2��}	u�X#������?�
����}͛K�{,'
rp����$jYhQM3��E�̬L6�/�X5<*�P���w�,�#ժ�~�&��Bug�S~E�ڸ>I{PC��ؓ/���$�T�� 2���ɳ!����a-�":���{y&)@Q���ɂ�E'��Z�F�R�:2m�q�BSQ� �EN���#�����s��"8-2� Ap��݉�$S3�8,f�N�O����`:��X��{3č���eL��1�h��ť77�]�1�������ȶ�8�ep���@��$O<���� �}�B�b;8CK�ڕ���a�>\v�[�!�j�q��~����	;�v�p��l�kmm%|����'s�K����nw��^�x��I����Aȇ-5�&;et�Et��M�Pi���`BO���,������{]2�����tV��2���Q�@rD�B�0Ü�#��=qߵ� �����[���%ѥ,e��aG��9f�0`6�v��N��e&��sG`y��2�~����1ڮ��u�㠮[��g�4�E!)�#���/�����i5���˒r���q̋2�[h^�G&(���� >�2�s>�Mw��`�w����N��e^A�v���&G�~�t괉���v��|��y.s������M��%A��4�P��9�keM��j૔y������g��\�P T�� �S�З�ܯ����Ij{�8�H����gO����� 'dEX+R�xG��;������R��>k@l�x�R;`�nKP5�}��!�>tº���{��o{��}>b� ����I$pE^�^WRc��n*�ǌ���6P��1Y�9D�#�62��{�;,J6��)����yW20�,�{C~�sl,!�
Xd��F�/>��}�����O?�} ���I�	}�@y���E�	� 7��aJ{����t咻~�Af\�)���!��>�5Y!;��`��d[�0O��2�H��op��� }d�a�I)j	 }�,4%2 ����0���յ����^�\�yr_�
����:��l��oپ������ �ŜY���^f��.�aey����8z5*Sy��0��zm*�!�I�͗bÜF��B\^
�ڹlӤ�(�r�#�ƴ/��:�O�Q*H�\�hok/{Z?��O��s,�����G�������Ȃ�B�9"��)�"}=�$�\�;8�:U{w�/��� ���4��WVLc-(d��ǥMݐ�XC�j�EUK{o��Q�G
��������~Ak�͜�bS�how�LIe|�K_�n
ʐq
6gXo�22\�H� K<��!�ûHXد�re��H�<a:����0�2˕5l�~IO��2@�v<Fp�Y\Z$���+�@�L"W��`H��@�8��SS<ϡj
3��Ty+ғj������^���
�
gj�Z�m�0?�������t� ��.#%ʄ�� �㶼����}LMCV�08I+t�?��C@&�%^���vׂ�Gu�,Q�ʀ��>o
�����W���=;���	��"+�l�i�>�<��&*]L�%K��&-:.����w�ً�s��U:�H�}�zS���(d�z��`�)�l��[���U�Pd��|H�i�`D������iw��,%HīN�����xN�H�$��4JeƮ�O`udM��'������jF��(��mt�8�qj[��� u�GK`M��a�����Joݴ]�Ԩ�������W��1L�����T����ޤha�DJ4�K	4@c,QI;�����C����&��_k��k����1?��b�ɝ�k�9�� ]Q֍Ѩ���X�#o����T��͵h.��'�e����Z�B���cuȆ/����Fhڢ���G����m�}-�#�T��zڷ�ٰ��W����x�F�o�����ի7$� ���z���.2�M)/��EmY w6"�]j�$2i�lU�{ZQ^@��V���#���0�&�rܕ1l�@��7�x̀xQIP�f���R�z*���q ����]��ۄj�xۻ;�w��q��������������se�r�/fĮC@��m;f�@&��O�߰7o���FC?/-]���Rǅ���>d��{w���l�C9ke �K�d<����)f�ڤ����a�U�"W	�E��]��{�|����w�᷒��`c��-!��Ő�!D�p�\�b>�\훚�IL`n�<� mX��	��������m,v����.����L�k��f���G�I}�Q	��&�̵T��6N���:��3�҆�ga$2�{EM*Ͻ�fa0_��v�Z&�����9�=���ǃ��7C���~ה��C5�\pN|S��"�w������X6��q�6%6���j�p�1��W:R>��Q����M8���$��f�F�}�����c~�N~�.�/���" 7_n�}��&��#D+xS?�	#'U�8��o{�֔j��ح*1�b'6�:x�B:Z)�T�;~�*ڦR���X� �q<$��L�<Wg���l����K$�a?��N^�_��r�ʺI�I���f�)����u��]JM$I�����/��ƾ�3'8N9��>�C�pp66_J�9\��+�t�>z�>Y�ЂN�a�f�#����|f,��("H6�5�6Y͋�A��PFMG�I-�JEt-N��Y�,&-�E�&�����&U6W�N�>���j ���{da�^�*�8�x/qq�{rСf�8���:�(H�p86�(:������"H]����/^`��ج0�*��t��-u����c:,+)�����.������V��ijfcKT�6[ۀs~;����>>�۠F��D�5���a����a�z�b���v̜�����;�"���D���j�x���:��M�Im��("p�{k:�\�a�r]�ڪ-g	��8�Ys?�Q`��������6_+��v��Ǿ>�xcn�ֻJ���f+)�Ti�@ﵬ�Ty����: �;�8���v��k9��&�$)���/�|����X5��1㱏m�x�(�s#�cc�������є��U� �]��њ=Y����E�pum�r hОfѷ��&k�!�)�X �
 ����|2}d���U2������􌶏���+�2�R���C0wa~���'e0�U��6�T6l��h��� ���9<p�fq�v�?c��6�zd8T���v_��+��,_�|����m�"i��FI@�jM�݄�qX߱?#8����:�h����'�̅}{��3�h^�AB[E�8�3�/	��A�z��5w��������q��`��e�kJ�o��q���9�W
�i�DG[)��� �f�@.v&m
ĬX�`N���B�b(��2�-�7~>ւ%�H�qR��H�kU�#��J#YGkRS�IZr-�[�>W��*�Jd�0��~φ��F�V3�lU��Ջ��v^�q�q��T���>s�8?�Py���L���`-���Ō�*;J�7�*^���=D�^ ��&�D#��JDXu�H��}��RYE��x�c�g,�т8�K�g�`̀.ި��s��b������h�ijF�/�U�����.�
%�r�� ��a���f��_W՘�yS����K�t��0P��W˘��#@
IhO�΢��h����%o89 o���^�^8=���������n~~�}����|���cIjt�<3=ˍ��gq/c����^0�������[��w�}����[t7>�������GO��ʺ��<p[/�ngk@يɉ,c�]�������w��Ҋ����ڠ����٥� ң?�����X������|���.-�)_�# >?9��m�A/���K�/���L-{ �!��2ׇS�MOqL��A��vt�*��J��Wg��}����L1��Lg/�4|P �X����)ʇyŪStX�|Ix��%D� wb��g;8��/�+	����%��gw�À����ݙZ^ie�i���2���-�p������p/�7³��&z3�o��{iU:�؝L�~[*�y���1fbT6G 	�X�HY��'2:���5�d,�:�n�� �E<;�{����8z1c�gD�c�vL[���k�GE�@NR_��z�3� Z�@\GS�+{S��
���83�l���F����^�������y�<�D���U?���㭅2�K�{��!��i�0��*;!��gt}�o����	���X�`�Q�E	�2H
�<�6�+
Y��m�� x�8`B	d�@'�� X贾Ϟ�66��{���L){�B�-��m�܊��ʞ�"����B1N�� )7(�������L�K�`jV����^�[(�ɱ�u?5�EG>UP91]�p,������[���l�g0@+�m�YZ��C�;.��[h�[�	�ʘ��ˍ��C٩nW��Р���`жcf��?���aO���۷yo �i�PN|5l���@%0�)51=#А� H������ L!{֡��F�ӥ�J�G�sE
`�ڎ��E�d�����e2�VV^�FI5P04�,#���N���֙������`�|��r( ����D�� m��9J@1�m:*�{5�-�aNNO�bk��7�ʓ~$��>�2L�Z@O����;n�Ȝ��j��זeh\�=.�1�U�DY. =���L0̇��^��v��+d.j{��L�7�̯��{Sc�}��tU�A<fVh&JS����O6Ѫ�nx�K� ��c3����� ��`����!Zu�:�#��ύ�:�o��7<ꤌ{Y�jw*P�Ƕ�
T�_j}�2L�, �E�'E�  ��IDAT{��c ���yÖ�m���K�l��:�nݛx~U�)ה����QY66'K�`	g�!u�ڒ�����$u���A�eHz�g*'+j;��A�KG*80p�� B��� 4�� �I�@�#�@���K�7�����!@
6uAm�<;������o�͛��������:�)���T�L����
��̓'O�8# . ��C������O>v}�ap����^�L���1����h`1A3%�L�YC�w(��6
���"�43��<���>l���@?J��c�59�&�}	�D6�\��	��vT�Y�X�\��I���<RKRA"�7���Ѿ
��d�������!���w[���]w/�5����C>w��$��>N5�3���x;m�)Ho@b�����3[��v^$���s�蕆��E[�`��5+{�P��>���}��f_I뀭�@ׂR�c��2*��Y��u�bD.�c0���8�&o�5o� H�]�kt�}3�Y���X����+�.Q��9%ɫ��Ɵ�����V��Nm��!�1^�k�ߟ�3(G9��	t:ҟ���	e�^�0����@�M���yWI������^�W��k��>5mY�{�ѴU˴��"Ȭ���V�kR���|�3j�Cgy6�`��X�0���^o� ���fZ�~ [���G,�y\��9S�F�TǠ�%4^n�$0(Y7� Jͤ�j�CRr�Z�����Ǳ���( eUX������k 2�'#h`V�@"�y0�i�j�9�pq���`7��<����5��L�hk6���#�� �ɀ�Ȯ�朱��U�R{���:	�NO;dZ�Ӳ�:ʎ��=���y�}&�����ҝ������/Ť�R?YT�o��v��C-��k (�KAg�[�B���ݤ�(y� 7��uM(4�I
Vg����W��-j�2�I?��}�4��Z�wձj{�;&]Q}�����f�x���H�AM�"iS�X�k�v�=�����ٲ`�\=�J��zs����G~��8�w�����cW���]�?���XN���r�7���5�׊��W��P���ћ�q<��hU{���z�B�qˊ)eQI�^�AbH9D*��(V�;���1�5��!Ǫ�7�J�S�����l�cޢ���6{�~�V���0o`<�1C� �x�f�F 0�cʿo���
M֜f���Z?��O6�Td&�z��4g�p�>�T��`g+8��A�ťwi���Ç�w�����}=��B�Lg���ְ8^Yr�,=�

�H\K�uq�����A�C��f3|r��r}��[�t��Օu��F�9��LWYu9��ѿ�l�����1����@ X
I	8Bw�|�TQ���po��K�ѣ'R�,8��b�"? ]��
�86�qzf�u'�R��h*������wF�v���s8���X_ Q�:�EY�A���up~E�Usr�8�.����
.y/�kN6�QYh�o�τ��Z���U��ʮ�����]ʩ�Zy,H�$U$��ƹ�$[��F��`N����j�����:K��P�P炱���On�\ңư<Ϻ�2
blbM�#��y�g�����<����X���0����.,�� S�����#W�O�FG�!}�Y���y�`ENP��q���k���M,�Z�]O^��'��k��Ɍ;���=~l����Y��Y.�!<���H�5}��~y܋�h�7[���:��N��(e�z����)]Ӑ.����׆@
�}f��1��h�1��}8q��}�+ <�ǬD;Z`�RG(��`=���)o��y�+�# {�Ww���L���11c&�SI���6� ��w��Q�=  -��s�иl7�c��nc��e�ײ��)�1{�c��l`�rS`*c?��ۯ�zy�V�䕬�>�k@���(l�KU�� �B�����be��%@�^O�>@�)ʨϐ� �����Rzm��/�8�޾�q�`M�&��&�0���0$�����U]Y[�w�[�yI@�.���q���a�H�s8Um�Bu�i�eRWv�0 `ʆB��V{�2�S����a�[�U�8,E�����I5���Wc�[捁��l���i��5B&�Ӓ1����]3���}� ʱ�i��(�׌�d�T��5yͲ6���3��{�hoc;sѩ�;��Q��>w�A���!�q�4��[cV�T����!6�$A�	!Q����/'S^��+��{,�U��a�:�����j��IJ��a�����1��|�~�V�9�'L��ఋ~�h�\kL�Q����aBWE��AhL!�ب�K�ɰ�xl��q�b�5 ���hỲ6�ʢ�fјV�S1�#�3ű͔I1��xO0�4�K��i��0��4�m2^q�V�m�*���L'Ն;D�թ,s5rw��g�>��t�z��{nk3	����|��[��Ng�o��^,��9�� P:�yǝNJ#'d:�����Z�&�ӣS���#��b�����0����I�h���={���}�V����)����g���e�A��p�p�p΅�=P�gI���� ��%�c�Byi켜}�8� V�VݣG��:�j��*���S�ϖ`sZi5���%
��a�}������d�M��$���v�;a��'O���w8ܛ�m���M��&&�5jP��o�XJ�6�?��m+ `S���#c�9>�$�>�+�&�-A�{�������έ��:I� ʋ�e�����DB@�E���KV��g���)  s+��0_}�5@��2��!p���܍��ih��j5K	(��D�w�1���G~�m_gkc�r��eI��赞m����ڎK;m������= SP��1\���R6aYF�*3 ���lT&�r����H�U����.�X�81��{�}u�
B���vx�c�2�^SY�9���΃�i2
�@�yj~���9�d�C^$��+��w����@P&2U蘄�v�&��,	��� c���ۺ���� N	�ZF��8y1�XZ�}E �@4�~�Ȋ1�\{� 3�)l�w��4�o�G��a-ʾ YW�`Wtx��j����H����x��Jr!%�-
���ϖ%����10�d�J���d�k�VdRu{����r�l�/�����"����D���~������7;)$f>��XWH�u�����|��u*vm��/)	B�/���c�!3�[��A}ظ|��¥>�Lm�/n)� ,r���{;�-6R-��b���-�ـ����#K-n+�W��V�<)������e*��v��hcږ�j�5`�oW�1w�RlTㆌ��8���N{������O{�����ܶ� ��z�	o7P9il�x��6��_Pf�,_#�T���D����W^�{s]�&�{,K3G%�h���#���g �QW!����c�D���%;�x���4;�8�}�+��E{�Z�&(�0�P�հF�a��&#�Ȁ+�E-��tۜ;n�?�n���7p��l5�@�D������&���\Z$tʺ�cLɗ/7��r������V�V�+�:Px��YJ&28Ax�����da�6�4�KӏU��
�dÂ�H�3���(>���w��U7�ku��[X�p�x�Q�N0�o9qZ��d��B�pqh[�p��ʋ.�E�׺����uevO�[��f����3����<~����>�^r��tc�3�`�0���_4D*Yю���pZ��� �`O�p�>�����";1�{�����-�Y���Dp@)� �=8ك�x�����\�D�5a@�K]F8���}��O�~�������'ܰx��:ţU��`e���^�W�T\1H�@�e�1aŝ�q�eU�+���`-G��I�1#����Dx���=���I�!�?'��EDOk�$����x��f�����p�m4���z�ʱ�
� �(���V$�=�vn_���D/�s�q��R�@��8���ٷ��o�h�1�8H�OR�N�4����:����d��l�x�(�a�c5��קy���ེ��/?眗qk�C�'>�;��~vf���@Ic�'�,X��@��G/�-o���#/*�ll�ڟ��"X��uL�� ؔ`e���:���1D��p�.
�r��b|ȫ�w�����D������y�
7i�D�~ �c��f�)k�i�N�����`�.���"�ZѴa2ɲp2 FC��:�8�Wn�� �ħ�A��1������,���Ks�IS��(���9��U�	 �þ��+<�A3S�p��8a��e���~nE}1��i\O!�������s(@�b��G���+��U�q�V�,@�u%���uƵ�C[׹��yM�����Q�Gi?+��s2f/�h���դ���j�wY6Z�����u�+��*�E?)a"+��њ&�Q
��̲عu#���@��R4�q�^v`�����S���}���}�;�8`��}��{��w�����|���ƺՔ��ߥ>E�5������^�h2P|4���2���Y��i�m�(�p���r�u?�V3ձ{��[,��j]�*:ѩ����t�_��������
�ʄ(N��is�8UYIX�o4LG����B��=��J���E���
�6�͜i��pzG0��N��d,���#������sx(:�<����k��<T}e쳪�yޏ�	��ɖm��
M�M˪�v�i�`���)�sHq �V^�����p�}w��%:� " �q�����w��W+P�1]ju�����凙{��	A7 ո��V�Ky���m���f�½X~�^�<w_󕛚�"��U)���g�,eqv��=���Г��� ��'��+g�X�v����hLfnE	gf��B��8P� �d#8@�\�R-�Y�bѡ6�[�f X?77����o����[��ɣ�g=w��R�bjm�J�"d���n�.�s���RG����K��}�f\�)�s����5�ϛ�꠲?��+�bj���7��{��	��]�j/�Z��eQc ���V?r��O<í�m����>���h��ͩ��O�
���%��T�S��n��:��nY������ŏ�j5�o1��i.���Yg����Z-�>W�aXX��1����f�WP�bG@�I�t��d<�*q���l��2�D����� Q2)؈�hyy٭��P�:&�Rڼ]o3M�pՠ�<3��P�G R�іְ�H]�I�o�����?v\��z�~��_���s�����0�~�= +�F�;���`��+�a b_n��Q]݂�#�������%ڼ��kr���-�O�hWU��@Ke�z�H9TI<?�sm$��)�g�J������inߺ�gI �p�[[;�Bc_Pk�ζ�q�L�`�¶  z��g�U)) ��fP�k^��A_$+ ����X�|}��U d��v�ӧ����;���ӻ�		
!0�[*���cM�Ϥ�`/�e�>}��߿�>���{�&˒�J0�>�Z�V]-��h 3�]�fk�Y�~Z�����f��fc��4Ē ��jYZdUj�޻76�q���Odf	��@ve>qE��Ǐ��h�,ў0J��(F�t{��3^�MD�vf7I�C�_f��t��=>�����)��*eE�S��ѿ(��5��9��G�V��i�|������Tv��r�0�|}�Ѩ4��f� Lj��u��I��*g���M*dK��`k[��rqy�tN��>얋���޽�2;�3�r$��3�۲�����[so���Z;x���~���*A���M��8�H���#�[!��םj�a�A3҄G����y,�������fv�,-ע�S<�^���˝ti�l	�n�9�Ly�s����x/ﲡ�,��}K��d-�А�M���p`�3y�=ٿ���5������7NC� "�cs�Ԇ#�����Sel���� -R:�pP?A�X���TM�2�,8?�8`5�9�CP��'�95�REqp<D�X��n��=H��K����%��q�N�'k��V��ݭ۷9�EgO�(bSu R����; �y�nR�$�Q~�w�u+q�зd����9B*�ի��ȁ���Ջ�$�x�}M�\v<�
܋ni�j�N�^�|�	���k��?8-p�(e��qvz�W�p�M���Z�!�|:�.���ƚ���k�a�v������=�o�7��_�_��ݧ�����Pi�SY�Ixt�vwN�ut���{K,�7G�_��OȀ�g�8��g�,���xNdGEc�V��L(�7I�/8�L-�ȠFp�7�=�8�]�詥�@���\W�~�l��^<���o�D�|'��Ws�����y����M�Ww?�	hM�e��8Vq����!Y��*LW���hC�si�J|.s.���:�>qC�;f����4s�b��͏������a{_�ˁ�#p�z@�z?�}J@s�nZߕ��([O��4���SJL��,�훯�u�ݹ����<����Ӻl?v�)N����ױ�za.�,15`6	�0�x����X@�#���KnX�5j7V�;o6���|��1�a��|�����ݎ�sJNk��ɲc/�$�8l�� �?=+�ڃ&��[Y]a�A��Z��e1����
@��3`������B��ffa^��|�N��1���u��@tN����-���[;��/>g I֬yM��{�V�{���!�r2Uac{�S%��(c6��,�z��~o.I0!�xxx�s��>�4��Ց@0�*��S�i����W�����{]���p�	XW��>$�<PPX�7�y��%�E��; (���1�X��nޢ�BP��� �XV�o�p̕�.rW�!߃�%�dع,����Ȍ]YZ%(�������MR�����}�N�/į�}_�|����܇~�s��G������_��ǏY,�2/��ӓ���J�� oO���5ѥ� }/�z�Li�z��'Z`0�q���)K٣���������̱|2@Z�{�Ts�%8����04×@�������ޗ����7�]g�} ��0�D7��0��א����,.H�	\[wqY2�B4�����x���P9hzc�04�z�����1H�\�v5ژ+�'�����}E��0&H��:��g��Ƽ�6T���o��J���`��Kj�K0�$@\�:��\��K-Ӭ��ZG �]*��xjx���"����0/���=!�3j�)�3����Z��1�l�WO���������8o��c�����Y
v�L���d��3�"P���rlg-~-��r��.9�G�h���e�\��I������<��5u� �Tj���r`6>�S��M�0c�����%Na(?ڟ���ӆ�OO��i�<�T����c������(����xT,��7ޅ_J���e��-i�My�ʜ���bc$��N��� � 7&��C,�u��8�j]S�+z�tlX4�CGLt���N%�W7I�<�3()?}2[�+:�H����䃥ri���P�M�k)���Ud�҉��i�QtY#�i��V@�����&��k�R�j�k��B��A�$V��[<����脂u�sGGR4��d0c��kD��h����2#	�X��B����Ȋ��Ϯ]�DɋgϞ����w��]w�_�O>[w7n�������z��x�"\XX�ױ��bÂ��C�0$������yS��F�g}��d�F ��6���44�U�6<c8���0[��5t����Tx�C�С��-�&�1���It�k2��WEj�bu��\c:��E�z	��BH��[��ݭۗ	P�P�2/N����0e���������Yg죾��t�?( cll�%���<J��y�B6��%�ge���֏8��rS���cD�w�UH�n�X�-3�sWO[�?f��k_�8~��9B�\����.�}IU�7���8ް�d�K�A���J���S��놋���n�P�O���Y�td�s�>���eY��r!`V��j�)�.��29kkkI�����R%�M���p���S'v�����%*o�r�m=�5�d�g	� ��0��<}�>|� "ٯ%Ӱ�1c��X���O���)�E�
�Hut�a�}��{�?�LH�D� ?XˍUj:��k�ї�[>��9��8N���\VJܗ�3�vb��w��7��� S���`9�tE"ɴ��Ɍ}WX���;��&<�{U���!G��r���A
��n	��1���׵��k��##���8f�t�^|"2 <s9���0�Ah�oŽ,e �R,�� y5�����
#�	ʺ��,+W��[����%����7��ٍ���~QP�x�U������DO찮}�(^(Fu*���E�Rpl; ����O���Bp�����Z� ��"9���P%�B�ja�#ߔ�BP����A�ݧ*񏱄�I.����S�H���%B�T���׹�.��������]f)K_���E
ØȾ�L���/9�#rI�#�{W	x%���Ȗ�{p�Z��nd�ƶ�����G5�W���}�~
��/C�J���OM~Y�W��I����6���Ѷ�Z�r��x�O����?e����*}β3��-���,$1&�M0y�ᔛ�)#+?!`yV˓�R�@�+���Mi�뿕p�B�Lz����i���1-<�~�fΧӍ-��=h������u:��ޝv�&M2��[�E��4����g8,re@T�A�{�")] ��dF���%S��`1W���Y\+���'i�]r$Q�^3���
�J�-^�N>����Pa���3��|:YPp)�˩(��zBڋ� ���V�J�x�S]9_l���詗=������;�?��z���V�4����KG��
,�i:73g ��(�6���1u���pxר=-z�����}��c�������q�������'��.�?8�����p�����H�Rg��r>�;�ACǮԔ�ߍ��8�k����� �	!2���MO5����l�C���� ��>A�����^���k`�����q���j�tS����Ҳ�W�ˆk{
�tT��V�K�yb��̂�=��`R����z���M2-&��o����l��kdgvb �n'�^�R:��PpCa#>~��m\� ��Yn�6{��Rܬi���N���#�r5����:��Z�TN�nR8s�ً�E�H2$Z��&�m�M��~J&��J��?�|���h�W]pB��i�y�����5�-���T�R�p��j9� z�oG�/0QU���`�U*��f@0�-�g� �����R�]_~��FDs
FYVH��������� �=U��{R���x)��dp}d��s_���C�	ǽs!3� -���l���fNO{s��q=@�o쑘�]-�
7��� ����.���A������>�IA����H�s)����m�y���Yw��/ g8niqQ��]J_ x]][M�hd�s.$i����wqDp
��n�wH�lm���@VD�z�úNs�;�8Y����ܸG�č��TE-�x�:�u?z<\o�Д���sO�Z;
�H�b}�%�@�kB�g��<��`�`>U:_DR��b�<b@��q�-ձ�u0C���W���"�,�{�s�զ�u� ��jɱ��yQ׵0'6�{ ���� �55��(ǀ���8�l��\7�i�)�J��@���]+m��ߝ��fK�-�:��Ѷ��6�5�Ѯ����62��{�E�i��{:�t��I�e��Ym��u\%����ߧ~[A��9}�-��� �S>?��Y�9�ǀj���=�����OYd(�Ǹh�k���Ԯy1���c}�I"�	��ƥ܉����l�"�%���S4+��ZoO���Ý5�&��z�4?\������� �zr�by�äQ�����ͱ*���{bZ�,�E	{�*�3]Y�Ɍa8Q�~�8�д<99b���N���(^����jp�p����L�-X{N�p^�*�ҲT+��Oɀ���n�*�}bMI��CY��2�f�8^_�p/_m�Y�{�F�V)W��t8qܹ�>�a@�1�GY�υ�La��x��:-p�zs�L�� �Ci����W;���G��q��������_��#w�ڪ�ظ��Q�}� ��=F�����2
�2��g�ޱ-L͍C�q}m�}}�֭���+utM����g�"����b�%xc�QC���Sq� C�`5�D_��g�Wp� �<օ�s�f�tcui-)���gP|�mnn��y.��g5J�e똰���qU�Xٻ|͘��՗,H��R���K�L��%c�Q�)���'���`�9�'�c��B��<�jly�):M�`��񑰖1>$6��z�ʉq��!lۥ�%L%�I��Q�;M��q�)�{�>H�G��iQW��Ć�uŜ�����?����������:V���\�7�V�w!g���3��́�yM���z 8+�������!�p͘���P���'-X����2cq��(�A�#�g�{X/����e0��2��?��C^e?��.�' <�&��W �t�A_�	 *��QZ�%���=�-f�c�.ǆn^�n0-ў��:���xt�Y_#0$�Hd��j�v�`d�s1F�|���\Sl�麆��iA���U��,,,�Z��Br�X�hV� ]��J�G췰�`c ��:���)�R��@MѠ�}�]�e$#�y��A\�.�����VC �f�?'����!'��������8��E�"���q`O`]��3��`sP��.��ΰ��i���.��4fC����\[�f�f��@ĸCq��(�*A
?���f��� h L����2��u�1F �U�O�i\M�}U�1j ��-W-�Gf4�y�G���v��A�؟��J�ya6�ɷ��vѴM��?�&�s�f1��D����Z
�ͻ^�m<�9.�1ő�wgMa?���b� ��4�����%C���9���2�!�,�9��m>E�3���;�����5���?�.\\X�pg=�{1hO�)�n!��(�S]/�E{�M!��W\r�Fu� �@A�bR����[&��璣�t��n�,�"*+饵�\2K��P��4�ř��&�ȍ��׍�289��:��^I���.�� ���w���gt0`p�{���{�T�d8�)��Nz�.�*�d���XX0�3
{j�?0�`!��x.}�6�~�����"1p^�@�5����PEV��F��'c�9��v2���?<�1B�.,t�<����gn�RjW����?����nX����-�Q4dDw/U������H�e��F�߱*{<���nt�稛��T��@K�U��P�NTg�� �����N�J�[���x�K�y]�h�~_�Vt��fiW��c�t�9l6��J<i%�x�=M3�5<�N-��nV���������op�R?�#�4 3��N����o9X�N0�
c�*����`s��w�݇}�.m��5������w�����
(Vj�� �`k�X�R�qČ�\�3$�,ƨ��
8J�~�z��YS�TM/��j҇�j�pZ��N�;��KB���a�M+�L�P_7{���������k`��'�G�4�{��I����L=J��R�D �qn���la+D5�q �B�,�$�5]��k�����B�X���p��#���ل��,�0�
`)�S�����8Mc8�f�3eX�T��?/`�� �����5��I*������Ο�4) ۨL����FO,:�Y��~A�v;��	y��y�$i��9*�4RI'�������c^ٞP�cx��Ǩ�c�4��2"�3"�����6��ʞ�p����%�e&����2����T
�k#�ɰ�>���vO|�t���0�keT35�b�T0�}�� {-A^|��̟E���w%Z�د��t�����s2$���'�A)S���H�4&b�$�agw��2 �$�}���S�uBv�k`C�	nYuR�V��V3����f��{e�ؓ�T��Y�َ�����l��`+猽���]��?l|�d�N[��>�_/�)�|��]��������9� ��?��9�~����ꚛ�.����
i��R �ǚ�9�,	p����Q��3c��,O�şl� �g4F��}��Q���sd'�3(�op9*�Q�̣�Fo��[����:���}�m?6;���/,�����m���щH_����{l��*T?��T�ߛ�G]#�J��n��ƪK,���r߭2�_l_Z��
���B��`����s�M�"7 T���ʅ�(��B@��Q]ya>����=���kW�i<>R���ns�W�����W��t�b3]VY���f��5T������ `E�(�����(!E�c��Y�`>��^OfOt��v2�EH$Y��p0 �wo� 3�)0��0�s2-<:ҨD@yo�P��q}���	��������}��o����vW�]���"�Up��^J�3я�SFy���>UC�@��с o+�t���p�Lۘ��:rR�I	����šP���ч�_�����@#�+��:>bq?:��c:������u��/&֐h�
X(z��ע�	�=e�ǳEQ�C2��ݏ��Jc�O��eq�s{&+7�(����H�U���B�M}��}��������]�|�]�zY�7̅��}�y�P\Ӑu�����g0f��
֫�W�O�fuu�]��pχ��k�L���S������_�[�m16�:}p�[�P��M=�k�M����4���
Q�.m\�<���I�2�W�i�e	�k� [$�Se�p��m�¥Y@kv�t຾u|k:������=~����W��e�ɳ��~k���h����~�Di4ЯR�	ku�Ǻ
R��Y����j\�a%2 �1ם���Q��H�kػ�bo��c|{����Ȍ�9� �1��ZH��-��YU6��7X&��X�h �=zȂn(J�1k��°*��H���+�;�?p���ƍ뼾Ÿ�c�;<R[�I�e9��1�-���Sܷ�.~�jK��F$�K 9�\�E]�|�]�k*
�;(�w������d�,���2�e_ƾ��w�Ǉ��.VWWR�=���������T[
�-`���M�����N����4��ט��6�~��p3��ǝĢ�ݹ��J{lx$�I�s�vt�'A�Z�7�+�sx�T3��I�B
*&V�w�uo����؏��m&�����z�h�d��	�eb��K2bab��h��|���Y�{�{%(<�w�m�cA���c�e��Ͽ�<�8S�>�!��*�G�mNj�T6��m���9�Z�X�hF���k*�L�y��[������*�@�4�5����켯�
�c��̷��-�\����w�r�5��tK�v?�>�vF���vѾזSܨ�j@���V�aGd����m��ۏo��,��?���i� ��L�ǜ�>�rc��k]��
�֊m����I&�zԙ���4#2gq��k0���	�dӭ��j�Ą3�4Yh���)hѨ:8����3aV���R�:�iJ��t���	��[7o�͗�ܽ{�X�	z��q�j��$�h��)�'� R������	���Gu�t����$9�4���(?{�����������
ؼν|��������N�I�������g�}D�n��6�=�l�w�^8������{��≰��7X�7n� � �0�4&ŀ�蠒}�XZ���[��9��Ќ��E�[���t�b���H���F��x�#2�9^�l�%hL����BT欕��Xu�I@Y�}�v ˛/_�1u}xU�dCf�S�U��?����V�׀e<#�
�K�B�܎)�tcHU�8�}�H��.j����Z�����P�i���?�5�0S% ���"��%Xo��T��z'��p�M���ʕ+�ȊS�OA0�Ӵ���֠hx�`�i�*�&��}��\����o����T�<����ڙF��/Ԋ�K�N�Ә����Y:w�`?��P�%�v��[@�ji)I �K`�_(R�+'��NnBe��l�&e:�Y>~������厪N��7�t6pk8��o[ٞ��/����/�I�� ��xH(��.����NO�7�l,(����K�\�14���eIa6�Lj4`3҂�V��R���1wx�J�%4�h,�4�+R��� 2��U*����g�l��h�2�M��� ��w�cTAٸC�_]�YQ& ��eX�.����D�&vzݴ�c�D��(���y*r �z�s̚
�нvU�*���,�,��1�7�r.]��a�P�L\OW-�+	�[�
�9�N��<���k�n�H�����H��"f�z�k�o	HB~l�o��g����/
+�Y�����`����f� �M����Z���^�@�*�SP9�L.e2:<f�JW��\�ic�|mй���(w;�kU�Y֭9��d���	�،JXZ{
�bă7k��O�~�7\ʟ���WN?�������5�2Y��2��A���f��}6w1ˋv,���� ��n*7q��e��	s��p�]r/Z��6;���b�ڌ2�ٻ������P��̺��;��z�.����h鳉%Q�:YJ�SWv��NaN�+�b1Q[!{���3����O
a�xq���8W����^Y'd���qǍ�
���d�1}re�@+���ڣ�u�*�=�l��^شE���Bph����4�ߧtA�^�F���F�� eei��\�����\�B�ggw���p�/^���(5����t�.h3V� ��/p���vZz��\X���p��Rsp$����"3�P��܋����YL�����~Ea���z喲��s��ã��0U������d�Rú�b\�t��j-��4o��Y��@��OGR�=���?U�cĀx��|b���8>wP�������?-��Cq��W�}�����t�0��X�޹8&��R�Y5i8�К�y���6@�D
V���6�M�R.�o�q�1m������yg�Q��s�� >��x�#�4	j��h��{[�2�V�d��[l	�U~��{ .' �Aa��"��ӧO������e����$Һ�����C~�k����"cG����gE�c�%�� �5����.S��-.�����sa]�.����7;��t��:0���x��`ON�7=�F��bLʹ��a����Ǐ܃�7�|��`o>��6� �
0mn��� ��a��i����TM\�ż���L��ﶝ��=T�6A+�7�ʧ �.k��U)�)t+���~��#�n�zAYf`��F�7ƇӠD�br\ot�
��J�����Kq/�
?�@2�P��iғMr:q� `ŵooo����dE�M�v���R�C���LS��}f�,(x��2�h���V @_��`);��w^����pLɟ��3��ԍ; �7<`�b'�Wu���)㸓��	�_)����D[�ۍ���'���+�wYg�`}Dgs�W�-���0 ݞ?3D��-cC2X��w���[z8���hGA��,d*y���c���i?0/�+c��h�S�\0��N�sg�@	̦�1Ǭ���v ��}�V˒b׈���4Ο7�S��f�h����B��z�o�Ae{��5`|��h��
��i� �`�/?���?�]�_�|�O���s�T��;�.*���h���w��v� ���:�\q ��Y��J�-�/L7��8z�t�1�Ω��ٺq�|�i�I��J����=���~~�.���S�!���!T��+�V%c��X�IӲdy��w~J�u�PGʡ��E'�5���sۄ�3����� �`�S7/� �N�C@�"��Kt
PA^�@6�[(�M{o�C������j (>�>H���Y�&��W�^���v�1�GG��/�t_}���{�r�����<&���HX`9X�����Bv��	��ޑ�+�Q'9��ut���Vb�mľ�x������u�Wb�c��E�4+��{�SPZ ކEj �3�C0}��&YK�._rW�
�ߘ^48)΄&�p�(Ki��E4<;��)�E"Ź��>{8�賽���s@F��g�/U���&��:�K>wSW`���ٍs�r|}v�b������(t:����Z�S�Բl���&�:2	(�7�Gu���Rx��ݹMF<�1�Ms��O������
�����Z[]U�{��[�0^ ��?:����"�S��1�P+ږi(��װ2�����|�ⳓ�Ni�M��|(�s�{�S��3Z���X;-Hdl��
�u����y�UA$j���נ��Z ��Ʈ��r[�U<Pn��SټL��E�
�E��Q�W�p�}w�E�,�Z��>�cc.`��Y���q�������0�` �X��t����?dѴw��S;�Ţ��������Vk4�0�6��� F�Ȥ:�{�c
�K�yCj=��md.�恰�;�8�T�x�c�X�2~Cb�Z��4k�$�x��<r��$E{����
�|{�`�����rRq=���χ���ʐ�K ��\?Y���:ns'�h�A�_`���A�j_W���>��R	\�5�A�>cVT��Ɩ5` 4�!Í6ks4�6�o��oݯ~�+����?�]��}M���(v"����ȼ�zR�q�ٹ(��
�a�k+ ����{X[��Z}��u��~H \���8��s�K�n��0@�R#�-�Xi�I�f������_�y�5�3�t�	��`���%��뺑���j�[��F6P��s��*��ǉ�I=q�w�)Ar���.���h�;��>��S�̶������p=�`�c�O�B|��.�-������' ,۠x;S�҇�fj��,�Q;I{�b�2��J�;�˳Oe��MGM~j!��|��%���j}4ɾ���r��*����';G�[9}ҍ�f��r������E�a7q����k�g�ĆЊԅ��/�YKUwE|gZtl�+��׀�sPR
��5���(�~7.�a$v��CM���A�^�'I��4���R�e0��8���ֶ�ru�������n{��Y!78* 1]-,�����K��%.u�0��/�!%!��?w�R�@��_�^�x��Ф�L/U��^Vl�^~�OP�+8����!3 ��p�N�lY�o�c��� �G����yY�(K3�U���X���Φ��߻W���۷o��}|�z�L�"�O��Nt�_<Amaa�w�8�G�9^�a��rrr$���y��j�s82G�R�厲e�B �:붿PlA�2�p���#�}�#-�v$�ݨ�e�S��82>�,tR�i0l����z28���6���e�b��?�y����&��ӏ�G4aڋD��={���%{U\�-����T�����	�G���y�y��s�6�֛���+��/�Y�*�_�K.�g3j��^i5�:���	��*�� 4�BX�������&F\��0f��`E�qJ��-�l�{����. B��Z�O2�9"ў���[�r9��s���9�����c����y^+ S�?zՍ����{���իW\��?�6i�8���b �Iu4�1�d9��.�g��l�ſ8�����e 渮3X���Sa��"D��xw��naVz_�}k�ؕ���{ۮ�:0Au��Sު�1�i88��8kmc}��x�X�8�u��[˞z!�R@�
28V �xN�����$W��!� \U��2�lL`�a�r�����{����>仜wZG���ƵKf��.�a? ��� ��_X�s�k+����g��a����F����+�HD@�a8����V���?��\�UM�C!8+ ���� оw�
�4�g�?^�/�e�,%b�z��5�>v� ��Y��s���Qi�M�]- �5�Zh�������y��:�V���I��j[V[��lX�Ě�&}�}�L�ڝ
�al�O) 朮Yb�& ��̽���('i���j�������Z���M
������l��w��h?�f����%cN?դO�w�'�LI��I'���� Pq�.]j�T"�U��E�碯;�}0�Z/��������~���t��M�Z�^"�z���
#�i�cS�}S75�\��r�K�yR{��X�2F���	?k��l�O�'���\#�0�Ke��
.�ڋ�Cn&� ��,<o<1�tj͒;U�?�� �:�c�,��eو���R��Z�&�tA����s	��� t���k>S��]G�T��t.WV��6���s[[�ܥ+���O>v�}��/�9�o C� lW0���3F��$�ƪ�Zp����|����;wx�+�Ykv���x�C��j�d>���	�
)$���_�u�z��C?tM�W!��	�*πA8>]M9���.}+��h���D����2rO�=�}�	.�����.�;"�	�K`w=��=}��=�,���n�����k	� ��Z��Z^XI,r�H�Fc��x��96��>�=�8�� ���z��l��p@̀U �H߉D.F��C�3��X��F�Z��1�����iP�RM��;z��𼭅|�ߘ�b��\@m�b�Z�J�����ƫ��� Ǹ���`�E��h�
ۮ"`� ƽ{_��k��}gA�ҩ����sI�R��"�U� f�
�0U�����K�X���3 ̥U͵̧߃�����M�ZP�x�Ѽ���8� �;G��,�5����(������<�:-T O(���S7�-��h��!�p�,E8]V����14��l�*KC-�� ���ފ{�w���s;��L�����drj�UFP{Y�ƶc6+׋�	�}m�)�D!�<|��{!����9s{g[ /g�n�MO��|�{��g��:-'��z�����̚��Lo�9���5�b{\W��!HM>g�-3����� �dВ��^� h���v�.ԁ�U�_���t��,��4�-�@d�����x����ݙ�\�k�xF�d�(�=Ո`݀^���hԧ�px `0
�������:�d�V��c����W1<�@��a�l6\��U�a�R?��d�C&��޺���gq+˒^�D������\<��X�O��"�KP�����2����R�>��+:���9�9�g�?�<>�3�mw���`w�|�J�G�1�{)��v3���um�%���2���9F�v�9���m��$�e)(���i+{�PV�H�f���o��g_���ƃ�W�N�K�r��<{���i��L�Γ��r͸�~/��d���u���cS�ܱ@�T�wڱʹ7�]7�]=�o��1`��{�h��2�zs$���1��+�{�^��ȁ�?N�j׎����yA! ��h��+l�l��`���۟�I\TۜB�1῕��\zŢ�Uە*��g��E�3;J����]����m��E+�w���̆/�U3~�͐�5hi,+K�ڙ,Lmr\�ld&vFT�c ���ΕA&��X��	�lQ]=l��'���ya���h�P
��uq��#4"��) �eH�~��^g�D�οc�'���5��������/>��p`���[���CW����P�P
�aj�T�g!Aeh��X`Z�@t-����:�Ǭ��y��Z��q<^W
��vI7֌<8�����2�` �|����)_����RJG/vǣG����M���
|��G���������|钻�O8�� ��Gi/���0�%éƚ���ԅh'.��}li�W�\�x���y�� >Kы�8�
 ����%M��u����ú@���"�� vc,	X����I�.���L?���`e�k���7��.����56b񞱢D��s� ��|M��g
3�8F�}q�E��C�,���DqK�����S&"��8���y&�k#�:�SUM�Ɏ�`֑ M�?<�"�픊9��rQ��o����Z�ْ{غh�͎ž���/됱Cwn.�^�dp����kkH�'�P������l"/�Y�V� ��p�H�i1��gi�h�U��0 �׫�j، �������` ��q7D&��c-X�X�Y���f6G�]^Ui���"���+���V+�cݶ�q�����s�M^��|��c�x��UZX<�}
0u?�����Q+hW�=����C��c�Gߠ�p��?�{|�ǔ�j�N1��u���������X�}���&�ĵ"g!��G4��:�)�u.A����ܳmv[��jp�2����%Sc}Q�s��oa]鲀��+�z����H��.��)�i���-أ���މ�y��Q�K�ҖjD\'�/8��az⸷��MܼyS���k�����y�;΁s�^!=�|�����>����Ri�\��J{Ώ�:X��w{"g�~0�5s�, �����}��$x���s��cߨm��W��d��u�Zh��[	�n5�9&S��aL�� ��:�0B�<e�eP��L(��o{M^;�EY �	��>�3y+��lD�!1�:�>�CX2F��/����fc:�)��kˀN���ߩ��qK��%0e�7�]�����St��4��E;_� �g�1o�|�K��z7�|�Ei�vXju&�}I���
.�ל��#H�ﯾx�e^��[e���ʸ�[^k���K+n�D�}��v���[\�Q6��UR��V�p��{Zb��񢀨���+N�� ǘ�Y�5,]�^�5�6���|3�J��-�h_�����(����Z�P :� �4\�|%:2O��ˎ��9r�Gp�����k�x�-.=r�3p'(J��q+�Qd��xQ`,oEGip�V2�&�5 �CF;�`'!�{��:C��}����b{ʶ������R��]�Ժ6�;P c�g9O�a����g4�D���WFU��a�2iE�L�n���?��i)M�!01O�}�l�}���{������,����ή{�4&��Ͻ��L6"tf_��tO�>�y �ߺu����pY5�(�~|���<��X�egM�hӸ�B?��}��ҥ���ᤓȱQ�Mj�֧�z}7-���"��_�0'k�,��ʪp�3�S��!ӥhl��@����F�ם���{J+���7��S��Χ>kt ��YaYG8�c�r�������;�Y�/A�g74 ��L!�q��e�^��s�ޔ�f����Me������s�����,X}�4nT����Tk��_�ti�� ��,�65�rSև�E�{U�y�7���8��G�t��6�V+~�S���&��,�����IY�+K���YP���g�x��lڨ�:���ڲ�����İ+zd�UI�W�)4k��3yY�xn�=v�|��9��&�{0f%��U£nZ j(�kkZڛ]�D%��]+�����I� ���z�ش���ɡ�AO����6���)�f�5�Z�_�T�.(	�ibא�u�B�_'dĊַ��=�75~�=�Eا�' :=~�©�/_�z����X�����+�{]�R-b4�pQ.P�G$��	3�q�8F ���mu�*��B�1d��F{���� ����4�F�/�R�O����ᜲo;7`ێ����O9(�TP�0�b�Q���ư`[�A�k������C�u�bS!����`O��[��ε+�����\Z�B�!'���3  fAaӮV���H��z��JUivZ��b`7��f@�f� ��a�5'M���e�`l@����T��Yt0�i7,���Z�~!}ᝩ"�~����L`����؛ �<>�p��]��.}>�#�ה�3T.֨��_�˶��8j�df������l�h|���S�*G�����`�>�͑����%��_�f��~:~x_^�s�!t������z`��@v�S	��Ѯ�CV�2��w1߾����ҙ8��:n�)�	����8PG�ӂS�X\`aaL�^\�W.���'t�������1��63pZ�ߩ���і�0�qr��<�N�E�h?���^[Q]ZY�|UY9��:8 �XRGIӒ�c
^�X5���鋽��E��u�:m��4J}t����Q-��$��������PX���h���1S!�]�s����q���ဒ`� E�ً��f�=~
y����YpK�ҹ�/D��AsL�@���27y8� ��.(�9�Z�(HL���'��~��2h��}�={������,ܷ���VW��vV4उ# ��F~����)�P�ڵ[��������3a#��q�ymm��������%�kH'N;�D�i���A��F`.>�~|>�}w�Қ�}�����9�Rzoo�@���Zt�%U��G��3���ظ�q�m|�믿&�pZ�W�^糢c��q0��Y@G���t
�	�؀!�؟�h�]�vM�, �^��	�'�9?~Lg���:BA�#�y�������L:�<t������~�ap�Ps���9A�	�J�Z-?N?��ϏO��D7i�i��?��v2�b'���z��a�P�EǒYP)0��}P�Qmds�3ج�9:�w �2~�A�,�c�}��7����{rz�6��^����gv�5�'�~OP���A�z�ǜ��qZ i�"aݸ�������Z�9�J�X�qN���)���Aِm�X���.�y�g������9��*���-!ɱo��.�0��w�F���ܕ˗%{a}�`��>r�Und���+��7� !�,�:�ǵ&L��V�>�cC����#����Q`�a`O��-h��1�F��'r&_�f42���O�#�O ��[�����x�c��K�K�oc�;���i.�쐩}���WP��iӟ7��o���T\EL޵� ��u��"x�>B�ha�˗6܍�9~�Ž��q�݉������L��g}�`&
�~�����=,Y�ko��y��,d���͒�X��fa΂-����%�$8����d���h�8� D�S&n����(�P4H�֜�j��~�+����`�}�a������:�ѥK��J��������<���|������v��8�M�^��P3���ё`<��������s;[�����P�#Xh�_n�T ]�-4p��,�$�E��#�}#����E�S &Ce80�;���<�؉2G�v� ���[��OȊrNU[��k��JߌF�XG�	�)��f�5�F��Ɍ�Bѕ��-�歎�i/�rm���b��iM)�b�6@��ek�w�5�+�<��C��K���Ǩ1�t/��;m�8m:��8���|�s��=N;��`�<~�mɖ��
]�Jj�y�������y:��^̓��}�泽������oG�+	,Sʏ�r��瑡җ=���&�w��~��',�q��#`��yg�R6���e�唈I19����0e��6v	&�����kߡ��-��ܔ�~���_�tS��^�?�fU�ь�k�.��m��&���!)��z�M���7MN��J�!$��4�kK��$��du�;HU�?MKE����K�*m�TK8]�ˋt`�h��Tuj�=�� �zt=|��BB����p����}�V��=�j�f�K�F�S�jk��Da��5����L
 �IA��嫗�|@�����{��Kt�E
DAc�ځ9��X���B=�uw��ew����,���p���3W�9Q<p��C�u�H>�k{��:�3XHI�r$�����ncc�rp�>�������Yp0�!��~��}a �$����3ٍN���O����v��M๙������Աi��^/�}X��2���Z�`��E�?���g�}�����%��,5�g@@���98��@�{]���V���\y��Tl�Lڒm�9w�����q�Z�6W]~?�o��<��v�,�`��8���Z���Xzzv.\�J ��)������cw��m�V�'�=�28�v.f5\X�X�%=��kH���N2j�6��u�]�X��D�k�y XO������(A�k�Hfq�����Ҵk�,O���0�Λz�Y�B�� x �����/o���Li�����Rȝ���`�q>������R8�~
��_�0NYm^�k� ��
�b>#��@���&�cV<�z6�ǰ_��|
n�c��xH�&��F5|����R�Y�2o�Eb2J�y�u뭶$^����r��jg�Q����Mk�x����e�S����j"�в7,����<��-/��y"�8Ǭ�E)"�7�������F9's�`gU� O�ߑ,.� �2Hݗ��.�k�k��.ރJ����X[Y����T��e�-#e뙟9��	�D��������d(@4��X@�>�ϐ��~�����W�w�`�G������qޞ�,�� Z�C\'��g\7
&�<�}[�5�D��������y%���ފ�J݄n*�ɀC�9 ��SV+�&�ol蜮����#�I��
��2Ã�+���_���,�g{tm��!BjF]�V�/�#�y���v��iw*K�/�5�0m�t�$�:�t4��@,o�v�{B��\�`ʼ+^7	��ϨU�c�����%iR�?�����f��寿9"i��[_�#�����������`��F6?$f�}���@�ı���__��8h���ƏW��n�{.w��9j�)�%���/5dL��\��]���O؜W�h�o���6���Dӯ�Q�Z�T�qS�qY����H��`���^��k����r��R^өm�&Ob���T��=�IR����ج�9Z�V]i�:1xe@���^��]�N�c���L�83�=����Pdl�����]H�$8,'�[���GH���V0����Q��iE�d%:`���ݪ��6$)�[ۈNOt6��=>��`� :��)xY�M�l�ؤ3���L�ju��<9�&���.���Eg������
�+ ����� �5W�)��� ;������㟹?��]�F����|���b40H �����sh�B.$$�[u��yt��q*v�{YX�GG~1:�+d���5��r�E����(�s���U���ξ�3J�,Eܷ�몶����'c�9�ݍ�W*p������y��)F��R�������?H{����(+����em ���щWt�K�p����i�r�y�(`�������s��[I�������A6��l�"h:1��mD�5^=ok��`��qP��)R�z��k��ڷ.�����Ɍ��
����}�ӺjV�a�!����� I�p��X��T�䲨$��8V766,��4pe�2�k�F���9{�R��zJ��tT}�?EnR:d�Y'_Ñ �Q���^��ml��7n�)����� �e�#�����I���B�2���$ӻ�-l�q)�`ΤO�`���IX�X�KٓO�>s_~�U|^[)��Ղ\&�`LKK�"gc���_ɤ�uk$�}���ֽ�Q҇�S9��?����u���g���C����Ε���9���~��a^�4$&���o�o�=��-���ܥ����g��{H3��ˢ��g{w�s��H@4��X/�f����~�p0J�1�1cܳ�q�@.��+AT��Z�Y�Ч}p�5SG�+�i�;�:�{�g�����q� �pȹ� �V$�i��|��^��޻s�}��'��_�G����3J�w=y�ͯ�).T1Tn�� ����y�@?�eʡi ]�;���&��=2�M�lN��\B���!X �n�`��X[L�������`(�ؘӲU��we��邿��>�@΄��<�,(�1�	�6V|���Ƙ*k	ey�x�瓾_e�\^�|��6�گ��4��.��1d9�c@����ڂ��-�9�b�Ώ�!u�c���&�n��K��;���6��9�� Qϩ����t,��Sƚ��b.���3X�V�l����<^q��}*�7U�ݧ�L�����M�͛�e�b~Z�/S�K��D¨�M�MY���WM�~+�w�f\�E{�v,��FY�oyU�0Pg� �ĹW�6�F}�w�{�g�"��	�zESg�'���i~�~��Q��*UW�����c �n��/�|��u��8ׅ&�[o�
8t��BLS�.,��,�e�Z+8Sk�2֦C����@�nW�B� �l�'�{|�4W._q�66�����`�(:�+niyͭ�/���m���ž �G�����x��._rW�]M�Ao'�pB��^��	����|�˿�6������W���;tj�,��	�K�rtP�:&t��8����� ~��������]���⎢S���M���{w��:���w�s�|�-A�o���Z��bϽ��5����{�|��t�����º�v������w�w�8`d��������4��q����W���o �ׯ�`��Z,�N�J=�ɴ�{���znM�;�� `!jH؆�ʴ^uj�Y�����{��{��'dV������6�	N=��8����Hqzũ6GM�5 `j��jӠ�@-�E�?�mA�z.�瓃�ݕ�r�+�9�s�ʗ�����d(��=-�
DحL��y�fʲ��c8,�u��HN�� P����[�c���;Nb5��=�(_?�^��Ŕ��x��0��&|�����M ��¸ -���	�����'��(�g�4魿Re�C��R�u�&�6�7��:{ccnV�����p�e=W9��o޼N`#0c:�%s�lD0��s�}@`��=�VK����K{����'}�����	��#f��iԐ���Z�áh�z-���]���u���S]��T;��2�� �*��פ-:���s6��;s������g��ض��~+���*`�@��ԃ�}�&�Ǿ9�}t�4z����:>��g�E�����n7�dx��u5��P�:��@��n$���	
�ʵH�U�) �x^أ�Xh׊�y�Eb��&���`������t!x}"�d�`��N��x�W⼸y�Vܫ��_�VZ�q?�ٳ���_������ꗿr���;i^l�T��;Z�#�1[��eP(��c��/���>�srS���U7������B:>�z�6�)<f��=��Sq��{7ؓ�0{H��9Y�"���dæ�L	2��7c�@@SA��[�r��S�cu}ŭo�I�j��$p̠C�-�ds�2��o�f�kw�iA��ӓ�O�H�i���$���O�f\U���2�����)�p	؞��S:�he��yg���{K`�m�i=�;gw�6;S�3�0y,ؿ�M��1,H3��r�Ď[*V�|b�J�>}]��&mV�_�ĥ�,#�|��Ӯe�m�ֿ����	�N߫�/�QPyN�L`/I�	��b��E�'��v,��f�}0�l9)CeA�J�8&����Z�3���7>Os�^�)��]�"�M�P������6M��*eI��{v��^��QL;��Ęb�nY+������M����|���,�k��T�ƹ�8�V���� P�&A��eZ*X���tG���X��1�Vb�t���/�`&$Y�0�� Q_nn�}����CG�S)����Ft*���b2 ��7R3Sz��P��\��Y�G���G��>p���_�۷o�ׅ݉>A:�!��-�88��j
������Q��zE��������n):W�g�� �qn�{���ɧ���W��i360Z�����߿��er�nܸ���/�#u/q��_��AO����w���k�c)`�����Z5���Y>H��Bt4��)<��s���v����T�O�ϑ{��)��++�o:���^W��w|���+�W���[_�䶷�2c�k
���d�'R����t~��������TX��Yb_8sg��)楨�)�=�%ǧ�����-v6c$�l�+�}�bV���{e��;Џ>�0^��3����q�^I��ᚍ�
�,�ޡ� ���h�����iX'�=+0�q?�&��d�uEǀKa%f�$�R���KG���LJ��M~�xu⎍�'�Ώ1��_��-�1�������)�$b��� M#�:Z����2�� ���K��tk�ץ�	ؿ�I(K�� ���.S.��*�e	�t�1H��Y�p�=k8�\��+����̋����*�9�>�A0N�F4�e����7uj�S���5����zY�q�wZ��(e W��dO���"��@��#�[�s��
N�Y����>�"u�3�0 �
��|����KF��fw��xqO�ZQ�@J���/�}���Z\Z�X]�[����>��]��~�����oi���-���P�+� )dBu��q����T�9���}e�vT�a���d9�w����= 6����^[}���_�����GnwwO�6B������Բ /5��q�F����_n�OQd�RT��/���#�96��.�g�$����w(��l�yJmX�@���7n���o݃8o<xȵ���;�ȥ8	4����� E�1�Xu�&5m�4&I�	���� �"�̘hj�}'۽e��
��� F��3�ɴT9=*�X�2;�ډ�Lɢ/�a�]��H+h�rT�y�����ɗm�Qy��}�1�u�Nk�q�)��q�V.M���7noۚ�޲��?P~$�賐�c�Kp��z�����������/�^��I�L����9y�Ӥ,J��2��]��Ӟ_��m`9�ӹg�&��86�/:�$}���� �s��w`]�S���F���䗽��UuCh�\�j�*��e1B�h!������-��Ŕ~�h�E�hv��e�:�M���(A�,E�B�nc�8/�D>':{N���EK|=��SO>ް�P9�3�$��T��D �<�&n�M 2�#�)��Y��7V�I*�˕�
bT�.S���X��nD�0�ѱ;�kL�.�+xM�qY���k�m�Z��=˶3��Q`��qtf�v�܋Ϲ���g��#5�+�m�4*LZc8� ��?����W�$c�� >T'�78� ��p��@o}G�y=z�
�,-��c���y�4��^�t�}����.������t�,���G���f�ghI���{�o~���d3�|IV�X��[�����]#��@�� /�۝��Fj���&�1�-�I�z�cA�V�tbѧ8'@���]�wd�kСIl��%jl���?'���k��|�O��/��fls��s&3�U�ȥR�
�p�<vS�牽�O���6�YS�@��z�s��f�����>d���a'iz�}+��8�0?.@�x���N4@�޾�;	iА�a�ik+��!1׸�"����h>�1ps
��h)�)���hTP0=����=�Y���7�{g==��l,�=�W�&G�O����d0b-��u�؟X�;�>��������*��*2 ��l�V�P2�{�֢�/�:0�����뛭w�%SJ���j�6-���^��p*�P�@�,����JP���R�DO����Q��I�5(��f��N�-��9��d k�:�S�\:���{��#��c������xσ�1�=e�6ˍf���98b/�d'a_ �*@T�C2�/]"�k�����H��d+SB�S��)]-�����k��������� Q��'��q�5�`�뉮m��а�"�����}��%�3�Ml�2�:�z�C��ƢX\%E�0ov���B/�;΍�i8���O?�T5�|n�ek�e�=ύ�) � �����|�M���GC�ů�G��E=�\�P�O�E[��穃= ��{�u�Y.Pg�-���"�(�� @���"��ie6�w��5X�a� �I�)/�5(��E�5l����B��R�*�Iۄ+���������W�]��������.��(��@;�C�0�ޥ9���M�k�$g�w���Lio���}�p
8}�cϐ�|�#���igxkX�_� h�{�����1k���.*:�\C��p�7�[���?�>������a>��7d?��|��&�Th�GG�Mk�kI�D'���[�sr,��)t�f�`��[9,�E�bt��E�*�4�U��� z9�,F6���o�>��{�9�l�v���Z�~}Gw�Z3�������fU���i��/��w��+Fu�5����0ip����k�E)�D��@�8`�u��XAd�@A�޸~#�C^����0
`Z�)nc}í��Б{��~��+��[����$�`�6%#��	@�S搀K}���]��^�{�����ft���>��������׮E�j����� � ��� �)C�0��������_���y�;�ۋ���߃c5bQ#8���FK�&�e��ig�0�K�n޸��X\\���sw�����`���W�Y4����7�ϣ�9��+�:�L���O�>��F� �k}�;��v�A�3��[�� ��93]I4)�^��W/7���d;C�L�յ5�x�q�	Đ��!@�^o.��!���j��)�ih܂e���|�����>������݃���ޏ����6R�o8߸���}�e�E��BS���PQg/�������s��s�a?���	'1H�X6��i�y�Ϭː�v���q,�l��A�f����Q-�J_Г�E��ɶ�����y�YeKq���O�x==�\�ci�O�<a��'�A}��u*�0n��k)6�'��@ (��b�e�J�@����^7C�_��B�f˵of�ƺb�c;�OOq8��pf\W�]�ʾ�PeT;��UG�_��ਟ�`R*P��a��X; N�Y�O�.����]��F��^<�k�?t�q� ��Q�;d�r�k���h��ݜ*����\Θ3j�E��;w�q��畂~M���ρ�\&_$֢M�P<���a�ٟ�Ʈ7�\A�b�%�e��͞1��;q�:8�q����`��! ��Բ>T�	{����c���W/�3�O�/�NW��hP"g;P��{�I>:��n͜0�����)��m �	vwMx���	�lk����>��C�ဵ� 	�,/_n%�9΍ 42�@��x��Q[�z�]�E�A1L���R����ㅙOq��E����6�p/�
A |)��W�>����6�=��5/�_� '�g�����{kg_4�1FWV�'8@��`<�p$6TEPy��{�R9(�e�N
�i����p�A<O�������:�Ň~�Vc�"���W_�����#��g�`��믿�m��6ļ~������@��$'���D���2�*:�@0PH�|�.$m�T@��*�e>��m�W�Q(�ƧⲾ(������g��ޝ"99���0�md
�u���Xq�\��^M�FŻ !�x�<{��]���D��^���7_H���;�ؐ�3]����%�8�����ؾo��r��~��Ź�ݻ��Y@�F�C.�j��i�#�W*��M�2�/�X;���bß�H/�;h���Y�rnL�Ceae��;V@�J�{-z��D�-_�Nօ�tk,*Vn��ۥ�tʥ��.[���a�m���.�E�)��R���U	z5�4W�w�V�F�ъkr�Is�-�Z�]!�d#�Qp�)ҪI#8������*c`�h&�x�� -i��N�b-�΂�~�Ft,^���6�sr��J����=�s��;	��l(���َ2q}0�����s��?�3+�NŔM��(sٖ"a�xw���=�|������(�Q�{�V20���4Nz]�:*[+:��F4:�VW� �p����W���={F���ޮj����ݻ����u�>a�ùE_nmﰐ!�}p��ӑ���� l��W�ʾ�۷n�Z�8�'��L.<?�&ԭ%x,�-cJ�����B*�����6�]������ݗ
�'����x[���7.o0-�Ν[�Qqna��16��0)Dhp��8a"�A+�Dw��ؙ�y���M��$Լӹ�4�&]B����M�<3 v��S��3(�����'U�f?�AS�2��I790��4�Y���q\C[����ߏ���iM�j���7]S��Z�*&���n��;q����'+�K�>3Ze���T�@&��e�Λ>a�����苐��`�w�#�4k&$݌�Ǿc@~��FG��c޷�G81�$�p�uW�^�Ϻ����X��R��V 4��>�6s��D6$40������y�&h�N/e��)}t�5��Y�
hp@�n|ڟ$0�т��� 	�RZ�g�bږ�Q�W��"h�M9�.�z��/�~�֜�SH�����o�fn����7��	d7�X��:�>Pn脠.�C﫣�n�8v�+�`�0���t�G����8�/_��
�2�X��G��,��#����	� �*XX{h�[�lݲ1[���k�k+J�u! [��`3 xŚ��+Z��L�Z�����N��a/����XZ�>ďI��|�w�c� +1j܃����ލ ,�5�*��U����~Y�=���?��q� P��f'�����	,3�E;R,���I �$0p�x��e�i7TԺ_eP{�`i����g���}���E�]��l����7Z �.XĒ-!Ϯ�,&��5��'�Jd�[FM�YNy��C��?�)���3z3~깿��p�p�3��V/��[_�Y����_�8��0~�u��/�t����w'/��n#D� ��ʢ��{3��������M*�[o�9�[�.ڗ6�Jq�Ƀ��V��Y;a�o	�Z�>��d*w�T�ڐ��}�`��یF�4p�}��Q�,҅w�jȈ��v��s��E��'��p*�`)����3&�7FA֑j߹H��E���4)����#Y}�@jp% �8+ l��C�����I��u��ZSM�iD3�,�l9$��5e�p�O/��e� 0t�ธT��J
� ) T�[Qo@�0�������t�������wߏ�T�/���r
�Z�E;/�`!Ւ쥡 �7��&`���ё��`Ā���N �p�y8��8�̈W&pG��R��	��_���ۿ�3E��H�Yq?a[�D�L�,�t�k9:�	&�A������=�~��V���?[[�\�?��#j������z�j�`�56�Kh��D��y��<�/�����yeѼxmW�]#�L�gϞ�=�A��%68�
z�ܙ�h�uwY�o.1��$�3�j�p�����×�>{�>}��Ę��w�Riye�}��'�4hOg�/��g�_r��-�i����O�B� �U�w
@7���b�L���435L8�%�[Lj7=�TЛ�~��)��>v��4� �f��Â�1�k]M.��&I��#ս���|�K+��k��Zq}��V�;yf��A�cj�k1� �2Y��-_u-��VV�Șɗ���8�w	��s�/tH�6>��?+L�i�Vl�6c�<2�]�`)�Z���Z&Q�|dA��HGHqU��(�Q`�Zd���2e66�Y�k X��.Pbe��"�����h���{y`2B��޽/	b�5�C&w ��u�e���w�' ��c�N�� �`N�\��: z4���zo�dL�ݔU%$�R;mݛ|� �ޞ�N���m���gFI+�N��߂!d|]Ɯd�`y��D�\�M�_n�gϟ�CZB�Rׯa\^f`{*��`��X4{D ��d�ޔ�n� 	��TC�V�n����1��\ �b�y��|� %~G��஬����saGQ?A� ۅ��om�P�����j�#�R\�����}ptğo���{(2��G��v,�
A�ޔ'����&����,!�(�Kˋ��U�J��U%r6 ���n�2��Ʋy���S���CP ��3�{����9Fnݼ�>��� *#k
c�����y� .k8t;*eh�YIpL�f���=H��A��k)��"%S��<)�f�!a��J�>��x�H'�̥�yc@Xk����5v]2>���[vA�3��ְ���w����7�Y����@���o����k�m<�{l������TV��/M�ʳ�l�4�bq3�6�����{��:ݜ�+��g������N�fs[��0Ha ��g�)�2�-����a6��Ll/��&�|;ؙ.�T��w��9̾ �/�O��a�Y�MC )[���g�=�,ɒ+1�x"�֥EWU�j13= `��.��w��5���`��v0�C=�EUwu�J�u����7^����ݳyg�3+3^�W�?~�`IM�, ��n����+h���V�;��H;������J���thӔC�DM7]e�dL��r�MX�.$����d��n�}�1��^|�9�ʚ���d}#22:�j��h��-��_��722��=>ʨ����f��@`�6�ego_޽��2�GF�<�Ho�L����Y\\��mT,?�c1R�\ع��l*+
�/���i2�����?�����s�f�X�<�s�� є��Z��WM�v=�����}����=��H�3'r��e��4��{��LNM��\����4oeyE~��ߑ�~8p3�f��N1 �ŅՁD���ɉq����Q�d3��}ڈ�`��`q�V��p�w���Պ>���Q�E~ �@��	g����g����>�*���'K+�25=%�����_�O� �& ��t���%y��Y�fn�)�h0B���煶i��
���v���^�jR/�����#��7�-�A�W���8q�=������6D�Ka/*6�����I��`����I��V8�U���0E��ҍ7�7�-�w E��gwvV:��s��شc���Y_o�T��TdV�T�[�Ĭ0� �� 8d��� ���Q��I�1+��� .��)�܉ws�E�4�m
�`� �/tH��>4ȵ k5l�v�0�W�X��-��v^�9�,d+�V]k΅���$���mb g̮z�MW �����@$�����x��̌5�	��8�4����g�e��g���e������|��	�6�MOM��Ԡ�8î�!���?�d��F��eQAATق�y���F�5�
�S��>8,�|@�Ăc�< ��8������b���W`m�D��ߞ�;>x�/쳨C ����k��&����u�o���\R��3X�#�y��@ �1�փ��`Xw{�!��
V�NLL0�L$w���`-����x��=SU�vܾ���E�R�����ܲ"|����8vu|kq�Uq�ϸ�L�8;c[VV�t��zY�D�"�����ѱ�)e2Ł�g�׾�~���j���VV���V�.��� �;���d����|��5�t�2���O�<��nޔ7�|��C�6� �qO�󲴴 ;;[Z�g��nH��YK����+ �:�����m�����e��_n����YKE����d�����>8�램�ʘ�:�q�m�\���	��JK�!��b�J2;��W�a�����}t�u�iY��P��ug�F����?��՟�4#9��w��tLg��i��g���Ɓ��(2r&��HNL&��C�2�;͈���}�X�ڭs �'�Nc�V�6�FHQ�%&T����֗���%"����
&y3�ԧ�t�ʋ�)�����.r���o��F+;�X?���K`Rtpp
�l_tK9����Ag�`�cL�L��b�a��gЙ���AsM�L��ML&����x��j��I�"�`z��AM��#8&�[�<74�z�UU�S�;�zo�:u�� P�yK��#1<2蜺Y]]"esc�9#��+r��5e m�����,�EV$��qHZ��:�J���XU�z�xoΧq�H?��Wdyy+�����W�E��<h�E!���yG��|͞�b�jp(`��� ��5�f��4��ҽPv���MS uOO���i�Ѕu8�`��Zz��Δ��W��#�d]����)��;���:'s�)��;;d&����N�54�s�����64<��sc*cŞA8�n\�=
�� <��p�~����XG���ȭ[�Ȩ�}z-7�XΡ���4��Y�x�V����M�0�y�4���СK��h6�7sʌ]X@]�����:�܅����%��6�ćvy��ʼ���y�U--x,;
���=&P�Z5��O�w�LZ!������p^�����ey��\�zQFF�Vt{���u��큲�X�D4X4<"{��d4��~^�IT"���Kc�dv�C�N2 0c��E"5e\t�N$�:ZNJ?�ĂJ����ω��)��&!�,C �Џ���~J���Ǽx�w����Vj�oh���c��d?y�/��;�6c����={�V/$k��2���ϟ��h�2X4c�{\;���{ˣ9�$E�4H:��L��}��=c�g���������A�H���s)��-�,Y�'�~���nw�l�b�)[��K�|���E?�0҉5(��p�\���#4����;�h([D��4�j�wv�	�A)ISc�'�8Y[_�L��z�˃oZKF��Գ�,�A�F#�L#!��-$7���d���	:�-ˎB1ي[3�=��D%d�����ϭʘ�?j�c���U�}��Z�r�}���q�Z��{�%�Ou,)����g�[cpo j�?a�����X���A�xoȹ���	` 9�
d1�� {�;�n�*� �jH��>F0 <��*��Z-��Oz��>�~~�����?�����k�i!Dw��fp,e���d0�([Ф.�M	^�_��ِ����{���a��E��&�]��}��w�ǵo�� D�YV9���?�O�h �tcZ��>%�$���	Y��$����>�i6N ��b�|E�X��$'~�2}�$��������y��ww�h����_r�'���HgfK*>�}&�?O�����|Iǡ�sw�]�1��y�&��j*�pOb&)ֈ4�'��v&@��}�v,'M'��!�lƖ��)fX�&Y`F��_ofzs:ZJ�����Vͽ̬x������\N��������ú��Gݺ�����:yl�����N�D)R�᧙~O���{8>nǖ�T��&��v�$#�7O���)���K"K�Yi�R��ʩ!%RAb��]+bc :�U�����a�G����φ��N��5��-��B��ڶ7Ed�¨�}�.i=�,��AK�O=>g��~��Ss��O�OLL������099%33�d0=�X��O)Ͱ���' [M�� <[�1��Ɲ7ސ��i9p�&n:Z1Y�6{P��5�׳I|!F�#4L�7� ����o)�Y`2-l�9k����8A(t���?����g���M����gLӆ�E�4�Q�� t�h����Њ���(�-Mf�kfv�ρs�u�k���{���'�Y5�x�~n� � ��7-��rl\�p��1�/����ׯS@� �nl�0�#�Z��۪o��cP)O� ���6�a�n S�Q[V�{i@vs9!qq�u�M
�������~�����l�J��%2!����]C����xX5�=P�jy ��-����_x�`�ݻwO����8��w���E�&��=����xx��A/��?DA�>
��6kf:��� �V��Y��~���� ؂1�?�'��Q�k ~ �Rv�8܇���͑�fO��CN^���8�%���hZ74����=��G�%`��3��$�����U `�&qP�,H�@�۱V*@��q�����ڢw�u���n�\]]�'O�Rc�f;�� ��z��`�Tjv�{})�I�"bcO3mj� ��s�����Y�a������C�*�O�|RZ�kD4���-EP)�|���<��)����>-�Ǯ�Zd��zO�LL��  �ח�qt��;:6��\��zh����&N�I�|�2���
�Z�-{&'�T�@�����̠��׵j�w��R��xcn����v���*�ȴ������4DEf�e{kG���d�����,$+ �R�������eNT(��^�U�c�@��q���wd���5�����������50�Ų�:��0�"���ž���_�6 D�q�;�{�')�:���`�}q��M �qv_�k'>�>�d8�ٳ�|�������Y���O��)؀�V3΃~��i�% {!с{@0��5��lk���ζ��)�9�C��\I�!1�����w�JOК�̾�x'���o�2��Ij&k����>�}�nLc<����3�h-�l�����9,(�������&AP�@�M�\�fw5L�揁�`1��?���ZBd+�_'�'���������c��:�9�K�\ן_�Da벋����}Km}�Q���9π������<���q<[�na����s`�D;�0{�"ޭe�@��0��2=����5�Q):�� $&�8�<�|�$D���Ȣ�L�g��w�u�!���*敿������/��X:��X������b��:QҮ b�1���o��es8o/o�����M����H�}28�h���փq���s�+��Q��O��8����'�4��Q�eZ�G�����e!��ռ�,�S�Y��vH3U����b�� 0 [�v����d���H�\t����M���i�Sg�|���	JNl���1�6�cc25�����&�	�S>���2I�@��"��a�X�ea��������Ν[r��uw� "w�F9;���H�l�����<{�@�A,����r�(`���_�w�yO����^�{�dkcW��:O�jc '�
Z��#�f����Ώ�'&����׷�������s�p�ީ:�H��C:B*�o?��<�L��&��u�@vuF�d
�,/�i859)W�\�ÿ�zς�G�ouU���V����0� ̾�!Q6������]_�k�+]�U�U���R��_� 8=<<"��3���<����cw`�f b �	,��ƪ�021s*�$��aK��O�5^,F��Me��3	��9�U8��tl�2��-@c�aN{`6�[r/�O�j�T<m�=	��8����Γ8Tα��ڔ���߃k��;���ǰ����N���n����5(�27;��	�̽�^�����L��U����ްGi��+�!��r��%Yr�R9D�vl�Wm#V�e�����=  �5�"Csw��B�)�o! /� ��Y'�F��w�/�Ǳn��pj���@��Z�4�n����Lz�g.@��#��{�Vۘx�a.��Or=�5={��3��<~x��2�Z�5��Ç_p-B�jhp@��Y�c~����3��pc8՛x5�[���Z ޔ��	@"` ���s����]
	-0V	//����-,�#�ᥧ:gC��)��D�Ǣ���:�����8�://K6޼�/_,���l�A"��`�̤V����v-�����J ��YY�4}��3iz)�4$�;����׾jo`��X�@m�볘/$L?�k��"�n1
������S��clV�5#ãn��=�2�Li���y��ŅEJ"�.��e���c�̺�^R5�`܋f�[�D�t����|h����;{��iˀ��@��>�q�����07���s�xM6�t��m��<���?�/W�\��%�{��tLbEf�U�!h � ԰743Hܽ��	���y�2�!�����.]���뿓ZZ���Y��w��`�.����-�ls_�$�����c����dF��
k��(̽�q}��[%���ʨWPY�����@Qqׯ�/�"Z����.��ܿ�@��ĳ�uֱ��S���[���
0�6~�2��E�ĳ�Ӱ��D��f��֯/��	����9��k����IuH�=y+/�ǖ h�����I�pw���F��\��\� Q�545����o�����?��v��s���s`�D;���z�ٝ�[K����tƈh�"��dYd )e޴�5I�W�Q'\bD�bQڄ�����(��:�m="�]u�J'?�����"&�S���Ś�A����=��wi1�6����Zч��~��=@�@Nf��,K�WH-�/د|����@��[��R�y!�K��Cl����7�Sc\4���6�+8����+�'��'��4���K���fl�8s�6�dw{��wv��vKf��lL�ԝ�d�:�K8� %�����7�����2��u_F0�Z�8T*�nۚ���~n~>uϾ2M��kW^�7߼+7_��k5� ��5��8Np�D�� Ss�Y41W'O�5ȌJ�=�C����`Q��4q勵J=e�o�'��~_���E���=�ӟ>bjiۊ��w������̡�)V`�mRc��wg{�@����Z�� ��,neY��>Y\��H���ƀ̴�a~D������v0�����C ,rȁ4�=��c���W?/7��cD�Y�&eEs*��ۦ������kR�����f���X������10�ۚ�u�w]�;�*�����l {����8s��D|q7}vǵo� ���qc0��<��kM��z��_E8�,�c7�ebr��h0s��F�J�ŀ���$��L�~��.�5�� ��n���p2� ���f�3|��l�K�KȐ����>j�
���:v!�^(�a̻��g�i Q���d;�}�ȩ��>-=5��ZM�,<#$/ (#}�^�!��U�uL��=�
���L����?X��e�5�T��A��΋�Ki,�bظ�Xg��a�⋇�qU��f�)�`���p��8�alJy/}i�� C������	��*�!�Q�G�	�2�;��r�B�߅���~�gx��I���]	r$I(��ϗYa8կ�q�aL �;:�@)��&+QiW	�e\�k�u���1�� �mn��:3;K�eh7��0�פ�@���>k�V�+w���e��_ ��l��`��YE^��g� ܦ�F�-�n_B��7�g����#�n�B�cyiIf�}b��se:�=��ܾ�q�r�;�Z�pOCдjr;�.6�}�R�=�&l(�gL��^ ��G���I�"�Z�בTY�iE�;;;M�� `;p�&��˽����������=���aA��)�� �WV�djzR�x����������{������������`��es��|QpX-r%*��~c&�:�Z��ˤ0 �`G�%�y͌6������Y�7*��T�ߪ`���ЖQ�w%{ T��)�Ӱh�,O
e���~��i�6%B�?��^WC .�A��bV���rR��g_����܏W�/{�s��Gђ�;>�[����;�w�S������5�6�kK��m��ִ�;*]'|K�X�y��kY�1ꦩ\�U��s*'mt��˱�W�����z�X�>6P7Yzq�_�*��`ɽa�GL4ʌ�\ص�D�q�U�'}�P��׍o9�lpЋ�F�g%����u�O.��HelyfSH�I���[���������+�Q����E�'�a�ޱw�y� L�8�3���V	-��TMU�x2��K�JH�����C7˂����$H.$��C��6��� 0��A`�T�ZUL�#�4V���j��#���:{un�pb ݀��AK��̻z)�U�sO_�9�2>6*�(�w��^s�ɇ�������;�:᜻�I�{�-�W����BJ���T-M_e)T��ꮻ��H&2P��쮼}��;G`��ᖌ�����r������G��т1����7ߐk׮��Ɖs��
�b2�Q@
Z� jͩ��N�T���i��$�E��V�k=UD�| V�� Ϲ圻���O�ݣ� �LQ`_����z�2u��o-ғʄ{/��v����(���%uG��x��}�`D���R�,���	~S�@���³5�`���cJ��(�}/�@e8������s�qVf��k���d0�ym0�XH�Xu_��y�� ��٤�{�:�i1s1���U~S���t���4���cp�k�J,��	Hz��sy��� c� ���.����`��B����Q�~����L��8MO��J-�+>h��Mbz�&������-�������*��܏�/���uܒ�0��8�ww���:���
<�u�5����"�u�B]e`��\���5�#��4q�O�{�21�
<��^�.�,U��_�v |�.
�A?e��n*��(�fϔ"Ii��q�j+��=��/^P�ׇ���Hh$�͈w�RO�K2�K|����Yˌ�H��<'��/�� �=��a�g.vv�e}�Wh������Dt�v�o�)���;8�\��d�3�j�b�* �`L���w�5 y���s�Qث a��������V��ޱ�:��sM�_ݏ�L��0��*���
X6����z�
���ρ`�R���._r{�|��;/]�$7o�tv�3nM��ӣ������Z��`�R�Ýomuŝ{��M�:�a_a�Cm�؛1�1��qFp���t�o��Zx��fl<H���(��h��4bEJ�avHfpB[��Oݳ�=���v��w��vk����Ǯ�^����o��{������7�qϷ-fo˓���/��'O�
�"H��n�h�f�w �E��ۛz���@�)���V�$�����y��^�,K���G �-���XaU�T,�@ɶz��x�sb��"�m2h��A&;-��X��Ih��Dez�������d�/��^�%�����'�{��y;oR�����b\F`�D+R�x����L!��el����x�::��b��[IS��u�$o�>ϫ�+���΁�o�Ő�i��Ԟ�'!�4����k&�Oy�x���j�2��x�y��˭�^�;�{����s�U\��Kr��Ylʚz��G����Y�;#��2-�n�=�y�a�"9�� ������;�"1;>e)��MM�)I+�szGg�QC���F܃<7f���U�SDM�lcVk���o4f�f0Q��
]��� �p2��"X�2�8( J"{C��dų�����^�P�������G8b�������9Gj���e�v�Nǫ�/��?(��
������x��3��˿f�\KKr��-�����������r���q��\�67�{�����ewo���z�K�'V*���z�e�;&3��M)I�З�LM�}�-�wD9����E�r7Ph)��?�s���3L]A�4u ? �QE��l�}:�`Z]v�/d0�|-,.���6�
��__[#���~���{���1$q��9�~<b���V�:�3Q��Ł*,Ƈ������z��@k�ɢ������׃���y�j����a?�]�����z<l�	.�tP�Č��,�oo%���Igȶ���4uOKX��t��DR`H���2�͸O�MN1�!_��D�'AG$��/@Zh\c@����Ey|�����P�#�@�1;���'ſ��zvog#(
�qo���`.�l�7C�S)�>*�^�YX�� �ExI��N5bߛ���"R����L �J�����R��Y��Ɣu4���L�qV�Z�yIy��؏1���7�f�xQ�CCÜ����A�4?���`�%��`��-M�9�΍t�'����[�w [�#�a�H�[�����pص�q��W[|  5^�S ���)�5��@��["I��F�^�^�?AJO��g���)����e���n�{�/�G�:�M�Km�Q;����i &GGF�_��w�qtLv�;N%b-u����8��9��3x�`�^�v������̅99t��X[�,(7� ���kY1��`� ���� (����� ����������1���ؤ�Y��cݾ|tt@���2�����1�% �{ΞZ_[7�]����}{5�	�Kn�f~`M�X0��Ņy�w���_6`���8�  ���\��ǐ�BaE �xv�Q��6��ONM�\ ���ܭ����7��2$/��oz8�w��}���JAt��
�µ-I���0�����}�1�+��v]B=`����3�*>�#�n�Z���w��J�l���mS\���v�faA�;!�9I��;�3�`�g.�^�ب�����n��`'l�4-X���U���ip�Xk�B�+&[u��y��M����y�8QF�$���yn&1x$)�t������������ ��4��-�G�J��Ҡ5}����?���B���`�t^8���y���9���[� >Ͱ��es¸!�n^���܉������E�FNy���y+]@�F��F�K0��̥��ű�3|�|'P>���w�]"�C�/��q��/o��9'�9o?�6�ns���t���j��?'ǭ�NJj�Y�ANQ�zʦ�� �6�F� �N��Ι�f9�8M��Pp'��@�̗���f��ܒc�.�/ؕ�,C��@�A�?Rw��ka�Í����snR�׃�`�r~[j7y>MP�
�Ρ����Mw��x-��_X�����ugܣ�_M�1ٓ�ƾ<}���#+�)p�9��zǙlmm� ���;>���r��2x꽐�8f����q��2z�ܙF�7�3��I���`H���>h���4*�#���3Y,��\[u�����/L|�s�82�=!Kwcc��O?�D�<}��	ɢ뗙�i�>��RD��&cj��x����
SV{�386:���9�`dp�����=�H-�c �^r��v2-~�1<S��T}f����=���7.0.���[o��b� �pm|U����`��/^�;w���d�&ƌL���5u<���θ�Z��	�)�O���������W���0�mo_��ͺ{�y�;�F@���0p���(8��'q�Z׽��Cj����k�\�G���":���@���D�y�u�#�e +�KJ`�f;Xř�1��p\�(	���7�{����;T)5�+��d��u� D��d;�ZY��M2G��*��U*�\7�\ŧ�X�ി��(�$���<6		��d(K��N-� ���8�h@�p̤46��?�~��eq3��I9w.  ��ݜ?�zfa��H̭آ�cH�����qd�ϞjUo~�x)��;�to��!���?��&�62Ӥ|�������zp�g?���Ar�d�Z�#����vC�J��JQ�:c&������ޑ�Mb{����5����,�t�(e������ 	�[��$�6��ڲ���I��~����fjÙ������m�X]���]�s�+ \\� �0
��Y���I+5f���HOϾxe�C�Rɹ�a�����Mu���P��s&Q�������� ���m܋ ���()$
�6��֌��uy��h��c���Ǹ� �
�{��X�[���1���&|n�2.�q=8�=����\�x��c��x�d�����,K��w���Ͼa�D�T�R�lᝢY��ͽ+�̔/1ً$Iº�����Q1`�Ryݷ�	$%	(cl�-��i �ʁ�\FC�Fݻ��1�qT�r���+���ܳ�úXd����g/Qb}������y;ogi������fS��>�ڬv˚�{l��b ��j^�lWP���u/�䫟*��a���o�/Q���Uͳ<+�9��_�y�~�9��}�D�&�n�s����ಗ�	�,~_�l}T�� N�uĭ� q8�;2I|L4����	$�Ns��s�1��V�Ț-4�E3�.��ܞ�r]�Q��m�_'����ݴ���_�?�#����fn�en�0�,E��b���^�XT�U�P+\�)*�jvOI\l�ErT��$�Zvͪd�P�s�n�	&�1i���`l{��� �6`n��pv ^"��n�v��B6�s.��>: �}j��"o�Ӓ:�cc,`�:�v�!����#�w`�Udjz� %Xm��=JXlmn��J�U�d�4ɰӐ�A���o���sy����{����T���n�P����3����i�ޠ�_����^��p�,U��c
��(���9�
�C"�ʐCj�g�&}�'����c �"�s�9����x�\�v�� G�/d?�.��BJ�;�/~�_�޽Oyޟ��=�~n��z���;�����	����Ϊ�:c�� ���f����]��P���R�Ucy��_�G�)u����;��S@
�� ��g�e�07���,dt�1K-ي:u:�8GHK��'6�0430���v�?���[�J�mۯb���	slhp0Ҁ-�ȧ���KY�y1�_�gI�`��s)���
">y"W�^�+W.�O�w�	*ws�O>��~���3֝��q�1H-hC�����~�8����k��yg6��?O�ѽ���HMϗ����\8g�����^: "�AYŅ}��ᤌ�9�E?�)<C���K:�\y@e��P��,��5�u��Lw|.I"Y�0�[�E�����@��?zD@+�{X:}��S�Y#8�D�Wh�#�\�a��j�D&��*��Ř�xB?�B�i%
���Z0!�/��Z�YЪ��#g+TR_��m������ł�`�K�?Ⱦ����.u���&ʲ�mO�>�~1
�^�z��&��Q�<��at��4��%����p��L �6�rr{:�c�k�ˬA�̞��M��R�.�cA[����D�����Ξؓ?��ܾ}[.]�H)��3VVV�F��f��u����ø{Y�J/a�cng{��e؟�]�&�Ã�� ; ��>/�s�C�>��ghO�M��W��:����o[�mgCl�y����s�D��|��	�}��E�{�my��� �^{������;�F_]ݐ��J� ��w�^�� ��
;b=�|�㋩���_�������Fu���m���B9��f�U�$�[�5�c��&���,i_ XD�~d�E���@!��	������ȳ%io�k1sE�����>�m�:k�&�곭JQ�)8o��[nF'��#����>�k �SI�4�ݒ$�Ua��b���F��.c\�3�A�il��dT`��q�0Me��@��%bs��%�-���]�s`�+�䌿{�g-R��,\�ؿa<�hݵUS90����Є�8^�*>FϮ�hS�Kw�ͨ����K'К�LH*ݮO�q==V�����Ȗt,n�����_�}��l����o�y@ �98R���'�-���{����_�.c"l�ּᜤHP���Ŋ�0��%|�lO �ܔ��WQ���3 �'����lӰ�N/�pq�t �b;)�9�ƸUS+V�b7`���9���~��w��������IEӽQ�ݘ#����l�p~��284"SC���F �ʔ�=��^��aw�~���Q�U݇�#:朄��a��m��j�hZ�O�Z![�Z(����qׯ_sN�����q���ij��4fr�����j��g��<˰�%�����2�Ċ����L֢U������OY\�/����<YM�)����+�/�[wߒkW�����m��3���������_�W��O�����;���+WD��~EmD0��榩��g�g�+Z�S�(��V�����1��pnHn���+@�d��O�=�ݝ�z�*u����3�0������F�|w�K�dƐ�fb[<�����D+LT�=:wU�Sba>�u,x���%�6���?�~�D��.���(J�_ɂ�܃�Aj�M�q�g{��{+�c�`��@h�-UG�9��$�di��<y6#3s�+`�7�r����uYI58�Vxꙷ d[�Z�`�%Qq�(52���Є��1��s�m�����η9E��̅W�J�;(��4"�֭�>�g��F�i�M���z�`��x��H�UƤ݊���7�MDb����Ȧ�Cg��
 �Y[[��}Zi�k�r^'�����,����?�8F"����������
�Ѫ��K����Q+8�@B�;�X�DcA\�&�q��Q�֗�~�ْef�1�o0Nt���
���j�����l)��*h��5�#������=>P��2w�Y �
dX0w�T
�7/�{�+算��|p7�� ���Z�T�ξ���fPwc}S~���08{��m���e �5<8Ƞ�ȈV`S`�S��0}:/�� ,�qd�������?�a�'};����	w�����ް�Ma�Ĺ3f5������F�k@��
{R�ʾT]���1p�J(�Xk��C� �!��}��Z�گ�.ڱ�	 x��&l���q��Oޗ���:�͍m~v���s�.��F�7���R�Ldg/ Ў)LM��c�9j|��0���\?5+�@;��Re�{I4_���I,�`���b�
*�X�3���	����6I��5(s���ͫԛ��(��g�G�F?>nq���q���;SB<qE�t�X���]���v޾~+� �y�Hұ�M9zL!�-a�-���� �gK$"���'�ǋ�ⵝ�r�X������k��w�]%����~����C;��RK��ߺSЕjB}Vec@Zb�E��*�Md������j9R~�'����Ƕh�dI�
�c���p��I
c�߁@�Ũ[/��{��y��ob��.V���5��o�%~���''�0�8��R�2a1M��;�X��[8�E�:/,-q����>AZ��Gd��l� �������������ƍ�yr�x@�t�*��ʢ)�3�(�朗f������5�۵�N7004�,�e
��l�f���
���h�X�ǀvBݻ&t�jt�&&��Sq� &4|��3f��<"�3�z���Ֆ�զ�L�gFe������{@����M 7�^�G�U�f��ƚ,,���QFm��	Ha��N]�w�c��؂d���J�@f<5�{����"+��k*%��Vg0�e���������<�.<�//�_8gl�=����ơ�Cq���~��GGF�cI|�1�W��y����>�H~�_ɿ_�zU�}��k��������u�\�~��Y�n����ۥTJ�{�pX��[0.P�B���v�b;�J|���/.ʭ[�q`�.--���}�m��h���N�b����UʑѹD�@��%I�($�Ғk��>9��^Aޭ(%5E1��v��m�b0�����9ՔgeK�DxG-KV�^��5��f�tv7rթ=�h/� h���o��J߅��������vc�,-�������S7P9��.���Df`��B~ �6�^|�E�J KQt30��l����fz浬�p��."�\��,�̀�p�1�̖� �	.���7`t�y��l�^�T8�P[�Ş��A�m
����k�����V
�یF�̞���=ʷ��K�������*��܃�#�Е�i��ߓ�������S�~��eZ}���,��[�̋1��l������OAA� o�����:��S,�k�w�����ڙ��ZX��HԢ=a;	ן�_jA. �Y^�^�ujxx�{ص`��8J ��
���Px��ӊ��H���y���`O�\d�  ����/X��ƍ�23;G9)�087�h<�k��掙�m�ׂͼ���w�}lhx����¢���\�vխ53Ζ��p~e�Y�f����ۯ��;��:8<
����4�����$%��C��Sj�ê�qN�4�w�BzC���btd��L3�ܾ���A;{�40ˑ)�=6:JY!��O�Hn޼�l���yW�6������j���n��-��ឳQ��Xc���B��>`� � �6+�ݽ$ TX�ﮟEsg_�8'�Z�l�LNM�fo?09h'�V,����S��F���P��6H���LȥKs�8e��	����H�2s��\����)��T	1���|v������4����w�78<(��}R�Qf�삡\ή*�ӱ�+�1�j�%ĄKA|_S����`����Ae|�V�a�~��̰/��8o�`;�`�(u�4�c�e�:Z�.�Rll��C���2���.� ���yK	N��@��+�_xN��<�H"D=	�y;o�f+En�)��"�����c��8c� �Y;����p�n���o���I"�82<(�^�[�+����6�>8���Ρ:�����z���GZ��kH�-> �d���P���ʇ��[:c�t��L��?��:����B���=�~��O{�{�2�����}�SN�y���^@�=w����O��?�u�8���gRi������Yd�E�YXXb1�k׮˛o�Ey�s̡!�O��l�!�r�Ck1%В�A�Z{V�I�8'Q�Dp���	�������<y�T=|$;�!C%{f�Hf�C:�H'F�������/��?x��Яmw. �w߾+o޽+s���>�c�����l�w�����Ι~��N0}nn��D�5Ӽf�w����mVҠ��"�����m:�Ϟ=#k)����a�=�@�܅9y��^�-@c8�p2��7��1�'�d��xX]�=Ӧ%�}L�SP��e��d��}�{;�pp}!"���Cl���j��$��@ �^��\+4�=���d_%!S�W*�� �&�����EA#�Fa�4A���]�.{�$¬}�;�B�-c��:�##�J�f,-/�5a��h'��� �Z�σ�s�;R�7���`����!�� Ӗ�E����I�9��X<G�m�dC��[M�y���C�57���|Q����)X�E�����>�$�X�:��oܼ8{��Ej�c/P`_����D6a3��Ԋ���<�s~��Q`%ǳ_�v��K��X�dEn}��2٠�T���	 k����^h�V�X�haV|���(���7� ~_`E�T�GT��Ђ��bf���z p�3 �����)�i �G�9�g6K��n ��s��F��gW�V�:��4����$����m���&������'�\���s�اx��̵k��>�B�W���|,333ζ�������n_wc����؂��h�p���X�ތ��@������<Xym��`�OR��e� ��(nU옌FU%x���k�f���;dŰ�'�����i;�e�k�ڪg�K �:���o�}K���{>��������ߗw��)���+2?�B��4�Tƹ&]�!�Lc����j[}��$	%KY�B���Z��������
�B����cn��m�)���Z+��h�Ss>��!���epX!��w�L�!��-M�e��ü�1������E����Ĥ}:��.[�y;ogn(���Z@86�����S'-�N`6���I�ҭ�h�������t �����-���m[	��7�|�9h��n������gն=��lA�,�t�|l�ZnL^K)��.�h����'�ũ�l�O)Wp���9�u|����ƿ���M��}�-Զ����ub@��9�h�2+=#� ���&��T��	f��=o4����'Y���-i��s��JN���g8`(�22rH_�ǔ�q#W�����t���*�*3I�:����O�<��/����1��NS���W��`V���J ���Ƈ��u�ߍ�}����t���c��Q�^��?<��[q��9��ƭ���_x&k�tHQ�,M4ݱ�R1��ݺx��-Ǉα�ڐ��5p$'&�L�*=�T�Rlw},DV��[$<�tۙj ���{�^���&\�q}͂zα��W8e�V[��ZA=7Q�\���7�x�z����|kd��ϐs^!'�ƛ����=���3Wh��8����4P��6�2x�qҢKm�=�)�L>�+Z���O�z: a��/� ��q��08���ם����>����; ��t�#�I��3��v�
����0�RefV��xۜ��UwO���2`ٽ�Iw�z�j�ŷ�X~9���{[ap{��ɃTf�8'�i8� @2�Y��A(������d��H_�<{��F)���3�|F�{�`��(��qM��0;��a�[ .��
�5 ���\_�2c��X��Β���['y8Qbk1�D��=���8ϢsĤ,q���N�@���ֵO�����r;=�*�嶁��z0�{i��Qh�O�|R� ���l����qRJm]T'?|��ɾ���n�Q��#�iU�3���:���i��'?��ωIˍI
�h����y�|�Z�Y6j(-xH	$�+��7�#�OK.N���hyx���k������Nſ3����I\�{�&� =�
 �I�Z�C�J3� ���,1�	���e!�`G�{y��23�7��fK�R��
�/��`/�p�d}!�qeqM>��c��>�ӟ�D>�����62��q/��0����++�d�b��ݏ 0 �'�S����3 `�>{�\d��Ս*��:�^r,�4���D �!�����cEv=���A/��,�9��#�}��Mf2	�p>�4I���%aa}��a��~��uJ C.��drrZ�&f]�;�k�H��V�]�������%��x��fxYp����=/��}� 8�hT��G�y10�� ����qiAzosyy����pE8�"�_�#�DTg=��D��(�4t���U]_�����B*-$���uv�� k?ﰳa{x)O�(��^�U[3Un�R
@�%�V��v޾Z봙�w<ԀQ���QfP���+ѳ���G�y|qw�Li�X�L���5^N�_D��!�ɔ�����?�VLa�5+�L�Ɲpå�$�z��$o���������Uy�h_�U��Gҩ�����l��tky��睺/������Ͻ�c��x�YD9% �9�5�<3-I<h�>VԆǂ%��^���<��R��m���H��Wsfk�K�9(����n�����Z�(脪�I8�0�=3,Pe$��7��2�z2x�]0��"�fa~^6�c�d�9]p�����5��W�a�_�Z?�2L�Ω���]�V�r�^.��W���3���pO���������֭;��	����NNM������9g�|��'���N�T�F;���9��Zu��w�dsmU>��3jlNNN���� f��d��Xq���x����7u�[�c9n(H����?%;̥��5� b�D��b?B�c��#+��}��%��O�%)�[�d����9��}K�|�-��xQ����{���C�oܐ������sV4GUw �xov�$}QE��qנ��Đ��p�1>4�Y;"� �A���z���e猂�6���Ӓ_�zG.^�#`D�U�tc��{Jz�l��<��͂��T�^H�ؖ�A����� O̤^�m��!+���j���E�N��wu/B���8�D�}5�6�3�W�xS?��a(@���4�e8w�)�6���0��)��D��47B�жĘOM�@�4���*�s��b�A�����ċޑ!82B�r-���5�Z&(�����6N�z��1	 �
��I�y ��:Cw�qР�x��N�˧�E�~ʥ`�b�
� |S�j�b�{vf.���I$��Z��
��I�	��G2Н��A�\
�
�C/���  {���,s� {&al�)u���E �/Ƞ��2�O�ZA=ϐD�`���g�V�l�͑
��=l�,�JS�˘�`5��NV�x�Є퀚�1�}@�?�M�<mZ`����s/^���I�Q[[k�l�/H"���P'�����#+�Xa�6�wc�y싔�DFՂ� ߸~���տ���>c�������~"}��4��s��q{-���[�|�u�s��˫++��&&ܜ������v~����<ٵȆ���$8�bx�y��Ww}1<2��4b��C�{I&�驄,.�ߺ�Q�J�v�`��{B��*�5�������Y)����J?���2������5���x_W�\�˗/��f.��X�\_ߔg����f���^98r�s�EP�����l݇��%*yI0���#J�a|,½--.1�ޠ�f$�6u}�b-_�Vxnʸ5��i��JK�2Y2�� ��?��A'�V�r�ws��vm߸�W���u3Z�sm�˺�oɡ��l�zmt<�A�6"�޽dG�@�k)���s�}7���gc�I�F��[@���x�|��p/]�l��i�9eL���2�#j�H�"�bT>-+���A�s`��0!Y���4)"�	6de�dyZ��G,� YX;I�L7�@n���qd.H.�^^��b?��@�%���l�Y��l�N����w�8l���@�1�-B�ܔR��3$�h���>��k8�4<J9XA��UJ��zsÖ��̐��r�����2.e-��L�B�U� ���q�N�}�'��zR�5I����Xu���z��Aq6 6  �={N6���K���?�Ң�P,�biJ(*�nfi�ug���Lӑ[�o���������Ϝxq�ܾs��w�c���G�+XB��c22����߾��!%/�w��4�u����̽c��i/�qxp�Z�H��U֐j@��;�����q�WGX���C���)�ϟ�hf�qV��CP@�s�iJ������M����E���d�{�r��u2�V����|��'d"�w�/��ު�k �pl��
��pp����3�� ��`�������vt�}�:dQ�}j��x�7���>�\�7�X,k�/�8ंH��pH0��www��tȷ�q����{�Ae$�3�N��n&S
�W�i9@p ����:�㫘��LK�!\�K�"�_�i,֖���w�Tb��'�ju��cA����߹s��%��=��RGA�k1E
𸋓�)�������>k,1Z �ڂ�L��h��if��S��ȴ qpX:����Y��xyOu�%%���#$���,\��_�8w�1H0Ʈ���#,r���I	���m�l�$|�荲W�����^�̾6�S�Q���nHv�L���&/��)-�B��΁Qú��k���k0ἡ��ժ��Sc����Ww�<��C2;�;$b�o��M���!�V[�����5�	�aOC�;� �.YF�3Ms�9�s��>W���
�(�0<|�Xfg�8_g�g����ޮۏ*G6nZ6��Nk�U�Ui��@c�7��<��>���q�ֽ�/Ɇ�{~�_~���A��ܘ�g��s���r���=j��y��e�,
��Q>� s��F����%�)���_`��Q�������q}��p��3 96�`� �x0�}��i�Ѣ�T��b�]���%�s�qv��1g�$,���c�UxVd�΂|�_��_ɵ7�/�l�����+���v�l�+]t��Z��w�g3�mςW�bԭvXS�7#���7|?�\�C9p� [r&`a3��P�{�ir7��5�[���ۊ���y��H-�L�Q�@�����xP+�յFA�c��F=�E�K���af-���i('0+�E��a��TG��Wrw��y{e+���o�e����R�<N� {�E�J;��-X��m��z!� v�� X������V:�/$���A�K;��-Q��/hd��+#����AY^c
�ك�b��\��mz�+�岑_ gT��q��v���;0��n~z���K=�M���y�ﲁ9��Q4�*��ñ~\�q���\|��D�jՁ� jdVR�Q�N�IdL_GJ?�:��b��m���  ��Ѩ|�XUu<�e�)��.�B���|�^X�5i++��L�t�u����g_��|�G#1�Q)�O�=��i�H����� �*������8�#�rx�ɺl��z�¬�[uy�bAV�#�O��/���#�����tN�����tJ�
׻�z�LOL��7ﺟ�28P'�|p �� ��]ߢ���C U��*�j�rt�k,(]3���<2<B�΍��N�(�
� +���9�N2�pR�b�����Af�j^3�E9	0�~���

�9��ڟ|�)����[�Ȗ�cs��O���gd���Sg���s�gfg�0��6��pj� υB{x7x|�NFsN�uO�S��/��u�7���0SB��L����zf��@0	X|�I�+�j��8�`�ñ��@��`ĉ���g�ϚuZ,������.�]�:2�A�9�y�#��a�LN�'E�*��ė9s�%�$��,1��@���w�}�ՠ���W��
&]��ﵨs�qT�&ſ;��$���z�*|ѵ�k]���3��w(¥�m�-���h�s�'
ަ�i��rN���h\7���-�R�����~T�:$�lˌq��ۥ��X���`R�4�{�����}�j  t3��|���S���D;w�!%x%�'i')��9�XQj� ��4��hw�@���,�'>�`\�^�����gM��H�ւ$�!I�2I����������P؄��J{zC�a�	,��0Ȋ�N���$�oQ������lި]��{�`&oQ�iy��\D�ͥ�6�b��'$X	[����{��j�`/q�Z��Ο޻Op�Ћ/ğ=}*O��	�0-27�؛�E`tvfF��<��0�4���ލ��n@���E����Q�v���"n����ؗ�����5cy�^�-��L��:3�T����X�|`o��XðUZVύ�ǿۦ��@q���1��L�u�6�	�۵@42?�]\�r{��ecsѝ���a	YM���85�����d�_[��}����,����M�>��3�� f;m���v(Al��ݸ���{0����)y���1fgU���$d����Q��WP���W��wp��*�B�Le�H0��]k-��׬���4��a?��	�M�x���l=o��kas?M��M\!� Bufɽ���&긶H�/��0E ��S��\IC���j���t_E�;�>�α�d;���ؐ.'���`L� �C4�(Q��sUDq�b��ಁ�g��\��I#�˸��|j�$�u#x�j�͹����y�֚ihj�6h<���J���J�@2�*�V/A����\�LI #���E5i�P@����G��j��]�;�Հ1|�k�@�d*!����ӣp�Z�Q�,�-�����Y���J�P?om�R�,���!���[2�b�ڂ3��xϖS����麃����*����~C666�6�}gN�5(����'������O�Y>���lm��_��LL^��'���X�6�D���朡C�s�\�2-��W��/��?�gϖ�^��r|d�`2�94�N\o0VXL��^d{k^5Y�.��Y ���������ElZt���|��7HG�=�ua~A�_�*��yC�}�]2c>��S��O?����u붼��;���C ���O�7������ɪ�����8�
ĂE�n��n�� ��j���:Q����k�9�{����@g���?`�ݸqM�{������� ��?0������>�U�c
g}sc��<o���n�L.]���y�O �*���A*flR�8����{Ouɨ�
]�^��fM(�pO^Ö���J�?��s9uf2B�x��=[4I�"6�R��T��O�`� �e�U�9��}�UN�_M2�J��?��Dd�'E�`�/��F,��w���)vz�=���%4o�� @��8/+��S �6AwMG� 4~�v�ޥpz�C_�jqV���8�n並���?�12�ݯk|fe0#h4<<���n�6V-��B���I�_�p�����'V�S�G��p�j ű�­����b�����0}��z`�T��E���ּ�����xɎ��Vh��V��6��T����ʪ\��h��x�/ߤ7�y��	.w�I�(h	���d�+H8�׬�g.Ǎ���4@��ځM�&��A
�+N�:)�I�L���WJ�5��>�+�>+s�3�?��_�sW��<����'�`��0���8�Q�S�QԸ=npv���ۇܿ���'�7O�g����_����OȄ���e��4�1����ɋ�n��.���� ��?���N[Պ�������y��\\Z���e;�A>썅�V=����c����nM��  �4dw�)�{���s������-{����=��o>�	�����,kJu}�gv����4�������Ǭ;btl��FF���[A�j��͢�Z�Cm&����O��|��ܹ}[���o���﮻F���= �|�ҳ記��u��F�`�g�$��f���jUS+i%hc��>����aSV��ey�٠k�r��(�h�>l�t#M�=�HZɥo�G�>��k�4�pNc?���Sf�����`�2�+y/��"�Mn#����y�c��֑3n��������g���i)���He�*���/���9��#i��X^RJ����� �޸�B(�)�;X`��R�9����{�* �b��
S��n+UR:TJ~�ǖ��R�|�^輝�o���WE��B�<�c |�4�	 �)�`�-FJ��M �"�ݝM2;_�x.�T���R:ԭ��a��c��"_�4�O�)�����@L���a^@)�,���w��g�Lgf.,#��&����Q�'���s+��`�|H~P� ��0di�^�whpB._�$w�ve��!���?��sv���F�C��k�A��O�������~�sN��g�=���c�\�Z�0W�i�7�d�b}#3�
���>=Ρ�n��T����9�C��8FS�S:g��5+r��S_�~���\>��w���ϟ�`I���������d?|��sh�@�d��ñ�y��4���I�^ .Bró�����w嫜L��f���lk���?me<!�L���s�4��������3�p�ܼy�)�Jj�ꐟy���졐ڑ�-��#��.\ �����jl��QU�Wnj�?�-(\0�����g\0������q_���c��D�S| �{;h������xm{�=P.���2��I�.�U��跓�E��
'&f&��L��{��ۃ�������>I+5���ׯs|!��lK�(`g��:��M����Ԗ��F����7�"˨�;:����h� ��O���sk	��q�N���Y����@K\�
�c��KҬ  ���ɣ�X�����G����t��W5�YO����L_�(�cE���[A"��������5�;k���ǜ���隅�<=z�~a�w�G���>D����� K�7� ,ƙ�I��,: ����ߦ���(��#�����'�ȝ;�i���Rve�m�Z�x^"���3�[��r�( ��<~����o�e �]�-���N�cqq�=�e(��#<neu�{��׸Ǿ���	¢�.@X�	08D����b�����P�om]�V�AjYciZg1Zφ/4�Ҵ��M��<oi��4	b`O�9]���ox��4p^!�R j66��}�@-
�Ĝ ����5P#�����|�D�a��is����@����y��'r�V3��T.����ܻw_���y���������LLNʜ[�*V���l���U�De0*���աn�MZ�sd����jټ�����5��JJ� "m�<�O̦�r�]� �~��y���}f4��$��eǔ��]C���24�˸L�y��fFV'EVQ��NP�bYE5[3+�[^���/~��X�Ѵ�H���R�2�L�$����rm��Z��gI�Oy�3�2q���Xs�ˋ@i�؀�3z���
�t����?_g�۷�<8������MU�B#�ﵜ���.2������� �3(v�,,(�WwF�������a[|�4���iЁ%|t�:�d$U��R�H4
�Q�w���@����X�`��̈�.2�>�JdyeU:�>���a �n�he���5�r%U@Y��?B��k�Uh5U��oݺ.����g_���#��_;�b���`=����\J�  �1w?}��dz���Lo���#9>j����;w�U% �1˘�{HG.�Rs��l4�^  GZ�T &��K��	BW����Y��u�8?<@�E]�/�T\�x@�qlt����gO�����+�׿��� +���W���}��?��Oht�lo��Cn�B���"F��g#��� �&5N��ps8�4M+<�t]cn���nk:=�#2���qw�~2�����07Kv(>��a0� ���(ꧬ����K���ŋ���ǵEDJF�g1H�Z�7���c�\?�y�F6���) &��B��K��Cw�7Y��e��뉳x�����P/ v/�P�������^�*��t�9)^W����E��_���X�����i�w�B
;���Ξ������ SS<J�IQ^"-�o�#n
 |��D@�%`�/�G�h�Y1��J��ueʭ�S2QS��2I��ُ]D��8oV�o��`N��;
��g������k��㎵6��3�pJ��@�6قP��K���2�x0�
�s��H$+�]�'oŊ��� �(-���(�D�_�Uo����?��P���*,S!/����{�LT�ڔ!�Wh�@j�ѣ'���/�Ճ���/q=����Jt��g �	�X�!�4��Dp����"��k�T##c��o������O�ǔ��=|.���?uk���e�]��~��pY����F�W���ybE~����(h���)|�:7���S5�`I���n����J13S+�}]e�j@_�<�|�d?��/��_n�?:< �N���@2�,f$�������7��sMA"�{4X2�V��"�����	"�XJ������ǽq`���p����0���>,� tx�	�y��ʣ�(��ڼ*���a�J�@	΁>h�m݊dw�:{�E`�3%�[�g�&��vJꝷ��U�����JK�����=6>�w���.H:#���H��$}�"������r	A�P��n��>�Χ����?��7<�v�bv�F�����|.�Wp�|�@"1��U���I�O�X�[�;Y�|m��@Z�;�4�୔#m����v޾f�)�'�x�1
g�E`��.jC�|���N���Q@�5!�R�Hc���I5���%w�C��Ҕ�� ���u9���#e�z-h����%���$0��;HаB�:��WW7�u7ɪ���(�;ǲ�}H�����!s��	��d@�?�L��p����!�CΡX���E�.M����r�V�|�Q*�����������K����_�忓���Z7޴��	���q�ڐ�^�sϙ���C���ؗp� ��T�JJ��z5�7A�����Q� ��z:���C.H��H:�?��;8�#�㔤�cg�"�C}233��G�������X�9F3����6��7��{�'�߹#����?�I>����/�V���r��W��,s����� ���w��b�ø���"c`=���563����`8VՀ�Tuu���t���Cp8?��S|Z^�yý��7>���yH��V��r������V$��qw��gE�*��*�՘��J���Y�����G�y^|�-/@g�W��k~��ړ��ZI;��x\c��ɋ"z�q_�>�lw/1?;@e�4�����[I��Y�ʢ`�c�57�@����u�8�!�QKT�TF�������/��u�sd��݊���A�z�`.��3>>!.B�t��gｺ$��4A��!R����e7ɞs�{{g��_���9�2����L���v�3M$�P%3+�Έp����{�GDfeA���u�22���f�}�-.ͱL�0v�s")�����#��c4ڒ�tg4�%�w|��u�6�����7�')�V��RI�x���j��X`��������1����/�lT�{�+��%q*ܗ��pq>ȣ ��J�~�0/���b�4�cPv�Q���+�*�Peº�lS�s�Jw����ᜋ2UO����m�����~������N��z31qJ>��,4u�*ӄ�&��m-x��DC��s1�Q�,׭Y���6�G?�+Z�t���o�#ݾ}�~����?����O����.�'�����i�5�Ǿ���=x�9����sY����K�����z��� ���y\�NCX� k�&������>X�F4wT��]�33�Q�BT��Y������;��3�~r��!��R�&�#����E6�N��s�N���k<�L1̋KKK���� (������ⵙA�fCdb���u����iF U,�!Yr���J�J��$�{�Ŗ��{����=~�~������"M��;�4\���\!���|�`s45=#6)���������&�G
�6��S�!���|���T{��YvR�!�e��rЌA%b���p.�p ������X�ʳ_Fm��kg����e���-T�{�l�I0�oQ3��$��E.�vu�r��c��l�d���̖������5GZ�O41ꃽ
�h"�L&y|s�R]�b�_��˰	%�L�����Րm��}n��4�����0\���T��-�o#1j���AÄ��,NOs�
�
�4h�VԜC�X6N�d�NM�x+�4ί��T�+��`�l K�I����$ �V�@6+��fJ����zl\@f8��:�׶4D������+�3�J�l���`Zd\�Lq8@�AA�V��"���l�n޺읛���駟��Ǐ����G��`�]�y��Mv��ő�MN��;�G�}��3�p��s�C�1�>I���� R��|��{1�Ɋ��g��&�3c9���_�hg{���_p�'F�8�Ғ�{Q��q�����~�p�VVV���N���w��?��;��t��~|f}	e�eR �d'2�m&� ��2�[�Z�7pNHmitk��#��gf�l�|�2}��G ����{���E��x��9��;??O������тMJ�ɉ�+�ZtGt��l�����8��Ǟ���[e��/����hc��}�kFdiEc \�ˡ�i�s������E߫��Fʦ��S���Y����9/�=#G��3J�M��Ύ�EW��x��q���i��W.�E�p�4�~� ���Wg׼�N�"w�޿����B�Z	�Ơ�#� -t��;�Wy��i��b��0��n����*�ŨĶdpEפּ2�l65��~��
lf8E���hY��b�M	�rA���"�~���,g_ِ�wο���]T�Y��6d��}�.���)�?���� 0�QK,���m$LN���in�>fZ��j�"[\
flA�F�2d�.��988b�4X�WW5�u��Ml��A��ƋԮ�m���ݼyï���8�O?�����`�C���=6����Z`]��8>�f�	R^X����~�dH��ޡ?_c�5�ɜ��.�U
QU�Gv�*�pkhḝ�mfv# ��w���n��� 0˰�&U��Lj<K�M��b z����~�$1�5��m?�ccm9�B�e[�����)�Ů,t���	��g������O����_O���3�3l���F0��?\�ׅ,'��Y>$��mN�ҵ%i��~�+��kF��u�)�G�S�{�hgd˺%�߂�0vc��縲���gƋ?L��Q������>uf���}�Ƅ��4S�2)�p���?)Y$�u����ϢL�9��j�$�:joA�o]��#V�F�N��
���T8I�uqa���,�d���R�������m3���9��^�:�i�+�ɦ�Y�����r�F���M9���}E^�7�l�)uTP9��f֐����2+�� 2�X�k�̦�c�Fx&�X-@)T�+h�UKkq�{���!N\�nK�_�L0�����*Z�0�'Ƨ��ۡG��$h#N7R&?���TzY��毷��t%�S
{�(`��a���)��~��W�  �CIDAT�v�G|�ٙYk{�b����0��O����C�
��OH�s�ff��A*���͌��fc��/MЕ�'��x��$^^Y�TS�#6�L�˗��d��ד�� a�!�r�;؛���sĲc�q�8���{Z�p��M� "�p���!�` ���6y��g�)��:Q�f�;�����/���޹:b��_��g�����glT�g)��=�	���̴�k�� �)��3�J�`��}`I�`cWu0�uQ��'�н���^�����$�={��7�'~^��8 ���5�7җ%U7����cՈ���r�֑4�I��Ԑ��l_LS�ͽ��ɸtU4��|�憾S�� Î7�X*�vVD��ړp�77��H"Z)����{�9_�%\�6 �3��F=p����}/�T��͠!���Fl�e*Av ���5���Y��c�?Ҿ��_���y���y}����>�>s4��T���4P�L�[7o�M?��32�(\?��\5�x}�[�d��o$g�W:������т��d۸t�uC��o �d���Z쌵�3�eخ�Bq�~�	°rJ/�靡d�}ݭ
 :X��~�s�mLo0�p�������_�'9H�������<'�
�a����?2�d�� �tA%s��X_P���ψN:'�ӟ�د�Kt��z���� ��䵴�l��#z��څZX��4p�Bv��<�G���~�yr�޹{ݯ�K���3M+���	}�����M��2�Y��M�v2��(���3�4�b�q�&��8d� �c�G��:	�f���x���â���d����A����n2~#h��h�LX}��2�>{�,�9����8�%�W ��u˵?�q ����c2[��,��b'� f[WU���@B��˲e�p=PþY�������#�ÿ���<��8����DB�\[�ܷ�����0�Tq������eM���X��GpϫJ���8$�o̲?:�d��x�Ϙ�nzUq!���L�)��G��l)��v�yHFj��#4u�����b�d�u�9��!0q�aL�F=�b���:joE�okS&t@Y�J�0�K0��
���헫�-�`v�o�휌ꗏoc E��,�ݽd�}����̀!�%��7fK����-�Ux���;�X����n�D�E��dfVe�iy��[b�6����׍|��މ��q��'�ִ�Aё������V㆑��h)C�+�a;^�3u�����SHC���:fi�=� ]A�6α�,')%c�(����}������K m��<���℉CU�=��z��O0�VVޑB~'���}���7�AB��޻������>��O~K����1��_�O�n~@w�C?���ݥ��	M��j�T�i� }D׮�C{���7?��2(Gpe��wF�X������yvt����8��y��M�k�������{x|t�:�Є�����ǿoߺE7oݤkW�j�u���~ώ;*�߸y�;��� ��G���/�гgO�0�/~�fT������Y
H����a��gH_�'	�$<k���'0C���2�F����X��`�=��2��0�/�N���/�C����9�Ǥ�|��39�����U8�(��]�1�Z<;��`��������I�_�Ue��������Q�V��C���p�20�g��RTī�R���vS��V��ڲ,��T��;�Ů� �"��W{�^39h��@c���_+����8��Dr�
�F>C_ŘA�(�ss3~<=�1 �N���>3���v�Q֛:f��6��IG9��=��pAC�5:]ɋ���jw��@�ׅ `Ȥ�=���1��O1�(�7� 	$Z{:j&KL������/�5�����W��S#A\�O�c��<K������z>@1)�g,dW�9#�Zc�.bVi_������l�\��m~=f�"YC&υ�Y%��猩Vƚ�[[����c?N����~��������2W�_�*7p�RPb�48�-��OD[_�������f�>{���&49���˳~�^��?��5��u����咩� R��f+���,� x�Ķ�i��Sz������v�� �~���W��x���=�g���g�igW��a�?~h��SK��z�{�ѭ[�9�u��1ޢݽ]��f��4�����-Yl1��R�RTx&w/���j0���R RW�\e��/66��,�����9ͤ ȅ��q։[�M�]����_���眡����P�u�I��c�N�O�2ײ�N���3��V[��+����ާ������]���H��?�Wz�����pVX�V�<�ya�����,�[7or���K�+!���`�LQ*�%3 LZ:1������0�Q|�����`����̋9�4``��0-�r[^��2x�S��)2n��U�Q��)� .���'�xNm��e�Cx!3�곗r{d��i��O�%�,����d�<��Uj�d���p�7���巸�����cO�e]��=�8�hp��[�.q
����8)�uS::��gw�$8,�錻@u�qp��P����=oo�y��-F�W�_��`�����6����n)o��b(� ��{�@�`8;ֻ�SG�S�P ��P�<�3MB8
��\3\���
���<z�)��� 8�$A��t�L�`]Y	K�����>�ܿ]�y�����T�G�yɎg�	h���{���L����H�*�47h�?�`p��9����{g�	}��c���Х�ZZ\�y��qye�Χ����ʕ�>`�8\����_����t��3� �������~#Wn�U�)3raq����W�\��v`G���K8�vX����5���c�	����K���S����S>��c�33�����OH�E?*zvr� �?f��g,.48� �g�f��V��i}��L�y�;��;||���|���������������@�Õ�<�J�I!�h�&�Q����� +�S��"X����A�?ba;5�S����	�
۾d-9��C�X�`�u;�}��xԿ�^��<~1���>ƀ,��815�����@��.��0��F��X���)j4Q0t�Y� r�w�J
w�n"�i6Ld�X�ހ�<Lo�9K�W�v��L� �w$ޗ�j�-��Z!c��������"LIJ�����{�ItI5�d[f蹺U#T�fF �Ǖ]�­�R��/i�s�{!��V� `Qԃ�B��e١x���S+��).��M����{��hV�뛍�Hm���,yQ| ���>mݹ��-���	�����9]�!2" L�8>>U��I��܊�	���a-h��~.z����X �!ɥ7�ыk�����\f �g:9iRa���jb���Ƹf���� jG�C0��z��	�Q,�@����"MM7i��m�@��{Z��T�6��I�����T��=�u =K.�L�&X��W���Ͽǒ'���k�t��]����׏� �
��!���?|��G�����ݝ�ޖ�� R$���F�ۭ�����U�R߻��f_�l�0�K�?�\O�&Z��LeN�j��ǅ,��w������iow��4�W/���Y��&���k��=1>E��� �Iʁ�������p�/��Y6��}^E	�,�ߊB�DaR���L!c;���J�X�Yw� �*�Ȱ{����Z5��5B�F�˴ACp�zckq$�Ob|#�u��F�K���'��v����A��(��ш���C�}Ќ�����巹�cį��GX��x�lH�8����2Ij2����UE���Ŝ���\����ޙ�髃�Ό}�����
������ݾIW���,���1�*M��X���c��h%;�B�@�1q���0.�5�2���*##����S	�[���H���S23֛K��t�$�\R��̙ׁ&��ఁ,6�C���o�������H��!Z��`��[�2e&�K��5��v�;�ӗ�]xt�O�����c����m�����!=y|H��[�?�������ޡ,�:
Ž�.�+�Qd�ȟ4�)�n$�ذA���u�{�6��`]^�ʚ�H�E����֘u���9:GQ 'b�����g
����A8u'��o`�"�sgw��E��(*te � �q?Q����8��C�O�����+*ù�35�-�����z2*�3k�����eh'OOM	�qq�������,�3����3��������K�X7߃C���s\��)�R�}�T�`3�C�+�L��@���������6���Ft+J"U�?_&�u�`����k���\&�G`�B�rv�G)�8��?����`���ՀV[k�׶E�8��͜^od5'�!��Z��ӊ��H�Ծ8��6�b� ���+��$eY�;����m�R/�@APL��l��7�ߋ�w��Է�2$���ԶK�5FR�c� �d�_m�:����E4��x�\��Úf�%@Hf� � � �6!R���Ϋ�S9�(� �Hi�W�l�W߈,F*I"oxMa��k�/�&/��=�����@�]�@2�,��JR\���jG�WA�~� � y���:��i��=z����ڦ���żm�[���uxzj���LiB��g��X͛���c���*.zM::8�?���O��8Υ�9Z^����u:���k��@mnmr��
!�|ʉ_�>�w�p�I��LbdJ �%�T��~��٢-o`X�qNx �a?�������~������_�R��F�(��ի��G?�����'����Y6��Y^0�6������?�;wn���!��/��>��C^�h��ű2�9CbG@�9���$�<L�����ӆv=�
��y��OLNhm����{\$�aV4E�����B++��(5�#$ѐW��S�46I�8n�C��q��a-�B��8j��^AvO��%��6B6o�aa.�����@��3]��L��`c�Z�uX4`L��+7j���Z�����cg4�+=���\��4�	���2��H�gɼm	���uZ�8�6��0jow�oE;�3�Ō�Y/ �
5�ˣ�V����X$zx������Zj)��#�%�aSJ�<������fMr#��Mii��T�`�Ҩm��4��x�]�+'�; �nj�� ';8�"OQc��a6�g�J�J{9
�Ѫ�XU��W�]8/ &�#l�<�T�N��Ã=Z[y���e Y#�ɐ6�����;�S�=�r�gl������WU`�Ͱ�C�1M�3]v.���������mn�ӽ�3ޱ��>��;e���??�'~�����\P��ww��Q��S���m���˟�\j��+3��r�֞��bF�n��VWoQ���#��0���w�^��̼w�V�~��:�O�����N����g[���6���cP�5^Y�����B�&*�Ϟ=�{�>�������c<�68� �{��*թ6��M6r��xvE�P��k/>��n��
@��=\;d&1�R�я6v7�K��6��u����� K�b�.d��Q�����$@b�U��R#8�>uUG���.�c�ֹ~'1�źam�u�=�y�$����y} 80� ���״F3��؞{
2(<��]}� >SpH���U�ᅔagr3�(�P�}48v.�?����(2���/�jΚ���~o�kQJ"�c͞���3��^�	+�y�Րw��[�h3�R�9;R=V�d����l�کT����1&�1���e�a�dV�"�@i/��9�_���T�v�^�ؗΜ��_g��#����t���������3r(BF�X�TU�65%kQVp��!�#+�����~�������a�^!@���w������}����g\ܭ���I>�$N�\�5[c|N`��U���f�ƥx^qH�?�����l���MO�Д?֥�ef��!3��"HD���`q ���Ǐ���Ջ�-j�ޅ�7�T0� ����� �L񓣎�����'?�kz�� f����o�@���\�xan��whfz�����t��O���鷿���w6��(hnn�m��W�ҵ�W�ҥUZ\X��~��s���O�=����Z���r"�f��1*����۪m}�:�]?F�&!Ņ>RP��ҭk�t��m�{�gsA��p�E��((�aF�I������PXO�[!A ۖ�Ǖ��eD�e����c!+X0���3+
-�)L�S��,�1$�dlw�(��
� â����ޑ}e�u2c��̨��W�\�����_V��>g�KI��C6m����&�/����o���|5[-	�|�6[o\�oM;��'2��,��ы_lh��L ��t[
_e�(
���1����<T�L��l쌗�>�о��s�n���� ��,5�q/�|�^[sN�\�S�����cfNE�G�rH(,��Yv�J�`�Ñ���XQ�C�).hN��ɢ]��	�L�PH+���2����c�����@��\O��?=�4Jo|M�_G>s]	N�pʤM��v	~����������wޝ�w�Y���^��w,���GϺ��a;��#b���c�낽����?���=���wO�	�zi��<}����IEW�.y�s�
���V~��	Z���y��ӳ����SZ��������`B���֖�۪��af��g�`K--/1+���{��)�m�\YeV�V �� ��ʭz��0g��)��`i
I�=�_�;��Qh����ǹ_���
�������Juf��0�&�"A���a�i�΂� m��L�"x�iW�Vg䧠s�r5�+����.tRNqd�3b\����z{�sh������%s����!���;���7���R.=��9�Ә��d�;�a�<S�5�g���Lpَ1�yWj� ������v���_����l��4o4��*��qH�^�ـU�W���X�5��{ި�/�ϯJFg�* �e����5K�z !���͚
���+d���ʳD�����T�����7���e-j݃ ,�/c�� h5�\~� DX��qpܹ ��3gVh��j�U�]r����$5�%�/Z@7y�����[�����d�ve=�ʴ��e��8��U��F�|>Ȯ���t�<ߦ��}��?�L�~[c-��X(��?�O�{{<�b�DF�:^o������%�H3K��5l0�Y:"s�=�� �����?�����]��ZZZ���.=���?������	}��C��?aI����+�W�����&z��D`GB_z�=zȺ�8�Y��h�����5�(��F`��7X���Mm���Z�_Lόӕk�d����).4��Ӑ��us�^��mai�j֛u2�8���z#��(	�%�-�Y
hU�9K0Ȥ��B�s�m� ���o~��1��|�U"�2-<j}4y]�A��-����vZN�8䵞�f.�G6FmԾ�v��+���?�����*'Ap]'�1����-�b��u�]e-�]_mLӨ}�X��4��%�Ѧ�9�E��)�\�V�9ɠ�]%2�C�	&qBj �Kϱ����w���jZ=ߥ�2�m�O�-���%�+bJ�����;��XLSo�]�,��qS�;bV��9-���}
 �?��R��+�$U4l|f��2K�8�zr�8K�E�Fe��z9�6��V���|dqpȌkI����Su�3.f�L &��6�w���2=����+��w?��I����]Z{�E�}v�����Y� 2�EO�<��<����_X��-��c��8>8<��<<����}�,]�f"���#��O~��	f��=��#��>���N���~2�����9<�碆H���0Yw��Spoݼŷ���c����굫�>~X���^u4x G�L�ڱo�-�7����mmo�0#�!�ݬ��h�38Zp���)Sy��:;�`��F���a�8K��Q��N�su�X۲�N�:��S\��/�t�{'���O��I|I;�a�;Kֱ7��K�}�vO����`fz,�;�{�5M�)���pP��H����v�^�0Uj���@ɹ�9df'$ŝ�8�".|�������F���k��������}��|�͆v���i�BDWV�>k!4��06�w�Xh���r�R��ն�CJa�ѸSRD�㝐�yTt~??���<�y8u����������kdmA&�lC|���W� /�x���c rg5�c�[@]�\��~�e�]|z҉�M���c]E�vjj��`?���g���؈}�ŵDr��"�diO2@�X�L�9�{��b���5iyi�V!Mu����K�;�ڂE�ܯ������VV/3����szr*ͼ�wJ���+l����>cF4�ӿ�w�������O��� ;l�H�{��v�
-���s[���>g[��������?���L)�v��"]�gy"� �Ec�b@���2�� T�զ���E�{m��v�������[��d�=�B��%��+�K��Q`�X3Z�@�ӄY|��V揲��S��#��k@\�:L�����>{�m���?�}jfv��xN�cd9E62�(�k�������f�Vq$��ֶ��l������ڷ�?K� ���hwf��ņk� ����s�T��ۼ�>k��a���6�ߺ�o���H��z�~�FƒH�p��#'��&o��u��L��7{M��؂�6��UtF�*�HV�o	9jo{�b�t tM�<�3�%��V��J�B.9��<���8�q%�]��J���x�r�Z��*��0�vD͑�jc8��DΦMOq���þ�l���6�k/֘1��qZ���m�k���b��n3�I��@����,�����+o�xi�K�s�t�����lz�j����YS�b8�G�Ǵ����\8���`o��V���z�������?��%"��|����3�|����sHb�{�bf�a�⤡P�HptАJ�Iss����JW�^��f֟�ZZ��K���2���:�mږ�Wyt(O"�����N���TU�+�)�W�\����Ӽ����z����'��>W�rzr�YLy`�:f�M�M���t��1w"ܧ�T?(W��Tm�p5C$f&���0�UIJ_0|$;1�% �I�U��Q��Gt�*��-����7��O� �@4$$��g�Y�����>��}��2�zLU�,�g6��2�]
) ��$�r��J�Y�a�BI�88&u�X-^;G}#���,��%�w�wi���!е-�9�ei�}��;_���=g�C�@J�3c�V��� �_ μ �^%/�h�b���_�g^`�Ϲ�?NY)���P �� �{�<&����Z휖W����������� V[�1�Ɲe��i�� FJ_v.����о���J[�%�{�l����
�Y@J~G�A���'gրi�!���.��oPI�-���x�Y.��T]��px�G���힙�)�}������X��%*�������������D���N�Jl� v�n��A������:�Rhw�� d�n޼q�V������Xɰ9�D�c�Uw����+�{�����n�ǽ�b��㗿����#z��z��y@;�����z���ضZXX���K,���Q�?�-}��,񱹵��k;��5�JT`��!x����2��(0�+�\�2��]�7�����z�u%����P�ՎE�@6�Q����������T���L�JA�2�\q�)�Y\kPUC�i8���m��B@���z����Czp�s.���|/�>���!��Uj7Q���rw���̓c�t��sJ�!v*��k/8rxp�A"R8���;�"� �綑hNF����_���I#�R^N�����k�����8���R��%�<O���s��c��0�c9�f�����'`Mm6Z��< *���Z��#��o#`��l�����N0�m�"K�,�
Vi�.�Q?^,Db���/1��ڤ7�tutn4�����j�@_�^�>Y�m\���ʾ'��f��[�a��0.]К7�ʼW��NضV�����O
��)�jh�k)�`���7�����w��8W�y����È��FZi�(R��4fH3|?�դ,E�o�8f�Glo���y'�d{�B �(�&��| �F/^lqU����o���;��ށ(YR�~�9N�G;@�G����J��5�"˽cR	�p�N �(���������|��U��3�����<ݹu��/�!8��3ӜV��X���� ���x��R���;S&�h@�̆B�+��(��{�qQ�3�s���E��R�*	�w��@��>��5w�t|\��lK���)�o�́��㥠H=�����!��׺ ��X��̉�Bm�#p
:��L��Ck*ٍ��cH68תz;YZ6��k
���Ԁe�3(��Z(�����y��q�s��,{��g8x�����~Z��,���+z����:�xJ e���\E"��q�����n&��<�W�{�b2`)�Ǔ>k��rމ��r�QMʉXc՞�h����qF
�@���m.��9rvv��''��|�����+vç��Bo��_O���@]���l��DzM�j�9 �q��=+r1��% �@tE��]9�c^+��i3S��Hp��n����A���=~&�/./�\�A���c-f c?��)�G�1(pU�#0��XO��3��hÁ	ұ~7�;"�" ���^/�(x�Eq�&in����?/q�^h1P�����)��%���������?�bM�JF&d�=}N��n��:��и��Wnҥ�+��4=y��ۋ���'�跿�Ksm�k��s��m;V�Ys�a0�p�eNʊҀa����B�u�nz[�?���v̡�O`��;o���:[T8�D�8�x�<+HV`��c�jP�`	U!�|o�/�5�X�e)�-���F2��pl�y;oks�67��3;�簿�ǌ��]:=����݊֞��ӧ;��|���)��%蔑d��:�KΥ02����~�|s^4�qo�|��3�z�{��XbY�ׂ�66^�B5�'C�F��7�^f����/3V�ʦa��^��ž�P�5�/��6�$�6~�,3��^�e�����Q���X��6��Etx,:o�T)�X9a�,F�#���a��qR$X�������ڨ}5��Ѕ�np`\$N�u�J�
R#]�9%�h!����b\�z�@�d��cހo%��/p}�<�Nb�I�7X�mrն8i���rݧ�L�ru��Ɩ���P�(tBAI�5���eƬ3q\��@�̑���i�n�YpF�'�ǟ�ғ�R�����\��{���O�>Qɒ;�H��TW[l8y�p �ڢ��c��,���<��y�]�r������=c����--/r?��$  � ?����쌤��@s�>?:�J��4�����}k�;��� S���{���y~��~���s<0�dI�j������x�s>;����:.<�_�Q�]~�pҽ�����>l�!�@0��6[W}�<�*���>@��Rh3�^�\2�%r��{%= �Σ���-y}������苷~�+�Gr-�,�}���*�k���k�ebǅV�L2oR,v�� ��mX�2EJ� ��,��PUR�K�MvD����EJMZ��`����{Q�� ��{�G)"�P��ފx��2���������oA�,U�TI&\���d���i7�Z���좴UM�H3]���o��yH�(��ƻl�`}����ux�X �捛����G���G�o�7a���=>:���?F�`�OeP��g̞��s�vS%Z��,p�޶[cT�̅�m0�N��,v��l��3X���ؤ�W�˰�...�5�
5}'����l���8p@� �Ts��&���`&?~��������͛���w�Yuhb���B�1��m������կ裏>��>}B�~}����L&��-� �X_�g)	��x/ŀEcc�{|Bt��->��58.ηP�٭:�N���J���s�7E��i���l�j�L�"ԥJ3V�w�p�:�]���Nhg{�����=�`�.0�Q{ �� ���tͲ�,|��o��$�y�1%A��)����;��.�rKXwq��8%d�p-��� 1p�H޸Ws*���NF��h��������|ݭt-@�6#�]�� km�d��,�x���<����B}ߒEuԾ@�ou;o�
8+iOy����D���U/����;ۺ�{ޖ�*�>r_���F�Z:��f�/�.��Ρ'��>�,��j�֌��:f������)s΀h8�]5�/9��vSS�����i��2��PߵF0�"`d`s��Y�#S�I �<�{`y����Z{���2o|���1�%սc�(��%לU��'��ˡ��ҳ}�s*�O9��\�/�3�z<��[�i~�������{{,M�b}�6�������]�L0��=��bO%;K(�_�����T�X�[��g9�5g�TE'�ǜr����U�'�&��=b,E�@��-�&Z��SYj�)a�TAn�N+��a4����)����{'��˴���dQD}��```�\����ƭ_<J$�#�KUm��G9Xv��d��H�w�U�zY?�3�q��״x���x�.|<x��p������?b	f��Di�}�&��c���6+V��������c�����`F�m����p�y��q��؃���m����I{����a�˨����;.>8��\��]��7i��>����j�yr�C��z�������z��d�39d�JN�.����=^�U?��
�]�޳ '>4]�Jً.�f�ޗ5�'�h"�
���-�s]j��������� ��
���f'KN1K�篱��� ��l�28����VǲB��ـe^��IU���5Y����5��[j��Ȑ%4HA���(*zM��k��)2�~���m���� d�&��\�`5��^!&+Ņ�t�E���S*��H#O�b�2�����1S� �hFP@�x�iyy���s�=��ONM1	 ����h�|�����M�V��2��,$s��xt��ޠ/>�g���������CSj����8���@�<���K�ƀe�����4��R� B�u��5Ѥ+W��u}�ɧ�/��%�����HM_��	ʎ�u��Hw��h�g,3����Ne�0�L\.a#!�wqߐ��"��ǧ,K�mPS��~&y�R�����`�>�d�67���f$h���;wX���p���'{��^)�3�|��^`E�L���krYvDN��/^Nk���N��6j_w�%�Z�Q�Ӫ��k��b��@ ����5[,�+\�O���}�<����tԾ�6���v��U�1Nk��B��{)fH
.e�%��6�A\l��Oc��! ·��A�ВQ��;�o���$��+6��@
��&$@��4�>�Mf�(C�j��UV�t��}�nM���lP3����� Jf�K�c�hO��Y��@� ,� °���:�7!1�]�� ������!�����'��ە��dN(J�+� �� #�@�7n���4e?e%)��<W� �o�S(>�O��tz�J'G`�0{ek�w�ּ��v�v��`�OL���%��O���wV'Y{qrr�;�3̐���8��,���L&8q���j  <>>a��Rl�����l�l�1{�Ԕ�^��(�y�����d�����5~��ez�{�zg�2�;8t`�Y� *��"�hR ��T*����"�Q��$�=l��\�۹P]���2n�m� ��� Ϫگ�����F=
R��	�����Y�Q2�����>��Uk�5�M�-�k�9�g�y <D��X�LJ�'���J�'RM=y���;'��*80Y�XiBpX� ��
�Q]Fc��EɼA}�s��:9ډj��B\���li�g|������/�<��*J���n��R����`A��k�y%o� q ��I`��+ �����	� %���y�5�+�
}t�{Q�خI��7�ي-z<64�k,r��9���ɳE�QA���\~L.�?�/�s�7�	۶`]`8����޽����q��	�H�ʦUr�O�%�q҇�oX`�Z�]T3�Ți�C�$�����X�k���ff�ibr����+�@��M��ZbWK&HV��+֢oi�7�S�cH���$��`l�늍��2���#�|"L��|����������/ X�F���ː{�����i.�w��U ��B�'��t|X1K���^[0~����_���E�Hkw��&��J4��������/��ظ M�~悽�M�~166AKK+�ߏ�����?����֩�|��j}��B����T�� 'E��a%�"��[���������L��h��� �و�L��+ޞ����? ������c�&�fG�#kA�,�є�Zh��b�|<�Mix�uH��Ǜ2�0ɛ�d���a���1g���fov�ތ�s�����$�&sF��(������/��?�EK�"a�K_�x�MG��h#`�;�L����cY%)�5\�>�@�I�,��ڞG�Q{��9R}�Ҥ �r�+�Kz/@D �H�+T����t�=�	J�K8�?�T<ѕ��;��y6��RSB�`5mV3�y�הRf��YrY�����e/��L��k*;:�� U�M��.��?�V�n��m���8
�F���8�e`���$��ߏ�iW5�=�T\��c��+��`��/��W�[���ёw�������C�p܃�����emf��8W���g�h��*�T��
���>�
�H߄N$�.s���Z=Һᘁ�@Z2���2��υ�66���'�z�t�@$�Rp����*
�V7��T����0����b�Θ��Zs�����ɼA�0�����u���j�:�_���ތ��x��>��B���>�c4<N����stjj�!�hR��Yg���Kp$�=��z�o� �)�`leٟ1}��Û��u�3�����;8CU ��X�q^�{u}-�v.�I�1���E6�D�&�k��y7)b�Ut�IO'�G��a�(�y��k �� �*��Թ�5H��@��*)0��R3�A�2��GnX��*Q�+N���S`����d$���SW��#�\0�U�d��ص	@UNe�qM��r�:(������?C����i��hs�5���^��!V.����>�@��"��ިf��{90\���A���G��4�U�̟I�AE6Q�븉�8?d�NLR
kP�o.���^U��D�x)�BNc��_���b�P��5�pM���q^�)��,:%�Y���
����Ӏ�.��[�G� e�O)k��cJ���
�Y�A`�+�,�� [���oS�|�Ș��6���Y��$��ׯs��0�=}�Ei�EI;ۧ,��w��m�}���#�3 `s�/�B{8��i--c���"��(��ꍰfXf�,@��׮q��d=�  �!�� ~KPZX�y.�����o��',7�����⬚(�&�7cp��wi$�{!X�R*������P�`&���&'�m��?w��.��9˓�>���i&��~�Rݞ�f�J�0����#�@��@:�͡��&&�i�\� y�q�Q���9�Ax��^b�l�D�`�f����a��V��u�^;G�m#`�[�j.11�L<��B�-u�����Y����E}/b�+ r�r��h���؜�.p:$Ά4qN �(��6P����)k$��,S���
�C��d 8籰��F�s��c�^��N���,�p���T��#@�	6�`)FA��r�a�W��ȸ0l�t1kiS������T������߇���;8?)����V�'��
������|�悪 (�d��q0���P3?$}�w� ^��9�Q�
���`��O^�x֥�84���<W�?>�F��qfsa�,f@g����#�Hl�M0#�����:T����=a���2�R��ec�1�gH���;G'~���=���#f����t�}�}�&ݺu�fo��Yx'��;a4¹؝�!\��E`I�g�)��N^H�ϕuX��J����Z@z��<���Ϝhǚʰv���Z[-���%���'��e׌�c��F����а<m`�Y˼|���`��b#�D��s��U��B��$���&l��#A� Q�E`�G�6|"�;�f�Ek��d�od�W��*��c־�0�nV% s�O5�d�l��x[j�X��]S"����TG�y?eY~��I�8��4�1�� n[���X�:���l��vAZ'�ұ�k�ͭ�*ks@��������m�#���M�UZ�k���Ⳓv�EMyF9Y���D�̔x{"���SՃ�!-��R��z���k6R5hW�Ь��u(���)�yk�M�\2�l���?����G�l� ��)�Xg��4�� �M!�9!ϙY�,;%� Mxcm�^�e�����q��?�sP,E�zܗ�/+�rP�V(%��R�M���ˊ�Y����c�W�*Du
������l��k�5k�Ap�g �X��x���@2�#�^8:@>9�ӓc-NXJ1���]�TD��"�����y2��' 0H��N���%�㘝���nmn3�z�^'1��x��U���au �5��gh�G�p%J�{���`�JߔL?-<zje�C+r����V���N.�N�jћn�yB�݉�g	jpˀe	�����j^;� k�մ����f'��K'����-Fm�B�1����'��L��j�5P9�ɂ�$�L�\�P�G�:��c~'�X�ֶ:�L�ꐥƢ��[eu�)��z���4�2�qL^���Q�R͉<A���yC�L
�dٸ�'  ��O n��q+�C�`���5��N~��=���-z���������L�+:������['������`8I����7���]�O~[1�� �It;��p�� �r"�U��I/6�43�B��?�J�4���4��H��J���iT�W�lU`gfj�WNR#+u������M���F= ��,���N $"��z�*�X�c��XP�j���w\��;{�q�y�=�j0H��=E�iE�h����s�}����� ,�Z6�����l�������l��3e��i��:\����#Z_?��s����?��wo1�ks�G� �1�rf�0��=r�q�,�R J���
���.��h��$߃�k�&�F�B>h�N=�ִ��������g��ढ�����$-�,ygx��gThq��AZ���$���ls��_m3����QI�\p����T"S���R=n<::>b��s*��L�-cg�f%�h'����-GI.���
`������L}��2�8d`XE�Z@Ԓt���,�"UaN����,îB���A��r���xY{�%
��)�osiܺ��,XV�EA���i:�j�j@����<#ԓ+`�p���,��d n`K_����t�	�@m�$�qVs�Q�#Ҭ�L-�0e��vxn���hr�IS�P笑�R�! ��BF���3%8)9�W��]�J����\�=����*@���;w/����j1PC.���:ra��$��H��oAg�ןG`1[�?")8i��gLY3V5tu�F�&Ƨ�]{�A�'=�'����6mn�Ӂ���'[<�>��Ò=�SPr@��2gU:��x�m����i��~��0a��:f�G*G�S�����=���v&KPAa ��rn����J�q�ׂ�^����fF�]�W�2{�������,�Z��6?�w��e�|�
��^��s�O��\�����E�Ӡ��f}A���3�5g�!_Р����1 � ��(�#,6o=��j�U���O���g�l>�dHUIڠͣYx��=��2=��PX5��7)�s�H�ى~�Pw6�Q�c���F�;�\�� $��oj�6�`F���!H��w��"�� *&���1m,ך��ɐNO�t-�zޥ��D]���W�vn�����t�&
,+�*P
��;=��>0�8���ta8R���D.`��{�z'y��%�^����ش2����������%�D�����O�-��,5c��z�uu��a�����٬�y�{�%
��K`^������wb�����kf�h����L_��Ĳ"��I�HGQ�#�JM�� �ﳖb�RR9���۞�lH�.;�Ʋ+��P>���7����±-�a�$�;0_Xk;�m��t8�ϑ��,t��  �q��9��5x��� 0C~��!��ܤ_������ϕ�ޘ�H�&�ˑ�XX�.��A�T�,cy�,i�.P'7��
��Χ R��β-(�����2#`}���[�\�	�2 �w������{��p��D��s���o�!�x�N��ǔ�^�6q�2����^AQV a,'͜�["y��,�Ա Rm
������c��53C�(I1�g�٧�B��6i�!�a^ ,h�)����N���eat�)�K�lN�N4�ө��mL�΄ə�{��+��0�-u�*;'���jЯ]c� ����`8'��L��'�$#�p���i�G��}-����8l�!�3^�;V&b<cY#��FU�Ѕ��9����#���i�� ���9^�1眲�lƅ0� �(�Þ��i^݇>��	��6�\F���C˼q���'R!�#31��Z&q�� D�i�H�D[���-�U��\U��WDva ��%��ՖVslg�x�6_lp��د��sS�v�#w:'�f"c��T�Lm1U�)��?��,# �e�Me�:^C 8O�{4 �߶Vc�(�Z�t�וuqh��y�-�̞�J�JZ��m��L�i��j0�e|�,%��E�A4h5�z�R��m�k׮�u����L�~;��2��BP9���b�����YJ�@&� Hd�l����&K�ؼ(�d�c��Ko'���[쾊�]J�p��e�5���eM@f
.��w�|�Q�"ͺL��t:/��"�612Sɠ|ɳ�=���w�����DKW,3��Qs]�F<��X)3�˃�
RӨ�������v��RU��~#a.T❷Eg�Y�
8���9�D ����ѩw�\����O�]�s�)�Y�"<�*�!`���k��Ή��$�Z�n(C���{�H����z�em���
GG�I�42 C3"rz�1�}��������)e�(�`��U�ΕR��h%���E;��v�Qa���2GpKqBE � S�!��=g�6��gO�Yl�Λ��F(�a���*}��:�(��Zb�T)��y7I�'�O`��X��
����?`���Xp ;'G��Ϸ6�������=4N�,b���Z���
�����G�gLU��/T�����qT/�*ϰb�G}NO����@ ߣ)=k������Z֒��a��`Cw��r���gI��������K抁o���F%eD�a�	3��5�$��Z�
� �ѩ&���i�p��Tb�]�^E��;�T���s�J8��3��-�
:`y��N���[�j�k XN�ci)ܓ�;d�Q����n�ڗ�>#HM�q�6�O���
���j`�}��Â	v'\�{�Y0j,�����<�7|��A�۫d�� W��p�A���èSp�},Q.���ي'�y�7C?���?�0�^�u�o��D��	�F.���V(9��̛,���%���6���cڂ!��xU.\^mLU�>��}�������}I��<�bi��$�c@�R�Gnnn��IPabr��������٪R�*S��R��(�lZ�BTtu��":g��0|�U�CH�@�L姒 nO�?�IۜJ9�k1������R�Rp=f�Z�V��u���xnR�"�u�sؑ"}�&M�O��3EK�Kt�����vÚ��/d�9��,�"��aH��좋�eN@�}8�
OE�DJFW���X�L�d��~H�N�e�2-e��]rm��5Z2o�Z�ԩ��u'G���<j��\���a�}$��|X�,�L�d��cD�A+t�FM�X�N�t��h�:Ox�!��P�Ʋ�rZ �U�9dԾ�-YG�p!"�Ƅ��a�ú��c`��aV	X4��G��<� ���)����6��?�{�=�/6X+M
\k�J"A���{Hϟ���� e!E����	ڹ��w渖�v�S�3�q��V�:���6�sNq����t������?���������}w����><���B��X1� �k)0l��:.���(� ,N[tr����AJb�NNO8��7
����M�|���GG �f. W��m�`f��*+�g�ٙS�h�����Z��*s�%�PV��t����vh�c�|�}��3ҁwvv��OK��h윬���'̐?99��{"O� |ll���� �ϝp�|��$�37 P�^�wK��\��4��I%�sƞ4��Ǌ4�LmgbY"f����@qCq��_Y�h��_x<<+_�<y�����H��8M?��e
{W�Ȯ�z�eݤ�D�ݘ����2wM2��]�3�}��m��Sй��H���R$3�Ș	-�2�����ԑ���>˫�SZ�C�w/�@�ȶu�>ם�����)>O����L�b�EV_��5$h=�;U���3
-ܗyR��4(x���|/�����먪p}�«�iD���l�9]�r��1�Ӂ�[~���S?W��4@�գ����Iw���9�~�� O�u¸�
k���wL+v=X�(
wppD��Ag����YgjkP� Jƭ�=��ac$�"He4��_֘m_���5_F�����#giuu�>t���H�?|���liq��gS[����,g��4�,�v+�&l`H[@���h�dL����Lo�Θ��*��[��Ԯͤ�2'P(ʋ�V���R��JǱq�dK^������&�&s1a�v���m�㴴�L�+����ޥ�W�Ѹ����Հ�>gS�J�fkN&�J������zX�"�_��ܙ�*�U`i�^��^��MV:��g��t���QfW��_�r�t�_~��ԧd|��nC���6j_cK�n����2t�$P�?/���ĶrJVѭ�nS=�d�4jߑ6���M')r��݂�/WID�0B�P���_;����nz�n4A��7�X�׽���t��x ��̔���e�={��O���IK+cމ)y������>���x�����m����^��[�0��LYM"�z0a�PS�@����+$(P4�bM�So�1�(F�S��9�/�,��B��tx�r��B���ܼ?��c B����֞�����>]�q�&'���pO���w4�3I/'���^�<d��J����O�ޟT�WR#I��i%�F��j8ǃ�=��h�&B�~zg��;^���
��L41��tt|HG�G"��$8�g��^�(�-�j��avyΕ��{��=���b�O����m�}�����+3�W?�#��U+�+���m�p8 �����fd��d�E�S�-�&ET{�l��5v�f���܂A�.ߧ6��0b�`~��|��yָ���7�.�K�~ff��ܹ�)�c��� �A��J.����q
��,�Q}2s.RI��0@8�$L6>����B�}��'�3�50�N��`�A44-�?@���EXNX��`��aE*k�r �&0}�6�>]��~3�zŃ���G`G�_��_�/^^X���d�K���� ��w.���>�7�yW
�
f�} �R�M�r�5�ɹ/��`�Е#�ד,�+kD:���`��@�zQ����~���(�LU��|gR.X��M�y���w�ҥK���K�=���?d�/2��MaHo��P�S�Y`�j��sNCZ-��6k13����~ܯ��>S���tN��_<�����V�SIv������/�.����l��	I���9�5�v��q��,-/��t�nߺE7nܠ��9��L*�ׁ��sb����W�͢V�T�,Ǳ�r���()�s0�Ml:G�\u�/�9E0���G�:�q��ٔyq��\�z���Q{�gqe���h��6I���iJ�c'�c�Qi�3��6�����#��F�"ja�JM�2:�!�!�n�ˋ����+��Fm�^K�3�i�w�N*�R%��$��'ިg� �"�LI'����0c�=�ꝁ&�z��s�����W�av� n��f�d��lE����)�(e�P�_DǦ�E8s������2��-��8��^�c4Dr�ApH>t;4=5��Y b�}+�S��_�gkc�hMNNK愛�nw���64�[`
�p�H{���p��(�H<2�`���,�t	h��8k fY��Y/�2pX��(�Ț��;h-�7U���c�e�c�ө�+Z�y`��yN������f�	������]օl��03;K+++�zi�g8���m���J�
��-��;�Yx?F%�e�Ϯqi�`���)2�C����[ګ�a�u��"JyC��(��<�U� �����֎m���\="(9y�?r
<���FG0�ep���l7I�"�a�':��������e��g)��]M/f��N0)Y��ϛN��OR��{�����6q}���b�l����������p8��O�b���
 v�B\:�=�����W�BEo�F�Fn5�Y��T�،�a�7*���,n־�l�8�T ?Bc��Uf����+yͲ*���Ӑ`����f�z�/S�,�r�u�e]�Jۉ}�e������� b���82�����t��*�ȴv�;����k�_#/q������lӱ���>B���b�\���XCع%���Z+���N�����ZX�$��P�}ρ]-l�3K[!�Ā|�}v�*�n65���5g봼��:��%�N�|2�` @���Ņz�����k����coEyBvW�u�ι.y��<��	)K�w}D�>b��<d��VV��,7H��t�U0$j�j���>��ٕ�����ّH��N��/�����.��ƴ`���/7dS�0��-u����Q&�ĥ�rPgX�u�Q���l�D"F[��ȱ[�x��1�,����ES�����/�6�ڨ}��lq� ��f�Ac�V�f����Alԃ�g���פ^��m��z%��s~O�5�MNW�Û7ڪ��\ӏ�ae��w��g����[\ .���r�I�6p���3my��Y�ƪ鬺Z�|�3I�g6���:IIn�b	�YEǄ�u�u*;%}�h��צ�]^Y���y~`�S>�Z1 �e��E�by����`�^u&�RXD��`���M1&i��?�凬Yܥ��-xgl���=z��9����B?��	Re1߁m�1�r�Ck)����d��& �q��.2����>K]��ܢc�_�'�+
1��wߣE�PfGK�ቩ)��4TW��S�fZsĆ���.Jp$c�n6;��HT xXJ{���l�R�p�n����y�_0�ڿƤ��*g��P���萼>/�R-:�gY��Qm-��%�=�ag� �\� ��,Ϫ^�"ǵ���i���Y���Z��$g��k��ķ��>��L�7�)�9޳�����z���������m����{?����W�����E��A5���Fp�߫�_��W��z0
��!b�eF w>�Nj&DĪ�1_R]&DZ�o�z��Y!��絰N�z�2�+T���e�7��W�7��|�L��E�(��ߤ3�ζ ̴�˽g�H�É������lc�f��n��U�sJ��ź�����^��Hm��t��gy&;9>A ����i^�z�n�~�vw�8����g���3�!	{��5ia^�"�����{��Z(EuM߽�9ef3-�/��XJ�[2�p��pԚ�g�l��,Alo�Aϙ����{V�ve��F��S�`�s�]:�=d�L��3 _�q�n�K�f`oc]�TW���oǓxUYQ��!2?�Olέ=����Z_�1TqnK~d����x/c6�3��d71����ں3p���.>3�x[1���#K�D[��y�i�R{�?=j������ӷ�9�tZ�yx��8��T�nFm�^�F��w��VMPUݢ���~��������h"�7�%����`P�477ïa��"7�wO��� �9��ީVc/i~^��N��OBw���B"�J�8v$��G��d��y�0F�W
�D08~7ȑa����������*�Elj{�NA�,����D�q�
HH���mmm��ᡲ�en�����<���A@����o2+W�
Mu��2q��Sg̊����r�?�nO�M����: `�Y��c�s�D_�0����o�{�i���$�UD1>0�������S) �KK�4;7�����d)����ܺGzV��*t'��z�� 
Ҟ��J*ʞ\�v�-)������QG��*��ȕ$�cJn�u�~e��9�s����+��o����c`� @i"�|�\��M�w:����tu�E/)�mJ~�j�Ym��9o#�T�� '���e�|���9}�F#�XP��]%�j��I�I��VQ߮��c���n����ه`ư����:T���u�f�$�$��}��Bح��D���Pג�/@5l<�3��[�:{���i.yޡ��y�u6<k�yð������I�Օ��k}��Mߘw��{�#n����s�o����:Ⓘm�R\����zY�:�XC��v�*����igg��YWr�c055��9�:������'��� .��h3�p<c���Υ�4r�'(��P�Ҁ{L+E2�Ԭ�Ԗ��Z��Vã�?S�ArΖj�8�>77G33Ӭ���N�3s4;;�6g_�LG\S)�_N�q:��2����M~��gjρtb��Чm�@,"y{#c�D��Ƭ~�u�ɱTc��a���ZE�+�>�l^O���aU�ː���o�<k�\�%�b{�oFmԨ⌖��a��=j�6����Q�ǌ�\��ԣ`�H_����ф6j�|KA.3��pøG&���]����t�q9 %efU��x��c�w���j��z�����3.  "ugf|�Y�x� �#�CM'����{�d޽`l^r���q�T����Nȸ$��/|����P(e�ދɸ�ű�h�S�VǬhk��V��������l�(d�l�BN������w
�}�PQ�$�_�|A"��!��/�����?~�6w��B�+ �WL: i�ގ�l���C�D��$0�4�!�H��ק�>#����� �>�F��5l)����Y��9�u�JP|��d2���l�$��C����/���'T�['�J$�n��b���-q1��AZ���F��e_�&!wzJb�&ďzf�&��痟Ɏ�KNˣ���Ƞ�«���s�����5`���$l:���"dqH��D�6E��c�hcr9��?!�5�,c�R2F���"�>�8�F}M�\�(�_X�M��j����G-.8v��w~�,������83yfn[u�R���h��8�G��/��z���f�H��1�s��Yޔ��.-���ve+X���A�k��F�}��ߗ�]B^x>!�Б~!��v���b���[n��kQ�b�6-X��� ��+�o�@���ݜ�����Q8������������s������OA�)(�|OE^F����DF�U*��F2*X��ƹHb�8�؈O4���*� ��A2�a�ǁ �t� $�)L4�&$~z~��(a��wu����ܯ����������������--܃��(�@*p��񼈤�E�I�A���������9i�YedwA���/������9d��D9����bd���qO�H�9�닾�GJ�fQ'��K�LU\u�Nmr��7�LA/�M6�%r���ZPI��ڇ�:0b��ȃ
o�n��뎗��hy�CR蜼����k2`�`0���V��5͚]ȷ���Hhi���bEaF˗��m6��[�!�]�{��Xn�24+��� �&~���d�vF������>+�rA,"}&��=벴0-�OZ�*������	�s��w]�>����
� ��ۗ������3*a`aV�@��{���m �q7`�ܖ������s��K�ҺݱώB��8, ��,��壵RW.(l?���l��X��[��S��*����7������ ���������r���ʀ��U��o��b3t�����Mi�%�qtz��8w��{\p�][$�TR�̇����N1���\��6N�U��y�=���E���$G��2�mKҴ���ǠǁS��V�����*1NYyquJ�+*�"r�,Km�0�"�|�+	�TϚh��{��'�~�1n�?�����T2��gR�&�}�r'+>r������SQj-!r�2��T-����.�vv�2\3���b�/G�E�����I��6�������|`�8{<�� _Y�y<��� y��Qc������i���"�Q�ÊqO����p7�l��]�����6��}���o����׿���׿���������'&������[7O�����?@b�{'��`�|��)���d���'����V��䬴w�D<�'��h�(kue~��@	 ��r�U@4�f�&O���E9����p\�Ï�?��]�����a@&���z}��~{|�Χx������?�V���r�t%���W���p����}yޕc���_]ʘ��i�hS�
��<fpN'�4�@bE-I�s�k�k�*��0����e�Au�G$�ߥT�Ҽ)�qLsw�]���r_�7�C�lPȃ�XeVN,)���&�#�����#���1C:��p-�A��@Ē&��
I�q5GZH�I�B�A��&Z�)V�[�W�I?��:��WJN�iN�%P �2xf
��b"�$�J�(��B[>����;�e|�ӭ�y`�B?<Q�A)�`P��99�D����U@\�c<7*,H�9d*ʢ�rH���B�v�n���t�� �F�!��SJ1�Z(S���N�5SlG8�kW���'$��]}��[�����<~���d˧�:�履q��)�����f������C���#�.��MR�g#��dz�f�[enRْh�N'3D��*�,NŲ��J�,9W���:j�^)��"�����pp]���z%����W����!
m&�5�D�Y����5�H\e��\"�R}��.������T���gE\�<�h�H������A*ƫ�VO8������[x�4�}��Ψ�_�+����	9�*1���S!sT[��!�p8�q(#z�;'��!2�,"�y<R�w"G]n����5�?`~xi�3Y����}r��y\we���Y�Ӽ��XA��<&IYI~�m*y!���_^W��r�}�kCĲ���Nd���Wj�j�)=qG�S��!�p ��������^��Ϩϟ>����?��ׯ�c�	�q'�B��(b���̇�{�.j)n2$���m�b"̐���=~����?�²#�����oW������(#|�dXH�0Y�������p_�1��(G��.��H�llQ�ri;�&}�] ��B���F��^��w��S9wd8Vxu&�Y���b1{�=��S�$�VN<ܔu�"]h�ĥ<.����Sc�М��R��g�4����7����ˆQ�!X�)A�9�^ݬ(Ҷ�ۉb"G3�v0l�5\5u���(A��-Y�� ��*'�ӕD֑��Wsl8Y��Y��ٲ�pSw9�Z&+	8��"c��iPV�A�OAH���$�z6������窌�`�u{zy�=�b~h>���v���'����w"z;�J�A��!I��@�~����}D��G�����p�ށeOKJ�YM�?�����WL�d������?>�����6�ާ|�X�`5d��?����)�`]��?~���������ҕ	�[�%B d�����cH�ZiV�=�^fwu^��zW(jԶ����g$m��i1�c"	�/*0�
�x���^)�j�Hs��u�
zn-�>OOL,ɽ�\EʢPK���ZQ��XRn��c�*���M,�D��>��:&bYBo���&��7�
�0"��"�s��dc���Xe�V��6K[�Pz�?/���=&��-�Л}��4�+�r�%��-�ݶ�,�
�"�u���W�����o�����/A�MxI	V�6}�E���1�����be^�Q妅�tP��>O�(k��^�G�f~�zj���z��Z�+Y�$�H��]�>\;�~��\�����=~��?����!��ӣ{٢��h��B���������x݆O�~��y����Er�G0D��}�� �~!��O�:����i�	���l���������?��;���_~�X�z��50��Ӌ{~zAO����=%V���D�S�@���~��w�[=��Q�{ӭ�XtP�M��!�urdk�rQ)*�Ll�!trLq�X�e	�\FK��p��Jl�,�Rx��k��C���^@/�K�g��X-������'���e� ��J_[/�pJ���rY\U��!��c�5��Jõ �M,�(��$&l�9ٙdWG��QH��%b������	�R�� �j�Uvq�9�~oB���S��+��I��H�[����L�.
{��h�S�R}���r�u����+�d)�_�*ٹ��kCϸS�=>b�o����gQ�~w���{�E�<z~��q7���cp_��\*w���bH�����}w�o����?���_@v�q  ��Ͽ��n�`��>��hE��Iyz�p��#� J�\JV&
��E��=�jJ��h��t�%��D�qޥv�Ib�c�A��-�ˎ�I�7�\Hu�d=�:I��ظ�ˋq��xe^�\�]">���ET�#+��Hf'�pY��D���\NI�R�T�����6�DZ�{�����rh�y,8�N)�����'�aTT(	�Y�"�3����	��v�ڏ�3�D�;�����Y��,��V�s�וsNS-Dx����i��X��MsA�Ċ��^�>K%A ֤��R����MH�e�"�0Yoòܯ$��|(�_��0$�z՟ҿ�͉�h��������bUS��r����}��8��Y&�����4h!��q����������g�d���+���ƿa�<X������b-�������X��}��;z]�ɁæS�W����?����O�&���f}��wH*x�؝�e5b.s���C�d�s�n�&�b[�2�ID�g���z�a��;/���p�1�8����~C��ڿ��a5�PԐ,��|��S�	�c�<W!����Z�Ur	���O�c��3&a~yI!���1��M�(�wk���`Ĳayp��<p
�@���U�4�K�(VLCū���ŖvW�4�J���JZl��xZIW<8�/�z3~��"a�?c�21��$��Y�Q�d�ޠ�oyU�BV�ˠKl�/���������Τ������^)�d��C�8'D�(����ڬ��x/�upV)�ݎ��a���o:e�	��K�J X	y�1��et�I�(�l��<�!�ѽ?��"���A���Ǖ�嗟�*�G�����G�~^�6hy-e�8;��+��H�EM"�==P�2:� l�yG,1�G$�@X�#)�I�'b42ᑲË^X)��>�&eN\��
֧��/�j�n��U���O�J"{6/���(י��%	WP�?q�e�Ǘ�:����Jg﷗t~:�����N��G�Q��^_���o.Gջ���)�j����'�>�Öu�W%�)Y��_�S��2Zn�t璵5-��`\�A,�]1.�,��-ӳU�jߚ8uѕ}����Gr��萜�9��,؉�R1�le��U�K]'����\��m ����cDq/.�����ۻ�b�@�����/�¸�tr���jwOH�g�v��~~�	�!L�_b�F����r��00�E�����G���X���Cb2p���֜���D��eLJ��C�k�B$�v.��c+f��ߍW���Wb<ۧ1/�ۥ
�#�HrN�R���8�Oד���ʣA'
���-��k��,VB�DY����bc��i(��� yD��ˍ��p�l�V��X9��#̾����ܩuY��I����׀(��/j[�-֦@���#�ƷBs��D-�ш�&e�Ln���,%�Jn��C��)�~�[}���¸J,�z���PHdTڑ����v��\G�>;kuIU�o��?�8މAn�������(���--We\��ϟ~�P������C0�z�@��H����Z�Sb�[1��ww��e����#YA!�ㄌ�����24��/��#�|"ː�	Y�)����������t���0P-N������^){��11����+J,̠�a���r���DuȌc�B���HQN�c�G�-�)D�K��/�@Q$�D,+;Eս+B�"ۄ���~�� �+Z�%�=�q�u�?z|��s��k��ќ���X�Θqъ-�c��97��dE�%��c`^͹�o������X
��� b�(l~7,���{��b���o��<�H����՞F��Izٯ��#��R��m4�3B,�rp1o(M��X&�P�te�s6�v/���[���i�`�c'[���O���[Myz��z�-�����Ǣ{y�ah.��9�s��ju�bH ��<�	���;ɭ�]ӔW-��p_����詊��\��_��^X��^��</0��F$�"��}�LMD:�(�������})���&��u���ԐdÊ�V(�Ř��t����_�p6oF,���Fu�D��P�0�P˴4mF���K)%�b��i��)�������S����IM$N,ƀ�]�U�_� Q�#���,� n܎��V���oh�ꂅ�d����%Ϊ�Bt*�"���B<+��-+�'%���Y��|@:�Nm������F�B@$B}���'J0X� �,�f�mBP�����OϠ04�������[p9NlD�B�EYM���#	M[|�;��0�R��X%��I!�E)�K9y��-�-�~fb�ˢ"�T�#NJ�$b����x{J��I��	��d�+��>� �,l�ċ$��Q����U>?�޵ee��"!u��X	{#!p|�R9�H��wm�&cB���������P�˪�t������0U��Q�����#6��c����?"��Y��k˸�H��B���&��@�`X!$����t<~7n.�"Ϋ��4�fP���[��V�/�g�AjL�\H�/;��q߱��:�ܘ�D�L,nz?�;@O�7Z^� Y`����,X=�@�[�)�o����D�s��g����e�]7����Ky2<x��5���wZNt	Q(D�EEه�QL��d��+�a^_�#��Pz�k��Ҿ��C;InK�M��� �c.�(����Ltx���`CtР�;^_yPy~)�#�d��mp��D0WO�=,bn	�e1�ڞ�0bٰ�����&y�L��=�tK.�8�1q��)M��0EB���Z�U`+�Qi��@��P���^��{L����m����.���	a��L�)n��d2���(��dq�DQC���l��s�W�N����&�-K�+������,8����1;��Tה$/��m��aM��a!�T�<s����VĤ�8T|�KRy�I	���U�ړ7��f�vA�2ޕ�m��Ҟ��uj�8?ײ~�%Y��Hm+-�?�¼�^����BrpLLKh%w�����O�a����4-,�U�'b�Q�sn��
c�7�����T>�S���u�fg�)�}�ʫ/�,ґD���s1��'�[6@�
+��X ��i�ɂ�XF5�F'!�$4���@���l7�b{αs{!/x>�}�e�)����{+����q�g8v{�5�}[�{
��ʅ&.�ł�)�.�ʜP�Q>�ef?Q�l�sMoׁo.{���4�u�n�l�lMK���3��kq}����=�`��d�d9h��!H�UP�}���K$���4wPh�:Y���x,��A�_C��a�?�-Fzm�YO��t�^�����UƸ�CǍ���3�s��l��m�͞@zųh�]a�Z�	�v�,$w���&�	�;����ˆ�����+�*��7�A	b�����h�"����&�� b���Z���)���P
��B0���E�E	�����r.%����G�*���	l��(qk�B�d�!�h.��[O9����J��#�fM���@���k8��|,�U�Y����� �Y��R7M����3���~&3�})|Uf~������|���]�8���>2�Ǟ]�A���?��N%(J��T�.�G�'O�� ��o�T���ؑ���G��6�r�*ڷ��F"����d��1\�թ&�y�&K���tD�h�^P��@�R"�\#�Z�D_������=d+�V�� �e�H"k}[H2�.
I�Or�,$������!�+{�vuZ���]�7���%ܘ�����G���֛
�#VA���0�p�VsH��\��0���+�Ю!�D���P�l�^(k�9q�~G���ip(�I^��x���Nb���+_X ��Og��av0lF��ez�r\�����0ϙ� �r���@5j�o0� F,�k�M~3�m���}�/Q�a�$��j
k@QC�ן��X0�w���P���z��L S�Cb2fa9['7N�X�d)Bq�(C�J���c�,O���-���Zu|e��0:��CKm�%�)��
\'��7E�y�鲒�,H�TIZQ������W�շd�V]e��(����F�dٝ���cJ�b@)������A�j��4z���Q?�j��w�$��c�-�՚�vi%�%~�LP � ���o�ܟ�SC��t�Z�֋P���glx����11����´���J���ar�I���!�#���ר��Kb@�G�$
��sV�\��i9���P1�/����>����m]����-�Z�H�*y��i�wh����SZQ�e\p:�g>R��L�a�
b�����l�\Z��C_�Mߦ�R�ļ�=�6�#��q�6����B�&F'� 2�ľ�ۗ`r��(�Qm�,����c�P�q��h]�X;Z�z8�-j�~���P�$q^_?����RS$k����M�~6�29���P[��c2c;�
�R���,��b�r�*%`w�j�oaк���ȈW��y~>���b���˜㱽�vk����S$ϒs���r���%�lm�O�RM�JG�:Y�����1��!���2��#7�L��P*�Qd� 	��Rw<t�s��E6L�d�,1)YYfH%E/$�V�9�"	�Mh��Xj�"#&2(Y
��D]�\�̕c�]
�yG&v�
KZР(�Ȃ��WJk8]�����.��~|�ӠѴ���~.��8*N���;�O�c&򓛾����{g�3J�c��.Ǌ}�z$�Z�:dr.*E�1Y�)qs����{+�ҝQ?��/$~'�\
�ላF�(H��BZX"�B��M���띕��r���2Y�G�E&�~�yT=B�VtN _�%ոT'��{��d����Q���5e��`���<އbAgnԲY�9}����@�8�r��T�i�Z�$�3�F}K�-����K��d�����J�֫u�O��ƞA=D}������ɒs����������my�!QB:�ˬ�OH����1蔯l�,Ii�ؔ,�cL�CZ|R�&��4��"�ȃ�9�V̾?6��2��I��D`��uR+='�+��>4�S�e�<�P{�X{���a�X6�4�i�j(�6�/&R$F�a&��^�n����̓��wH �'��I�S���E/1��	�Z���!��ĵ��l�(��>	�:�*�A�l�r�e�v�,�ry��_X�F���,�#�e ���-�r���λ��g��ݺ��G�z�l6��æ�{*z�3��?`�Ae��1��:n���^��?U[�r��/���"�~�L���	$}�d3�t,��@,�Ǐ@��J�kq��c�E�Y�H���|�,n������S��;���,w��D�Z�#���],[h?)��1�X�F�Y^�)bY�� 5y3(��blBY���J�ʆQ%M����0�����9�P�т5΅k!Qո�+p��$�L��ϿP��w��~E��1��1�<e��G�n"F,��2�E��$���_�b�Y�/�F�>RT^����ʪ:�Ǡ�7r�`0��X6�4R|H��E���'�.IyY$0N�p<d��rW�#������)�v"�X��l�-|���_���ʨ�|��-Ĳ�i�%}&�E�)���n��F�J0N�r�/��5ќ���sYDw���'�c,�~���S_�[T.��NvnYw�Z\�T���G��\��5P��q�sb-z`~l[_I���Heٴ�pU�Q1�b��B��;��mIa")������4j��Qoc�U���}���XW�U1������L	���]sq��c��W�.�g.[��|u��z���\O_m��/u��p�tm@�l���I�8�}
�]��D+�A!q�c-�:�ƈ��:t��bɈ���	��R�EU�9��V��W�K���� 9V+���Szl.����p��������2��NT﹖�sqb��u\�X�ݺ.���NǤ�&���/�<������Ob9g�T�:����߆w��.շre�$��n�~��Q��`8F,n�P�BU��HK�g�4��ѣ����!���V�)5����r�"�a�LՒl+[)��rI,g�H[%	��?A�����DA�5sHA���8yn�.�H�I����9����G+r~�q�����2{�Q�hAn�i�s�=�H����=�Ȗ�Ҥ?4.�~�c��NWQ�L��qI)��r5��R�)f, Y]����l�r_�^����=�����U�q�q))5q��1+�S�Cu��(ʹ)\�>���(����ty<Nd85ҹ뾃1�#%���(,RLc��D�;�$���t�����<֛���1����h���ҭ��a�r�E��pr��
��� [�^8X(�8Pgu\�~���.�6��6��,a.�+������+\������%?�^@.e�M#�Bi�7.���Y&n$�D+�+��7f26�U{h�;}�is�L��>H�. �!IWS%�R$SA2�U�X�J�N��^��1�R7M|��Ou}}GC�a?>�����#�����;���B2���pW&�����X�U�ԘE@XO����{$�d��Y@�)Eb%yW\W�ZJ9lꅏW
ID�OM&��Å#��"K�U��Y½8�/%,L����娉�>�L�Vн]Ga)�<�c��9W���
���$��ȋ1TGL�{���K�@��nw�]L������I>w+�uZ�w��ܬV8V����j�ȱ���;��|�:���e�9�P7�4ȫ[,���"r�f~F}������r�Tt_���3%�{7����A{��D�G�C���o?�Xc0�F,���S��l¥ز#�_�1�{��+���(���7��O�I<�̘�䞞-�$��6B��ƌ���@�D�&����jE�%�>���lM�g��\���u���j/4F������<��wmA�)�,����o�ħ�?��d�& ���B6	�Y�ʲ8Q�}��F]~i'��<�">& AP/�Z�]��w"�c�]�4�J�+ĕkV���p9N~/�B7���Jm�&Ž/�_���5�u��!��1ʻ�^ף�8K�t�>���#2bu_Еv�-�r�D��4X�?����T�x<��[�w;�`����	����p�Sc�P-�s�;�]u�����2�K;3���ng�绔�0H,O�uIL,�(��yz޺�nG��[�C�aba�?*#��'�+��>5��U#��ÉaĲa��"m>��B�b���|C���çy��嗇$c@,�lI/q��4[6]�k�d��v�b9�+ !��j�!/ N�"�����#E��O������@SzL�о,7���(�%�֫���cIJ�����V�p=
�X�����0�������~����]�x���1�z*��lm+E�]����Kl�OVb�;��NJ���N/�S�v������yM_Jr��p5�U.�������s���"H(�k��0DE��,�+���^����~{.��P�����_�/x��˳�n�#y��ᥲ����W$�c�2(yu��asV�M
���]�M<�y��a�e:v�%p�k_���{сXf�9�Ĉ����W��	`��n�ݖ�8L]�R��s=��߇)��W~IM!q�d0,�ˆ�&2
R��~JC<�5(4�A��B<'��y�jCE��D�v��n��B���j�hmԬ�RY�d�S�w��2�H�rEʥ��1C��ʇ�&��lSz^xJ�4�3Y�}�a�l�>ӂ�����s\�jkRԆ�����R+n���|�j�r��@J_�>���� ���CB�Т�ڂ����^o�i*�W�NM	<Wy<�?����-d�Ō�k���R�E�r�4���\�B��#�f������;�	��?�yܠwK�y�����?�j�W4�&��/$��X���0�þ��_����[F��y�LԲp���[��7���6�n�g�W���l�qb����m_v$���J��WC��9�� e�O���1幀�cϴ�uq\�b6��hv'�5��b��q�i��X6�4��i�V|������������8ib��b@���/�!�ւ��J�\цE�G~�mS�
0%�Rb���-��`��͢k$27$�zz"!0�~r*�5c?��೙8&�vug�_.�z��M��R�{����9��@T���N�̕�kE>�X)[1eA� �G	E�{�����D��wQ�����/��R-7�LĢ�'���tw�}�yꇲ�*����O���2Ļ�Or�!���c"Sm䤚�W�ӊ�޾p5�+�k&�C�cJk�c�id�)?c���DiI��j���`]9;"��Q��I�LG�Y�"�z�'��X֋+�Py������:�R���֭>�a�O1����h��q�R��ԯ���1�H���LT�	I�(/L26z�o�ş����/��+vĢm�:��s��p
�l�iH�I��j�.��c��5b�pdNO�Bb�Ea�>[�0D�53X6�6�;�I!��2�ö�
��4l�ܤ0:9_YS�*�i��A�j%���t���j�$�nY8��{�����+���Y���g��ßK"�������k�$�}q��\.�1��U����5_/_k� ����9������:F��MHBmb���k����m6k&�x�H�i`�8� J@������P���I!��R]j�&�-�G��qd��U%=n�q��D�c��MdKe��@"����W}f�� D5���8�	�٣lyN������GNe�ɑp�������o�8|C^��N��x�[Lݦ��i�U5å���؍x��#��&�c�|D�TS�Y�l0�
zZ�7.��	�����h@[Ee�-}޼��!d/�dE
�@>��N��P*Y�|�׫��J*�rwI���
����R�j7���'�Yw�����{*y_>3.eh2v<y�1d�.��H�9B2�븱C�6���:M"��GL���`.V��G�ɖz(��� ���8iլ0����[�W�b�^��;l��/��i�h���J}ϲ�<8��h�`�؛Q�o�������W5���Z�m���+IBz��à_/xf!5 νdQ���;5t^�ɽ�E?ëƒf�I���9���`�w�^^����Ӽ"��s~��~��$�X�}������6��7%2��ˆD_,G���:YX��b����*�'b1dkc�����
A��-�a�X�]���!'�K!0B&��RzX �c9�3�8+��|o#1[e��^EF'��vd�,�|]�FI�δ�,���5�+���΅E��YI3�p�ȱ{븯�"����[^\T�r:��osn�ʼ��z�r�N�����7t �u:���~F��B��Y���؞�W�A�#��#��B��A�_��w�?�T� s�7�+��-���"K������z�j�$�{fq��L0Ϻe?R�`-R��>�����K����s����A���H{,��U26ʐ����ͻݎ�-�c��u���;�]F�`�N�Y�N
#����D�2�:��ր�$"��z U�k�md7[墯��Dqp?��x�D]��2��p���1��Cnb*|�� �G�����3�DG&�Ʊ��`©�zM(أ��OpL��
��{�s�}�%�C�@���Uv���r��Fٶ<���y��D�M�؅T.��j�x \��[o����g���WB��8��QH��n#��y ��Rc6����]Z�9��q(B;�WXN�C� ����P�=���CA-%��o�Λ8��,U<�b靑�=)o�ᚰ�1ۂz?�lʆ���qe�{ j1�W����k�P�uO��n���1np�H��OgxU8�Ñ���eÍ�F7�×B#\�\ƀ�AU�(E�%kZJ��ʐ�������ݡe� ����sX=Ԥ���e���}*�??�������?�c���>/�F��.'�{}(�(���Z�8�Һ���������h�į'c�Y�ƏC^�{c]��oU���<Mֈ-/�:�Ғ�(%�|��#�9�Ǽd~���|A�%�.����[���>f�f8-�hO�Ϳ�P�_�'�n�톌��[��^�Ns�'�Ӄtő�zN���D��{���v`Ĳ�`0 ��[�l�BCD�^�Iт��������fC�v�u5s�O ���R�#�υ	��F�PS.��7}�gƑώB�����i�;��W&��^�]�w��%��yW�3�(�T��1�oӌ2Z9Jn�+�G�jr+��8������d�������1�&U_9�i(���˚}�^�[
�dAJ��I��a.���Ȝ[�M����F.�
#��a)�X����)��,��%�sR?}	� 9��Ã�����f��5XP�$�6�8Y}��vl=�iU��^ĝt�9��q2%��k6�������C~g9vh&Yh�p����%m��⹔	���\��jz҄��(����P}fΪK��ƞ���-��+z�pL.��C�����:r����^��pmx�Ѹ���~��*��oG�M�Ob�i������mY��:b?�s��F�:�e��`8i���NQ��ː�O�5��ظ�����'�-��x8��~�.a�N"h�2��s�z��w/�H*Fbn�Oo�Ǣ�i:4,�� �aC^.8�(+�j�nT�>d-��(��]{)$��;�^nY�����wm�x�}�e���r�ĥ= f�(0^��!-gFN淛E�9�`���������[�F���*�0gĲ�`0,z�F���W�!	��H��-W��]�}�|É��%���'g�=���z��y�)mn��E_;����sNX���uۈ���Xɑ�|��"<����\I@[_��Q�EO[��l�$yg��oo�Ke��ҧ.�x�Ic���ϭAng����ɽ@����-�w�1;��X�Ǒ���b�ѧ\
6v�"��}~�q��aĲ�`0,�%U)�+9�[y�pR���LطZ�]�T��b�,n�O��+�x�j�:k����ۨ��a'﹡!N�8N�ގ�$ǚR$/ڐ�a��2��զ[қ(�n�����gA���k\wjP;��ט5����܁�A�!N�H���8�c4/G&��->M�{.{_z�*��Y��2���9�
�ث���yb�˛��+�D5.�ƻ,F�:������l'��9�u��3��]K"�JT��P
E�>�P��z��=���E�n;���e��`8
���Cr�m0������߹�j��̃�K��"��kǰuեH�2����z��Qj�p�c�C��ͳj���[{cJ��<طjuy��V�VN�#�4d��\+�޵
���/�P&*���g?��qh<�y��ʆ����~d�9���|�f��y&W۶u�b�g���-uV��c���k� �yq8����p�l0KA��#�'�V�e�_�~��߻��;��ܹw;���/L�5'�G2�Z�>��5�����{&��kws��P�Wx��T�	��v1nppbY��Ir>>���Y�q��m�n�qv;Z�2K^��3+?��h��t>6.#��at�d y��lg�X�B��
��Wy3`nt.a������ۂ��ͯTo��,e���ۯ�8�k�җ0��0��d�%�Y�������b��.�ܼ���0qCl�6^!\���`b�c��Io�O���-7��{G���Z���Ã{z�t�Ϙ�/^��I8��03\���~s;����I���m�q�lx��Q�V�g�	+���Zy�C��q�mB���`�<��m�?%�H��6|��u{���$0����K�/Q�~�%���w��_��R[}J&վ�'�<M��0G��N�s�f�[$f�7_����ʂ�yJ�	��=L
Z虝l߬p���m����/|�]��빮1�Sۂ�k�G���憍3N	#��H.D��W�Ɓ~����`�V"�^�X��(��Q��v��Q1�����S�c����nq�ս|���r��a��ЃX*�1�D!��lFû�C��T����k�s�n�C����pY�|/�Z;4\F,n	�}E�n�Aa�|a��Ŋc�� I�Ư4�>�/�x��s�zQ��#���
�&���;��pb��տ�7-̞��W�?r��.s֋Ϲ҉Ɠ���>�R���ʉ��CID�Er^KK-���_�բþڮd�*S����r�V���s�y�e)���^������7����$���
�ӓ�&�C?�%.��)ya� $�Āݠ���+�D�{���k��y^8�u�^L7����{xxp����v;�����>��:rG��6M�Z'���^�!���󜷬�������'*o�D���ea�;W���l a��5+�=+��xm���aĲ�F!"Lξ@ㄫ�ȋ���O�|�Ϧ���@^<�}��;�1�!�;�ͲQ�cA��nb_u:����8��`W�U��5_������r�<�����7zr�$��ıQ#��Q�c�}3����"�x�%�n�*�W�kn?�@3A��,���_}���0pNnp�Rx����eO�,���1&���u9��� ��C'w`��񪜈z��"����Mc��;�!{�@T
��ƒ'Y�J�-��M�y�8������?x�mAƸ$V�<'|�����C� ���[\��>�sY�l�����m6n�Y#���~�נ�0F,nB�ɪ���86?H$3�cCj<�����4ao؇l�b��V�He��p8H��x�2!��!|q�Z�`,��:���R���1�f��X/�E���o���qY��:�DXu�$[O����`��? ���v��V1���L��0�t]����d��4&��H��v۵�m��#c�n�f���6�%�gom�p�l�y` zT �o;��b�&^^�����S���$��̋ nH@&c��;��"7�Cl��(1�GBH�	Qac	Ig�Z [��pƐV�{#.�G"N����}��E�a�`0,����䲐��C���3:�!�4n�5�,!k�WD.�W+�}����F:�G $�};X�J�2��:�M<L�0�l	[}ͯ�e���o�_G�)al������Ƞi���S��~|3B���ˆۇ����W!�E�r�a1�\^Lҷj0����=N�i2_:Ĝ��i`�3`�L���Ic�!2Zq{K���YV�"[E��ᱣ���H|����e~�k��s�a��r��I�^q�>,��~�u}Y�q�۴5m"�������ܡqĘ�a&�<�%�	+�t?O�3G��/�)��oqb�P��:���0b�p�@K�N1�f/d��sa�j?��	$I����w��_4Aft�����&4h����Vta�;��c�q���#��.�i�td�H���6kZ���G���p �`���mp�vEatpi9�rK�>�x"���g�U�</�t|���N`�+]K��Z��Ś��P���`0g�ˆ�p���1[cH8�	�?��p�7�t�<��=B[:q��d}���z�G5C���Z��p0�����8)I&6i���|�/3�˶c�mg`�XJ�	1�rLvg0Ί,3BH����"O��D~�O$!�\�t���]���'�4��sj��*)'���!���697���}��`x�փ#��6$T��pA�l�q�����Q��ғYF�B(C�0r�Jf����Ka���B%.�"
�r Q�j�bES�Y�v���uV�!�u^\ץ��9!�'��x���N�OD,֛;���CkI ��>`�b)�F��}h��`��: ���yz��1�� ��ӡ�Fm\1Ŕ\�ƃh��`��,A�-P.#�7���4L�O\��At(ԃ�0A,��%��e�^^�Qy#2���t�e^���s�e�Aί��ޮ�'��.,\������~mUH]������"�1I~ ��h�=�S����v�k�ӡ�G{a0��j0b��
@�rJ��x
�1hM6`���~���PrC�{�P.X�;�L�����؁X�謍� ��z��B�l��k� Vz���v�~���ƃ~<q�P<�ȼd#��`8���8g��`0�ˆW���ɪ��w7H ��>��@,b�FJZ������0��GO��!����C�����Sj�5?���HV�0'4.��zę�z�8���k��4���H�sh��EO��p4Ԙb���aIw�`Ĳ�� p�����P��3�5A�gXr��G+�t&�ʂ�9.�i �o�uB`�7���`�*bH��T6N��\\��U��e����?��`8l\1��pY�l�=���!��Z���\���VY�Ao�U̕�Bj,Q���eҧt���Qa�B��=?���PA}��\)j ��T���sM�`�!
�Fۊ���!I��E�*��w=���^���G�7��`8�@� l�b     IEND�B`�PK
     #{dZH��`�b  �b  /   images/3f9b3f3f-db41-4a6d-b13c-7e86a7741a7b.png�PNG

   IHDR   d   G   ����  0�iCCPICC Profile  x��||eU���4�K�ҹġIr=g��3�0D���d���B&3�F�� J�6H���U)RD��tA@@i�Ҥ���}�>;p�{�{_ s��Y�������M����/X0gT5I��[4�=ybuϽ����j2���l�l�?�pAKWWG����ٟ�O���f+���Yw��$iX�_1�`������.Z@�ĳ���~��a,��D�r���'�7q<�ݭ�S�d`���!Iƭ�?�ha��������sA
z���w�Ag��3�dUH$�5g��!��јs��>7I���xV���=��f��[��&�I�K
:߯��uZ�ؽ�RƚS��L��uRu�Y�����m��d�6ei:0c.kb5֔i������);�u����:{��l�tE2-�JX"���'U�)~YҌW�Yb�ڑ�&��M2+L��w8J�m�&�+p���	���@2#��\��,���5x���o�k9c.�8K0�vh�M�����,<h���_�txh��E�h�`�}�@���'!Y�m���|��_z2�%������v�EIҶ9w�m��$��$Y��ض�N���N��� ��)�J�����������i�y����������ÆU6o�5��phÙ�5<�����Ge���:l�壞]���F_:��1��sƘ'�n:v��+��c�wԸW�h�y+�f����x�-W��ʏWX�����X��v�z�j-�ݺ�^��5�Z�5�\�k~�ցk}����[�u�Z�����{u�ÿ�ᗮޠm�?mx�F�lt��{o2f��6����=��q��-�-no<�˭�O�ݖgm5��v[��͵��������v�4�nީ�^����9�/��]�O��9j=�t٩�w}m���qh�w>��g�\>���&�}��ڵ�}����η�n�պ����z^�6a��=��s��S���o����}����;�6���l֑�ٯq��9�����C<3����o����6X��u=�;kv�ky���s����{_?᱓�?y�)��z�gu�g�朙�t��:/|���_��u/}ⲫ�8��}~�r̈́k?���~~��1��]o�����|����u����{��'?x�Cxt�.z�wO5=s�=��S^���ޯN��n����ķw~G���?�~��G�~��S�bE�W��h��(�v%%5�6\?j�QG�zs���>c^{�u�ݴ�����|K��U�_��ՎX��5��y�Z׬}�:����^_����pˍv�x�Moz�f?����+�ɗ�4�i˖��m=k������������jO|�����C� ��5�zzc��m�~��e;l��.;u����9��֋']�v�.�O~y�w�1v�M:d��S�N=�����~�w�������=���G{�������o�}���a�)}3�.�y�o�>n��]��5s����濵���Un��i�Kv;p�.=��C�:t��o����=w��G�rT�hq����y�������N��K���ם��S�;��ӯXv�?����<דּ�>������s�>������hᏇ/:��.Y𓹗�\��e/�抵�l��ë>��㟍��r�:�mv��?�7���q�7��b薅�<��cn;��s���k~��_���G�z淯���=����}����^x���=��#���]������.}��'~��<⩅O��̴?�?�ӟ�s�>��_�a�ǽ4��ѯ���J����z�����ߘ���[K�>���s׻Ͽ��?7�`���������>y~�w�'�jأ��Q��:fԻ��F�4f֘��9n�qw��`�v����ݕ嫜�ꉫ����k\��kݲ���<��K������6�����I�-����S[���q6ܲi������>�.���۝�����n��}����5����j�+�U�ۯ���w�vG�S��S�����o=uҏڮ��7�����ww�tl���)�St��������<m��-����>{�����꛿��?~��}��o�o6�6c�`�̡Y�g=t�~��Ü{�>=��ko��-j[�ǒ�|�	K�;��Cn?��o���_��͎dG���1��{��w�����;�֓����'?s��p�˧���3���;g�w��gp·?��������.���O~��"��O���]���n���+N��諎������Ӯ9�ڋ����~�����MO���/^���|��oo��r�:����[�&�k�߶��{Ϸ�uߜ��<�߃s~7��A��ѿ?�ѓ;��?��ӟ<��{갧?3�O��N��n���|����~q������{�ѿ����������/}��7��u�������#����7���õ>��/�q�'3>%$ё�0y�aR�����g�=�����4���د��y����Y����W�p��*�]�U/X����Y��5/[뺵o_�u�^�o므|u�)/�d٦7o�lu�[7������n���m^�����mڮybm�������旈k�m�^��y��u��v��:;m���zGˌ����>��_����o����&���=:�N���[���ݳe�iӏ���=���{�����-�5�o�>�����w�xh�ə��zq�[C��ڜM�6��i~ׂ�>b�E�.�Œ��Ao����������_r�)G.?ꎣ�8��c�[��	�'���yҞ�8y�)�O=�CO�����8�ǜy�Yǝ}�9����sO>��ϼ��|�Ew\|�%��ɓ��q������^qΕ'^u��G���w͉מv�9�����p͍7�t��w��[~��'o}��n��7�|�W�z�]�;���=�޻�}��?��Ox�����C����;�������ǯy�'/���O����gN�ӱ���#�;��#�r�G��ݗN|��W.��e����]{��}��7�zk�w�G�;��{�{�޿��7}p�������۟��ӏV 9,��Y^�2I&�+�zŊ��In �]y��X�ƁI�J�r�I�����/I2��I"�a��G�lu0Ǫ9.͹�g�[��1������Ã����&˧����,�wc�}�J;�]�$#��j��::��&��F�$����{_3�m��u�:�����W���u�� ��};0{�^o����+r�����)E�=�?�Ư�8>=���z^�3�b����F�6���������_��S����|=���+����;���^���h;s�{�
L�K҇���������%�����Rp�8d��-q�~!8�'�������}�[ ��@����I�ecv��2��	iN���V�c>�~��Y�b���E�$�A�¿Sѫ-���c�V���E��"7R߈l��R�ԭ��D8�en~&�v��d@ݠ:�\��1�K�����T�2r�����>��9�ƚc����܉��rO.æ+l�4�ɠ	|D'Q{��ɠ;�F}��CCsI�K 3�����e~��ɛ4J�OM�i�����D�9���?�I��f�K���s��)�Jad�H��J>Ӈ$�ğ7��6�s �m��9��|_�P���Bг�ۺ�S�_���c���3��B� K�9Y�w���j�Z�Lj�i�n���]ml��tΜjk���}��͟W���5��:0�xQuh����s�?��������SZFv�1�p��`���Jkw[KoۤjcO��jg��*3��n/�����@#�����������Sm�����ѲWc��}�䎶�I�}=�m]���pS;��&w��U�a��i��u�S���ۺ��ݓ'��7Vz[�'����O�����6��ڸgs�Т��PV��%��_�5<���:�������
�Xe���޽��0�.�m=�V�L��_&�����c�Yc%N����������#��1�R���cq}��:Y�ъ��2cҪ�5�5ci5Km-S�2�X�2�����}�I}�S����ҴڸW[Ocez����}�z�Z�0����}ꔾ��==�;�<SebN�bث��"�Ꞻ��4/�60����Smn��WBI�Vm�Y.�Q=ph�� LS�5S�5^�7���|kgO�ղk�6w�0G���J۔I�sW�N�i����,��p�� ŉ-��a��{۔�+�������uLkice�v�O�D�♋�}=�^�����9uj�#��Zz[w��i�}Z���8�����}�1F��)X�E*Z�2�sb[w6�K{[Ǥ���"����ҷ�Vo������)ib��w����$��t������	id�s����T3-G�Qɠ�1~J+k��\����i#L���k�^ӪQ��ǫV�O�*V�¤������a?Y�[�VFd�qn�`�Ƭ4iEUY�M}?V3BI�5ոVFq���LY]�U�~a����LUeM3�-�'�L���(��~��ha���L��b���IU������Q�Z*YZұز�5�	a��B�X���J6Bc
��Ѡ��Y���m�Y�Ѧ��P�BFEG��ܹ����9�,ȸ�Ry��Ŏ�f���F�ʤ��7Y�����BǬ�f��g�3�lUԌ���ɒ�/Zp�f�N_gF�vjP�D%S%�X,^��2LB�X���k�Ӫ����k�X'3���괒!bߩq;�<u�zf�x%�d�q��,SnG�'�&,t�ɘf$%e��*��ki6n�v�-dꦖBFgj��SO[jݑI�2C#hK�
cU[3)�d�uؤP�#n�V�XF(�!ѣ�l&3R嚐q�[f�d�B��L���|���Ab Ў�W��f[=��5�j��j)穵8�LèI��	Vc�hk@p�=jJؔC�X���s�#�V�T�t���3ȆA8-�IE2�'8y*r��a��Z�{���9�:B� ʤ Xʍ�E��@9df�&$w=c�%<F��b_
��% h8"��Ba��B�T�����KY*l�c��9� ��)'�j��E?�L�q̎�� [&qPB�W�;��4�;�����d���d� ,RK��:���º5��4�� [
�0DHÍ�%
kf���ּ��yF^���[XGF�ь8h�&�z��]��?"w*H���T��#t�f�`cF]�p��@i�ƒC�*>�ђf���Z����j�6�C	]`�P�`uذY� B�pR�`M�*���*,D��o~/��B�
��YT� E�JK��N�L?������*ظ���S�:f�8F�PV8d�?Ο���J4��J��NW�v�G�TR	I�($���#����a���� �T��x�x~@��_�?����$oKl��T�!~��
�e
�!UCH.������掟[�*�X��E� M�YO�L S
���ʤ�����ai��8�=��j�F�x�bh=�_G��X�!AG��=�8�
\��F*]O�_�ʪ�L4�R*%:�q��C�u��J.Hi-t#E@b8[��A�g5���K�0qR�h#*�mj>��1#�
�����(��U`)���f��4�����eI�d*#8����0�#\��(RUǑa�:s@DV��A������Y)L-�\ ����j)��i	A�s��l�"�fkLW��X��#���O9Kx����VTV�H(,if=�I��;H\��W�<LTUplG���X	��!�1!��W�a�ȴ��)X=~��q��R �!-K3f�Q8Z;�:�8�����	�����T�]->Gb�<Ӱ_K���#�a5 �J���� �����p!��L订tI��2�
�ǂHL��A��V�$k�3"�"_�(�XC@��U�-�tbn{j��'�2�'�Y�NK2��#�I�ӌ2(#,�4�9�0}G�Y#�i�>�I�֜�
�]챾#���52S#�@�!G~W�|D�V���4yE
��^����(bG]vD� Ԟ,����@��;"�"�3�� T����G�V��f r��S�=DNxI(��%�c<J��g��C �8d�
�E�X�,c�Ȍ3�!Ht��v�+�p������� �G�)���O"�Ü�w���T	y i;�SVǉ�w�PC�GP�����XMY!'�,���:*	KhP2a��Da���52���
�ft%��E����F��$g�h�+F�LU��t��N�G5
���J:�� �q�+�S�#�*Rl1��u����#�� �I���"	�5i�TS��8#8r2J���w
�Z��g+��[�r))Ȼ%՝�g�����;7,�S�CV��蘕t��E�-B�ȕ��(�{��8���+Z �U���92J�,�#��K�\���!/�����ci٫���dq��<�"ˈ:(R�*v���g�W	Qc�GDd��C�xŪ��q���3��U@yKf�t]�Z]�G* ��l�Q��Qb��8L�{��  �0�ܣ!]��RXA8��=i9`#�9(�$�X%K�JN�`�6�4�0�Q�)�0W�K���q����*y��3���e*$UY�k��6-yEr@���E�'/�Q	�R��3�Z��SO 	�S�8ר��ԒsEz��
pU�Ҳ*r�
���Uu��"�p�!_�,�#=z2 rIՙLH�:zB��YVI�;W����hW?����LQi�,�%=9e�j��U��L�h��<���R��!���^ʹfM0������U �B0����Sp�焝Sϲzr�I���&�[ 슞6E����@� @��S8l���|�[��%&%D�V�Ef�jZ�:/�P�e�SHq9���ef3����YS��$?��XC ݅=J��S�t�� ��y:�)S+��|5�S�8̸OlN���Z��*�L����\a�>E��)��b3���%=�gJ��$ y0U�e� 
~��)�H`  9-S"�b�*?�
�J���UX��Bl�ʗ��7�m�X�׌�-����΁g�8�Oդ3V�T"��|_J5ɼ,��<�A�p���������T�cT��2(�S�x͸OE�{�}S�P��˩�*�Q�YXJص�:�q
hK:�t�׌*A�A�aC����;$z$[S-��T-Ȩ��<�(B�`z��W�ȸ�<!)F�;�88'��iLaw�)�r�%�m�M(�A� q��srK���䯩䋸B=q�4'+�&E����+6���O�es^�腨89h���a}�p��1�Gb�ěD	QL�CaܥS�K�M��"�/�Br���.�͉@���e0:j����8���BZ(�WK�_���C�r�*�ܳ��sSŞоT3W(Fz	c&}$ᢧ-s�EO���v%`9MVj�S���x�
��j��,S:�0�Ŝ"+s�&P��N��W��,�4'#ۣ� i	���˥$E���$�P��*T$�W׸Z�;º\����'7��S���'=(b����$��0Xz�Z��G[!kԈ+TK5�x%�7�C�,�Q��3
�b�=�R��4ͩK�f�}8Ah�
zJ�����>iNS�3��܄_4RN@z+l���O8W�Wm3dEyOC�V�W�FR��t?��!�T��n����(*K�=����)�i\
?$YIςPT+��Q��|~GB��o%/��'Pa�e�OY�����
:O)J�mѓ�H*�-��~���S�e�z���Sf��vi(�&����*�7L��S}���sJ�td����9��� o+M�xx=M���=��m)����%ϟ�k��rD-��'���?#����z*	��Ա�L@�F� �S��2�ZU���2�e���
=r�\O	���e�4bO(�v#�g�)��ڧx�>?�M�>����."I�>�x%J�m�Uc(��b�e�."6Q�$:D�hbȳf�8�(.2F�UeIU!3�-��r��I��.wP�T]COK�����(�ʷa��iʂ�HM ���%z�A}ᇔ-a�&dT,����Hm�3�X��t<a��wQ�L���f!!=B��{��P�E�[1��srðOw#�\��OC���&��4��ㄤFV��{RI8e�e��pW����޴(9ƸO��p@'��Ru���a�?�,E���e��hW���_tv�������\��YԿh����g�~��&�a���&�60�ڼ�]�i����<κ�<3#z���fd���.�Wm�"(k�A���DS�=m��F�"a�yOZH_���̞?ܷK�ܡ9K�����9�6V���y��3�,�$)J.I�u������:$����AqG��/"/�3.")�P�D��I�+%���N��4���s���
G�	N�@{T�s�tBrOr�kQ�J1����s^ʋdn~�����
�bD�Vѣ=ת�ԅ'��V���xΖjp�j`&6_��*��Z������"���ka'Y�*nf�"�"0:��VpOJ@��D���/-!�[9���9��y^F����[%�Q �bgN���
Z���I���\Ⓔ�`)���)=�w�6�.<���� :�|\I7Y�٠T�I	[�I��+�N�X����ړ8,��"E�o|7x���D�|�*?�j���y��X$j�K?���ڦ�T ��lVӅ�ub�7D7И�$���f<�p�p�g�y23~9\J!�s��µ
�$�=��S�R�x�SʜA�p2�d"��#1i.������nk��ʲ|\K��/�.�z��T�oSЅ��
�ΜB���B+s�c���ɒWZ��߬ĺI�s^����z�/!g�w���*I7hB7�p��(�V�a�He��F��ש�k�0]�y��m>?�N��4s�3��k	F���.ʵ���y��qG���V!1H���ޜ��W9���Q+F�{iSF`,�y/Xn0^x������x9�/�ca��=���n�:�vG�cR��0׹�g�:�
Я }���0t�����$l"�֑����l�6��e��4��5S�,r7��Z�7D�L�)�dΫ�a$>�d*�'�]�mf-B��L�3�M��.=��/c�K�&+H�ϋ��x^�_�r�&����l7'�<�t�U'j��f���%��$+t{>��M3o��OrxaO^f��r��d e�I��k�BԊ���$�?OJr0�7Y��t�/Ge��h�yU~+��;Ox�б�e� �I��#@��ņ�lP�p�Z��D������o5�ҁ޺q �Q:^2/�?A'�����ij�>��0A�#��:��n;�1m:'S�f�(����"g�	��Xa�] ��q�EC��	`�	�؏_o�����If�m"�k���aTު�WO($}�$'�.��-��3���������8�u�3H�K�B��a�o���/���ɃLM�g,wQ��4~�Ț�' �q�g�P��R+�R�Y|B ò�/����@�ԏ���U2���LN"��2�!L�j�w S�!�x�͡�k� ���]�yE^|u��e�daoPz�=�.>��$P���nd����=����l` 8�,�Fn���G�v2���x^�q�IN7��@��|�:����d�ې->g��'�I��Har��a-�Rxs�Vi<o�a�+�d�H���[`�z��-H�M����c136gl�'�"����[��`-�����#�!P��=��x�����_$���Ъ����pd_ގ![�Bk��"���iV�<dV�E�0�
�ړByA��>�GC2l��ܜ�{��E�s8�c؈ិ�0��O���!����GC��k���M
?n�04��K�PoZ����f��H*>y��`�ګ'��29�,�y���/eY�J!9%�~o�P�	�H��i��e�-0�A�0�)��4��F���JA$���Y�0T^���#��~�Aw"��,�E"S������p�I�V@�A�HLe�-0�x#�=�@�H��+"��4�_����$�3������37)������r��P����W��7b,�y�J��.�n ��[`�6`9څ�d�������i*����,ƍ:���d:�Zd1|�����0BF��y#�A�-����@���SD!)�*(y�D�`��FP����@*�㱈F�-9�)����*�Ǎ�4�)��$f���>�C]�����y���)�T��h�~����j�L鲤�!1�T��k�8)a��"���y���. �O�мJ*��]H���-0����"􄳠����-0��"����SD#�"���ҝQ��"bZNx��J��""��r���R7�������z'&`!AS��z#��r���	��� #��/���,N�
=��~��s�Ҳ�MK�d�0���Cf�WK*$�� #���jH�}�L�/�Kd�0���AKp���31ր�AjH:{�[`���*{B�r��R�0��a<�3_��HB
~op�*�@�e<o�a$��F�,'1���X1i�L)
^���[`L�y�	Rz�̥����'Œ�����,"��x�R���I�"����t ���T���LF#I~i<��`,�C�0p�<,�"��Y�k��;��6Hﱲ�Fҧ�M ����RF#��&�Oh�$}3�?��a�jø��ae��?n�0ha\"�{�#���g2b���1-H�nR�5D�V�C7(�_}���E�0�B� �����qHE#)��k�\�Ӵ�ۙ�-0��)�@�l^�r��Ak_@%!�c�`�*bEϗ�'e��L�����n�R�|�PT�����0h�60���E�M��ME�V�����+�:��-0��}�I�;�4��51�b�� ��5D覥�U��a��7��>��e�����>��ɂ�`��1�B���Kc{Ni��g*bzt��>e��L�:��F�"�*�~\A���Qݽ����Wi�㨈a�-~oT,���|�FQ�xeȥ������Q�� j>�(����,bE�H��sR�1��;�Y`>�S����(x#���>��ی۵>�@zg�7R�V�|#�Q�t�,I��cU�0вP��Y e�A��a �{U�wiC�JE�H�K��}8Pp+���#����>	�rU�>���t�0��B�V�sR��L�y��r�kH�L���mSGC�"�����ߟ��Fõ����z����!u�0:+�6�����I1�~H�z��`��T1��;<�Sa�_���#����T��9Ĝ����u�0�2_/!��S��a4� (*Vx����5D��t`0�q6Sޟ�a�ǽ�k,� ǥ��D���xՀ�Ɋ���"��{>��d*���U8ވa0��,Aѧu�?��a0����3�� ���[t�0�By��]�$=/�y#��)T�U��G�
�at�0`�M�&?��K�9o�0�"�IMR�:�,1��>k�;�wC��"��/T�PBC�܌�>���8P��k��	��� S�����G6��1�h���n��Ve|2àU���7_��{)a�à5�=M�DњW�+���*�ޢ�L��u�DC���Az������0�����k�`��M�0Ԛ^���'��x�DC��Гh�a���k��Z}�0t��OAy��Y�0����!p, ��#��a�+���+�7CUO���a�*}ܐ���5h1��ų�����F��̃S8
���{�4�CX/�C~
X��C&b0��y@=V����a�|B,Sa\j
&b�T�wW�N^�4��Fc���npaǀL���a�P(}8!���-0}����@�#$=��5&1���VNJ���31�=���N��!rx�c"�C(�������5G12;�i�1�p��ڲg���..J�ڕ���z��Ga����0`�a�t[=o�Y�-0�!ǔy�,�P=�l�7b��1 �I�5�וm�0��(/t��>I_��ㅍ(����R-�J����0H+C�e�{��l�.�y����=��Ґ��`�٢��RӰy�_}0���FC��s!�����6b�!�����	�[`K_n�7ρB�l��x�EC��}������Nů7b�d�+D���c���0�*�ab@5/_��?o���	�Dz�˼��xc�K7�
����'m�0��f �T�����:��o� MW���0���P��ǥo2��1���p�A|p<���gB7��AJ؈a���8����89����a��o���{:�H��F9o�a,=D����@��g��ۻh-��ņV�R�x�;I����Q	�/�   	pHYs  %  %IR$�   �eXIfII*     (           >       F   i�    N       %     %      �    �  �    �  ��    x       ASCII   Screenshot�j�Z  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:exif="http://ns.adobe.com/exif/1.0/">
         <exif:PixelYDimension>1018</exif:PixelYDimension>
         <exif:PixelXDimension>1430</exif:PixelXDimension>
         <exif:UserComment>Screenshot</exif:UserComment>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
�v�  /BIDATx��}Yp\י�o7zAw���B���
.�6J�Bɋ�vj��.�l���j��$���<(yɓ=IMeW�$��Ȳeylٖmy����(R47q	�b��ro��?��{�� h稠�o�{�~�r�.���8E�\.O���8����o\U���D�ٹ���10p���&Ȳl�
Gi��~�C��5�^�͛��F�����Z7��Ys^����fx.�'�7-G^�o��5�M���Җ�[h�ރ�<�^/��stm�"e2+d�X�E�yi�͟��э��J�y�yy?�+V��x������KK�3'��!3�S<����jY|���O��F`Yaiq�"�*y����ޡ|.'�(�"`�HD�X,�=���J�lyyY����4���5��+_�Sfi��5��ƆY^����$��d��6K��M,�qK����!�-��/~�S���'�+Ą��Ǒ釵D�B�0��q~�-:p`?E�a!��x��4=3#�p-����0_u]��X؛[�Q�����M�BQ�3rs��=��V!_���v:v�1���!�/..љ3������d=&,�����i�u���%4P�*Z¿���ѻ��ڹs�0��fH6�LWޗW<��%�+���÷XSF)B�"[Z��_~�_�
�Q2����_��k:��L�0��ݻvR,VE�"icccl2�d.?fSV�k�\Ő|�(fI��s�g9����4�2SdmlJV�9���r��~�����499NW�����%a�ѣ3��?������%�����e޻ɺ�`�/0~t�k�C���ޕ)�R�0#�[�$0h�*�+n%�J���L�$�k�����slS;���t{t���y]z��Qں���y�$Uǫiv~��i�yD]�����V��ߋF#��Y�u���hX
컚��6��^��&�aƹb�!JcC#=���t��Efƿ�ӧޡ_���4�Tӕ�W�w�}���o����s��_��y��/,P�5�-��D�h��/aZ�l���-���ǖ&t��D��d����E�fn1ff��Ī�����U�>����k}�_�˗/��������eW���$=p�քq�1!�)Չ?������A���1�b���R]]Z���&����M�3$E׮]��g�1crt��҃>(�C������z晏�k����<uuu���{��7OQ�ۺ��~����տ�7�����Ye�A���7��l@�1p?�1��lfʨ��={���W������`��oX�ރlf�"Q�r��H���	Yd�\�PϿ/�4WӡC����S4�f'�P}]}���oG�#w��x�>�����kdu�����E��Ps�fgi۶Fָ�����;4>>%�F..eE�H����/
c���VJ%S�F������ԇ>D���ML���,��7��{555R��M���'����R|�M�R�Ï�"��k���5�-�����2FHq|��̷��c��)%3.�f�]�8�N��ȎD7�0�ͼcٶH���_[GZ����ӫ���w� �q�������J�����-�|��y��(Kp=�+E	��)��'����uo�"vff���*��?@h �`�f��X{�htǎ��,��Ţ1�k��W��>��%K�.]f�7ѓOc��o���mv�ﰙ����i
#�"�h^B�5��Q��{�6����QJ�ֲ��]�!cc�b�I�h2pN!�� ���k@*|Xg�T3l]	�^{�7t��0����j;%����K_�+:�kd���fėī�l��X��x�͛;��_� ��5R!�� ���9�Y���ť@_���b�(��Z�_�����3Q���ߙd�~��az��?�;���#T��e@��5������lP�k�l��\���(��,��������Q�e���@}[��MNαt�YM'����.��MN=��MbR`��M��=����-[��<�-�z�����ʚ6B�w�����-�6e��}�Vho-kV*���=�]�.�q��cF�P�B�0��Ba��}�������2\&ғO>��������f)�����$`w���N^[���)3�*�^���uuu�u^���	�m*�%�F��9�4[8ˎy)C��,,̭+	�r��H&k==JW����U�>8H�E;����ut�3�}�N�>�����Q"eG����:�p5�%���>p�}�扷�~7QkӦf�q�kתhB��\[{��*��q���i;�+��]p䚡۷h߾>:п��:q�M];���n��g>��eA�E�/
������2�t�* |��!{H ��[��\	C�А��R(�J��`�I�$Z^�j壐w����kW��/���<]��>���H���]�gn�f��G���g襗~H{������K>�;�f�_��lR3e�Ȃ���L5�fX�͐M1��t����"(������ʗ�g�ѽ2�09�m������Rg�f:s�,ղF$�_=�Ѓt�<��ۣlژ���/�����!����t:����<Y:����R �����I�ji�֝��+jR�H�m_8TEEy(%���ݼ��o,���=�*~��þ@S�3'�ё�G�	{��.���"a����mJ������v��W(x�#���k_���'?aB��#Ɓ�I������K�=>��3�a����ξ=�ŗ��w;=���<���]��.��?��t��!I���#+󌵚$�ƜA�jY�d��d�Ѧ�t,a����J#��Hv��PK��rn����/}�^�56'��ܠ~�"��B�l�^{��4ű�֌���TY��9����om�D���g����t��Y���� _B��iS��\�Y �� B$��*�H�1м��]t��I��9s��x�ZF�};�$Az���l���h�hZ8�� �}����srq%���r5Z!k���-�V���Ǐ����4t�&��1��HRVS��Nz�x����>�]2�+&����Q���O��a�0�Hn^�fX���,� c�����`�`��/I�|��`�&V�'��r�"?�oK�,���xr�)�o����{��=1������[�����t9:��+Kf]]����K.
/Y4�3�G)��I[A̰"2�@#¨�MA�J�@^`"`�L��6��zϠ��H��C|Qώ��P��A �	x�R��$�/ {��Uw��ú^�&�KBT D�E��C�ZU�4v�9v����'��I1ψ��u�C�� ���Zbz,M|��-GC�pH���Bf^��RF IGu���# ��PA��D}?�l+x�AM�FC\������mW2�����՚��r�z �c���$]�|E�i�ozzvQ��]�3���;�L��Ĥ�����"
�iΛԳ�p��G%YOW���:�H�ʕ���Bʵd��恃R�n�x��c����|��j;妶L{
�b	S�͵���a��l�V��>�������tgl�c�IA�L�=�K�H����,����E�(+0�����~+;e�2���|$��*}&\���(��ς�rPP_�Bp)�9�o�{����&ҧ�"������k]�F��?a ̰1M��l���}�	ŀ�R�Z�.?!�������M�!�JHU

666S����"��i��mԽm�dyU�H�|!�+b@�-\�6Sy/��$E��;w�H,*y$��X<&H�{r�	��okE��P�)"�7��mO[�_2�T�������c����3]bU=į*	'O�H)�i�����O�x�谿sl���0�����LO��k�����ws4=5+վ��EFX+��O}��<�--,)������`%���Az�F�@*��(T';;:˘��� ID���t�7@Bs��,�Db�:����o�|�((����i�s`�4M*%�0��V �|G�a�&Ճ�	3|#�lȣ����J��L���)�J���&��ͫt��Z^]��:��JU.��iq%����4�R�%��N�֚�B!'����,�\_eB�y@ T����LE�ڵA�s��LfY8��{�6�����&�,0Q<^�K
"�s�Ht���.0Yh?�k|��ZjS�
x]G�GR�vP�Kѽr�byl��EVêdz$G�>J�c�i1?CM)�y^�^�!]��y]{F�H]bLH0E�
< � v��#���|X^2�j������
�h���%�)iT@��R$b&���HRq=��ftum�&/,�A"V��Q��p�\'&�*�[-�ebz�-[�k��W�����;t��g�9�A�[��ۗ&dFp*W��E6C!~0�Jcp�*tiG���*�n�x��T���#�j�6����D��C֠W/�JJf��*�ڄeE�1��<�U�Xh�9�l�qF�a�ĺ�z�<�-�P&����)�D��Hf��ŵ�aB=C���a��*'c>v�H��8����M�6��_�Sj��`,�3S�"�8�a��ռ,�B��c!���u�&%�c�Z%��J�bF�0���scR��u��KPm�3��h�J��d��:S�>�~,/�����=������!���`A���L��OU�]�0�e
����H����T3����&hp�ev�i���,��LfIl=�2̔Y���N>IgG�#ݝ%	�6����h���ڔ�-�d4�eh��Z�Ԃ��P�|&�t�ҋ;�b�0%��3����1�b�	�lso���(�"(�t����իW�	[�m��&ʲb�`�IQ�F� 4�=�@qD����PW���T�݀�YkOAj�wxdD� z{{5S*3���[�6gh˖-b��gvww��|�F<�9����o��߰_�J��{���Xڤ�3K����ч����M�X�œ��&O��z����N�3�|����-3�J!�T��0�%]��W�\�g��^�&$���Qq!
 8����g��01(��4�bb�oϾ=R/��B�,�̇�	ʾ�}-Gi||����4tK٠�r&��T�Ӑ�#C�ch�OV�	8u_ \��=O���(��Ч>����Til?+�nll缜Y�=ϾczfR�Ǻ�FA@����D:P�������|�m���?�nApzz�	]M�l�PC�
�R[���\�Zk $0�|]6��F�Ef��, ��2
wkQ՟<����
j/k�+V٫�CΙ���C�=;�,]� .Kx_D�ꑣ�
DE�jJ+T�@*- ������@�WH]�a��s��FKK�4���֊�C[�&��S�P �noo�nh�� 0�*��ϫ̻I����8qd._�L��{`���I1����[O�Z�g���{e���!0)VHl|��&�B?~e���,�9�a���*/P[����!W9"�FmJ�6 -!�J�ⶈ��rP�D`8�'GM�E�G��X���t���A6R��[�VU��}��oni��53tƀ X^n�$N
fЌfj�`"�}�v�' �"K%Vmχ�!2��xB/�L]�B�*�6��P�����9*PL5T�)�b	L��k�%����r�c�U��ƣ�����!�`�nũ�ӂ���!�;,�N�?պ}h�}I}]��4�5�|����I����$Aa��<���%!&j&�<�����M��h�yE������_ ���"\-�I��5&8t}��N{�f��VP�����/�C;��+�#�i;��Co���P�Dؽ��L!IU������ ��HXl<�eb�V3�K�Ԅ���Mr@�u�V10Y�!�v?���%�k<���0+���I"j8z�� ��!< +�;k5,u֤��7ri#�#����ZhjzZ�3�$�h�0o��h�-*���oh�N���:����$�iw_-M�Q�Q�3��Tb��Z ��2A2��9�B� P�e�<�2\�y�
T1@ ���)U/��wgE`@TH.$��f��C���kDCp-��## m�s�gb*E{M�x ��)P4m./Im�P��݂��ϰV�O�6����Fm}5�,N�_׮P!�@�����O�'&���_#�C"Y��ٴ����eh	�D<p�:Q�� ۍ~]8}��Z%�":���9˲)�� >L���+�J���+�������l��H��0�ý��iU�\�Ĕp8��<����K�р�M��>�ӗ~MN8O1@6Ǩ����7_�_��wbV�lӟx�=ʋ�gB�Dʱ 䦰�xC�[�8W�0[���M�L
���@x<PT�$i>@��������M^UiUm��� �<���TY�=K	���)T1��e���'���	Z�*�K�j�hvc��4Vh�1�����k�%��c/E��k
~p�o�����w�jv��[��#~q`�
������� ���ʰ�����q�V�� (�1���1�&����8[��������@����}����Vd�H�#$�h��&%%�-�iY���Q���Y�[���g������,J��%yf!F����t<t@|�(Kl祱�!L���&*�~ ��Gy��Y�"��?��C5AX�P@B[��+ƾF\���_�c)�T�21�,ըᘧ-��a��Ip=J��ؕP��̋��J
#��W��l���v��z|�e)���{nf�MQ3���*%��Tj>P-aa�q�����t�gs˲h8�|� �F�����Q'�TB�43&�D���1y!�|U���R*��jS�/О1��ϐ`�Z9a0��-3n�d�';ZY=6n�1�*v�_p^�CL���>$A�Sf!E�^���R��Z@��b�S�����x�ԭd��:�������#I�0��
]-5��a��E�d��s���bVr��Xֹ,�/#��CpkA�A��A�����uW}&���b�Qv3 <&��g�\������l�,���J�oMR2͑k,,�q�Ra�U�Ԩ"bi��䲩�I�D2!a�b���D���HsFv��nP��"����HE���`(3�#|�F��172�x� �
�V�͛EcTS��W)m� �4̓���F��%�F�IM��0���;�M
�4�r��*����l�z��q����|F��N{���@,!�(��|N.��,ŧdRm[F��*�D�]R��ʗ�0'���ׯ3�N���Lή���A�p_�&P�� }��>W���![�<m
�"5 "T\��▙�Y����%RZF{ a��������r��Q��6��N,P��B���/����?��46��*_dy݉���*-,��G>���V���������.M##�,u��.��,���a����Bp@`�[�� a�������h��o�`��1'�V���0[Аt�8wWy>Q t`.�z:̷��|OA"�|>�*��"f �aJ�����Z	�4dͭhsS;���X��Գ��U�R!KrD�y��{�?�C��"��'?�T]W�P�ue��6#��%FE�1�-�qE��i��
t���z�r*u? �M�9�Bm��Y��3l׮]�a"�����#�mQ�f[2憙�꽄�G	�a!Y��4M��U|W�MaS�IiW�9������ ����|�]��ʯ����̐���@͕�#�H�o$i�&���� �_0�ss�}Vs
���g\���*�u��-Y�B3I b�!��iS+�P��t��e1�z���6������ΐ �)�����xL�7�=q�Av%��X����Dh*����(��pAO�!Ʃ��=��U���Y:�� )�M=yz����XJ$H�yB����O_���e�5�K��&��n��}*	�R/��)�����BN�B��~��0�C:@0�Hj*(^�P����P�8�Ô�1|�
k�,g�33Ӣp�ذ�u�{�����*�m��5Y~��!��VC�S���Q8�(��c&\pYp��덇�BɄ�Bjy8�duBc���Y���\]m��hcU�T^�*�Z�jݏ�zA��J�m�K���(*�@�}0�æ�+��8xE���{@@��A��rn�!�.��>SK/c��4�_�Lo�X'�V�ST�ht���t��jhwO?M,]�ɕ^�_)�#R��s��fE��|X�l�'�����I�7�Ʀ���@f�6]�T�֘��g4���`�O�1Y�A6io�U5�$�&O�	̅k⚠�����(�㛙-Kw�佮��J�b�!�ܩ ,*m��ʱ��~��3����s�Ԇf����(p��f@[��T$(�68_�	�l���Ķ#�FI�+�-�neTE��6^��ߟ���'|��]�D��k �݇	�C�k�왤u�h�F�%�^D�Ӏ�|�&�ҵ�t��9�s�gS��7^yB��\;mI�� �������~[��R��&&&�u4��B�����t*�"4�c{�"h:_�9r<��?b����������]���XH�:��u��dT%e\L}Y�BgQLl��I	h:C�~�$�q�=��WW88\踚˲?hdiv��ɖB���ІX�Z\�t�M_��\���
(��A�����3�emn�һ���=l2��D�� �588�k"1i+B�Q2�f�SGG��2CL�DP
8�.�U�4�ՠ}���˫f����A�o�J��0�a�h����%8F��6^�ی�(�2�\"�U�"Yd�]�U�4�f�"��^K�T�Z���^�(�LK��N>C�����&�c���h
,�R��
q �\@ö87�#Xv�ڼ���##5}��_�(�2��91������Cv�b�����at�@�{��m]�����*פ#Q�-5b����z("y���ײ�l�+�?x`������:�WVZ6 �����AF?��BR�}��W= �-:P,2f�r�N���d+c�	7�DE>��j���� �d�;sUF2M�H�m����f�T�	�q&��>:������f��&�9qg�ěJ�($`�Z��|�,a��o��K����)̩?����%Lc[��D4 )"VI3Dv�3���G��AڨRY����0���B�Qlc�7����d�d�m�rd��m�E�s̨E���$P�gr)�k������%ѐ<��x\]������>�QLAY����ڊa���t�L�.��X,"=�.��5n�	5�*��:���^���;���A+К���"���|����Q��pӋ�*�H�Z|���I�^
Q�9�W�����ÑG^�>�IG�|�;^7����D��t���f��A�Q���+��z%�c�ض!30�R���
EX�ZN�}"&�i3Q��֋`ѣ�4��H��S�I>��Nx�tn]ݔ���N�I�zBU��Zm�QZ����e׬e�=���|�,��l�s�΀�戏?u����:���c����	ܐͮqn~m��2��->��/\8O�)oܼ%�"�Ro�ڽg7E�V�W
��W��x:55)��!^���c��.�S(�~�z�+y��:q��)G�&��| }���wg�����?�)X+6��d;��bd��71",�`�x���ܔ��"�Hb0��J̔:��w����B~����H��K镟�L���9��˿�mۻ��_z����?M����z�e�@�|@�P|��I�sgX�`�Pa���0C�Ξ��7��4�/��g�0d�.?��?O/�-��g��x���������=LO=�a1鹲�7w*���(���1��~ ؐ!��4>1����᠘��<��|�皢{Q[�~�C����_��2�46�cǎя_��[��.*ҙ�ޥ����{�	9i��>:���{���[ζ�6x��\�~��6��C{8��˩�/��}�+M��햮J�s3�`�����NC�X�z"�G���h�(��R�Ο������?���N�����_d959΁��t ]�HĥU�|�a�?v�6;�,E@�|||��F�a��"�8������~��o�b�/�Fwq���������&&����M����@�;;X;�$�r��!9���>��w��mff��&�Q^{�m���\��-��_<M=�=t��E���{��7��m!�Ґ�0C^z�tm�*U��nji�x�E�@ ���9�1K����=��裏�r�����83�]L��Wd���E��Q�8��\
q�[B�馝%h��:N9����� =N8�ǫ"ձ�����ݼ1JS�����O�	��Sr�/�S��E�XPS���_�U��C�Ϯ^�D(z��5÷n���<��.z����o�O��L_x�TXR3n�;o�!DA��-�����Z�ǟzR�	H��� 
�r���^��=�D����i�r(����j#� /���qf�;��x�t+��>�D���ͱ���)D�,}����3L�_PSs<���o��Fo�R�:-�Z�z����.T�6���^���9{jvfF��m�6��U)l�CS7�u�'ޢO}�S�2A�ӧN�)u��]�����4?7K�L8X��՜9���LC��X�C�`����bV]}�4slȎD�:O`�8�lm�\�\ÐTM�g�{^s��fV�K���eL(]���h�����9)�l���vt����F�
D=ń�f� ���"��n��L��^`�<*0�{vjJN$�|�~G�� '���j�!�煳��P�p���[���#�^W_�����kT��B�P�����S����)d}��7͡r�ѹYvK{���$���A�b+G׶9�|�aT���Ul0��'"\9V�����A �2W8$g��X��#kg�084������O���qq�ȑ�4��QE��\���ր*���|}�z�ȡ}�u�f�bi�36!SIw��a8�(����	(��rˌ�q+g],��d��<��hk��ԅ�mݲ�������^��ke��hEu���2-/C�^M�=�!'d������-���F�8�bB62S@+�Ƣ߅W,�'�TJ���������&j����aw�?L�H��)��Q��h��������D*Rѳ<xH��}���Т���r�#���[E#���ooO�@؞�.�j��Ժ�tR$�FS��M>.�������jAzŢ�$u�6��R��H������k`�bf���h����DnW��<�+_��\��v����%�޸k�^W�(�F/.�
$2m�4��𳫖����!]�D���d8��g����	v£�s���W=[�t�A�	iñ�9���G9&������~�II��q�N69��8������0ML�K�̬�{�Q���Jif��/ӥ���(?*�Duvlb�ɱXv�����.���2�(���|S��R2�YG����M�we�QN�d�%T@�ߵ�h�b�v���v�"���'OR��C���L��jSL./� t:�X�չ<mjk�Vj+�Y�G�0��C��ޥL��9HL#�����nA@Em}Z��*���ܲ��v�����.]<G�&�w���-����v��5�(](`��`m���$A��u��=�,�p����	)A_�S�&�=�	�ڹ��R4Bj$�D�Y�hu�3�
I�ND�T����l�q:αYF
;R�E����V��bƿf ��e{&0wǎ=�,]fص� ƪ������X�,]����U9��,�3ȓE/���oJ *�kN���`��rNp��FX����z�������/X�9v�,��g{_�Pi�$�E���i��>
��F�<�~S�i�uF�KR�)��Ըl��爴[Z�ş�1���Q��r�B�W�1��Ni�2�'��/���U��Xڜ��lm�w�v����-��ևLFb���iV�k�,
��e��S��#:�J檴��k�D��ϵ�Y˕�`���Ťl{�}�����YBLU�    IEND�B`�PK
     #{dZ��_mE E /   images/28139415-969f-45d3-9930-3634e76076d7.png�PNG

   IHDR  �  �   ߙ��  0�iCCPICC Profile  x��||eE���6�ѫt�q�"�����ٰD�ݐd�b	!v��X@��)�p��)"ME��   �4AiR��=sg��E?����d�y�3��)�s$���?��j�̙�p�{���{�U]�d4�[?�l�?�`~KWWG������K���f+���Yo����$iX�_10�����K.�O��ĳ���~��a,�;D�t��ONo�xz�[A��[m��L��}��[�x�$Y�<M���>����4����93f$�j�H2s��9C���1�.�}n��9za���$Y<{�u�s�A���M
<�t�_��˴.&2�[���5����jG���3�l�4I�4m��t`���j�)�r~SgSOSvP��Ń�v��d��ɊdZҕ�D$~wK��S������Ġ�#iM&�u�df2����p2�$�$MhW�L�_F�ׁdF2'��YR�/�k��Չ��r�\�qc�m�ޛ��Y8x�Bzm�7����Y�-д�j�܁ZIOB��ۜ��yN��DlKH/����m0���GIrŃI���m�N�5�I��� ��)�J������}��c�Ӓ��ɵ�m�ɓɫ��6l� vmا�І3�mx��Qk��FMuب�F=1�2z���^6��1��sƘ'�n6v��+��s�wԸV�x��+�v�MV^��C�LX�;�<Va��+�:c�?�ֹ�]���~�z����r�s�Zk��������:��;n�3��r����^����F_�jö��с�������M��l��n���U[��|��ÿ�:~��p֖[m��k[_���_���/l{IӬ�k�����_�{��؅�$q������M���]�W�o���v<p�c�vf�eom}t�?v^y򖻴�~��]�w����ԍ�Zw[�}i����O���5{��k�7.��ߞ�w��o���i3�ۗ�<r���5�?<�ws7�w����w^p�	��?h�%KY��Ӿ��a�������1�;������=i��ǝr�i��?�QgN8���{�J�-����w~r��=?]o��^y��W������_��uO]���ˡ_�r�6��~�;�y�λ����;�������#��x�����#�y�u�������ze��w}m�7&������/�k��O|�����+r��FCF�+�(�����Q�:b��g�d���؃ǭ7�ƕ�]���˫�\9w��W;b�#�8nͥk]����ܾ���y��6�xõ6�������N���[�_}�1���7Mh�r�V3�^���_>{�˚nn����W^H��>�be��Z_ob����m��l��v�y�������#'��z��������/������i���mʜ�'t]�۽ݯ��<m���>k�c���^���#�|�[+���{�����2�7c���}���Y��p����z��s���7�2��M6-�~��u�В%w�Y�.��M߽�g��U��-����=��uܢ���N�����W�|�)�8��Ӯ:�򥗞�������:��������?���;���pя�d��.>���?��l��_:�/_���+>����>���+׬{���m�y}�7�~S�/�n^�Co9�֓o;��K��׿��]�}�Χ��]o���=����^������c>��}���[��џ�q�c<��'N��O.xj����������-����0���/�~y��Vze�W��{�ͯ����7�\�֩����;�y��O�����}�ׇ��G���s+Ƹ�8�w��7��t�1��=4��13Ǽ9��q���c��+o��?W���|�3V;q��8}�ֺb�׹g���{q���0z��7�z�6�}�6;i��[�Q}�o}i���&4m��VS��{��_>|�S�~����-_�7}<{�����Vz%��]s������� wl�i�׾�2o�᭧N�q�5;�v�<��ή��/v~uJ���]'�vY��=/M3}����{�C�Z��+���o���o�=��}��������h��Cg�w���Ͼ{�Ss_������¶E�/�u����伃�:�C����}��U���HvT�ѻ3�{{�q���/=��o9��<r�ӧ<w��t��K_?��}�g�w���|���������.���+.�/I.���-���?\z�e�_~�G_y�U��섟�v���\t�����;���Gn|�g������۷|p[��;���f���ٝ;����޻�}��{g�7�������z谇������)<�������)����=�����f�_v}v�粿6>��c_x�����ˏ���Wn{����������eo,󊷮���8�����{o�k�k8���Ώg|BH�#�Q�Zä��>����G�ї�i�_{Ӹ�ƽ���+O_e�U^��n�+W�`���8g�׺t�k׹m���{j��o�𕍧l2ӥ�ݴ�3��_ܪq�/�;��	�my�Vm��6o�^Ӷ�k�e����Dv6�D\-oU��G�3�o۽�����q�N�k-3&�z����~��&��>���j:v�\2�GSo�z�{tτ�I�����{�f���Z��M�%�=�o�އ������xp��}���¬7�>��ٛ�i��㼮��0|Ă��-������A���Ρ㿣�����_|�)G.?���?�c�[����'���y�?8y�)�N=�CO�����8�ǜy�Yǝ}�9���sO>��ϼ���~r�E�_|�%�������K{��.?��<�#~v�Ϗ���kN����~�ˮ����n����~y�����<s��r�w������ѿwW����Y��U�w������s����`����������cW?~�����'�j��'���g��ˑ��ܑ=���^�ދ'�t�����W��ο?������k���[;������9�ݥ�-�׍����?|�߯|�������@��,/NH�I|ŊǮZ�b�����iW��+V�~`Ұ��R���k�L�R�H`�k��$[�̱Z�Ks����#u��xS���������k���^�������ֹw����%�������������8-I�w/3������u=���������x�ۿ?���D�̞l�����񊜡�!�*n�Ff�����+x�G�����D���W���������M��Fo�����������oC��*_��'���c��㎡�m�W��#g �N��޷S��a�! �~ �%��C����x�-��|��_ �y	�v7����x��k�"�|�x٘.;�LaAB���}�A�U�����߭+Aֱ4�m!�'�,P3��T�jK�$�����o��Ѝ�7"����T>ukjA>���AYƀ[ǀ�	��ݴ��P7�N7W/z� �b��!�)U���a��&��u6~���EX����,w�����\Ɠ˰i�
�>w%Mu2hQ�IԞ�m2�N�Q���c���\��bȌdD��q���C�&���Az���>$d����fh�Z�b'�E�t|
�RY�,��b��O�!�/��Mg�5��d�!e�l4�W�1�� �L��6n������>��m�b��;��bNV䝽�Z�V*��zZ�ۻz�vW[�g.�=���?{h����C��V{��g.���^X����9�xcejw���)-#��Z0x�Fc������mR���a��I��jf��j;�\u�SOoom�k�h��6Nj���hٳ���>erG[ߤ�ξ�޶.�Ib���]}����,�0@紎��:Ǝ��}�m]�������+�-ݓ�z�ڧ��vO�l��[mܣ�{h�`u(�Ng�/���Tm�7{�p碹��f�2_W_�]mw�]��S�~�/[z��ڱ߬�'���������ґw��	�M�α���I���hEMe�1i�ښ��������)e�i�L�����ѾWۤ�ީ}{�eiZmܳ���2�}R�Ծ�i�}�`�����>uJ_�Ԟ���m��2�'�1����uuOݙ��T�W��Um��6�b���$Q���,Ψ8�pV�������ϝQ�O�����jY�5V�;q�#Bkc�mʤҹ+S'��uOo��d�g}8�i��Ď��]��vȏνmJ�ە�̧���ٺ?�����K;Χo"k�����H��،���:�w�L]-�������6��Rm�����	��p��k�,�"�L��9���ٹ��cROU{Oj�m�ۙN�������ᔂ4���;���j�}{��t���4���9z�z{���#�d��?%���Lh.G��ִ��Jصt�iըZ��U�j���W�qaRU����������-h+#2�87D�T�cV����,즾�����j\+�8��S����L?�_�j�Y�������L�BTL�^}?Jf�?���p�I	�RS�q������LrN{QZ
ڨU
-�,-�XlY�τ��b!��V,R�u%�1�h�Q��`�6�,
�hS�F�L!����j
�\WEZӜa�d\a��D�bG]��JM#XeRZ^��,CGQvv�cVK3EJ�3Йb�*jFI��d��-8i3F��3�i;5(�Q����c,/LM&!U�Pf��5��iU�t�q��5h���	��KuZ���Ը}��:C=3��A��8G��X�)���`�M�dL3��2RfF�5���� 7\;�2uSK!�
�35�SЩ'�-��Ȥa��4�%e������[2�:lR����T+R,����QA	6��rM�8�-�Z2^��u�F��D>CrM�� 1h��+g
[3���� ��c���`�����
�B�aԤN��1i�5 ��5%l�!U,�����f+I�pY:UV��d� ��դ"��<�F��0���T�=B���!j eR
,�F���{��	3]�������p�#�f�/��4�?��i	��df�r�Ff�C�Х,�±l�ќvTG��ʔa�s�⢟
|&�8f�_G�-�8(!�+Ν|N���T��e�Y��zAI2C�%�R`���Ra��L�YO�-�Q"�����5�
WUnk�~눌<#����-�#���hF4^[=Aڮ���;���a*�
�:I3�	�1��f8Ha��PcɡV�hI3�	�K�`���5Bࡄ���i��S�:l�,Y!]8)r�&K`CV�s ���s�!pv�,*�Q��u�%�D�Z���
SB� �Pl\B�©t3Q#~(+2����QT%ie%Ep�����#l� ���@�G����d�ď�
S��}�r*BQ���� ?����/��
D��f�m��%�zA*�?ً�[��2�ѐ�!$�D�u�WLs��-Ij�S�Ȁ"J�&ͬ'`&������	ieRWpFJհ�����B
���l5i#l<p�?1��#�o����#����J�T�RS#��'�/�LeU@&�P)��
�X�!�:�� %�����" �
��Vb��� ݳ^B˥d�8)X�X�65��I��Z�YA�pv��*�d`I3�	I�FXNQܲ$I2��U�b��.K@�*��ȰT�9 "+�T� PJ�u��̀���t.�L@�K���@�Ҵ� ~�9Mr6\~�5��+
lp,����G��'��%���� T`+*�Z$�4��Ф��$.�ȫN&�*
8�#I��	,����}ુȰTdZ�Ì�� ?L¸�[) ɐ��3�(�a�A�ip��H��V*��
�#�z�iد%���� ��R%YCLt ��}	EH�KX&tWQ�$k�Px�	��cA$�L� �Z+S�5�X��d}�!��H�*ʖd:1��=5h�C�ʓA�,@�%�Nё�$�iF����y�`����#V��ɴK�$TkNY�.�X�~U����q 萉#��h>"w���d��"�rJt	�Z�{t��.;"u�jO���T���D�O��FV *�O�dn�#r����B3 �G�)�"'�$@��1%P��3P�! Q�?2�
��"[�O��Td��$�p\;�H��c}G�Gxأ�Saj�'�*f�
�;J�� ����<��Y��)���s��C��!�#(�A��p
����O�FA��%4(��T^�0Q\p��ymyJ��@3:�C��ʃEǌJ#�H�3\��#K&�*�C@�@y
'գ���Q%G���8��)
�K)��UȺ��z��@|��$G�]�隴X�)�c�9���@M�;�D�bl����J�Q����ݒ�N��z�Y� �ȝ�)Յ!��jt�J:�s����z���\�=��
�s��-�ʪ�u��u�Ɋ�%^.
P�Ȑ��@��lV�����U��H��p`V�e��`;Bs��3𫄨1�#"2Uѡz�bUIǸTJ�p�*��%�B�.t�.q�# KE6�(S�(1
et��=FM  Cu�ѐ�QF�� [��������n�j���e%�h0TEN�(��D���YIϸXDRE�<E��Ty�2����ĵ~j����"��k�	�"ѓ��֨p����V����'���)J�kTጂ]jɹ"=�m���ziY�X�pv��:HB�O����/z�Ց��= ���L&$t=!��,�$ǝ+J��{��JW�A��4z�Ւ����A5U�Ȋ�@�&c�Z[u�j)m��RJx/�\�&�^�J���*c!�z��)8i�s�ΩgY=9�$l�l��-vEO�"}EOV 
M  `p�)6ygh>�-z���j+�"3C5-J���P(z�2�)$������2����Kَ�)��D��IO�!������J:DM���<�㔩�yq����Kf�'�������sB�M�`�TV���q�"Gٔfg
��z
Esڒ��3�T�D�<��D��R ?��`$0�����)�d1h�N�e%S��*,H�!6F�KE��6c��kF�T�@Z��3m�꧌j�+{*WA�/��d^su� z��DI�HP�x�rZ��1��P��)K�fܧ��=�)��`C����S�xͨ	�,,%�ZP��8�%b��kF��� ٰ!�jh�=��)��EO�dT�F��~��
�=m�׌�`d\t����J�����4��;�g9���&ݠ}����9���ST��T�E\��8J���x���	R�j���S�'��9/S�BT�4Uށ°>R8z��#1Q�M��(
�ҡ0��)��%̦BO��ω?!9���f���D��y�25S	JNp��r놀!���􌫥�/H�!g�l��	��l���bOh_��+#��1�>�p�Ӗ�٢'e�F�����&+5�)�\^<a�G�r�)�t��bN����B�|J'��\O�Y�����s����X��R���ckj�ag*�իk\-�a]���UޓM�)�R�ؓ1`	R`� �zJ,=W-�ᣭ�5j���r����!z�ꨆ�
�p�`�[)Be���%X3�>� �E=�`���`�4�)��Ien�/�)'�����ߎ�'��ͫ�����!+ˌ+j�)yj�|�C*�a��J�m���TIz��ω4.����gA(�@�
HA>�#�R·��������2ʧ�����e��%���IQ$Ж�
�T?�{ҩ�2L=b���)3�a�4�O�VA�S���gr����N�V�9%e:���}ҜY^z���&<<�����ƞT����fd����5aj9�Tߓ\@�Οsz�F=���Ti�X\&�G#�D�
�)��bX�*��Q�T�2Iq��f���W@ϲK�'qV���3��Sv�S�d���&H���R�$Rh�%�6J��1�v@1�H��(Y"� 41�Y3�Tf�ժ����֖�c�t�$us
�;(]���������ra�R��0K�4e�o�& `���=w������Cʖ��B2*�K�J@�6�Q,�e:��u�A��(_&]Od����C�=�~�Ƣɭ�T�9�aا���~�Cܧ!�F^�Bu��~�qBR#���=�$�2�xi�+�SOBoZ�c�'��8�JC�:z
zʃ���o�������2Y\���M�ϻ;ip���৮��,�_8��v����V?{e�ذ�pe�U��Sm^��4���Xm�	g]m�7#z���fd���.�[m�"(k�A���DS�=m��F�"a�yZH_׬y�Ϛ7ܷs����K�������4V���y��S�,�$)J.I�u������:$����AqG���#/�3.")�P�D��I�+%���N��4���s���
G�	N�@{T�s�tBrOr�kQ�J1����s^ʋdn~�����
�bD�Vѣ=ת�ԅ'��V���xΖjp�j`&6_��*��Z������"���ka'Y�*nf�"�"0:��VpOJ@��D���/-!�[9���9��y^F����[%�Q �bgN���
Z���I���\Ⓔ�`)���)=�w�6�.<���� :�|\I7Y�٠T�I	[�I��+�N�X����ړ8,��"E�o|7x���D�|�*?�j���y��X$j�K?���ڦ�T ��lVӅ�ub�7D7И�$���f<�p�p�g�y23~9\J!�s��µ
�$�=��S�R�x�SʜA�p2�d"��#1i.������nk��ʲ|\K��/�.�z��T�oSЅ��
�ΜB���B+s�c���ɒWZ��߬ĺI�s^����z�/!g�w���*I7hB7�p��(�V�a�He��F��ש�k�0]�y��m>?�N��4s�3��k	F���.ʵ���y��qG���V!1H���ޜ��W9���Q+F�{iSF`,�y/Xn0^x������x9�/�ca��=���n�:�vG�cR��0׹�g�:�
Я }���0t�����$l"�֑����l�6��e��4��5S�,r7��Z�7D�L�)�dΫ�a$>�d*�'�]�mf-B��L�3�M��.=��/c�K�&+H�ϋ��x^�_�r�&����l7'�<�t�U'j��f���%��$+t{>��M3o��OrxaO^f��r��d e�I��k�BԊ���$�?OJr0�7Y��t�/Ge��h�yU~+��;Ox�б�e� �I��#@��ņ�lP�p�Z��D������o5�ҁ޺q �Q:^2/�?A'�����ij�>��0A�#��:��n;�1m:'S�f�(����"g�	��Xa�] ��q�EC��	`�	�؏_o�����If�m"�k���aTު�WO($}�$'�.��-��3���������8�u�3H�K�B��a�o���/���ɃLM�g,wQ��4~�Ț�' �q�g�P��R+�R�Y|B ò�/����@�ԏ���U2���LN"��2�!L�j�w S�!�x�͡�k� ���]�yE^|u��e�daoPz�=�.>��$P���nd����=����l` 8�,�Fn���G�v2���x^�q�IN7��@��|�:����d�ې->g��'�I��Har��a-�Rxs�Vi<o�a�+�d�H���[`�z��-H�M����c136gl�'�"����[��`-�����#�!P��=��x�����_$���Ъ����pd_ގ![�Bk��"���iV�<dV�E�0�
�ړByA��>�GC2l��ܜ�{��E�s8�c؈ិ�0��O���!����GC��k���M
?n�04��K�PoZ����f��H*>y��`�ګ'��29�,�y���/eY�J!9%�~o�P�	�H��i��e�-0�A�0�)��4��F���JA$���Y�0T^���#��~�Aw"��,�E"S������p�I�V@�A�HLe�-0�x#�=�@�H��+"��4�_����$�3������37)������r��P����W��7b,�y�J��.�n ��[`�6`9څ�d�������i*����,ƍ:���d:�Zd1|�����0BF��y#�A�-����@���SD!)�*(y�D�`��FP����@*�㱈F�-9�)����*�Ǎ�4�)��$f���>�C]�����y���)�T��h�~����j�L鲤�!1�T��k�8)a��"���y���. �O�мJ*��]H���-0����"􄳠����-0��"����SD#�"���ҝQ��"bZNx��J��""��r���R7�������z'&`!AS��z#��r���	��� #��/���,N�
=��~��s�Ҳ�MK�d�0���Cf�WK*$�� #���jH�}�L�/�Kd�0���AKp���31ր�AjH:{�[`���*{B�r��R�0��a<�3_��HB
~op�*�@�e<o�a$��F�,'1���X1i�L)
^���[`L�y�	Rz�̥����'Œ�����,"��x�R���I�"����t ���T���LF#I~i<��`,�C�0p�<,�"��Y�k��;��6Hﱲ�Fҧ�M ����RF#��&�Oh�$}3�?��a�jø��ae��?n�0ha\"�{�#���g2b���1-H�nR�5D�V�C7(�_}���E�0�B� �����qHE#)��k�\�Ӵ�ۙ�-0��)�@�l^�r��Ak_@%!�c�`�*bEϗ�'e��L�����n�R�|�PT�����0h�60���E�M��ME�V�����+�:��-0��}�I�;�4��51�b�� ��5D覥�U��a��7��>��e�����>��ɂ�`��1�B���Kc{Ni��g*bzt��>e��L�:��F�"�*�~\A���Qݽ����Wi�㨈a�-~oT,���|�FQ�xeȥ������Q�� j>�(����,bE�H��sR�1��;�Y`>�S����(x#���>��ی۵>�@zg�7R�V�|#�Q�t�,I��cU�0вP��Y e�A��a �{U�wiC�JE�H�K��}8Pp+���#����>	�rU�>���t�0��B�V�sR��L�y��r�kH�L���mSGC�"�����ߟ��Fõ����z����!u�0:+�6�����I1�~H�z��`��T1��;<�Sa�_���#����T��9Ĝ����u�0�2_/!��S��a4� (*Vx����5D��t`0�q6Sޟ�a�ǽ�k,� ǥ��D���xՀ�Ɋ���"��{>��d*���U8ވa0��,Aѧu�?��a0����3�� ���[t�0�By��]�$=/�y#��)T�U��G�
�at�0`�M�&?��K�9o�0�"�IMR�:�,1��>k�;�wC��"��/T�PBC�܌�>���8P��k��	��� S�����G6��1�h���n��Ve|2àU���7_��{)a�à5�=M�DњW�+���*�ޢ�L��u�DC���Az������0�����k�`��M�0Ԛ^���'��x�DC��Гh�a���k��Z}�0t��OAy��Y�0����!p, ��#��a�+���+�7CUO���a�*}ܐ���5h1��ų�����F��̃S8
���{�4�CX/�C~
X��C&b0��y@=V����a�|B,Sa\j
&b�T�wW�N^�4��Fc���npaǀL���a�P(}8!���-0}����@�#$=��5&1���VNJ���31�=���N��!rx�c"�C(�������5G12;�i�1�p��ڲg���..J�ڕ���z��Ga����0`�a�t[=o�Y�-0�!ǔy�,�P=�l�7b��1 �I�5�וm�0��(/t��>I_��ㅍ(����R-�J����0H+C�e�{��l�.�y����=��Ґ��`�٢��RӰy�_}0���FC��s!�����6b�!�����	�[`K_n�7ρB�l��x�EC��}������Nů7b�d�+D���c���0�*�ab@5/_��?o���	�Dz�˼��xc�K7�
����'m�0��f �T�����:��o� MW���0���P��ǥo2��1���p�A|p<���gB7��AJ؈a���8����89����a��o���{:�H��F9o�a,=D����@��g��ۻh-��ņV�R�x�;I����Qť�   	pHYs  %  %IR$�   �eXIfII*     (           >       F   i�    N       %     %      �    �  �    �  ��    x       ASCII   Screenshot��W(  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:exif="http://ns.adobe.com/exif/1.0/">
         <exif:PixelYDimension>650</exif:PixelYDimension>
         <exif:PixelXDimension>700</exif:PixelXDimension>
         <exif:UserComment>Screenshot</exif:UserComment>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
��^  ��IDATx����,Gr&�Y���F` r��!�<�l����������5;�r�C�� 1�������U��BdeV�� �� �uwefdH�Ͽ��hY���]�6�d����K���|s���r*F�l��镏�	�Q�}�o�$�{��ߧ����n2��m��n�c��ߞ�+,��Nz֜�D�|ߧ������}�>}��Oߧ�F�� /�HƸ&�*\7
7��|Z#O~��I�YK/0��S<����!�� �_ן����o\��}��X��2T�,\�k��.3Y�x���3|Ԗ���-����;�[���n��5g��H��ga��dx�}m��Ar��.����l�'�}��Tm3^t�O%�{}i�o������ﾾd���iE��-ɣu)icm��+�:]Q�]�s� �\�6������O��e��y"W"�X��ԍ�S�@~F��+#QWI+�`����4��yE��������D:���fSY�?n#���:/���'�0�F��8�l�:��g}��3avi�A<�O�.e�g�����w���7 x�*��Y#`�7��~��B	�_�5<�5UY���+(�oE� 2�l �$�Jea3���D��O5�ʧ��r-*g�֗��h�z��R����k��IB7o�alC]&-5��/F y��AK�8�-�O�A��Y�Y��A�0���W�N�����Ǔ8.C%��k4 �
���}hL~N�����k!���,�%��sz����ad��Xk�k��a�g:�F��J��2�X2Ɯ^Q��6=��},�3H���`�@c3P�G�H�`����x�68�4?	��9����O�v�E�3;aMl��E=����R����ƌ���|��	_E����)ɧ�@��1��~,�T����J�Ӑ�u�A�˃�A2��s��[g[7j�i�.[-G����^��1�$�M������,�^�ؗ�c�WS:E�����dD�O���(�̐���Y�
7>3?������1���	eC��Y׎JĜFx#�e�/��5��^�e7�o��Z�@�4;0M ԟ���%���}]
����`��F��S�"�&C��*M���R�+x+��"�nPa��2��;���^:���-h�Z��ޒ�Yݯ��\i�5������I�@*�ˢҶ�ߥ�7�7BL�&�lu3�F�a�_d�҂�&��L�\�Ψj�+(RF��1�����J-���>�
̖�N5:@���j"R@��S�-�x�[;�e���<nQ�iaUH���@���)�2���tw&�X��������h�KM~�I�*����0����r�&%�%u�#̸
e�@��Ku����L���B��kC�>�O���o(a����]�ט��M�V�F)��؏��~��������7I�,E����9O2{LVY��<)�	x�T���(��{�rN��y��dy�N�诘Б�r�}��*��Yr^��L��L:��;�N�0&?�XK���`�:��n亰�V&ד��$iQ8,��@�V��Hޟ�"���V�ɲ ��#'�-'��k!�C@�^��4^j��aHt!�Q yrdQ�ҕ`BGE)e����8<�vm��v%Q��ǭ����wϞ��f�Z�9�h=H�(�D�U��н��Q�")F(��0a8���>�`p��SG��"v�bTrgZf
ʬF���b�)+x���G�m��Ԙu��`vn�gf`zj
z~�]~O�Z��u`��l��I ��(B��*����A�I��)`� b�(�1b���p{�1j���1�@K��EB�@���+J�x�)}�V�b�Ҩ�&U%T�֥㸬��4X�x�B�}9H���@Mb Q��k�+)�O�x��H���)��eb0��ȧ�\��6���T~3�J�"��z����'*����K_;<�R`�Ō��B}�N�ƒd�.�*�~�[���=�>��e���B^,U e��`�Fˠ��~kM<^�%ri����_��aΗ���2��l@��f)ER5�-����j�2����;h��Xv���6��Ѹ�"S����J���)�$/���^��������%���*O��)uy���w֑��v�Խ��?�=�Me�/wƘ���
Wo]�L�O�?~T�7�~��)��\l#���d���+�ј@�u��#ճL���qKm�8���沢cT6�.��N�s���k��E
�ulb��虜v��v�����C��v�-���9����1��j�n��	���'�8P�YS;(M�ԗ7���#Vw�������&<z����'�accv��`��Ё�C|��5�H
�'(��K~T�&�V��y��H5
測<VrD3���g�������R�7.Xb�= 	�1#��J��'��J��x��-	�1@�����@d��k�dG�SީJM�W?�OY�BiP^Z��X��C�0�yy<6��V�=�*�J"�Om��O^�F20S����:��bEc��)�,c���*�<���b��2�V x9�Y�OƏ�: n|{����ԩE�'��5o�������'�WW^�0fE13�b��&�X�GW�������S����ǰm;�����,��{Y�mJ�r��V.�} L���yVoi�bf�Բ@M${h�T��]�
)N�{:�T�`��5��llEu���H���K�Ȁey��wr��{�\5������r����i.��F���	�FLk�r��k
��X`pSz٬�%o1�C�P_��x��^_ed\�{�"�SB:�r����O�o��i$������񧲡�P�r���v��{��a���C�W[󉌑���:�&��-c��wb�ᅼ�6��qP�T���H��3sї�ѐ�5�o��_(����♉�ṫzZ��|��r/��͕H���{� ��S�S��,1d�N���鞙����yX\\���p��:,--�w�Y���]�Wg6��I�z̈́k�L� oH�f�B��HXj�%�ZZ8i�#8::p ցٽ�z��?{ϟ<���Ã���[[�������D1��<�r�:�(9��C8�P�v�*����Ec �l$hZo-�����n�}������n���2����C��L�G��X�U /���YX���;����`���xOc;q=3�:�dy)�����J�L����x����슭/���z�"���	���U��N��<�JU������;��װ5N�W�nnp��^�����i��oǱ�Fʩ�(��[	6z6�ň��?��z�V5��ܧ��JN���
�(7�>�c��j�dC����o�d�q{��mV�Em� j-T_���X)��cw�\�;�J��	���\�q�*aeV�I�N,Q���b��D 4�*;M�W�A�;��k�Wѵ����1��m�����Q��eGIlwu'�~� �IU�gTLۉ�]_ΘV�WWKVFF��҅eld����~��1mc0$Gp�!C��	��Օ"��ȍ2�<b�"�9
��b�ȯ�u��"g���5l4�jL�ۑ{�Fɶ 2���j82��|y�R0ȭo/��܏d7Un�dE8ii��5n�rԐ(������ڞ�TRy�{Y��`=YB}*$	�nc?���=Q@$WQ��.�ǃc?>��LOO�����������,���
����w�g`jZH:�FU3��ߒ��TC	 Fz��¢g3PG�����x���w�����K��.}����@�2����!1pE�>��1y�>lU����:#�h]'���	ᗰ�!U �V�7S�)���!�I:	s7H����;^XsYdI�XQ�Y`X��:�	��\���x9S�	��.�`F�2���^�H5Zni�%)�X�*�P
���
_U2�D�m�Jm9Á>,�c����k
ǟa�V�N¬"um�����X[d�I���6�]�̌���B�zν3��P(U�E=^�R��� �UX�.
]�ä��2(�ߡ؅1���۳1y�,�^,?�vi����	�x� 6��0��ϕ"��]��'\עd��kM)�m��ev�^:��oP6�ǫ��jjo��2*Ac������Js��Yx���x�*�5��Șvb�1(n�!m*��b4��ܻ)�-"�UY�jBcm0y��Z��)�����2���v���S]S�ʎ�Z��*Ӄ<f�'2��[�"�GV��JY�"8}���c�<F\{G�$�S���`�w;����X�C��o���W��D6S���[�f؀�"�͜�i[^��.���O���(�`@���Q0(01k�P�>O�  ���<��*�w��e���`������ ��.�2��(Ï���x��su�	��$֏A���f�[��Q��M�L:2�x/���<�f���	��]8�/�V��|vHF�h�{��4�F����`{{>���������%��p���z�ܸy.]�L 9su�zBv|��k�&�����d�դh���,�����������ށ��-�x��߿w�|Ϟ>�/�;[[����:��,B�L<�\���.]�Tx80�u��D��E��gD�ui���;@��	T��Y����H�B.��(sͻL��$ �'s���"�#9��V��TYa r� ��7����.(H$oR�\�`֛KN����g\F�B��h��}dFM��N3a��S��OC�m�L�H��ovS�	^!zV�Z�?Fm��H�8:�)����Z�V�U��ra�l�� �����+����g3B��sA���F������./�<@5�l9�1�hxY��J&���֡ȨAK�g�X��2�g2H�VXp]�wUib:U�d��lܜ��3�v7�2G�*�2��9ӲFmА��tW��cq�.5�P&�9y��|�g�Yd>Q�dܷ�;�rkt؎�I��.G��4�t�zZ��Ge���h��Vb4d$r���<�)�^S�8�q���*]�ou���9��dq�@Z9aC�6��4����eC������H�lF���m��%�Wow�������z�}Au���ߙ	D@�F�/�~5��khf�}�_)�����(��d�{Y,B�g�ZV���֜�U���P.u����]�s��je)}�{�t ������e�uC*�֌�mVd��׻����z?@�o4ywf�N�Ḏk/]�����K��@�@f���J�h	� ��vƮ%C�>az��q_鲲�!�L�WÆW@�����~���П�����.�t(ˎ;�������{�,��L�j]��0xV����s`���]�p��=����`uu`yyV��a~~��&�!�c|�#i�7�ΦnE__��o��R _�0d��`�i�ht/6^��O���{p��=������m���Wpx�G�� ��X���B_#ƌ8񽰕����|��3hȎM��rѪ�Mo���^��6�D�������X'�CgE�s��C���xyA7!0C���f�@��8O��Pb!�Q����Z�G�NX'4�����huW'+'��Q�r@Z�}��hWo�ꡀ��D	������ ��U��| ��Y�1#��A�2%�*�z�0q����0y����	�`�Q�)/�`rw�<�	�e��+��o��� �N�ڔ/	rϺ��@�P�!bհl#�ލ�֗SAe. ���ĭe0<�,G��ƠT�@j3�W��>��і��N��"j�Sц�0��������V֦��>�`�/�Y��տ�����*@���@���Kr1l����u�W]!"�Y�b�>�����Z��?�aV�,kz��8Л(?�_�hN��S��0r��g�s��V\���vb0$�T��]�2�ڠnl���i�Lq�uH���ep��a�������L�+YY�z�/��
a�Ș�w�a���A7���Y�.���܌���|&�m�v�h�KhJ�ͺ�m���V��M cv���ۚ i���Y��i|��TCˆ�� ���3�̑�
�5H�e�Է��*`�Q��VX�4�r�3���ќ�f3݃��|fe��H t�����+~ekTR���W�ߧ���G�Ӗ~G��ƶ��膿�=�va&Z��F��K3��s�-3���}� X����Lx���C����܃Z5T�khV%*�M�v�o��>��^�2r�#��<�Z���K�����孑�m������o܄7��sb}��ew��k�_��Y�>����i�K��?,Y���@P��s�
�i:����܅/�����6ܹ}�?}欌m�	������[t/�N��..��@�w�g������q���h`�r�,Ic�ڴ�3 ROX����#����p�@Fy@���%�cw��F�$+!͈�%��C��`G|([�y�ftcSƜv� � ,YiEԛ�%�6��)�����RPݙ��V���`��Y]hM���%�
�G�(���n#��X.uu��D@��$����
U}w��ū�jٳ�U�D�u)���G��cW����+�'b�_t��x�T��B��H����L̡G%� �x�E�C��+�cĄ�m/�v�M��{����n�ԕ
�'[���oC6�(��=U�Fƚ�me�ǒ���[ʵ̰e#QA�D�*df���b��M�mm2�eHKÚ��w���+^�	؎���65c��k����5xC�.�򥚃���d�m�jP|62Ό�J(o�˦� ��32V�|r?����	��& �d#��� �k��GE�"+ �Z%Ɍ\Vh쏘	�$��LY,$�P+��F��h��̀\�l�������<���Y���e��-y���R�
e0�{٧ �6���}l��*��l6:�g�a�(�aa��B2��@(�O0?�#�Ap��"��6~��(��2��Ѫ�|ϫ��x]eT�8Ӿ숁�׼Q@nX�o��6�.p!<B�p�re��wdQ��o��qO����kf���g�%�d�r2D�>�;����އ/����\���o�͛7���+���L�8���_ki�9x�+ΠЉ�;�d!38���.lmn�}v?��Sx�����W����G���	G�0<b����mg�8P۟�Pg��S~����4YL�^�����N�D��Z-���	_6�c
g6p��p?�=��|����}�����3�F +|���ўb胘w@�f�d3V+g_��[BX��Y<�x�f�Z�C��ӑ�C$0%.���]�NKo�ƍ�0vaSB!��ay(��;��z_�fA�BA!�O~�hՊ�Uل%|'9�o�%���3WĊA17HC#²��<�x#7�H�kya`��-fFԗJA4>BG��+1�._����z��w�+�R)��}�k60�;\3Ġ`�xcF�"��"R5����'J9�d�Z�<~X	'e����8��x9"pcLs%��M���4D��XA����X��d�w� �ī��]�(i�y�/'�G�+rS���������|�"�DY�M7�鳥tY�BZ��[�Q*�>5I��4��V�}�ay��g[�V��ZB����P����1�C[
DZ��Mm���x�xۉ+�2� 6��ǭ�!�β�nc-��x�;��	�H��F����'W�Ck4�*ƃk��a	�T75b�h5J�d^*��{�2���>�2�Qp���M�*[�EϤ/��R}�rYχ�3j�K���WSTfYӪS��t_�Ob��X'!���d�-u��(�Ql_9I~���܂cY->r���2T�֗ƅQ��uJ!�F��F��A���� ^^�e��+�E�wX	�5�#��������=��]x��9lnm��'Oac��}�^�J�wfv�C�u���������� o��x�D�8�q�2��`@��~�|��'���ݻ�]#>�x��P�<n$�t�r�r v�Y����p_}��?	���1������+�.�3J�5 K�h4�����������6�x��:��c{� �ݝ]�C�F|Ps^Vd��v-p,�dk�P��NX#�3-y�g�x�%�idx9\Y`_d	�U�J�	,�R��
B9��T�ͬd�)�YR��Ki��>ʜKƓv��Ň���
�CQt����^Q�	�Δ�WI���
x�!���jg��H��1K��&K�H[���E�k�}o������ӫl��５i��m݆g�AɓR���i��a`��/0n")=�3��,�b�q�I����-C��I,�p.�=^9F˃OzF� M�ƞ�:���@�̰�im��by(:~wR��%_h1z�]ӕ��F�����f��֔��7�Ɣ�e1��e^[��{��v��ɇ�D���7h�&�]�^�#c�2m[-?����nU��$T@��A%]�r<�t��*1׉���tU��a�@�W���)b2��:�s^��!p�J#[CusJ.F�uX���z M�-X��E����*�]�x_Q8�~,񗃡 E�]�lS���:�w�g��u�b4��9��'0
����2FT*Ġ���D�Z�>tN(h��-�~Z!��[��,�聀��������2SлPk9������7�F/�A ��ƓݤZ^��Q��n��,���xD���24H����P�ū{����ySD�t�+s�f@�u�Y���<Զ<�SbIWS��@��O]V��B�J�Tq��,,�����`gw������)��_��׮��#�v���{]�9#�q"hl���*���
K����$Nf�)s�&�������;�����࣏>�Ͽ���>���&�(Cl�N�K��g��`nv`f-���Ӱ�0���0��@0�]
�~G���l�_[H�
�r��d�%�L,E7��%_�q!��C�{���[��8Ћ�w�Ŗ���`cc67�=:�0j�
���,d��\;d�`�!�թ,t�Z)��>(l�]��,uBLKc�q`��j��uǿ2��H� ����2y���acU4d����$f��XaٮV��L����.��T%�iF�M(�E��
��$�P|��\*�PX�ů Ã+;��%f|l0@�.F�:@ĸ�OmK� N8�H���gd��)�Q�L�� ><7��[d�?<�d��
�ɰA�@�6� �c�ɓ�!k��U��Ҧn9i��	y슒�0`���Rlqţ�J@�0�B:���
�;����_�N6�F�%�~�}�2?�4�%���"�G�(��e,j=�,4��Hwk�}#���ħm��.���	&}���̃��^��zC�x����%#���H��o@S�V�ص���o���,���5v� �@��Y������L�.�K�EV�T%�
hl�4F-����8s
���bX�Q��}�7�Ʈ>����$�#;*��Yq����iv-��^�ɑXp�EQ&o����d4_��� �+�G�W���d��g��a�g�|PpPf�J���n�A���ɟ�|h[��h�G�r��ْ���l]1��o*���>��@�%+�~�,�ʢ�SШ6��`z^O�!3�ǧ��J�Qx�m����/`�Ϥ���<�����Ճ���R�����9����3xp�\�v�_��R/��&}:a'�v��r.1�����R~�I�=ڇ������[��Gx�x�76��u�7�pT@>7�;=�,��XZ�s7��05Ն�i�1�:'���҂k�E���	��.��u��сC��|U4\Y$+�&�	��F'��D�0�R8�������<s�����Sx������+���C��-Y1���(-���)�T��o!(o�Mu(P���K9 3Z�0�2R�q�N��^���2J������b6u�P����A��y�0T�R�	y^�\�2��22֊;���,��0�i<j0��Y*S"��b���/q�(:r�τ���d�]C���KK|���l?Ux@e��l�Q���n���ns�$�a�Շ��x���
$�7���n�X�Z��Q�,[a~ː��d�D ��r�ft<���c]R����IX�y�����p���cd����ě**o;Ej�U��+3F�#ـ�>�M1s3�H�:����x�uF ���0~p�,�l��I��J[ ��@�89�qB��伃n��X�Eㆾ0�x7�7,%�g�-��p`�A��DsÊ��M�)���h�X�8x?�|�󴌎�_ąn4�w���~c��6��/S}���1|��i5J�%2Fx�;�0����pH�h�_0��+�g7)��� bZ"�\�W�q����`,���n� ��W\�+h��l�~��_N?�I�ng&+�¼�S}M�#	+G�$cىl�nBϺ�_��f�����]���.]��7���N9�8�E���c)��:��" 6�D(��??��
���9�y���d��đ��t� �8�9�᝝��C)s����f�aٞ=��߃��{����?����'o���S��^z�NK��R�W��bzy^�l)7v����<cf?���������>��?��� O ��$�������unv�g��C@;�,�Yx�g0�i���ޛ�C�X�.mT#�.�1�.�d��!\:.��,���,�� �@�,�� ��Ŋ?Z��K쀹���6���K��p��E��؆��6��� ���'����x�A�G�G���̀Lc��|o�Ś{��y� B����ju��3��g��@b҄!@U���J=Ï
����!$�:U:	u�HA�A�U��������"�>a%��B�C�/N"���A�Q�	�X�����v�A1�Ɍ�
�t�Xa<���ZA�B:�+�yn6~ ~�e�K����ՙWt�J]Ã�#� x�ۏ���V�|,��Ae�Pu܎�,���uɂ�f�f���uUP#��+���7�W���Z#��w&�E�J
���7�\�W�l<h,ٸ����o��Ё�s���㕜e�����x�~���e�K�k�aߞ [?^C;�'>(l�o�Д�!Dr�㴤��U/�c���;i�@�i��.��'� x�x���p��!2�Rp�k^½�v1�`���O��=�Ȃ����>���±��6�����(���ҿ�z��~!�hՠ��ˆ��8��hD���h�Yխ ���v0��'�j�|��M����������|o���$ڿ�hl�AR��p���(: �Qy�s7�2:A��р�����1�r��H��Am��c8�yØ��ZO��,�$+ϐ�UƋ�!#����"��=K�ƀ�/��.//��n�=X[_��,;<|�����p��M�y�����_���J+⾓y���y�����������Q�<m�ݹ�~�	�˿�>��c:8����C����wdnv
V��`}u	���aс]�9����sq���BK PrP��^
��;M7D愅?�a�)%F Zǖ}����m�y��/�&�<h!CQ���uZ��~.s4�Ѕa�|�8�{��{�՗w���'��a6�����0$���\@��`V�(�4�R'�#1uU��0��F��El-�L'R&�g%_K��YT����BNe�nC�$cBPpӓe>���M��e�;���kF�ݗ(PA w+���̨�"�JY��+���DUf�G_(�_�N�+�����%7��-���k��eL��הU��S��>�r�	�P�,�6����*���`7�p�t�+��)��ՍMU��A��|:���IBU�l(`�� �z�!y��ZVZZ�P'��0��fI-@�Q��[gq\V�6�?� �8�|�H�gOx�����0?p�6�Ն������M�[�ؗ���d���>����潵�IdE�lj�_�I�0aޅ�!k���V�Qp�RP^��dh�(nA�OQ�!�������LO�IX��ۃ�J���xf�Y:D��eƿ�Z��&+�_����|�wl�Od���X�I0����Y�!��A!���^v�1����~ѐ����7<��'�;
'���X�jX����πD
`�		�zɃ^1de����?^E6��08.�F=�����@�s��Ns�w�/U<7Ϟ='roc�9<|p߁��� �ua�,,,�>�p�r��E��h���Y@��g�t@�&ZuH�g̮�� ?�}�>���[���;���U|�v�R���Me�3S��4�,��ps��0Gn�+��EX\���i�r`��mS�d���FG�/Y�R'1�n����2��l���������m�.�$�sb���;<5�ٌ��0��,���W����p�	��.���aɁ�W/�?�<��������A��9<�E~�#<)�eߦ3�[����އNT�Nt���%���v���U����Nbk� �ɚ#�EDK�F��?Y-z���BN��B�D(�i�f�	B��Y�@Ձ�S�[R���'o��32V��[u��'U�K\7�w�1fߵ�����@Ϥ:T�7v-��%������Y��&�@z�4��QO�.�##���&�[a�`��e���p�M�<��o�dh�`� �3h��!�R���������-,@�2)��|̺�`7��U�<.N~ߞGY�>`cCX}jcCd�qR��X���f���~%�$簤М���Z;a>�����A�˸���S�AL$o:v�)��"��L���+�1�B&�ӕ!�G!��$�D.>�Vò�<��X�'K"�-y��_u��O�ku�d}� �W!�	�j��p�&���m��ۅǏ��6<�meu��˛�ݠ: 3|�0����>��#x����|�x�?���y��?n}�U^m:=��f��G��q��O���}��>|��?�[��w?���c8�'��`N!�0z���k�EtW�]�#�	�..�����.�L���G��p�V؀���V�Db�la�h��� �Pȡ ��"E�����p2[�4��L����S�����,��%d�j���g�;�<;݁����勫tf��˗���p��C�{�!�pF��� �.)^!����M��N�9A��N�?I�	�$��?�2"Ь�T�'K������|5���*����}u �c^�$�@Rk'�]]�b��"�H����WoOۢ
z�yFP���9I�|�I�G��,� �.������ʜ�w',+b�qkHi~�e�������_�{�	��o�hC��L��5\f�Vuaa����u��p1jt�מ�>c�ԁ]��U ^��w�:�<�M1�����ߒb�kT�PXKrR0n�+6j�F{��/�N�3����[rsU�N��3��K��pTnm���% TH��0��oI��}�x���-+�k�ɹ 	W03kZF�p�\����͍��́79�jMQ&����V?��K*��؈�4�Zc�=�ݕ�T������܊�St���n����C��m���\�vVWנ��c��06�l�穇Gu�﫻���o`I��a�P	<�w������_��~�}�°����N?�o�Ȯ���]]���پk�%�r��kz�ajf�N��h�� 8���xpEYpx�p�H�%���N�Q!������1�x��'���=�GJ����6ag{��=���]; ��ʶy�ű-�2�t~��T|2@|��wz˰��
����p������(�>��s��S0��C����Sٸ�Y�ZÛ���3 ���i��:��g�~W��0�>a�I����*[��`��h7�. ��x�l$���9R�~f9o)���i��˲������I�I�����0s����i*����	�&�1Tk�30a�C�eƮ2�l
�G
��;]*��7�ed����b-:3�ɇ���y&ʚ7��B)�I�S�(�$������$o���y�@5�\'�#3y�N름@��Z�b̥rՎ�O%$.����L��z�YI��'���Y���1�3�7���b@%���4�m��G��1k3�F����y���[~��EH�>�"r�P�uN��GX�o�x\��B������قg�ٍO7o�1D[�%w���zO�=�Օ�r�a�U���a߁�G����_��;_�_��/�?�����[��� թFI�3�$i��d��7AH���@	��(>�w��;x��?��� n߹�/�R���i��[ ݹ�.,-8��؇]����Hk˰vqf(r�YZI ��{݀7��0/�ƾ-�yK̲��pXRL=�����߲]tW��Aoj�\2	 =��{ۛ����6����hg�g�������df��Q�`�Ů(}�u�O9���X^����aݵí/���O)���H��4w� ?���h�5v㘰����Q��M���D�U�~�[�F�yDc�}�e����ZN)�u�.��l
b�x��Ż;<@��|�-�Bk���}wZ&d���IJ�,���I˕�:c��D���m�t�A|�N��\���ś y���p�Z/��m�f�7�T�hNe|q�&9uσ�dc.�X�Z���a�i�X�1�E�[ꕴ�����a�/ƈ(V���M�MJ����3� \���S�BZ�p�Fډn�&>�ŔU/k����VL4@��R��`��I�M�Z)�M�qx�~6��+尊�T�'<�ʥW��UZ���JC`�lLrs왭@ӿU�w��PF��e�az�S�'!B�i-��� ��&5IWue�}�?G�{@����+9`����-�	}t|[K��,���,�'C̶��<�b�;��ߧ�����azf�ݾ/��Pn���}�v9�ɥa��&!���lm��/>�_����_��w���8�="���@.n@�v���b�>�̴an��kK�~a.\� ��[�'֯� �#l���S9�2�~C:Qh#*7���B�OLÍ]9pCY鬉yX�[���+0?�y�C~�\K��Ӈ_�����[ﻼ��\�V�ё�
��i�ۇ�.=�������s��1��x��,,�`a�*�|�2���W�G����+�p��c��A`wc�˓<������K�c�h���:GߕA���"7��u�q���q���awu	bm�x�T )���9���BY���.���4+�o�%UP�M��'��4@(���'E�ƌS�Q�.oc�Q����Օ�B���o��t��0^Y�V7Uƪ(��?�����%�~�\�ÆYL��%�<H''љ���tꖜJ	�SJ����$~l�ܱ:��DuJ��UF�	|~��3u�[�c�Z'�U��Gl!%l�v��
�9���~����%@pX߄pq����Ad��W Ӽ"��7���9[Nr:k�7~7>�Y�D�ԍ��I�#Z}�۠ڎP�K��AoK�m_<�͟�'cχY3�b��4��d~u�:Ty��iIY��a�LR�0��V�y'��٣�]r�|��)l��^�	�?Z���n�����w��އ�?����L�{^�8��H�qxX�/�l�L���o�C|��waɚb�Iȱ��]��z��ͯ	�~�ѧ��l��!��0t��++p��*\t���o+F_X]^���`e}�槡��Љ"d)�0q�
���)YHlX�00�V��xK�	�H�Q���Ȟ��3�ߛ���+%jyZ���7�ᾑ��簽���c�P�'���V�x������>
���xr��ȧ���@����,���S�p��x�����ný;�8Bc���o��@�8�x�2oe��A����X��{��G*Vj�~�cY����o����E����/���w�81�<w�>�ƍ����!�c,��*���r|i�e�B��I. �:51��o&�P<%����?����ޜbu�)1�'?2<���H��>��gxǣ,�����qwƝļ�x���8�����_���p;�M

cS��,�SO���)�SН���O�	�4�K���qYՇ�vm3'.o�R]gfg`nn�6��)VX>�|Hu���wm�#����t��!Gp/���������4�xu�i������iMU��(_<A
ˁyjL�8RA��Ӥ*c?��{�����a��'�� �+��#}���r¨�o��F(�8��!�ģDB|@�-����8��{�R&�7)���]y
]���aC��؀�8�	���i�䪜lZS�J�LyB���8�<6j_ߵ�R��%�?��h!�$:�3��,�o�����2�P��D�C�*|��1�>Q���\Q^%k`=�Y�7,�h��,X9�#�X�XY��Ɂ[����%�z�2��/�O�|>|�n}���/�O>����/�?����?�ٹ9�:�)��졊����a����}��;�6K�?�a=<܇�O§�|���o�W���oo��)�N/��)�[�v`w^��L~����)���X�p���1Ęick��B9B_]va �� $�qK!v�j_���%��)��:�dzN�8e3�����	�_��pP9p93��̝y��<z�	x�Ɛ��n��A�M�#Ċ��.�r��#���@k��f;NH�p�KxZܜ3.��M��t�X�gϷ���a�˒$uWD��M���ܯ[O��Ϣs$�fA&��@0�pEO�Y���B�����x9��qc�Q@}�N�X��$Lm�nAy��k����%�:�+�����g��e�Ӕ���	�Py>�=�������z 0�-:�C�?x߳g�(\�Qt�<�'��C��ދ�W}z�R,o�'~f�hM�Xw��F���.�tn<��YZ^"A�e�wc��w2���#����%`9�:�n����X!�Xn9�re`�G��ɍ.���=�q��X���K����Q�M����6�0�>���+_T�j}�\�
�/_ruX�=z�(F<]rgw��"���x�����Xl�E�;�G����`�ٱ��qp�U�Z��s�X����(ʢ����9�'�Ռs���k�Wѡ2����W�/$��.H�1'Ĵ�A8y��y�`0��z�~q����d�x�K�6J?DfP=�r��j�]�9��b|k)'��}Ta�K9e/�\���<J���S�_�2�u�TA����3�?�,S��Dĕ1�+WT&=�4�&�k�s�������m',ܸ����xý����/���m���"�w��k��~���4Dj��Wv�甦f�Ö`���o$X�-�� ��;o�����G�����œ��c�u`wv~�	�U��/���,,��`ǈsp��XXY���:1�a�gn���eׅ�ttE0#Ο,���@$4"�;�����?k2'���8 �Gs�? 'Q	FA�W�ՅnW�Q�Ї��(T6Aa�\� �$����=���H6�ɩtx�
n�����9��,ӑɿ�����9����`'׋� �V��-�[?pýM`�:\N��	t�� �2��iZn��UӪ ���$ƠZ�Il?\���ؤ�����eu���6�������i������"PR�va�Ϳ�E:��h쪠B_�0;Z�Q����X��6YX�O{C�R����wa6K��X�t<�&�N�MGr�;8#H?�=��<��m�U�Ӛ2RhX1���}&w`js�++d�1�z�´2�:" �4D�3�:�u@��@.���
�'MM�H�!;�!��_�t	V��A�wwo��H+I.ۨ��L����MSf\�(0��|�"(F?=�e��2NN36'���4i<7_2	�����0n�c����b�)v5zU��w)���o`���J���	h��Z��!k�&O�����* ��U�����F���,�� Ǫ�
Ī��5J�'�ɻ��f��^L�Xo�1NB��r���{p������x��9��b�~��-x��ml����{�O���b��c�`E+�.��>��^N'��*��8.�=�~�����~������ų'*lj�EKk�/-��k�p����vݧkk+t���:�g�\E��䣋����щ5"�B)�c���}�Z�Tb����y2�v��B�cm>(�w�6����߼Ճ�F�X���.�Q)��ۆN����V�)�J'Xߞ�����N1��0��E�D�;��4.ܺu^����va���[˧|i;yKH�=�N�@rH�Ga����2���Q<���2Lr�y���$o1��BU��,��q��շ�w�IYh(���\�tn޼I ?
<�Zjȩ���y�3���W]#�o���=0Յ�c��ZJ��V�Fw��q�luc�1�ir�@&�ŧ�a�q��-:�{)�Î��Ȑ���f��#&X
��q� �c.S�ʁ ��Iu!@���wkk�ʎu��:��9q�?ty@����-���<��aE��s��0 >捪߇nXG����`�ʀ�aݪn:��X�s��<K:��	׽r�n�t_I�Oݪ�WKL���\'��ϻ[IU&`��l�#5���
�L�>IU�� �S�k��˧0*ĸ���Ȱ�ط�J��\Q�ͯ%� ��4���E�BPO*k8���6ȣ�.#�5���툄���#�BCx4" ��������"���c;�λ���[�~^�M�r���q��ޕ��S�܉�7�r,���C%\O���ϟ��z��?�7r<��zA@�?����\�� o�q�\������,�,8%v��נ3=͡6�}�N����'� �2�袊�F֙R���+q�Z_m{��cV��:����o-:�&�[�X�\�$�*�9g�,�^y�ST�fɐ�lە"J�3Z�d"��A�wV��Ð�P9t�յq�߂��X�1���������"��;��3�VW��}���X����#!l�d��>��7�abk.URu���N.��x�4��	��ʤpC)B�����-f�M�i���4Ϟz_V� ����
�������>��O��G��NH^z���*,�XeX�o����R]�9k�]�;��"�U����`<O�,���Q�@��x� �����`O���n��סu Yh\N��IJ(�J�]����dv��C7��!;JL�4���.}q��]�mYD�������]'�%>>��ʀ�K�$3�źu�%�����>��rc������xS�Ic����铩���c�ń�"V�?>��7D���7��U��&e��e�>�j21߳��o�1��R���I@�&�'��Mz�0�c�j�<��R\Mf�V��IޯT&]ȭ�qn+��h9Q�O9���<�=9�5|B,?�� �-���↶����r�(�}��?�K�.�K�'�|~�!���.�߹qXhՁ�i'?��#)n��L�%��7�<'x�ǉ</eӕ���Mx������o��7�խ��p�N7���0737o\��WW`qi���Y��pi.\^���8۴�mX��4�-I̮����$W�F�"��*J��!�V�%�ъ�����F�*��U���~(�[�Y��F�� �8���� �i��:	����R���ЕYiӁ����z�GCX���?��<}�����	�r0�,m�*�F�k&��&�/��V�W�U���{��x�*eK�/��yZ�z��h�5�DP]����I��$�NciwX��~~�_����_�/����h�����^d01��/�w|[���s�u,���D]��M�!��#�������Y�_}?mY�A����XR�hD�,3y����hJ�(�0�ܙF^ z�51�Ȯ�Q� �*xżu���#�D"ƻ�~$�}�*���;�څ���< ��e[�!N��|��ͣ��.]E�Y�c�$��͏�5k>U���`͓]2����#`��a�k�o�`}5o�&V�N��)�Y��%+)%04�'�q��+���7�"���QW�Iz�����V_˘������8y	��7RH��;�K�4k����LuΛ�軽�Cx��	<��9n�G���'���{��W��~�7��),.,99c�[|� n}�5�Y`xk�K
\���h�爎~������/�����~�(�䒀���N����ܼ~�__s����l�W����u�x�"d�y0T��1�A�'�ܻ(Ʈ�R��F����L�����V�i;���`����/]��\��5G�|Ȳ5���.=��0@���9x���Qf�K�S�0l�+Ѵ:�ꙅ����k�avj�6Ϡ�p��	O�2�rԥAenGsM�)�:Y���X�*�<K�g�#;؝O��L�i�Y��3��Ĉ�jv�)��*��0;	�&� ��Į_���?���h3+��Y=������>��_�Ǥ�T�;��
D�)\��2�,��q��]7���_XA�֩��p���#YA���IT�V�ST�
Pi��` �8��x.�$��3�q�k	���l�O��.���B��Q��d�[E�K!\�\[�����]ݤ68vmq�Q��o8>�C�Ǿ��|'��h�\;�?��3 BSt�1�n$o�VA@
^�G�@tCs�ԊqN����l}S��� ��H��>����� U�����}���h�Jȉ�chkH@mz3�[c��Y�����D��1�[�
�"|�Îreys�ȷ��7(�9n�}��7���+N�v�>�?��mx���`~nVW�a�?��H��wV-��6���z��X���`��ާO;������_��w`og:-�nf�0�qe~��˰�6Cn�S����0�����vH�4��O�>��?*ُ+��Yw'�)C���W�ژ�'6-8��ʆˉ���U)l�	�Z��`��f�X�t����<&�d|��6PQHPhe��"�6�1"��\�e�­�-�V�vMy�)�.d�.m�;%���6?��?�������~�����]^Nm�c�r�[��f<F�a!i�Map�mp��B�Yh�)��2�'������d;G�̱�֟M��N��(cp��kĂo���T�jYNb߫��֏��s�&Z�?����7�7�?�t���_�3g�a$:R�	K��c���t]�=[��P�X��cE��
�'�a<�ؿ���	��]l��eFs�F6�墫����\=�E�,4b�1dYY�e��6$�;�`��V*�H|؎�,�Di� $.��BB����K����e��Y=M��mJrc 6�T���ZJp?2�>>� ����������I2� �UϏW�BD�n<��|�5yʑ��)8i
y�If��2�Eʪ�Q����S�4���Q���D������@޵!Z��3�y�>iD��1>��_O9�h^��,��\d�ı�S<İ$��A�Th$)O�E��ꨨ2�x�E��G�d0L�7ȵ�7�P�<l#�\�~��&�Ꮞ�p�x�������נ���ҥ+��b|q��h��i�k\4D���r���6_<�?}�.�������>���-
�9A==5���e�ry	�3-��{�~i�NM[^[!���w��1>�C\�/9F�p�~n����/n�0
��"��u3@�!Kk�� ��qx`E�O�jd�Hd��h�]� ��g\[9\|(@�p϶��fU!bI����&O�ga�1ޟ�0+iir�&RK��,ſCf��@�}�S9��t�Sp��2�u��a�[/�/�Ã���sq���"��]�q��� �g���y��C4	<��(��\꾫Z�'�:Lbm����I>�ߓ�:-��|x?{er^�����Ӄs+�ŏ��P4�7�|~�ӟ�u�r��޽�Nn�J���l12�`�8,%^mI+$ ��Vݨ��W��Ad\uk����x -����P�N@[���C(�� ba��X?�F�����3�%�7�p� �9�G��0Nb0i�A��5*)�ب�:��g�s9�G�'}���c=�ҷ���ʒ��1�y�m�����O�fF����ts̏�WvO��1靵���o����"�z#<�T���J�h��[E�-+��;vuB7��xڕ�&˘j���I�T�'&*RC>�-nm�ރ�4sP��$�J��B�ň7	z�FU��˒	��G��<u�ZY���1���i���1Q�
�#����,�T��'R9B���%E���<p�f�fi��O~�����y���]���%?��i'�척t�� x!�DL������S>wn�/���᝷�s`w�p�k���Ц�ܼ.`��fgz���Wn^�y��PXↈ��{����9>��
888��0�L���~����[��O2�&4p쇫�+	V��Qi��9�����M���,t��Zds��ϡ����o����>�.���@����Z�	F��[�x��`�x3#m\V$E�|�}��П��;0:�uŝ�Ψ���̸6���?���#8�a�҇Ҙ�:��L�h�3�e�
��D�R,|NZ�?K�z'	��`��㓺�tVpX�M��c!��q�&�&�^�O#Ŀn���I���y�{��Mre��7n�{��?~D�8�p�߃?a5�����T1����3O"3�a	�cථ��X6²q�c2Z5\���d�p�i�_k�F�
M���t�QO2B9��*�|�'+sbC�y��giY��jP������,3��l����d��J�D��	Ó�d���U�\�8>2�(=���Z����R� ����י��u�j/�&���@B���W~Γ��wj��%̯ɭ�
vOC�`RcX�����|��y��RGS�U�R*@��v�62a�Y᧐�D��[���2������	E2R��<����E�eQ�{ ^���8ץO�<%�����K��?��#n��
�~�c��:w`�ۋ
���^�,��$J����o+2+G�;��������O�R�0�V��r��W���%XY����>��-XY_&���i�+�b���%��Y� ]hwg��˼�.2���n���!��"���}�v�w'�ƕ�tܝ
iq�{{4B�}]���<|"�; E��"G�Rv�C�ny�~�g�V�)�!�!3�*�96=[j���� ��`8t�F흽#T�DÃ1��0=�'�K��`|P��v�Bg�����t�k����˟£g�a��>��6lllp��LM<���Y�&(��>��[��.͊]�8�uPMZΟ�l��
�I���g����'�ʓ��t��Nc����KD���b=������y�l��ӡq�鴜�>�d���qCFk��؄�/�IE�Wt-B� �x�h
�����1�_�{Ť>����q�!��e*k��#�ˈ_Up�*� �eƂ�*#y��$�h�˝�~:]��~���3�#�9�f��q�ܠc�\F�6jt����R�q?RV�Gd��Ɵ"�qd�ʚ�[���2��(��+��dܿ�,�D_gj�ׯ2�&C1��M���I/S�I�
f��']K���~]3^�ez����{��[�����N�S��@ X)ؔ*|­���@�%�d*���n���B,�&Nt���ކ�w��
?��ኟu����gp���կ~����7���c��P�����aɨ�� ��v6�|��__}u�w7���R�t¾���ի���0S3m�ڰ~i.]�D���G�|�4����=�
ۇ��y��[���,m���#x��!ln>rs�]���0�&Z�60�j-�;[D ��igx�޼sY�u���9��K���ڄ�]����h�X^�.�K�m���Ħb�~iUcEX��G<r����<}��}s��:wс�˴�u���S�O�ųm��v��1p��r�e;�03�+7�ov��6�={�G���XG��%��l�E�ʊ���	�-C�:A0��_��Ͽ>�����i)_S�`��؎&��e�35qR�U���Y���t��i����&0����:����a\s�`�����
���EϠ;��n~�Q�3ΐ�ey_� �Bܬ
���N�q^m�xcZ̦J�2�J �򈧕&��Ѱ�tFIA(�oLd;�����g����W���22���Z .$S�@##_��"Pn@
7w�!������'>�N�X��;J¾i�i$����'��#�,W��T��:��ں���T�u+B_�l�D|]��U�I����u��Q?����~��9^�2��W����C7C��hA7�n�)��x��_`u��`��
�H��5޿� z�.�����:�;��q{�>{��O������k�Ϧ����l��M�"�Ґ�����
�~�7��[o;�{���-�7rJjVW�a}u��z��氶��o^���e�#ee�5AP6,0�yN'�-,����
�-�Ӊf9���������`f~����x��`��4ː���°�xB�o1<t�{����m���1�A>u�Fq������=��L8�kv߉B�d

�'�}�D����S>�dwg����
�_�	�s��wufGn��ԑk��Ϟއ��ǰ��� �%�fܩ�n�/,�/��/�ɳM��?��KZvm�Z\Wٕ�H��+<����A�9�I����xU���PMU���ϒNR u�7V\A �I�u|-^N�����1O8�ߛj��V�����qs��|p�S��8��5�Ֆ%o�J���iCa�~�l���xD�*Q=�"^>U�3��;������=�h^v��o #�ڢ����}Xq!�pe�`o*S���&y��<�M�@��]�3�%]�\Fq�G]��e�ˎ����b�uC���+-���CoLh���;+l�F����6�3�&��o��<��['��d�Y���Dx�����ڦ���ʩI�Ĳ�NT�#�L��V�L�1����T3�14��}�D�%n���I~���8G�xq��'ݤ��8  m�`����6�1d/����dGQa�x��9|���p��X�_�0�O�<�;�����S�}��_�5\�~=t'�#�vGt��>�m����ֽ�x�����Қ����ze	V����;���
\�v�6�.C#�E��V�Ѕ�� ޚ�aa��'�l���������}}������p8�	r� �a?�L�qJt� Z���g���d��v��;�Y�q㆘V������)��~w��쐃q&���F^(dMeĪ��B��)��^�)�����a��ux ��,���Q���<��,;ea`� ��`;�v�=�Q\֋��}�5���r�d ��l�I&�).k��H ]�PБ~�Ȭ��Ԏ���u-5MJu���MKcU�v�DL�XH��A(*��Ь[֬
���WS`?+S[��j�V�L��/%�	m�1�w�(��xПuO�޵r ����?h��,ڼ�{���7^f�kz(������u���a4��5����������\PT��XY�@�3������l�:�Ydz�8d<�}�I���lDeV@��c���(��"�@��d���`Ơ��G�{u��wz�r<���WWt��r� ؐ�;�'�8U�w�*��;>�OS���Zwo�ZgD6�3��Iu��z��gM�������k��2�M�b'�7��~���lʫ�����@$&��l(W"����d�g=�e���_Ui?_^#sU�9e'u�r���>OO�i[�p�gz��f^�q�Wޤ���w��<;=5Cl/t�ܣ�y+���G-;�4�{�l��U�z�[�[ 
��]x��6|������ ����A�a�߃��i�rq���f�e_���%
�U�r�/�P:CS��vo��5�K��?����д҉D}���d0�w�T���x�(#?��C���3hg̾��P�r�ՌJ� Z���,Ð�~<�A �.{P��\�dcD���1���cG�4�c91\���3eBز��-jG��`x#K���P���ۛ��BކW~ K+W]{̹�u\���A��:mh�S�r��6=��!l���6���>m��{�?�3:���Y@��|��}�0�鶙�!�X�|Fc˟Y���OP��O��I�,L�*�.�� ��\,���~�����ى���}�P��g�i;+TMU��,�	hW�+(�n֋�Ӷ�C ;:�Sw���f�d�Z?��>.e��Vvu$!���4���;��ńsAs�)����:2ʸ���f��O�g�����ʤN��!v7y�xt���Z����bg�����0������K�tQ��Sd�gff�~\������<肆'����dli����m��1��X�u=�N�@̳��\����:�)j��+45��%�<y���黛�ث�eu�i��I�h��W(<����M��b��C�LʧYƝ�F�*��j!��؎7�s�4Z���ӷɘϽ��a�=�ٖHA����@C��R��07��49'i� �S_�Ԩ�Lت������:�W�P~��x����۽�����?����v�5�����t#~V���J���<nXC�]���ǇGԸ����{=X]Y�Ņ����]]]��Kk03?K�1أ�ʂZ�۟sh|�}��F��v�a*�*�WׁZ�۝���pv�+�&tG�9<P��f�Q�>m�~}���.�np<��	�N��@��Bb�I;�ip��l���if-�P\�$&���8xY�7�|:� ^���gw����[��3˘;b���}��N�ӳk�ʰ��v�x�����f�VV���7n���w��=|���a�h$�r!���F���<&cV6����'��('��xg�'�3��[�M���j�־�7/���iU���`��lb��ޣ��yš��T�L���#f$�1�E�t�ڀ�cȚ�`(;�M�4�![(/cc��`th��h��o�`j|_u�q-��� t�M}e-o£ӈ��s/�U�G++a~�}�������Ǭ�8�Q�����f��%�����TafT�^o�@�0q�P�[ۀ7�w�бD`��8'sS�!b֜ۯE�vœ!*L��*�g�1w^c��������JR����\���4�t�n���Ӿ�4��Y�wV�֔�Y����޳[r�� ��ޕ�vd[r�1z�H����Ғf-I�!9b�l���U��� ��;" d��k���tg]�	 qv��QZ"uퟜ?�R�nAy�_%�� E�{�Q~����G�g\s{x�&�p����M�ƥ�_���CR�k���L1�v~=��ϐ�sf����;-��Gf��,./����_I;^�7���Y\X'�&������B�2���*��;���a0fa��v�r���,va4SY_[��w�des= �
�o]�16τ̥h��VkA����.�nYZ�ͳ�h�K�0@�Z�-K+TL8=޷��zdVb�^�ֿ(����H5-�"�O��@�I �*����
�#
�k�1C��p�C"�ސn ��n[Zaқxa�u^w1v ��'��U֘m��UQ\��DaK��|7�C�8�&�@�OX�2y3�E��FwE�׶��u�%8"�>%�P�����֭5�������%�}�Y8�~X���u5�0wB��7C��;|?��M�yڍ�g��,�eF��:����%���4]��ŵ�ev���9|��N�$9X�'Tf�g�3оO ܡw#�;&�J�ID�4��͒I�"|��r�]Wg(���*�A��1�%��D\t^�E!Ur���z=�k���f��X�<ꕹw,Z�Vf׼I�r�`ft�Yތ���a�c:���������\,�� �HI�ns>�������D�6��z,LSI5�Ӏ�Ǐ��#��g��B~��W��IGwڱ,�geF뇊�v]G}������|��dlӎ�n���p�}\'�u�}L�;9�Z�Fv����O5O�����,��l^l^ѢJ��ɖׄ�J�#�?�,N��b���]c�$�'8�fB������]�\�QG�
���du����ra��s���o���D�Vפ�h��@�	Lm�<��
@�І��A8@���CsQId�Ӑ��l�vdu�^ �����"5xY�z�X�ňiB�Zm��X����hD�Gd�խ��[Us���(nhւ��p`�����R]��D�����ٹ�����|@�[v6Bh�Q��b�\��%�f6F�`2���El�_FN^�Y�����,/P���l�E���h�%bs!q��o��<�
��Q��jN��ۙ_TrN8�˫J�ݑVw!�_����i%v�Z���ֺ�쓏��?�����3y��i�7���U2n�e�%mK��yp��Qu��<o���̧AR9�?��"2���������7_�n�y7@`!cwf�	���D���diV�F=g��3/xyX{�Z��Z�����)�q&�4R/�?�lh��X��&hg^�֓Z$%6M۲awC��-�� Wl� ��
i�"�WiS-�XP��H�I`��BC�2�`��X2'1s�C��鄄����h���\%�\Xap�SY�vX�'_�Ԋ�+Qޘ/� ��}ف,�l�O����,K;ؙv��n�~�|�(��I2"��Lsbդf0,���[3�0�#7����iq}_-����N8d߇ͺ���s?�^}_��2 ~��؛믽M��Q��|��s9 ���ɨ�{$�:�H��)��r��/�g9�Wt��>�m�l}硳l��gܳ���q�G�Y�{�l:�)+E�h34Ul8������ԛuY�.6����6>�B�6oQ�7�m�z�h�V#Zi��gh�pvv,����������ؖ��&�VWdccU6oo�r }f�J��hzAd�_P��5k���3��E�Lj��<�"- ��I���Xso�B���� ����DN	v��b�0��)�	 qA��3�J7��fr&�ޙ'�6K�>�B���Ka���X�xa1���s����4�!U�{��C�4c���qJ7D�s��VV�Ӗ� ��8�NrLv)�1�2�䣏~@�H^�8�gO���)@э�<W_w��V�H���CVZ���Vf ���x���9��6k!�z籕���2����{&5oŜ
��9(�"m�2� ���g��=�PQq�x�#�s�aY�5*7?�{���qb�!��9�� �׵P-1V/�$)�5�����`jLe-�(�r�-l8�;0�d�Mu�C��[����dB�ȏ�Vc`Y�5�k�ƥ�4߶�96�(�kjl<?I W�JN��e�z�I�v6�M3�Y�q%�Z�&_�v�rw��� ,�16�\ZZ�D�v2�0�W��1���t7��^�W��N�;>ϱ���CI���z�h��dֽ��׊�֑:�LCI�������s����4��i�ee�A��F���]�^��p�ϗ��M	����x��
&����@�����S%���8�1`	u�rj�������ӽv���ϝ�̡��[y}s�ӯ�98�!���rt|$�npăc��^X�����+�{��~i����{q��kU��v<
�m/ �G������B^�|~v*h� �`smY֖P�e�-�������E,ORt {.^�x
��qj��z�[$����M�@I�/=��R]`( �g��v|�������
��{�C!���4;��ڦB���%��[R�5���;O2I��-L�hp����i�z"{�/��h/��Sy��D^m�z����� �7�S��;�n�7�|�<5�A�/�t��U��0)�G�,0�[�� �T��uO�aLhe�)��������<�B���	ԛ��h��"�]�9�Q1~�KqS���:LH�����t�u<���.�����Y���8�~-�[c�D�-0��>��	�����=��s�v&z��j�V��-���y�y!d� 4�EG�,qՏ,)����ec��Ui���Uj����%�k5Uv�P�3 �0ׄ-�\8Ӌ��UΑ1��#�
~�j�+dV ����px��Z�7a�y�s�Rd|A#��砎��"W֏]����"AJ��Z=gf`�p����}�M;�Ws��ȱ�y��u!�}4� �]^�V �l*1R��)ۭ�د,��x������/�����>�g��;����˰��+�*�q@K��<R�6����D��=
^�)*G�9���ΒXޢF�
Q���a�w7��6�i�z��~��<�_��M�����9�e |:=�uS2���@��9k��{��a�	�J��ec+��ҹ�H}M����h���.x�b����;�u�ҿ���3wOy�K�ų��y�|�*�v]#Q �E�b:٧�g��6�g0��RG��I���9::�xQ:���I���R�nщ���@?�F���Ky�����;;�Z ��v'D}�u�ڢ�o,Ӡ�0�9������8Tj2`q�AW�`��!�"/��j#xt�#��b�D�e�@+�F�y�`FC]�C��frz>�� 7F3�6��v���@��]�� �����=(q��b�ɽc*5@� �@���s�N�����I� x�v q.�(�Q ��p��U���cAS����>g�M�/���iK�!�?��P׃1��-�f5��z��r��-������a�'rxp$)rM%!H�i��xv�f-*' ��\���i�4��M{���T���w�ٮ�jL3�o��b�Ώz�ޤ@"�΋qy
����Y6���嬲$g�DM~�t^nX��T.,�2�(B��)$�1y���<lVn';4� �/�l�)�Sᰎ�Ġ�*,�$�����O}�
�1�HJ��"-�ZS=\��rC
�՜�4��e���he^�!68�Y>�"�NW6���\�"��+��>l-�s9[[�U��]m�(�C���S��B��(:�-t���J�(p�dǦ���ծjLxL�B;��!�4�{����\���<`�2�ç�5���]�����gzo_܀�U�p�H��#|��{�b�j��Q(#T\Mm2��*�h�NDĢj8l���Ǚ:�i)**@����pv�곔?z�g��V5�^�����M�\�^�~�{�?��J'��~.��_�7a�����:�Ĺ�,�\�柏ģ`e���$u�K�[�U�Z��]	�m����	Yy�����3�HU�|�a"��b�3�h�g�y�6ϔk��_�qU�f ��=���2{
ۃ�{���@�ΌK�|�-d{� �NN���N�����?����1���^\F�@/�v۲��"+��%���.&�FT�-MRK�����)����(���J�ACŋ�q,eЧEt#���,���R�����`xAu� �P!��.n������n���&;��Ua���ox�M���7;n��W*4���K]��ޒ��0���r|�#{���Ip^�x$;;��D���6�Νu�uk�ǌ�x��"���Ӻ���s1�͔dv|g�S�/�'�3�%`�+p  <�@�!��@#�|Q��@���0��3��'a~��1$Xh'ކ9_��{?�J�����A�UFn:,5��A+�7aS��9o�B�-<��C4�=�*qΰ�aK-,���Iz�,����6�`��XQ����ſ6$�p4�50�ޥ+�
��;��L��c�8����hJ��ek]�
E><X��:���8�3�ar(���U���"�0�x�}FWT�[e+TY�v�%�9�����15���y�a���v�0�Um9[�ي�} ���u�p��b�m��j���	��j�6�NGn߾�P��~o�z�����"Tp�0Ͽo2b�8g��T�P�
�0�#%Ya�wk*ZJ����g5�|e�Q�!W o�n#-��u����rp��ݓ��� `�����a=8�jp�eyeU�nݕ�͵p�|�{5��g6��󝩺X�2�Ͱv ��Ѭs��)�b)e.����p��������R�G햇�c�sH����c�s��C�hD�"�s�U3]#�b�k�Xh/��W���6�\�94�����f7e6���e�7^�z��yv�l����<a�:��O��!a�����iR�U��9ٱ�6�##刎6�T���t����-R���%z��Xt�ɉ$s�������2�}�>��ؙ�����8�R̝����bO�q����ryG�ͱ@��B��=���|��Wi�јbiiEdMr��q�*���rp�+�~��|����?*O=
`�8,=6��tڲ��	�a=���F��!
Oƚk�t���Zu3�`�!��"-Y���i%c�Kʦg���H_��d�pR��$�bxο�)�ӓ�!Y��Jmߵ�eY^��V ��YX�Nw�z�W�A��Y:ƬEYq�L�l����j����(����lIw�.;��x{{��w�+�����)�v�\ݖյM��R.R�V�0�b�z����yW2���9�b ��4������\u�R�R3��ك���н&��ܻ�)��G��{Df;o=�',�]3�?'Qp�αAW�Y��>r�����iC|�g���.�M�f��K޽z�7����6��A]�ի������°��yT�BuskKVWט�	p�|S�x��'+����� �����
x�5�~c��L�1U��k�Kl�gf��c#�mf���B1�(<��8S91����1�G�=�l��QcH�Ҁ��j^阀:+��X8�)@V�]a�Aj��Sr).q݋bƻ�����P��`ߕ��k��A%^c����A/Bk��mbv�����������*�3�j��&�$ �V�j �X��Kas&ĺ��3��4�6�s����"�To��܂)9 ��/�2g����,#%�� �3@���o����2s�NO�xN�����Ѿk��
 w!8H�@��+U��cEu��X�&$i�G��S^Rc����Go��sIcM��7�Qp�%1�/Il2����60a�{V��[��گ�/ó�%Nۆ7Is�v�灿�����❷O���u�qA�Cm�l����{a?So���d�J�93��	Y%;
H-��1�4�+^�*�ڛ�1��I��8�Y�r&W.�EmmTg���a�����?�n15*�Jc��q6����G��C��Bͫw~"Ϟ'�.k� ��D�RF�Z��y&���O���������Wrvrx胰�Ų��b*C�U%нug��R��T<�����Ԥrh��aP-Z#�?f���h�q�;�)��t@f3KO�bx����c�g�P���ixO��s��]y�du�^ ��a!��ԁ��Ī�E�r!����%����z�PU[l����]ٺ�P~�~p��w����˟��o���i��H~�]�V� ���փ�"��b
�[�ZWEs�BcAP7RlY^	���`��ݖ����#��r%(�#Y^�;�yyxG�>ݑǏ���UodŽw�s$�>@�l������2�3����GyQ�'��c�� ����������ɯ����g�_�����p-�P5��y�kk��:�#��կ��wecc�����=ޯ��R~����S���g���V�i0�P ��RU��6�ĝ�L,�  ��+e�-%�M��`dk�� Q����]����X�Ԅy��� ��D��絢+�L�T���P�e-6�\6�[�Q�-h/|vv�����B����*%;�_���sc�.a˻) ���h[��GG�~��ll�bZW��>86��9�Q���G����n?�0�k���j �i ���}=r�����	N��:�`�2I����LC"�M}4BZ�2$]�:���m��;����h �"S&����v��	�N��V �`}!tvrJ���H	�{������m��	�kS
F�@G��*5i3'�x��w� 6*�1fo�A �hHǄS7����� ���q�%�: [�JEWQ����3�� ��
�e�`���unZ�o�z�6͆^����R������0���|KMe��H�z��u���\�n�i`�%���!b��e��s�2.��so�|�4�+�ҿ7�2{&�EgY3=���cq���>O¦���\{S�XD]��2[��'�����5Y�u�[H��<=����`G�\���6��ʢ���?����}�=IGi޼�?���������"k�벰���ۼ'��£�(#}�8P/�����ZfR���GY�`�a���$,P��`��dp�~�9�?��Ӂ�UYY}(K˷���PV����z��[�2��L�����c0-W���囱�����U&;
�T���>�j0���������7��/��'�.�eeF&8�?Jy�F`{��0$ �)�z�`l	~����fQ)=%2�#|���,>�kM��ɫ�C���o�އ�3�V]�jv���l�����)#|��N��o��bnf�!���e�V�H/[�L�R�������_���?}�9�P,�0tO���粷�c�5i����9������(�)���%��v�����7������W �����g��0>�|����Y�� �zg}���@��pV �hB�BJ�6M�#�ɀ#9���<����a��9UE��������dt�P'�!��]���C *��4��`���j�Z��:2����j���v�[a>0�(xx���l)�juE�wU�!QvZ,w3.�Ւ��4\���4);�|2�׏�H�ʘ��B�Ŷ��Y�b�9�q-�v.����&g�˼/^�ڕӓs-�B�oLuscm�"[��8��f�Bj= ���Ҙ�HYj� m�?�(���k���y�����>�)Ϧ�ְ��E�L�Hk
�� ����H*�U�:��M4���}�Y���
f<�_����M��l� Oka��P� ��ÀNM ��<����\f��,x�읲�����m�4�칐�<_��-f�����y@{<���{����*jV��u�8��	�Y��M����>w��� ��A�����<��i��k%���u�%�{��OC�ce|���6�`Ϣ�-����Y���<�V��iI'��fD�wN^�H ���﻿�J>�bLb���]Y�.,��{�O�<��O�"7�R ��z��කhY�`����*�|,J��(dd��V�F�b1 �`��6�@�(��-�V��U͸�
��(���=,�g\�������قl�~Wn�yW�n`�\d�n�D\Lr�k3r�G���Z[~�����q��s��lK{aEV�7ü-�(,`��2t�2�7�ٔF[�`d�t0V�*�����z�� ��jvK��m� #<��Yna��� ��U�}��s�߿Y�Z����FŪ3ÌGz�GE�ޥs`��}�P�,�x�"r���%~��M��Uǟ#&�Pc�D(��?����?����,�[��d���=y���l�b�+޿���������k�s�LV]�w�Q���[o1����#_~�Up��������ꮢR��?b(�ѣ�t.���uk�!l��j(;�4�fô]#�eM���s1�^��gO噠����2��Zu�I;n�b�.��zp�ó�j-K���"�GT��P�v��	��S�T@l��ΊhAwQ���:� ������.tz�4V�D��|YE �������r�x�g�+�sӯq<V���YF68b��������t�vѦ��O�Y�-ű���&8C0�Yj�n2]4c�Gl^c�d.�X�h���EɄ��i]~M?wl2hj�`�2cK-��s7�̵$���� �\H��IP���V����ĕu�`�|0�;V3�y9�skk��,K+�^*J�LE�p���P��us��� �N�ΎJa�nmm��u	\q��^�C�3���$3��h+�g,�E>�ҫ���9\�6����J�8�њ���G$�m�t��ei��Rn�>L˿�_ӄ�v%'�r~֘L�0�[fs�	8��0���}n���S�nG�&��i*DL�f�S"9��F�Ե��p�rl1��i�N�GL;J���B|q��uR����k�֨4<�w�=X	� �O�U5����Cc����� �:�ܥ`�������b����|�]�;	�I�7^!Nb.)Z {���(��b�	%n��!@�Z��4,�G8���Y8�[w�}K����,��e��(,�):�y� ��������i���z��'����pME��[�֕ŵ��'�`xoɧ����o�,_~�XO��<��o������bU>��XElq�t1BjI���"�����q&������G�������޻����������#FC�:!�Y�]&b��y����6B����s���}�P�<c�:����>�+<ȫ�+��G�[o=��"�u����������_���Y�V �Hex�w���{�������  zq1��࠮���'�|"�'Х>�Y��<�w�ܖ����G�~^�G|�v@���]�d���/-hp�F�E���vw�ѷ�z�̏^�i��6nT�1F'�~��wn��*:@�Ւ��w��dg�\�N�d��|�<�	-�e�.әD��q���Ÿ��������x I�̞�����*��@���y�r'B���l�h��^�O�oS�ǌ��U��3�%�͚M� ���Fb����)�(cA��XIՊ+�����<'�pV䒚ݫ�8�f� �K-/5a��FpސV[]]���uy�j�cq`ٜ�}]\Z�s�;��R�7@Q	։͇Hɹ@�H�����=U�d���mn,˃��=�A8�2�p��pm[m:ap^p�c� �".H��_ �/^>�/����=��Q��� no�م�bp�ʢk���{��""�����?�b�(��E��j$3����辩�xS�~:o���k���۟���ŗ�$�M�(�k���kl+�z�خ^�<����s��=�0[���U#8N8���m�V����2��%��EB����>�RO	���{���u�D�׹��U*��55-t�Yq<�E8;=���v���w�ރw�jc�1f���d�2"䥅&N,/w�U��x��򈣉�@C��ӊZ�S^���qXpÂ�zu�N��cUe@�}�} ��,,u�}[��������J8V� �n�?l����4��\7��t��g�w��@4��d�Z�^,-,��z�����'ۻG"�}�!��B0��.�:�>T��XQ�� 	�~���E�a�D"]��o�y�yk\Å��i0�y@�����/^�)cb>���0�48�^Q~�y��1:�	��3|��Y�e`����d|��0��fyQ<S�����'���N��� ��X]Y��������[���#2Z���X�g�4x���sX�?��C�O兺lmn��/��͖|��Wg��@��N8�r8���,��>?�s|k,/�,�hU�*S�R��6�?�g IQ3��8�S�y�$OV��m���'���Ԑ���g䃟��Mp+��>�(����ю<~z ��y��d����P��,]n(��O]Xh�A톯�om����9�s��	7c�$n�K2e�_�x*�/�y&`m�E5����H����^Y%��ZeI�5��Md�p��h4�f9�F�j%O_��*�kݯ���0WrRAG˔�T�.��+8!�'Z��{����G��:��LX	�Æ��$�%���y���h�GX;vww����0zɵ!�$���ݺ�,o=�%~�n�����hzX��T0��0�H�c�1�T!�5����0��fg������枂�E>w�1��C����>	�����lmݢ�{���������Xƞ�v-�{UJ�ev�T���}�(Yٞ������U,��
�M?��<�q�>��l?���7������3����8���/���E�F#,w�o-���A�h2r�T�}��I�T����������ݜ8g7�v����f4��������ޚEN>���f$t��dee�6�>�?���:���g�;�3++k,��Vk���fGG����s��m��j9��U�� 4�(��S�N�ǡ�^�V�XS��I�!$�<�,�H%��v.�ZC�:�x��C[B�ahyb��YZސŕ�r��{��y/�&�h@�[Kڨ�%Q��4���r�y�*��(��l��� ��Z�w?�'YX[�A8�o��T���7�|G��޽��B����`�2��@���}�z��7���[h!*�&�{��`�4���ݺ�!��O� O���>���A�/�3N�4/�s����ɵ�N.�*�ຠwָʿ�l����R��-��Z�B�x�N��}��{��9�d�'��aJfr3 ַ�~[���K�����=�;�'����s��������w����M�·�ł0 ���e��Xc���v��A� 

���X�W5��:ڑ��Ƴ=��Ќ�N ��6�� ��ؒҙc�"hH�٘���jK�����V�z�p��}Kn�]�'�����j8�� �頂;zD���ݻ��� ���8�\;�\�լ��_%|�����d��U zパ1
���Th?�̔(b�y�}�I��0��cHSe{`��ƻj���ի�Mf��xf*L�˹��z^�'�Hތ��J��ZG7�M��h-��E�_*�2Ɗ��9��?#��hq18>g�����m4�������T�����"�Q(8<{�\���g�ǈs���Lec�%�xGn��
��=y��Ep¾���3:Q����ll�ʃ��������*u�c���4L����L��ڱ�#J��~��&A)��v�~��<}�����.0*�:|s��^��ܹ#���/eccC�߻/��/�B���a�U��Ω�ʲ]�f{�3��e9���L��^��i�T|��)�\f�n�͚��څ���.8�N
�U�掮����&�˩�t�:1.��>���jdF�����ͩR���tޘ�M\��7o,�D�*��y�"���h���ĵ)�Vx�:�N�U��j�d�y�Wi⩖� �'����Q���iS��1��u�}:���E����b�B\��z�W�ꥪv���/s�ƃ��T��jI'�n �+aq�T��Nf�mv����B��c�H'�ջ2�4�!�x<��Ef�=�,)��!w,���&˷e����Y\�i�#� �*����g�Nݔ�_���z�q�|ߖ��W�h+��䓟���?R?�ų�� h�PU��|���1�n�]��9YE3���>�;��*�(,�ݖ���� ��:�ʹf'��?�~��d��S������+��{�W��W1��0�3_��XG����	􆬮���۷��ek�Lk �PՎB18IH_�C����3�?�� s�����/���C�vmĐ��g�j�Yg�4G��r�=z�#�x��]І��L"1�Ώ�d������D��
�*1D���z�[�=�;=dj0)���d'�FU�L�+�BZ-a�S
u�����A����8����Չ�������8��3�UK�b���h0�N{��d�n���9�n+���Z�Q���ng�F�ҥ��l!��� +��+a��s���ԉE��Z��p<-b�>s� �F[����`�ck�A��xUxi�1�O�`l4�eCګ�yķ�}�NkP8����jDv���s����p}zj;2���u����d<<
�g1�m	@9`:��zp8µ?8<�:��yu�f&*�ڛ���i5��y�~��2F0�Ŝ�	�ݩS,`~��8�Q��J	�~�FhGZ���ur�j8���� ��?�s�ep.:�|����r�o��_Ƅ���,��|�i 8}�7�&����2ȾND�[�����y��\�7�3��^g����?��,ϻ�=R1ەe��:\o�y�����N;^T:���Q"*�e�;VqT]K�"]<��&UG6����t�B�����v�D�+<��s�x��%�`�$W�ܪd�Ox#t����9ؘf0JMYe��%�6�8*�m��)g3��� 8կ�P=���1���TVT&&3��`d��z��������@��M�4��a���zP�,���P�<�(�k�o�N{U>�蟸`AK���W{��hH�9ͪU:i�4n�ZU����^����;t��5��n�.���9���Q<�D.���޶���1�P䞽:�N+9��ݱ�ނ���\'؀N�7��s�6|n߹��]���y'�����)&�ݿ��� �sR������ =��Î}"�(d�0�х�Sa�eì�A���w O�}+�{d��67e}}��a8_���oCt� ���&������B�z�1�V!����V+��@>�ý��y� ��t��)A���6�n�Mc��I�k�X�<RtfDX9�ʜ���~6e*I���
<�y�b��$���ГeqZ���k�茙�Õ�� �8����SK�(�^e\�p��Ue��_l���Vf`1bԧ��S�B���4�{��ol0�
Q�"����" �ۯv�b�x�H#R�v g�!::ܑ��__`�K�6N\֔p��Q����kY��Tk8 �#gQy")�W�I#��_D��ż=2���"5x_��b{gO��x��@UI�5���p���`�
,������2���q��P�˕�6���q�,=����ϊ�\��˶�s+=o��sN��7�1�RBe�ZRD�s�53�0*����F�[Y���M5�0v�+�mLm������3cvqN^{��"8&��`��y|�ؠ@�M�I�U�jb��Z$��X��z0�����,.��2��YZ����LRP�<��&<5�	y������F&l����E<�g���K�����L��aU�C���P����|��_O�%.�.|#ۅ�q.��'AY<��jl(�kp�Z�xG>��������ٗ��w���^`1�$U����ɞX{N��c;���L&ZoX��sȆ P�d���syo�ޒ{w����<���#����1�yd��9���9����Z�SL�}ne�#>fn�Ұ����p��# *0��H�C�o�qqa���Ps8�����2��ڀ����>�H���� ��~%a� 8�3y����w�%+��fJ��0<]X0��α4�
���m��n F ��rz|����������)ȽE�WX��p}��1�C� �3�^8B�8��l�AM4;=V
���҆�1�8�3�]2���\�1��|[�B�,-
=Q��*
H���l��|�뭓�׵�}
�HG	U*B�HZ��f��ﬀ��]~)\��)%����,'O��{�(�c����g$yȿ�8z
W��`�<��v:2ۢ�ED6~<:�8QRaX��5�/RI�p��u�Өe̺0��^���u��#�Y83�zƦ#�~��9���X���!R'Z�`{(Ѕ>�wZ�������W�q���x{��w��9�³�fN6�ς38�%�_�P4����i_�5�O>�#$(��=��ga�]9����tC��ñ~�9o���k{�87�_�g)R;/nj:&���G��hm�ԊD�6�,o�dI�&��J�Jt��g����ʹ�)����@Y���`S�h�~q^�3���q�RE��#�4.�������sfm$|Q�^t�Ӥl��bW��6n>X!Z�8��yF%�g/��Q��V8 ��[X�}�HU؎���`:C��Hf7u)3�Re��XP�Z��[kb|�h�&�lЛ�1���X�PU�n˻�e����`Gz��gll���s��J23�\9}~GG�1O�����9�*�6�^'[�ֆ<xp7��|��xX����Wo�,L���oo0ob�/+f(��&�������8��2��v��5���qjp����S�	�����������ԂJa�[��}"?����{���!����3����b��W��W8мs,�� ����[�i��o�!�{��m���N�RwHm���C�K��뇐2��!�?�+;�En��W�1NB�\�__Ѐ�׭�q��ǞW����4��}rz�м6�L悊�J��n�i�s5�.L�"��)�v����yQY2g���݌��C~�.�g/S����v8��B/Uo ������i�9~JT�R��0UW7e��xb����y�^����`����XGn?�nj$,R�R�2�ش��}�"s�������.�{��sQ|�O4mh(���ۧ���Ģ ��t8�}��gli�0�+�0��U��!��������_4�@�� �o��GQ��$(3�{y{g�ǁ3����;w�j���K��i��K�����sU��_p޴@�:ۅ��5��iW�sL{^Z��'.=fN��/�S�8�y�7�S��(O��3��+��<�^\�ce�d%ˣߔr~�Oz��\�SD�����q��& k�!�VM�c�{�]oT5pdJHU,r��{��ּ�F+������M�4�K��hD^_�y�1�T�K�<�,�x<�j$��S�0[���hTa�G�	^X�Ʋ(Y�aF�go��B�tEa���򵮻M��l�O�#F���?�fW��w�����v �^|+g���r��wL6����jؼ��Po��h����8��6���"�|��Z��޺'�~��x�V�3ͬ�U`�?�6K-���	�@A�� ���@,�K���R2�`H�m0����z����_ʫ�]�㧟+A��7��������o �oԜ��������M~����7_�Jt��U[M7J�x���&N��) ʨ�?99d���:���( �P���7Zw	��� �C6@����P�l�$�زh�yg�R�I)=<+��c�ɍ���3���d��-������m]ڪ��<�,�����E�L���]��j���8l%�㭉ǣ8�.�1Aoj��D�M4�kLF��0���;ދ&�f4�!;i̷6�д\W:+U�/���pe�Q�������T���l��`qU�053]`�~�Z�b��d^�6$�u��Y�������{L��0w��4�x u��nHܬH?8m�����C(������M�s�6�3�!tO�]XZ�V�9P��Ġ?V]�Xs��+9S0w|�YR�7��Qp�����(q����r��}�^p�Рiee�ree�⯛���H�U
��(*��f�Wy�,����M�������6q6�O��dO�ݡ�Ԧh.�3���+}6���} ���6`}�Y��l��;��y��R�W�R����qe�u�$�8�� 4@��%�Ы]��Ŧ�c6��,1�l2ɴ��xE�"�Ű �.Km!�W��9YZ��C��~!��T�Tf�-R��|�d�#��岒C�q$*~^�v�^	��=��.�jYf���'�fyrd����&~�N�7�����F ��Z��q'8?%qv�-��V�gY���(TRiɣVТ�6��jg&7 Z��ׁ]-�n	_�cݑ{�6eq�I��8J�i�9j���)��s�� ��Ѻj{��\��n�����7e�����ɹ�i) ���u����5� t{r���}:x�������|L�R�<y�L�>y���,/���®k?����m�����~�����M���KV�C��C�Xd�SM���2M'}�7lo�d����ǏB���%#���Q����K����:��'�������%��e���qF�T��~F����+|@���=�S��L"{��QJ�`��+�T�s�J�He��&��j��9-�sp���[$OD:̨�x�x���f��(k��v6Jy���'a�Ga��s��Ԝ	s<� ȴh��L�����F��zF��i��$#��|�����T׭�^��'Jep��	��NF�jA8\c i(/,��� � ��MN���!UgL��c���ѱ���9��8�o��I���A ���Q���ۗ�O�C���}���P��o����}^�Ęb8RP� ��4����4�W8�p?>�Po�AG�Z�X�9�ZR��z.�6�47��=��/����\Y]�=����T
I9G���R�?@��/�[ q:���]�U��V�e��Ο�us�ui,R52�K;��^X���4x��O�M�î�+�\�̏k�X��ƥ}e�҉:��d�[�������IK�;R��EQ)��f^������t�i>9yj󄱀h��s�uX� ��$��h9"�00$ԓ�5��k�����4���I2���|���E�U�<�X���S��D�L�yt@�~�&V���b�փ�j.I�&[M.���TZg�o���i��EVz��㩿]c����,F4�.
J/�n��-����~1bG4�:a��Ũj�,�T��<�X��#-V�����ӥ�!�P*�V�0&k��Ԗ�w KՐN�{Bj���5��T��y��nΔ_֛�z0+/���eVE�U��}]u�YW!R!)4��',�R�0�FÇ��Ej��W�����	�$}�w��Cm3�P�;o�-�w G���8M����׿&����B������o�U������)��P/��1���j�H �B�e[�������(��1m�J�ZѢLo�
 ��{,rr���iK���n�G 0����3�A ��rh5v���P��;�Qø��xʂ�� �����r|f��]�MŨ��[ ��~�#2�t���"�_�h���VK�<�d�������U�F*+2���זb�z�q������`|�\�O�"["����Y����]/F����S���7%����1�}q0D.t�8
���X;Y"�B�n���:����1�lթc���'c�#�_g��45V)�s�p���=�BG�<X��.O_���*8c/�}� H��� ��C��?�e{w_��ڡ��˰Ỏ��H���;��C��4���+��)o�ڒ���p-F.�&ǪD1�Np��`U����CL�r�?�?�!�q��_^^aa��o��S�7ɓ�~�P�u@�U��M��ň�Ik4ѝ����`�v����yÃrDv=*3���G~,���7\��Z�M1��
�ٸ���]t�
v� ��~�D�^~V��AS!��>/r���#dq���b`8k
�KmzD�'3�ȵ�9�����\�5��x*��r���oj��-S�6�d"ULǯ��DL&��ex#B��a�d��'ob8�Y�q�J.�h��ߣ\TV��(�I^D���-1��*eҠӈV��*�R�uyF�`l�����4�<E1�gveu��Âqz�4�َn�B�M="��s�JEj9(���Êz��})�4��`��:faL�Y���%���� TP�`���� ؿ�vH��o�\8�������E~,R~�w�'�.�,�����W_ɿ��������G"4B�����{��������.�^x��VG����B��w�ݦܾ�)ߺ�{"�;� Vv�6DkU�=T���E���pދ��ZpD�mԇ�aJ���TV*r�V&�iXaؠ�
 ��l�_~�����%�� $ؖ)Ta����Y �۲��N��w�ȋWg���Xc���3�����R����3偑Tn����#jpc/~0��%��j�4g���f��k+�\���G'��W��a�?���N�Ҵ�C�/�0� d}csɤ�g��t�V�$5pܧ�9HHbх��i��*����~_�iSQ��H��i���e�ω�=��T�<}�Y��$���8&޷����%0�CԨ1����C�}CU�Ӊ�D���X-�x�p�}������2��/,�5��$qK�5�ܢ P����ա�����p.i8�N �}�N�����9ܩuws�;m��>��fy� l`���.��*0u]G�M�rT�u����x��۴��9�Vy(����Q��j��9����FE)��Z�]�J�]{�J>��b��#����Apu��C�� �J�pdG�3��'U8�����p������v\�����������OǓ����G���h7��|��yD;����k2���XCᨚ����9t!��ͺ� ����{��([���Q����M�GI��}���Q�@��X����6�8��/L���>�dr���V�iP�Ţ���`��\�Vx�<�RH�d�Az�B�E��[����H�ɔ��4:�1<9f���򒬯�R�ro�P"��:��H�Y�2��`�=�P0��zWePɫ!s';a���Ç���|Ďi_~����_+�����`,rQ���BM�ܿ[>��p7E�c�pF:��a��gg�������   @����m2(�c��R�Ls}k [H�l6�0�U%��]�02ί�<��(�����D^=!�;�$ 6�p ���l���ɹ��6�g;rt���X�3N��/� 8-D��=Ȣܔ�כֿ��e�V�l\�кHTZDˬh��(Om(��rH֯ol� �i44�@��gO�����!10�"�T�3s˪c���tq��, �">��7 ��Xs��&�,���Q��CV�9�#���w�)OC^��5�j<V���׵�q�`|P�@*MѶz���R1P텙�ȝ��8���ީl�ܓ^�ƭ�F����X-�Z�n���E��'��"�j�2����c���8Fa#�[-���Ë�¹�1��m*F���,{b��|����j�ʱ!��),�U��Ѣ��^'��4Szr௹�S�Y�������=Wn�����tg{�4��YR>��i����h�X���2�~W��wg�Ko�au� �v�	���vf�������Y��RAn�4g�`�E�sήzu�q�VT�9����`g��������!��_AiL{i�'Q��W)�tZ���5T��?as�E&-.�2�i�o��2�&Z���&�c�O��z�c��;����Z�����%Ņ��%�u���7z��Xx�8�qY��p��Rƃ#9= a�	<���R�)v�E�T��9��wo7�7J^���|����BW667���(~I���.��a�k��?���e�o�$\�+�%l������D�{�X>�˗�>�y�� �G�=�b���}�s��HCȘ���Y揧>s+V���'���w���W���;�o����_}M��C�f�l������1�,���g<fU<�f��5HP��>x�C�QG�=-�Tc��wHnoO�={!�o������s*�EQ,R��Ǻ(�kR�ޒZ�+�q�}z$�q�y��g���V v'Q�D[�2|#{1����2���(7��"U�Z��B���*�SU��r����GG�m"��������j+���!�t:�4�p�vf�J�& zx��>�]�Pa,Z�) ��|���"f��0��c�)e~;j�X}��Q�vd) (6\XPE8f �i��a �ϟ�
���9��z�^?���
�զ,�ܡ�7X�g�^ʋg�ɰ��%��i�xTc��x\�� ��vp�j1�
�����=^�Ws|��5R`p#�ao�H��ϩ��B��`�P�����V��Ŝ ��w^����4:к.�:)���i���1l�b��5WleP��*�n��.;��<z3���m�`q�������5��$d�\R{�Wbv=�`�B�6|���z���Y��۵�r��֝z#+#�!��b:;�̰���e�B�k�G�o�9�V��_皉�ټ���9���Ek�
����-op�H�Z��E���A���%-l�qgØ`�<��.h<�7��d@Q�@[hk�v�؞&�g�	7���B(M�UB�aAY��1:�37�V5�\���ע"�`���
�4b{1��إX۠�1����̂�͓a>w՜A�Y��Mo�r�.;Ƽ��k��B�	@Pp�^�(��+�3�S",���w��� ��?��L,ڣ"��T\���C�F��?������w�糡�N�9����4�L��`�Q]��3<�  M0
H�x�2�޽ 2��5�>�X��AsW��tJ�1h梅p;�d�#1�V������y��6�� h�Qd�v�0��a��zpn[�R	�.����
@<�K�є�֤r8R�ԕV�]׺�qɲB�T^h�c�$Y|O�k��u<�l�u�7����2�6����ňM�pC%�Fڂ��J}�>a>�^��q�j�7#��F���]���d;L���2�1Z���N1S5"e���v�s�(�%��#��8��$}y�jO�����)��L%�KH�@ Ib*#�O�u���l�o��]�o��@B+w<��y���,�|Oꍚ]7Ua ��3S�27�j-�	�I�xT1�5�>?0���0(�\�3z�*QQ��4R��f�N��i;�}����x�#%����i漜�Pv.fus�.��۬���)��H�������7������(�M�<2^
ٗ�M3q�-� s[�10�y�&a�oi��2��(Ή��;�����:6�i���68��\�Ή�J?�A�y��O���i�Q>n�RVr��/eycv�i6*�̡Of�1�#g�"1�_%���Ƃ��ja� ڭձ�7�w(�����u0��Ҥ �:�qi_~�?r��-q���2e�i���@���Tz�'�DEؘy�4&�LU�gk�F� b�P�S��2r��(��, /:Y�o�v�-�PE�}�7��y�����cd���)�K�-ߑ�_�k] ���3��b��}���������Lm�t�},�loo�������|���.J�]�;q,D��	kg�� ���@}��#9=9e�(�z��
�{��!���3]�p�!5p	���F��� �|��Ʋ�b��0�_9�©@%�7z�S�!�q_F�G��׻|U��6�Aә,���ZWVAR��Dh��TblM%�2�#*[X�J���p�Y3���^������B�r�Ūo��t"e+�k 
�,��;�>��a?��(6dBU�<��(�Xq��=V�vz�tlH�R�G�2��D\� B��vϾ*T\B�V��^YY�.��;��=�ƈ���sc_��	�q�GΘg��!#����h�S�8���ѩ����y/8h��]X������zq*�����'@�k_�^�����+Y �~���ښՠb]�Lۋ�����2�Q�l�u���#B!�9C�����ʅ��Y�r��c��MoȄM����M���rfmަL�G`�)���e�	L�j4�^'9�	IK���b{���!���J�]��FS,vT�=�Ǚ�%�9���~�!���Z��Mѧ��i�Zqp��AJ�O���I\`̂��kmdtY�Q1e.y�B����"]E�Z޲�&�k�.?E��;,r��Ҝ/��kubb���e�4�k/9`����<ot�A�/�$���BQ�K3�S%���ht�X�%�$��0��0u�n��������9i�����Z��,I����<��X5�^V�(m9�E��؊+��[	s]��z�9~dp/,&\߀N�t;��0��!Z�ud�ryg��_w���~��N��M��>?=�	��D����d.�}�H��Ͽ`�x{{�M��EڶF-`ힿ|%���	 -M��+�W3'I3YTy �M�8�{x5��{|?Z�"}rg�K�����<z������AL�F�����ۢ�3f'��u�6��}�;�[�-l�+ឫ���Tci ������6H  W�Xe-�*�� �6�.YW��z����l�P�ؼ���8x�T�V���.�����yg�c�y] �����R�(2���bo\Q�̯i�":� ��B��0����Ъ�E�*c��*{��A��0O�@D~w��b�m�Ր���^������y��ݽ�0�,� �Ƞ��o��Y��I�<���2��<�{ڝn ��8�l�(^����̔!4�Z�l��]%v� q���q.�ᙍGYnh���3�&Ff)�K�����%�*NJ���$h�f���Y���i@p��ռ��ڵy����`�ئ��鱕�ѝͲ�XY����/$�N�e�t*�U��^@�Ux$�	yd�s29�b<��r�)��N�'����\f��4��}GR��#��|nDJm�K�e�R�>��{���'kN�1ET�@������V?�XE�o�qd�	U}|�~��J�������7NkU.  D`�Rcx�_,��"[��rt2�눆���:����X9�Ź�	{o��Ҩ8pF�&����j+ॄ�2�ˑώ_��{h}��:[�/�~\��@����)*�{�i��x�"��8F*��mV�w��+�5i� /�-��&@�$ o52'rc}I67We! ���)�k'�v��P
�^̗�Q|�st�t��{y�u���[Ӌ�b�������>�&���I&$!O�E`K�$/�� �����D�W �e�P@�b�ʕB�$��  }�Vm�5q?��O��ޗ�ť�춨�{^x�b�v�*N4�A�g���;cS1�9v�
��Z���0~ I ��j�d9k]CG� N;���^h�����`�Unb�
*̓^�H_��Z�� �~��c��P^T���ŨK6�h�pX�:DPi׃@X���T:��6�e���Vp�C[91�5��ExTk�v=��,0��梪�nK�b4�I ���
kk˲��(K�^�����C�r����vምPMS*l�q}�!�*�"�q'''���}���>{O>NV�ݑ#����(�ǫ�j]�Om ��RS��BF4�B9̓��97 r�u�"��H#c�xE���ٴ	�����T��Fg+�9/�|������5*����{�e�?&Fc�������?SΗ/�ͷ�gq�8��>�i�l��D�?2���6��;H����f�w��iZ�l�B���x�$f���A�;.���QD����>����$f��j�����9�ֲh�> �϶�S�~~���a�-�޺�;�����k�v�T��d�Q�oRD�7�������h�\�tc�u�	��$ ��H��t�K����ς�g�4�~��G���Y��?��Y�!�����V�-�Ȫ��PL̓���H�3��"[�ZT��.,��]�o�����^A�����:����M�|���:��t���Ѯ����ٹjU贃��pr�^������j�V�F��F5��	�#��I�oW-�X�����|�ZrU�LN&�:֤�n0�7���W�Z�Z'��q�<KlR}jhG#�>�wɲ,Pc��J.W�)
nP 8j�5
P���n�Rg Ih� ��)�d�kt���j�����#-�<0 L��^ �Zю]���%J_��1}�䰴-d�"LY^x����n�A�`���f��L5?��O�:s��y�z�������g|]���`X_����Z���]Ӵ�4� �tp.&GV�5�n�@g��D�7S���A�Ϸ���]2�.��`��˫�Q˵�1� ��nW�c�# �lq�766da�C��Yp�y����Aѥ����#�ߩ�*�[��C�)��:�e/�ϧO���{w��ͭ��SG��(�iIT�B�'��f�{�t����Shp-�#.�
lbKI9߹&�@#/e�qQ`3H�bhg�o؜�b�d�u�y��&a����:�ӟ/;��U���W~&���7f3Ǟ]`j�����$z���A����?��>��T��� �ˇ�0��}k�[6ά��H#N _J��,2:*={��E%+]_=g�!�]�o�qH��u�gH=�q~`��L��D@5�*~j�Z�&�6V�p��٥�9���X�p�C?y�ʶ��^ lIP=��տ�'�r ؠ�����(�9`�z�R�&���l�DM�H����V�&n�J�d��]��H:L��2eyyL����d(���8/-m����,����?�$��������E59�N��"�v7����F��F�V)A���tq�R�[&���c�^�^�o���ٚ934�p{�@Ș-eT��i`׋�TiC�X�+Ʈj��o-X��S��
vE	I�u5{I� ag�%���{8#2��A���.��P� 6p�l�A��͠j���!��2.�pe����dc_��u���x���0�O)/�[����)W(��E��&���agjZ4`��pqLg�ʅmz����=v�bs�b�QU'��ut6l��=p4"K�r�����=����[ܬ��Xx���.--�5S�j�BM�h�$[���1�	�d�x+�*  �c�M�[^Yfz�q�xn�+��lLf���rx��$�+���j)��M �D��8���q��2ZO�Z�/,,��P���})����a�,���g\;�5&����M��5/kk@��#NFM3g�`�����U��}\w<����ol�g����ihW�[��W;����7������{f{&౏��S��Oy���l��Qj�_p��~g�'?Z0�jil��<e�%[{�u)������g��9Rƹ�zT�[l]+"u��_e�r8������5/�I�k�	zk����&i�*\V��Ź ��K���!�β4�BJ(�'�;ݓ�W�eo�Y ��rtzF/^�u%SJT'��P�{�!�'�̕sXv�&=���ɏs�֮aQC�oԖ�i$�a�S�pp�Sg�N\��7:��aX�r��[��'�k�,Xx�=N���)�Ί<�M ȇa�!���ye`v����rJ(l�
��	-x�A$я|b�F<�k���҃kB]Tq��D�}�>��� �8�Ұ�������h������Y���>"P���[64��6��5�A -�8�`V�^�V]�;t�. _%p��-Ea�L=���JƠ]��ɉT��F)6�m�}0(/���}�'Ӊt��1H�!�e��*�9A
�p�$���u2Ι9����j� �z#l1�j�|>��ۙEX��A�m�Q�b2hB"�NR	VW�e}mқ��K�7� ǁ�=��ի�,NX�8UUC��
M"V����(Y�Z5�HA�X��8>�&vΎty�a��j1���h
��Q8ƆC��ll�;s[��2Ϳ�D56���ٗo��N�>
�?���#}:�O�GP��5�pb���Q����T�G�:H����`�څ-���Q��������i8Oe���EE#�i�Qw�ˀ�B��5Y�낵�x���~_�=яȈ��U���]�9���������{��k3���{&����҇�������On�\����e����J�n����Vi�ϲ�:E%�8���geީ��=��G%a�9�u��p�"B)l\�li�il37�3�o��M�����y(���d��"��|�nwC:�d���Ԑ/Z1��Q��~�T4������`�p0 .WZ�Fo��{��G�9lg�.f(�֕`�q(6��|sA�5ټ#B�㲬o�˝{��֭������a�<Mmw�Et�Od?\3T꟝ة+n��•aa��`�cgx��Gڮ� ����b~�=�b���W^�9�51s�&	Y8>��$�W�d��邭���!I#e�~(�3��6~}��A���V���Q>v�zWU-$����Q�s��V�x-t;������{{{rvr,�d+hL��֌`FL��|����+�;V%��2� �/�H5�Co	�/j6�Es�IpP�./_����� �Dh�]���A����;����t.��4��� +[��ŋ���K9��___#�ð�4 JF�@�JG����v���V�\���<�4+ev��ed��֭`����a�B���9r\�=��̼�cdjfj%Uʝ���cS��Zeȱ^S� n���W��T���zo���Ml��=����:����Ԫu�cRg�Ҁvs�9���h:��:fpֽq�*��/����.���}���1l�c*��>7�^��vlވ�.f�.��ҟ�-@^���8~���ÜzEVpV����Ĝ.9%���e�pN_Teп��D�X=���x?�|_�F埈�b�Z���@G�gd����u{��4x��(*���+�n����$`S�Ҩ����}Y�7����"הb�)kt�$[uY^Y���{�.I�#Y�#"ufi�U�D ����{������gg� ��P �V�eVꌈ�f�7"2+����P<8��N:�5777w;֕�A�]�0@�r�N����K:��Ծ�Y{٦c��*�����1deuM�4��])�:�t�s<��(��#7�ޓFs���{�,}���Ud��H	���o�-���;�0L�����Aa��O�e�d��g�~���*��Ե���&WR+ބ��=w��M�þu�J�ق�� O���w_���lH𚪦3
�ժ�.'�ؖ�f������2[ռ�"���
}�3�̼^%�D�ݍ�y��|�����'2<����PkR2�`A	z�Z^7^�d*��]��6VVǖ�zT/e���0:��ę����$^��� Y6��'�J)P��m>|x_�<y�ϋ�s�E \�_v����\�O7�8g����3���0�F�L������ٝ�g��;[k�E]�x,����S��ޚpxPM˧������q�Ι�I�<����%2�(d������-;�;TQ��ϕ�(���qo5y5Ql��Hi6A��V��A���i����Cc}̃<��	�d0��*����ӛ��HIm0!����&���J��&�ȫJn�&���y������e�w:(Q�v�q��M_�Y)��� ӣ�$4Ί�.�!�-M39>�
�l|��K�*�Ϛ�U ��.E�;������{��6��H��Phdgb�}9��Y<Z���&�c�b��E��X�2�N	�%�9}���7+
��)�8-���eBV-��	����h�ܦ�We�;�����'	��.�������`ZX��[�xA�?p�@
�JֱH�i�$��h�J��8 S^*�X�'�M�߼�c�F%�?�u.�E⾻�{��9��K<�	4� �H_b"d�ǥ�[��,��4/Z���ɔ��?�^���h!�
#�L��,��0�� h4a�f�ive;rWsT
��;e-D`�	�9א�۷dmm�^� &[[o��B*�e�����ek6P�ԐF��47�1u�#z�bA�*&;�La��Ùk��oc;� ,^�V�ݿHɏ�}�K�Z����`yK�c�����h���e>�����K���m�,�S� �}֦&��u<ۇ��Á2�`Pv1�h�ͫ�a��0ާ�^c�2 F����,/��-��� d\�uj@�Z���BDd�V門m�o��ʱ� ���Fr|��~ʋ� *9)W��,�]1�)���;ޑ1�v<�m����=�g�b��<~��'hc�;������)�b��fW�W�|Ay����&%9�F�$	1k;p�<`{n�\�Md�-���2���~��c�b��v�������Ƶ����R;:8��՚���ew�5x�}Q����k�}�/����*���٢��������e�t���������ټ�u��/����dc����<#�a���U&�3Y6����l��Ϧ�|/�A>�y�I�=���������'Z�k�ϡgd}񬲮��zP|	a�s�׊<y|} #���<$~Ȟ�Z�H�FԐ��W�ku2Nm��B�
����.�'+���M�}�(&  ��Ra�&s�Knp]�����b:pҳBV��Ur&
�	>��9l�~-��;���Ɋ�R�>:�[+��cuw�[�z5���׈�pkpR���ښ$������f_�Þ�|,�Xg��	�{S�Y��m����t��b�{�V�~�ʚ�����m��;d������/?�ɏ�]h:����U�]-h�3�u��@൨M�6n��O��裧l��٧L[��
/-̪�������Z�0��j�y�S-�l��� `l��F��B�?�ƁV��Z,��);����D|��9 (����(��ʩ ��J
�w��Lh+�^-�@���?�Ё�9��ٕ/��B���lr��^� (��ۛ����,�_����}���rC�W92[�,��C���L��EƗ�c8��F�N��[�l��hhc�rI��SZv��WX�6�%i5�9GL�t|���� ����0�i�������;��º픤ك�d%,��Sk$���w�":�X E���;�8ck�ؓ��4����Ҡ������o�1W��W�U�l�|ڍ-��F�
e\^b����ZGa�M�yH� H��b�[ ��Qw<?7�}�rv�f�=��[��$��,ӊVa�Y����x���&
�/��W	�߶�����wW��M��.�⹜�F�a�������"�=������� �E��Ɨ����w��2��Ԁ^xr����ҜM�v �g(P{D4K���|7�퉇�H-�:�6��#Ź��%8mf�P8ݗ &�Q涃q.(8���2�%- �.����
����`��V7����l)L���<�Y�p�!5��	1J�+~?�!m�Lϭ���߯%?/b̶�R��Wjڳr	�f�&��M=��F���`r=ٝq�#0Mu��[p�o�&����1�ظ���
�drJ�[[f�E��b	�t��t�,~��E� �\�*e����W������?$���*�������Oh�s״i��)��,,�ɇ~ ���/��~�Cy���'���P���KN��uQ+�e֢���ܖ{��;P�A�{�9��R��=�W���� *�SF ��,��J�d	h����]T�;�"������i�q�6AR9��~�ƈ��H�.m�('�6�$���ڊ��M�w��,/�X�:���8�Ӳ(6RX���*{���Nv�*���¿� |Ѿ��l�$$��Eu�A�n ��kp���W��i�x0������4�):��v���D��XKl��%p���M�=g�E���F�X��J�1���mb���eb���B������@��Ô�<5[�q2RKJ^�Kf������D�I�s�w)�����V�"�x�� �+Z[WY[P%�ra&���Q�KLXTg��X���^�Ǡ�@��2�f��Ň�R��]���520[�����8o�n��2=v���m�4��Ml�:�U���qO�g�ݜ\�����������c:	����o�N�~���S�7ML2��.t{�����P���( W�S�i��2�yw�٨��������2/a�ό����~�	˻mҵK�f�/���(�'b�1d!�\]�p����T�6��V.��R3C����4�?g��w���h�D$gu�5��9.�����+(�赐�V��4k�e>��]����M
��՛ިj��wr�6�� wNp������Fq��5��^���lQ���O�'?��ܹs�zDL�;�۲��Ǣ�ݽ�Xk��}��{������_���Q�;���c2[`8ն,�  R� �w�l�ӧ����mug8�ȆnnޖUJ���,4�����:[����/�����>��֛7���+���Kv@�悸�RU�벾R���4kc�W2�L�����.��#�p*���Zuw��n�q_�s��1�5}ks�c|���Y���$碢1zV������v�M4Vu�hk&���ynY,[�j\P�1��:Q  ��6+f�&V�˱v,��{�xB�[�_�r�AW��7����i�f��g�6y*�H
�;2��f 7��l��H�tNI��Ԫ��M@Ue��p8�FH9J��ۂ
��ݔ'|��l�Z�8OIR�����qM�\3���''�dmـ��H=�aٶ���1ڐ=��@�8&��"H��e�2K�y�g��X�j �m.�`�"@z�1^t/";f�{�}�!�<Y\����;�.^��3YS�_T\�ϋ=����������*3���$oA������_����$���IL���$[+��=QC`�=ජ�,ne#��E�z�:�ٕOS�YG���Fbt�z�l�,�¨d�BaagS	
/ �p=y��dĂ#3n�:��r�D`��}^Ý�� vn���\7
m"�ϼn���*�R�5$եgm�1�!]�.m} ���\�f�>.���v�Ӆi��WY���o���@fmuM��{ O?��d�.���5y� ��c��o��+4��u�޽-��O�����������͂,�V�XӁ�Z�N� ��`��7����cj���g�v �� ����O�}���?�^��'߰a��ũ�z�R���?ʳO�"�'C�BTS�:���e���u�������ݏ�@F��Vy(���;rp�v��P�U����2R��`VCyJ����Ae�����!����� �8;;s r`�i?���NU�S_l-y�=��y�R��a�ף� Bp�;d;�+Zbcf��!a��~ȉ)Ό�u"Q�V�|^��`�yk՘�U�8O\蘞���+K��b1%.��ݿ�V�V���D�vma<���i��8�t��<0�tܕ��U����b�r���cz����0����� b��ʜ���C���k;-x�kKdؖy��:� ����v>YZd/�)���\���G.�z���-d#x���w���:V��ٻFh�Z6�i�
`�����: ��˳��E�uz���-.�j8�ʱ]X���=1`|=�w��di~�;:��Iz��S��e)���6*���~F��q<C
q1��2jo;�I�8��� �2։x��/��HUҀ/㜠�dlQ~j�6Z��/�zj~��N���50��<͋�JR��������,�}���N��S�������]�4��Nџ/����?:�!�\.c�͓՝C�?B&�-j�iQ��A�u	~t�0�V$���Q�4S��]\n2y�nq=oc
��ݻ��Hn��뉢H
��B� �4i@���9y��!��ހ1��c�n)�z_^^t�ߓ۷7�Z�h��H�O%��b�HF�`/R�Ht]���zK��X/��+n�hQ-r�oK��ut�dx�ݳ�����2�ޥ����s�;/����T��@�~tO��"��ޗ�A*��D�H�S�?hL{}e�q?��9�C�Q�W�Fr��-��E�:뜲���YT�րEa��2���b�d��t��51�� l�*S�0���k�4.�	��1ґy̆�§a�����k���:.$I��S�W�`v�'�|2y@��|>�xf&(��sA]9k�m�v>�eq�� �	�pm,w�6n-�n�Y�����]`��w �ov�`�X��n{��\Yi���!+�r�72Q�O��\쁼]�К�`,�c4�� ����:�s�{ l�0���xڴ���8`?�LN����3� ��|�M$YS���r�N�]���\��Β'���E��wx\v��E��%
�h}���5'*,�nR�:̥ٿ/�Fa�S�(����~��˹�~z�����(N%��/z-����!�4��F�#���<2�G���6�F	�0`��T�¶`A��N���(r ��&-7H�Q�`��Ā����+-v���[|�6U��{���D��ҥJJ�%X��� ^*��i˿�$С�i�^�j�_a�f�9dw�gU�ܲ)���oa�*Н�M�p�]^�*%f�=�2���ݥ���p��nV�n߾-����^��勆�酮�ѬR:2�V�rl���yk��N�b�=�%��@NN@8�ۛ����{�A��p_FîB�h0}1A�X�[C��#o��Qw�ysMN��}� ˋY���B�"����{�)��,��`(ggn?��ޟG1fÍ78�Pv����U�Mj���iD�����`ڸ�B�y|�� rG�OTZ����U��j�ԕO���������8X|�;=���s��O�.��u
X����hO��}{(�<�ŧ�e.`ß8�g�ZfH��ڼ��u�����x��o*5���dg�}� Jʘ��w+�+�0y����Y���ꦻ�6n-��ݓG�ߓ��U���z�%��g����6�YT���tU�h),&cf
5��/��y��/%m���nŹsu">g]wux�����~e��*T�f�O,�@c�ܢ�������˴�_���b�o�L�߿(���Mv�=�s�;\���#��Rܖ�[�X��O29��Q꛿\�x� ��1�_M0�!�e�2�$=�g�^�Iѽ"�x%i�e�J ��z�҂���U�n`!�d7Hh0�F��0I�Ћ%%Ֆ��I	),h�0h��e�/-�H7Y���u�JcTH��M���{d�F�H��]d.o��I�[�W`���9y��=w�{,��k5dT+�FU��ef�3 <�q���'w�:�@Lw��c�d�FL���=mT�zXm�}H�l�����|ߗ"��h0,:1�M�{ɖ����=c�]�;wn��G��eN7��	��o�ӧʫW����iC���/^|I'�U���S����qن&e�xcEG����xa; m�8߻[����@NN��Z��j��R5�a�͖��jV���AK�ZJ�^���@�J���c�� oH(����;�=�w��I�W�ӑd�HzlU����� �۷���b]=����@^��&�}�[h�{�����s]�v�Ŷ��A%�n$�('HU��d 8�~��
@0���aA����x��IL*��ep*Z��SV3.�<H7VV e2/:�#�ESu��1C7f�;����ͭ5 I�m�����2�M����������,�O1	��x�c�<^�ۑ��mٸ���r��Ct����[�{��w߄����{ �z"���҉��)���8�����z�(��5�#��ۋ)a@p�h6��h0T_�`�f=��4���R��Z��������rU��U
�޶�����A��e����?�^�rl_��7Z�E�eo[O�aE}�
�(�R�O�+��yv9_��M�_6+��b`��\�"ٳ�1Y�=%�<dOnv�UR�;c*	⻌bY�8�ݗXm��1"���ỉ��o��~4o��+%`�Xc=fZ��$hL�ݏ��F�I�Mb.���I��@��h��t�"s���H�=J��}�Y�on���;)��yn��?u��֫����vS�ǣ��?b����)q�D��bLve��d�[@&`���I@���������;|9�2q5a-��]e���ޤ�%g�FL���˽{���v��	��ĠV/�KՓ�ˋ�/����?��.Eb;�;���w>��s\���<ASo0"Yp�ѩ�c�ӓc9�ߓ��Um��Ƞ*����*�D�V��i����X�Eq���Y	xj�X�DZ�D�>dB�������*��:��U2���R��T� v��F�P��ݹ:��Y�^��&�ŀ �� ��u�����:ک}��+��d.����,����1�DĴ������5�Y����q�<Ɓfa�dd@O�7�0أ�ʀ�����
*�Rv/eщ�ƥL������2�VV~l���pN˦�#�B�م�J %��Nxlew@� 
�q?��'�`쇾7p�H�Ҭ��5��n�%i͕ ��c���3�g𴓞�C������L�@�*v�`��l�o�h6�������[vg�� � �Eo���|���c�� ����
�`��c���g����k센��&뻂> ��#+P�($��>|�l�S�j����J��援�L�kr^21{�����{X� rd��V���c)�B��Y��͏F	��(͎���p�J�'�:��"mV�4t`�7��*x��+���ٍ��=캍c`���)t�I�>��#����H{��^/��S��Ԉ�|0�Sk��+}7e�0�b �G4���h:�D � �8��w����z(�����YL!��f���7=�\��%/�ß n�}���<~�P67791���ի��QhUoT)=���{O�ȣǏh���g��	�.����#(@Gß��g�-	��8���4�rf�U��W���VF������� $%�RK�c�
dl޴��1�6�B2;��: 6����.�-hr�R)�߫���zE���{(2r ����O �靰�#�@���zömρ��]�w�VWo˭��L0%����pޱ���]%�\t����X�2��
�5@�  �~�#����'tǣ0͂ӘAi�ce!���6`38x?�}hP��?~u�ж������u�s�5	�,��}���c�{��a(��+�s�RkCt�J�M�u�fؾٮ���.0��Ղ���$Z���`������M8�T�ۜ��PT+�h�)��c�c2�6����>����M	���v�ñN�5C:��~ �2�Wl�����qYz�@��w�S��"��]/7	�o�݋�Ħ�sU�����E�1k��~��]ZR�A4���lԷ�A�:�A~�}�|�6��{�>�ɯ���}.�e�������.`m�,v��a���*Uu�l%<�`tǱgTǋj`�����	dpp�4�P�Xl�����x)���%���3�g��W���J�w��%�A=�[��.����t���G*�oNh�?R��TS�%�4P�="��&�r��(��rS*�(ꎑr2�Đ���;�q�k�����H;d�zvSkq��>�d����@[���*��e��.��U+�g-����Z]]��>�H<x��``lqO %��<@K��҇�?��^� �	����������ky��3oِiX-���.z��{C��lϠ?��� �b�,R�`u�m�12q!�v��MW2��- �l��ZCǮ�r}�5�W���bN/t)���*��AB3
-��Gu��|ρܣ���s �/����$���V��z��ޫWo���/������b
4�~�|IxiOv>��!X�8�A���$�>�z����@���H�D�Xe�'�v�Z�x�I����V0����Z�d��*�F\�� ����V!�M};�� {`�M"��d��^��QHߨc%DF�*�<�:��r�P�c�@�~,F%�ЀY��!��QE��|a�hM�q�m����Í��F�1�7q�U�}s,�9���Yъ� |�i?�9��-�M� NoK�_V�v��cؕ$ _����ae/:�����r	.|�+���fϺ�����o��5M�ϭ�������6�q� Ϗ�E���j�rܑ$������^7̟i��y�,#����~oĦ����CKwÎ�H>�����6dp˕�h�/h�b�ˢU�q=w�t��M�M��1]�L�+5�N��R���w�޷���+�%HM�7bu< j��xi_��n��FTK�;��Ћ��� ��7p�`���j�F� �3C&(�9kwP�h+���1'=g�����}�l�5Rm�����t¾�G�M�b1�u��ap=	t�{��]�8IL����A�ډ	�r���_�E��������Ng�7s����!�H�ͣz1C:����� ��jt��76~�\h+� �͂���E�`�|l��/�h�A-t{�32���]mk�JpfǇLX���`.��u�����T�;��>��q?�R�7�5P2���������������Ng {�G.h3��6��(�����7۴�"X+\C��"�t�k���x�SH"�uC>���B�z��e�|�.]SD�Fd=�K߭�,Zݬ�e����}<H� 0�^J�~�z�ȃp�
�H��5�Zj�0��,5'ũ�Q[,�����kJ����c9���&�������w ��y`?�~�b�0G�~T[�N1����9�PF7�֠�pq��s��m�;�f �MY^i��?�tda�)�z+rzr�]g��ؘw��A�hВd�~D��${Mi_�M��]o�*���q_��oK��u����\-��U�mwaN.]{Im��򔜭������Z�A�[ߔ� �Z��]�[�0�i��� f];	�U��[���2��A�ۿ��k�L�3���u�Q��8��$@n��j���-�`���Dz�J�B!��(%�+#�Z�60te@+[7��|1JO�b.A������Q��`�u���6�)sz ��/f��T��wsI�^X�!2և�B8���-��.����Qt�BB�gd���-I������L}�Is��C�oׁ^�HwϮj�^�����Jz�IcZ���5 �`'ἀ�h�3@g��!+��hH�l���Z�l%�.���cy��ܹ�)��G�z�)� ��$����`�j<�O��n��7�K��r�|������@vw������,��LC�� 4��FMX`���z��S��}�z�-'gy�rO�vܱ��BGN�Oeq}OVַ�����7ۻ��w"{g���7�u,�:/ ���/���x��j L�J�Ҫ^��������0�� �+��v��ޭQoh+^�.�Ι�+�5hO�8��G����.pұY_)C?����c�{Nm\,{V�7� �j0����5�-��KV��� �  ��IDAT�`�����a��E���(�l�2IJ�4k/�X̀�;�� ���h�-�q]�8T�X+�Śr��Psn�w*�>{�,���Xe1"�#w��V��?�x�͊��C�w�G�9::��㶜�v�~�Ujc���[�1�?���!ZZ^�ͻ\����VP|�׉�;t���MN��>#�yvsǎ4;'��zyw�շu�����Xn�Rq���|����p5F��&g{)E*�VyV+)$t�����t㛃��}-H�P�[\%?�/���2�p����%�q�����x��$�m�𦆪Uڐ�q�z70�1��M���?"�Fc���`7,Ռ1
�p4�;����g���ǥOS�]�pVv�z�d��TZs܎��"��;_��`�����-�k�KOl��z�t p��4D�7q%���o��=	��f����P2�xl Y9���Oe���ߍ�؃0u��� w��*�4�0�]�� u�㸊����{�_Q)���I�0��{�dss��bZ�v��پ|��9�%��7���5�VKr��y���ܹ��g��@�_=�S�j;V!�fb�X`)*�����i��`x��@�[�^��B�
o��}�nU���e$H�E��B˨�Zr��g4���d����w�N	�j�]9p�wO��V9���8�{([;��:P� �JS���w	��z|�!�h�������XGq[���ďck���7dk�ʘ����D6��*�t�Y��ِ�%އ�t`����VA_���!�(��N���5w�N�!k>�J �Ke�8�E��1@#Z��WW;������6�sNHHeY��� �K-�v�{��BƲd�KQ)sm�ma�)��Y��$16�dr���E�-�w�7��|�R>�l�b�rIY�5� �[��dn��H:ݱ���V�c<ᘤ4Bs���h�"&b؍�c��w�?���;O�{v�����]�7H����T���m�c���>�F�T�q�\��a��6.���	�&+��/��8,h6]@�f����a��ڬ[+��$��NLd��aXC���D���7.*|���٦ȓ��5E�V��!P�qh3P� &��u% ' ͊~�Cv���Y��&��,.��}��b��[���ut֨<LMw5�dI�ҊR��L������݄�"�������4j�^���2�Ad��H��\f�<���%ow9�C~A5s�B�!*�G]�S�ㆧ%Xr�_Ҷt)�\��=�X�640-��^�+����9
�ܪ�+��Y�~�''
X�z ����*���Uoϛ��FdzP���-V���m��ş�s�L��	%HRq��gQ����,`��]y���������j�W��/~!���(Zۤ&���Ey�����e�H����� JTky�p�o�Wb1O�ہ����_|)w��"���o�9=���z�D�
��
S�j4)�!�H�����: ���K���o��L��`0�������pВ�\S�æ��C��Jí��F5�<�}B�Z0ph.X�����&��R�J���U�� �NLs�;����\��?O��K���#�F��S��R�r)�N�fρ�V���z�0Ўp����ˀ��Ve1s��$�YQ�������~��_Wp����z�
�c�/�S��v�Pju��1(�}�C�a�Y!>�:~�y��iK����!�9��iwe{�%ІT�VՉm8�U&�b��`�֗�0����h�(u	�*Y�nHl�?N>;�� DHl�0�DZs�`n�֛m��ْ��t�tҳ�mh�n2��/�)z�Nۓ�gh���ʶn�ܴ~`��V<��$�e�o2&�T+|� �������2���T�fgÆl2� NХ��-�(=��O���@��-����<����/~�Ks���jP̼O6� ٢Y�5H��Q �K
�T���(�;k�M*�hX�Q&ۓ|L�N 0]��T&�j�G�j蝛k(��D%W�'MYXa:>6��4}�����B`�Q;Y������  # �XT��ݤP*7��1�~����9ŷ�����%d!��-j݃�fE25-1sj�RKu��J=h��������*��	X���A��Q��
��fN�Τs�VQGzS��1b���&gc&zu��"�;k�h�7),���qZx����s�U`,���_������,����.�����n�%4[s�� ���%w�n��V髷2��R�����t\�zJ��X���GW{��_���yo����gR#��z2��+u2��d�AB��U���PT���� ��M���GGrvҖ�d�W}��+�,�J՚/w[z�
�H���:pH�����ś��r1Е"-���O]<�X��P[�z9 8�C]-r'/<��2�Y�{Ѣ�=_��=>>!��9���UH����UL3�0^�Áu*g���fPr��j(ު�م� �9�G���K�zg�iCk׮�s:�s԰`�Cg������_X�d�1� p�āmsB�����y�zK߁m��F�]t���o�d��|/�.�}�Q_�m����\�4�}n��ݢ���0"؆����77ɵ��gw�g��\�u��ͦ�x���w�r|z��Zm�N�a6	�)����e@�����_���� ��,�m�r�c�:�j�݇�,_������s��֍�|�%�R �<�-~�o߳����q�h0��<����+����}u�M3���}��m��]��|�t��Ԉ:��(&
�/�����,dCL01�ɨ���!�����Aaá!|v���81͈����u�
�i�E鉲��lt����V霰��}$-X���2�	�xZ`yM�����2}Q�Oŝ�8[	<t)���8
�j'�W
���њ'T[#�z��&L����^�Vm�Y�zk��r��;��r(G��rtܦt�PR��w�%�*)����6���ޗ+}/Q}�Zj=h_��><j�ϟ�o~�[����@v6`���?O�Uw`��lj��f���H'����`�	'��Ե�9|g�.��? ��6ՄH��
�F��__|��@���T���������z�ZS�+[�&Q�'�R�F�����UE�%n�$>�^w$ÞV�S�I4'��T�/��Z��SwB�\!s�vm{e0 ��%�Z�X`Kjq�S%Y��p�A���Ҏl����n,�ؖۧ�~d�q\j�K�U���Ρ�3��Nc�F��I���Q6��\P�Z� '4�ew�p��� ~�E갡�X].���S��(K��Uъ�V�W��b�.Ƙ
�V'�Ԫd�q�''G�xC��I��Gu�O��`i垬,/1H���e���[O*ՆH���m�����1[?c�<��V�k���Ȱ�'D��w�u��Q�r���S�a^!=�hc�Ȓ�^i��zV��E�j1�~��VR��]|'4�_Ӓ�D\�<P-�F��-���Nu|I�dh9�~MiV�f�$�R�[�9�`z�u�������ekc%d���`���`���� �B&@'�4&h���[l�=�a���ׂd���놴2e;Q=+A����[�*������\��X��	ˠ� /cx��2���A��ġg�8�݃�c0P�6����z��.icv�b��Wwmh\�J�F�]�oČv׍Q�e굧����	}����u���gd��@Q��������4[rI�t���E��֗bz�n��,苗���ߐ�?�L����M������_��t���ݗ?��/���F�����쮶��M,���n�l�'�|"KK��w~��3wͷ��暼7��ű,.-�%@n�͖���H�R�����5��r/�y�;�WkSJ��9������ I������� �/K5x��y�w���@�uP��\������`�/�6�n�Afz��v�(��c/�����x@�X�fW���ڲ�}��1�GR.��rd�WH��1Ϛ�Z,�/�k����rtk�}d����82B��c�����^ߍ��nW�0�7v�KU�CG]�F�}n�^k��Ϋ�ձy�]�)[P��:ٸ�
�-�K�����@CY^Y�;|���t;ǖ�	L�g}���^�(k�jg�������H>��j�^t���MŤ8:>��S~�L��E�4����|�*�I���K�f��-����%�ٷ
����"�_����$V��e!�(�ջ�oK����ٽ�1�ƙ/�{1�/0�r릘��y�&�� /��(2[g�T��@�VFu6$���ӣ�Q�z���SI���"ı6����R+��\C��rr���e���-��8��� Ɂ��6�dd�������)].��EG0��	xC���`����X�m���Ô�mS�D&���X{f2���Bc�&��Ӷ���u��'�n"�6��$�~00�Q�� ��y¿���"�[�����/��r����x��ujb��r����O���������_���-i���"�\�gN��j������ޞ|��39>9������QO����w���Ф�q@vk{�����y>A����G9�{?xJ-+��ׯ^���/����Ta�{	Vw,��NT���6�I�nk��Ra}N���č5�t|&b )�#Sn�b��ۏ�@	��h��2�� -b
5��0����	��|��v���2?��貭�P|Q�/���@��%VDJ���!���@�K������@rL��u���O�ѣ(/�*j��1�ߑ>ơv�#�'��BVz�F��01�u�q�(k������;uHQL�,���H��-��w��
-�R6"��yh�\��������(��V�jI���ȝ�J�&}w�������s��aC���?~��*g�XJ�J1�@b����Eu�ݕ���Hz4�g%7_4�1��`���2����k�1�B!NP�q��Ly��o��o�~Ѣ��W�Ƚ���RDd2u��%'&� + LjEb�<�q0�Ս+֤�B=��xnB�����@�銳-S�*�kk��ܢr��2+G�tzM{�$BH��1��Ϻr�&S�9��(�P� ���8�Yj���#ɳh���^i��~2�&�5p���N�]s�fD��s�����k.��E�b�Dl�<`W�a�-�*�W�� ��8bNB�'�������#,c�9�y�1�UL v��ãy� ����&�%�>w߅����_%��h���kr(���o�8p`u�V�-�(}�~ �����gԵ���8p|�>��@Z����/���Z[��~��0�w����c��~�v���|��G���t���.�Z�{e�����ճ]��bE]Ql�~-Z��3�pL���P&S�aG6��� ��Ju(�j��\��l�Ѐ�"�ڛݼ�
��#L��0c�l��=M�q�&dC�exS�&�(;����GZD��@6�,�eN��f���ȴ�ٺBh�Z���H,��˝Z��L�O���l�^o��<����;P�g繈ޕ�W��w�R3��ȯܛ]�u��y�Bc�qfF���л� ���g�{�lnޑ�8���5�VkÞ���U\x�y���؝�DA,]X����Į-�j�e�Yu�zO��$�\l.��,-/�o���oy�.J	fm9���w��s�0�|��T���_�A�������&��D�e�|���� ]�Λ
�2n2LYԛg��t�x����*2�6�����
�ك��B�^��J���z�`d��������-g]5p�g��!K?R��3p���l�����|��8����#Ԫ:�JH����XT.0��{��>ȿ!7_������
�ű����8�؈��^0�q��j�l?�D�SZ��ޚ*Im��LkhE^:��|��Ѱ��:(	e�N����u���=�u�o~@�����'Q���vvv&ȔM$
��J��z�����ۖ���Y	>?��*|6�5���=��Ӣ�Rx�H�?�Hˣ�F�<y��҆xCA����ShmF����,���3`B[���̵y�GsF�q0�9hf%��V��V����Hi��(V�GcJz���:��9��I�3r
�BO�`eBf4aQ��q^�mWlv\���E<Y�y�^�Ԏ-&�	v�����#�<�����%���kx��Ն�0 �8�K`)���3V:`p@}/Y����\]p���>~�r5�±a~a����ٵ��������Ȥ��3��%P	����ŵ:3@2rtr,ɗ� f�T�66�?�ED���ɩ�JZ�����>��)RUǋ9���^��a��a>�e�oV�,��"�q�����b��E�״�j:�U���Ơ˶1볯2�^TH�u��f}�u,o�^��>e��ڨ���yӷ�1AxNo�������w��&�Z>��okǈN,V�kCvd�w����� ����q� 8ϊX&.�����`V�I�f�&��R���P���4�Y���ːt|/�-��� Y�H������+�v�E���r,P�����F�G�� 9����M��\��P���&�4ҽ��"ut�:>б�^���J���i`�"�5}5'���$T�Y`�n�4�nTVWZ�?�1���ȩ��e�@�H[��3���Sbԓ�N�M�CPv�|�R�/��G�&Fj:�!-��w(o�����ڗ#+�B!�Y�Mx�:����i��;\��Ox���&�=��N11'�1tܬ(�H?Lu���xS�5&q�ـP��r)�'ʲ���YhJCk�K�,�>���W�e8��_t�����i������Z�\ώA��5��! ��c��r�P��H@�2�V�:H�1��lI����-�V�ZPV��oպ�Ś^3o���
l��|Rѭ��}��R .--ql;�̸6+��A7F�g�b+<�kh�h+�&�\�E������沱� N�EH�nA,Vc��Rs������C��҃4�s��B���L8
��s�a�9d籁upt�ŭoiyс�U��y_VVVU�Y��j�k�2�1l0���c�sU�Ӫ�zMF\�`��L9�{ߞ���C7�����P��j��iE�̹�h\�5���j�}��I�	�u�ʰ�wþ�F#Xj�]���v�I�?�y�Q B�㒺\��^ ��)҉�h�����U�,���q����],�O\��.����K��x��/j9��l3>�X�L����~\����ˉ��/S3^�L3Rɲ�ib6d	�GXLRr�g$oy^b-h��3	�3X���УS�XKY���!U)
�S�w�^�Ù������}+ 圜&ѧ<�����X׍3�-(�3TR5_ ���F�v��.�?���Y[;�g��<��o
�&#��㟩.��q��+�4fO̶������ =�Gn�D�ĉ�T"������7@:�_��^�.��p:}�羙]�4��0f{�a�Tb�g��H��Ѓ6
�;]�����!T/�� ��"(�O����N��
�rtt"{��n�9�	n����>?�ّ��gjzP�,��� wU�d��/�]-�Gv-'�c�b���k˂���#[��0P�TeRł�ܲ�L��A�^�Q�f�m����>C&��f�067� �F+Oa��Ø� �
j�#r)��0 T'�C{���i�yy�?u�/\2f�zL���1!�Y�=��bR���E��x�U�g`��A��F�a VY^M���fCh�̓�,%$#g�*�=h�eՎ�z�^���'8X�����`�c��dA J��D�M��Cp�/=t!W��Be�	z��D^v+���ꍡ�F�k41ټ}K�W���{$c4�i�����ܧ�����c� \�KZ���M_��W?Q�ڭ������ε��lͷ���{v����ȓ|��R,EY�w�5wMj��]7�o8!�ѹ�Qo����'����"9�E���Y�h�-o�o��gW�|z[�Yo� pֹ��L_g�.ڟ�u�m�{��)�IJ��M��֙f����~w%�{~C�L(���QȂexu�)�@���]�V�%��,l��k��#&g�W�)�JN�>S:���\[�������,��S{;�A|N����Y;߱����T+����sg�P�� �j�1�6�%V��j�/�9㨋������YࡗIir7`j7o�"�:F7X�9<>$#��-�{�y(�@��r�%����6�.'����ƹ���9�A�HJ��*.�8���BjFX��6�� .�0x�y:8��i�O��y��~�}v"o��eg��EOa�bg,	�)�2��<�ږ�N��2�_ӻ8�Z�][��jt��%�s
�5�v��:�����"(L}�[�ɣ!��RKMU�C�E�c՘�����?�x `w0�g}�4�%Y[]cC	��Ԩ}Ģ7�LyG�a?�eD�3�}����1
��J�� �<���0��>���	��Rl��]�����\dR�R�V���~h���~��j���^�~�y��[��8��j�c���sѝ$�i��p�Ӷ�(��p� ��J�a昀ˆ���4�-n�s�~����H��;�U�c]�;���F���Zt'��.72��$��سC^�������h��[|޻w_>�/���KL��X���б�_�>�����,�/���/6�8�O�u�Z*3��M_�q_=�>Ӛ�]���f� �����a�%
��\b���#5���=>?ƺb2���� P��.�:?�
 '��[O�Q�|YY���8�"��ll$O�����g��¸r ���YL���|�_��D�����}�m�~�2-Y�fy�Sn3W�v��)6)N���k!P.慯����[��A3�RG#�r�V��e��Pӥv��zIno�ȇ�?�;�w��n2:xg��Ѝn��/���7r|���&4%���43�iN��]OP(���Y�?#%�yMeL��¬5��� ��0�gS�?�BD�K(�IaIԑ��3��e}�퓴+�t��D䴭M	�Wܲ�)�n9��Ȥ^;4��r�%v��6i��ߒ��5��k��+˙��~I���J0�%�՞�D��j�މ܏���qOڙ�ǔ/��=�p��j��l��%������X�dBj9���I�F����T>�vWh�)RkVX [�`vc}�W��x|%�vb�ްA֯<�]���դ����T�'z��~pF�t>���eNVWkƀ&l.2D!��C��N�T`���W~ ��2�T)��ş����J�4� A+l����VK���Y��6�����l��:vh��(
�X(�%Pp5uC�z20�>M�B-��Alm�m�����ۙ��>2g��Ǎ?�@��Rj��@���->�&c���Z��$Q��V�I�H�9�}�����dN�q�pN��U׌�r3B���5�1Gϕ︈�9�'���(N�8�TeyiQ�ݽ������S:vx���7���}SqAs�R�+r��]v�K�ޓ�����:� �0&�j��Q�'p@'�*[��u���C���9P)��VǍ�\�;���mdq�$���^�v3���'R��2I����}Q ����EnE�T��Z������Yr��f���L��Ϧe���6�}U�M$p�`���^$s(^��딌X�؇iv�2�L��K�˚ �	kJ��H��-l�bamyN�֗����#�s��{�V�37ϧ��j��;oG�x$_|�R���?˗/^���)�E(4� �c�(�=��yL��
$w^֚Og�W|}D![0��P�}���J�n�[^Y�A'����uew��^��1''�����<���3!b�����3gKS 12�l�/tU�� �K�:���,�Y{$''{�~��}h��
Tft����o�r�[���/�#��:�,4g��w�?t��]�tGh-
�"�$ ;f���@Ӯ�\I�UH��5@@���g�+�F::~+��z� �^��ٳ�.C����̰Q�c�KZ#���R����\.�(���毛�q��@�mK�cJ@� �-`bAqPܓ9Y��?�%��[-��\Խ�X膵�-GG�n �jsQЊ� W���'��FY�	�����۰l���q���|@���p< $hQ�	�wwQ&��w��,�K�3e_V6��p�
zGY�T<��R
`Řo��3��6IV�V�k�5b��(�m���6�H,@Ӭ&��X�`a����5�'�b�l�4��_��[k��B���_�]#�@��,1Y�vD���7��:�}��`u<0������cDН�$
.Q<�.�H�#�ٸ�N)�ƭU7��L�����>�W�^�ՁcC�^�U������H~@�wk��26�:Zz5u	�̊�Ȱ�q�8�j�8�7�[�g,�9���&e��6�x,.,�`o����40槧�BM��u�0�f�4�/��5��R`�Y�iv�3�W�5L�s�ߧ5��c�e���"�w�>\��"��%阵��sq�qLK��7t��z��1`�1�~�I&�;w��䞝L�u�8Y�@�0]b���ܽ�"?��G�ӟ�T�=x$�֒����,=`e���t������	͆n�@��S�fl���U#�Rɟu���sѾ�,_zM��+oDB!��YWI1F�7�ɮΎO:y�2.2�ԚRͻAx��S988v���M�82|�`6�J�?����w��i��Y�t�^e�\
)����v�Rw �Y�+�p���ؑ��=i4�dР��^og3��n����������"H�� �hh�z��7����YO��,we�;cJ�9����+sDf'�KX��''������mط��>�P�Rm�*�0��~��M�G<��&C��d�����,��?M��6� �����'��?��#��O~Bf]�����_��o+��qr`�Z�H���,���  �|u�}��E���������S�]�wa	�t�EQC��;�ɲF�A&A(��B6��з�f8�xŅ��`�p�#}_)��Ύt�J�a��D[l�S\"*�:����V��8U2Лd�����Ih����^f��	��N+0)�����iU�����,�-�34R�K�^���9wݾU����g��{ w�vMw�p�677)m�s:�����',��Z�`�|�c�uX\��{�D>�S�����A\����:�� �v�d��+`_�1�@����c�e{k�m�B��FsNm�$��j���RA�w��"�����ʑu�D��O�tK��������B�$<��(��ɻ4�xL��>;e������٘�X��42�b��,�u�XĊִ0s���9p4K+�����������m����n���"�|8�\�d�z��6�vֺ�p�7��)�f���Jg�!.v�8.۷i���M��`�/�`���O�/
FP�bg���K,6߬��ڦ��g���ǟ��|����e�J͚��Pg�����<z����{�D������R�&"�~\�S�
�M�x���*��XT�acB���[ [f��%*x�J���� �����yȎe��-��G���(�+��y�C��@[ڦ�),��i\n����}�=�1��I�"��G��A���lm��Vu���@Z%eL��A��jE'Em3�+SyNJ�o�h���N�)O���{�ڧ�݇l���پ���0p��EL ��e�d�&ޮ���Hg�s����^��n�죊�s����255�<� �n�{��S�&�{y�Pݸ�w"�^���aX���l^��?ɋ��/7<.�D�����%���-������R�܆p|����������,��t���%~��4�ڐ逵��!~�T~��_��|(wn�6��X������{2����?���ɿfRJV�� ˁk�v�HnN�'h��b�������jIU��;��d���
�a@���Y����{8Hۣ�`�����|��0���<ا�I#_:1�B���,�+������
��_�~��c�=[ơekʰ���@�"��p�8>9֬R�[{y���`��/aP�@�ZF%xK��6
fqss]������{�!À�ڝ0�p�s{Y�ݻ%�n���\���.�Q�RjS��/^����_�A�A��{$�6��J����@;���RģS�L��v��MH_2(b#�x�P��z���>m�}�Hk~��\c�o(k�F32C������S�����c3�����[�9�Π�L�:>��"��5��jx��� =��j:�6�s�V$5Os��YS����y��k<�� �q�T`�3���}�������/��L��a����ǔ�-Ӏt���4�:��i�8����3�B��(��o���������?$���"�W|Oǉk�C�e���p���1d�?wi�Ng��XV��>JI��-H�qlY~�1�'���}�ñ9��UM9��L��r�%KKu����tE xx,�[�?�lo� _�U�,~JT$Y�x�_޽'+ZS݄���T|o�PV��dqa�M\�r|ڕ��=wZ��2��(v�g���|;�
v��2�N�5��[._r��
�S�~��!|wOd��粷���l�x+1�$�f˭�"�q���������F�L�>z�:�LO�pేҷ�ne�� J���(X9���-�0�v�>��D�V�ɻ�����#7)���ng}�R�ϱ">NG�B��o;�3�H9��V	d}u�M�MM��Ff�N�K�C��I��ɳ�^�g�o��~Gӛn�8�S�`�����\�L��t�\������/���l20��H��Ž_�����~����?��lnl��ˋ���sw?����m��723`c?��c�߿������?d}}U�@�wm6�9`�,�=���B�x���|<�Eq�̵V����w?�;2d_~�%�t�ZY^r�rɽ?O&���cKZ�f���Q����q`���W����׿�������}>���Uw*V�������@��`>�}��{�1�K��� [�����ȓ�ޓ;w�r�q><8$Ȇn�C�ٔ����֎���|��'��Ȧ&�U�2l�hA��" �h�=��%�gQ�x̦9Hѣ���ڊ��-��SV���A���xT�:�L����A��R��uOKaM(����z5b�,fc�m�M�&��#}w��B���0�Xp��������Y��� ����vQk���H] 䂥�/�T����f9`�1V!-�0�p�ލ�Q�u�UH����Y�/qZJ`@"���)�������� .M̛8P)�aߴ�)t ��:�)΍���h�ޘ^����!�w,4t��C�{�YL!/�y��3-x6pܸϋ���,~4`Zr�z��ⁱ�+@.e]�x/�6}�
����af�Vd��_����6.��{�k�'8:>�yG �s�[��L1������Y�u�/^t��%���En��*�33>,na�#�8�̸<x���׶p,���TR`Ǐ�5�XT�,�x ��@�%�wwE��?�X�ܿ%a%d��z�4��KC?�!�,Ck@��.�ZC<�%���?�	�O>��,՚�̜��*O��H�$3-f�ra�Y�-�C֜$�sKx9�����`szz���Tj-	�U��pg�H�wZ�qk�d��xD�7�vP
����]w�ȭ��X���U�_\u�Um�D%������'y�ꥬ��ee햠�N��C�ۖ~•��X�4ܱԴIE�m��;J��[p���lG���̼'�UHra����������Gnrs �4v`7�FU�;�x�9G�댘�æ�di�4�B�1G��$ph���l���Y�-�3Z/#]Z��B�kf��S4�/Uxn�5{��y�j��daY��� �`M��@��'߿�0���������o�~������S:�脬^�1'��[LsS�k���`^?|��l��[�)��&��[����S����K��Č@@�ٚ�v�ӧ?���/ts8#;'���ОԮ9�Ѝ� +�z��@.��+l������2m�ķ��G]�% ���=2�K��Ϲ� =�ԳF�����)}p_�_UG�Ӛ<��(����X���tq�3E:v����c��d}m��
��/p� J�%�9$`r;����;w���'`��C�M>RKG�~r�ۡ�E�@����:8��6܃��L)TVf�&�Q9eVGus`�S:"���#%���	�1
�(�0�8��������j&M���'D�8r������$�]�Ŭ%�+����i��]`�ܠ��1�ӡ�E���<z�.O�"��#b��6�$�8Nܹ������G���.�{x��\��o��xQ26+8�Q��v���~-�}�)Y]��Ƶ��8X��{�N諑��<�Q3�>ӹf%��}��2����n�������.f+~w�U�EM��ܟ���]6�u���+f��� �*�/n�(��>?�\޼y�1
A���y�^�� ����-�h�/_���@���_��}˾^D����������y&j�~IS����C��Q�w�R��c��=ؔ;7�9W�;�s�DЍ�  ͷ�{9��1�������C7��<�N�/t�}����Ė�r����̥Ţ~;~=�c�jWY�Emzʪ�t_>�t98����`���ޮ���*������Xh���]��*[�h90ZYp�Қ���[ϒX�8M章������
�O��2���|)�ϴgm΁ ��|�Ԅ���VCZ
�u����?Q0'ZХi?���)��Q��lL`b�����=�^��p�]���ڗ��9��=�����eg!7���iDU�,,ߑ{?v7�"*u!	�1'G;d��^.;�=9i�٭���@Ed9�gk�Uᗠ��C��w������ ��͉04ɇ�������]^��Y���te�>���rn��$�
�C6 ��E�,<|�P667$���Dh�����chdO��ٍ�L������K�=t��;;����޶&�P��G�Ł��ei��g��,:�����G���O,À�@��~���aL�=�޻'�V[����Z��s�տ�b��������dum���� k�)�����mw��8	i��o�Qv@wY66֤垳W�߸����や��hC�&���G.���˗/_��Sh�#��3Nri ��A���<�բ\� TW)��%��(�U�sh���G�N�M<��%�z^�d�w"^V%�]m�.�
��5Zhi F0�� �P<���DiM\�å�>f�z��\c G���X��ԍI�!Ʀ�,̭ˇ�ݖ�O�|�x� gۍ?Gm7ٝ�`�����yy�����?�'O�����UV�I.���CQ��X'�ڧ�����>��Y@HI@� P=����� ��f���΋�΁� �(��)�h�瀚��(>�ә�Yl�g��{E��ĽU`>�P>�4�=������O�o�P�?$$�ŀ�9)��~���8o�zF������L�>�Y`�]�ޛ,��n����� 7�(�o�;'{�^�j�9�I�B�8�h{�>�k�ݳ����۲��Z�8�Ű9�-�}�Ț�����T�\6/�\`{��]�n�gj���5�2��5�)��i�����"�N���+PF�D�R1c�@/gc�}ʉ�B5x�n��7;ǲ�z�����<S��g=:��;l�f4��R���Z_�z:�&��9KmF�F+��Ts߸�ukG�_Ȱ���7R����:q?m�u����,9C7���)'Ǩ�R	M���X�Ӊ�"QG�L	S�bX���Q6J�+��7���R4�Xh!U�`�c���%2�%��h͜���[�V���"���|[��y	��:��;�ֺl��]�����Kw���:4��/zv抬�h�I^x������K�)��ʕ�(>��V}�˷��~�K0�G�n�7�ը�-��$�h�{o����\$����'�Ǐ��� ���ە���O޼~Ŋ�_��W��1�4t�����9`	�փ3l�,�� .
Q�=$�G��~�D�~a(с~3b�_�5����L�Y�����}�*gGHGK�� �	`xw�*��m��LșT�S��e���f���)�����C7�b@�J9J�}r���?�_?��=Gr���o���:ٽO�}����٧d^�������$������P�~W�Of���`�����b܁.�d��Q��LH�����ln\I�`d&L�|Y�F���k7=ݳ����~��߽��{3����(zS��( �����ȼ QII�R�K}P�
@�{㞈8qb@C�Y���甸�Jj�Ӵ΋�@o�Pe�ƕg�����ٚ�@хR_YFpf��t�0���bJ/CA�����a�4��@���_z:��sp����EY9�"g�v��4/L�����>ښ7���"7n\	��B'i^�#JS2:�Q��$Ȍ���s�P,.��ի�,2T����������>e�*ɳ��"����>�OX,w�u~���ߪ����m�9��������� ���D�3d��q��$�n����k����1v����]�i���~'���!�wg�A��}���n����m^5�g\_n@�S�]wnߩ�A��R->M3m<1֋�&)I8����C�W<+&VTV��IY�lta��-��]�xA?^�z�aBE~�a���+N��1�@1�;vC�G:�bl�W
�h�Ǭ��g�z�)/���H6�7��K2;�b�\��O7� �[9+KK�X�#r�d�"lޒf zS� f�j��%��V����X��bt�ܵ��7?���� fQ�}�c�G{!�g���" �>S�&/��I�V�ЬN�,eC�JC�^>�{X�`���^X��'��H����f���4fVZU��R�� �ٜ׶,�+�.�>F��4�#��(��0�,�	�rt�E[��v^��;����w�o��g�#����;Jkz!�Cbϧ�
�Y�-��e4�C����AP�����p��%��D/�@ �B.�˗y�w�A 	�,�a�P�xRp����OA(9 ��+W���"����L~�{4E�!�C�<;Dy�����N�s{a;�iC�����u��Deo#��H$e�:�� \Xi�ՋӲ~���G'��F��or�LSڍ����,�|j�����̴���bÙl��������48Ϡ��l-��m }�k�ܸ~S6��e}sS���6�l6�U)�Si�����phų��EF7���F�� �"Z-�G_�E')	�7C�,�Pyƺ�1���˥G5b��?ǥGkJ����^���yi�c�x����7�9�?o�x ]ЯR�+�z�F&GG��$C��p� ���$�� @禛�9k�17'+������0N۲����Ax�5}/^\��疭{ސY(&n��x½��L4��l���]�|��Mp��"���A��� T�Ҳx����0^��b����Vŷ�ь�G,����-y.���矟���6E�k3�������G��8�����ƀ���/��/~��t_����^xV]60�&9���������$�W�K1
����Q�磑��g��w�]����Mo�9��;�-��¾��!Z@�[G��k�\��2�e�b[Ap#��s�V�a���1�C�Z7���e�}n+'���uP�#l7����x���UrE f0(^�x�,;.-� ���v0Ra!;C}Fp��P`���:d#��jS�ԭl�"� np�3����@gA�3�������G�n�D=rr��yf���6�n�c��H慶��^C��p�a�0��%����Ĉ�Ȃ3��: OD�����Mi�;��@��0 2�"�`�?��C�^dK�P�H+�u�:���j��L�j(�q�X:sQ���Hc��n��z?��4����ᱬ>ۖ�?�/_�(mg��E�S����)y�?���f�8���;{v������V ��t�|��Uǭ��c��~y�+Ҋ@� X`c� �vwA;Z��&���g�"�tC�� 8υ�v��ؠ�Z��1C��(4@-a�v���*8uY�c'�Lu��&��BW@UȚ�,,�A�dz$3S���S��6Ab pI��x}pBA�k�kJ��l	[`�J砪x&������qX8�/.����:,����+�~�N ����9�2��
0�R5s�I�<�|�3%����V;7R�ܢp�iE}Y��h`�����}1����k<z�)ʜ��6�������d$V�XVP_u[\@�/��I���ST͡�jƈU��Cա�ӆ��7�*��`q�2_s�UQ���1�`H�[���c��g�L�3��[V��Ngr4)8V�hep�T�3�� �ϜYdpc����<�Smf6���9����ϋEJ��A��������A<�ǹ�1������⤂��X����?f|������9�?�x1���ՀE�'�rc������|��7w��7�	�bG�u���:�ro/���݇ӭ�bpE*M�vc![��ڭBs��(�YSQ���J?�B����E�}��T�P�*5�, (^�$��8xOF�˪���1y�{3�zm�%u���#�(�y�bQCT=�p�{�h��RXX�R���`��GO��Ⲡ2E�&�Xt�ZD����������/"I|i�/x�`��dn�4]9�?V�!��yR�H ���C@������ueSZ��B� nn���$2:������j��$�&#�9�C�N�������h4�~3��A���ٚ�`�΀�t;�Diz>��m����9.��mF7�8d�P��X�B���F�Y > ;����F��$#�zm|_T��m��!8X�o��/zo��ͫA���F��qɟz���%\D �@M �}��4
���oip��+W/�x�����r���u��^*T��}�qO���8��L[\X�����E�`:!@ M)P��b�@RZ�&�B��ʆ�?pS�1�L�l���1?�99�����p�Y�O��F�/M����L��	@{��q�Ë�k�c�����ȟ��h���6݁��5���y��e9{f!�SH��[o^���@�NpP��?V�N�b3�B��|%�E��Y�:��{��B+��oj���,��*T�SG�f:xh�Gey>(�+����@m$�R����;��,��.��o�,��鐟�	�A?�.�X4�@�����r�ie���Zi��&Q
*����"�(NvP�G�
���(��$ܛ!�+��$��Vދ���n$5C�]a
y56z���L5��6�4�[�m���EOw��(x�1�t'�Ϗ���ދ���O����=�M����g�w&��8���I��ϱ,�[$ (N %���c���#�[e>���F��km���_����e����Q�s�zN!�i��b��҄�����0��a����:��� ��4E�"��Q�5��
�&ejR�
8](�����m�Hg���xA<UU�����F=z���P��CN�h��%E�ۙq�T"�����bמm1J���W�������֡ܿ�T��87?�6����	#���^�'����W���ElqI�@�^��Hx a��E���� aj�%UD6,�E8WmD�$��i�OL�)E���M�"O({�5��n�)�`�r�������<
�.)���p�=�m*�L#�4� mD�Z�E���T��1�^Rzg��
�S_7�c>�~��n���gV�L�
��l2�͝��/�����!G�t�`N�t ��x�˳c�%O^z{�q=�3���6/�'����;�-��(!�4Rr�9��ҢF~]1�����<��կ~!��^ ��_�:�G>۔�
�4���{W~��_��B|m*�$T�Ȓ&)D��U��0	vPk�&����wO�ik��`�a|��t:�pN-v��F�CWI���%���ez
��6����	`�&"�3��Yn�y��� P҂�ZZ�;Mtz ���]��^��yK���6��+mPNlk��X�����ȵ+�ewgWf絣8��=oܸH�����6u�w�w�<��$t���������#�6�;�eU{o���EЌ�E*̹�B>�b�4�gk -&8��uR"q8���P��%똆�|���<Uu~ D��Ұ~�X�|�xx�T�vT�gk�lа���B�,.Y\��ɣ�O���5�ۻ���M�iv��p�D�d	�N���`w����U
8�m9��x���]� K՘�{�1~���"�4
����l�~vf�zp�HA�x��t��Ժ0�JbN��:���ո]��q}�Ǵ�
蕣�&ٜ9�~�I6�U���1N;���������8c<�=�^9���'�M�1��q�y]��֭[��j׸D�2_v]��I��u��u�_�@4v��h�"�u�i���� �w
T�V�9M���~ �Gj�*u�l5�e��V��9�<�J�&�X���\R��`��H;c��Z�݊�-Z��vueA���?4Z�5�H�*[�u�]�Xi��p"�	�ȅ�<��l���c���3�� ��w��t�v ���M�*2�F^��q�n�f�u2aqfD�"��X� =3�]2R�R��A[����H�P����6�]�,�
߃LY �iN~���Ej�2��Ez�� >3=Al���=vQ�v��.$��"�a�"0��G��H���q5t*]?y�<\5�*f���١-M�"#����� v��_>�;�6�ʯ�R�7�/���+,�)�Ҥ�I��u@��lm/�7?D0A9Iͨ�(��~-���|�}���Oj����H���{r��y�RgtK#g�y�U+��7���y�� ��ݫT�x���nM�!��J^,д�jdn��n�ݱ��8�1���g��ߙj���o������V�9��%��!#ht�V3�� �����Ӱ���$�*�2�A�� ��t�Tװ�.c�`��X� N��u$�6z���:�ctg�(�8�}SB��&���L�{�H����L��������I�������������Ϫ�z�Hm��⮤Z0D�sK���*���4�qMu���>��X�a��,�|X���gHC�q�V(W���cu���|aHSs�U���U�T� �a9�$�t:f�c�� ��'���&/��� �^X���>
����v���s�\B�9�3�L^��YEm0T@��Q{��EC[&O5�F��ɽ��O�{��8M�ю�a�C#��h�]�Z��6ԁ�XK�847����U�p�:-gw&}'֓��x��4��*ٴI��o��h�{�;��0iӶ�5%a�E��A���[
E<�0�W~Q��E��:kJf�T��ݞ;��RKϔDa-���������oo�y,�a-�����\+`�Q�
���l[%���?$?~B)��TBT��&~�Q�1�"��J��i��ygcY�}��PY;�p�` Q|��p:�ϗ��j2��}9�<'�g.�ݍ=Y}�N鰹�Y<;'K��b��-�FyəUc��Y�u"��ʵu�\��*T�6����0Yd�PO��0�1Hӧ�)34�$|����N �pH�$.3�� r��ݏ��L������  ](5�y����D��!TQy�E�6��B��vLS���(������tZ������	�����Oo˗����Ͱ�LI+���
ynNwH^};̀���3?������QD'��t8j�@
/^��ǉU��H�	?���T_@�e�
H�pM�Vꭢ��[o�I�

u��u@���Tp.�������)�@P�6 �I a�;۲�W��k�`�={*��V�p\��;��dѾ�Np�:q�Qwɹ%wU��A��{������µCm�@�L ��6:+�qD ^���;���~,�ǲ�{D9�A��Qp�7�������AIR�^��Xcss�_\>#�� ��ޅ�36�PR�����#�3��a瞒W��hE�ł�T�I}�=��s�ؐÊ��&�@B�鸻O� [�y���@��o�c�ɲbZV������w�������pz��q0K��yT�|of��>e����3<_ ���uv�kOM�(�SUT<K-�
���a�Pqw��`#����g��۵v�3k�-�i�� �=Ή��C�q
J-��AՋL[J#2ݠ"I�Z�h4���i���f �Q�|�@Wm�<&8���Ms��;���D�����h�.@kR$x�/�[�}��[>�ٸ�o�^�Gna+�����Ηvq�bmP�Ƌ�&�����&��Oam�9�8�s�
�g�'Pr49bw�U98�y�6a?��#iu��$2(MI���l~m�U�c}Q�k7<��t{}D*�j+l�ވ�$KR�H��{�͌v(L� �S�1]�Һ�ijL�/Rl;���P��ǔ���޺yMff�e�@<���N�Lɍ���~NTF�d�)1mND��Z�l���iԌQ.
���TX��^�ǨjB�W����\t�!/�40�:���<�%����VG�B�}(r֬P�����!Z�/r���h*�̈Rh�3C)"�I�
A��ʯ�ZCv!i�P�2�7�z0����ݵN�q,�:�ۊ�@|�ɓ-�����G�â�%�m�X�4��Ml�N������X}�x�L&:���_ �67�0�4(��2e[G�B�?!�������g���ׯ_g�Hx�xވ�8�z���M �``--. �cE�0����s+��EǬ�-JA|R�Խ \�������LOOqnB��wrL'�S����<=���N0|��uI�����d~vJ�.ͳ-p1�1�f�gG��{��v��ؓn +���陹��dn�4���s�
���Y ���" aQe�����93��Ȗ���<�ht�2r)*�0��f�?�K�n������ĵ6˘�,xuZAZE5: �*,�D��p�(���	�0	����{l4�ḢZ������V��1�9��8צ6[.������4pc���#�b���aWt`ꞪY���n�\#A~�t���c�Fe�\C�������fQY�4ޑ,8~}��U9��O��6罳��{���4Y�na�Au��pϺ\Xw������t�:�T� Q��ĺ����g��j��YL��hq"���T^����F[��x��FW��q
Ë�1~�m������ޛt^�|��}�Y�Cg�x��G���J�Y���@����;t�/_�"���Ͻ{��ѣǕu��Բ�V��/A��^�R�g�:��*5���֡v���hվ�����{�CY[=$5�3�k)��  �#gi������X�a����7w�	�d5ع!�K��R�����}r֡��i�w��u�w���W��5<��7��iw
�\�粵�K�sJ�--�^��ܽ�*��ۅ��Tg�d��9yhh�>`��� ��cQ~b�&�,RJD?��� /z�� F[#�M*/��-��`�&N���%�.���1�M���h�Մ�o�Kҽh CJ�G��4\�"+D��!]IuO��.�{�#"�dJ� P�îfiѤ�d�F{N�t,Ly���F��}�}�|��C
�C��f���Z}����%rz�\#s���)����x���a�$�u�{�V�q|c���@i/8^����	߹s�����[o�-o���i&�)�tp8��I8EH�#:rve�\`pH�?{�ʥ`Ȧ9V{�i�>/+�Y�]dgX���(�H����j��Ϲ����`�RVSP���ޡ;3Ւ������Ji=��LY#������e�)n���������g�.�тrmmO��>	c�C%�&�W���퀵N�`�vd7�wm}]�ք �
��cQAw�jg�0E���"C�sҡ4�W�˾FBX���3����pp������,�����PQ�۝�
�Ѝqg{Svv�i���m�gљ�(e�� 3?8w����2���J�À89�ňc�c��Tk31�ߍ"��T3���ō��袆�*c#S.u� �AJ4)�#Z �Qx��_[?�V��Rnz�#:l(t&8[E�l��=i���|��ӧT;0[Uu����ͨ��n7l��� �<�U12�x^l1��l�s����l�Ҽ�@�ռ���i@�mA����?����V��ۋlߋ��6�"���u�۶�\���}X����%��^�~xM�)I��P��G���bțo��~@OBF��&B�0����>��i���-��Ss�ClXvwM���s��u�M��١|}�iX�:�6;�a��T��5�H���JY�= n\[ې?}�L��_�8OQ�u���U�0U��8 �L\�ۻȥJ�p�w�#�n@�X�aH<�!�@�Gl��[���n�]�v�RX�ߗ?C�0,��~v� l>x�.���RCTо�E��V��6���϶���,ӯ�',�h�8������K+�Qh��F�}����6��^V���e����ӹg�a�Y_S-I�Q����_B�p=3;C�ᅹyi��j礴i@R�
K/� �9�iO���z]�fk�j�vx���E%��,�q*T���p�B��NB�_tn�<6�p��O?�F>��^ (��:��(��;3���1V@ᩈ���+O�шF���L��X�؛�T&�r;������;w��1����
|�.�=.S?�:;_}[����)~�G������L�����:��,"*�q��;�.-��o��Wr��5.��ϯ�'	g	�6���,���H�	>�X^'�Lww@ޤ1T��aEp�j�@;�
6U`J���b�u�-z��O.-=�%#��ˋrf%8�S�273E�}oДã0��Y�+Z��`0���
"�h#[��M��lh�A�b�4f��
��;#v���Y"��Un
����sP�a/�D,�/a�ЩӪ��#���@?�Vq^���+2*��0h��d*�	�0����� d�h��Q�(o��ܤ�0��ɈR	TzR�|��aeC��N�,6Â4ՙ���}| �ܴ02c�(�C:tЅN��a �ᗙ�6���y��Zx&s�{�y�,ب6#Ã0�VJ��ڦc~(�K���Ea�WuCUm�Y�ԣ�9�G��༡��6�6����{nU`�y�M��@�	��u\������bp������/��*�}�1���ȵ4�� ��a=/*�^�@�GdEj%���1 �� 8���b�޸yC�}�r{�e����l��pߕ����e��x����ǿ�)@,=��$#��2~kk����Ōtf�i��h �6�$��>�D(��q�RXc��WU�>)�&^s��B*�FA���/�����G���i�ӆb(�U����V�)� f�Tբ��Xi%����*���V��VCbT��;�$�Up{��"(a������,�-��̂�]�ȅz}s]n�Y%@D�Q������l}|ǔ<+pנt���v��S~^��"����Ϩ0 kj7Bu,m$�
l�7C�=�~����P?J��2-� ħ�av	��)/�q��0�C��H@3,�0�M�`4�kϥbj��q��+�'^y�G &t�
?S�1�yFxб��Po�V4 ~�6�'�����򁱸�>ے/o=���~&���y�S�2�?�h�
�{�X�! cw���������׉ �Q
_�|����: ���?��3ޗ�#�N��a?���������O���i=�����p�e�7��w�(���orn���	�vzz>�G����3���<8E�r��]���Oe�ٺ�&���o�o�@Y��� `�o�xk�H���̮ L#Z+��Þ�8Ca�I���k�~����!�Ɛ��T@!z8�v�]����2�G�@W��0?���=��;(*��4����jCJ���?�V��T.g�:P�]��4��s�ҍXो2�o�ν.����h�����=>p�P�����:4a��"I(M6d������=e����nN�B����2�:8<�Ϲ��0&
�llO���E��"[_,�js�6�q;T��sҫ�9�%#���;Q�5� ����ذ��sֱ��y̡L�-�tZ½����ӵp��`K���P+x��%�Lϩl�^�FY�ڂ#H$\/J�����r�_�y�%w�y(����F[Q �`U�ҏ(��6��0{1:g�+\���N��Gy}��zFc�?�6�U��xd:v�c��ۈʄVיG�w%���R�L�Z���Ұ{�׈߉1�
$F�想�H/N�*t�D]�2�8l�i|Γ��E�8%m|{*�_zc��y	/�9T���1 ��x0���v��`�,,.Kw�X�gt�������x��]�t�:�SZ ݰ�7�Z^j0E��=�ӟ��;�<��`�,|�e6�QX���RǛ�DM4"I6~�����5r�#(�57Q��uAʨ�b8�����ti;˂���`�P427;/����b�?�i]��Ɓ��꠶��0VaA��6�hg��R�y(b���z�'$ϲ�(�O�� �8Q�2VA��1���o0��\5k��;�Y�x���yFf�΄s]	��\x�ӌ�����Sy��^X�7��}HO�3;-���f��
�4~Xb�]���F���)�?��k�7p�SnSU�4/9�P�	��hn13>q���$�C���?����?�?���wwS���2�:�EZ.��|>������E�w9�8�:�X�Qd�I�ߑ�������I��GI�LD�g�W�J� �駟��� L?�*����v ��	.�F�T/�.���~��S��L�b�-++Ka�h���ERz�� ڸ��L���|�����������lo����G�����C�I�FF�����Y� �~PsL#��0��{�l�: v����;2=7�������9s���9w���H��=��^��D٠Ҋ��.�:�f�mi�� "��Q�g�oi2:F-���eq��U�	��oP{*C���Xc�T[ ��ea i�iz���Ʃ�R�{~����ي�*	DF~�{0Г��KfMRJ�Qs����^.-����8k�.�]8DI\U��@����74�=�3^�p欖#�cW�>���ʪ��g���J'=�q�VձP��G�m��`���_���˹����-�}/��|����1��F�$85�Ɏ�>֨;nu:3+�<�m��":)��G�ᚷx��� ����C#��tŻK�~�^�X>��+ˑԾo���=窞�y�
|ϋ�Y�GQG�_��ݎm�x+ߗ�]�`�m=2�Q�ԴQ9�J1e%]��x>����s5��/��U׃i\��xz�Z���0�����>�����d���[�!ߖfC�	"�b�Z���k~�[�0đ���?��NA��Қ���W�~�3|nȾ!{)�ťꆯ�m�a�����[lվ�s [o�ʍ�����/����,�Jp�s�&r�����������3܍�YS����Լ��;Ej�{C��GWR�Lc�[6�:B����:;Z��@4K��2>v*j�ȥ��x�`\�z9x�s��[��!O�n�7w�Z��ϟ�d.�_�1�T ����FX�T�c�d����!��S�tIM�`<(4ݧ<=O�F��AMu�ؽ+t=���et����� p�es�Qx�>���=9�^Z���v;$�n��d{0����w�xN��� p�##�e�=�Z;�ROhc��%��"����+����?~@�C��(	P)�g�ʭ=���N�Qڿ�6���Ћ�����6D<�q��������_�߷o��r�/���\��8���hw�>���_�E�<y*+�Β��嗷8I��{�w��� �W����G��{w����ǲ���f  [/��w��f��ڄ�LMiĒ=��L��1Q�+9����%�h_v�ߓ�����9�!�BJ6��gh���
�cn~If��H��81ô���Z G�j{bPE-� ӡ+� N�sʳʭ�e��ة/���Θ��&�|/�&�rb]Cp,Z�"�w�*��Q���)�������\�<Z�hXݮܝ"u�k�)����)d5NLP@Pa���6���ܝ�Ն5Cq�^!�T�vq�{�n ��|�m`GG����v�Dd��KPt��"b�ޔ������8�t�}���f^V³�~���-�jMv��h�)9i	�b�g�{3��ߠ��U�1j�K]�a����YḚ�?6D����=��Q`6/]RУ��E[�^ό�؉�S�>�yϨ��ەb�g�b0�R_1����4;�s�Ś�bc).̭�e�W�uh@8�愧��V����������-���� �K�j��h��/ϵ�������=eG�!�1>�g��Ȍ)Ţ��,�৒�<m#�t�. �8u�r�_��y����o�Ӈy��������s֓��� �8�'�G��vx<v�$ �M��`3�i����tNZ��`�gdfv��	vE;8�՘N�sD,�~W��1�G}=2<��^q�%���IU�d����Cn�9����~����^���<yTʃ{�XnH����tA�K �d����46��Kz���	���Y��%�i�F9F@-#��m�i�r*Dj
L�]&�~f���ҙ�잓���ʕ�7�x6,� �HSvO�e�ۓ��c��
�u4���D`�JH�s'���T�������fX�����ʥ�O	�\�!��퉜���H�v��zr[>��|�ك�M=d5$��=��
�/�y����b������U��ֺ�5o7�&���aa�s�u'!��� ��sÖ��f��)@mx�=�s}��Qp�X�5 J����H.]�D� �A k���N ��?%��:	�q��̛�r!m�I�$i���KMA;� �M9wS���a�sF�R5.)���S�? Ѐ�Yj��田N�� J��F����ߧ��R�������gʿ�F'*J�mVG�`u~�J��;j���MiUx�'�/l�˨ܐ�kN����b/�Wp��'�L�Z$R�
\x����c);9"�Ig�&���gO�%0#��Ѻh3���"�<Վm(�;1Z�3��v;�Z��$,��.s�%X�y�����MX�&\R6�u��y#b4���q/,�gde�<e��><:�B��к���
}ە��dU��E���y�E�7huϮ� �Sm���^m
Ҩ8�H���
[4�?�`�#�n*pk�v1m`|��-T����������N���ǀ�4[���j���d8n�&��{Q^�f׉~�kh��TC��]��c�9ɬ۝��S�ܰh&��]@��ɓ�������X��Β��P��t�??�jԏ)��0IA#�΋����:���7ժE� �gno�І s9s�\�|5`�
nP9h{���յm�f��M�xr�T�����vu]���=b�����@u���Yb*/�u���=ϴ�#<]B���nuO����n!�� �����p%�����ee�h�������޺)g�]�'xx�)_}�D�EC����9V��}(4(W�+��A8�&�x`г��賯sZU��*	U��_lnԆ��X�A�"�F�#�-�Μ=��"k�����K��t ���Y9��x,{� �X�TvM'�-4UU�R)���c�(��J]6���ZKQ���=����tY�O��P>|&�������g�du���<
�u��s�_��o�[o���Nz_� %~�#)�	�XH�h�hh�೴H=��
�@+\���>۲b��«/��~@��=a�9>aQd�@�@��5��e�5��z����U���Z���h1��m6�hhU{ ��|N�'��JS�9�(����]�>�z1�X��������#oPt��<��zQ��~�G�b�'�Qe�J[���A@�{E�"v=�[-Au\Uü�%T��0ha��*"��� ��;H%zt{�XC�,���vuZ�V	�oƜG-��8Z�]g�O�wDJ1�p��`{ 8!��k��2�iC4\H�gZ��� �(w6' A�$�v� ���0�d m�����r%,�P%�z�Z ��(Uwl�Fbsl0T[�z�NWH�rP���:R�� 3�^�,\�Q~(��1���6���"��Hj�iu:RO��fb{2)��t���b�#�7��i[��	����Ɲ �1�V����8WPR�g���w�~�����ꗿ�ٙY�$��?:>�[���i��.Ӌ׌[��=�}��}����2B|��}�w�U�����8�����8��1��Ӷ�#қZ����`�c~��Y@{�7���7��������l�!��T��7����i�i!������
?؝[���32;7O5"�����[�i�GjKa.H��0�(�Z{'>���n�Iq��h�z�7n����-�Z��-��t�t-����b�S��>}0ܶܽ�L�n��������V�� /�1?�ч��\�t����u�NfQXأ������xpN�Ft(}�j>}�ʹC
���VCK�, ]2�NϜ��g�,&����3�,����W���CQF��_�..ԹR6ʼ�Ni����H�����U����c�����_�Gݑ��E�9T;���~>`5���</��2d�o�x��~� �e@�}?.Z��6��8���>�>�@��0���A�1^]�TC���&0�Q�|N�y��eG�$���Њ��xj�l�-�G����awAp�P-�Z�U��tW��_w�Q;�Jg3�	���"��Qe��1x���yC� ��6����]��9:朮�Z4<����6,�?k4\��(W��6$���Q\��M�:���ZXj.�Z>ǯŀ�J*�A����>��i��>|G�V�!Q�ߝ|�$]�o3SM's��]��T�
>M�o�Ů�����]/ȴH�{����.4iZ�a�3Z��=m���Vj(gR��hd�� HI�ϘJ�s�9�;U�j��F�\[���-�c��w�p� 9#/���8��[eմ�P�_��=*9����9�5�,*�[��"׉��D���T8:�m<o �7�z��Zؕ�V���DQ5B�2s}с:A�a���6...��o��9���:�}m֢�}�3�-���{�}��ou����b������U�GY�8ӄ{���Gl�����\8�9��
��<�~r���W�]��5!ݭ�y�rA��Æ��@��)f��au�+�:o3��AC��u���þ[��/]�C(^�����X������~*P�55����=����n��-E0�뫩<~�&�� �sܥ!;���(�!�l��a�J<�EA�VE����!�`���@�2�(�h�h�JyF���j�2��
���0��N�BG��]t���` ����wI��\7�bF�K�B�.wy&*�,��N�3!�Q�{��O}-�����<|�}Ex�;��P���eA @����m$�T����Gy�d���ёI�$1?/�X<uIq�Fʌ	;u1F;o_J� HZ5�T �$Ҷ�w�G�iJ����s.U���$Z0��
G
�cȡ�Q"�\�ʂ�pȨ�~]�M�$�*w����~[u�����ܹs��S b����t�B;`���:i"�E�D"�ü��noٌ�o��>�R��9� �v[�,m]G)hIâ	JJ���YU'@������$����/z3�E��AI\�uSt @�A�e@A� u�R�Zh�R�.����/m,���d����*�Q��D*>0^�'���6���M��m���f�7K!���=���h��F���ɰ�FbQ]\K����nPxVh"�S+����>��M���4�L1�Y�̋�lA�tx}�y�C��ƹ���jέϣx\�;����8c�F"�����%���1�?uKj	*?��NUEk��R���͍\9����ޤvE�o#<���������YS �ƙ��L��ʝ�&�qwI���qrjZ#�)N��򗿢�)��Ws<�~$a<ŎQl��i���笠)N+#�7a�.��G�Ԩ��1/����ۑkW��;��L�~�]y��_���OY\�
C���k�n8�����]K���Q�r�`������F�ux׃�^8�K#U�Ka�ԊWGp_Mŭ�b�	���@)��S�����W��"Z 2d�Z�PtZm9s�2�ywp��9�
�ݸ$/�!�FY,��Y�1�|Q�v��A^�3P����U����D��
�Z$�����W��|4P�M�x���y��"�Z���%f��:UZ�F��.�Z���f�@�Fݕ��"A��NA����P�ɿ�������'�a@�2�p.�WUk@�#�/��N�*���C�����}G�'��Ϥ�cP��E�/�םA\����2ݗ0������w��#I=3��������NөȰ�<0o9/�t�.4 �ǻ�M��%I�}������4m�0-��f �:��*���3�$�d���,W�\�>֞��ϴ?�Y]{��J��]fi�~2��s�@'uj��o��Y ��

��
}-��9�
x�jN'8��J�M+��>��PE���j�K����Ms���|դ�tv,��V�e����+ kVψJ"Yj�t���ŃsU�ĚG�4� ����Gv8y�"8@'|f~SqO��;�_2˖��IP#��6�J�(�}ri����Y$�;|Q�H�Z;7�� R@`p&�j�#�9f��h.:��q0�|�������'m�v"���cz|?�b@g_�o���;3U��?'���	�	�zf�01�U�g�2�	��йt@���ҥ����o�����ȃ���R�U)�aU�-KQ��ߡ�V��;$ �M���?�� ��v��2h���a�dL��q��/��:V��~�-Z�����a�H��6?l���?ؓ'O>�sgWdiqQ�V".����+��w���2�v.�����t�o��/$��ܬ��V��ؼ�Ӻc��(�)�.ӎ=�S(���e�uB��dd�$|P$Q䋑K�:����p���#�Ϟ�����#Y]��B��I�J��Je�UD�S�Z.Q�&SP������"�I�P�pI<�
qel��$S}a��ld��u���n.�d��120��4�:3���X�C����k���"U�"��(��*��s���@��ԧ��4��r�+��ؠ�����7w���I"��e�_\��n_�{'40(>H,5���G���Dl_���ۤ�ø��u��$ 4��˜[��hqG-)������Rj��Ws���+�!�N�G#�_� ׷�H,=������>��Yt0���6�>��]/�!�B���;���={���T�=���.;"aD�kϭ�1~�LwXu��W����^��8���(�ށ�H�y4;��i�8u�$��<v�weY� ��UB�Q����M3M:��#�UĮTǁEp�
��|�f#�4R����;T��|��[DEU���:;�9�+��.�"��ݶ�t�L�S���"��½x���<u�[Rg�ԡ�Z%��[�3�Uf �)�p�7��&���b1e��.%�ʄ���KiS�"���|&�C�R�}=l�!�[MS@���Ń��լ�����6.+g&�W�[��i����M�_�viܡ~ѱ��eg9�>�ң�l���ؑ6)M�ocbz� :w���sT��W��o��3G��J'�uM/�sgϯ���v��B��W�����w���Ę���S��I�����
��}�Qe1K対�6z��Ĵ��<�A�E�<a��Zl���ln����
3uW�s<�,.,S?�)����)��T�9f��p(�F]HiAU�H+۫1�l��^��TF5���1�2�A���0���j�5�sT�XDJ�3(GV�������k��]lv�r��}9:>
^A��n������m�7wWi�v�w��wn��K��Ml�T�EhX䪎i!��b����Xj�=={]|XU.V���rps'�KjB�e��-�(Uj�&�JӚdב�^a5b�(t����]���.ԩE9��������m���������ϑ�	�����i��������U&Je:�C>rj/z�ֶ׽�������wYO-:X����jݒ�gR��F2���T�IF�8�J���MZE���,��q_�_Xa��{�}��aή�6j�SO�>��w������0fW���pM��4@
*��Fw�|X0�ߵ��̅�(��ޱΛ������+Ы�/m�w�H=�T'R� *(j���W���B=�s8	:-�&Y4�S/*�rI�Ӑ�B�6�? ��ܑf�t5� �ɣ��bb���[l���8�$�ך�euS�3DsE�1��*�&����:(Rу%��k\��N��7� ܳ��jX�_�zUnܸ!7޸Am���uG���+�R62鵗���X|���@��ǋ�ˋ��9㯳�>�<~^R���;���9����'�L�������?��7ߔw~�.�I��޺��lnnсIS��j&�ii��Ԋ���@)�o���u��,��C�6p�Y��nG�^������l��W&���
)G�}�8)�5RE΀x���ޟ}$��N��Pe�D���<(t�1�1�lzѥ%2Oec(uh+�sz���g�O�".�X�{�Se�yׁ/�k�%O�9�w���q|��O*�('"����w}SyU��,-�ȅK�Io@���̀�{a��b
�n�];f禩z��u����)T1�z�,����n.����9uvؑ�꒔�ǋ�
�ʹ�P_jhZ�Rj���j<!��{�|����&58��+͗��'����5u8l�W�~����j�̏���j�I{z�n���C�ښ��ur*��1n?$��l�QD�q�6�⹬���m�f�M�G�=E�F33�sFó7�GS�v��A%��7ޔ_��W������|�,/-��~�'����ޔ��Y��?4�3�m�����	J� ��Ϊ����PH�/'\?���y$�8�
r�U�$f��{�(�y�u�j�PF�;�s��ו1Mj�8��sЗ�����]���>�I�K�Fq�`���ުs95sĢZ�^���'�k|���T�"��Tw,ꔡg�2.:�žPZ���l(���I�L�Q�����H�6P:BEY�����_�����˛o�E�{��OՅ�_I�zRE��������YG�ynRD�lRA���* �4��Cټ�گE��S�����^x,�W���:<ܗ�T�o.�{p��ө��AP��5I�*����yp�|q|��9hMZ�ŋ������2�(i���?�H���������f ���� qG;��AΚU�4n1��xr���K��#Q����N�>�t_�dt\�F��YQ���Q�=HL�7�j��NDVzyI፣����w&��&�;���\z_ɕ��wޖ�Wo���(w��R�?X�ߡll�z<��޼&W������ Lr��EL�h*B�f�����b��*��!x�����?P=������Ԣ�g��55L\�WnmRjռ���$�-HQ�huIZk�Q���\Q�zIö����ڞܽ�J����ʽ�;�;9�"����R+P+���בRE%�Tiӏ{�ī���w1v1�%?��aD�O�h���S��k��x}?c�p�I�5y�տu��oL�#"Z�[����8.�W�&�^�z]�������?Seev���_���ٕ�0�ޑ�3�ne�����IXȦg�8���~�]���Ao5�=���96T���v� �Ŏ�����!u֏Z��Ғ�Dx����x�*1��@�C-0+N�
H��<�9�5�cZ���!uA�-��en���b��� ��˚Z%�j�j��J��j��j�6� w�8 [��E��c�-?O�v�]��Y�B��t��^�G�b1�Ι\�̣ۺ_�Y��=�?�+����zu���ka�5*�qs�� ������}���� {����'��V�����yJ��;��6^�=���l��Ҏ��O3����ܖ���:B���i�H��7��� �)��7/o�����w�eq���� �?��Z�̾$b\n�[=�宭iA.��|���25�߹s��,�A�O�(�n޸���K����P�
>�Vδ��Ʀ�e�|���`�5�@����a��
�u�N�;�W������ei�^�'�e��E�c4X�Ю�X�_���{�X�C刔�����$ ˾� �dylKr���Ӟ���]y�d;�[���'����.��Z4�����>hu[�?�bV��PCU!��M�&R�9eю����f���lX� �ϮFR����8�� /޳�{�`7� ����K-��^Kt'	^��
�v�ރ-�{o]�������H�Tb w��Z@�V�d�Ϫd�Tu��;�㉔�T�qj�2 �/�.��I���>~�b|�p��ߓU�/�룑�r�3�b�]\p�+�G����֎I.\�����z��2�C��lM��?f�Q�s�.�ܸqM�{��������}��<��tVE� R��=�.I ��< �iV�+߲m�_����O��(M��2@�B��U>���5nGc��i|���TRYE��g� ��&rV�k�UDKY�V,�q�S9��<�b��S�~\�*����[��B�T�^��Z�5w	.�u��e%\ά�9�5�>39���^I��i�R��w#��:�� �4#��=�4��<7�����7n�o~�����!��r��2�&�4!�e>�_oћ������z��!�m�)vr����Q�W��~�|��b�A�^��~+��{���bl��.���V�8��Б$���!9��gS�Ņ�`3ޠ"��'O�^n��ZYTA�8+��ll��=S---�;�[�"��q����o5��h])�gK��
X1i�{�.���΢������>3=�6W��b�nG��Y�a�HSe�_&�o�,�x���IUJ�{'x֪AF..
z�Cף�$T-���7�8VZ%���
c���M��ٕ7�!{���z�rr|(���L6���	�<x�Dn<8'�����go���@��Vہ�(��@@Y�F�������*Ћ�Xxm��q�V�;�wt�k�B�J�����-�͒�p��o
�ܤ��$6�r�%����%b�
{�/d�5;8<��߬ʭ��ɗ_��w[��mI�W���체�f$kM��`�~�L
Dy��-}q}��{{��6�Lb� u���8�w�c �����>_gK��؞�F/������>먌�,`��z��������oߐN�@�|������G a��yC~�޵k�T]����~#��O�֭[�c-iZѐ:�(h�Q���͚t�[U�G4��㠭rˊ��C�s@��E{��� z��ړ��5s��&"J�P*V���QѼ*L�Gڲj6��i�e�fz����@1�6��R#��ZN�E� ��{��X�FH���+����Y�P�}����\��E��PZDG��0�+�4�w�{�)�(C�b��nD者�xP@Ao#S����8f[A�o~�w����$���_����_\����U.����Yyl}~�{�tqp�g��>���B��:��~_۫���I���'VV����H]]���h���g�q�:���":����t���]9#����`3���^����%h�0�a7��m��c?�����s�^���'����p7����z��Ҩ�^���i�W1�g}�u(h���:E���+�Q=r�fn#Ίj ��F�r����A����1�� +��[G��4�$�2d�3g���26Z�7m�'�?T}�d�6��ቍ��a�B��<�.^���9����/�����ȝ�۲���ܹ�!?����^��W����l ���O�=�8���	SwS�Ąw�rؕ4L,�����x���-�>=���nT��>�f�~u�s���L�
��M�Q^Jb]���3n^���P�4���C�wo��;w��	�-��;r��k.�"�M��Ux![�.&7t&qa� ��5�n�Km��^�{/S5���y9�@���1nq��_,��4p=A/�����vO��z�&�N;3�J�Q��NRb#6�����!�����E�ݙ��.��������E��֗_ɿ��C�ÿ��m���y(e�AG.]�̈�7�˙��3K� *ֽ���Q�6���
1�ۭ�������B��߸�H_"e��9�"�9�_�w`�y�ړ�ԁD�Т��
�4�]R�����|/��*�FR��2k�*�Ｌu&���a�I1�U�4���^eE��1��*�$M}���F ��
���F�Ȧ�Mh<լ�r`�w���v���+,��a�|�?�կGj�;\Yz�O��6�w���|#�ӌ�]�t^����gND�9�!k���!`G9�hQǵP��xv8е�=�zꤘ07�����w��_�F��kԮ���wd*z`9��p�/�9u�/�6i����S1H������'�5�:��]�&���oY�����Q�����iK��cܧ&	:�ݻw9v!}����Q����خ��^�Z������בi���Z��̓�
�&U�������f�i��pb��*�`�L�41�<�+<F�ގ'� W�7�@q�u���M��
N��X����UӢ5��JU��]Xj|�F��E�^�U�%Z�PG$l�{z�t"5��sr�s�J��1(7Ic@��R ��/]���,,����ȳ�'��x�l7�m�xwO��â{AΟ_�����r�fq���VW�����J�[��|�7a�e���/�oꀯ$��
 qR*�!_�R��kS?��C�����TD�^o���p}G��ɮ���_˭�˓�lǇ*�V��dvaA2�ǣkP�gQ�A4��S���܋���}E/g���<^u�:m0� }�<u��ix������S��|4h|�yѽ{�y���8��{���%���:���A���˗�| ��f��ܿ�@>��+��/�=Րgk�a._��ʙ�l>��,//��$ZC�QdJ"K�iq�V��\FR��B�8"9�#��0e�df�,D���T�m`:���{C�r04G��QE�'�f�FHF��V*����b�6�&u;�ئ�\jW �7<�%Ԝ:��/�.kT���XK�Ŏ�o��������"Q%��7MqIL �ǲGpk0=
"�ʂ����lD���6�2����n�T[;�MQw7�?���}�s(�jn�W��|5�w��{�>^�Ɯ���W�󣟟��8nA�;�A9^Rɲ�%'Q�xb�L�N
V���s�v�ǲp�4ء�INbc3m����*����~XOK�i:���[����3=�,���I���+�?�����0��g|4x��sz����?��H�>^��+F5��Q^:�C�%�t�C�ϯv�ʪ�5���j��a�Y��>�0��<ppo�^yh�T������%#O8�pvb��[�����aE�1ִ[M�!����*���]Y9��s�ƛ���+WesmUv�7��k�4 �Ͼ�'�{M�|�J ��Ͻ&Ǽ�H�
ʠǛ���� ԋ��B9�y�8j��
i�3��E� � ݥ���'l�� ��ኧIx��iV�q�0ᶶw������>�;w7xؑ��C9:�d�L �+�@]h1�A� ���>5K1au�Ϊt��j�����&�O{sN#E���Fa� "��J�ͣ�����T٤th�N�1l٭^��n x�T5A�
������t�m����a\?����N ��2�(�h��{tt���%s�{A�!p��9�u��O,� �T]As�nݞ9���wl���=�=��T ��8�up����������PS!|�c>���P��G_q�?�-�0����GYѾF�`M����Q�&��^0�l��a`f\�B�ݔ�Ţx,�s���ٸ�,��!x���������W���+t��R�(��I�鈴�ŏc�[L����J��M;
��R1N��������r��M��K�ߏ>�H��8T�6�ӊ�ˮh�11��9�n�_~�%3oW�\�_��\�=~L�ę�i���opi�΁�K\��E-��:�0N�)�<ʖ�����M4ȉ�6M�w�9��t�ڄZ#�׆�{q�%
��	�)���*{P>��������m��)d�R�E��V�:���-���
����ݣR�����2)�O������Gf���5���� ӳ�r�RB�� O�{$G7��ccO?ޔ��V��Y^������NO���ч�(/Ύ��M�_ϯ41���X�W��k�D��`�@� x�N5x�In7U��Ћ�L�I�i�H)'H�@|tԕ��=��ؖ�O���*��}&��l������9�Ӽ�;3�nudhi�A �b��R[�v��>��;s?�m �!���.@�/�<u�O����=���I�I�I���ȑ�2�%T1��^ɬ dqq�-��n�(N��OL~�+��\``Ц�SR;� �� ���ϡ
�% �I��1D|�޹
��so���@a�#M�JC*K���QT7�RED]m�'H�"�"��f8��C]d!�a�۽j�y�YA��Gq�i�^||��k��|�z�֟���Ϗ���Yj��R�P0�s.͑O�kp9������c䧒�;}<�ʾ� ����_|I��'OS
o:��Fc���e��#��=ϟo۾-Z�]�J���η�"R�,4��ϑ�o��l�Y�/�mx!S��8� ��ۓ'��P�W@��G0 Q�����Mz�\%�P�Î"G��S�0�U��SKIȘ��	ous���.:���xv*�����~c����eü]��C4-{SV���wڰB)��iF��$�3\~�f}Փ籫Ʋ��W�>�y�*{��͊�4����{�r׈�7P���!#����V���[k��H={�*����=�,�Ν��W.ɛ��W�_�UTn�A���<x�*�|���[Y��ϒ�p�����9n^��ὔ�a��h?vH���� �^ ���@*e�()�  ��Iu��I��4'L҈"aa��o?nMˬ�n��G��>��㧛�����1y��΢��/`0������� ������-MIV3~����W-��Kn1H�H/�����
؋ְy���(����Lz��m���.�ݮV�,<�D3��s�(d��K	��;Z{^�a\N�E�b�(��f�|B�Ͼ��|��F;P����M\^+��b6`g���P��9�T��=#o�kF;� �R��N��正�V�bQ�v<��Q��������/w�b��#�A�OA������i��xc���'��+�p�YQq���7 �G���ǫ�d�_��>��M�����*�8��Ta��}��������7w�p��x��ϝc�)ڍϸ���	��L��ktn��)�Q�I�s����z��dc�FⰩ҈Fn�VW�y@D����O��O���B������e�44�)�%5CSS�U ���(�}�IdC�߻�1��o0����� �9���ҟR���-1�ϳ4�)��`3�)�e>��ʆ��R��MF����΍x6X4���v �S}.r�)f *KXZ���E]XSU��
q{��$5j ��E��Q��~'U�������4�CU!H��P8����bʉE|��)�EnJ�P;��F�҆G��	|a���{ L=���ųҙ����m9>�7�X��rtw5�=���c�p~F.\������q�]�:3h�d*�B��d���Br;��۵�A���K�nl�-�2L���^0�]���v�Pv��d}}O֞i$ww�@�Pp���"��g�Ͳ&i�- �;I���q�F/�jR�	j덗�c{5��Oc����<���8u�-����WYt_���|'|2�B�?��ʺ��HU�B����ɬ!�ؘSe��I(V��[�x����8R�ڹ�nv� 7���*5�k��SPІ����"�1
��I�G������K �W_�V�Y��k��x�l�w��i���Ť�Vf��T��h먝�q� ���F��Z(�ϗ��6;�4� x�=�<�xW*�~;��w�-�\�M�֪��������y>�U�H7�@r�׶�gv�=1�V��)FY'F���:��q&�>q��&g����T [=F���
8X�p��]�Elׯ_��1��=�o�(9�#8F˚�(666��|vf�g�?�n�߭ZÏF�ڐ��-��Ng��Mk���Lp��ř������ ���**�MR�[�-�n��_��Ω��{b���k)�v2{�*��Q�A���
֏�zGm�s��6���W�[��^��n*��.��L��������q�.%�Snd�`�Ems{'�֥ b/ȕKW�+7��=:ؓ��gD>��g����u�te6��3r��\��$�.����W�̙ *�;L�΄�#H3���Es�Py]��&R���D%4�Fn�;yB�;l��{$���r^OW7�����Q��p� ��s�!��hA�A�0�՞�0��o-���d{g�I���*����W�uY���6	h���_:E����xq�m�c9nH�}[
4�^�_�9�����#�3��^yM��hB����"̇�1<��d..���Yv�q�o��&㋞j��RSH�B��e�yA��shR�9��&��y���,�H	�=*L�V֦�Q�|�O����4y�N���ѣ�q�j�"�*'���wf�֖Q�}9(�S���#�1(u5o�Q���
zDT�y�A���v�\�g);0�PC�7C����%�[ xѮ�����8@l�<����J��$O�ƲgN���L��e{Y4��^e~��]���`+����I�Sߛz�c;�kDQY�uPP��W���kO�Ђ���v�-�m-��:�������B�Ȉ@f1ˎG��ߒc���q`��В�Q�fڢ�x�)^������r��I�*6��:Q��� �S��j+�H�(<�)�h��uTX�+�FC�FZ��/]�����V�Ee�(��5L*W�Ӛ}淓*��W,2���ɟ6y�y�,����tXb�_} �.;�?`�ww{O޿<��Lw�ҙ����o��˗dwg�����'��遬o������=�AG��B���ZDu��(ܷ�apd�Q*"������z4=��p~{����nn���a/�� W�N�p� ٲ�/�3TXP!�֜
7��k?���?
��cT[�>��(��&*�E�j���.�N����`�&���5&1��#Y/:�_b�����{Ǒdg�7��	� �]��ю�#���j��G���oWz�y�hL�tO�Mo@�e3_|�ƍ���*@�̜��"�����Ȉ������ F[�/d��]'<�賢s�3�E�yzδ�.W����� ��캈Y`��U>����5mL��a�*Eu,l�\J��*�f͂A�&��Z�E�@�����D[�[�q1K���⯯�o�Rƫ-QŐ���J����R ���Q�x�� !�i��7|?���na \��
B��H'�l��hπ�Y�$
��f�Z�����b/�k*>Q$,�������3�(t%:<���ׯ_�KB;^�tӓ9"�Ra��(B�K�FZ0�9i�8���Ғ?�[;����z���C�n�u��.���jB���>�ל�6_Y0��j����_���^�J7oݢ�w>aw��������!�ځˌ�u%�_V�߼Ya��9�~�.LŖ���1c��`�����$�톸����n�7P��E����l��v#ʆ���x	J	 }�r��iȼ�o1i�_��F�e&�V�DeK~�%���i�] �1�$Fj�*1�bղ~I ��X�]i:2�@겐F�[
��!#�}*`9M^����Q눃�vwv�j5 VTR97;Mc�NLJ~��������]vy8<B�\�¶Ă�E&���*G�#/���8� @W�W x�ˡ�� lG&�8&�s굦�����}q[����7�s+q��N'V�� 6�A
��V�7m��"]
3V�U�����~��^LBr�"�W^؝d�v�6�<��vX|-߯<;�v�ą�=��[�
��)�n,r�?��i��Xl".��ngw��.lJ�z�Brrb�A@)�!����+���cD�}dC�Zf�S���^�O��ڒc5v"�ff�iĮq�Ԯ���]�GN 7��H�N
Mx���uW6����*������`4�䢩�˳'jbAl��
��������SS�-���Y5xC��EK7S�<�����55u
�:?�+񁉃"���C?�P��ʝ����e���ێc��yq�2��X��"tu�}<�9���D��sZ@���bgorv�t�S��j���Rkw�E���Bl�έ�����%�%����,�M�;>;�.���8W*�����n�^��4<�.�Ơ� #���T7c�Y�<�{v� Ue$^8��$�k���e(߽�������<o�a�p�G)`��O��Ӊ�d����+V���;3B�e�ߒpg������4(%-���l�A�x��fE��DH�!�d���$o�AaڌDYK#���Fۂ�G��z���ݏ[a;n7�ё���@SS��Li�Sl���Q���vH�;[��;$�B��憃�\9��!J�����W4b��o�^�	����U,��9ֽ*B��\m>�{�ŭsY���`�X���8�gȍd��i�E�h7|���]�~��hE C�j��ߥ~'4Y�����"���֍U��{E���� �vc}��a\�a������,���  ,�<wn�������=`_����wXH�fJ��0�Z P�h�,H�����Ji�&l'J���Zx��E���ӂ)�t%�[-�i d*�D��A0���v�4���n0��F
���*E��z��	���e&�X�8�:<��`��U?f��1�$��T��ʹ�� ����o�"�rnb�C���)�ss�<'����Ç�����y�1f\�� ��ד����?�k���Tŷ|`@
c��%���Pֻ�E�}��ܲ-\��g �L6�MK�/�Z����Ν;���@�n�b�q�ޏb��K�J�Ǵt��~j����`X�w���ރ�B�^�]�K���5KI]�aP/�����PF����g���@b���2\�(��թ� �ā-��(7������,sA�>�)���;<;ُ���<�!��2T��\�>��ڍ��Y�8�UP06��6����:8<���1��A�P=�T���=�Jˍ���n~u^��PRc�J�{s��ח�;��$�)��H*���Df���R��Ʀ�M�3.�Y�IZ�5%vF�\	���1���8��m��{��]�4��P��U��TE��6����~����m��)ӡ���&L����ڠ�K���re�nB7�I\ZZ���9P�۵�C/^<���u��+���ag�qހ�:8<ds������hff�E�çw���X���`��\�2���@�&��˵�$��
p0�c��!�o0r�2\���XL�������ww����T75��88��'^����y-�`3���i`ϱЮ����ޝ%I|����1GW�O]�=��CR�\�Pr��Q��a���b�p`v777�s'��]�*��Wr����"��0�y�ͮ5��������RҤ�xWr���-����"�D2�Lf~%��%���_���{�H-�250(�
V�je�ɣP֦ 7��q�8N������=����2��Eә�xX` �rM��Nm�g(��Y�1 ��[��{�!@�e�R�S�(�Z�ʎu� �)`IU��o�pֽ$�W-V��r�:.XW\s�`B�1����a�A��V��X&.���F���~��A���!�)���k<� �c�ì= �@�@ L��/��n8�G6�6���j��l���垺jnj&�M�f������3�¾�uI.~o�#as�W����S���xҦ�2Q~	�e4�����~��i�p7f�}k���)�e߱�:�i��y�cɻ3_�Q���nq���5-툆Tx(�򆶷7ٵhlt�K�޾}�����.�ӕ��fkG�v�6���G�w�v8P�x%�ȝ?�N�L���ܖ�����������'
A�"�X�����J8W��aq��\`F���������/�upeK'䷶�8����6_�"d?R���,�H�e���hF|׆��)�S���x�~x��|�$��7�9�LM�\X�Or�>F�]n�|�2ΛX���JDAJ7'�Swag��pF��p%��+�ɓ'���3�c��%�ώ}.��چ$���&	^��ܗ�`��)�s��`��lh���9����aZ�PLf�m��d��֕��G���h�<Ŝ�ڽ|��]#�����rp��r,]�*�CE����n����{R�	��Ε�W�r��^�]�!�*�2��?A@>+���7"S��p���K�C��Z.嘳lUK4H^���d�]��r99�W�)�>[�O�k��xH6�r�(��As��9$ɽ��S$���՜�S?�sgr忱q�+�Ai���m�7���Mu���W�(��$�`����Pe$`	$hM�_��K�.�v�M�Ƒh�~����fU�PQl�ɛkZ�NY���__s�
Dk���b��/�;KP��4�n�:�Z�`�ּ��?���� �P�~P���A�a.h5�^@����_[7�-���ĭ!as���>�_��W��W?��Wop�ˋ�������1���=*����w����-�'@Qŕ�LY��D�>W%���=�w�>�lose���9ft8p�ƟsE5���`	�$��s�*%�>a�*��
PQ� �ׁ�3��ܰu��sO�i��
C�y��JA�n��? x%�v�����< ��U(-�S���坌��F+��b�+ ����@��2s�H 
�L�g�3����f� ��Y�)эNA<�W�(�^�\�u��I�MP�W�8���l���of�������4�����ϛ!�YP&�2�����=�?7G[�d�k��)ۚ*��US����U)�gb���U%24�G&�d`I�,Yc�z��}|���q��p����(bsf*�B�"Ʈᰊ����Jz��k^y�fϩ_vX��Q:�L�o\Cv��4.�AɊ�#$[-�i|Ò[\�bJ5ay�ޑ��;�e��P���l�,����a)@�Ϻ[�����t3���L��b�H�۷B"� �O�̝s��CE��a�ӛa��*�R����kH�F}�)k���q�&.#܊E���r~s-I��H� �[�KfyX�X�[0�6%��B\"x\c�.��g��v��Ӆ��˘t�ǁ�~[? X�^�����:�6&�e�]m(E,iؗ��l!X N��ز @���`��-�o�)4<x����i�E޴�s�jҢ�Mz�������A1c����З?��4�������������ol��5�f0$9w� =�A�́%O-XZ[[�H����B����WTC�#kG�m�I�ݥn�3ŕ8p�\JYV<3�4�]<[�A-݋�Ѕ��yIj�t���{yY��,^lT�Kx��]��wvX�h~M�
�Li�k3�NnH�s�` �?����=K�:9W���uL���>�ꞡ���_ h}�+�����7\P8�>|�<bf�>+e���
�{}m�^�Z���sVn��,�.��7��(����q� �hM���O�N���<�> �ڔ�5k╪���Z)d}Wy~"H����j�Sfy��+�k�(:-\��k�ฏ���I��5�69�c�Π֩���ӭ��/��B�����J��4>�>4.Ј}j� q�%�E�fkh3�����^�P ��Y������w�(�����7���8��|G�V�㡳"�|6
�]���>;J�����|�Z.��Ic#p��}�SƑ����j�2u,5u�^;��Ç���է%vw��/4�&��?*��+Fd��
G(��BSF���`N#,�=O�ۋ��׫_�Ρ�B�Y���]��楹�4,k����ks���0V�|�H�@�d��?fo���}G��
-��$����]Gk�������Q�?yJ/�[��._^dS8��S���}��w���c$X P��L�JpW�7k�g�
��H�$������7lA��Bc�2v����nz�*�S?[��xA��9��>V��mp�	Ôqh{�_�Y��1�?����?��玗V$R�F�fM�t ���ɕ9��z��넲��3�n��9/Q0�Qw�`�aef�k:���h���`(�xz-㬬0�%(3l
A��Pb!췚V�//�����cc�t��C;�����J@F$&��=�%����?�5����[�Ld<'<Y�6���1��͈\K��]�uX�(�L��7�+Wb-��*i���߯�ߊ���w�oJ��@-� �����kI1	W��%Jw��0I~sivC<���@8���b�
s�k��SƤ�|�B���*xv�"����~��큫�ű�ȋ�F�XA�~�W
��8>��1���K�c~E.fD}��ίT��s�k��.~.#��aQR��O/�y,���~W���0�4�ۓ[,0U�^�21�&�Nx~P�u�2�(:	w��W�
}#u�H���_w:]��EG�سdL����<���½��Y��^G�-�^5��T70�*Bp��T����\���z�ku;&<.{����:����������
���ҥKt��eNK����zh�.~b<��Ίi9eQ�Ϛ�1�+q��@p�,����a���%���\#�	�޷^r�orr�;��><8b6T6�W{��� nbb��6!��Riɶ3���g��y4�Y�-v��2'j5�g�Ԩ��}u��ɐ��౑�l�B�ɳ�F��ZA��+6�_�n��o��1E��=�$��ވVW��?ܵ�w���ɓ���K��C�)����گ��o��j;��6����Y�������
��62���fueS��t�L�z��)��(�Oؿ�ߥi�
����o��SY�@��
�DB��]��Tg,0*#T�S}�B�x�1�2�zm4���c�ʠ5	��*rAL�L��!GƉSxқ���a�eL���h��@��}K�������P�����(�{��&�TI�>�|���5I�N���N�̡����wd�����K��;J�KWM n��@�'W����A =I�:Ѓ�x�v�o?f���Oc��s�u�`��6�W+j�Ӊ�0XM�r�߮�9i��
��{:����9�}v���DF`��£Ge���:n�Ny��7���)�H���B;E��%��-6�U�l�WP�(\��)����d�ZX�!|.𹆛č7(������<~⿋�d��S=N��K���h����x�jr:a�ż����ᮀq��� � �433C�����7�}h���:��sa�!���M�h�Jy��v�Д?:!��,2���z��9��(��nZ����=&z�^��z�;N���ue�q�/�_1!st$Yo�DW���i�~Ο�;�Ԇ���'{�?�����ؚ�X>t�e���(�u��k�:�X ��M�����،�4�0���ݞ'���l �n���d%�&��q^wf��=O[��S��s�I(��q�M����.E+{�B@��H_��|M��X;�/v��lW��Q/q�X�1�JԢ V�}e\�2T�Ad��p;0`K�M
?z#Eۙ���~���1s//x���}"�B����"G3�����{�0w�>3������`��]x��5K��F~�yW���yfV�ך���C`�5��Zp�2��w��iǴ�gs���gҿ�yE�@נã�(*�G�r������T�]�����8��� ij:�ط�:������ʘ�ٽr�
��y����F�;`��s��Q�� ��իt�⼘P)�>a�͆��� �4Ҭ�j.L�irr�._�l�"-\\`�[�"5iZ2����0�����R���c>��I߄�fν�\��0��s��w_�|i��8n�������fB����e1��8�K4�\zV�LH��A.g���m1Ƕ~��w)s�8�q��~��>�5 ũϿq�FΑ��WK%���^�p���%+I�G���$�[��Ž1�)u�Y�K%�Z�`���&����O|'�����+�͠���4ɺ�(I��Y�\��} ��Ǥ�ֻ@���r/���O�#���1�Ki�1��O x��U�7$uT�SEډ�DI|O���3��.��$��	Cp)cZP ������,&c����P�~亜�����;��/S� �{���[�z[�q�4��,��7ej+ҽ �h��;��*d�CV-Toh�e������*�P˼���#����}΄捀.Ai���J��f�I���ztX� T�A�^e(�������(U�s����\���>ۣ#tn�ݲ߻|�2MMM���g7 �����c�����G���`B��p߸~���{���mq���?�]"]��/^pa�Y#�/^�H�o�����K��F���N?zt�~��_K]�~��nʨ�6�@Y���f(I׉D�s֠8q�`8�#ROb��׍�8ͺ*�W�s�)��m��K���@#e-�����9�`O-a�� ��x
��2Ә��;�Xa�O��v�]��Z7�B)Ӽ�F	GةkHX2���)
Q0��ua����}P�T|��Ԍ���9�M�����'�ҲgJZ���cv��vtoA�[�ȩH]�p�(���K9v>\-�M�k�=�v��ǘt"�M,���S�-��L�s�Bqg�v,��7O���j�a{��Ur&�<�
�`  �Ů�X���f��
]"NzO�@;��9�.e�	<�i��ds�(�%�����S�A��W�<T�-�|�|X:��i
f.qEŞ{jj�._��E/�V�`E��'U�@�)ʛ&�*���6��}���n	P��#��.��k>�+���8�R� �@C�*#��5P� �� �?���w�Qp�f�!��c'Y �hbr��}�*������C j��O:���� 8֬3�g��s�S�LE
�qw���e��~ZQ���}����)0ʿ���((��8�e�q%�%����#�An9���
y�r�O�K����E/�O���s���YI?Pk0vx&e���Jd�1�/�VFŚԪ���b_\&UB�h� wf�\Ʃ[��W�����Xb�$'Td֊����"���n�쾧$��`4�Lae�hv-ɐ�jJe�$�sj&q�+3A�+t�`�܆��F12<�����V�e2?�Tk�LƐ�����:ݴ�����I�#�+ǏK�K�;X'=�d-D�G/?���^�+b��
 w���3�E���!��g�ht��nc���~�V������q|�8T�9��)`�<v* s��rL\��rR��BSy�_�{H�UD7���p_��+�. ���x^ ������q*2���*K)ۡ�qc������+���`vzz�_ �W�\���w�_�ӞUʔ������%Ba��K�.�[@�Z�_��A��Z�$� ,��޽�}��}�5^J�Uן;?�~��߼a�v�(�}��ql��Ӧ���e����ү%��J��p������d�i��.�y��9{�ɾ'�J�I�}�b
fR�O��_�����J$�G�3P`$��D��HM��-�̊�i���g��R����m̡�>1�G��"���i%L�����7Fp�Y�"Vq�Ǆ"q�5�N�}f�
'�,]��T�{��� �{�< 9)Tk���c]o�=W����k��`���W~n:��?%2�ax�1�vY��uq������KQ�	�e!�$~a����{���N���^�B	ȳ\��+r��1!�;zw${tG7�I���'ky!^�����FN
�1�����1�{�%��C��6�;������ڴ�#4w��Ǜ�E����isL:I�G)#��H:'�y*�f`Qݫ�Ҭ
aM�<�ѱ3���Jc �`H8�=N��;Ȁ��wwv�;�ǔ8o$|��j�̜½���̌
X,qP��+W�歈�6�ڵk>�������?~���3�Y��f`�+��k���
��������������������l�3�D�\�@&�D>�F8�/�� F�����IZ/%7\G!�W��Ӵ�b���n��cb�;��a9�N�i�X�x�l��9�+�^9� �ǳ����=qJ��)�� X��2�X;��רǜ���N��-y���5QA�-Q`�+�Bz�F�M�5p8��dQHp���R��X�1��W'�$X'�)p�ѡ9�����9Y�&$4j��BRP�EŔ�L�YcT�����I�&qb�����s��чX4I�p�|UKM/f�>.�&~��u�� �a$�l�ɖD�5˚\�*�.�%�fs�wce{Y	*K�1ۺ�r>Iv�.��(E{Iw� �a����s�W�~�ʿ^#�ֺ�]��A�]�B!���󜩬<� ��4޺'}�'g�N���Ns���)�g�ƫ�e��^�`�]�cx���=���H��P�\��~�1���!cVp��Y�U?X�w��u,5;@�d�̈́I,�fHy��w��'|�"1�%~�]�v��op@)�Ǐ������M�L�5ff�1�� �_[ʹ��T�袄*Ϋ�T��
w���/�c�̺���� ����ֹ��`{�<��
�1�=G�[�Ֆ�����ko3����
���;!��oݾ���E�gL>�k��Y v�\��֛�.��!*�|���
�II���#5U+1�D��@)�����Ȉ��;��G��J
Eڌ$d�JS�ѱ1���`RfZY�ĥ<K� O�}�"+N��<�fBR'������sU<�k/cقdM��q�|����ūA�����nk�(q	�{b8i��l%�{vQ���3�q��9��P�2�z��<��F�,�LA��d:��o�c��m��G����"7֮ty�~d�.���L��� �\΍SMЩZ!�u�@�Tt���+ ���!N)[=�۷���_W2���cmgɠ���{\?� )ʆ�A9!�Uƫ��λI���Zy3쩙5
$QǲH����uGQ��g��bs��故?+���i�\�Y��[��xHNXP<:6*��$�_�H�#�p�%\ P_�|����������\�z�.��� U��0� /@-�^�zŌ.�9�x���*��0Cz5�_�鸪[C��!�kq��t������?�_�n��>l���쟠���ݬP�OL���BK�{���.M��8P��gLW|��9N��B$�RQ���R�PsuSK�&��" wfz��>N���J�^�r�
Y��RĔ��Dߐ?|pH���upp�~�X[͠Į�=�!GW��%}�С(� ����<nZ*��N�*��B�$E: /���C���4lr\���_�`�����/1(MF�C������jM�C��.��e�HeG��ݓ�S�ΑV�,ϑ(�W�s?�ì����0����`8�����K��/�X�r�Q���ZF�'\��plϤ�o��#���'鯧bI��y3��O[�-r�}��5�^Z/��ms�����%� D��Z�H����=)�=n�}�C�}�DG˿�\�p�|J���0JXA�
bd��.L��/_���� L�[��I�-���������+�����Z��0�ۼir]z"�yk��#���ZZ��W8���i�������Bv׀?/�Ǒ���W����(�� �!�}ll��_��د4��F/\��;�����A` m�����aQv��
�L��e? ��|���������ߏE�?M�~������8���:�n��$��jYU\�VT�Rf~s��s�ud��{q;qnm�>߁��J��ZH����u�.[�N�VK�k)��n�/< N����0�[���y%�`%��Tf���1�{������=�c����jd���Ix���8fߗ�i��u_�>f�
��4]ÑfL	��ڱ�lK�l���>Iyy�?G�kU��!���ʧ�����9�$pU�aMǴ��%�$(H	݄SJ���2� �-Gv�1���4m�
\pM��H�wY�$�ò�jV�.n!m����6r�����2��I�KZ@>C�s�iC��[1ؕ�q0���=�g�8FG+�᥀B `B����!�
}��9yOڊ��~��,�0 C�(�#���|��]B�����O�d�ltW�^�+W.3�CU�}�/�A��F����y:8<`����e;�'w�^�p~���q�1�бR\*���E���
t5�6|�3`�$�]�]#\c�A:.�R6��u�C44<(@�2DW�^f6
���J����4�����t���p_H-'E6hoσ�o�G�<��-ӽ~%���Y�|l���Oz���u�9�s������O?�������?���&��`P����Z##����0�� Tx�?$E B�]�o6�~]#�
ʕcM��n[���J���D &� R���U+�a�krb��Y�\��~oߗ�V�ZTV�����T��5�|q�Z��t���ݽ�-�~��ɶ+�Aη��.	��K�+4����Yb|�o_$��8a�+Ғ�s����(�U��rz7�ߕ�r��jpZ�_�ޏ>D��q��$�WB���	e��N����.��̎����߲�l�FG��U�b�5"�lsY}q�f�dlJn�속A�v��`F{j:A�;�|z����n��;������]������Ճ���C�T���R��f@��N(�R�Ѽ�^��O��G�?�yא���)}�����~ �3o���Gً�ן�lH�ք�۹�9���h��������fF!,�, � �:�Ag؈��_�y�s���.�r�
pV��0L`]�&+�X7uN�f��k
�t \0I;撹z?���窨Yι��\�	f�礍x�Bp���4՜?0`-e`�l�he��|�� )߬���To��}��?EׇbE'��$~�r����_�΂�O��J��1U|� A*s5б삋L _K>ST�522�l�����6@3�����ػ&��M�W�sE]�ƀ]�#����Y�o���`hK��$z���Ԭ/i�O�ɲ��dh SЧ�JM��O��e�W�?j�0���)�`\��Pf{��i�Q�B4u�!��'=��,aw+.���g���v������OB�F���?��@uo:V<w��v&H�v,.6��}:�߱��+~���PL�eG� ^#�P8�:�:`F��q�,������d�z��
�U�vf�DN���D�tO�9y�}1sXH��c��6B���fL�+��/VJ2��$�T��<
x�:�μb����M&�
iN]�
�ہ �]��)Ai��C�=��~�?���,�'�{Dx�{}�Lhm��E��En =O�� L�S����Ņ�J �].na�Н�����z�Y d_ �<~�A!2  �-~���Ħ	�D7_��Ŭ��u��Y�H�dg��݂QT{�,�F��@f�9�,�PH�%sd�wN�H����_Œ����p��9���F0�<HBPD���'6y��7�nnn0��P�&�Ӏ���Bm?�4���/�h����|?}���^��i�I��ҽK����փ�s�V�����:w�����c�"�'V��23wxXcŬ^���E��ٵ��_`�#�u(�=%~����g����$�r�T��#���Ŀ��85����I�J�>����=�x�#((K���Z�����<$��r�h�|>\j%�)����'�b �`���%�NH_&}�>c�z���͸`A�l�5s�I��
�dk�g�ߚQ��4{�|W�+\l�W;:��w�*Avn����G@$w�OtI4`@y�F�@(�^h����[���u�5�Q}���t�(��<���o�y��NӁ�r��_��7xȮOE�<v���LГ3-��9�1��K�����p�7��5�����<x���\����nd곦�^G��E���ҔY���\M{Z�*����_��~u3��Y��7�0�A�G���YL*d�m��K��PDL��NQ%�$Q���/[���I+{a���>~��\�j_W��_��)�(��[��r��m�a�)\  ��,�Ե�C�x�:H�FUb�I�I�cx�Ɔ��A���iװ��V9��\��	�j�m�z:rEM ��|}a�k��OC����a��W�6�f�싔c�],E�z���/%�-xAu9$��Tˮ,�0m���ǰ�i�h	ϛDP����-�3�����nѹ� Χ�Kɳl& /�{��97h�1����s�l#��쇞iM�@��-���Y��Ak�봺���{�k�@^P�`�����ʙI,�k������5j�+ �����q�2��o�������22a�Z�c�v�()G.�C�d�U�4C�e82��4zWuq�{�a���Uٛ�D2�"�p�/a����e����/�����<����������J������>o�9��v�ʾ�D����\~�t�$�~����r�JI<�t�S��0�S�NR.���Z�Z�`��e�f��;�9|��Ԝ�U�1�����Fo$J�K�Җ���q���'	~�]�~s��_�@�����? �?o��w�R ���i�
t��-6A��.���k���"�!�N�7�y��R�������M���4�*���6 బ������m�u�~���������{!����P��t=[��e�KRq)#<ʀuaᢸ2����G��J�>K�~r�mmI-p� ��>������.���Z���*������ ��qް�I���{Շ���즍�l"�Y�§N����;7��J����y] @,��������O�\��)69CY��5�ڬ�#\>���BM/�c�h_�q�õN ���Q�y��K��G���q����]���?�r?�A��4 8�ι�*�5��\8���O�MJZ1���ƾ�kO�<��_����:R�!KXߦ����*�	�a�N�H� N�$-,^�5:2*�8:�w��$򠷤���C
P iɖJѫ�@�_�,
��W�W���@5v��5��m�As6s����cM :�M}v�4�߃c��*�|zm����X_��#�5�TV��y`Ͼ�mǖ&�B��������CG�e�� fJ�BM����{6z;��	Q�>���Z����"~�b�c�9���� �2�0���F���K���`���G�B�T�-7���۵h��6�>k��	v߾���T�HT��j���E>�r�A�;Պ�8�*��w�����ԔYш{4�ET4|�հ���[�F|�b�q �ӵ��8�G�VTz��]����?� �~��_W�v,"�Q�4�BP�� q=���#f,�H?��W�kW�)���l�s��r����>�=�
"�����477Ͽcη�6�l1�֭��_����u�^��n�x���`}qi���&y>���w�G��_�kmE4��1�)�<~L��o��};V�ĭ�:5�A!�~��@ �rI�q4���-k1��������zY[z��g�6�[Q���NZj"�p/��Vη���HJĲe��8q5����V���ݡ����o~�[����ѣǜRogg���kl)����b���Z=�;dwxd��C�mom��+��g?��.X�����.������äo쀖��n���E� �c��g�j�����)�(�z��}�c%"��xp���O���p��o��ى<�\>��rʮ�@��j��5Pb����U \�ݤM��\��Vi�Ö�K\��&>ﱞ_�s�2���dn=��Ay)��kx�6�S�f�Y�!KC�ɆT�!Iܛ��v.
�l��F\��G=��� ��t�=�K�����-��`��>��N\��E��;�'�XL��P�A3���+�:8?itA����:��t��>�EG0����5U�i�����W	���u�m�Ɖ���V�o5�Kꖦy?�~�u��ގ�y?!
@X� �;���9/P�w��t�;w�n�hbr�����å`�n���>�,��]��] 
�V!��'F��*��1X�|n4j�[0�t�>��K��>}�}@���?��7���sT��_�DG�nm����&3�񍍹R1499B7n^�Zm�Mrp��An��|qqI�Y��ˌ�&�������8&V�)��W�����*��v}��/���A-�?�R����g<}��ܑͣ:��4'KrJ)0��o��e;[�5{޷������K��u�R��#.���ϟ���Z���o���K�[ۜ!��/\�"-Ƞ0>1� !W1�!GkGG���kU�߻���q�U'	$*�(FM�Ha�j�oXtH܈4�m��1�1�n��s΁T%��c��iйr{&�<@�	�J)���ڼWS0�z����Y?�"y.��y���H͞�����Gw>��r�֭�4=3a�|t�|��-���B�b�}�o޼��(�~����`�����au����/����.)�`8��m%R��8�ŕ3j�}g� ��Q	�;��M�4��I?%f��F�)�M�/$��t@�A	�Dfr?NǴ�ة[�p��d8���w?yx⎷�k�C�In����	Y|��5Y�a��2&�֐��/
���hM� ���µ��V��5�*���5�	u�nXE���,��Y�+��[�.Ƽ������j6�g��x�]c����
�k@�(>}򔖗�9XkwoWrxVʜ����[��8ir����$��M��
t�6�c�3ӄܾ �����O��_~A�|���3��U���ܦ�/_��"6���N56>D7-�5��m7!�p�����i~n�Y`���*VW���q~n>H	ຎܺ������������<[X\�c���LO1k}��67?~���@�1dj���������۬��W��cc����An�潵Dw>��^�+OF��h��Q�<xD���[���W����F��l�Bz���}�6�>3;��a;O�HJ��]>k\,� ��ᣋu�^�v��{
�0����(��i�ұ�$������B��A1J�R_`0�-�<	�lH(I5 ��ig�xx�4G��H�D�v̻���r�Y�`w|l�~��/�u��-�N�h}%i�KKf
.�A�ւ��(_~��=��?�/��C�~v���Q����$`n���M����n�?Qe�2�lS7U�g��R�=�(�ց��P��CŌ��E�!�����ǃ�J<:gu��q��&Pvs}OAS�����tE���^��<n�w���9��������9&")���D��:&�r����B�%��n��4��dTC��L�K�� �?)ӻQa��:��L��j�����@��Z�M+8�q ��<8Ⱦ�hX+  ��)kI��b��,����'���֧�{����h!���:F�.�M��4�[�`W���hE�6U��x��������/�r~�&�YL��⻣��W�\rQ�m�J��M-K��6�-�>��3:?w�n޺��@Vʁ����M��>~��~������|�b~��^�e�u�]\8o7�[l�X��?11i����Y~�L��ߧׯ_��\d' ���6�Eq�)1[���2�!1̿�R��.]�DϞ?���@���t�D-���6�g�5؏o��h�*��1���2)�ҚMa�pa��n�?������kz��9m��p����޾C��/~Aw��a�r(�CÒqAK��l�yc�jf�_����|ԥ��A�Y��5� �5y*W\!w~!j
�����L~�����\!��w#�3��g���e�*oSv�+xv��˾D�{L����!�ҽ���nĕ�$���N��[�SS�Ĕ$hN㶘����z�j���������{z���6�֩�8dvr�\��@��^
Θ| ��c�q�5&�A	�bx��*��5V�٣�E���e�dT2���	�=����kSu��,�RO�O�&�Ʌ�HOtNͰs:��Z\.}��׭���������:[�3w��	'����y��I��̎.i<
O�~�����x�t�H�]t����+
~�$��7J�@����u7�f��S$V ��9��85
���I�c���
�n�����G7��TAm��bPp�8Sd�<�_�cw����[���h��`4D�ҕ��G������Bf+�*i�ޚ}Z���~��o�޽������; ����#��8��w��2�Z5:8ءݝ}��{�#Cb��י����*G�cK�M��{�ľ|�L���==}��A���ml���İ���=>�v� n��9z�f��v���`����o���޵����cp�8��Q�<;TåA�&vw������+�?|�����c��B  �bFn��ʚ��s������i>���|���5{�{����$���fwq%.�Ⱥ:<<t�
�}`��h����:{@�������k�h>��({c���D������뿢�>��._���p ��,n9�q����fXnF�����ݘ�O��SC.U
_9)*�")�D��R`6Y��sr��}��.M)92��v��4�^m{���X ȯZ��.8�� D'd_�`ֶ��V��?�jneNq%�E\����RO
�Q���Aȹ_@i��Q���ۚ�K��rŰ<�K�p�Ќ�b �����~��>={����V���V��_��g�fg9u#
w0��� ��x5g`l� ��/n�#=S�ǥ��g�e����-~��x�+�fH�FxO�{=��I�6 ��E��#~�����:� ˑjYQ�jg��1>gŜ��(�䀅z\k��H�u�|��.�W��Wľ\]B�\��$�����t0Y����M�x����w�0s���b�/��1�NR|�.��R�6�~(0;��v"�nbڜtz`��N�I�R$���":����:�^*p�c�e��f
l��|��2&ڎ�&��_U3�9H��B�M�K�^ 5�N�i���t���j3Ue@���c�J+��<����V���\�D�o����~���׿������!���O L�`z���\���˴��a�9��@WW��slH�#0��g�\�Be�<vv�S|5RyA5��'��L��}��%MM�Y@�EO�<��s���q�
�`zq>D�W- ��pXs~r+<���Czh����R����-иG�G�ݕ�U�\X��J"����l�&�ɝ���b�ƺ��T.���y��{�}\;Κr��������h�����i��[q�(P�g�V���*�-�;A�5�G��_M���oZ^~��5P����_�����7�7lU�08�5�����]ͻ4y6UH�&�Wax�?-��'���v=�l ���p
x�ŏU��+�X�x����C�î@����P%�̀f}��F9r��2�m�%P��(�
q�433�J3�].K��\.@ž%�/�jGV漶��K{�(MY�2�Xx{E��(r�t����Rf�����m1k�jtlإ���S�ˈ#di ;�$M+��ij`�U(��J���A�ʖ�����o����_�X|״��(����Ol�:<<�۷np���4c>�����z�Ʊ R��q��Ǐ0�Zn�%.�	n�����s�v�J	�����5��Z)��=%�����mфbW�Y�ܸ��vRMO�Ҕ����9���{x�J��st�n8�e�����V����ڎ]۴�j'��v��!�e-w��5������vBƎo���$MO�Y��53`&<w��$��S^���5����b��y��4%�~�1�����V���!ъ+���>Ow����L�ZM8�[@x�”��Cf�kV#F�(F�dپ+�[�P��n��n��2J-��>�&�#�����\5�g���^w����h-����G��>� ��< &�2i�w~�Hz�F0H0�C�݄o,|������`\0�0�n�������&���2�D"�Օ5�i��W˯mv�w���>��s~g�߷��k�$U��G��qc�^Z����Kz��9�y�j��v���,�9@m�͊ �`�p��l��g�ܘ�*FD���O�^���ȯ�{F�(0s�$J��a�C�W�N:Ǻ�^롟�����cX+ǵ�Gf��O�le�����Mh����w߳%兝�(m���/җ_|A���7}��'49�&	[W8V������:W��N���hmf]�� W� :c�՞]7k����aM��%)�������eZ� �Xڼv���y�&��S�|�.�>}��/�y�a��is����7$Ob����E�ru��_�jA�֨��$�! ��/���������4mq�����_��.--p<B�5tw��+VA~��'���L:A���իW-�>g�s�c�q/�^��o���ʸ5
�>��&}�ŧV���㆝���������ѯ~�kz������X�*A{G��?���_���]�N7�X޸y����bi>��~� �/��u��e�q�*����e4$�"�T��r��<~D�_<g����-��鲗HF
%H��7%�ɀ�~wi(�fwvn��\_�۟_�s��426h�O�5+��W�EjH��Y�Sg�f�jF�Z[٤��W�'���~@���ç�t~7! V��0!��ӵ��I1�M?��ˤ�\O���,�b�tS�ܭ�PSV#t��Ov�P��j����3���s�l�%�n�+�hN�ؙ*P��*bvn����|����6|d�hp�,��YU C=�Q�gg-�����'X$to(:���O�uc�t��wM���>����*�87�1�"�A�\y�~�� x�B�����镌{.`��d]��&�>��n7���M���P�lr5"
W����8o�-����[0�(׻fA/~GP�����nn�fiss�n-�O,�D�&?ƹ�9vC��͍M�{�>��V�����42:��А�	���,�\v��s����$��b��Z@��X��1�ّ��T^+96��RTǳ��`���ۀ�~�T���{?��gKT�k�Z�0qE��[#�����'L�f�Ō��W�\�����KC�+�B0M�Y����'�z��!q��a��4���~*�`�[`�F�����:~�
/�433S���	�����#V�^��kA�(ݾ�	o��Z�0���~z��X�ž>2<�A��#孭uV�Q�:�+ԍ�-����[K�_�DRF`���_�-��?�3W��q�U��hb\J"��M�]j��@���Ϳ�������b��1��g��M�sMQR�cQ����g������ϭ��{<�rh���/��aߊ[�!� v���w�bR�v�ѩ՚���#�����}���{���kO�ly�j�~�˯�ߵrn���򦕳����Xf�p�qg2Ա�`�77v�����~������嗟���O���d�1�,I=�����#.�Yu%QK|R����9vb������t��<-^����c40d� ޤ��c����:W��FS�asi&�8�ש�ͤ�Z�e�l�6��!I�KF��B'	6;�yr����ۋe!Y��V���8�V
Q��I�2��d\,T��1]A_w,�*;I .���@d��3�xy��ݾdA�4M͌��g"�OR�o�K�"u� d�
m/�_��V�!Zy�i�]0�c��ݦ�NmIs'z6�vq�?\+ژ��j�����9:�Vz��KZ��M�4��	�ggg�G9;q,��s�ۛ$οĚ�8��� .�C�G�.��f��R�n0��4����P��,(�ѫ�.o���f3�W����/���62Ze���l������} ��� 6f�0 ���>��\�;,�'&�� 秌�lﰉ��|	U�����?���e#�g`���R�x��nr$=�����S�S���̑�?wQ˯��`x������2-��e�W�}�.��3�v��{�V̱Qd� �g_~F�n]����چKP�{��Ǚ\�3��{R���(�o��[�:`�����,7��]z�|Ղ����:+����ĭ��/�F�d)��s�1#��磬�..!��y��1t�\q��f�-=P(��x�-9;;�t����F�&�i�>��k$댁c���v��� .����-����K�)���n�v�V!ߢo��޾~� �5�7��\m��N��IR�JS�g[  ��IDAT��(���-�?�ҥvU �xU��s��7U*�p��nf����V�]�t�.�/r�9�=�yhЎ/<w�,@~B.�ZY�s�`�.<�͖<w�,PT�E�o����G�/��ꆽ�>�{Qvʜ�F��2%�F삱.k��RT",S&�����y�PϏ���0���̐�V`�0[	s~���l7'6>��i`8bW	�G�B�3y����4l���tc�r�)	T�p����,LTF��[B]6��/h�=eLl�ֹ�Q�g��&D�K�^+:�Q�>5��]�w.���$�MZU�xU�����]%��m��؞Y�ۮ҈��QBrsc��q��:~A�GS��K��9��i��AU�6�~����f�.Zx�D�X�\�����U�lG>�^0��
�W�3 v u�S6T<Rr����&��3��e�3Ջ��*p��$������2;�zt���ko޼q�B�\�I�A�^$R.iyQ��Q��}�x�Z�d�_u>����<�p7�<�(j0�������-��8-�S*`�T�B�)�
�!xe���\aw
�3�^��o��l2�pWn�I��)�۪�'�3?I�7ȳ[���rXrt�Qѷ�}��V�yh��k���-�)��}y�53�{����a����[7iii�A��!he�t_I�>���X��Ju@��-*�8#.8aʞ�U��[+�k�m���V���m���z��	 �MN����]�|�/ۿ��H�F������%v��_(�zOMOҤu ��(��;������<O_�[���lC� �m���쫿�}Aᇈ�<���8J�O����n����D�|}��r�}�^�988b��~zLO������MZy9�V�ёq�����J�������ꦽ���ӝ�=���R�O��I�s���~����V0��B��ٽA�H933m��
]�v��G��c�:�y���T��������ne�5����(g���ȴ�����O��mXLQ��y܆�F��t���X��'-��[n��eM�'#�S+�f��d@ï�9�LTi�ĳz��v,�6u�4fm_�Yn �e7�Z}�
�=~���	�d*\K޸�ș@-�����#W�X��:�n��3�Ʌ�Y?�:L[!��u���y`l:���v��t^��Cl~z����`)+�@�7�H��ɩQ�pq�����#T��@�q�v�<"��%a �z�]!�e�&�Y]���a+�8��'[|��"�?�&ѭX�|��?�Qϼ0�Y*� VҔ�ˉ�a�D�[��	�0�_��M�(�5n3�}�xm�����F�w"�`u�k��:Ǫ�{DQ��5���u����B._U�c�F�bX|C�rx�el�<���{��es��M���u2/Q?�������E�[�R��R�)c� F4������>޿w�=zľ�p�  0NӓeM��q!8��u�8�;��4n��Y�~@�Y�E��](�l͍�z��� ,�3++kv2��y�Ԁ/,�������T ����@.�˟�@�M�� b�OOOYy0d׊�޶}��"sTK�*@^0�d�\��P���$����Y�_ӛ7�r}�.]Z��7n� |aKd�8T����W�����/��&���4�sti�3�� ���m��
��B����	�n�ւ��WoЕ+7h~n���F��U�<mq�+�1�^W��R/[0
 Hȹ����O>���o�}x�e�E����022ie�!���[�eE�����e"���?~�d��{˂�������.r�"�K57+�<�=w�w�?~�E+�������Vkdoȗ!疕��^��_����W���^�z;��X�+L0����y���F�CKӤ�@���@��z�}8b6"���h���پDR������N�.j��4v�����ʆղ\@��J����s?�&q[Ӡi
"�)d`��%� =(���!�B����6~#9Yc<��~W0���ߗ�s7��l��-�'6Z8�i�ʀk�75������-~$H�_.#E	���0�$e�(2xx�����Tq�}C{�`i��K�{�T�����]���Tv��9�6������!}β�k��.�\�`e�q�/�b�8wfЍ$L��{|����m���߷���&n��XG軫i��
#�f�Vwee��Pwuu��'�g��U���'�Q���i�>O�3�m\�t��Ո��L��3=���.�i�b	�5䁩�7���9H���� �G$92��~,���"�9m��h�]�Ф:�m��瞦σ��!F3��#�3���ň�.V�Ϟ>e�e�9k��&�:�Uh�Y�s'�J^ޟ���5�m�s��4Li׫�h:wK����e�ݾ�ݓ�g6�����^���[?�tS�c����u��D>�̞�"m)���`���[���y�����֜W���%�:�$�4F ���<y�U��5�����6��҉+�t���:;w�}_Qe��a�41�y�o�h/--��n�m����4�%��V�H����2��+rL}�C�)���	vS��J�����^�57݋Q����.�1[�r���u��>b���Ӥ�A��*�Ѣ+��v��2c��g?���K��S�I�[�k�$�Kpwb��ri��G�&��B���s34??')��M�3�x޺u�+9�:���#%o�Ǐ�`�_��n`d,>��=�xp��ZEI|vu>J��;�ㅢA�E�x�&CA�~�--]�5��dP�I�rϩ,i#H�b�1(�sH8��}xe�6�O�Gs��bvM	~�-1m��8G�s�պݨ���t�"�5z�|�V��G�F��{S�5�ɂ�pbi���y��O���*�����H�u��8Oz� ����
�:>Ϝ+N��<��|��Ut� ��vJ����A�j�;�`9�	�5e��Y��&��\;B@��5��%}I5��GT8|E#�42�0��s�&������z����ۛv^%5*Y�0P��H$�/W������m<�`?-f�����)�������>۔�"�_1��J�y�C���j��p�η�6�z�
�i��f\ ;��1R�^���F�8f�%�9!5�y��*v�k7�=�;n�U��x�J��HInH�� �,<Ỉ�:�(	��?��6�RĪ�F������9}_��i�bV�%ײ�q���DO|�ledu\a�U�c&."�%�o���ܹ9΍����~��_����ͥf�~0C����%T�¬����R�y*��K�IQ�B�'��|Z�|�4E9�4�װOx�ϡ�+>�>�.�oJ���$�ǃb�a*������E�W�=�,��њM�*2�D
�G��]��Y1C�;�m�2�<ϐ��l��Hz�C�ْ=	iK����/C�߿�+\BT���2+�H�����@41y�����S��J�I�	��J5������/���-h��fw��L]�H�Z�Y�mI�a9W�R��|#=Tr�b_E6�Ú�Y)^�r㒭
L)|�^��c����Vᜟ_�|��[v<��g�Z�If���K�mlѫׯ�鳧���� c~�*_��+:?7�i��p�y��ܸ����?L�c��*KqXh�r�u$�ߒ��;?��U�8�??c�[g@��gN�[��1:6N%;�5�w���kEHtJA3��
�Ȕ��ϝ��p�ݸq�����"�,��� ����W�x̝��D�JDW�^���a;pDV˪c�@tp���e���jV)�j�b�8q�#�2)�W9��߬�BK��. C���W�jF,޵�J���X[c!�2r-�t�����~-���Yۜ�m�̜
=�U T8	�u,`,�h()����;��&��.�=�}?y��SJټ)D���i�k��owdj�f��`���v�HS֑$|�ώa��4�µ�[V�l�b\���� ����%���X{��/�Ұ�ן�at~�n �5�.44�ED�Q��(s��y���A�����,#�X" &4��i��l'�P������}�\�֠�,�t��"�1�$6N�]����c�L+T��?��c.�� (���1i����#�+�&   [Z4�M�Ծw�-o׮^��\�@ �l;;ۜ�!d��5$�Z��4|�y����^���2v��E��ȧ��
�]��ʮ����f���%Dзf:RT!�$[������ɬ|��>��l�>y���`��m��z�4��+�J
>�"&�7��()$�=Uc ��˯�o��*��]��j�+2H�?~a�2��Bf����`)��BA���}����Ϙ!� ���;<���D�Y��e7��ئ�Wo��e���
=~��~�����w�ҁ]?\ #Rvְ[H�����)P�?~�y���v�-(ܠ��9�#Ϝ��©Ǡ�nnl�>�X"ky��y�*#dW�v�K~�o4�YQ���r��G&-7Ζ#X�1���+�p��{y�D^Y�j�s3�ͳ����*�y�f���խ|��I��/��Ȑ����p�HBQ�V�q�B��[�2?;ٮ\�L��aZ�ܧ-���| �-�����3�/�H�V�>o�XljK�����'m��������D�K4R�f�� �R�޸�d܃*y3���n��iP����r~v�`�%ſ�2��M���ʑ*�>r@H
h�
d0`��1M\A������,s)�b���g>Յ�`�USi��oRS$�� `�Cj�4u~����ma��0������R}�Y�ĥ����7h��z�-X��,-��r3Xe�u�fK,�mp��!Q�
�JQ�����{P���%'8�kƤ�����}>� `�$5^�Y��Z��"ߎ3�~�v`Wϣ�V���`qYɂe�Bs�� mkk��u��K�W��A��!Z�C�n�=|_?#�g2��Ǚ���&ܜȳ��TA�� ���ڶ9�.	�����Iv���46%�.������d9�����m�����Y��G�Zx=Hw ,�z���^GM92�=~]*m��Վ��b:�bd�ч����q���1�
v�hR�_��@MI&.:	�R&�k>��GN�[������gZ�L*a^g0c��z����>o����G�ۺ�{��b
xՂ.�L��k"*�MM�ӝ;��;7���~��ǘ�)���z������S��)&��@��?ϟ��������EO�<�Z] 90���ٲPr.W�e����]�zU\���~��5��ܫV	��R�&�z$��(����yi~'&��ʕ��Ҁ`TqeR�,��:)�<��<h���ysk"��!X��K<W�%��|���&����Ϙ�L�L�ŋ�ta~�^�|�Vެ����#�����`�Qc��k.���Kc㣬�|������Vk[�f�sO\7�/�V���7�\�O��Yxpؠ}��-��'5���E�a�Y������@Įn4�Hb�$Z�1Rn��&<B7oܦ[׆h|d��'id`�J	��o咖��7K��MD��t����O�!�\J���0o�k0�˶nr��� ���<�{x���T	�:�Yw�S��$鐡*h�=�m���h\�ax��أ����;�n������{���%�JTg�0��ي���~l|��^;G��S�,�-���U�A>��-��]l��?���_�5ݻ��$�`RdC�?�g��t{MѦ��g-������{� �cogv�se�I�$�5_����A�>�1S`����S���cZ�V;����tc5�ٛ��ޗ�
����Q�W2	s�������6�<;;[�Ï{���3��?L\�&�-��@���W��~����϶��P�ϵ� �^��vz�7=F�C��e-,\�E��#H��_T� O"�u�(ێ5<�i�+-�i�b��9��������+�g�bG���Y̖�X�3R"gr1��;95I�_qa��/���&�]^~N�	��^�#����b��8$~�1S˼��uD55X#�wirr�A����S���"�M��F���z�k� d|����,�E�����e�ָ���Qx��ox�*����ȥ�x��x�*���߸q��.��G����U�?yF7o]g7F�rQ�bW@�j�i�*� ���������%�
k<־41��o���5c9v���r�1�j�=��_@����!{?��6�3)���5CCeZ\�g��{����� 𮮮ӶU��8CV��	Uc���ڪ�IO9����.,\�reKիJ�t�\a5V:P@�Jm����y{3U�7�tX;d�ۊ��S+��T���8
���I���Fƹ�f<���! �����N���y�s��,&DS&$E,��f�+��D%��@��f�
�ԅ�k����t���ԌP +�W������Ɠ�%��M�Oh<�E*���g��93P
x�:+�*.Z�Z|��a��o�U�҂5�I��6鰹c�7�D4\�N�����Or�&���b��E�������kھ&�R��"���at���]��`�^]��.5`��y�%�+>y;=1N����r0�x�3��P�7�a���m���$�0�W8na���c�ǃy�{ �,S��j�}��� }�C���nX�c��C����B
㌪Tpa���cD)m{ Xԏ�o�v�����'������-
�eA������� xay����BN���ލ�s�B	l��.����y{��q����=	�+�K%��8~$������~�!��ڮ�gRw���Gt?�i��E����<��,`����W��)N��%fx��/�f���LO��7��u��H1��W���Y/�@MKi�|onnp�XF��]�!U����{�c�4pe�ˉ�\9rê�>K�۲w�L-	�]���s4m�����v����������X�O�>� _�A%90��~r�3�`R�ei�7���/�C.i�2�����u�(��@`�U��B���
��y�N&p�DtJ�U�%{cc�^�����
[�FF���y\�ѣt��];曜���.-rJ8`ʴ�*cҀw�AN�lʦ��[��Q��o�2֌*���dWqY �Q\��w���t�������D\+�O(:�����А]�x��n�3CH�~�S�h�h�`��j�*8E+c�� N��I�_��N�i.���*y��G�����E˾�6\2�`H�4�J5�,ќ��B\�O��,�����׵X>)�B�;�)�p#d������	όD���{�79��J�Ff����@���G3��M�W�o�ӛ�J�Y�C���@����xq���̮n��[%X��2��a�=q�En��8�y5Ԕ��b{�sAv���\� �&i�?C���4ѝ`���$ָ���SOR��@9zt��"0��`�a�
h��p˿�d�Mq��a ��I�xqxƖ�%P(^��������y��nNk8 �s ���a`rc�-�������:�6k>�[3*8>o�2����r����΅�����ͤ;㴰��Gn���9W���<c��ƶ~��	w��{��u��������so������l�r�Y���$��(#�ՉƜ�㠾au2��?�e�J$ �qZHV21)!i�<f���c̀��[I=�Jad�`naa. �y��Gv�7ns�"�! 'V��r�,,(C](iT����,#(Dv��a�� ��DX<a�Ko�s2�!�>xL�}�}�׵���!��(���";}.�/0�BW��K�s�����>�+�ӟ�_�V4��+�;��k{��h� �\`p�r"	B�����_�AH��cg#� �4��=�,]��o��0����:�M�# �Y ��p/Ir�����R'݊iD��r����䨩�$4�.������~��#�s�>g�;y�4��T�����ߣ/��B��[�t>�����c&��Lf�t��2�]�}�А�Y:E/�h��0~�r���j���F���p�{�R�Wjhht%$�
�m��IPh�TE�<N(���fs������v
�C��ZfM������=����6k���j3pk���i�ά������C�;�Eb����|_��M+�M[�6!)�O�����.h�$�$��HX���z��=hy��ȹ���-6�=V������ݜXY��
Vy���:���
�W�
*��kf�M�0pf��`�� &������V�%7&�/ �$�	�ۋ\�y�*���ϼN &t�l����&$ �8��j�P���ۦv��L�8g��������� ��l�̂ԛ>~`���z���}?��A|���9/�l�Ru�YB�D�9��Թ#��A��%�l�E�3q���no��?��jΜ�̥1��~u�:�eh�hV��a��Ό
k�}ү�=���݃=x�6���1�mm���#��vnl��{���@�ɔ��1��erb����}������Sdm��R�.��¯a���A��=�����2G���^@=�	�8~�N�8Is�����Y�%��Z~�����h�?K�+k-�Dǝ%i�j��ٽ�l����:�-��L	��č��3hq��.©�l����]
�	�bV��'�f"�\\�'~��:��/�/�ݼy��� ����`�m<G�O���s���͐x��?a�|���p.���R#\�z��Ƞ�Y�^Ɏ]�/��k��)�x��,(��E$�g��0�blC�p��9f������X\v���'m��v�r��hX��b����-��>�m)3b�7/�q�`�,�l��;����[��A��I3&�`����o�a@���C6X��}��EZ>�L.���k&���g��!#�* ���������x�� *�f��� �0
��v�2�ـV�
=.V9�6�n0�8osYh'�A ���-�\������,Mj�bb�����,y�u��` ��Đ3�V��aR���������ք��a�[������K5��j:Ù�:�"�آ,<w�
������7�50nؠ�T\�R�X�k�ka|��:��1�(��C�Ɓmh� e��To�i8ؕ�@=LDS��ۙ�h�f�<��G�|l��ifv"X�{,��0�UbbR��ߓo�JƯ"�eZH]�������EZ��D���b��(��.�A����x�zգBr&��0?,`PW�4k����u�d�Ô-`�R�6@L�I�	N��I�$O���ް8�/� '٧�2��MV�u�v�k�C���3��l�2�QϨOc�g0�0�P�&���a<'E�3��r�_�,�;H�5�����o^�=;�݋���#ח�i;��.^�HW�^�ͳ��0c�{nv����#2l7o|�������,���6�7�"�a#0�G�ºZ��ąE��.H`@�>�G�r,|6G�Z6uT�~c<���$��:%G�A�f(kc�u^�:3� /ك~�������c������<`�Q�i����g���k�ӟ�L�����k��`�������H�/_�ӧ�p,X�:
M�����￣��8&�Hs�:̌h�j�s�S/^D|�#�j޾u�nܸ�I$:�I�u���~�z ��4@��s��=��i�� ���uꓖ=���N��W��%��>��|�?�c!����Y�`}B{͇~p��1z�����?r�D����uz��cz��v��
Nf)R?Y[�o��}xF*b�&���!¤�FTu�� ��K�W3�'u �r����� J��*�bM�V5*F<"-���6�`� ��:aM.L�m�1�	��Jy� �7��P�Z�
�����S�Ol���@*-�xy2�)5
5ni���x	��bm�ȡ(u�|�j.���N��>m/y����z�TFX2$�p����ļeξ����![���9ꂯ�̀ ���Ψ�� "!n` �!3!xX�?�!�G���^g��7j��~F�������(�7ǈ� �V�\�fz�� `��XV,c���x{�vۋ�aǫ�oh�ai;� n2�E}!�hР�4� ��挹E���h��Wb�L�eL�(��-�T��U�v4��}͌�s��*3jh�j��"��Do�р��% �%1��\��8�vM{�?��������g� ̍ɼ����8������~�n��s޻}�6ω�N
���J_~�ݺu���pT��T�,y�J�2�,�m��|��:N����{{��)(�,���R����i��QΦ�x�1=~�Ëݽ}����Z nt��II��d�w�0��nq��B��:�.�ו|笣!����:����I�F,G`P�v�?��Ĥ�%2��� ����($�= ��~��?������e����?��C{��2��� ��N}�r֊d7���n5;��{2�!��ѕ%�p�\ �gy�D(�[�o�g����;�=fv��gv����?�`�!,S�w���8���Y��MĢ���Zg'�s$Sh�k?��0�s#&G�׈0Y�{K~�|��i_9���'��ۭ��������t��]�<�Y���O��'V� C���_h;M������Mi�ߚ�F�I����A�d��U�>m����Q����z.��4��>��Q2�ԑ��!�l���H&�Qm���@��N�f����a���� ��%D��.'����_��;o�#��+���t:h�U����11������ѶP!��Ztb(F�iJk'�.:-�tk��+gx�`����:�~�57~� �b�w�`��z�HD��6���4U��	��4�0��'�T���x�lź�	�B����+#n��d��)��El�4��b�b"�I������?�x���_r<�H0�`Q-������!Ͳ7�v��ƴ���~U�p\��j����P؊-53ҁ�7~�6%H�����>�:�q��sm���<׾�n@�~���$#�g<��������t�mvv\��k��~f��c����e�������~�[�˼p�M:u�$/�X�nܼ��H�����Nx���3��lF��Gr��-�z�#.��-4.���=�LgN��{wߡ�Mɚ�����v�.��&K���2�A���q�1-h-)yw �@����
Տ�M��H���a����8�f�>"`_!`�����Y�WH.a�מ<cF�����ycd��"�s�2}���o?|��������$��E �u��0��Z�N�����p�Y��2��?ҍ�f ����W�0�EZ�~���c^�x�Mf?�̵|dI��I�v��45��{.M�@�4�#�.�T���s��9I3�{����?���ꃥu*����↨&ǎ#<ى`,.�u�qX��Yǻ��#g��3"Ơ�gg��t_ ��k`��X�0������A�-0��2��RPT)�5Ұ,.��K:GI�u
z3L-6*|���M3�-Ę��^'-���DVU�Ccx噚�V���& ��f
I�4��cgv.v<av^`R��?�o�&V��[���W��}L��<��W��@k�v=o0M&�����4C��,�* �*<�����m�J�mg!elR��h�8L���SB̅_ã���v���㺅em��r��U�D%�b6�f�����`�޺�@��V���9j�b?��+���������j�YD7j�=��w���k $O���m�t�j/���K����EdKÂ�{��9~�%L{�ﰴ c�L�ھV{K�e�j�g:l����ɓ��޽)��1���OMS(7�_�l�W&;� 3� t�(��.�7��a�;�H���~�g�F>�Y�<n�����A �v��q�>g�Ԥ�݃@���I�m�r�9@� ���&}���܏ b�A�X�`%��ncc�C���C��\&�K���:0���<����@�AґTe�W2qFg��Ң�9*k
�1V/]�H��8G2�	�����M �Lo_���i��$VI�, &^H�;�1�`W����g=4��̯�B��k"��w9�
'�Y��ݎ8�I���땸aɫ⚵'�t�΃0�68b@��g-��+oP6���c�D���Ae�+ )�GTgx���3#%aL��_ �A��Y�]10��d�����C�a�c��{�.3��V��[/�� "�[X>R9�`ۑ�EH�PGX�]y��~�E+�>�8b�#��r������fTIr�/%Be�[�q��sA,�'�a)���0f����w�}���o���w�&~y�(�!������|� idf|pt�.oY3x�3dO�5*��M���j�aY ��+ k��Բ*U`�\��JF�O��#���� 
H��i�!�H�<W��@Q�Jf��Dņ��� 	�&�/cR(���j�y������4�u`�nr���Pg�e�����ً�3��}_4`팭���39lA �k�b&Ȍ~UK2
ii�� �-�xoR����^����ZB��#�X9�f詘E��%d�#�:���� ���Һ��q�ژL��=m��CIll�,���P��u�j4�h�F�6�B�-���|��8P��R�W?r� �=g�Z[��9�3Fh���km`�/�9�f�~x:�E̍�c�y O�8�FН�w9���c헴��<��;��c���0x�+<,�j|s7��E��7�4$�m�hf�q�qP;�+9�|�>����F��7.|X^����a�b�8�k�Dh���������_�|���g��շizj�� e �H>�˃@��X��ghO�����_LZe�J�'���e�A���U<G��y�������7oܦ�kOhg{�V?�k�~`f���:?�fhzf�AM�%^�E�� Ѝ���A�âP�ɮ�2&�]��v0���D��I�L^�,���0�5G �f>Ӱk;�;��h4�d+g�i�d8h���Ky!a�$�p�s	���ޮF;�TfP��Í9C1��"C�ѓm��N}9�h�����o���E�@(�c�VX� f!�,���i�;�#�΀8�l�)��.�������i�~-I��4��<�~���h��ɉiN "I�l�U�S�#0�p�;�Z8;"�Ç[�>d�az�O��>�l��9 Y��S'X�\��R������EcP|��=y?���9�J�Sl��t�|H�.�̴��]��¶���\jDe���)0D�H��0�� �=�V:j�c:��J��  ��$�ť�*�A�q��WD���G�?�#��%�Oږ���Z�zqब3f:u�D��K���Lr2�x�����=�v�<����5͢���}��G�AuJ/��R��������rM5�����]H0�a���rwX� X�k����Hל�(6G�T�+W{�5��p��Pb]���n�l�$��i���vئ<�үq<,��A�}Q��U�D��� ��5 5Խ�~2v�<B����O���m߃�}�`W@�0������S������^�?62��:ZVpq�>Qo ��<OMNqD����LX��`"<�����9\�}.Ǳ~jzfKՌ�pn&%9�
�h�}�;1���qX�q�9��P^�_�����E"x*�݇����V5@^cп<�MO�<�ַ�~�>��c����SZ}�����/۱h;�4ϴ?���<F2��E;2�5_e��F��|A�fi�G ���p҈�������6�>�a I?]�@�;'=z�$���t��
--��Ԍ$9F�`໵5u�M�^�F_~�5���&YL)J4��a-I�:��Q��H	"�tƉ�� ^d��{�G�`Vv@I�z�ϱjEAj���(���F�B��p��L|�P?�I�� �� H��(��.�N�Ij��(���[�Ⱥ��Q(�ӽq8�L���I�3#�� ����pJ�vá�Ys�:��Z*/���j@[�pf��*?�zy���r��QW'N�ƍ� �h��#p����ӥ��P?w�A�޹K����у��l��K'ON@4��-,�3i�,����C�4�W�݃�"'���Ȗ�"c�N����T��툰��@�^*�*-�t�F8�
<�B+e�*u*�4���LZ0��?ӫ���RU!�����{�$�L��-��յ˜��H�R�6����&zg�g�'�Rn�f�5Wt��nAN=E�$ܼ>i{�;\*�<�h("'�����(�Gh���v��N��1ͺ�}�N$��e�Fɻ���� ��4��^�Z"�&aw9�yi����y8��7�ÀX���6�����w���&r�Nɕqk�X� ,�� d� HĀ%��`����q�������ȏq,��0�V�(?o�8_�^��9�;/���"�A�A�a�iF�y
��8�-�xn���u��d"�ݸ��|��x]��� �e�ܥ˗�{�	�� ���aڿ+�}D4������lǖ���p:��wy[���z��y���>��S��04P�>7�y 6��߸:��!�V�6��m�����kssYW��\���>/G��k}�z�4�_�'�,��0��w��|��ҭ�f�7�?�pND�#��_�s��`׬~�;hi�[��̘4G$��j�s����0���}��uv�"�U#�K��,�Ω{�%��՜b׺t���<�.�k>�ݺ�3�*{2ܢ���{�{�	�L�����,�I8��5�FB�m����ѣǴ�l�ׇ��^���C��:E�JN�5�L�;���x洿��m$Z`��6�'&��r���цo�;K��.ݾ}����Q_��_��K�<Y��1�iMNN�{�	b]1��'$�EA�l��L����c"�s�p�1���t,�ޕ��8���iX���B=.r
�c++��c���/EI?&*;�0�7<�Ɇ���N��;ʲ)�B�B0΄�����~o����������&mo�w���<�;�t����f��.\x��%��P�CM������$>���Y4��"������9��&i�Y+T�S�G(��I�?������pZK�E��@��i�ȵ���$�7
.�z��XR�Z�z�S�6����i_��P�}sS{h8���\ŝ5g"�_v{d���h���^�k�ɨ�T���g��u��ڒ�����I�9祂�mV1c��EٷE�{0,E��<$�'^�CފUz��H�m6��a|�e�#��@��G�[V#"e�cC�-b�M!�No#����;����CO%!��	���'��rV�Yo�$�;U��l0Xr��<�J�����m\[{B����	�tDx4j�9�������Y&���y̷��@�/�0�H=�ߵ���2�'K4a�7����J��{X���v^�2F``a��/\�@�CA��.m��כЛ�>Ҩ?�\�������3�1c��^��.���E?ǁ����s�h�ɵ�y�������i�ϕ�
�A;�m��Vo��|��˷��z+c�w����g�Mg��$-��pM`��]�+@���6�1S+aY�̙�t��EZ�X�����x�r�|��]�&]@?��E۰�s�Nڜ?ۡ�p�a�LCjk��k��P�B�ȶ����vv��Z�>w���T�*��I`����i5<��l�&��4=;AS�A�z/ؽgss�c�ֺ�Πsr��X�st	;�X���e຀A������tB���ݑ�G�eh+̰jx%�� -�Y�n�ڵi-� �������a� x�|SvT�x���0w ��Pc/p�t���$�@�
�$$��u�Tʂ�.--ҩ��C������fZ�nx8�gx�3,'8�-�h�_�>�97<�Ζ�Ap��3;�s�;K*�j���#� �3�s씇�";�Oon>����;����ޡ�OvB�W��z��e�u��};T��@�#U0�~�	:��Y�&:�zKt��i�kA�a��0NP�\�vW��E�lW�q�S+�t��-�������x�9�e�5��܀�H�C���'��i����T�����6?�$�U���OaP���0Qޤ1�Z&�'L(߄�g��~k����Z��}��Jm���ts�����,��ޘ�JBe���Dx�aAp
���`d�G��E�b�r��i]�h����uEjk�2Me̟�yj�D�쮗x�ȧ�qX3R�X���Z�U�9FR�fC�u��pX��l$Lh��S�n��s��q��^�, �T ��S3����l��K�
�Sp��s�Y���=���U� Ǳ�����u�_z�<���@-c	-�2���P8�ۄ�9��S�S�J�e�-�X|gsH2�b� <��-t��q�- &~���qa���c:MNa�2[(�Fv�J�ʜ��yvn;O����Z�}�,����v�Y��b��1���;��S��ȨH��M��~�n���~K�Wq����z�K�;�\�W�{�y���/���{�[��h��֩�nf����!ڒx�7������.�O�����,%,����Z/�J�d�6��0�x�`'�F��i�ݧ�.é'9� bҊ����� �k@϶8!A�8#� XP��{�u���x�H� ��a 5`��F$I��tJζ������+��1;;',�����~5��h���vB�����N������v���w���7�����/����ٳ��ի��O>�� ���;7?Mg�8E�s%����E��G�jhA����?�_a��
F�9�/���MYzW���}��2]�|!\�#�r�JX�f���Mt�xs9����bD]��`�����%�A��2z͒U��0L.\|�=|��'�[�+r����\�ʱ���~���"Ub��� :�/ >џ�c�Y\�1�If��l���G��}.���P��,�oE��9�)�l������w�����"�{u܂�h�["���I׉c��#�\�ea��x���B�1���]��ɏ#P���aqȗ�e��D�m�PF�� ����-9���{�R�Iߎ��)EM��j��ps�jaJ{���i�V2�����g��r��`(e3��EC��W�J'�O�.svW^��$}�2c)������8�5&����F�����T2��.W�K$3)d/�l�d\"�a��YY��-��gNѥKy�:}��"��Ir��K!��hHB�����_.��t{�w�1�;����/v�
�{@�m��q�$����az���:��S�~�F�jwv��E��������$O����v?�t�t����V6@�9@�q�bed�R���)���b�����Ǩɸ��{�NN��&X��g��9r��/gA-B���R�fk�
�
1nF�=��)�hbĆ12��>Q�p��+�(�6�cfڗ���� u4b7����D�;" Ϙ�`�`k�-e7>G?0)�a��O�Te�q�9�[��� %ib�,�H��ɓ+L8��x�kLW���G����=���u�����u���Zg�4�$�9����-mH���^�r�P&Z���9ۀ ������?���w/r��If�]�	\��y,�Oz��n���o�U¦�G����� �%%oő	3���q�[ �d�GgϞ��>���%�s�ޠ7Ν�H��&��X^�~e�ý�[����=���#s��qfz�C����;t��
���NmBf��x��P�c�u��&��f��Y�|�r�+Vx���48RE(��t�"}��ǎ��ǫ���E{��-�$V��_�S �f��u�-+&Y�=g6�=K�4�΍?gϜm?�u�t�Ku$�U�����Vw�0%p�)�Q6����%��(��r@c��f,���9���pT�Y������m��k#ߠ����l� S���3��l���S��cI��,CF�3��y���D���y����-����|�\�]�N���2��8+�2���'����v>˲&�}�zka�GU��eO�iO�F���X8���4���YN��1�i�v.�u{�؋��=	:�l���t��C�N��C ���e�3���&,0o�}��}�m�l�,/.I6`�B�a��O�}�-�����d�	�L^B�XL����p0���^�1�m��Z}k��@݋9�t�lo���a 9M�� �A/����N2�$�	@e���Kꧽ��n��Z�����$�P�d�O�� �C�k�Ʊ��G��ƁO{m��y٭>�L�.Bxa>hg03���g���h��l�}b��Lg;g흔�sS���neRf,yb�������2�}��)=[ .�C3S�<T��ph����w�^���%6H�E
�j�Uʁz���kc�d�'F� 3�`��ga��цk���X�X��>_�A��d"��EÔr�^K�M�ϐ~ ,4���$'z�}0�g�������T�_{�C�y
����O767�,,,�G�l�w����$�ѐT x��ˬn s��2���ʕ��I����%�!pdy&�����2��6t���;B�q�0��%�q������7N򼰾���`�tbzf: �#t��I.�;֨�>{��޾�G8@81�#�/9�v��x��X��� �|��i0�gi��| �ﱿ�� \gP��j�#��`��鼴�,��{.;}������^���V��}��� �a �u5�z&	���Y&��gf��I���x��1=z�ʡ�`�9�b}���'� ����u:3�p��)�����%�؉}��1�a4��	��<3��0C�!�В��StI� �vQ�v	�w��IRZG�I�9�	Z*s�";�ke�kM�
�IW�Y��ƥ�5;.�]C��~/�Y�X�y�\��dM�g������,���e89=��9bcz�X���GQ�]*	;��Zs|NMO'���5�#�%;�������*K��al�Zo��q��n��}����n]���B��J� &s��RG(��비&�;^�ܸ]!,oڊ�y��d033G�K��#G�y;ZU����L�P�~��b�9F&%l�}��t��������g%3W�Z��g^���D�y�A�����xM&Z�[.����1�f�߿Ƒ�N�����A��u��w�/�����@p��=~����av���e��σ�*��=��k�y�$H��?Kh��X_�^��<y��v���,m�9gR+o�5@�o��v+S�@�v��o9��ֲ��+��k|C�\���x�:��\���ݡ	xC���7\���q�YHaL��T�8�$�X��J6���}N��e�iw�Q��d7������~j�C��g�Km�ʟ���k1#�,t"�����NҲ�E���'=��5	� ~&� ��e�6�4/� �r`m��� 7`%��9���n���$;ZR+"��c�j�2��H��l^ F`-���yO7M�ʂ"y���Z���0�o^8ǑX�%t�~��a'68���og�#�DUY�� \�A��k�i^��w�@>��Q ��4�0�l6�q��U�I��_�s���(��5��hX;��ۅ1�QGХ&�=f�I%�q���k=ϑH�$�c
�EdU�/���s��"��8�s ���e�ҡ,Et�YN��n8�m�ˉ���!1I���R+e,cW���̘?��� '`ZW��Z���@������b�-�)�
K>R.	�б}8M2�,%���FG��Ǒ�Nl 3s���t�Qd>G�!{�9��G�8��1@;'�W��� �g�0 �������eJ�0�55��ե�W19t7���L����e�1���@�f���y��Z&��?�ƨ�88e�9�Lm�K���T��^����lsJ�9T�Q ��t�`��!9y�4]�p��z�-:�B���H�@a���d��v�%����=~��A����������=ݹ{'���j�j�8B��h36m/��w��me�Ysj|6V!'�?<ek���NE�3~��x{�D���F��ٳu�v�D2���G�)�4 ��_�@y ,l���m��! �5�| _ `K��@��O[��;�oLm�o��m���6�dX_�uƶ�ޖ/��D~�6Sk�Pr�5���v;�u� ��s�v=�T������ 4���������.]�?��a�������H�3�Ѡ�{�m@�����@|�At.D�,��b��7C ߁�A��j3�
���f�X����C����6��B�J;�31��%U�r�AX�o�\��P��N�Ԭ�%q��q-X[���t�^bז�Ā*ư۷��7g}% �鞆�J�Յ$#�T�!.-yUɠ��T�0���$BZ����T'���*'�W.��<�r�=�"+�X�j�^ar=�87�p���nru؏ו1��1�l���̫�b�g�)�� �R��~4j������sFLI=�����d��p�E���H��U;L2�|(���(C(�� FL�P#Eu���K��o>���O�$Kng�R��	9+���Z�i>�;��1�*�cF���E��cDVV��\�pХ��"�:�4ع��E����Ŵƻ�V�$���][�h����b�8��L��������a�XGZ���@��8{��YUl�FX$����F�j�~0d�̝`��؊�b�7�m󢣌��'��9�h�a�ڈ�w�GV�5_���!���x1�]�m�B~��q�j����5T��>j��b��E�Sr�;��Őp
xYo�a���������}�]�|�
o�`[D����f�p������@R�^]]��&d�Ȅd���W�/;l���Ųذ��pZ�ŉ����':ZTPe�u9~kgKY媎V9���р�I�=,����v���LV;9Bp��V�e���}��]�\��P���Ptª*��j�S��qes���̫��v� t�f���(�$��h1s-���+3��������L�À}{�;7�Y���I$��=�C�$��V�|��
���P�9,5����*�,/�:�[٬;Ž�$�D].@(�E��%Z��9s#�Ǵ?�����_qh8�?����^�۾�}�={������������V���@47
��>k��n3�m}��l3�;��$��,KR�.K�k$t�8���I׈�3ɘ�5�Dl!)%�jA���\4��B�h92�!��
Nhd}J�����hr���{T\��qE�-�ܜ���ʒ�TG[��TwZ�{Xv(�6&��-�J�O��+g���p��H��|�MH3�C�#��sW����~�d�/-Z��K��R��`N��5�W�%^�k�S��l�Ï�W�:��ßՅ�掆���*.`"�H��vJ���[��k�����u��\�r��/�뗯p�B&O��"���@����툱{����t'ԥփݑU���l�pcy� j��x���qp���m|���2��:@��̫����d��I҂�z�q���d����c��*��x�~ኩ$n-�"�D�_�i�;,�9�<��ҥ-���N��!���M���p�� �H+	�d8�^���⢫���0fDi�1�>��V�X���1(��j���ƶzt�A��s�<�d���i�7@��8\rI����1�fB�B�:��|�(G^���ʌ�ٳg��P`���'���s���w�u����V �9*��d	C��1(:�TDYy�9��Ǹ�,c��-�zI�� P�X����c�u��,R l2'#n_�E�S�['����X�_r���>@�w7>!�8�"�1�����Mq (��W�~l]��;jY��"�'/.� ���`�P~�E<�����3�9Sj}�E�>�6�)5�{��c�.�K��<:@~�����#������������{�/��Z�]��Hh�M;�x�����gΜ��o�g` ���a�4��;a�AW M/�,��#y��o���3j��8�k��n#16E!F�l�[�Ǻ?lY3s��_W�
۸������L���έy�2-���Jݒ���s�4r����][� M@�T��}d ���BC�k�M��ę]����h�p�sٳ}ç��흳��"��6.O&cK�a��{>ޔ�r��}~V�6�G`���Z_��"��NP�e1lG��S]���d$s����0X�@�+촮s��������߇�x���t<�����իt2���W�dh���:����7� �r_2��]�V��z������Z�[45�k=(�o�g�Z�ȏ��YO�H���	j���bb�
l�D�ez�5����Uvzԇ�hb�f&�i�?�451�EC'"�*�ǃJ ���Sz��F[Oi{�;��;�~7N����u5�liZ�W"��V�_X�M�qk�9!����,�}������<��)�����zaZ}�܃�X�5�YW������t��J��PV�LcH������?���������}�����d!�ce���<?_؍��'c�,��9sciw-%eLO	�[oSS34���c�x1E���7�99��.߳1�|M���f��9Df����j�_���.^�m��cu�� �[� �phh̝��}_�1���@a����H��� �*�nl�1��L�ތ�Ł~%����ٵ�����H�^��>5�^�K�h�b�l��j�qվ����X[��_��/lj�����s�,�k��,�l�)3��m�W����ݟ}� �������嘼��h�?�~U������_�D!�O�澇�#�6�,����yc0�	Ǧ���v/��+v<+�����w�4��h}��k�:���$��(�]�����
�Tg�-�e��Q�hg�>[��F#X�{�('0K��5�ի�����m�3n��h�.��Mn����]�(Rs-�	���gFU������1L˭�}E��ꠋD�pV�����]��� v���O���e@�sl~��'�態��PW6vs��e(�&�����
��������#����TD�i�G+���Xf����`kr~k�f젲�V��)��l�BwU�DV�E�uh^� ~���b\hjaL���'��©烅�H��V���ݙ`���y{k�S�|��)�h�	��b� ���Qo{���p~��]��*�&,D%����R����e����Z]�tJqM@�-1 sv7���q���K�"(�v�F{�go�Y�������d��?����k~�
�Ilafl�@����}DX�mfC	N��"N�dQ����{|���& Pm+֘�H�3|�h�LIl(I�
8Ϝ9�;�!�!�;w�r���38�mR�X܅�L�!�ªJ���l��]H_�����k���[j�w�a�J����nF���V���l2���؉@[�?#D��$3h[|��+��G��o�KƳ��\7�{��wͷ�Ǳ���i\��n.��Lgs�����l�j�V�qd��[p���3���#������p=x����q���=^�a("���{s\�X�!������O��"}�/"' r�y��%�`�EO�,�;HR��3�]��=^	��FܩEbWb-*4u�]�_[<v+���d��]eh�'�h�\_�#v{ۘ�](�1*����1�jr�eMG�=���'S=cL_��<�F.e_j����.��D�A�}ͷ�	\Vάx�� �5�7����\��LЇo ����.�i�����dR����?s��O��|J��c~Cv���b��@����ìV _i.��*˜�H�UҐw�| ��Zۯ�M��(�:ETq�*�%H,ľ�7k���}��$KQ\�>,`{���*}'LR[4Bpn�x�v0�E&�r�:���$��)U���U0cx�lh�N8/b�v8LF����Y;!!2x۹�����-��\@�M��D�1m�������60�8���6��,"�+��2��e>��Nn
��0iT�KO�&�F�ٶ)����_{~i3�܀O2vj�4�)�\,:Xh6hg1�q�5� +�>b���?y��l���9$gG��|e�%�	 ��d�^�B^�a�-�pL�d��h�iZ yN��`����}�ɧa���������7��_~���>z�lu��=d0�Ó������0�lo��8YD���W9�Lg����dK�� c����s��X\�G Jc?��[����T��M���bi�[�,�7�=!��ֹ� �^��jeE�2�7�f3��cNk�X� f��=��A�����]��^�$>7b���a��8L�l�u� \w��mb���cQ2#�$V���`؏.����������)��ϩ��퀶�x9w�<}�ч% mC��w'bL`�|��;�!Y��n�,VM���n�c�'�p*ag��Aἥ������"y�7׬$34ws�y�N�F�OJ�P��V���_)��Ȱ�V>%�c�l�Kr�t��R361g	�wjMGm���2�4j�����n�a��[�L�U~�7�_��A}�}�|+�o���0�a�XF��������s��O7���;�O���y����G����y���U���������0P~F�P>�	�G8�q�� /i��d7���E��:e朳�m?��0�e�f�Xo�q�臘H�N��<��VJ��Ø���po���a���^0�C'5�D"Sc��맨�&�g�l��'ip�����U��Dx��Y�ه��$�,XX0y"��J~�r��;1{���:��峅r�Xf�	�lo�y�I-�f�?`��W��^-a�bșmw3P�ڱ9���}'}�8��:��m�܉GiQ�(T7Y
u ,$׾�F�V����:~b����9��Q��G]:}�����1�h��X{��chb�[��S����}"x݇ձ��<ӕ-t *���c�,:�E�����V񱕣�L)��{��?�c�w#�_i�`/�Jƒ,<~&��k�=��k����=�췎7��kIڻq7 ���J%���v�r�#{m�6.��/G��;=i�1���_�~���>Pk}�2�������/8f�sK9�����@؎|W"�c�o^�<F��M�˒��m���9��V�oYH<�|��<��ڮ�lO�t:�7���O?�/&�`����gV�|nzk!C���Y��w�ҵ�ѭ[7y���C-�#\�����!
��-�8����}�������qXp��S����b�9��͌�4v�Yv��L����`�o
uN*���|���ʐp�ќ���>�.��q�q�����0Jsz���x���X��+z�Z�|"/���xcA��;�':�c��Â?T\f�h�R#��l��O�oП���06n҃�����U$�8}�]�|��������}�����!c}��C�(R}3A�!��	p��횸C�Y���:eS������]��mg�vG���Ѻ3'.��9�p7�|�����`]w�8�*�.��#�4�ar�3��l�a��S]A� ���/ޡ���������QP��-4*o��}�p�|8�H�8|^N�D�ǁ���WФ��hw#�{W<K������v8G�y��?|����� @���־��.0��:֌�I��oy?���0j����dlIX2/r��]k�mAıD���t�u��9(���.-�;W���ƀ �޽�t���t���w�>�y��x�����$�?�N�����@�ܹs���o�&.}�3�C{��@ǂ<��E-9&��cGii�;��jv���!{c#�rܣ����Qԭ�-�o�aa�)�3¿b����{�����dX�6��lA	��5'�9�E~�׀Sl8�Ӏ�p���,?�M����[�h7 #��lv%]��	�� /������ٰX���5�ɮy�T�@Z�x�c�v�������-���1'5 ^nGv����0�jS�97������ShH*c�0w��1���γ�x��%�F�:���!��X�dw��a|"��;��I)`Db[�>Í6���,c���m`�뽭����	1�&�l��+��R��*�Hb�*`5cSds
��� ���/�y['��G^�3���'M���.���m\���jl1����H������W�qU�s�o�.�o��KhQ��d}V޼\i���,��wڼj�MV��v�!�*�¸y8�`���Tj�o����/������;�wÚ��B�㙙i��c�c���X)�� ��()�O�����9������g���4d�g�B��VW
��e�sp3�j�v���x(�M���<Cyq��|:��p��Ȍ�����0L>�� 6w�T���'� h;%��̇"N�����ߡ���7x���9c�^��� B��d��a�n���p��lb؞��2 Z.-q톃���a2Cp��&�N�^�� Mb1E۝����N�;����6��&����e���"8(�b�խ��%��Q�ڛ�tŚͺ2�U�O"u���"��K�	y���pu���d�h�4��튜�S�" >��/�����\��#_}�5�'�����ɓ����3���L�s����O�\��.�Ɏ\�Abk�~�o�]c�x}}��R3�_�% g �4�� a�`�p���g���|'�xgϼA�|�1;�,j֤���;���x����EQ�2�Ѕ�����''$Õ�m�ɚf�Pg3���D�Ͽ��B=���d�p �^1�!q�+��lv�/ZGyx;��S0S��*��7dm�{�O�����$��PY�vH :�s�AV���L��� �ـ�x "5����� �,5���"V�m�m�fl.��,�/ �I p��&� f�E��`�pX���M��n�?����7o��@w�=' �2d�_�R���cyY鲲+
Ͳ�[ۖ
_'6|�[���T�(��I0&?��#66z1���%���
�;�Z����~��g��~܌�b�a�� ��Α'7�����,�x����7�˽���2�NHf$��y'�t�%���|[������6�k��k1�1L��Hڑ7R�\25ۺN�r�T˰�Q%l�(Ig��kyՉ�d�_r����p�׺y:��u�$�u�y-��6��k7����T���u�D96� n�z�a��J�������R�T��i-�����u�#b����1rty��}�=��O1��W'N� �B�]|��}^k�2�a�����͈o;��#�$uiy��sϒ׺?��4C(ޡ^����e��kZ<��|�����ɧ�"^��[S��`���)�4`�	C ��`TH'�c�4"Ͳ�~ ���.�ʙ�X�Y��#(5�mv79g�N�;���-� ��/���:.���t���N�G��F���M�� r�Na�E��~I�Pg�8E�<�!��G7��n�
d)�;���$?�ڮK�z['N�[��Ξ�q�͸�}�i�8H��n�5i�k��	�e��ҋ�6�%r��ʾ���[�d�ə�YN+��� ���?�S���ɓap-�L ����<ē�N2�
���l����y�v�]�E</���#��nL�� ����� � c ���ǿ�a�0�	���ެO��^��p:��RҘ���D�E���_q^�ҏ���g\04�{��Q�]k>������I��L]*ko4�]�kΡ�[0���D��3�l��"�ŗm3�9s�c��,;Ec����+�t..�!]�r�6��_ۜ� ftz�@�1`c�d{ƣ�q� ��eX��!ki_/�����8� (��%C�E_�y��v%%�gjB�K��ɲ>�) c֕5Ħ����]9�c�i{k����s��{�mW�޷�E��wu����ϸ�h�{s��Q����<������i2 x��z�������.$Tfx滳�\H-y��Ǵ��R��@DI^�.��8��X*"!��<����8�	����R�F��:k5����ؕ-0���<%C9�^���G$a�(��lb�k�z6�%�#Zq4*��6��ު3���I�Y�QO��t��R6��<��:���:=&r>x�7�d^�&&i>�j���e^���jo���x� ���Ts���Pvx�ҫQG���y���8�4�=��<�F/�Y���l�b��.�A�Fj|!��G�%�?��H� ��i;��p���wh����^�u�X�P�p.�r�C��:>ѐ����:� ��Vx�zF{�[1��@@b@����b�ڛ貦	*ʢ�޽�S�415G�������. l�� �2�����؎��h3L� _�	Ifa�T2n�C�\�d�f��~�vR@�iu��6Ih�Ĵ�zY�����d�d�����˾{�`��x�%~Y�Ԁ�s�u�d��cf]���:}��wt��9��D<��'��5)��X��0KG��I��k׮��mWJ]��7��˩��K���;��yw��G���4�D�U�.iUx�I�#NdDT	ڂཅ�4�<�Iv���}	L���$�zG��!k�]xsD�1#���2�����J)�-�y��f!�lێ�o���X:������my�Oƈf[�98oo!���#�������r���R�>��Xخ��a�3�YDK#��������2��G�0ȧۍ�9<GXx��X�\%$������VQ*��uץ`�M�eG3�ssC�D���N�sB�=Z}�q�A~��[a>A�Ql��.�KI2����*u�����W��W�ٚ�> �]�f"1�-+]�l86�>�u̱��?-�A�҈�|�����I�{�+�t������8t��@1�%�����<�cN��fV��	H��ZV�����9��t��.���P��`���Pc٩�eogW��v�Y��F�="]C��i��XccM�����+���E�:���W�f�� ��{):p��J(���{�����[��/�r��Hj�
���P��Rt,��`ӡ�H�4��۠�=x��S�Y�(�^�t�q���s�z>�s'N���M�seh8MV>�/�J0��v���5U���0�:q�_̇1�.�#�Xxn"T�$T�M��-�9lmm�6 �������g0+i%G�s��/4�(�g��y��&{4=�L�� |�3�b��������|�D�3%�o�kn�`G@;!KMM��O��U&ogG��������o
�c�Gz�����Q���Ú}?i�Rs�)�r��b6�ዴ�s��M(ԙ!L�Х������ހ��xx��1[��>9~�3�gN�a�wZ�����RC�c4:?i�{��"�fi˓�k�;�����{�_���~�.\x���L�p��d�,�j��X�q`k�2��h���w�ɲ�u���AZ05A�N���|/Y��[������:�3��Z��!}�y�$/2$�H���i�= ��y���aQ���IJɜ�I !g���Nھ\���H �Z�A' ��ɴ���4���w���@a�d�J)@QV٭,c$�4X��q ž�gE3pk��m�+��c?h�׵f�r<7:�9V���3K�,''�I�C�ֺ��	�ݶJ��$�ɐF�ֺ�0��+�y�!��9< J��斐#UJ՜�ε�z�c�Ӗ��C�w�|$���l^./s�������ͷ�X&����̕�^�j��t8�IG�$^۪��rS��*�˔7�)�J�d�9�͡J���{����<���n��w�X��8��H�c���X�P��F2�2�5���@b����K,�:��`1�-�T��Zf�
z�&B���t^WG�Cʡ��2���ň�U�VtRl��itP�T����̄�E]���R�إB\|* w�=މ�
Ɵ�*��:�yk�ī������5X�A�v!G���I,B?�����F�돩w���ga�_���E ��"��FD��5��!ׯoz-ʎ��6��K�o��`��)
���:dA��.4���ʥ�n�? ��׵�����3W�a��S �����E�i|G.@/fU�.!��^hx*>��V��4�u4=գ��)ZXY����	মg�=̄��poSa O0ܣ��i��xB[�����kXp+鼥T���k� ]���W���z�Vidg�]�vVn#[=ꦕ��voN
z�j�ãSJط�P"m>1�R==Ӏ�5 �=}J[�н��s����t���x��9s:���<X�߻O�?�y[A�u��e�t4-m3���%���x^�l�;��s�К�zťa��l���s��a�A��4E'[�e�F�[J	�q"z��,k�+4J�&���t$p�9�t��r�e��u�ԌЗ�z����f��� ����h$ �6�m���3ǀ�Y���]ҝ�Z�|����R6�=]D�A��� ��`�H�w���x��eI�b@�h��+հ����x7='ʇ�ja���f-�U����q��x���Ƥ0�!Ŋ��F�W�*�CĖ�܈���na����!�x֨"].:��y�A9�M�Xh��ܹ#��H-�����u�Q���/�y��e���&w�|ޑc*���ܿ�ߓ'k�o����tHa �Ϙ|(8��́G�T_	&���v:}d���y��mo��Zɺi8jNNM4�O�x��g�0��O`�rGWhcc=&�B�J��q��X$ �C2�:�$��OQ�r�����z�j�Y����ǼS���z�T��`x�=��mѰ��Y��%��J-b	'ܪ$?A���9��P���Ѳ{��t�O���0hp��@�@����6�77/̫��v�fT8�<�;�/���O�i�=b��1L���_1�"k[�_�k����������w"�>���y�#[n�/�^*�M�'�����!�B�	@���3MB��T�`MTؒ�T�֨���ŀ�#�0��]��I��kL]fp+�����h��a�1tb4ܨ���r��Сm{{�փw$��P��a =C�,�*\o�`8t��#�0�&V_x�v�5�c �+
�̲�\��R��9|@��oeD�Ƶ���>��w��n�c\;'�%�Y5;YU 6��W- �i��Ɏrႈ#+1!�u�Y&ǹޞ�	�+� O0�����ӷ�~ßcK^�7~�����3�(,,Z,�,N6x�b�e�i������<	@R �:ϱ��d�� �]zp�ݽs�z8�u��o����&&�x�v�9�t"keِ�p�OA���O��`*��"6[����P_�d����BV����؋`n��<���J��$������e���Z�M����a��-���0JV��g0d�!�EJ_-m#�;�oY3�c.��,,�i	Xv<��e�JKÛK�A���xA�*�`��{�fx5̄=a���^dT�ÅvpM,�	4K��Zk�n��$8���|��	�Tj:\�����;u��nx������I�v ��1y�,�;���#�ۈ$�����+�K��`\�w����-ެ�d�$�w~U�$7r��M.��*~�pz���Zӵ�`��0dc $ ��0G#�|/�u�`�[EL�Î\��՚A�i�a%_��������9s;��b�Ey1���'s�v�D����P���A��G xu.u^�k��W�R�av��!���|��/��^e�����n�q�7T*��%�.��i#�-�k��1b�O�2�Nd�e~�5Ki��qE��D�H���5JO�Jf��#괵��0�@�Y���b�<_#��w׾c��A8𗯔������bαK��eH��#��X���0�7	���p�9�[y�6�#o�2�fe:�KT��<��m�7�b<"=w�Kn0���	�a���R�y�۱�B��`��v����zR@p �`ƺ]���vX��ڢ@�Ձ�&x����K��3�-�2]e�.�Мh��	���p4Z �;�Q0 �XM`ԝ ����e7"l�rOM�ɸ�Jaig� �� �6X���L&Cp͊�-�v���?�ާlL���������{�e�-Cdy��6O���s%ЋA���*ٙP؊۬ۑ��:"��ggf魷.��E:vl����ЁH�^1� Hܿ��?x@�>d��fsk��ן��E�e�H�������CJ�l�ӗ�U����!��/�;쮮ާ��:������bڣ��i��;&�O�Iu6 fq�Ը��-�k,&&x��>Y�v��壻4=3ǋ��d,�8{]���f����
��a�2v�)[�,jǶ�Jf&J	�Wh�*L�� �����,��n��ЎO�9���K�u�D� ��h-|��n�u˗��Za0I`W����D
p��q0�o�ST1#U�[��q�������`�w0!w;zj L���Ԕֲ ���R�HrڇZ������t�灸W)c���<Ҟ�����#3�S�|���W+t�ܛ43��ѳ�z���<x(r��]��^_�`��b��D'��- �K����FdQ{�����0����w	~	o]3�L�co���/�d�Ԭ���cz��.'`bg��y=L��g�Fu9�[�w�$Ӏ:��� nt��baA�s�[l_c\ ���R1���I�-H�}� �l;$#� c�To�v�ȫ�f�r"�`]qi��x�Oj���RH	��R��n1}�6}�\���0�<�uM׋݇�)X�+�*�y��|�S�ܖ�v�q��}4�/.Փ�w���"���'�ԩ�a^��u���U�m��P�Q����DFXq�X��KQr����	d �*9������8���+}ZXd���(荗Q�L�W塄<�E���U��Z�1�V"_�n�k�@*T.>���\���\x�|�	�z�T �=��^�
�s[��������P��a��BӃ��ya��ks�sy�yXU�_rd�.�Lw��Ba���M�`���a��C���ޭG ������4���<}�˝v�8�� D:�>;�F�6����n(_0�=�^�.�Aǖ�aϾx���%�թ�4A�8��ĝ��ɶJ�
�wr�K?a�#;��zIf�K�L���7�މ%h,!#J1�.�?��Cz��w�ҥ�h`�{a�0�k�b�B���FX�~��:}�ͷ�/�gND��t�LcvrҐ:Yu/�%�t�u���$�R���u� �ùwX��d�.}�k�˿�/�w�.��n��ܬd/B��@�D��=7�������A�f���~����*�y����۴��Bǎ���>-gX��q�t�߈��-��(c�%�}t�	]\�	���K
@B���'���ũ?qD�E�����W�gG��c��̱�a�i�s-����ŀA�����;/����j�b�w �`,��}-�-��t���>�����	��$Rt ���"�@4��.�`�ww_�c)�'�8����G�z�����w����� ���ꗮ���5�����/幣�����7b'����P;�}��GR��~C�S���ݽ���������?����}'����4ݺ}3�����\�>�{/.�x�
 
F4��wX��<p�^��cƊ�M[c�~�yG{�������czs���4�찈)b�������*{#]Q�����M�I���4�������q�	 ۅ�^tT�"� ��!�#O�����I��Ϟ1/R���R��PpJ�R�u+ ^�+OמHjq�M�1����^;h��`��,��y@�h��J��"�>%�v��T�N��aG����&?�v�9��O1; G�vb�z8�Z~�9�s��ڕ�֤�i������f�1�ȸ���ܪ$��.�8+�-���EN�r��Y:�r�:�	��l�}��猝�#KXb��a���Hܠ\Q�'��_qd�����Z cu/̓�{�K�S�K"/���I$b}'L�=��	J�>Cm9��0~T�;.�S�M	z{����Nj�m��˓:�!�R�Fx�^*ƅ��<LqL]��va�x������aND�<��T@�`	 �� "��Cx3':�Z�?������Q�c��ǂ�X@���0�C=5�1� *��' �\�'����a�T� �w��9�ZI��.LZ ��,G�6`ߝ����Z�jj�}?��O��`M�X��'lkѨ�	kdk�/�`G88tގ"Y� v���r���o�����
D0a�VkTya'��ՌI���G��ʶv�[�n�}c7�U�`('�_���H�&	���	��$����뇡A�ؘ��׿��?���=z��o��V���cKڢ���r�.OT��͍-���eƴ�lU�wC���B�&G��Ȩ��n!�ˉSg$���Tʂ��NIc��!�=��*a��('��P�=:�� ���Tz V�{��΋M( �AL�<	ve�XF�xb۫����فhlw���m�_f$�Әe��H�D��k
h��S�B��1�Bb/��PKedZ 
��D\h[��Q��y�X�V�<�P��6��r���M�2JL֒��](0f�H�|d�Ξ>A�<�/v��aL��]�)������1���7XC��#�'-�񼁶3��ǉ41�����p��狲��@o��Yl� _�Z�2Yʖ�'�fQ�Z��_�4"�g���1#�A����4q�ϟ?ǡ#���p"���^ �`O /�M�y��$���	�;v��ŹK��:KQ�9��0>�����g���U����A�gy�$x�U-�"O��q�z|@o&�8����w�؀i:�E�������w�9�F�(3��
�$�^%��w����ɐ@��"��	B@�� �O��^��2�O;/�?��Q_B�,>�,�q��q�u�	�$���k����h��ħAd'y��]�S����-�SJ.�,<�_ +{s�)��7����1b駶��6pt�@� ��\YT o;8M���<Qt�1�yed��B�f���%;��g���	���H v9���1�[�ك���D��M����ŋ ���l˃!G��1�7g�/���T~8=X:��az$�"	�![��gI71����tCFl^ё�S3%1���tfi� .���,���՞HJ7�:�`��d���F���������O"X���$* �휂Z폵�k���P`g!u��b9��i��laq�~��'���ʱk-�:�B��lK���%���y���Ko]��.^���0РG{��!OT�����ˬ8@��*͊����ɜ�RF� �Jmgg#�ӂ~��{�y��0x�� Fd6�xr�>pDGÂ�� c�&/� ��-��/@;���� NU��Ϝ�k#���#Kt��)����2@�����^�,6�چ��Y8�*2M	�:�C�>V�<���������rX�po�^����&?h���{��%�yd�Ff�m;�=�a� ����.�����ΑV��hA��3o��}��|߽��W��ffA��$=�2?{#�ƍ:zېխm� �㕬p`���&�Ik�����Je^�����K�����B)I�F ��~�n
<4k㛛9�J��G���5���'"�0PX��χ���1�x�<Vx��k��_
-��_�|��ŉhԢ�%��&��	��^ AKa��~�2=�4tjTY[�9^��yql�P�n,Z�̥����wh�y��_E�>s��>p�����,��'��;yϹt�ѡ,����k�7��m D��gr�Ν0��(O��hM����k�
�sX#�n#w��X#0�P��?5�+�XFi���_	{i��!���� �w�����[➀5�ń����tJ�{�$~�Z��hW����ϺVYĈ�-u�Ǔ^��)����I�%<�g���f�)X�ݨ�r�{��CϷkp�]���y�W���x�a��%��%:b=�A7R�D5�ܝA�T5Ǒ^P{&zNU�xy�-|xO�^�l�V�Z8|���Ȩu�8�49�\�D��F!A�����c;�G?FB\9Q%���9-��FD1�*A�Y�
����ԝ-s^Ù#��V6YO���z0��p���	�����v��RℲa��f�T�ሠ�"pR�8.��[X��R)x��䑠�[�=~v<2=��T;"���E�]4n�����є���+����e4X	ײ��NUc!-l�,4�"@q#���4�_x���X���K���/�W'���Z�~_fy���\FFk����Y촏�~�9N��,�(�"���r3��0eKj����T:L]r�A� ���r5�@_��O>�~�'X�?<|����/�Y���Bh�]�~�<#��v�ކ�������f�򠰂ɩ5#�m��4�	�eX���5�&�^��=��(Ϟ=X5X�VV7dk�&>�M�K��.��R฼��0N^���JX��!��
��t�K�� �&e>��_�(�cx�?���p�=fO�fUó,a�Q�V ��-4[����i&�&�gzr���,G����+��Kkr��uzp 8�� �~+o5U��-S�0~"ee	�nWSF|��@P;k¼jU�0��H�^����n���D��uo"Λv��U`��Bz!D+�y��ʴ����,�����z4T�2z|`t e�3�-�����#�yw�;�V�(�Kԁ������<��uz�`H�5! ߯���l��2i��_�6̽�a]ؐ+�>	k�=��������a,��q�g���vQ㲌Ik�9�q�~紣�!I�Пsɶ"SIخ��^�P6!e��ܗ7/�������'��{���(�&�mU�7�2�h�VF��q֘c/_���׫C_㾴X��Zh$7�D�`xbMA/:�0#����#�Q#� N���N(��i�̜��>�Y���r;�{~<�~\���o�x:=ZZ�fY�G������{�=/kQ�rÈV�;SC�Ա�RH�Ds������%<���z�7�{���!�Zm)JQ���������R�����3�T)��[Yꤺ�d])�0��Ү[F'm���Wt��fo�!���h؟MH7��]M<�r�Y�~�E��&u3�|�4�8��MGsռ���(��Y�cSn�r��^�@7�N� �6	��B�B��@3�6-��PR��[i�FYi�Az�[+PiZ
����њ��C�+�KT���'$�bX�5c�9���6T��:L�++M��N�͊u&S�}�7lR���¤��V�{ȩ�����;������:2���E-3e�k'�'an��?-��zM�o��s���Y)@ҥ�qV�t��+-r@w= ֏?�HP���t$o�hщ_��W,���#��	��I(8|����Gq�.����W�?�T���Sz�>|�I�"����bH���'�a~ɚ�)�d����GOh�����6���ާ'��x��j�{{�2"L��䳶f1t-�^tm��
av��5�\Z^��K[᷏��G��acXY�G��`��m�ͩ�PpJ��FA^������-]XV�W���[���`�K�+5n� ȕ����3T�Ӂ�zlUk�e G�B5A5�д��W�����Y3v'�l�98�G�bT�0�%�>�u�F:&<�AZ�eIr۸J�$�F�<�JA��[Ohˍr���HǨ�؇��g��p�Z��`AO4��٧����vko�W�`�#;�����B64����w_1���߿%��������g��_���"�q�K*w7�T�?�����qzμ����3W}�߫�-����;YĐD=& �:r��%���{��ؒ������a�E��%&����c;��}ɵX릖��k�7U��ﳪ���i�Kk�	�k��t�Tc�K��X#:�DZp^� �p��qGհ���������t�͡��2�,��r��\�f�f��E��rU`r��mn{������ES���z=E26����y�����@k�Xtxy��%N��X�l��;"��ص�t�TF��uV�S�E���ᭌ	��U�9��i��H�	k8��ϵt��)�k
1C�9���+�Zy�T�N�}�����������h�ϡ��>msz�&SzR�ZE���a�*h����ܥ����T��>
C�`���2�pp�	�	?5���U�pޡf�gV>QuC�A�:6������$,�9�|sLh�'<�o��!|���c�!����Q��jc3F�f4e���3�3����U�[��|)�:Ӌ�qAJ��8��֒�πs�|n�pBh7M��R�2��bR�f�v;a�Z�K9���DzT�[^]a�8`+�l���{��{��/)����<
`���B�{��L<y��I�Ȟ��������·�w{��|����aLg��i�p��<��vW��D��`Y��:E�|��8#} av�v�� Ć���fp|<���hb�����A��,��<n
K+c����O,����6�&�j?����t�QHvH��{w�#�E
$i�k~�ógO� ��ޛ]���A�ra:�sQ�惨Za�j^O��p�a�N��y���&�%(2	�1'��Mhx��
����P�m,�����(X1�pM�� 5V��\U�%ͪ�tФ��	ؠ����J�)0+�\�m��G��u���=��4�W�c���]篥{ٿ�#MNı��j�Ja"<�%zd���[F���f�C~r5�+����;e!�9��o��_���5�ExoG�w�k��w��)cIR�.��8�����i���yS.�"<{^W�q�;�1g�q�j���+��P��V#y�Q�W���D�Z0<�&�i�k��Y|9�:����|sܰ2�������Bg�j��cT�Yg�v  �=�%�C�he�Ɗ�m�X{4�w���zK�6����-��x�ȫS��,ŌI�&��Q���ݝ�<Kw��Ѻê�u�wSi$�UM�qU��]��	D�����	2�K��X�l��y�Ҁ,E\K��as����drr{e�KZ)��v��/3�p�b�y��Lk#��^&>F�h��o2�̌�ƪ=�V_][�C��W3����gs�#��<�VUQ��PehZCo�M��q���`�,�x��טg��2����`;4�~ �G
D����5�P���a�s1l�h@㎀GZ�<j��ȁ��6D]l.k&V�0�.�� C����Ct<�#D3DGc8$H�n��y�fib4�J<�k�T��%s騬��!΅�H�'黱C�1�g�����G+��u��}'S5Z�U<s�d�9��F@�x��"w�D�K�}���0K�h���~�9��%�z�d��x� ���*����B)h�
EMo��FZ&T
9����>���)<��P�:�%���2]��/¢��Np߆�-U@
ٸ�)7��r�3��CMjҥ;B�Z�����:jV1���;�ͺ6�Ɍ���+W����O0�p=��ȼ}��'�:��vwwv�@�o��G?<�|A�!��-���$ri���u ����������
 �����֯�����/���W*��P�2�Ux�I����nH�<Rq3.�����d�@���I5aE�7h�x�U��ֲ�Xbx�d�O��J���q��o��QY8��[^Zf^J0��7MJ�y�S���c �#��mOXy�#��8G�)b`,!���뗔��۽�]y���_x�2j���c�h ^T��$?�B~��_��W�em}��
���8��%&AVp.^��&�J�C����w7U}p�;x���j���rA|�6��H��M�,�Uw$��a �%�,%5�X(;s����(�������֘nt���FA�~�֤h)��fj f���A�d�( �va�_i���E�wǤ�h��\�`���R�~��\	�c!��J�D٫�YUI����k�bF/�+��s�&(f�7����?]Gç�芝��&�^�;79�FyB�&�R�X���JEi��#�!Z� �������M�4k���h*M�{�>��(��vD쭹&v��,>|��zdM��<���X�J�k1�_A/��9��� �ܭz$�`y��U�@�V� f5,Z�t�
���~_�ǵ��?Kz�9+�e�IB����J�@�hc�l�ȑ�.*�SF�:M�Q/O��ئL1h�����z�t)߂+g��S�@f$<�����	#4�h�Y�X�A�owk�a+&}�4�\&�y6ͮ��
��
bٌ{v&rϮ�]�\[�Rl��L6\��q�T��H`��D���1��
��b`CZ�'�ӍF����w(W��YD���^"=����Cy��F���r3 ܏>�HVV��*T���4cHj���m7�/@hZ����������޽{1�I;;�	��.��/>��Sz���s��E"ڲܼq���i�u])}��dai�\���	n��Ƈ��rVq񮛄y�����&��e�����ڊ��ޖ|��Oeum���������o��2N?Ћ$3�s/�fr��� ,|�} ��̆G��+���
�]�^�
!������c�q�@ub:�Ns�JD�E��[�̏�?�{�`&�$	l�:��o�	��� ��5������F��WP�R���E׵p1_���:�i�r��oS��v�
r��e��
��{ld��û�?��ho�&���PZ��<?��f����b����{���{n@�y���C���>\�{�7hN�q���k��F#C�m��������y�\ڼ�Hǣ ���/d�k׮��.����!y��������̋y��XJ6��4r� ���y����d�g3�t�C��gQ�����Ttf`	���J���@!<������iS�*�U3�z�4��i�.�ُ|��k��ӱXK���ܙ��Ri%*���>���m&�����+e�Fl�Y�xeXs�P�<�g���w��x�.q�4z�y��ޙ1 ���.�m"�"���<�^�6���s z�Md�n�����?Y��9�h���1 ��g=ga<���L����T��%J$zu�ᜀL iq7o1�0��g�QX;[b��ԡ=eퟳT��ϵ�\C�u46S�с+�Zq�e� �p�(2���3�1��@��e?4B@��,��~��K���詚N��`?l(�0����X}{ό�xa���	E�oZYҋ�Ӑ�e�D3��:ht�9�aю����.��:�J�ݕ���¯�_E��fEh���6ɥ*���Jzh�iF=a���ɋ��q��cfX�}�N��l�gO��B�IYxP77r�t���(�%�̪c)O��*7��^��D�
~��(;G��I��z�ҳꋠO $�ke�̛�� ��� �����d�\�`�B��� ���/����˵��,�?�m;��zJQ�����ߥ����_рi3�x�%�U�=���Ih6!7px)�x�J����*�1-4Q[��(��%*C`����WϘa��@oZ��p��֢��6y3r/b�_T,cZ����p��p_nݼI�<�k�H Z��#�bm�z����[��:��Ą�B�>y��A �#^�&`���zX�"�W��z��.��P6Y��o�p(E�`C�����?�8��D/�Gl�����u�Y�񇄴u��?UE�/1i�f�/���>0���Eh~' _��~���5�[��|������w���絼rF}��`(ݼy�����D���<c�� ������y��O-�m�,l����ø�w�hX]]�W$a]>:�Z^0�0�.*���9B���c!�׶Q�g4�� >�`V�pXl<;Uc��g����1����g{uk9����>I'�B"���(ő�� 6�i�~d�K����%ǺJ)h.y�9ثX�J�hB�z]
��(oI'P�^`�Ƴ��m �{O����п���;O�Զ�"�X�>�;EV�;^��m޺ǝ�{�]�}��9g�����"1�$�n8�g^�%����[;{»*Ut�S*���(o���>�ܺ���h�,���Pea�0�+�����~�E�C�>�79o .�#ٴ-��]$�uȑ��	j;���ًp�[�m/�*����g�d�t��_�?��/���@Fa��fx��Al���S����5�fL���U�a����!ת�G�x$>6�c��ӣ��ż� �T���l����:c9� ⎏߰�XF6\[9}#X�c�o����[��h��ԋ��;��Žh�Uޑf��S5�+���T�j�$�ǆ\���B�I�r6�^x�s�����5p����p���D��z�ܛO�so�����O�?��?�)?�&Op2�~����޽��.]Z}��y��({���5�GO!����&G0T#Z4%�<�T<ܞy�Z��]�eUՀ%L�iH�p���%��Ge�!� ���%&�ֺ�0 �6�峟~����_|.�|���  �D�Ƣ'i\/�{��G���Ͽ�f2��V
���}�>��Z���93�|�����gy��9�Yy�L���f�wD�2[�ܹM��[�n��r_����vG��������?����������P>��Bp&M%:����4�<�������7��ս{�.�h��'7��t6C{��e8��������p��l��Y��.�����"��E���C�(6���w�����ȗ����������'�|"����p	$&(�'V�Hy�����}���)P�7!i�Q��c�u���/��!�C�b�pl����}���e)$�$����0_��G9}6�z�5�T9���i�y]��E߃���@qY��E��j�.V1�3M�Zߋ2`�'4��m
���sytX7�ӈVk��Cs����h�z�N��[;(Ϸ�����zq�Ѿp��'x���u����}�������V��C���pH�d؞<}LcEF o�;O2tŜXf�9��q�sg���PQr$���I�%�J�Jhb����mV?�w7����o^���K<���`@�Nȉ��Q ���zج���ko��! ɗac<�8���}��>��Tc�bX[���n�|�l����,�E5~q?�e���m˔o[�wM��U�j��dtD}ԃ�C�c�4����1��j��Eqڠ�,]�gXH x�6v�Y�+��b��@h2,ssvP'3���l3��9���KN�jff�ϖm���B�R&lFlO-�xH!�^�#z���|/lf}�����[&|���C�'�t�޹s��JTS����"|�ڭ�-�w�P��J%�g��
+eu
r��q��'��׿�%?�� ��V��|��r��A�ޝ0�i��
cṴ��T AbK`'��W>\t,A��U��  r����5�f�8�Bd�p�<~�����=�ݖ�jG�=�!\�S�Q�0�Fr��u*;�e�I!���~� ao@/��Bu�d�X��cq�$"��nn]
} �˜�,wTL^(M��:	�a����DX�( �4�Mb��.��k��#AԠ�Ҧ�.-˭�WB�,0���kM��oQ��/8� �����oׇ~O��a���H¼�F�fs�����$���Bc��B1�9��~.�G��z���p)��-&cT�ϡ�`�t\?:B��^n���}�t��_�����M�Ub��t^��ۗ��H��/�/~/O���v+�7�?�çLJm�`�:���9��mY�:q��F�8?��/_ȣp�7��v����!�!�׷�9���y��i��Yæn6���Ϫ<�PJ ���Tf1��Ѐt]oӭmj�'皹�9����6�H�<H�UHՁ̇`�WbG��Ӫ˫UD����a��zBUs��%�|a码�S�[�U�SO�y=�|1q��e��s��� |�Ip�5��3>�;�P��v�|�Q02	�N�HV7��FL8A�ժ�����1���_scc�b#c��0l~�&A.�*ث���1�!�����C��>�vqcHz ��^T�	�Q�����~M�^?
��l�~�{Tх'8@�^�D�{�)��\�~Й�ɓO�(�����Ԃu�Cz���[��r)�
�ݝgj�j8y@�䃽��w�����jrJ��Щ��7\$8�%�ͥC�:�אgc�v�;[ϵ�L��Fl��{�Ě-����ܙ-9�d�z�-�2V�����΄�����0*�; {�Lm$���!��hx���L�� Fk��É�&>9,��q�3���*����5��3��Y��XS2g�B��*����Y؈����˿��<x�]8�.��/¦
� ��6�r�X!�^=����BSB���!���[t&�,T��b]��tɒE��ӂ|oH��x��<z����*4�G���5?>B�}j(�~����*gG�G;g������dK�S��X0��$�^���=�+W�%2ǼV�Oõ�B�����	���D�!֖��;e�Ci[��o*J��&ѥ�˘	���	��	*q���ܯ�G����f��W�N�A�߄`Ŵ~e@�[��� w �ݰt�<7��7���rٚ*lX���=<��` c�F�eM$4o�h5�����]�)�����������T,J�|��W_Q���߄��&�ە `W�1|�k�d���^��amV�iה�g��(�~�r��5�;��e�j�lo�h��X�ʟG�gv�}�����ohO��Վ��ﳏ��ip?7`�t)�}y�vO�����Z�#��<�\V��D��6�>}z-}^��H�A&�c��hݰ���������^"���u�k�4��^�qठ���dћƚ���p�i㥜5Rkጏ�yM��p..�E���ކAIh= _p��阢MeF�˱6ҫLZ�-4����-�d&�^|o��_��.Z�A��#Ϧ ����:�9�Ș	>9E����9�΁�z� ���CYZ�Mܬi�>l�Ka1�Q�����BE�k-����IEK�!�7*�]c2c��r�5ym�% E����[�㙠e�� ��\c�?>:
`�X�PR�8��E�+r.����,���R� W��
1y���%i�j,���Z��c�A���gͼ��U������
 <k$r�"�d��P�f��)������ӊ �	`࿪����|�����o+x@��p;8Z��u�y����O���(7P�E�u���y��QV��c���Qn�õ^Iǐڪb��|��/�a � �W�\�gw�f�� ����ˡ�*���?�8������Bb~�6�JQ��7�6�9�L��uUkYI 4]�#�I7������ Ŀ�l""�ފ<y��HD`e���h �_��O�/?��Ka�х)�s��(ߞ��0��+Zw^�ӔO=5Q�곳��t��Ə����D�2������;ryk+ ����U}LB0n��yg������;a��J�^�v�G��ln^�e��^��,�!��4!��n0�Q�Y֙���Ϟ>�A��R��g�&�N�N=���u��v�ʫ`�C�nyiI��Y�����|����.:.����e�谐Ʉ���������*<+�P��g�ςg�M�5��L,ea���,��5֯Xej)�;��f�k1���.��J*A����zj��IVeM�̒�\�E�����*
�Ŝ���ݔ"1��8߶��'\��������RQ�.��ň�ל"�I撹g��&��k��&F!=�5�.VF���Y�=���[0�?��p`{�W3i��0��6EHY�,��u��r�t�G����j�/�63>.�L,���Q�5]sꅾ�z�x�`���ׯv	~��E��ll2!���P�YV��N�A�m���K;�l��T2�C���m\kh�Jm��)f��Ϫf�V6*l6��2�`"�{̄�� |��x*Ӫ�d4���{emKֶ��?,�OQ����Uټz]��\ ������zE��&"6ǪU����D�&�� >m���V�E�߂!i�Z�Y��KwB[^^e����po��j/Yዖы���w�!�Su�Sl�3��✟X>��X��'-�ƩVq!��`F��ٖU�j��Ѐ��d>Qk.�;*f��YM�G��W��Dx��EF��ƚ\��� $w��֡|Ѻܿw���?�ɇ��-� ��������VM'k�i�}���F�c�Kyl�B_�|!O�=��^ڝuNH$�!#OK�½��@��^Q-dwZ�Z�+�����'{��t(�����D1T�5٩ɜ��y�Nj�����͸a�G -�E/I{Ҧz�1�����?	�@� �s7Ng��h���Q�_�Z!���Ͽ�KOVY=��)��J	�p��`��)io��C.�u��̶���HN�D��-��������Km��}2G�aL�J��Z�r�I����tiS� x�W�e�cF	�^A�7��t]����:s
ZT��{~���T���6";� ����� /����q0���Ɂ�QXi�d�}?R�_���]���[e;RۂQ38ړ��'���e���ۖ���s�!�2�[��E�{iZ�0����<ؗ.",n��t8Ug��my
i�*��������}���F`R�6g.NSI��""5��K�}��f�w��&EZ�I�J�Q���T֞���ص���ĵαFf{�8��V�t��Y�(&J۾����ZX[�����ڱ���'P� m�6���4�mr�;3�=c���2��5��Ϝ�"�W ��[ Kl�Lf1��9�:�i���IhU�ʆ������B��k.U�j�h�F�4�^�һ�.͛_8�˛ZjIY5�d�E�|f:Ȋ�S���"rK��U��d�	��!��ef�~� ¡� n��&X�A��_=)�¦u;�|+��E�5����dc�ܺ{W�a����p��X̡jOZ�K�2}��������H/V ��uo$�y�wZ &eFE�V��hRa#,�5BvZ�
�K�e�҆,��B��J���W�H��8��@M��{�$���<��0�R� xi~��lE���2�	hTzY
�LE�� ��ъ�R�ٵҘ�-`�����s�曯���'�����V����䓏�᣿��7{Lp��,x?��_F&	��0 9�>��7�����y��M�V�(����u�Q�R*�?@���~M�x����<��q+�S�~ ��9��f	��+z�qs@�f&ɃD<��{���t�R+��3^�I(�B@�2�,�ܺyK�ÊU�T�N=�1���Pv����p��&�y6�f&�<CQ]D&e�Z&���/s�}���ԸE?C"h��{�@��wW�Q��|2�`�mn^�+Wo���ن�B٠��9��L��9���y��߲�0?���X���iH���Hx]�����)[���V��ޑ��F@/'wCX�.��Q�E(U���#jj�/�Mx88���^f�~�=�h`4e8�����>sVjJ��H%�e��5Eq�=%�2U�W�	�cFIV���F�r:����~���'���s�0���UD�Z}9�M?��]�Zc������j3�Pa�]�{� �l��h� g��Y��#g��`^�,�|:V��}���l����3	k�M�jU厠��)�S-C�{%D�V��Iu�����L���5}�d��6%9E���^<�˂�1����q]!��E�R>��`�E�Y��[s�M��u����ǅ�_��Xt-|;q�����ҁ��'�@ﻭO�qGR��˹���`aM�9�!�HM���>�̦@�y�%s�������"��]�6мg;K�?sZi�W��X� ���ʽ	7P���M��p��AGTH��Ģ����;r!��!���)��E��� i��+���Xt"ˬ�g�ٸ�l�����+-㔢������+���xu�����-4u�1�P.T!�W�µ�/�����7�ݥ x�+�a^!Y;�	�	@��Im��ؼ�ᡡ
$��pj��M_dz����'��_�Fa��\��N��u�}Qγ�ZC��hE+��S�GnEC�?~�D��?�3C��	�{�܄MpyeE��{_�7G4BZ��@�><:��(�RĿ�/~�%�_�* ��Թ��7 �͸��K^�XX���̒�� ��G���y��	��,\�c�d���s��L��l�x}�
 mM�����U�KZN8f�6f�vL��o�M]��\�u��5�2�5,H��R��73�
�V1�I
����T q��'�i�cPP}���W�'p�}X=�-K?<�������o�ED(��R� �����օ�ɺ�uIz)Y���aN�$�h��X�w�PE�r�zx퐋,��sg��+$��!�<�_:Љ���i�����F�j�υ)��_�ɪczڏ��P�@�c�x
:�R���H�|�Q��&=9:�e��1	��E!�Yf�,-90���� ^P�:2iM��X�Wx2q"�d$]}A��#�:��M_�TI��������j������[$u6�{���n|���l�����*�zt<���)Z��XK�������7�*��<�9t ���{!��OK��Y�e8N�Z�vb*P�p�����>�����9p{6
}�#^�<��O`����3�=�"Dv�Г}�$q��pʙ.tx�;.4ܒ����|/�|�����<0�v/�Q�M��3�f�%�^�$ݟ��kњ(��(����\^�$k+bh�����`q���2D�\ެa�4�w�P�}p�+�^O��Rx`G�x�%ȕ�Y
�zY2&�r�S1=[��*2���p�b�������m��3�"�j�b��lye���E��h�4#WXj@����=��):H�gl���+t�mSt��R�E+�%>�q�������L�A=����,x$*�b6��)-Y�z>l� G0T �����6$pAA 0����۷����=�o����cȚ(g����������o~M�N�)����R[\'8���c�3Iy�J����5��^+\� �Ⱥ��GѶI��;�ѣC�\+UU�d3���z[(e��kR^@��䛌�)��1!�&�Ԣ'�7��cV3,���^�� ��h@���_M��6$;����|�	A� {-�c`�PK�&�}��U�V�6���kJ?��}��6����:��3��kÐüQ*seޞ���i&��HJ�NT�	pcQ���h?�p��	��#x�����x�-U9�,7�� �	m�q�ú��BZajL�2Z��&$ʮ�p�1�ц�:$-k\�y-(��FXq�Ll:�T�+��^�ҹ����T����&��фm�7�Z�����N-鰎��,��
PHS�T_X# �7B��Z��uJ�1X2��<�@��"���+����W�Z4��87��@oz�z'�|���{6@U$������MK}83Fa^����(Q�����h+�V^!L�vŪr9v�j����k0�H$��<&�	��`U�iy7�:���H�*yo/z�FĂsg�~�>��S���r�h�<�����^�p%��Ef��c�Re�qX5*W���5U L�W��sϽE�[� �?�(�}���5L-.����9�����S-�|�&�,lJac�Fr�P��+Knӡ�ګUX�F~��1�<�K˚��Ѱ��n���*�O��p�>1�ʫ(նP��I+���]K��!j�Nm��o�3\��B`���|mM6/��&e��N��f�vj�v�[��V�H�k�E�p�������K 6��ڀn�yz�3��':�]�ڔ�� 8����+1X���v�@"6-k=���lZ��h(�}�0���[�JD��u^[]#w�`f��~�YE���O���}/?<zDuxҘ�_t���i "E;=g��g@�eܗFk��G���>��ƃ�^X{��ݕr�Q-;�u�|�^*��G�C������*�m+�Ƽ��ʟ��ՂWrj�9T��V�cۼ��n�l\��v𒍰Q���pP/Zz�S�4��������* ��"cI�`���о���!����v��ݺs_6�\���-�	6.i�X ��#9z�+Ӄ#z[���&�K�I9��  MƐ0����p���ЯK��qU>��?�{�ݥ��E�>{�4̭��b���p/ZD�ml��\bJ������E6�x�2Za�B?Re�*���!��On��cc*���C���-կ�X?���Q3�U��_�z�K������ ����게�e>�(I�4p�����4mk�p��mu�<l�am�N��0t@�iu{a�h.��H �xj��bg�_�+���䱙�X�)v�680�p*�KA�Fi����a6�9���C$��]��'�IY�Ae��74� mȊ��+����@�V���J�u�#�%X��`F?�n�iTvj:�*e���$��Z0~W	��Q�]�3]e�8��O2u���̓�?�5$ג����sr9��.v��8���W/^�����|��sX�L�'��s5r��+�n�A�=	��V����5}���V��IbR8o<x�߀.����ۥ	���(le7�A�
�a�MBL���C�+����<d�k�v!�_�/Hm�/��<�T'�z�-�rCy��yX����=�~FI��~�$��Y
V2S81/6 a�f�v2cy���h
tq-���#�Fԛ�R�w g�	����W���Q�mOt[
t�q"Э�'�o��2��<�׭������kf�z�P�v
���F#�y��Drҫ��Y�
$��KO��;�p4;_�z@ؐ}�n/��S=ыY�Vl�
�{՚ҡqqF2�`d2i���=(g��9D�,�|e�rJ��0���:-M��,LSS�HeZ���fܔ3�l0��ʳе]Fͯ�U�
�l�avx��E�L���9�Cm2>�-:j��&Q�a4T
C�J���P��fx@rؽ���g������}�|kT��>��`���?�V��8���m�h x΄���e6��J,ҁ9U����{r�އ���=�L����a(���<`w$p��`U��f{���ra`��Fp�d��D�<��^��P��y�o�i�&f��r����U����y���p��_������OFy����8[�ؔj���$�-�a ��w+���u*s�Ko���|Vt��>��?k�R�#���ɸ�[�r��3玂����\�N��{z�c�ǘ�쌆y~�3�z��Jd;����}=�_�HFB,
�Э���u�a�����;��_(*xa���x#x��l�*=�HSGQ�B�pX�1����`���a��e�EA�z�=�%O���'���=Nis�|����Zҳ�%�ԟ�@��)���9 n="/�� r��U����)PW���>�P)g�'�:z,��R7V�4Z�ݐ�pH=�	�5|����7yX���4�R�3�>����"#��l��&�%��ln]������!L����u:�d�r�u�E�-+��\�c�/p�4�e���3�3��
F妶:�5��kUY&��RK���I�z�ڬj��t����k�P,N冲\둌��o��y*�E�q�U�%3u��L���{��'d�<��=�{�B�x��,����+�EX	a�{վ��O*����!i����k�>��ϻ�B++r��]y�j;,���ٳ�Pt:Z&��$���e&�h/�7��d��Ĩ2nv dT��rzHW�.�T�(,�c��iei:�X�o:�Mf��T�Q�Q�U�j3>j����DF�,��k�Gǵ4Z�p�b��QYV��k��������Uwv�������� �����d-*��7�������Ln޺�*e_}�����c�&�S�Q�:��L������	����`�M�)�_�[W�޽�峿�� �_��	���`L�����e�+|�%�!�Q�BQ��t�K��g�����v�\�A��q��ܹsWւ��	d����{E%,����3�U���r��B��8��v�	�J��~�pl��k �����$�����B[{s}U6�Wd�R��u^�v�Ɯ�ZU�J"���!V��?� M&E>����&֖�`DG��$�݉�H=H��"�'�X��M��O�7�����_��û�g�6,j��k�4 ȼ\
rF���=<DY�=㡬�-�v��X�z�������"k��:�J��L�ȫ��t jy��P�*)Hd�^�&a?mk�h���+�?y�-�G9�����{���z+a^��E��9���򵫲���$iy�6�2�/��C�iY����޷��{(g�x��,�'Ķ�+ⅰ30��z�$�`o��k)i���yM07���ތG�� �X�l8�F��si�Ym.����]��WW/�ڕ`�c��b�AL���Qf�V���=�@� M�Q���yL�La�T�E]�j-HF�t=�y��[��Q굞0L�QI� �=C�9$btTԟ\��U�c�<\�!��(�=V�q8�1����ѐ%�8՘5��Ӗe��6/��w���kzo��ӱ��0�m��V�`U���p�T븑t���� p�z�����!���q� ��<�U66/�իW���kr��,L���Vv/�&0�4ؿ���2|����o~KO#����u��s"6�F���s�0s|jR9��-�ä߫�'P�;-�L�؁�Q�9Ӑ,���}�N�^ڗn�ef���ܫ�i�L/��̯��Lm�-Y�{L����-M�	�GE<z�C{C$��_6p��al| ��f��B�Kx�ɧO��>y�I�yˮY�ڸ��T�ӓ^��nW����xv9v�鋪|~�Q/�9�pM�6.iu�,g���n��sW⚠�e����e��:��0�oܼ�(�n0�0&Q������@�m�>ȒS?�)ѵ�S-��u�@j����^z4���T%x�KZ0���˕�K2�q5�|��I��Q�$+�#�J,nmn���D��1�{֤�hY>񒹬�TY�����o���l�\$1�"�����]7���)�tq
�/
xO�|O<i�vg�v�9&p:��%�{a��Ơ�F�]_Ls�k���f���w�0f�K�B�{/웛�ub��զ�תt�ڊ�8�#�����Q�9�+$/>ϷG�w|ON���h����-r���E?�k��ed3/�p �%��:�G�X(V��0kX�*~7����.+Hu�뛬/"�[��a�����*�Q)��]eTXx$;f�y�z�0IF��ԏ!:�ʰ����ޱFK�c7ג�ܴtcq��篸�N�w�ˑd����|�����Y@�	�a�v�0K��X4��d��j�Y�^�G�[+��&�364����,�����fЕ �V
��T7gi��_�V��r���@"���#d84�c���1�*����Tۤ��@��8�U�PKU�T��̂�A�V6!sn��2/b����w�)�O����Z˔.8�H�P�=�έ�j�WK{��r���|���_���#�pOn߾�� T�¹+�o��8C�͖-�}�������_�J�<y��>Dgxj��k�N�:��M��4`_����+jM��<qp��[�H��dNm��*���=}��\�H۔}f�̾yh�T�mUG�4�Q� =IG=bXh�=P��C��:�	�d�~�L�#}�� �6	N�&Y0d���Ő������y��a��y.�`x��G�ً���aSe��0t�___br8�X�0V�����>�{��; ��wn�͛�y~�'5٣t�L���z�cq�\ˏ��;�\�����}���/_�`x}+ ^<0><|Ȣ׮_�k7��ah�W/�e? ��/_�q�+$e����&z2���{ͻ�����*8�s ���h_n�ؒ�+[��O?���ߨ 8�2!*�F^gf�7R�b�*�v�5DЇ�x{���up�1��3�"�MHfZ�n$ʉ.��{b|�X�!}��;���JCz�цິۿ�?������8�ft�M�4?wv��ܖ�ɤy-�"��۞��\:��ɢ�k!=m0f�1H5��`O���kk[���EVA�C�w��s���4F�J�24k�_��#���T�p�E'�L��3�w�3�9�|�˧|/�uF=�u�X�l���MI<?L}�:kxgs�Tř����fI�T�%�&�o����i����_�,.�6����:p2�8jf,��(�	?������A�&B-ʒ��V�Wi�_�ޞ����ٖ�R��0	��¦=-�9��f�k	ܶ-���.����:�N��[X��d�T��q{̊ȩ��wz,c�d�Bt_*K�D.d PF���]n��Gm����n��*8J����푌Js�~�3�GY{���s���k%.��LW����J<�Sjk�җ�Gޓ'�A[�x'Ta��|n�� �HY�����3����L~��� kk��0T���pwC�������I�qЃM	V�i&|S��P�'Kx�7iUǶiY���Ϝ��u��*��_��s��p��ۮ���̫5^�t ��z}����<���N�#ʛM�ƙ�ͬ�&����6�!��7n�����r�@�_���m��j���i��� 5ŕ0@Mq�1�˅f��^�|��g�o�kow�Ɋ���b����Q�۷��u$����r�aa���]�}gNx��G���k<'GG�T�@��!��B:�n ɈR\����:@~\k�'�r��Y���l��8f�����۔�r�Sz�2K�L�.3��,�0�����,��=�ȡqL�I����xfBb�r,J�S��;9ڔE}�[tT
PK�Z��{C�t�u�*��Xp%���G<���,�^T
4}B�H��~ :B��^{����������$�����5�v��zMX��>��9pAn�w�}pf����_P��̀�,}����v����<�9ǏxO�p��s��G�r�k���bё�y�H3��"�����ܥ��{�J�SR�9a
;<�X�&�(ǵ6��(��5�ր���2��K��Jh�N8_K����M�� �Tr`�p�"ٱ&��ic��'�� �>\���� ���*���л�k��6=�˹VZC����p���]g	]pw��v�<�j;z�n���yN��U6e-��9�:k����^j�20�Q�`��f7?Ӽ��^>�є�y��r�2��ݗ�O� ��ͧr��-& �'�`�`sh�XI� �j 23�P^�zI���y��� �I� �獂{�.vj�Ƶ5�R����(K�5o��E�b�I�"sx�2�p�����$K�H�X����4ٍF�D�<Q�}���S�T���W(hlmm���� CNf��^7x��D~ " F��8�Tjȳ�v�]���ͥ�K|�Y�8���7,Z12�3�;��{�؀� �����Ƶ%�F����%�4	* ��`��	���A٘�'\?�)��Ïem}��W���M��=��n��L{����#G�{XP�Gj���j+����f���x��ݸ%^4o��3���=�z�^��|��j���è/����C����>�H�Υ���� �M�P�u�-�g�%����<�\c�}���L���G�W3j��L8�k��>�ɕ!R�[D I�pX�0�ߋ$E�����2u��i.b�g�{�����`�58��w��Π��?WO���_���^x6g����3w&��V9����*�fn�"C*nxo���=Do�S���1.�&��	U����፬ljvAg�^VE�e�m��``�C�S��
�i�:��j�"�o���?��;�^ ����I�L�%����o�lV��Ť��s�R`�QЛ��C����٢�1��V]��Ed�C�5�g��v?LH�X
���&8�^Z� �.I1 '�ln�����+�7OȌ�[��:RR\o���>��3�S��ն2�{U�8�y��=xbU��@��W@���v[k׏��_�~��|�������������~ (;���cz��#��r�4ڔnH�����'�������3�}�R5K*�˵�[IMK�ZV�D4�h4��L�K=���`���[7@�IbQ/n���>b�If��D�~�n =J�	y�vϵ�� ��6�����,ͨ�*q�W�W��������ɷ�}G��L�v�ܺq�:�߅�vvv(��a��k�"���dL*�^�q��*F)�.�{#�	�-P*�H��W�{�Ю������YDN������ʣ�˦׻��"�����mFl����a]�����g�3�=&�W�ڢ�i\'����1� ڔ6 TZ)�F�D=���8t9��p�4~���O�:6r93Kud�^�3U�ܟ���\���S=��(�k����'m���[Rro(.?�z�,�,	��SqMmG�
� ��V6��5+���LKg74J�~Je�m��7��)��6,G]�~/��7M�-�Y%F����y�SÝiu�x)?�	N���c����^jo7O2�u6��3���2an�Se���~���Vs��>=�=;iN=�����=�7��W�*z�Xx��j&��CI���B֘,��p�M+?lt�o�Ti���
a�/�[j����KK�$Z�e$3��}�V�+��زBU
evP�Z¸�	�w+;< �T�G	,xr�LL�Koi�%EṦ�!�{�Yx��N�*�X� '8̨�[Zg��ΰ��5`�����*�5}~�����������k���l��ן�.���49��+�;p��<@	�.�f�������} G�|�~�2&#�fKb�����"'���ٓ��}��$�U���oy�G�t)��<y��75:D"���G��G斃���CsR{ۣ��Cl!~C�ғd��"�m�ӚkK5>=T�B0b\�H�H�H��]�N)�͍���5R����m<���	8ax Q�Wb��k�v���"�6�kt~1�U3��txȂ(c�:�����S�h/g�|�ib�Y2e,�1�IB^f��\C.�����0�}k�
���i���^����k�wṽ��*"Y��iz��T�Uit�&'iE�_�1�2��]������bI����N��jN��5���(�����}%�y^	����^��R�9���!�->��O��R��|��>�ை�|GB����w�|x�#������k��R3BP��Ïz�>������7.ro��9"�ܩ�8m}z;\�[g�]/x��H�M�k1�K<������3%f�����\��K@� ��OT�ۅ�ЂV~.=����6����PC�J�k
��/�yv;�h�&K˗(y��(��ת�R��e�Q���&'Q�E�B^��`S3�K�fO(g3�{�*��Y��24#�o� ��J-H����0�2�TV��aa�Duv��ڕ�Q��P_�*]�穎NA�Zh8L��Ꞃ<+�c����5����QEO�k�z���,��ܹ#S�0�a9��h����w�;y�k׮2l��eD���k������7����K*q�K0���p	_G����Ғ�ftS�rvL_�@�q��䢂�l��S���w�h$��\Y��H�ʞ�6<�~)1q�o,�$�����9���ŝ�n��~�po�ʳ|�*�4����K�? ��{�5�b���KkP�x���x <88�g�}�� �0���,y�D��6�V;HCg��+��7�|#ϟ?�B<�7nܠ�e���.�4>}����[>w��oC� �����cP'\
�o�~�ʏ_clc�\�|E�ܽ#�n�
��5&ʾx�I{�(Á��z Q1'���YZ��>��N`U�0
`@��QzL&Kt�(4�ɔ�s�D1
Q,g�����W/�k�ࢥ�'��K���*躼�ZMf{�"�yj��=t~�s�a����;�
�o������&b�#��jTa�QYRƵ��U��d�x�8O*w��U��;p��(舭eu��Ɵh���f���ŤF�[4�	�;������8Nue^���P'����f�k�jW� Ͻ8��1Qj�R@J�U!��QE?x�<�~�;���j� ߏL?aJ�xQ	'�66P:�Q�)<�f�&��<��{�����j�l��ư�Ӻzx�m#�3W�]�~��@�L^�s���F��*^�N�^C��p����oI��Dx� �����$��i��*��lH�Ѡ%[�����3L��8�_),C
�Y��iK3�g<�M�sɽM�`�X1����٬�����W��͹,�l��8nM������)2xr�_(ʥn��h�"�]��f\<�ؘPP^���]�>[ٵ�'$��]�&|���a3�D]�H��vS9 z �� `��FM�vWG� ��@�`�����'�U-c��w�	��w�����a����=�b��8�E=f�m�ܹ҅*����0�97|�	־�4t%\D?�#B����g�d�<4xQv��Sn��<w�"��r�M�<��9�]�g�>���Ғr�����|��W���u*+|H����6�6~�	��e�����^&��   ��� :�6x��ެ��@{�{�t�{�ݗ��ˌ0����0�$�)	�Is|Nb�B��G
��yZ-�_s�������NXd�VXGѮ(R��}9����,����UPdc�L�q"d�g�����V�*�L6����y
3V|���q�J�E��5_X"�n�N�݋��ٝ��呂�/�b�MB����ƃt��6��:�!j����V[�I�R��s������M�c&��sm�}���� 7�ut�vDg����|���}���d�Yt���w�h�E����'�"����)7N�h��o��El'<�uJA��ͫ���y�5�&7󴉓����I�-�Q2t[��U��->kvL��Z���D�r���v��Q���A���`=������M��[�5{�((nw��ܚT�-���v� ��d��J��aF�]*�@÷L�`-��i� �P_��j0U�Ɛ��aS�J���_���A��@'j}(yuE��u���z>�q=PK\�n ��UH"}%�9όƠ���ךx ���̺}*��� �P���Z�����8����i��%�)pCߣ�-�W�#F��LC�hc|��h�s/�m�B�^��1�p5ʊ��Ā��|K�v}[B� ���7F��ŋK�x��Od����
]�0�F��m7&��ڋ8��UP?V���K];L����R��Hf���=�����*�uS&�6�.M��E����HnZ�Y���۞�Ԟ���3 �L�[q�a3�|�\�q]�^�JI/�/�텇	^���>�	���Q�o����d�^������5�-�N߾}[V��h���>�o������{�-h-���+/�<y���s�	zJm��7ovM��f2d�nߺE��7��W_%Ϟ=gR�-d��?<T�B�A��P.��a�$ �{�缂���DϹ9��4j<�1쟋`��M���?:ܕ'OJ��{�%ׯ��RwU9���4��o�F8�.��]�O+	�t�c��}α�}��]��@أ7M(ff��������Ӣ�ta�3�c �l�������E����,���ޯc[4�Lq���[k�k��2�zf�;b^o?���t��������f��~P�[�1�e���ds���";v�����W�N�Z��-�;�_��[�z�s�o���~=�w��ŀ�>.�J-�����E�=Mx�sM�3(I�#f2F��������z��Pw�IL��G� ���e��J/l��'�*,, ���	lQ����j�������)
Hkw ���qh;\ش�pxk�Ji���Pn�d���|�I�����h�Y/�o"!��8H��8�x�@i�"xmt(��^��{\�ǚ)|��5�r��Wץ�Y:a�Ϗe<�o���}�Qda�����H�/��q��A?�Ƽ7m��q�vi.�#;}��A���b R�5�ĮLbE���-�
T�{���^x�\�u�Vf�Ix��5�d����f��I=*�}�mR����Ϭ��&|Pz#�_5<gf��b�,D����А���p�����\�k�Cs���f#��A.�U ��nnl�?Y�F2z�J&`�h|B�KϧF	�J� 2ߏ����Ki�hrbG����o��w��]0`^���a0 p-����cK���R��� .^<@y8T�wye�T��~�)��-���{��|��:��Kr����>�uW�7ᜠX��z���I�h3��wq�y��>/ <��@_�~�saM��3~���І��>)�&>>R�bD��l��D�ƜKR��B�?���,
l��fE:K��}��2��o"!��)�}��@w@=��`7��R���nɕ˫\�'#U,���c�
�I*��)���,%��L-�o��RE����6�R�>K/�-����~��׽���	k����xH��o�Q��xJ����c0�&Ԍp5���`�,6�w�h���0V&oY���)�S7N�q$����;{KI��gzA�G-I*녚>�?�ߏ�Ș���ӎ�5�>ZQu�g�#L!M�Z��z�5�/v�����LV������h�μ�Є��#��>ߡGQ���<�3��r|\xxJ� DSߠh���e�2��"v��DW�_���I�j�y#�մ<�c�n�;�bܒ�J�b3+�&1� ��z
���	�ѧRO��9��p_G�2<|#��{܈�wr�?�q&�Si/��@�K���6��u޲�-���K��$i ��L�;��.'��t�4�{���R��V���A"��f\8�T6]V�T_��bx��߻G�ȫɋ����%�Wj��A�*�2I�s7��H7�l4��p��f�r��:g��$�%�}�'�];�j�z������f����mc��$^�~-׮_'��IHY���UAGA���z��Hi%~C�Fw;�o�0_�}���_}�������	�8�Rꭚ�'��L�*b`~��I;�b��H����~��^��Ź�i����oՕ�"N�6Eф�I��1?m#�G��E9XV��"�訮7��8/t^��_�v ��`R$]+I!��妑��@s���sg���H1^x�ݎ���	��Aoe�+D�5�  ݑ���6��� j���NqQ޲��� �	���PR��;�6����9�;�n�i�3�`{�Fy+��n�r�kP��@x���ӢK���4��|�V]q��[�-oY��妺#�r૨Grߛ��̺�΋ ��Q��<�|z�̀޷��l�l6g�]�����6�Ϻ��t��f,�3d/�e���3�Y�eߠ�Y+Q�.��I��P���-��7T�<�i�TM|R�\�f/l`e �ْ���8�=�p4�DŃ��M�^]�ͨ����x`#a��I�%����2��֍��0  `	�r-1/a���P{+�"�*ݫ	�����+��z��a��q���%����h ���~���ݝ]f�cA;>���ڠ�+����ƕ��B��/� {�Ah++�{"�d�����n��'�;R�>_0\+w�m����ә�cp���8�����9{ 4�BOd� ������0kQx�1>frd�<���|���Kf8S�E�77��M��{�P�{g�6)��@)�=�qsJZ'��U����Y����N���YU7􎔮�^A�hCK�(� �hiYϘK0NA�<���5��-�54I^d5��P�>���ՅwF ���/�����cax ���{}�@;wۊ�T���пs,3���z'L����|�  �_��������c@4�^�|E�M��0���b�������U'�>�"�P�>>>$���?<���]��������_�#)T�?|��t��>�L n���q�뚖�������[V�r�9��_�w�/�,P�?�EH��h�V5AE��^G�4E/|���f�0ÒY)yիdt�c���E����7��֤+��mS�Ud�l�X&��f�C�ko�����u��/�����i����B��q���UO��it�҅����5�G�.��,k>�;;?S5���	�N�+c��x�a�<��\z��ķ���Ϸ��x8:e|:� Z_�L�}X�E
GN�N�l���F��a�� qqG�mB9h,����F�� r�uQ7�R)&u�E��[��gKP�K�X��`/@BN@���"l�+�9��V���*P��PFYM�U.��$��'����T�U���@��"�$���R����Fܱjm��߱��L��Sl��>�J����p���9 w_�l������0��g2�2���J'+����Ό+�VM�h�4�N��Ļ��{m4�t�,x��D��׍�ϒ5e�[,�hܷңsf��%�Xh�:��fM�����Z�={�r�H^ø���O?���;wo3)��RS��VD�Bm���aTx����`���*���$�L�W�*_�t�";�+쿯���{�Ƭ���<)Y�3Kê�ԍ�b�����9�N�J���'��ЄM�����������K�HJ)e��͑��� d��5�з�=�)�W0���Se�x8��[X[E�-/�\�����E�- ���_}%��� o�����@w<�?ƱF#(�
z-��!w�]a�G�s��7��667H���/(6>�/����'p�w�\���%R��k:m0�p:�$@/�k��@y���d�����zx�7�]��������5v�>�@GZ�A���*O�]��Ϥ�P��Ί��n�X�sM�v9��
��)'� O�<�(ߌe��R��O����si~es�%��[�������u/��|=J����H��XǼW�T�G��Z�٢�M�������d9M�o���䖐X7������p�_s����*���5�9�8�3'�K�c�i�]$9�3�ŗ9rk
Xt6�D���&���ט:xκ��3=��5�9��fqhxā���/�I�x��y��^�.C�!���Zxu)l8=Q璖v�
,����;X ����)�zPR��]A��2:�-"X��n쒻w7����i��U>�MOA&��Re�%d�vY(I8%�B�bѪ��6��W���y�jOv�d6�rR��o�C�p�p����(���(8ޮ ��8���ӥ�wQ9H3��W�s��A��iH�nL��^�t�I0��;-&�u��\����ih��UȢ���e�P�h�)��$T�{��)=�}􁬭�r�_[] gI����{�.I�#;��=��j_PX�h�	��4#�ht�����љ3�4G��M��� K��ʪ\cs��5���{FfHt�����ʈ��׮�]���t>b�<@�x<�"U�p� �Ϟ>#0����D���W�H�b�%�P���i�\w��kI`�[��i��o`�}a�|Qc�8��N���֫~ף�OS��h,5�� p�".�.ɢ�
h=����ѱ@?L�ޫn��#�?��͞�m�g�{��2�@uU�ܹ-��?�n��_��Mmb�	 ! ��.� �f0������+�!6�E'_��o�y�C*E�h(f����{����2q�>@'C��&R��B!�-~��s�B9�W��%�]��W��炁�1w��2ˈWެ6�i�9FA�����<��"�d���y��y�q�z������׈ݞ0�L��2�6�_��M����%�2(D�	
�|�������-_}�9�1�{���;��1	ȊƱ�tV ��W@U^���Ó��ĵ䠕��y?mPF�Ism���c�e�s�i�.��(��vtлZ�f5��!e\����8з�h��*���=4���x�RP�	���	�/9~���&�/x��b�>�`2v*J�z߼ym��~Hd�?��֗aL�U�=\u���O�^?OS�C!�Vl�+��9��x�b��o+�X]����mG�H�G	a_�\D�aE������ي�ؾ<2�ڿ=���]��-!\`<��c\�F`��ɖ�p�#�*.@�n�c9=^�8�tk��A��@[w<ۓ�F�X^>{���G���Gps�);z���	pA����9�[MȢ��j����TX��� �<C�H�n�*�t ���q�x��<�����o�&����6�}w��6�W�1��U��	eW�:s;�c����,ڏp9oZc�|��`��xŸEoq��`��2�7jY��H���2���i�E �����H_Z��f��ˑ���v�]̪Jm����'�u�&�>�����,zH��\�R�������V�|t�ƍ�"6N �o~C��Ʀv�-q-X!��U���b@T�;��� ��<���<�;��e�I�-3}g8���3���tg&���[�Toa���2n�gg�����&��1.��[r��]XE`{Hc}s�޽\��8�7����&��<h���(�|��y�
��1Ƶ��={m�Q������~������m��Y���<�Io��k��V��F�W_~-�#Fx���VrCl`c��^��'�ߍ �O~�1�5�\iB# =�c���f :3��J�h��  ��IDAT����[�[qݛ1�06�W-Z$����c�y=��Ձ��2�q��R�.zv��3��,$�hB[�}p7�����t>��-?י5��/;R<�j��O����!�1��ן}��/����V�[�4W#��>�`7�����"t���U���~a�B;xa����r�L�H�����_o�>��y��F�g7T�Y����H�B_/a�7Z���ťTQ'�c���_�N�����.<n��Ÿ�G
�`�ȵ�ErRp��}:y�K��X�Ǐ�c�}��g�����4���⻉�����6�.U�2���k���΀.��U�J��b�^�@ap\�����큚��¾A�B�md��H�h���Յ3����-���@)�\\���RF�4�����`�^��w���.����U����&��E\Pw�q��2Il�I\Q5��Y"�lb�@Ɋ���J^ ���)^h��C�/J�Vu���k$���:5 D�@-�����9���n��-���Q�>�����Oef8D�����Z�&.B#�0���n��Ő��r�XrJ���{�Z]J��1��?����\��UV&8l�i��d��b-�W��+��V���I�F �y/���s��'$�ƓFnXu�q.��T��@H��Q�.���SV��������9�� #I�8[�P�
��GsK�e���1C��,s��^�D[%�3�F�Ϲ"^M2�-���\m"/����0��{�� �a�d~����U�³b.�~��ƒq�d�D�T�? ������oӾ���O�|޼q�}�dԘVs<�$�r��߉��ccA�+
Hh��K��q�U�(B��;���}�բ����`o�P��t��M�RF�C��W���=-d�_��Rf�7���*�K/�D�H����r��=2��P�u�����k�քm�i\Sll,���/��@瞚-���n^忝�d!c-�a�`\���y�;�K)����~�2{�T��+��ߐ����f ���S(?���
d('�|\i���al�
.�o:���������\�	BjU ��Z����`I �ދe���	W�^�n���M�tlz^���
u������,�Qm�����]�O_�I��d>�xq}�A�y@|��:PTlX��¤���]�wZ��<�:0����N\���� (g�[�8_���1�I�1� o���ܷ���BȄI�[�Be�M��
�gi�}��V(��@�b_�.��-�R^���s]6�F��o:Ebg���bٰ�3����H�z���H�|[0�u\�jMTk�da10 ���I\,״0&�=i�A3o!Y�Į�����K�.�Q��T]�,�-�l��l�q3�LX�CQT�	*c3n��$���Q٬������<�^&�t:�j���l�JV��,�f7��I	G���y��|��G���k�@R[3��5�5��E$⤉��a�m��$-���@�#�?� N�W���p�0�����Q	��H�~:��ZN�M��l��	��21�W>�����{c�DpcAC>����C)�_��Lb{�衼��{Hl�?8���Z��	:�
6 ���ى|��o����EF,E9��g�w�\�dcYY�o�Xw�:W��fvǭ�!#�C㛫����j z�#%��D��X��F
�.b�Ѯ}��������'�ȓ'O������?b!�)cc��w��۷ͥ~n6�w�} ��O�$����1�(аi��L��bqMf(�@��xZZ�۵���(��q��Љ�銅��b��B�T|�懘ܽh<Cw��x�ƫ��]
m�Д���bsоy�:� ���0	\���B#v���p0�h�����r�P(\$F�S���ޞ��,	k�@�3�8���r���	�`�[?b����&x�jR,hF�G������8ƾ�Z�#p��G��zZs��Ǖ\��ׅ5���SW#Ȑ�z�rղ
&B]g�}�!uO40Aω�/�+`@3�E��t�7�?��6�����c�˰����'�|���Y�V5��\4,��wsM��&�K��G�ò���ca�USvPШ̾�ʒo�2�q"[T�qC=~0����`�X����pQ����D�ٕ���:+��B���j�x\:L�:�Y����� r�a<�����4 ���K�C�]a�y��;7l��7�vu5,��}dN)3'�nb u��`�d*���w٘5�d������DΏ��6�ߐ� .Hq�CYI��̢5��j�פ�E�����5ْ�z��d\ 2��vwE����"8�Q��CV/�jc+�D6Z�=����K^{�xA֡�x������Wq�[�)n�3��� �0�0���.�h��^�����rly�jD.7����C���I.>��Jm�$�.�Y`�4JF���6N%ƪx{QR�*��-��b0f��
k��_�|A�_��ܽsG�ܽ-׮�`�#W�]�ܔ3Lͨ���6�m9;�'������&�0Ǎ���q)qbk�O������"��f}k��t��� ��9�!?{��E'�T���cu�ca��5��,�- ���m��''�G���,|��!�2��B� ��S���B�/��P���,���X����@���C�y�@��6��[��D-��FV��,jC���8o����w2�b����T_�J����G�F��9T��,��8޴��3��:�kȠ����
���xĽ?��Bm�����J+{��3��f��d5��*ǲ3����R-#�s�W�e�5���PC�>5����p��ۑGp�`G泩z��l-�aI�JRo�BDT�r#����Zd<s Ua�[$B��à}~�XW��N��c^os�ֿ(�5��/ �+>�6���aS�P��R��UV�6��b
���V��-V|�i$��X]��Թ�^����s��S�1���&Y
�-K��C�֐�d�,'�4̡�
<�H��T=�Ǩ���:Uzm{�꒿x%ݺ��9k�L�jo����=_���}��I���C��1���q1 ��k����B�)JJ��X�D'�����z�c-��E��*nL��rt�TN^��9��4��`_�v)�ǧ��{ ���h�ߎ�s7,fq�d�������/��;��X�B�]7ܤ:Xex�x�d��{�֨��AV�4�j��Z<'�а��!n��{&�'�������$�zy��"��.�x��FPs�Ynx��Q�q�L����M(�F�m�;��p�7~�� ����Ti�ɵ��E3][냔״m$�Z=0����REv��X�������\F7Ng���KM�u���`%l�]�F�2���!��x�L����nݦ��D�f�\Z�ڙ3R	Mwnߑ��=��Jpio�$�ƁY�q����!�O�Z�j�g��S�+H�=D�Q�/��Sg|w����z`������3<���|ƪe���
��iL�&�"�U�NO�巿��J{O�����7����<�]���UI�ƞI�'{,d�����o�vV��PL�L~����{H����t��|�#�'G��O���d���q٬Q-�8��4�Pg����X�Y ���c[ $�x�,�%�0���ޙ�7IEa��57ޗ/_�a4�_���/�2� ��Y4�js��kX�d�J�M��ͣ|����#�I�(���zR����p{��zAn�;J4C�ށ��3� ��z�#�����h���i�q[�[99�R����C���.�N��,��ntn�s%������P��ˀ*%;�z�1�j\��AR�3��UV�14>��=���~���Q���E8��^#Z�K_=_`��(�d���s#�t#+�:H7&�<���ת�^�Om����/�|
��CH�Ե��TZi�eB�'Coz�����	��(11�UŞR���9�:���|�9{̰2���g{8�҆ңXǣ1�3��N��'On�������W�4�Y���q��g�����}����b� �w)8���9�6L�\Ԧ���K��8��Ϧ�"n0'��l|�[7��JkFX\5naZ�w�`W��(s0��u4ZE�[.�1��W�Ll&���gӠv���	dU�C001 6\��sY���R3�+���H�k��6�#��:ep���Q-T�v:��8�����f��'۫*�-T���Ӏ�W��Ux�:S��7�$ƆH'��h��cx#�ٛj�_H˱���@��D���SR��`�2�ݡ�y�h�Ou�T쏒�֤��VjBuKy,���}s��'?��<x灼�������ɯ�tu5��f�i_���,۬Ie�K�Y,�t��	/�	��]��V��z�r����Rm�(��E��\���]d���	����q�''d��ߨ����q@|*�x�ذo޼E6IY���/	\ ��ݵiQE_�Dk��q��M7��������?�W_~׎���t��b���Ԯ?B�c�(ON�����F���MIB5��Uj3*���*����X�������s���L���B�XA�D5�ѭ���>��g�XsܭV-�6֧1c����X>	������\�p{l)���0gU��؊�HOnK�l���L����PfL�?�J�:���ׁ�z���JhԯtDc�d#��;���]�oXmZ��ϣ�S��(A�I�_�DkKC������-��a[�ۆG.u�܃A�=ǘ٧j���㥿���o��h����M��Z�=jR2�AZގ��2	�N�~�&Tz�ru��6���(h����qZ�ŽM��j��cb��?��d$��MV�2�cm�|ؕ���ݺ6d�C�����w=6=���0�y�χ{�w�Dۙ����{^F�.�qU�p�,�����3:���
�(J����M��wT���s=�o���4;v:�X�����S؏������@ǅl7�#A	���a�̧;���Ԍgc���xrzD��cE+]AoKK6��?��%6I��Ѱ���[-�j\T�#&fa�Ԙ�7�5��ݥ�OhbD�[ `VX��[����������.�C�k<͉j�g�R ���vs��,����]�Ps�B����QI�D0�\]Z:�B-�챔�gK����0�uּ$���$ON�ڸ�(�f��|Ȟ����He֨�a�� "���U�2B�%�1QA�Ql ;�c��13��?d6<���匇mR��&�`R��'�U�H��6I��N�Y�o�lY��{�lAN�u���e6�t��ٛ��"1X �M���B�!lD]�U
?!3o�6�X�W!!�X�2>'y��� A�!�3d� X�޽'�؏/_�����ɷʵ�7�oݺ�ji�8�jj,�Ʀ�ub:,�8�|��Z�`]aB�uܨ�qĪNc2z3xz&���9=9���G���� �F�	/	+1 �B�q���gϟD@w(���|��',��7(3(��a�˳g/���~Ϳc�#9v��&���|glp~��ȳ�������Ǭ� �w���ۍG�����}��r���X^�h��7zT�,�ٍ��LAi�n�U{`���+a� A�ŭ[w��>��_ˉ���!ZI����2���~KVs�-_Cux��}\I�l��`�A�8 v�������.�	���^)���Fu�s���Pm^/(�P'�q2�b�Z)�!j��+ �=��j鄹�f�t �i^�gW�K��\��ǅ�]��u����9�@��\0�~s�0�5����K��1v���T��4���J�]Pp���`7%�e�滭Z��WE	�V�Q��鬤��}.sT],������n*�H<�M�{&��8�2B���00�FĢ�?n�{r��Rޏ��£WGq`4L��z��Q�����q�<Ƅ�mp��	��$�ݸ`��ą�L����8�q~,���&!^�	���MScX�-�Q4I����gX�N#�>�ׯ7l��A{���K�8���3��0FX�u��TI5�@?uV��dq���׸�M�n�>&�R��I�T��tc���ݱu��*��g�w]c�3ɯ!�gl5˼��p�@�<2)&�/�Mb�"1I8� �lnm�� �f��7'xB���w�1�"��G�Ѥ�!=��ꜭ[W�9��}�ܵ��x���B6kJcD�c��_1W��+��x�w�	]�O�;������l�y���Z��q�zxF��5&jPT���ʽ����I"¹�b����=y�Z��޸q�U�nߺ-�}����7�ˋ�t9��P_�O~���������;BT{[�Ĕ��d�T��Z	:�+xT�Q�0�1��}b��N��'��v&GG��� ������BP4D���P��0�����'��d6�;>^��M�~�Z+����ݹs��v�7�XU����^a�&�.YB��`��%����A/4���`}]o@`�cQ�w�2VkL��b�2�q�c�t<h��HU@�,�X]�J��p�ќ�.H���A���_΢����6��َy,�$���{�͵:1ʕ��`�h�\��2��6����%>']����z(�W�+Y�K+��7��UǛ�.;.c�q�	�HA�8Vq����䰬�{c�8�}$��w�6��} a�'ٗ<v6ɩ����{��nK2b&L�E�Zxr�>>gњ:�d��E��������*����Mk��K�xi�;i#U�\g1ɚ?c!��S?��F�d5%|�!>�y���m!����'�8OS��dk[�?��.�ý���Y0�}��A��ۍ͊p����;�'c��U���Rb ��B�L�ƻE�[�����;���"����A\qci&�Xl�H-֝�2y
�^�:hU�lF��r,� ��ɌNfKYǉ��}}v|H���|E�1|n�����>����p!�ad�k��ez���w�s��QX��1�hvԱ�f��Y��YK�n��P�rɸ-�3gnK�=w�se�ek�ߙ֏�v��,ߢ��Gx�q��d>��bR�ids�*71 o�����ڥ�}�j�^	n���P��U�2U�����{�R����U�!y�ߢ�oA��DQkFE�f�>�ø��x{L������,�X�}N�쮶�I���b�7-_��EO�$�	ֳk�T���F*�2c�J�{�K�x9���v}e���0�	V�ڵ�d�CC�����#Ρ�vQb%��{�=y��&#�ꆕ&16�i0�h��s��sH���s�P^͘��$@��c���&��M��6�*��(1G#^wF&���٩��Ӭٚ�Ό��u��x�e*k_���rM㳍zB*�c������;az�4}��A�e��6.�f�8���kaD�	@����ڔ��uL/�S���7+�xE���:>9����J�U���L��,���є�2tY�ݐ[����xOPyA�=	��hdY5�2���Cw�T4�U���Yǫ
Pc[�'�^y\�@�Z&�i��:�g~qU�����{�]���N,xRXr�;�L��B�A��ѓ�Go4�TYʱ�F6�Wl�E:�k�U��AN��^z ߛ��L�]!�eͱ�{[k`90oGU@p��㫫K`ôOߛR�Z�P����s�֕B�}y�:���fK�O���L�����&�5vd��Y��i6UE��Oe�|R~�k����i?��JkfB��Z�lP/����U���V9�B.y�? �R�u��:R0A�Xz�Q8�k7ߓ>��\^�<cц�|��颪Q<�tA�,.�ؖ9f��`�'��*F�#E��D㙞��(1*�u<>z!ǯ馠]32I�ƪ���U}Z׬��rȡ�ݽu�D׌U���|�&�ڈ�7���+�M@�Y�H�¦:�)oR�����=e�������7aC�S}�APUX�>&��[���g�d�mS�uAxF�b_|42�~�� ;~~�H�������tRBr %e_ K����&���4�������'*|�����<~Vl#k�9�/�iq�\�q��K��Y
S���U~Ց�}6N�wR��WA�	�8u�d8��ט\�n���'���=&�|�/2�+M��ڴ�p!��vHA���s�����O�bұ#� ��H�/ˇ�|+��}̲� Cw��ar!b�p��1�X��c��[SV��!;SVu�����۷nQ.��O+�Ŋ� �����9��Q�!�;������*)�rrrFm\�pgyNΊ���d��V
w�ľ��ʊ��=��W�Ѣ�H�'�UiD	#&z2Yn��%�qE�%
%����!훏r����+�� �X^�^~����y�P���>���@���g�~������v{��5��2��p����E���f@|6�������a��)qC;�e�P��ޓ����ap���� �F�ؒ��J��$������i�w�z�-�����A�S�Ot�rW�&sա�+���$�/���b�Uv/Ϙ��_�q�����	��N
U�s58V:O3O�$���2�'Sz� xk'ڐ�� �7d�H ��s��ܗ�޳���2���x�*H��0	&���'�zM�(�y�ClcX$�N^+AI&�"��#	�%��ߡ������\ m���-��U���Z����+� �y��ZC`9�zM+��[������t~O���F�/���h����XoN�� Qm�<��U�;7�Ohk��馦�4n���I��J�K���6$��q����E���鋳c��U���{��U������H`P�V��d7F$[���,�2&l��v�0�	A/�0ࡻی_Lk�z��t��Irk[g$�����i�3ح�pH�vȣ��VN׊N4�P�k���{�㬿9:��h�5V�#H������{��j�&��=MTx �h����t��Cn��3��1�~��vXf_���!!eB��T��ͳ�nTZT^L !����qv/m�%��?+5 �X�t��t��݉�}b��;�@��"L���@�`(u,θ邑UM�1�^��|{ߙ��?,K&���_��'O�q|=}����{A��8��?}��կ����	.�1��;xK�+��G�#�3j����5.�|ָF@?;��.֝�Oam@"#�ϒz�k�;0�&��R��e4,e�:�f���p~�kJ�\�i�Q���x�w�Zo��K�t���m��?~�9�'�'Z���`(1�#)��%sY��/׬���k���)	
��bF{���#�Z'A��v��țΤ!O��}zvF�dP�@. Cgq��j[�A��C�N)(A�>�k���=���]ˊk�.�����~�ch�l3b�{�.��I���QN�X��m-;<�~�d�k#
�5���1DDC��Y�2	�'.=*�6%�-E���5�
�4�v2i页�$��
̺�mr�P�4�z.�&���X�%D�xP�3� �~^U	H���*�''�,����>��__׻�<W]��OUA�y�qR����A���$Û���D�xّ��R74c^;W�rfa����5��IT��Y��Ds��WG0A��u��۲�J?'k
���K��@ņ�\�@x�����'b	[Y-� XG�r��S	�"n���w⠙K7����t�}�B�9��T�	��9KP�>k�M ���p�F�7�,�ɝ"���=.b��2 � �� ��8�	�%*`m�~�X��4
�&��7����`71�E_�qt)�ff��-����BB=r��� �-v������c���c����,`���_0���]H*�e��0��.6��ٙ��k�4�`����F�����(Ֆ�賧|ׅ滜p�,E�ܨ|��(Ÿ�f&}8i�_ҭ�/��[�	'ٻbQ��zNw�����7�P��� �����<l��2~v�X�Yd�����/��:Α�V@��4b|b�(D�������=�`���0Ȩ��Y WVw��f�7!1w�+��ۯ.�9 W��È�f�Y����0*3�<��y������c |40����7(m���x����Z%�)F��F"�|�����Z��:a�G�8]��,��Q���pS��<ā����_��J)�W�bw�7�7�<��o)�%��b�2N�/_ʋ���ڌɮ�y�L繫���+0@k��<����E�#^�"wt�*��"y�:���0�C�#�=U����v������T�h�G�o�o��R�����/H��7�ߢ�.�C>�o9 L)#?Ky�ڒ�ض�+blz���a��
�]�����qL���Z�0��!�aZ���iE���������U�0��\m�4SJv1W����gW6*m�&$�a�j�_�-)�*��@�Ə.�瑪�Uf���C��KM6�����O�:��:��L���n�A�3w��U�Ğ7�JL�������7N��D�B����mZY!ɂ��p 3�CR�֐�"� i_��A�հ& ��U��F�������ft�d<�ȲUU����&��� bk���f���9%����E5g��xY��J�����5{���[q>���@��T�㱜����^G��vʬ��x�F��0��VY� �$N�����c��R�W4Χ��d9-)�Bυr�II��ٺ$s$Tz�si�b���CM�"]ml���ëT�X"�aB7���h���@���2�?��O���	T�@o����{���G,�������;;��=��x�m,�	�<;cY�BX��&��L����>ҷ��m����̚�_^U.�O����������?�!�(�b�aw��x���#�d��G�;�ܗ���y��5iit���q�^қ��R#ID�7�T�� (O�`/������{��� �|���?�W�_(3�"����Q(7����J<�Hx�
�@F#�������Z���ގ�{}W=zL�D�̛�φBڨY��GPjl�������YR�J�a��������h��c�����D ۽h !aF^-E���Wm2��RHO���xJAZEC0�gg��׶V�S��ZY(K���B �R��I�������c�CJ`P�A���&��C������(�BZ�B�,_ӸC�p9P|��׳�
zk�_/���n咹�U!I�1�d�f?���G���󮴐Ȧ3);�L�0n_C�jXW��7 ���A��E6b2�/H����B�G+�V�(�6)xl4�� ���N��>�$���|}�0��iJF�=M��{�5\�-����U�Gr����r#.���	s�Z�Ѣ޳^�J���&�f�8�Y�`�2��1��\��R�;�$/n���q��1���*]�,��Sz#H�7�i��Ժ%#�-e�bc�ZrWP��l)�U��?�b]S1@�~�4[Wl10�%%�B��Os�nV�hs���|���(1:�(���J_ۍV�~������zM��n�UTL)*H�
J+��2��e�b�X��#hX�l�"�jQD0�gC�*����=���e����޻��Ƣ��k�3�R��}JǾ�֨nTcK�ТUc�MU��`��}��ܺ8�&Z��'�NLY�q�܉�$Y6�� 7
��x��F먥��T�\9{��pR��I[����u��,vn���Ϋ���5�nÅ�T��k�m����{�pmZ�z����6�`FmU�ժ$2��<l���c�Y��Pqt��l�
ߺyK>��c~���K2�`7��**�����|6�9��Z-��b�µf���l:b�&�}����pJ�b�Ó�ЪS�*P]lT$��FUEF�]�Xh5�TQ�4��-+���ٳi��9����"��E?tu�{0jR;�j���x�&{����81� {H�s0��K��<�/qT��X�>�'�/ �#�nC|=�� z]����s����̭�_�t-���o��� ϟ=�i��h#�OL�����M�0*a� �[�yp�7 7A�>����_��>��z�/�˒��%��p�w�� �um�Fy��}��{|.%�������O�A�J�5�����X/��.���E톾�Ӊ-�,�1p�	�.��A�}��Y�����SO���g�2k����7�c_��r����*�p�cmA>	��&3��_S����h�����Y(bm�Zs5R?UF5&V��#\A"�$_��*�J;�iE��>-�/����PKb��U򢤶��]o�qI�[̶#�',��w?��ǈ�lL��B�u�u�q��P� o����"k���9��n)pc�L���[(��� �ڨ�B�Z��*��C*�0~Wf����d}�a��W�E\��i��Y�HF�F�o��Q 0�"H9�.n^u �=��3�:N���q���]�s��n����d̍h>A(�ٻ�Bf/^��h���ٮ�m;K�k(t�'lh��Y�SV|�np� J�;{��޵4����Z��Ӛ! �I���OeK�b�V�Y��5�#��NH��R�A\�� C�s�l1�_<�JC�k��~6���w��=�M%�E���hg��Z�vJ��-��:&[����sV���b*��l,��6K$a\C2�,��N�
�|
���x���e�T��O=`9�{ͅ�*�Y�R��!Z��>ai��l�p1�����+������vy�δG\q�G��n�u���`]:�����,rg�;_2��v��B���|H8���/��e��?���F ��ٳ|Ub
W�A��)�$J�e'��� 	炋��� µ�f@���ܫ�WT�x7�������Ϟ>�gϟ�E���z!��ф�6n��s���9 {�s"� s�nw�P��G�=N�V������ӟ�T^�|�r�'l���%!�����W��n��1�st�M�򏎏ا0�0V� �Y0<�@p�6Q��� �e@�_��u�T��`���zL/@����-���=[��RGm_���?�1���|����|��soD�y����d��T&����L�dR`�d�J�[0@��N������y/ �A�˒����?�Tv~W���~gZ��j�l}�MǾ�ƭ��+���O^��Nϱ���g�g�K�4��x�d��(+k�7 �㶡�6��3x@�ձ�A
�,��၁��4��0�k]}�x6*KF�Y�J^���s$���4җ�h�K;���<��8>�,+�l���Ew"F��xqx<7�2F�,��|Kf�q-x{��0��02qV�oW
�+X"!"U
��_:�Ir�>v�)iܡ@���4f.BU�:
��0@����>�9�K2����ր$��9d"��9�� �k��
�Z�m���5�wU<H�j�zC�w�����������c�kT��5�6������������z�����P~r�>'�]/�"�:���L�x��ӓ�I�Ŀ-d@
E,��uiQz6L�|�bӝ]�ٻ)��^���S�0��d`0 �C-�F-Sl����p<8�K�vk���|g.��)�7��X�w2���F���c>���)�~SҺ�Jw���l ���|�|�ԕ��R��9�<
3h��[J;��ul��"`��~�6 �v�!��J���?�7o����%�\L(؅q�2�����	:�@|��G������T���UI�]�[�@XrE��->�tJ�Y"E8�L'�j0깬C�#�^W(C6��l��]��-~��߇� )���J�Z3�,~��]!C�터�
� ݓ'Ox����.��II�)V��y�ႈ��6��Y|vg��$"\k�5T�}U���$�Ύ�����D �g��-L�y��
���긶�A#n�z�f��_g;��b.� i �p�cS�`�� �:8؏c���T�A����i`���h3�d�[�=��;�&�$�~CŬ��m���(�)���ho��SV������]��K���_�v�J���6e?|\WŽh�>�	&ҚVY��3�C����iO�b׬�b�,Ʌ>@-c|���%�/c��~u�ͦ���,�$�9{�t�khx2���:��e0Y2�=9�������,yM̆��+�����yx�-��E��h�/t��ЎF7S(��t���'��+�ߛ���Ly?3���Im���I[l)gU�'��+3���qS�f���?�{
�1<ƵѤ��&���t�8����r`dԹ�4���Óu��Չ�5��y�4��w�%86�[gr���_�yݓ��ڼ5bds��Dʑ��?�!�(����a�'���.���/$���Y���󿊎� �jb�K7k��9�$uH�E����ӈ$���D��0�A
z���&ʤ4Z�q��(��]&����`�p�_�.� �E������JO|����k��M<�T��h'Z��<��s#�|:� ��ܺ���Cĝ����#��T�Ys��0��p��T�p���^y��g3�	���C6ƚ V3���]3P����w��*�u���F�?��ؤ�e7�^���
+��جռaҘ��h���5'"؆�G�rr�Z�>{�gN6���ʰ��-�efAc1����ط�t߼y��wc�7~��"WL�2>8'���q/���Syaeʤ��%�g��e��<lG�*��H��j�k+�Fډ�L��fnW��:7l�^R�#m;��3XY�M�"��؃���A_�)�\Y�X
\��E��}^�8�����_��Kka�c2)�������c�^ ^��H޽w�@H�M6dR�8��(��7i��`�<y�{���v��H�KQ"�`w4f�!��믾��x�۷�����;*-���x��&��u�q]g��-���T����%�ccx�m��5�����Ѹ�<�������u��7��;��2�M�u�ca]��J�!dR'�����������C��g1�9�����s�5�XKRBl�C#��ڄL�D1D�RZ��O�.�/ J��X�Y[Q7ޘ@j�[N2�;ֵ%��b�H7�),g�L̲���@�M��P�y2n8���y|��-��
�>`h����K��$���|߉sjOvP��QV�kT��Iy���/�:�KL���{���M��N�汈��w��7��U=]��GL�\S�_cĽv./�2,�A�"ժ؃S�'�Ǫ�n�H����ַK��]��[��F��`��ij�E^[첈i
������}�[�7��|�#��)*�e&6\�������6��'�%�ʅ#d˽�j_j�j���q1v�XqAd�^\��qvLf�`�*N���j� N�u8A��,�vt�J�^���=����lM�j�B9⸹�[y���\�&�n>��w#��U:b�띸Xܔ�j�����']ӭe��U�01���kmieռ�BE-ȉ��x�@fUq�Ow�$C[8.>��xG��P'k�oeVS�b����#j�uћ�S�*���LdD�<ɦV�%]$u�>�dA���^�\	*u3���6&�O��U�Ԛ';܂i[G�s��r���:��)u\0�2 ����ܓ?�0U'��Ȳ?yNlʈl=QL�$�-��E�z���y���h�mU��̫�V503a�6]{�d���7DUZ�l�ٺ��s����6�?�c�dP�9(0��F�����JgՂFԣ����T���+ޕ�M�]����&�V6k)�6C*"Vw�	�'J9{E�@
^#Q�#nu L�N �������2�ʔ��5S+�iH�˗3^�ޛ�1��e�VJ ��]��&�8h����4��,@�ϑ2�ʟϟ���|r�턶[� ��K���,�o��؊�-'i�Y	z��_n�p�lq��e�V��nn}1�=�Rv؃5.��bE��q�� �p`���'I��z���θ���x'�3㿬W>��\[;�%��u^�l���3�ɏ~�������gO���!����#A�h�8!Qtm�
�Z�T�)*& W�jƜ��5n��W2��ƈ]}�� �qh�P�c#XXjd�B�x��U�+�_;o��6c��9�Jcщ���\d�{{���� ^ʼ������"�a��+��Z�|�8�$L��W`���p�/�2���D.|��+U�s]��}��T'��o��|��-�V+��h�PR��7Ɵqp�"�99:�u�v(%YUq��[J�%��Q��nV2����x;�����H�=yI�"ȓ�s�	���l�uܰ_����{/"��V��k2�;�î���Ɂuz��S9=;�WG����Dp/T�D���|.��*M�c%�����$����l�f<3�A��w���I�}�Mܕ2��@��M�`-�:���ISve��evP@��N�϶�Q�=��	�tMa`d�i	��l�J�I�x�����G �5d��,�g	�{V��ۚtp~�ᆈ���?"cvpp�.m������6���rbZ��J��T�ʤ��a�9EǄǌ�W�W������M�;m�.䐆�!�'�>��0�s��D�ְ��k��\,4�J79�Ж�f��&������~}��d���8��΢�7��J�	�]�р��5�xg����!>�~5���&�)���s2�0@����7�I�� r�\n�Ƣ�9ϩ�!-�عƽ �jz��?��Ԯ�� �t[�����=����ʸNW+(���L���V��	��h��R��,����I� �_�6�!��;h���g���_�"��.+�90�X]7�|���^��l$�p�W�8α^Uuksk��59ؿ&�n�漃a	��`�%�`!UQz]dh�xH
�r]�����g��'�,wYeF�_����L��n����\�ߋ��Z�F-��[�^C���:~��K&�XuV�tfH���\E�Ao�`V)����Q����=iGU6�+\��
:n4�c F�ɼo�h�����[_n����4D`�X%p�|���%q���uk?E�ͳt���ŏ$M���4�3�h�~�����_�~x�BW��-���o��/*9�!uO0�~��ws�&k�[���K��8��j֮�U[ot�w�5���|�BkV��֐����lI@��C�_?�ӓu|��X1�ՃJk` �eI����Ͽ����}_� � p�pXe�޸s_6ݙ� o���#�FQ�i�lgu�V���ɝ%���-N��:�_���,~�\e�%I�d���Ƿ-�U�K�4�:aKϖ�_���w貣�Js���1��N8�ۙ۽�����M���f]�5ީ�kg���|ϟ���-�Fa.J������������/~I7<6�QxY{���.t����ژr���W���T7Y��������<6��2��o�5�r�%�i]��W��sa[`
�ۚve%U��b�p X��f��.�������Ȯ��b;��>�C�e�{�Sġ��x��
p��M��"���ף��j ��nS\����Q���Y[ y)�����:(�4Yr<Ob�v[Ɩf�M�ZJV��O�(����?7N�@�ecrx�1���6�9<��џ��#�!W�+�*�~�Rwk��keyOÿocj[S%poT��xo�d�������U�9J�`"�v�M1GǠJw�@�x������!w��� ���_Qc�DC��z�ZR�뚴���%��C?���1��G�T��[$I�Zq�?%X��P���/��B=�R�x_ȽA1��fIՖ�k�2�u#��L^^-�e�
rv�G�  F�+(�W+�b�l{��b����ђ-�/u
d=�r�c%�;c�MS������1����n)�&�W���!�d�9�֪�3c�"t��j	�J&Xz}Y�\��q��ժb�&T1���j��U�D��
����2����ǥ+�a�O�Y=��1����<�B`R⥾{4o�y���^<UDe�̪���6�$AB�����H���5�L�o.7���-G�:C��:q�Ir'n�qR��<'�.9Y�"������|�h#w߹%7op��}.@#lr��܊w����(�z�$���h4�+�J��&t{�
�%��p�ϱ�+R+ͤ"���"�3��������4�҂*;gkW�k�����œ�~-���:���P9�PI�[�c�X���tZ�P��S�2�61j$,��Ve��RA���s#6j�>���#�����<{��n�_��d�4)�]�Wl�l7<�e�(d�R���/7;UOh�.[�v*�ǐ�5S�U��̀��*>u�hU�jOH�1W��v��JL��-���,�]TPCh ʔ����uukk��إ.�����	i-P�皴2�.��#�E�Sp��Y2��G��;ppC��4�uNy9]�ُ]�xQ��U�L�B�������!����d��aխ�˺�����@mɆ�?�C�]���s��ݛ��cxo���q"P������o�fy��_��{��e�38�����C��{��%f��o����?CC!�7��ާ̞�l�������~(���_����k7y.$oC���a@���]J�!9F�I�UV��UF�^����D�kC[�<'�	�XHZ6*_��D��u��x_��+#��;�L�.��4�z݋sux�j&/������#�u���GP¥"1��H�]$�|O�}������x�'c �^�?�ޓ*a�����jM��Tm������b�*�3�ԓ�No$J�]>�p=K����Iq�JV!t�L/����l8*1ѥ�ـ�dh��*)��oYO�o=��doNZ�72l�ˏ��W��}C̕@���`,�µ�UC%qY5-�Y-8�ɔE˯[��o��L֋���ǲ8�dU�滲{m$F�wpC�?{*O�>���esr�Q��(��e�УoF�<��]�ؕ��0�V������i�/�~�*�K�Xcl�j `Ю�J	�� )�����h��[�e4��7j�!O'2�V�8�&30�#�lT¶�X��r�W��ew�q^o�n�ġ7$���~��ä2Fέ~?������sfwk�xZ�JS�х�S�xPRU�W�Ƕ��5����n�����jI[�����E�ӟ�.vWߛ6lg��Fi�j�Y�J����gbr|A����$��"�V���
i��*��n}�\�.��N��a�X`F\x�*�+Ƈ$��'��$���Z��%5n�HgfIu07L� ��u����eV�Y���Чr�̱�j�偹-�$��L��ƩZ�Y�?�z����g}��ӲΞ������6?�L<5�*�&�^����CpW~��}�Jp�sQ3C�t��������<�h�J��Ψ��d2g,�c�|�{���m��ai(dF�"3><.7�m]���::~.w�����N
�����0�ۜaV��C�e���o�����?���D�os��b�����O�u�B"��C�<��������O>�	e�`��<� �+���CV�s]W�5;;S�{熼>��ngN� $Ւ��-�7�t6�#4HU[�E�U���v�񕘱��%p���z�g3�M@�rwW泑����ys/���:��}�ɬ�'��>�z�Z=�D���x4Ṫ�J<��aUb�,ט���F[o/�E}L����$�,ϦJ����)��%�Ly}�<�Rϒ%8W^u4���ͤ�=�M��8��8(�,[��R��P�:�+z���>�kKV�|�*vum�3�^Y2���u��}-xXC	rK \��L��Qe"��G)�,g�!���}Z�y3�-O�"��V��{���L"V�0�Vq\���
�q2̘^sc�À�f�1N1�as-��趶�5��SU���E �{���pkn�D0�d~����5+7��*��I�6���n�&�%�=�͗q�/��t�$V+ł�*���.7'|�)/]����I��ԥ?���!C=���M}��fZ��+���!���jp6Nh&�����o&��
@������8��:�n&�e�o��F`��&NMB�d
��f; ����h���^d��<#6�ѣoe�檥���6K!%�����r9X����d/�vvw�|q�7���4��S�5O5L�A]g+�Q�e��� �jH?��һt�>�=qA5�\��Ҋ�ŝ���`T*a8�v�ѥ�K��C[�U������bQ)6����rp��{H�4ߓ������G������(�*x�ظ�z�+AYy�۾[n@C@�c�߻����~vv���1�os���!�~g�Fos�����gO���m���%C_^w������'�|"���C��o��o�	@�ڵ~8�W5��b¨���U�. >PH������k{�����o~���g�@F��˄�Ϙ�8_gs(�Z��J��= ���F-B�@$ >�VCM���k��=fE��B :2�;��'�wmz�P'Bx�!;6�8c�8=>����I�~���	%*2�hsc���Z�3��OY툀]�ʽlt���r��0erT�o��w��J��VF��{�:_2�)0P�1��z+���`��m#2B����:z�2�#�Q*)Ă������Q�d4J*"y��Uubq��CAMb:�Y4Bv���֐�*%��-/Pٛ<�\��Su�I�!�_�G���/l�)c��M��#[-|��)ڢ�h@=j�t���,���h�<c��;�C�/ݑҏVG�� U�PxEA{�`�q=�]��S�Q'���M �zk~Gn߻-w�_���WT~X���2���i��G`l����M��q����L6gp���_۩4���,6�]j�O\LV ��cY�xOeݞ3fw���ga�R?�;��`z��kB�%����~o����  ]֣��ps������ĘO�#옳���E>\�,!�CJ9��1@�<�\]�4J��Y��e]��d� ��~򓟐9�����?gV��qd�(�z�op���xݍ�6 Y���kr�&��rx�<�;*O����!��M�.�&H68��� �<7<ϵ�G���Fj{\b��91�7�bLU��[��-�U){�ɔ+���a<^ӕJx1�Y$�]�*�(<!��1=G�f|�鶾�"�ȅ�Ǉ�ֻ� HU	a�絵��(��
U6
���!{x��6`m���/۾��G�����@�3�CFx���~��+�s���6 ?|�4������r<_�� �{�'�*���sC,|̔��7�(��駟��	�o����z �8?��"�tI��C��c��h�Jy��f0;��_��>X����_}!���+�����\�pH/Pzo_Ϗ} {��)��ʅ�
jܟW�s����6�!�o�!�lA߃w# ��w"'�h����V�Ը�//�prvF/ދ�/��,%��)�5�BX3��~��+3�fg��j��F�l���$�.����4(I�rP$�8ߏ�s�����zo���w�L��}k�p���P��,��	�	'�\��ng��@@Oo8o\�I��\�`�Eұm���r����Mttïo���5�����*�>�D�^(�P�tz Tڸ��B�Z;�6��P)�3Z���]�H.�J�WƆ��$��A��D:�t�4�����*N�6�C�(�U4�N�n
��@�H3�Y�"�Ƴ}ُ�x:��ȵ��e�E*V�d2�d�w�����t��F%�B)�Yh���=��#VWY���Z�n�Y�P�|�0>w�����Р:_�U*3�'qv�[H�Cb�\���0`?��Y0E=��&U:鿟7��g�:��4�٦<���]VyB��tɦ�����+��Ĵ��q��	ȱ�n�޾sW޹�@���-+p�>x�.�a��_��[f԰h��s�hw��}�ɚ�]p���h�u��0����	�4b5\��±�ms~���׊��C5��	��ޗ�<������u�d���2ל2�y���H�kQ�M�:��D5S�W5�A+�;�$�kAOV�R翵�����QY5Nۢ.؈�ԒC|.?BU���p�"�y[A��s���s��6P�-b���]��R���b��1�۞�|�mZ�Wo��^�]_��\��9�|�}��/� u���{�w����(�`�� �������bA!Gy��{ʬ�������������r���C�qU�4�ⷿ��@�o��ʵk3��O>fx*�j���ڪ�,��5Uj6b+��V���k���~{Q�� �:-�rpmO�y�^|����o���/������P_h���R
!}�ř�d�:��>�d��)�z������a\����r�q2����ؚ,0ԉ�J)Y�-!���/�dG_l�>���l�u�}��J�\�8w�j�E>$�_��>����J� `�+`x��7��u�e�s��p.k-\���CkX␃hL�8v���K������?-����3��	�(m�ŧ��˕��]��Ð�������`78��R��Tn2�B�
�C����5'�2��#`õ�9� D�3��5!W�����4v�L�	ͼx�������f�ఒ�׏�� 6^�d���挲gRC���6�������xǯd����Z�^$�Ў��6��v�4���/��i��*�������
�[����=�*����FK<l��C�]�n(Qe�Y$�^��y*j`�NHf�� ڽ�G�9��E44�1E[@貳d&ev}vK*����JD���|��O�"����'�c��.k��%����6R_���Ul���}u��b����-�.��O+��\ڀ6#�r�Q���Υ�F�����x5i������{7ե��$�k������3�;����"�M�cq��od>�aE�������Jf�U\%�(��@ȃxxغ"�!(�(|�ׯ;�p�r��M��xW�5
�;�	��֒����.�>H���}?��u�k�_�Me�k��,9�M�g�K��JW<�����.�ۂ�2�끖��������\���&�a�[P\��Q	rg��B)?��"�o��cy�;wn���˗/�n��C���uZtc�eiUBp��Œ���@8:~-��k�}�:����ܸ�+��F����1u]�#3&�wN����`{�~������Lצ.���b,�1�$D����Y|�;��'*��n\�w(7����Z|�:��#��r�'\����#�ݗ����,"�=���&�x��Q*i Θ����YJR�Pt�mU�͋S��`p�[�g���tpd���2���p�zc�)��N�v�������~�*���S�mI��8��lu����kk��b~3!��/q�{c��]�ȂJ���C0*q̠�䲂Z=ZǱ����g����F4 [m������<�-�h�F-���p���E�e]�x�"0B(ܡ�$���4F�Cb�mC�L��K�(�4 kY�K9=?��+�&P�p�Ak%�թ���r��@wq,��#YWH�9��z�H}9��$�ܑU��c֟���~�#��H�e��+���e��~�Xy߭��i�W��Qr�*�����r��y��6\TC���X%h:�f��.[[�[��8 ����c��������t4�����S��>���j�:孤temy~6��ْU�۶I3ak��3Ӻ@j҂��u��ܟ�y@R� �c��:�H�R����Ua�������dB]���K9��b���.���F�T��l.��P�n���>��Fȟ�ٟ���.ݠ���/��������'�J�&��(+�����Z�{��$~~�VVV�F���Y�4G
���a�6���,�Hua��کhCv["�6`V���ۘ�Y���c��(w���
wvs�0L�+�?���~�YC���?�
_v���po�]�<��Rq�N�;,e}��C5!P7�Z��|��F�y�����q��˿�s��1ؿ��1u�KC��cD�g�7�4KO�N���g��_�6�k���"�<�w����k,����K9>>!�uo����^�����}�m΃��w�jV@�dx}�J��j��/>�^ל�����v������\a��L��ʄ��Z{���f@ @��������Lf��V:���I�0��A#��ޯ��^m��b��J,"����)���Q�Ҏ/��f|� ��HfX���?�r���4~���Z�-]/-{zN�9��~x��\3̣jX��o�E�-����c����0�w9B(H���e�'\����,��ef�yc��r��W* \��T6H�J
�0�M|��5��Z�f��.>f���8���F��4�&�0>�Z��*!4��T7Z�5�"�u��U\�Pw��&�A�- �i|/Z����O¨� Q�6n��1csG4P"O5Am:�xU�AL{yH��A�-�oH�*�u�ϥ<����6#��ǐ�X���gЉ��nfq�c!�_ ��U�W�&���"�b'��!�ͷ���|��+cW�2T�~���Ï��"	y�媍�L>�ླྀ���d��*M�T���\4�?*��3�V��y���mRJ(�u����m�̼���W8��9]xܿU�z�������`�]\�]��e:9*8k��X����O�(��؃w��_��O������D�H�<z�M܈_ō�������}�k@F!/`����`�ݓ��KmSq����1�X���߻�o*��^%<�T����םB
��rIU�g���Vɚ:�t Z2�޷�����c�ݕ����W�]�ku��!	C��V�ʥy�\ZU�˙�����n	x�������B!���2�yh8����vC���=-�c�څL��A|�_�~�����������kr��-���x���R
~��E�Oh�~My0��01^<\H�]��A�\+�<�{[,�L����/������ʻ�#�ĹIv7����q�Dq�M���r�T� ]('Iw���M?J-k��b�d�w$���/
�T����TPd
�$֛e4\��8�\PyPO�E(��Ξ�$?�)��^�I�����;��O!�9���v+��!�f�	 &��"ε
i�u�!y^C!���#	L�j����O^��L�G�X��Ee������9�*m.��}(�����ﾥ��}��(�a��-c�����L�+��p���TJy�oo;gI��4GWb~ýx��E6�7[��
8��/�[l�ۮ�w�_,fqB�͕�����ڎ�q�VbH�~��%�ް�D+����vE�1��`Q@�/H�@�Cy`����w\PF�YL�0\�4CQ5r�i�\�!N�*�詺w��;Q���\k��r�,ؑM��?�5��37do���:^]'XC���D����\Fb���b��M���ed�g���B(��JBS�4���ݞǓ��A�
��7�&u�k���;��P���J��歛�iŢy10�X�=��V|�������j�Et��Ԙ�?��O	�>|H ������e٬KZ'�$�m]k��%3Ĵ�T�e��*͗~���d��$6�*�_��%���f�}�% ���ƞ@}�N:�>tm��F��7'�m4��Frc�/4|� T��;����z�u���&���q����΄�cKa�[Ѱٓ��q��G�YZ��>�a��U9p/k�,�/�3���s3n������PV6�A2 	�5 �yw���#/���Δ0�c�Ѥ�7n��+*����h:0U��8���{ϒ�S	&}�u��+cj�>/�VA��� �����X�� �H*B6���(��Ϗ��l��p�aXŶ��m��	z��2|�۵L���,e�p\��{��Ӝ��x��A4��y�������!?��r��=2���p���@A��͛���s�����<q(��}D�E(8<}��c�/J�C6P�B蜁~6 XTbݲҙ���q�0����#�����'�E*�6E���B� �=h8�$΅1����sZ��E�@}b55+�Bo�je�<zP�����e��9�,���<:���9�xo�7��Ym �8��JO�ǹ<��q�{ �q��b?�1<��͈{��ݚ׬L�V�F���̄C���xغ��;�1I:gm��R����U���_��j�5֋k��Y�� SoV<�1��%V �P�^��U�M����n�%HQ�*�."�o0������}�r��!!�p��DM����M{~�׻�����b2(��=u�v��/"�[4E�1�����KA/	�*V�h ��iY�!L���V���1C$�����bE0��s�l�O��j,��\���m\<C� r#-�ʸ]lr�1�׈ x�����-ʻ���du{�>+;����$�x������-nƊ�=�	c��XZ�j1~�@V@�O�U@"��W:.�+�h��x��u��f�iu6��	��� ���;M/k���7$��ot`�2�'c4��QY<s���c�Fs�Ɵ&�$T�,��[��������WB���9郧@��F,�p�w���J+��A;c9S���ܺ͘<݀�������ɷ2��H^���~:9~E���[r-����7��Y�qx��)� c3�	z���m��1�
tr9W�����.Y���JAM�'�����&y���3e���mj�p T��]�oC��koׁU��MoL8��"����)>{ �X�sz"�G(��0&����X�����Ψ�*���g����J��I����h�E@�7'󉐫M���ơ�GZ�h6�2�&����"�(�R�6��5�_C�&�|fB	)Hx<N�t�z����U k���ZV=�U��bY��ڋ�t�/Jr��5�'n��1�q��sJ<^����#I�s�Yh�3����CJ��D���;G�����۟�i)Q�n8޵C��Q6c�&�fVV�顨�>� �*3#���~ם���v���<?8��hs.3#��,٧WR����T��쐸�>�AyEd��?~.������6 W$�!3������#�9(sk^D�~(g�i�ݨ���g -�e�T�����)3͋8����&�]��w':���=`��	���|��L�\���u#�x4��U����N�'2,Ο�#k!�q�+���D5#�2L �U�`���6{l� =�Z�Kv����Ƃ@����Uê�0�(�ۓ�Y�R $e o̾�I�]B5=l
 �����+U�Dk`�ipل��i]g��GKI��^����Αk��F3�rD����Z7ʀ>�AUH���Ţ�5��������+��Z�0/ns-61�<���ϧ����F��uzz����ֲI��^��;m3�Q����MN��<��]�_U���!�PX��g�~�kX6�R��:�n�Ul���'-���!?����/�%�Sl
~����^cH�._{�Uz5����=���9�-|��GI�=es���v/Y_҃�^�����OBpD�����^}�����T�a��ؽ`.$@WH��k�����b��I� �j,�{�1c�&<x�"�cT��3cR=h5� -��@��\Z[p�m��c�m��Ԓ�O�i,n�7���U�� ��g���u�3D���:��j�Af>����]>���W�
��U��}��:k�t�{�\��N�ǈ�W���씉(_V���@��>�5�4��E�������E�� ���5�q�&�o�̂^�ڕ�gJ�?�� Y�HK���&v�Z���+��[��=?�ؽa4�r�����IG�(�<;�"A��`BTմ��ɀVܐe�@[�/[Qa!Z[�'��9>!!)4-3�hmO�Ɋ���,謀�<���?�F�����Q��pˮ���}�h��E*f���7kսa�d�/�+�z�uⒶȰ.����3sf�}��M��T0KuWM,1����^���+��4�X0oBz/�(6o^���{�&���&$���HՒ�!H@d�%�(� �PAn	��h��XW^����K����o�3�%`��lWZ�V7J��x���H^KCf�14���yƁ7�a^��cS^�Y�IRQ��g@^ ��#�<]��a/y���*2�>�͋��9%�z"�� i�I��������+w������){&���4pb��xMYЌ���}���/�믿a������K֎+(6-���4��x�a&۬m����R,�V!���CH�=��E�iuB����w���.�k�fr�+ �ĵ��`�ƣ3:;E0�s3CP�?ٗr�iLF��N�,)#����ۇliAc\ x�9y��X��X��2�¤�c�J/L�V��|�=�iH������s�z�,�8���a���c��� 6���%\����/9W���>���K�M��E�X[{F�޵ ���׀z[���6b�ϳ�����<<�X<�a���»1�:������2�����&�ӧO����I���Ν[��wc��z��u�f&C`a�*�Q�|�9}��g\I+�iZ;�=�'O�����^|a��!���Ġ'lmE�tco#Ϳ9=y����O9�
�Ys�}�8wm�J'��d���5^�	l���Ql��� 5�b���xJ'�;L<@�^}rtF��أ������.Otso�S�m��ei��Y���\�i.i� ��/����Y��by»j� bdZ����W��g����ۅ�?F%��=�C��%�*����⯗]9��~������y(ë �uL\4��Lj����0Л�-d$h��Z�u?��T����**��۔2�U�zd_����E9c��W���S�7hZ")��
�.J�eEu�s�|��z��r��`9����`���� �4/a�
�m�E�a�����5�w"Irmw7��@�1�Q��_UQ�`��L�/ٜ5��P���O?���+JJnmoq���v�$��x�&�If�%�����(l���������S �2��_@������	�����%{Q�$�Z�e�k}+�zɃ�*HVD[�����ήv�֎�j��ōaʁb7o�3%��b�kx
i�N�8��!X�i'���u����1���c�+�$���_���qONϘ�B^e�L�?ժ�I~\��0}�D
��p�����ګ��8��;u�ԵK��j���5�Aۼo���֖�G)+:�O���aײR�޵�>�mر�ہhy\]�>� 9���~^t~_�U�޶2�Ϊq����G��z���9�����+�飏hwo���"`����6�탼����_}C���o�_~�oim<gY�93f?��35�Y�F�U^���٠��Az�1��z �"��\�j^]�_�7����h����K�a�L���DH%J$���l\Kk�;Q��@a><8�ԑI��]��a��"&����8�28 �������0k�ӳ5:^G�z\oȹ漢�Uk�d��ƴ���eV��D<����	��lj��J�_�/�C�F�[�=]`�5�
��o]M<�cEZ2c��uI��b�H#�L�����T0��o}!h�R�
Zl�d��w�I2jY�}�㩧,�c�DTZn�:�[�}���y�thr������̤���m1�9(���"�q�ڍ� k�	������xԼp�@3ë��F5k'���^8p�ƙ�I768��N �����U�c(��;�Ҿ,�k	"�*��tU�
{<WA�����\K�ӏ*�\�?d�/>���� çNn`������J�6Ȕ�xbG�4jIܦ�*�s� ��.�r١��G�ۋ}BS?��c~.T���7������OO�\+u�+f�q�zR2��:+.�?a�

���#�`���޸y�vvw�G�;t||B��z҂)�t|��Ҋ�VЛb^�iҟffԧ�2�g>�91:���_I 9�L+���,/X	`�y�gT��|�����3(�B���R��O�c>3����������N{�j�F�<ų�c��m��[�����=�l��U�tӧŌ�g���+p���ϑ�\;xM�x�L=
-���LS���-�ʃT������b����W_���gh8<<rL{?j�
[�(I[���K�6y&T#��>���d����X��o�����-��o�u�b��"����&�<ܺs/5w m�8 ��*����~�b�`b�&\�8�t.�l\B~&����(e�cIG�@0�5��ht���8�����G�6���	��ӗ_~�A��{�ӳ����IR�w�:&�N;{[�l��7F���r[��p��,Qޏ��k�0�g�4P�j���X��"�K{�Y�<L�+���1d v����/�ْ��m dX�,/_0�j�r�8�"��� eSF7�L4ԏؾHCC��?S��|W���w6:D�[��Ӿ�,�EP�I�7WR	0j��clɮg�h���yi^��	 �B��}[�p��c�vl�ݫL;�ۜ������<��)�/W�̆0||c�5���Y�l�Z��RpB�����6D
�2�Ȯ
��Yi�TQ��GKW�3���[>oe΂D$K�/��m
>y& �^��ok�n��.p*wb���8pT���܆i���	.����������o��?b1o�3cЄtIb����z�li:��u�ݺy��r��z�fc1`� ��V�����	H��%
��b�(D"Lz��g��T��RI˞ó��w��j��{������M��y��y8Z�>��
7���{A��8,�������p��a��,�0��;�9u۬pWα����yc�]"]_/cb�z��s�k�߳v]�n��e��/S�0?�/������7�<��I�{����h¹p�<~���SP�$��[d��Տ��+'i� j�����`���/���g�t�}�����) �1�;�� 7W�+ng}�X3g�Kժ��%�/��`��l��x������� ����9���h|1�a/�1k�=��)����W�G����N@9�Bԛ_��<)��Z�e��%�+���e�m"&�ĝѬ�~��\S,�{��������C�$M�x�w;ɭ����[�+�^��qm�
'](�6����eW��V\|/6���e@��B�Vs�/��9�@�� ���H�ŧk�P^�Q˖*7�.����n*�1��X��0�{�IelT�9��d���>�+���9dC~�����+(��gᶙ	_,LB���v�tR��=W$�w����3�������������_��(����z���5���Ώ��eɩ�++�$}0;�o0k���J;�t8;�I>���R�<�vP��gN��ls�=��-���Yux��#�`�lg
�u�Ms�2f�C�)�>z�n���+�1�n��d-�<��|�R���uMx���ҥ5��#I�{&�y��!GU�J�^v� ���}�?���V�7hc}���a������w���~�����=y��>��SN�tv~�`��b�*�M�}�y<����{l%1˛��Y���m~#^�������`L�6xl���oL�?�Ky1��c��Ƹ���z�]|���������}�<P7F�γ�� �Rv�M�0�����2�k����R0��2��&l+ ���� �vo�b�?��9�ezO�4�qh>y�O��[cn$�{x��9_{#|�gZ�R�[��������X�BH�>d.���m���ލ�����O���0����=?<��x�9�H9��\��M��`�¾g.: �l�L�`������'V_%%ԛ�g<�ކ ��$�G��A` uϛ�kLf`�gt��?����3�%�{�t�h4@���6�i��יh�Z)��h�(�b.�)i�4��"�L��ؚ\l��X0��%�$����D� �+��[ :��u���׶6�Yai*���_T/*�c�g�
~�Y����'
�7�3W�}�hg��6��Kl7�.��V��-�]M�E�ꌁf)Xh�<SAx����vv����1����eQ|�uYF���-�������<+�q�g�ȪЩ�h��Sɕ�N�b殐_��CU�rm��6`�MG{F���y��\�趵�+���v�rf 1� ��}˽[5�O�TR�5��Y�� }n3�G���1�~/]�'2I�����̧��VT d�@�	��܂�����k��oҽ������S�%ez{g��ܻ�B����=~L�GJ�����O���ӆ����Q����7��m��쳕c�)��}�ߣ�7P�]���6��=��_؃�vp�/&�-oUw��.��v}���L]���AQ�]v�b���Ϫ9�~���=�%e�*���_���Gz�w���>?d�+�i�+ֶ�ظ��6Iv���:�k�!g:O��a��A����#�M���NR@o�Fz�]��ץ�%gXH����)[ep �U�������끦��i��Y�5/q9�F�[Α��w�ݭu���E���J��R��~_d�8���B2������z�&��Fa��`@�H� �%��dL"���*�#��W��
��6�a���2�����Ul�h]n�t2�A�$H>}L�{a�*��е�]�ܕ��-��Qx�ܦL� �&��R�7��\����R�Y�im
������j��Ƙv�6�c��D����_�$�wkˑ��@���h׎1��1Z��`��ȋ�E�E�Z�V�d�Jd�dn1�
K@�J�ٹ<\l��ж�ź 1KW�$X�_X����w�aV��1�/��^X����h5#NKU˼ �ثK1���|���`G�M�Z��ht�)(��F�5�).���	k>�d��,�a���/?+���NF4��W=N���tr7�^V����tf��|BI�f}s3�Հ�1��iwo�}�������t�?�6A�"p�B{���IMI�
�t�;�ٲ�{��*,�'���z���6�g��l���|�v�
����sH����y^U�Ҏ�,�۾�d(�V��?��m߾f�=�)O�sp�yS䯹X����o�o���t��}�O೻��S�1�8ה��䛵��N�q�5g�e���_��B��LXS���gH���#�9�G�z�~:g�+���c8`��`�T�"E
�R-9gy���E'�W?����(��⇌@56��QRg�h��l'�y��޺A{7wh{s��Kf��	��]LD��p��{����k���(��!}�}F��[Y�\\�8��䈕��f�.8�B4F����/v�谯n�Y/�׎<"#���˗lᓎ5�r>�N�h����g��Π�
7�l�k{�P37��b8��lEÑ�4�r�l���nh�k�ߠ��k����]v��V�P(kb�󚗈y�4�x�PF�ߪ��d�8��7����͒fv��'��Q�S\D���W�o �ٷ���2)����җ��TYy�&e׼4��~w����h�[J˚2Ľ`^7��l�C��V�^�>��W~�x�

RUHSI]VS�\s"y�ͨ+�r����M���L������1�,$=��N�>|=R`��p��C:=�'DP3�� ���+;{7���@�N&�HgLHI���3JhY��cI�d��8S���Ŷ^�h�[3Ś�Ϊ�s��rxS��2��.�����x]!8�;̴]&�*#^��vM�n��w��8�
�W��j) ��Ɔ�P>9>� �ãc�Sz����j˵��
��,8��3͜PY�I�����%�~��===�'O�ҭ���%�btN����Gttr��ېN�Ƽ����S���'#��s���:# [0 ̙�Ѥ~�Z�E�^����-��1���+n?J�_�����1gf��f-y��
�~��	��߾)�Ư>x@����g	L��7\〻��9����wB��6��	be�o�sr��ղ-�W��'!��)vJ���Wt�k�j�+7��X���bы��k��;܁^���֪���+3���(��x?,L�����ߒ�JĲL�.E���l]'��=��۲?O`;G���"�I�'��~c����lL��;6��-��G{�Uc�곗&k���B"���V�jƪ(M�b3P����C�>Ǖj�����u�9���Y�_�w���6��:�G�۵�}Ϳr6��2��nwm�E�����y����p�R�󛱏&�m�v���WS&��>O��$��!��}jv�-Z�_/;F�3K�:&9C��S:8�yݣʚ�zx��ڢ���M�H��<F	������J�7e%2��x����E�� =��kK'�l������בOk�@o��a�m�ў���"��� ^l�`�eH�X}�XA���ql���e���fz���_]�̽c�Y��J�+|v=zB�Ϟɳ�-S����!����/�%e��Q 8ww�hzp�) ��)�cK0R\FHx���*���%��S�w���$2��[�;D@9m!���!��-���L:��c:>9K`��sn��5�:\�}�9_��7���e��O"�����b��=ٳ8'���kZ���8��1�Vp�8����vL��Li�;�H�|I����H�� x�C}�#^��C�3rB��_2$B���|d��tsx��,�|R1�C�K�fŅwH������O͘�de�h�?�r���U&`����$ӱ�[�l��y��� t
�X �Qp@�,��{�BG�����A+�QU|A������6�Y/�-2�m ����6׼��
|13����s��{M�59U�O�*�;�*��;hM|mE�5�������<��6���8�&�3�*�,��U�Jei)�,;���3%j{���YX�x'x��ܮ��/��������g���Kk�z��7�ߑ�??�E��S7
_]�E�G-�E0d@��.����EY���������v^���a�����+�\�b�F�틋�����]J+{h�Ժ��Â-��2й��m��]���Ï_i�X@%�u�ӽ�R� rТ*z�3��)������l���������}�`���c����Zڽ/{�V��|���(�:���V���hl=J�u��ɄL���[l�9;��3xlTS�BV�z��S����D{��$H�s��O�u�%��}��-�<&��=ew��fiG[�C��+7�/ S��T���^�w�Zſ����K��j�^���+��e����b*dP�[�]_�ϸ*�Ccu���)Ha&�҇q�b�e!�S��������g��>7�`�����{ȶ<�I
�]'�Eb�G�(�ށ��_1�!�lR��m�t�Ct�#\�`�����"�V��&#�^y0`�(>�UU��uI6��D2 �슖1Ā�1�1v&,LH,���/��.��/�7�e~~����f�h�;��Q	�>�=������$W	pp��2Nu��t�O��>�p��a��>Q�ca���dU湀�:��@�o�
Nz9�O!��UqIk��B���B�R�$�8�����U��e%��D�*qT�LS��y�և�q��O؄E!�����9F��]y���z���*��Z���r�-�k��V��p)���c��js��}��k�	T��^�g��r�gn]�up�ش�]]��;�H���M��w�gn��X/�XҠ�w-�.�.��kl+��V�NI�F��J
FJ��n3�?] _d�@Q�?W��,�յф����1gW�ԏ�K>p�3í�����Pe�v)__ҙ����{�����gfY(̕�6�f�t�݊�Fk\2[�rd��X���b��35e��'%�|h�'�,�f�2�2���jl��ے�ڥ���������?k�?1Z��f[l+e��P�\����*erE�X`5_B�w�9� }� =�Y�4ZA"�ğO#�9��he�����,]6�����uw��N����f\�W����_cR�ٺá�h�:�G[
K~��V�DA��ϲ��GcS6:��HTM[2T0XÏ�4%����"u���Y_�I��i�ҳ�x��_�mJ�pt�b�,�(�ܬvZ������:}t������	������d�����L���Ua���5_̺�n���%x���p;b]~�躪�:�_jQ��c��7*�d�H�l1cK�5���WnV�d��URi��t��1D����jX�`�8�X�< u���tmTٛ�y���Sw!1=�/�͍u~�cx��.��K�5R� ��|=�k�k��Z�m��m���n�3�v{�J����%��W��)Q�]vH��&����I�eVh�]��]��ʴ�R�}�W�=�+�b`��e��]֠n��l�x�^_�1�(�-Lĥ >���9I����3M�8�Qx���,)�0���k�o������G\u���t-�9o�h"
@�u�����{N��o�.W��U*KLE2[�A���=�]� ̱2ە��=~��1�1����k�\��!P�iРX�\g�n�
y0�[Q��	�-�ْS} @��l��;0����x�M z�#u�j���J7v���-'U~�5t���뷾���q,�F����*�Z{��e_4Ǻu��^��h_'����9$�wǗ���5�M��a�A]m�]~~|O������&[J^WI���ak�t8�k�f��L��q->��(�jv�.&;�3JR����87���^ژ/4���P��R0��ݔ}[cC�U�&P�`���-�5"z�aU�L�ql���7@4^0���s���$8z�$�`�����, ��,,G{��\��hkc�+�:��4�-�g?~�kԟC�8a�?�����'�wF��دz�@��K�{J�?�.�|��֗/�X�C��Mޤ�>
����2�X�����7���e�=,lx�{�+��Ӻ܍��!U$K�X�[W��w1�]�o����\�j����Z`��n]S�<*�{�Q>�@T�67����'���ʄT�`�����2�`�������7�P�?�Y�(WD��"&n��P�����i�G�c��T	��)SqA�MX�����F��~I�{�U��E�.1R����`��}�zmmps߻��2(����j{��p�����Ʊ�]X���U`����_�����1�џo���q�?xt��И�N~]�����;���p����4`k�3G���i��JQ�v�_���.��̩�=�6���%ea"�5�$�
�Ƚ�&�9S�e��3"��\7�6+�n�/0��������x��l�i��f�I#d������� q�:�ꅙ�����=+X�<���j��=�m�R�����xGttxL��	��L�o@�p�Mۧ���2�w�gߧ_����mY֞k�{�o�%B/�^,���LPh�W.�Ҕ���w�������p]��{&�2w��J��ǻD؞���5� O�ڠU��[
�6�k iV��
w��+���
��t��n��"0s�
�0�u�wi�Q�V4��ﰺH
Eɳ�	0� 1ʅ �g�cݍt��v*j�t{\���ل]�~���,�^*e�z(�>�)*�&���+�{�>[���^��ec�ߍL0�+�m��H�б�4��2���S.�b��#
���u��k6�P�3(k��p���	�_dɽ����W���>< �����e}�!r#��~8U���+��%�gU3V����n_�Sm
d�+��檭K~_<���������me���E�� �l^��j��͇컴a�i�:�gSČX�zo�`��&i��s�6�*E�L��sT�l���K�~=�F�"���LMP+���0Ʌmnn�8 @�޽K���w��-_} AkÜ�)���ܽ{;	�*)�K����"+6?J�]��>��z�@8�������U�3ĵ1�/Ud�^g^\E����׳���n�Z���(��DD�Q�L\�r����i;�E��(\u��V�b}�}_
�U�U}~�z�}cG��k@��9�{��&,M[Z�������V1Sj��-`��8G��SfuM��QT�-[sd�$s��g,p��晼�)��%�OO2Q�Ʀk��CR�X|���ڀ�h55g�X��Ŏ�UNɖ
�H�5�Α=Y�E��Z�!�ߦ��r�z;pIp?�K��lVĎK/;B�g3h�!��k�f���6�Npk��%�w\�-�E��vM:�������}���� w�e�cUSB�rZ��W|W|#�_�`p�	��߿� �9x��12��}W<�=m�qsG���r;U�x4��s5�I�k�9���9�g� 	����ZJ�J&���~h�cRE��M�dԫ�5�,�?=L6�¿�3�^��(�F�J 8! ���w�Bp �ߢ���-���lon��;7�]�����
����+D*����$�I7X��{�5��4�F�i���)-�_҆|7t������7w��V�4t�:���}���6a���d�5]9s/;<�پ��f��6��� :;oUP��̳�xI�r�$����y�lo�U]��<g�1ªX�H�j��d&!�d� ~'j~qu�0w� 0<!zQ�{���{�AtY���� 2!"gd`���f�/�'L{�8�i�o5��Yߞf� �]����H9g��b���)�(�7`�Z~O?w�!��ugN[��ئ�"��X�����6R��˴�޾��WC^Ι�������ݔ.�$G_�{�����e�������M�K�Z=��C�&�}}�g��I�&����y��,H/@ҭR�jV�0]�O��%+�b������B�U��-% .|W홄egS#����7۞D㧽�r�
lv�vfE�R ���eG��SP��P���n>�^Q
�\0�h���0�	|�!ô���Ay��Xn�4\���noѫ��B���ѭ[���e�K[�K��z(A:��d����k��B�sD�?���3�L�Q��r��#�\�Gç�����e�X�vZC����x��1dV1Є�a���d������J~��(�/[3��07[�v�����U �*�������T8�/�;ѝ����
�5�+Ђ[��A���ӵ���u����e��D@뚸-���j����-~VTD�o��`���}�wfb�V�z�~#KP��i�]_G~gH����T��z檁{T��h�5�#^��,I�;�"��Ot)�]rߒ��s8E���Oܖ~��$I>.Z@o;
�l�՜��
N)��%t�� =�Q��=�3^���ZG�[���
�*���uXc6��yگ�O.Gk*f��H��:��`w]��ha����i�8��+��E1m7��B�PU�2E��V�O������R�6�Npi�<���uʀk������nn�K����m���ˠ1gC�ܨ �������1�;V#���5�P6�@U�<{��&U�m�[ �1��.*�9���L�w��\�D�pS�i~p S����^���XC-k�S��w�WM�&��Xh5G����C2x�츳�M��>��l�&���>|��c�)jz���Q�։u�n�K3����-�+��GX���(���,�~��ſ,��/�9>�$��-��|6/���L����n��l/�B��.�ej}E.*�㵘��{N+�b��Ϳ<�mX#t�6���v�*}��������o��!0j�s��8��,qk��Q��?�<��Ɓ�	�t���:�G�{���4_f�(Y'����y��"�^����1v/����s7�rO��g�� E^B�P	GU�-�Bc�)8f�5=�)̩�-�Sw��}q�$�I����B���<_I��/�����Rr8�#�ɰ�YA�<׊���H� l�ț��t���D(�.!�KZ�S ��B��~�!^��f,b5�+����.�v��*�/�����6�����(��	��*�H&��=m~jԗb_̳�bI}��i��x|����+'/I�h�y�E�ZU;\2A����:x-�${�C�+����-��j��c\х6�M��5�.=�4R��X����9��Z䲘� Vf���U�KJ�L��3)������*o�e��RA���>_�vh;��m�m���g�F*�v*y$8�T��H%1\6H.�ӣn�9Ou^���˖��_�~����埳Ar�����5@eD �V^#I)����Y�&� �e$�wT��%,�3m[�-$Ͻ��Ak�7is�}��tr|H�A��&MK-��)1<gc̅Z6��9x�e�J��w��Y��<�6��R��A����+�m�"V��gU�&��k��BB`�M�S�}�b-=�A�T
���VCNΏH������,W���KXc��u���HHEI%rS����)�"4M��`��2�� �6f~LL1kKמ�]��z��m�Rh���V&���	0��4,
Q�.J����F�c�LN�s��r�sk�M��.@��DD�1+c,t���[ X�R�+(�L*������959Ky�����s�}a�f�y��ڲ��yd���ݯ��A嵓�SQX{�<��ZK�����b��E��O�
=�@Ef�K�F`W��hI�7��R���}3t߿}4Ғ��b�7�p_�X�,89�ż畁(Mh�9h�_|���m�B��f��g�d�K���`���}�ړ*��<��Y��Fv��(����6��^��e�_�4�Nz\�(e(IǼ6�H���N!�t$E��$UU���#s��C@H�M��[0�Wt����n�F>���0,��rD�����g��VEpŬ�Y; Pp= ��-1%���`������/=2����.ݠ�ubl��MUp����L�v�������ś[%oO��P�Y֥�32*@��lV$���j@�7���9 ^x�̾��JU��upD� �ÂU�ڍ����|ծv�V?mN� �������O�� 0���E;��ؤ
��S�)���n?;Ǌ	�ua�+F�����UX5d�@n�w�y��z�-:K �������k��Ʈ$H��3�Y���q������v���.�����@������?M`&���E_¤�W�-�y6�5@��=��[�n҃���7o����t|t� R��ԏ�0��y��e�Ux�H��'s��i��e��}��gc��w���3��?O2����i�)�rڕ��:�J�y��aJ�!.g9S��8����\��c��X�> nVYN+A�
q�l���2͉^wN4f�B�W�=��w�A�(Z�s.�j��ca�cc��ݽ���lf����M��ݺ�W��Mq��wdkg�,�Y��f{��憖k5�b�:Wj_�E|�c��څE4��6q��v~�L��	E)"/�1�ht�����x��	���������F�ᕏ�^�]-������7�(!�r�����fj/ ����0|�Q]Zr5�(�>�YfTcy������ϳ�^g j�2�Mϭ	}�6�寓ͺs%�5�T����f�nU��#��n�IV�r{ܜ��8�Gv�W��P��7�͕)
��z3苟�W�
��,Wkm�À T�A��6J��> � ��5�{��m�]�V��
C�m.h��cU�|���**<��8��
��{���ߤ���:<:f��O>��NN�)���9����F�w�F��~.��Y���y�Ъ�����+�k�{���#�VP��8�����p���kr�/c��9��w��r��$NtD��� >��f�^m�2��r��	���^�6�z��:E��W�D���*���5Jk�_95dY"r[Y[��OP��m�����+:����g�F���#��*
���Ar/v@w Ey�%��:?��_�n�^T�
���{�d��|�Ε�}�9��/��;��!�[�x�e���$&_@�sIvLo���ϗw`�-D���B[����1������DZ���������W1U\r�֓���a����]Mˇ0�lү�f;� �~;g��t��-��١�3a�O�6�UL��m ���	��}`��L�
���@ww/�vw�Φ�\�!3{+��캼�e(��5BV���8��tF�ǩ'��&�����?8$��$����l�1�i /���9L�S�8?��uq����4@�����k2�B�-g�tN�	�N�ɓ'�6^�H�*�n1P.�U�؀,eQ?��������l��g`Ї Uh���!��e��ɮ)i�T��,^�����vj�5�<+�UY�����]�3Q�0��n�o���iE�?���-�/���7�>���4�\0K&�I-�Kʞ�[�5���=�-��-+"�w�@������B	
��$,-*𝞝Iѓ�d*�s����?b%�����9�9��8�1`��J�Lr�>{F|/|kq��;;�g�lkۻ������� ���t�����K	�*Ư�}��-'$�B�r�n��m�Z~�n�;���:��Pd�d�`#�:�#)nn�<�z�T���>�4gn	`��2X�}b�C�,0�xq�m�����4��7*ђ�Je?~a�����lG�\�� w~5	��o8F�)8�7;�RL)�z�f���,��NX��q�i�h`e�]���x���{�c��Vd�|�Y���o�|�mKN��P�!hz���@�hNe��D%�g�T }���5�9-����N��$�k�`��&V�~�r�jD��uccf_!�=�/�)|@C���IZf^��x_�%L䗕�l/�e��8�1�m�6#��S 30/c!�=���S�6�y��Q��?�-q����X1�B�"�^����L�=l*M�3Q6��E���4!��{�'��4��� L�����@�~%s?F�2�]��?z|rL�>�6��S��#�jb^dK�<h�{g&��k�`ct���S?�w�+^y�z����}NO�>��E�:4a~X~T�["�? �ww0����D�\����!�F�n.@Z[@Si�,�h�E�}1�>}����ɣ�	LN���0�O:O?����~�P��_`{/1sc�����á8�¼����z��k��67%�l}���`LƩ�?��{����st@��x��ʈ	�"0J뭤lC	?9=�ǩ�����S6aƪ~��&��i��,��!ʚ(�AP��m��sɿ�y��:Z���9W�M��w���^�J�s��Ow2�Hj20��[gXuE��`�ǉY��kmH�阯����6�Oi�d�oKC<[��C�V]���ڧ���p�~����ƱpN��Q�k�1D������k�5�ŴH*w- 7�T��uS��Z+���%����LS�bݵ��0������Ll ���/�hf��������P�=
؅0�.Ğ�dUrH�� qC�����i���j��_j���f�DHb�\*�����l2�5%�m����h��iɪ��i5`�	�u���t��^d���o��Sk��6�_�Ȏ6��`�"K�+&�M����	e���+��*m&��)��,;�51�W�K��QY���`A�r+=?F{Of{)`����<����e�6���3�m�{I(ݠ��6G��w���Ae4:І{�C�gI�5���lLȝP���s���(��-˝��>� < A� �'�@�� ��Y��6E0���:�Lx��-��@o��ݿ�>��C����-}��G�O�G/'��qf��@��W��t<�픝XA��y,�}Qţꉢ�6��������!m�����kf�'��a�8�_��W�T�b{ڡ�/�3����͖̄��y޿ѷU_����ꫯ����A������믿R�5����*)%��M`z��N�눦�1+e=�����{?z���G���'Og�}c���#6���-��j0>�V�m��~�Eᰗ�w�*__�<ZA�R�z	���8�n���|��⌭Sh�����KH5J-+���^_�Ȋ,�.��H�&��Z+�um��f�sp'v�~��y2������0fX����?)����ީ�t؋T�<�t�t]����[Ȱv�b�.��>Bcb�%-7?$��x�@� �K�� oGx,�	j��i (�*X�Ƀ�G)ED��"g�@ E�����؅�P�I1N�|1w�P����K7%��+e?/,k50G�n I���`)f�Ϧ��$�]�trfwKH.>�ӹ�����>�z��	orlrV��es�M�ż�1���َ�ik���D�j"EЭ������D	��5`g��Cn���� J�$��l���>�ނ��3�L;6P�?-�N���� �o�K?uM������  ���°�7.���xJ��+��5X̓x��ޝ����yVm=�#`e���$̃/������*�*I��h�P�<����
Up D�_XYl�� Sxn ���r	i�]M����tt����7^@��6� ��@^������x�&@���@$Mߜ��p�WA-j��*Y/²�9i�p�w�	4E��O�� U�Ҝ��k����������@��W�gV��r���%��NaQp,�z�̜��)�Hs�0${ʭ�7��{<6��.����iwy�� ��O�>����,$.8;;L�p'�;IyW�ϊ�6���(x��'�����^�;I�9{�}��g������tMo�m�����7ᗱ�t헱��[�Be{��A-�U�1+�Q��9����ʷu����y�����ݭ4��ϖge�;Ժ_Q�iW
�<��E���:�`�⚒���@��"[_ָX=zX�U��un�}D��#s+�gHa)���!�.��9pF<_�l}����1��2�k�J�>�
9�bne�4⏻H,?�-��T~���}����kΣ�K�ᗗpC��l�"L�o� ht�y� (�{�6�`6G��<t`���X���� 3.�(��sw�)�A���G����{�
���Ȝ`^�� `���d�B�j�s����u�#5VZ��i�٤��˅�c�&�t��i&!ɋm&>E�𦅗�\½Q�wk^J&���g�.�����ҕlwu�g��k٬��KNu��TЉ6�Jl��� 
�-�@j
���?O�}�� ��g��3�A��`�Z���&ij#���A�׭ ey=�B�h�`��\����	6�c�%!^k�P��v����ns�@o�~�"񽐢�3���)[��<�'t^s��) ��,��e�d$��g��0#�DƋ|�k���u1:8I����o&0�&K�H��XK�B�p�F�@�� ~�c6eל����W���b��+�OsQ��\�R0��n�ה��J60�o��&��ƛi��o�0l#f"O�o����O��Gl_[맾�A��ݥ�����'�$��w���/�8t<_�W��=uߨ�y�h����(6M��\���b|�D����'}�w��e ?W�{���F2M2{��
�������FN�X,ײ~)��i�Iv���������O~�Էл����|�-��;g������y�}�ŧ�����VO�]�[7w$��(E��|:��@�=z��70}��?����Dvh;`�����t��Y@�Xj�<���K���e�2�%�(0��������E���96д��{��J Y�c���t�s\9���y�s&�eA���ϵj�)e�fՊ꧍�Y5��Bpk�g���M[IqI;�5r'=�ӴO0��C ��6�L1p+��Y���#P��뤜�q��G���v�.���.������ -'[]�-+L!��ɗ�us;�H����	�H��lP������,��=�����V_�o��A*�H^��*��^�=檎�v�"�]���ϼy��� �#5�¨95MCSl.N�\����u���I�A��pEZ����"Y����:�į���f��gxG�s::9����H��p��S ���i�k��fE^�d�)QB�ͭgK���K9�kc״^qZ(A���"]j�� Q6q�O������}#�l�i.�k�dVI�
�ۉ���Y�f�@��JT���Âil���79��[V�B���)���Aq���򳀵t[�� �>�,���솑�
����13;��Lb�d\)������e�s�6ݾ}'	�n3�7r������9����n>�,x � TfS�Qg�N��|
bj�ݽ� �;4W��'_�W_+y�<��g�ӖN�2����̛ϟ���E���/�������/����������{?p�����p��$����'�' �����^[���$p|��x0���ߠ����7��ۦ�տ�U��0I�9��T��[��f'~�����)�Ir�����9��M�+�4��D���}fl�����[}�Y"B��q�NS�$V�9��<2	 �넴��o�w6����O~�>����U�{�	pMh��*�3@��X������4KW��%�S'����4P�ϕ���27�"��㓣4�n)�,�6�ukA�ۦl��`P�8���'[�ms��T\"��Y=ܷ���P�/�Z�ў����uzd2V
������* *p�Ԃj=a�<�g"J\��y���\g �
�\�T��-N�m�x-�*�����Պ�Oܨ�i]�N������%+,�ќ���!����z�ͷ�tג1Ș�(2[u �1��kZ
��\8M��<c��]&f_"Uby^>\}�Gfuq��c#�
�
��X8-�_��2o{IA��nUe9e7�yo�6�^}k�b����ki7K޺�y�g��;�	�K�u� xˬ�,zI&��T�`2�+;����j*���=�>�ZO�Gd�:�yS?l�b#����6�f"������`?��%�{@'��#��,.X?m�2��2�~����P�>hEXۀ��c����r��fӕǩ\!���ָ����{t�b�jт̈́t��T�g��H��ې��M^�SPPf���Ӿ��w�Q�P^�'�dY����1��5�msc6��*\�p����+�؛k��TB�r�<h`�M�~���́�ڀp]*��vQ ��U�T��%�Q�  d������TN�8llnd XKW�Ӻ@��4.I�����6����pe=��j�VB�$����V�l+��M�5=?<�*JI��M��m!��e����U�v�O1����`���ӷ`o��6f��	�D0Y$��	i�F�ܮ������S:����<g���iI�Hu��ܹ�x<��� ������P�A[9>�TP������}�/�[w�����Z�=�cf� @�s��aS��X���f3#�F`��Y�/l<*.��M��gԙ��� ecwv7�����Ř�����nk��e E�3]�xd~��r�dB�	���ܬ����~0�����j�:Ο6RC�n^'�u<�j{�(%n�X��54#��;Ƃ5�gFc��~�3�7�-�\I5(�m�[��&p��>�ȳ��#���L�}I��X}�N!�pc�A�;�:?�?�̄��)���d�2�H�%��In�>� �����O>x���o?�����$��������4��ݹ�E7�v�\vc�b8i~���W���-�,��P�%�+X-B���+����v�[���m�I�~ب�f���v���kȿ��Z":�2ހ��\��H5u����X��*#m�������)rK^FI�3W�6��)AiZh��� �&�[S�����cz/$�~<R=�|m+a�$d�.U1�����{dy6��1m �$��Fۿ�6�}�<}L��7鼚����dtNu�H�M�D���ד@�mQ½	�����V-�S�㪫���"Va�qݥ����b�ɷ�K/��zU��s�4u�&l����������d�ؾk�,��]f����.%C�0���2QqQ�c� ��}�ekg);5����9�{-���+�_�S��*��Ϯ�Vr�T��L�+
Rfӈ�[Auv�`���+�o��%��.c��\D���ό����'�"�� �������"{���`��~FZ��w^��$�������q���j(��#�H�occ'�#���]z�p�>��kv#(l$�L&�����UyTUA�Rrz|��:x��F���)+�k���u�::I���s�/��/XH��5Jc�@ؚ0�'�!�/��>���}�3ڑ9;G��I�#:�8ePUGI+E�;����ʡ�|�>������Pk�6)�IBmS�}����+A�Q6O39XI���ɒ����*W�{�}��K�4�2L�`Գ����'e���4��Қ>g&���R��w����i�&Z���3VB.Ώ�u�~�9v}#���t���:K-��)���jg岽�3���'��"{�\+ɕ )�筧uTq%Ê+8"�˲w�
�����[��k� 냴�\��*�����o������b�����٧����& �� ��8�5��@S��xd��H{-���Ș���I��s�ʫ���6�p �M?�^Di�o�����f�o���<�C�{ki�\$�{��|�~:��io�Ir� ��@��r7)�I����q����y��w6e��Y"*s5���ls>/�[��: �_���U�Oq!7��2Oe=�us��\��J��,�E�JKkR��cDV��[�KC\��:�.k$פ����C�i�4AT�7s�5[����u����9�̪��e��L� ����~[v���T~B� V�zNSG�'"�zQڠZ@����
f	'=<���)Mc�8�9�
�a� �hF�ɜ۶6[�����{샒�r���J{p|�\k0�z������o\��Y&ă�ڙk�o�� ��k����{�8'*�0�`a�>���c:<<�<�x!����r	� AXފ��H7eϴ��ޏ�|{'�>eAf9E��� �����\�����;c � ;��*RHk�Xv�`�֭�첖;���f�j���9%��߾s��*��9�5Ez-�':�J���$� D`�Q��0���t�A3 �s�D	l�8�O���kf�u^G���!}���'�����~�ٜ��+�˽y^|KCS1����$��>���_ѳ������~�'�����g�嗟I��X� �0��>n.#su��� ��bN��BYشG�)x�AYj���):�t5@W_�2(~f���������ə�Y��X�@�J�g�;Q�l	�.��h�-���nmn��d~����@R��n�z�5э���[ז�_�Nfb�RP3g���|�B5�  �0`ˉ5����-V|7���'e��]J�̲�̊� I�����M�e�2�>���3�!cz��nr�;�(�899�?��c���Gz�����v�P����vv��������?�_��	��<��|�ɠ�c߄������U���=�v��{&�e����8_�X۰�#��92,����B���p������72ف�`� f �����	4���	��\�ǚs ���&�_=�����N�����i-	�Z[������Q��L$�D�̫�g�E�#��_����q���'\cJD��Qޡb�>�h4��}�\Z���Կl��{ąS���FoW�-=�i�����HP�}���b��O�ֲ`xc���3���2���~�}���O������,iIßUc�����H�:\_�����U0�m�+m%�K����6J��N��o�����6���WpS{���6�8��#�Mۙ�'��y;����
u���]��|��8�Gh�fL���0e��D�@�2��4H��Uh�M�]l�?���g?�Yڸ��m ^�щ>���'����_K�1}��g���S��%%T�����P��[a�qX�F�!�C-�pfi���A������C�!��N2#�\Ng3��~��V
��:P�Xf"���m�]I�c}dx��)9N=�$���[I�����إ��Gҗ��>|��������V�Ǜtt|���y}A��&z�.F���R�@]zTr$<G��5�����ӿ��!�{�Fj��[���6z��.P�'���@�" P��?�?�٧�pYk�p��	�?f�}��Qv�98xƩӸ�hO�'懔�J�� &Zv�{#.d0�J�Je(�� 3��(Ơ��x�2#���RK�f��
���V��{P��B���(9H}~=S�L���U�ť!��z��dp�m�q�V�뻹�1C��Ρ��5�N`?��a��ي�nA*�[7o$�k�������~�����a\�Wܸu��,���If��ɘ��Z"y��V듹B�jkޗ��0E�������歛�������:�&�Y��{�ϊ��"�#r���.��7�^,mV�����w���IJa<66�8�|�HOO����f��T�xXS%�(�v�X��`�`�I7���k�;��D��jAש|� X���:cp:���@!�ys�^}�vz/����t���t��n�HJ�ƀ-1��U_֟R(�x�DT�B�Tl�X8���_����-^qa��o��k4��I�f+����3r��=!�B���U����7��(�X����,6
�])hM-Z��|�֦X&X�L���*�ئ��V�k�4��6c�9#�|���bV7�i��!N���Mך��Qq��PS�P8O�3�Uz�:�j�H�S@�MȌq�I�#�aƞJ$�d���I3�hs��OLm���&�t���Ӵ�N�溎���I(�$e��$���U�ZTeB$r��$�oum�,�m�]�w���oe����DNk���A"A�����6�]����q �NՔK�Z�x��Io���>���.�]A���X[T�/��������_�����a��_�럙9Ae,� &y��w�Nabp�k>�����e���i��r
� �ך���ݣݽ=�0�f�����u��m5�P���3��f�FV��!ϺIc`�pϽ��TUU\d���sz�����X@�Q��`w(���[�F�Xܜ�+ *�af��@^���2�66�AP��������!m��_��|X
0c��}�V��$�ۀSIF����Ԫ���z"��jV��W����9}�0��z�h���Al{��{vz�,�l�������W���-�C��Fg|�o>�\�`� fF�1�cl�L�DV�{����F0�TL����[��L�@J�F*���<܌��gc3ϧYa^�s�G��~�`�VLi�u����5����
�1� s֐��	U���J�B4 ��>��G��L��p�^��:��=���Ѝt�g�}��v�@ңz��^�{�;�ޮل���>�2�=gw�0��uR�����I�A�'y�e��L/!�"ў����	x��,�Э��~���/�~���	뛬p"��(��;��Qe�Gǔ��0�Ä��*,��'�y�&��ݝ��č��O�D��C�կ~�k�-e�+��=9��ҟ���|$���8�3�p&A�P@n߾%�ZBL��5�mn~�I������Z����#�2),(u=`� �\�]����qZ�Gi���%�戦i�!�v��te!��.�U�[V0�����RcYyh�U����O�+{��K�@]��:f�ˇ`Ki�p��n����>B����@װ���\�C�U���[��˼�"���g����^��p��3@�y3u>e�N���4�G���O��Ed|��_]�9Mk�v���0�g~@�{�� ��\@�|�.���i���4I��b �������i�%`��6�}i���x&�UgS�!���Nm����`�2�bvȟR�3C���sud�9��A}1MJ7K�}������ih����������b�B�>��2�eZ����'��R��U/���涧}�i�9��ܟ����O��O��;���D�kp��<M(��-@	��z�mn5X��>&�ű\� MƢ���� �����ڃb	����1* 6�[	�ol��@��f� >�%���9=�yю̈́�����}�g��_��ߢ�?��Ӥ |M��C^k�P������M}�����g!�3eZ�"��]�AG�B�G*9�G�)�0���5�3ֳ�/��곬s\���0�2����J  L�f=ɿ_�%�mϙQ(�y�-�sz&��������3��ڞ*���S��g	�BQ�����~o-��N��ՠ�������߲����'� 衬s�O�b�\׫�����5匕��J�Dg)
�A�-��8�`�քg�U�<k��MU��Yz,�0 e���^�G��ɸېX5�h��M)��N��3`gf3}���3.�qv~���n��]:}k���()X;i�ly;x~LO?Ks�h3�݃��7]��ZV���ͷ�x�=Kc3a%J��94V�c\)�F�d�e*:��H:e!�\�~���ϮZ �i�@�6�d$��vmf�H	���JxUcO�u
�[��w���������?Ԣ����7��Hٷ�J9
4��d.H=����_*��1\��Z#F\�n���{'��7�|��޹C�I���4��W|�	��/�>ak�x̬�����l�O4+ǀ]�$�X�v�Z��4� ��/�W9<�ܘ�z.X{�W��bx�#��*���uY���Z�5��&e��"9�6���	��w?��FO&J�L�o�#w
�--�2d���hu���hrh�	���0�`�Z����4m��~��،�O�]�K.9 	��(	��'���$	�#JK�f_�AOX�Ӿ��C�I#^K�pc����b��sN޴ُ'HG���o�0M�$�>�iJm��	�TS�Vc�=M��}��D��eP�[݊�f�BW\�p_�rrM AΉ����x3�a��4�W>g���/��s�œh�f�8�<*c�.\���s�.�e�@[O�������'_~�%���� ����u&����@��B��9�8?Ov�r�r���e+���oj�m͌FT@(��������G����"4�R�C4f��J�ѹ�瑲�7o�ѽ��Y\�R�tH��w����;o���$��df���]B�/�V��N�vR�����o>��}a�6T��yZR/	�O}:��w�@����[�ME�vೃ���'釖���.�Q\R�zXJ\�޽�� >KoN���1�S5�ԆlQ`gOr>�8=޿8;�/���n޺M��Ym�I��_~�V(:��,^����b4���X[A���sgζ�[���`���e^�<o�+�E7�k�Qݥ�}�م�d�Mv����\��R� }�'V��{MU��{]�)`^s�1EP����|tF_������C�~�%ݻ��3T	�"������@�i��M�g<~P>���c�O$�m�>����;>:g��4�u+�iۜ�M�ͧ�k���&���PM����� �yyzD��6�`�U�K ��@����g2�
� ��?�?��<7q��@���ŮL��D�ff�����F�}̃��͖2mn>κ>,��1����i��^"��&I�]g�׻�Mw�ݡo��*)+�p ��T�q@��+�a�K������'�/�ulc��'I��_�`���Y�gxM�*~��Y(*��! �/���68$����H5���H��B��}o�Z$����b	��V��b�B�iC͏I�2`a -F+a��B9�ؔ'y=�d���N�ٝM����I�PC���)�����N0N����i��`RO���E4�"���:��_�M���f��M�iC �4J`��{uL3�ԫuN���֓`��)O��$r�)��|Ĕ<矬ku�e�z�_k��r�#kT!��J�.�q[�T�E���Β��eo�+��:W`�B��u�o���0<`7�w�}��4 �c.%�5}�6H�=N�� n'	C����jzݼq��+���{�}�8*���	�Z�,��1�k�ܼR|` �k ���a�+� ����S6*���6!žl��i���a���;�UL�?���fm���1K�k"�,����GA#X
��H� ���}�LRg�oy�3���S`�~0�N�&��}���L��cs-҉��D��5�f�Y� ��i~�Xq�k��L�ٱQ���1mQ�o6;��p�2��hun��?�&�,~b��5����g�8�͔������Ey>�N����$+�K���ϿN
�����8��7I[��ȊP/��¾��̀��w��B�R��u=��_��s�C\p�Z��&V�U���l|�+�%�����'���r	\����J���	n؜O�
���G�,<�3��ӓg���}����+��k��웯��y2���;�q���/�cG�]f���@f|c��8\V����ӮM�6�l�z2�0��춚F�����M��M7�Y<�v�G>i�o�~��g�l�����̰b3eS�9(�܄"�)ե�!���/A�
xa�0W�Z��{J.�aD�Y_��ܹ��p�]�ர�@����O�B���A9���$�/��	��Y�Q�6AO�Ù/��}}�1[,��y�^�X6G.�Ҫ������b����;��ך���[�+�cv�C9����ƴtp�*\���%m�x��7�e�q��K��G�n$L
g_�ܩS��JR�z�ˮx�̏j>Fn�i�b�6���rvzA���^`1InRCڶ���1H^U,F��ͭu�w�&�L���/0d����8�.�+ ��&4_�?3� !=���D�ƙ�WCf�(��{�*bՋO��,f�r&��>e�t�BnLX�����Uk��[>�icc�l,~�k̜C��S�����7ߤ��{��d1'��r�~��_Ӈ��>��O��K�u���M�A?������"�,����o�_��� {N��ެ}Z�U�:�k�6�]�I02���M&I�"_{�U����O�� /|D-Eٔ�I\�T��@�(��J5�kal%��|{�޲G�<������� ������v����>H��F`@a�����
�����������!૟˹��4J"��1c��Կ��)=z��}!�P��.Z3.2��WI!�����cfw0X��=J�J������Jm���9_�O�[��Y��@) `{���v���$��/(�^��{K���ň�=�\�����/���#�f��?�����5P.Ӎy7(eW�3��yI�ֳN��suC��=�Ip傃�A���,
�+���� �v^��Q22T��d��"��[�>N����y���b����ɜ�m1���V�����i�ʧ��~�t�	��5����Cz��!]�aG��Vs������M�;>��-i_�$Jh�<�Z쁕�MvM髟2��߬>�hwɗd�\�ܘ��kZ�����~+�k�\���#V�}�썛{��!�knp�<A.���=.�rv�g����H9�\���(��,�楰�*W9��IHQ������u�?���O��t��<��ꮾ�A�(������_F�_�ٟ�%��G��ﮪ�;�_���=��� �Q� U]�����gf�Ƭ�AN�l~����)Gj4-�[7����u�D`p�X#N�N�|rtL�����kh"�0�1���a΀N��,��0H��!����M��_'�M��\Z��(�YyTI�e�[����l��d��J�f���>�n��<O�,��{NоU����v���ޮ���|��/Ic�/�����mgq�y�����F�=�c��������8N�h&g`Y�0��H$Ig	)Z�e�hk���_�s� 1֝��99?�\��b�ZR�VC������|L���˿#��kXH�,;C.,T$ݖ���|���C+<��_��c���d`�W�޻F�/FC�  k G�3��8-ȏ���4���o�[��_��}�.���� M&#2j�g�!��g?w}�S���3�=�������OK��!7����TϞ=#�k,��n0�
��ϝ,��(�D�1
�����{��<^3 ��u�3�$�jƯR�bɭS�Om���;�0�����c]%Xfr?4u�J���H��x���sw�{����=��hH*)�A��L+�E�`��,����+��|��6!�-N�����;�-��I�;#v��޾�����Xh���#�����0���q�P��?�|�64J�{����m.�%}�	�:_H
A3)���\���#���[�H������&o��7ϵ˓���O��
��{��6�¬�9��(LAg���UO>KG�-J�FK� ��������L竒�e���Fv�NI�����{���B���^��+in:�W���>���`l(��{ɵ��m�D���v�r�
�:�u���둼y��H���F[6��?)��i�5@�1���:���1�|���g��h!���������6y?�ч������O�
v��%�>z��8�,�\�Kc�]��C.�8)�+-�|A�h���9���+��2s�o\c$j��>S�Lah���b�SR,]kG5FP�[�Q��2P�ſmlB}#ڨ�'C_��j��$ x�F�)۞W�olJT�¹�؛A��҂�����t�o�������y4>��DF�V�͖��O���Q�����D3w+dcђ6I`�$:�rq$D(��f�L(X�6V��΢���
������$���t�����BRW� �*NV�C�<�`��N�R���;V�kH���K>Z�ۉ�߮��'V�C��9M�� ף��S7��Ӹ��l�1���@������Rޔ]�k�1A((��;�K����]��{~r�.v�#�7&�&�rk7-o�E�Y��UҞR�D�R"�V�����o~C�&U�O�-;#�=�~#�wށ��:UP�P�|VTi��X����+p�9�2��Ў�|r� ��9т�.d�HC�z�(z�N
��6y}��M����V����F�\�_�OY��wя����YB����.�\1���������<� ��
���O�j]�L�
�C[�
2���FdM���'T�8Ǯ�=��X4 �9�S�}5~g�
��o��~���|v(���4C��;��sT����~�s���2g��|�#�K���RP֠Q�8�޷�7ԕȽ�AH^PVI�V���%�DjQ��p)mr*%�6( �����u8�9i���:˅�ak3טݠs��v���XJ�GxFҊ��7z��<u���F�TTir^cc�+e��1��'���D6��STU*Q�A��X�E��T�#�s�U�^:ޱXoGS䨂:��%'������-�p�/V�.k�ʥx*�g�R
�H�ձ]h�gF��x��1z�.���>W5a�-�]];e�y�����}� ����m�1�"8�O�<R�~�v�:3����8�Yt&M�m��*�9F<٢Z"+8GDy�Vw�5(�E���#���z�����/s6����ebPt��jF�h���n1�
��X��)<]��{��XiN`^pھU*��[/]V{��P��_��I�m�-`�ͶD��\2��W|�Y��/}_7�*ɞʳ�1�&�cӳe�x�: ����MV�������A�]·0�a�g�炓�`wޑ�u�h��r�dY �;����Y�'=*�gs��#5t�kh����<���ɐD�[q��V�c���mQi
Oq�a:�M�A3����(0/8����M3e���rf~0��HG�:^�ܝ;M͠l�V�bqR�X�.���4��.TzʖCW�TVM
�0M,R��p�I�^�P3��c&,� 	�Y�?�\��ٕ.$É�q�,�����35����g��<��������(�`Z{a裂Y�D��'���_An�A��X�dL$�S�0��i6��.{�ީ� �/���y�Ww�����y��>q_�c"6��	xm<r�x}�2W:I.����@E�5�-_V��|�4��F�ZAΤ�<Ўs�m��B"��w,Q �O?�<.8{���۬������� �Њ�n^�HM3��I��L�U�q�錍" n�H��[[�d�2O�O� ���]�{�UQ�h�aZ8)������O~�n߾E�4��#MŊ	�y�5�3�4o�E�:�Z��5f�����6��	�è�|!P@;��Vc�l�h��t�։�|)^�0(���ť��퓦,,_c�~R� {����Ls|r�L��L��q��˧��$K���*�6�����*��Ҫ�~i4-�0.�"l�ҧL�r/�N��K����J�����Q��	�kz��+j��BB ������:Бɇ-cKm�����N���e�qY��U�2:�HWXU�� ��)8w��>?[��l�%�,�ړ�Ac#s�6�*����?���Y,�����q�D�y�At������Ś�`�m5maG��v�9� ֡Z�c'qѲxWl�8Vm+�s-s�e���k��=��k�^H'��{��6�Z#b�c!-CT�ZY;ٱ�f:�ڦ(K`���R��ڀ�Hw�BY��.�Qg���xv�{y�/iʕ@tZ{�����a9%&��������]N���u�V�[��_V�=����9-��xY�΅�NTέ���y4	�{@
x��1�$k�� �=�P؍VW<D_���_�?�za��@����P�&l.�Ħ�򩐔,��U��@r+��	RC�!(E��h8���؂�S�f:g�h�V���L#B�("K���C���`��	�ù�JM��̯��s�"0)�nB=Xp*��Rs	;�-X�FoϱX����6)/�z�$�����{KN�qc�z�͒?����B�ҹ�* וM ڶ`�6E�U ^����EmhD&E�|�1�:TiaC���V�{RisYȤ5���E�k�[��hIN�G�c �C�_e~o</(6��w��ZA��Ck���1��4�4�ŏ�d��I�B���{ݟ e�J$s�.��ܡ䶁����۷w��l�"� ��������;<:f�([��Q��M����!og�C�;��}�8�Q��>%ũ����yA�80�xF�	f��������5����s��}��Z�P|	@�uN��u��tS	˲by��X;XH�n�,Vn���nC�����d1~�x��b����D�>��z�m��2з��Lb� �}��V0�C�Wgs-��Q�b�Gl�y��9q�(�	��eG��DA
k���rZu�l�Y[�P�Ӊ%vi\;�c�Y]{)�N�r� h�zd��ݥ��,������&s�]�:�t$�[+�c��	ܩ>�9FU0�&[g���*e񝶸͊lv���tV^s��u6�^j|[�b%��:�30�y�d����*:������, *�������цn�2R4�(3����� �)�eN!W?�T�T��qN�h�[�d�n�M��f/�{���<2�o������Ax>�ZCK)A6A�@|�%�j,�C��U�oD[1T,"�چr��t�s�����K���D�/��]7{N���^z��,�&	V�uF(L�a�P~ޜ��n��m��)����Î���e��K:���h*|�y3���@	���s�D�g+�b�Ep�C ��3 ���A0�XHY 'E`Ζ4߈(����$��v���QR�!�L+Sf8DP�5�����"�q0�~#���ժ��@wjHɀEPq������aEp��|��d��� �s[�Ŵ%k��<d"s1�С-DjX���	NF����}_~I#R]���͇$�Nc�P�F�VW��k�2H����E
^ӂ��A/ �le��V�� ���L�.$�ДB��g�Ves����ԅ������Js�w�K���β'��{>G,�H�.U� �l���
@3���^bߏ  �Ѯlۋ-�n �9��ZHi���Qq�U5���n�Z���_R?s���oG����q�&s����{��?��u<z�r` �"p�H*�M���2".�(x�}'p���)�c*��A��A8|x��� :�������������'�w���(?�����{H���6U���X�F,H*J�X,�g�����*��4@���
&���<��47;h�V��DzM :�5�2�ԩ:�.�ISuپ��h��F�(�K�\YLV|)9e���g���e������Θ[p�=C�4/��0*���u�h���t��o�]��"R�!6�����A� 90ߛz�I�H���=LZጞ�y�$R�E�ڋ����u`=H�l o^���XtIG�t\���T��!���ٖ��ݦIo�s�C���Tgf�,2`j
������YD�I�p��O���L@��͸�mo]��[�W��י[_O��ٮ-D�攽`��Ev�'�-��!F�
�w��F�v׊R���4��ǏFP�%�MZm�2tn�5bz��ɿ":��L�]6n�Ts@�����h�v�S�A��c���YtZӃ���>��maՓ�k���0�2��*Rv���� 3;�orN���#-�բ�DMdn���E���I���-�a��NU2��X�(U���ͧ-Cd��!��|��s*#�:��w�¸�5��p��|@x-��һ�$�C<Y'��03Ri^�!�Aw*�v��!|٩'C����~��Z`�q7�� �i]a�H;��jj�3Q�`U�PY�ژ�y�gi�����W?�W<���$�'1G����.BЂ*_�K�ZU���R�R/���bCxr��#`��ل��P����-s4�X�߸�3��{�}�@`r'z�`3Yذ��v���l�"`�X��P�SY�����7�)�:�6a2jek��ʁ���؂��HY�����r���i���A=����(��^0�^tt��bll������b��Ϧ�0.k�@B:!Đ���o��pa������p�)/������e��Lr	[��mEE@)�S5[ک?!�(仂%�È�X(6�sCj
l 4�׍�"���R,�[�H� �.���ͤ�쳥�n�����Q���6�k�{۲ 	������e�Y�u��(������Ō}	 /r+��h+�Mҿ;M�α�m�S
Tj/�ʡ~E�κ�3h�uI��5B
ejY@�Ya{�l<���2����{߈3�Tb3qLk=�;��,玿b�b��b̖�vuBf�=��ccƊX��:����/FNNC�t�|�\�Yc���5E�� 6�\�]i�DF�:9E� 9�O�=�S���*��}1���{8}P�� �F���D�D;��p�^�.:MYݜM]��2?�u���)�8�ݢD��<:�_��L9�?z$i^���:޳ć���(��'E����(���B�󚉮���љ8��t�ƃh_`��.�( �ɝ�t��va��"�%��#�K��ǎ/�|�H��j���]�u����vcʡ��b����t��v�����/f�L�����UTc����D3d^.��@[9L�<`Jv��ðc�#��*�Ӳ�m��<εDAoP]I3$�V"��6 a�7>�LӠb��e*<@be'���)�3,����.jJ�D��q"�#_���Q�F^q�{�P�F�*�<oz�U�!�LO��˟�s�B ��.�$��[0�q��T}OY���7�1�s�_]%
Kk��)<���`1 F���gO	R�k,B�u����{��t�H��Ps ;�"'����]w���H � u�����&`��r!�b���=R .��V �Z��AB���� "�Z�!<l���ѱnL ���8cP�6J�/�"�����!	Y&���;YK\���� "��z<�R�HS��2kj�e�@ׂ�4 PK{899���*����Ř�R��A�5Oݧ�y��k���x�q���yطo�&c�{�B;�l'[Y���]dIz�P*$/j���U�����3���a��>����,jE�`�Ӫ-zM���aKs��j�%�eiA�?kj�l�˵K����Ė���^�2�\izB��(V�#޺��9�oru�rkd~7X��u�{�騤>�W2��9xu0%uG�M��Q�+����BP�BTQi[c���蠃	F��{������[�,8f�#�_�ݷ(M�j�cU:!�&�=�y�Z,W���z'E�3g�ز��SE�	��RP���"Sw>=�Ǿ�����C̷���4��{��ێ�]߽��sw��-����ٓ��j�T���;g*�#x�T=�P<��u}�������?s_����=?����4���#�Q�|�j�I�����T[@�i�?���c��Nν�~Ѹqt|�b#:����A=f�U��&����^c+svՖ&�kxR�d�^� ��G��v�U�`l�g��I`��f(
*_>W��o}+���FJ�\�A��8�����BB����1 k6��ĸ�!�A����l�:�+�FP[ ��9W�i�XYȸ<K�jr2��n�p	_��@�o�1�;�C��8N���W�o6tu\<&0������o�7����&5�{�b')J�32l�YY8+�4��sF2�d��~���а�nJ����-]�M>K@a���ag%��p��R����PP��!5V�������L��g������ x �4��(h �El��E�6�"F��� � ���`���/��T�Qb�l�i*Q�@�U�c1A+al�{{d�j����b�~���L���)�kh�����!��k�T%�z��晿��N'����l�������0-�ތ`���'�C�!�+��S:��M��N��uwk5o��ʕD���c��fSV^O�@L��I�֞�Q��J��F/"(��c�b�
�%��n��C۵��X܆�ς9����O�2�������y��Xx�G2
">|�g����oZ	9�:�	�u���m�c:P��.�:S.����,��S�eX0��+��pɒ�灭�Z��t% ʫN��Q����#I50�H���sX��1Ή��v֙��/h�-��6��9��ek����ԩ�7odCt��#��P���s�x�c�)��SЍ��."<l��F��v���z�)?���n#:z(�D1����D�o�ھ�rsCƩ��f?��r�M�ݹ�r�c	Z�%�щ�=(�<=;W $Z�..!.�['�Y���b��D�!�Z�]Ѷ��A�N:r�_�1w�2����'O�����������m+�R�4�B���!�S	�������+Q4�#�3�g�XP�b�&m�8�����S�<Z �/�ߧl!���	�"�s΢�i/^T���3w�w���n��+�G\����ε�sY�8���d+ǫ+��ҡ�Įs����,��ۻ��K��[SΛ`'��EOe�Xp��i��_��D�7%�l;����Ch@�Bp��"�;�lv���\�0�m�
�k�T-+L���j/���lMk�q"��l(�&J��nP��^k�����E�D�V)~o9�X�a�3�U��O��$ڥ�kc�l��^cw�w��weg�5�ƅ��-�{'rHHy�Y��N���l1�O*�0��c��e*Y�����5�x�LA:�8J�͔���r9��ڌ�P�FY�&��A=��Ѡ�8��E~��\d�Pl�-/w���?�!��X���FC�}@ �����O2�h`�c�	�
�c�n��7�,b"a� d�Ҋ�5�{�s	[^�Sɞ��4�	�G�ڴ������9�G�.�!��"s��=88V����s
�c���/���s���rN���4�%�c쩽/ژ��x�X���1�EZ��=9���͵p�����E�sq��
W`E��-�1��xJ`pA�!�ߜ��C����7o���3�����ҽt>�t;�s��ݘk(��+�{Fٹ3�n8���W�$�m��[o��7v�C6﫯���sJ�1ߴ��͹�Rh�{]���g��(��.)�}��~#	��)6G%�Je�t�"��,��P|��B��3pQD^n]�ޠL�~�c��	���qf�홈�j��ttt����z���;L]�}�#'h(t��x�.�D�7 ��_�6f��
kk��٢�!R����;���g����(�+WN��
�.��w�w�;6��6�]bg��̱�ZG�y�9�����>si� ��I�Չ4(��U�H�����L��Ӛe����آ��3ѹTi�#��mszt(�����0L}-�'m\�IBI���L5ˍ	�if�i$EȂ�:#C��9�m��0H1�Y|ư+Pb@]��Φ�,�M9��Z��O������;?��N����紃��S��)e�I��o%�
�I����?����)������}�-��9�E*�%'d<���=��s�`��_6h���׿�=kX��EW�bs��SޚݘD:��;aQ�DK��:�l�Ϊ�([D@7��	���0\���bQ��`͍��`,~��9�p2���n���,�VL��^�G��7�J�q��Eo����;�ݭS �M4P�S2
��nl��;f���Ĕ��I>Q;����E�u.��T���h�mG�}mw���Z4��^��x~�	���$?�����H�~�~T�V��aQ?�3Y)����x2��n���EP�8���'ֳ>�� ��o�"lY������|�Z�u+�M�+!�:u�C��P,)*���z8IndܦZ���� !2lV����0:�������U.�&��d"�#�_I�~}ն̶H*��vg��3¿�r��ꅻ$�0  ��IDATy�YE��i9>��;0�҆�HX�0Ò.������b�NN��Oa*$�0W9�y��}�S�5 �4�ckav_�Ȫ�^ �E�b�+`fpo��pS78s�.�2���L�0&�P&>�{����l<z��½�bƖ����L�R��`���4 y.��,l�_��-Y�
W	��s�2��;?C��e�n߼M\�_E�	��|����}�0�;���<oߺM���8����wܵ�����~t��/��s_?x�t�=|±h,^1��L+����'^�,Iȿ�oV�W�M�fa�V�ư�{���}e+%�4 �QDu���R��F�4�����ϦS ����<?��w޹�~����?�1ӓ�]ݍ�u��Kp|����^t0�~��W�`��G
�Ro�g����+�t���'���fMX������P(���� ��S��2�p����T`��<pa]�'F�SP� qF��꧟~��,����c���#�Vx�zAK[J�����`��D:i�����y�(�|qtH۳���y �z3��XW��JU��tұSH1���Q^��H'��<pa�%U�@��� ��G �҂X�g��lS�q;�M��$6��c��q^RJ�\:���Z�r|����n&�+X�f�oz�e� *f�+7_��og{Y��+�տ��y��\T�{^1`��1['�oGN�7��eeE�!��S�Ӟ�Z1���.�lJ�֭�n�R�7�v�+�{|��>,��SU0*qR8�4,�4��\cn+��x` �FS7�"�D`�ܥN'�I�8�֩gX[A^�4�#t&���J��%��^%�$�6^�J`Y�k����(w֒%B��v>�<_1�Fzkl�U�d�a�p���y`X�P���k�Rf�k�
U�́3F'���(RIe(�˃�x�%�tY-1��k�(�����t^�����V[�
S0���FBٕ
����:uW����<V�]�6�yR/^@ �=Jx��P'#�0��:��`�aHa\���Ë�e�2����Հw����[Ŷ4%pW>~��}���C~Ĵ��o�u'�[�7�ۄ��Ҋ��4��	�`���i����:��m>�1w)���p�T�5-�Cq 7�rb�^0��Ie��u]߹M����w�U�-rk�$��E
C<_\�ݻC\XP�_,�8���Bf�� #^%Kj'c,t(���"=�6�W ��Ǻ�X<���y7o^s��]��獽]wek�)7/^���mP��:`��#�;�U�8�h��"Kh߻�'v~ļ���J����\�:{Q�Y�����´�D���9K+p��bY�sS�,kV�6ɂ袅�3���i��]�Ht���\O�=����+��H�����?d�)Ƒ�d�̀�$��a\')q�ڎ{뭛�p`n��\e��JeΎ����s�"+���뷥�iCɡ7pgl���n�x�t
��K
F �t� J�!c�'O�����w�&�aoo��|��^ۈ_�|v��,�x���3J��F��43��`�vm���Aݼu3:n7�ĸAD��6mV"1`�{$u�߹�,Ih������gn���VL������ij��4Y�v!����ʒ�g	��8v�mD�?&Q�Tӿ�D��L�葐6�B��K���߾]��Ͷor[ے�]��;��������U.�/̛�g���Q��d��f6��L�ә�%Лϸ��dL'�����"��$h�R�&���[��|�\��G�mc���r��
��<��0q��,��<�J(��At=F�t7�~�E$�U���V��Q���Ai^��{�,P�!����̡��Z4h;W��7�r����+7[x�I�Ԑ䚜E��2;"-��C�*@7Q�BA�p�,'�K?��$]y��X\_�.f���u"$�h0 ����-FÓѮ� 5҅K�&��Z+�Q�C	0V��-*d��� �PH��q�@J�!�)l�|_AR�*�H,���J`�� ����~7��^H�5�H[�_3�X�5���l���v������]Ð�
��0�b6=�Dו+g\�����N7u�����OY��j������{��	P�Cv���.����,X������O>��;rm7֯$�=��v]*>*<E�A=�[n3jh�r��:( w��;lg@��cJ3㌂9��5����1���r�P�<�q)M�d�d?�L"���`�T���8����<��I��srsC:9�8N�v�q�w���;2� T��X��X\ /(� �p5���w'^���!��}jOV���l�w��/������N�/B�N��T����*3(iU����o�O-f�-�B蒷�bg
�z���4����"���u�nj)�D��7�3�	���hI����at������O���#�܎��1��e�!V��50�#F9^�}�aj:5�O'���x�ܔ�5i�b�Z�� ��Qy>9*!`��\&��oZ�%l�MD=0�\r.� ���uQ�l�) �8:�8�"r���&�0��Ç�5Ǻ��(���1�����:���g���p"p>��`��xiYh�1���%'��5�&�����2�6�$d���uI�.5=_���L���!��C]�$VLi C���w��7��D�_ 5�2u���z��@�x+�^�����A�ožu��b̽��T��n�������z��f����0vy�+��[(4$8��Uߥ��!I�Hޮh!B~�q���p;T�vq���i;����<� ��A`KB�?�]0�A4Cab�{�ڡZ�,>u��fD��&0�ՐE;:�&! ��V�O2d��Y(C8���Aaښ���f����u[�7�ϫ�n"�O�HRu��=l��şS�=�y�v�4߈��j���=]~1���-��U����)��Jٞ��#� �A-����o6��-m8�����.r�#���3��%MĨ�8K7"q`$�������ѐ�!\h�"����}��dL��{��P�}�#���������EyÛ+�����h�sUh�v�Lu ��0R 	��fXؾ��k�7���kLAhoo;�k���"�k���m��񢺁�̽�5�)>��x� ٹ;=;�u��p6n��kc�k�߻l�q��?q���߸�>���a�X�MH�IY�KC�NZm$ӽ��� �Q���䔌.��~�u��P,&9|C��������� NXТ����'�������v7������0���qn�
�5���~糹�N6,�I]�X^l���&�|����"0eAH�+�3CfZ=I��+�s����Bɶ�"ĀE��e��s����]�;u������嵄�B]��F{B�$��Q忋g�ۨ~RW���!pك�29�=��A�� %:U�������������b"@:�vt|����F�r�*0�)C�F��d9����!}Q~�iJ����UZ����W�~K��O����>>IMT��mA�55�Y�n��3������Tl����;�v��~m����K9�s� ��}z�쿐4���#����N�i�SF�����|N�sU�q)Γ��s6��);�N����u����/�k���j� ��j�����y���K7�&\���.8>��&e��TiX�N����n	�]��7���-2
��nS�-��.�
���t?T���E�7���%[�!�k<�<Nz޿� ���r���b�'�����a�>��6�Ր���~�*��1Z���L���8!p���G~]�+��E0����aai����T�?��G�T0$CsL���M��ǀ#�.�� ��Ո�k�&��6��Bq��uE�9�5�;�R�����,����dr���(�	��v��nta��`l���zo�0'�����{�����6ky�F[�:��'�[�[���}�3�[�9i�� @ra`!P�7��@��ˋC)6�q������i9�G��7X��7�Lɛ�R�������.���u��4���H�.�W�VGw4��sPO@ 
���� _�;�y�L�9Y,�?Q\v������[��E`�q��5���ml�@m6���[A�L��0c?~������?�������ڙj��~�	����a��b��"A*��q|S�@Q!
�����)5�)��z]�.=��2
�2:�#Hix�������^qO�<d^. ?�B���[k]r�c@ �i1��v� 6'c���[x8>�V�.)]:}ɖΥ����Z�F�B�l��)�%�Sm�*+=�n��(�֑���R�[!2Hg��T���dW��� �gfn��{򝐽�S�(-����耠� W�	h�iٌ�C8�d�ݹ���!����S'Ńm|Ώ��T���@5\7����s�ᐚr
6)�hQή����R |.(����Ed	oc|�i7I1�ymҽ�8ҋ �3rj��p~����ѱܼ�p_��O���q�O�N�3J��6����:�L��
Si�t�3F;i�{�:��i:x^�A��U�f��d�)m�ye�k �Fwid�.�{�4�ͭq79��7���Y���N�8>�8o��/�M0E�r���] ��$��w�����R0P�aaHH�-�6��
vƭ܊��e�̙��H�_*H�&��1��[2dN�\۶SY1'9H�F�ܱ�MD��@D�G�7���̹�8���lƉ|�ݸu�`�E4Nd)��&�=lT1f�]s�$��U#!F�I�Á�6L���
��n��������2Z�E�b?�+0�w�\�����Hh0 � m��y_��.��5�����EP��0���ǅ���w`|��G�]NO�
XMi`W�%9��X��.� �9���z��UqH �!F�i�h��TȝP�2�U��	Bb � �`b��.����q�~�]�������3C�����+-nE 
)O��S�i�B/KeX��P2^����8k(��@�����#"�#`���{��Q|�(Ta}�}�.�gg'\�Pp�����<@��ņé�/d�ű��Rc`,�o0[�"d������?d���?��q��}����d��)o���.���$D٥$��/xM���P�G�=�^���=a�:5�X9"�����$'aSG���O��?����|������yF�.�
��$��B#�g"��� ���ئ�͝耫:����i4	��`/+��nYWX����N K�]ŤÔ9wUb")������Vj�=�0˨)��)���R U�LM��?��b��h�6kMP���H%��!^���@����0��}���c�)H�an�8EP` �Sr�'�޽/X���sM $%)+���
[-UI��Yҍ�ָL?�u�*�dtV�\*�6�R�@�Ę7Y9���l˒{������[�|}�Z@z�O���?�x>?���2��>���0���c�i��vI�L��\�f*��U��i����N�ҥ��ŗ��!
Z*�u	�/!�432��u3tD**"1�D5�/��"�XG���.�]����V����1 l��~���\/�ث�O���ElM�|��}ih�X���c��U W��hi=b�c��5ڡ,lO x�6z��V�B��?ѕ�s�;�މ�4zuG���Fp	%��9\`�7���6�?�#���2�kZ���C���V��.3�[��/�j}Q;�j�;O�E)�`#P�2��YL�M�`�{�qqA�ɵ�x���L�ڛ��7�qFo�^e|��(�P������/�O�³�d��'�M��m����#�n�<U��i/�Y���61�zn��S��/X�	�z�5��	�}�-�ӟ�����Ь���� �9+�%���}?��lB�(����@�{p�"-�n����%�[v�v�X�,%`���(��!�P��0)�-��H�����������8�߶q�8Y�'��R#�4?���R(2�v>C^/�8ؼ%@vi��9A5JgԫD�)
�l\QމLP���辎�/>C�dF+�%-�������e���w���;Ho0�@��AÖs{/9�*WT�1�����hlHc��<?#}����,�I84h'������U�p}�m����nkk�̻H.R�'
���NX��?gnh��|A���c�گ�+�ƽtV���WA���(�%	!�l���iN$K^�&��8�l�y��Ϡ�1���E��h{a��hNڗ_~��U�µm�tJPຽ��֟��߇G�Ի�Кz���	��
�a������z����5�
I#��7Y;�4�M� �')�.�����@�������&d�,4��_p=�ϼK��ٸa�2�$H�a�=~�����[q�����׹F��v�����U� -�o�z�9�b$����Q��[�cۥqe���{A��P�[�D��ee�I�(b�/Z�"�'k5���d6�5�8XoIPK�n�ڿ�\�{�����ooo����E��2�b}|.��[©f;�v�-��gĽW�FZOl?������fmdB��8٥E"�u��pq@d�	9��x���@�A�rVwd=�C�噛�F���i`��e���h��h|�]��v�37??"��D�~<�r����G�qZ�f	� �g!���O��5V�!)	"tO5�!�`(0��i���ΚA��u5U������Qk��F@���U-�0��c�V`�"�m�+�Sws~��=v���`2�䊓��Z�`F�j��l�e�c>����|�y5R\�z��1�1޳�I��H���P[�
�������0&�0jN.��h<���������������~\��$L��BfH����p�cmC i� ������?^�E�U�S��a����~V+;�b0���삵}��Կ�|�o�={Bf	:�_����ۨ�7�C��ѐ���6��E��̐��1m�]P^E#ȷ��\�s�\�=<�`�.U���'���E�R�[�߷`<gY8u^sA��z�pV  �| z�}�]��xf�p����w--�@㲧�c-��YJ�-�<B�/�o8�K�J������i��8��qKG�,>������O�;������D�v� g�^|θ���z�<T8(tL�D6�uF:Ґ攱�Mդ{�5`8ʂ�g����=]"RQ���|�<�΢3J�i�_���Ԋ2'�RL��T�(?t�k�P�d5 c�*i����?�#�����U�裟���slH��A�Q��/�C�t�� G�ѱ�;L���5�
��	�}����xV�������~3W�#�N�L�1U�[8�4��j��0
53�-�5���e=kc�ߩaR�XJ]3��0���e��d��� �����H#��0t3C3؆�R�(��J
��A�X�%��-Z[�4rͰ�c�O�;�~��L"!�r�ӂJ�^�S���w�&4��-�8Fa��C�F��z�hׇɜ2�]��@��r��ų,�Ϧ�����<˿�/����+J@1�����6�����)��1�<?uޖ nr��u$�'�{�5F��{ښ;�-�O�Ի��M��G-]}?Q�v}K�Ho�TVƅ��;}�w0�B�= =0v
3������De��"������S �h�Io��)`�F#ZSz�0 k����
�T�޹H*�]@���0����d�Jk�R ����yLʪ�

�h2	植0���Ʈ�uo�I;Eݩ�0�ax��֔x��:sR��/k73�7��dd�֭�;��-=O�6�@X-�l	�ŏ5R�\3D�S5�ڛ~��L:NP!�w�P�,̝�^��r��H�����Jc�A��	:��B���9} O)#.F@]fH�Z���>��)p@�u*Y�ЛUm��9�8�k�(:%�;Uvq6�?4�n�@Su�(��-�(,���'��FҐ����Iק�d��^x"�%���Nqp)�n��3�� [^ �������a �{�Ne��Fݫگ�V���yG |����ۏ��T+�g�0�cRP��`�zz(��Y��ݻ�]�N�����(V����be<d��TbvL�����Yў33N�k���s�dJ9Y�_�ӥ����a!)&�7;V�c^�9��4Vت�͑)�6�CiE�vA��3J�%�e��m�z|�Ȟhs��~�d߽u�3�_|�9��~/V��=#s��6J���	� �ź���>��C3�8���,�},�^S�Y]G�TIr���Q�`�JWye� �ʭo�x���!���s���k��굫��H� ��Ԭi�|�Ӵ\����)/e>6U�\N���h0b��],r�t��ts��X���e������YrF7kYOjm@e9�ؓ�f���d��v��V��rK�]y����� ���ꑑɸ�˟)w��K?��(o��^ZV�K�����]�E�W�� ��'}��ؽ��tͻp�^�鋡�`^�@�ڍq��I=8?9rG�{�ڽ�Ѻ�[��3��z� �VdϮ��v�;c��x����y����6R>$�O�GC7��G#y&	��}Ow���l�&1�!߸VA2{tÆR"ڀr���`l���Ej�˓b����L�g�d��赾���b1��	�<��k����`m`�����a�L� A6��qɃ.@/G�J�	�ꤛ��c��"W��h�VY���ԋ�e���t��!��F,|�/���"��ϣ�H�M��M*N >�ҵ�kԝED���BS���))WUZL�/�y��b���5�G�ύ\]4�� ��������w�{�{�A��gҌ��f�f]K��'$�PX�Bb<3�l:�hǼ&������1�\[ɚ~�g��J5@���r[�']��x!����!���GiÐ�B��r;ޜ��s��}I�ɗ�ʀ���+��Oϴȱa�5y8f,�٘�\�rj��"��>��g��t�T0��7RG���� ~Yd��B����ƕ�%ص�O�4��
��_�U�I+Ÿp� <���6P���rp���g�x~R�d9���E+��(e�K�]�]*�+ǈ��d�q�glmj����Gǻ/>���~H����@�M�NHl ��~>I2��H5$���,���ԝ�[�%� T�򳼕�������sq�@�ԗ�������;�j�Y�8�gQK�ˣ��xl��VJJ�ʪ���@������^�3dsQ'W�x�|m��#' �U1�ծ������Fm�T�zb]Hk��s�f�z�e#.�J��ͽ��{�����$�����ڟ�-���v��}�>/���F�|���X��.IP�U�����4|��\2�χe�p�����t q0�+aF��G0u>u�Gg���I�S7٘G0<v��n�ͭݸ�(�
a���ފ ȍ��>%�]к�}��-A_��v!u���P���u"�Vx��*si�7�_1��t�&�����B�*�fMA��= ��L^H��x�u7G�4�h�D0w�m]���񁛡�5.  &�HB��0[Q��G��i���}�\.<���GQ`f�$st��dOL��U������!���T�������玢&7�;�[���t7Ù1�<[��Z����~��j�k4dwj>�G�����o���;�_�H�]9��#��+ld#�@��R����/���E	�� ��;W���*r2��D��B͆8!��P����PQ���� ^��;�	�4i���op.[̗SA짅z���� �������.�ޓ�����8�[�̂��m��I�i��^0�pЦsg�)��t�J˸�\x��0R�>0⫯ av,`ǋ��p�D�!׺;H.���d`3Eg��ҿ�̹�޽�����l�]�d�;��{����*�i��Vyw��ؐ
�p�x��|P!���]�i��C�%l (���؈�J3��:$6��zɢ��r�s� 1o%������.����bL@���SS��h�5�f��˩R������]�<��j�D4mo��8����x/�)iJT�5���c.m�D���=�u���;,��tz�c���2�B�Z�d����*���A�9?��h�:-^���������
po�;���>�KX��q~����r��n�{�V�l�
m�b���
�	�6}s��T/���^M����[�A��v^���f�Z ƅg�p��$N�S799s�ә�(�x7�gT]��Khf4^w�Wn�� �ڧnr6s�'�5I��$@�&�;�>a�0��X�+ݹ�70G��Wѥ|�d h�S�Ut]`�*���J�9��m��E���$�}8�4��V�#��6��5�nFp���0Nx�nh��z����:��T��[���(���a��k +(�#�ͭT�[ǽE5.�o��g.\�v�w�i����I��n+RX� �0�>gs����o�^���{�����{�؝񜐲�81������W������{��f�R�=�%�1�c�9�ӳ6���ڜBD�@�U���&��[4�(¤V,�*�ʾ����/F�3���5��خȕz��e�ղ���q3p@��4����d�q/�����`���r����2RV�M�7t	��WK���di����z  W,����=:}��3��h�m�s�&E�a��+�r�2�سHK��0�Um�-$5� (�ȫ��p҃Z&e�M��0`{a���ϩ.d����Գ��9m����@�+9�ǳ����b�m���t�&!���2i2 VAzU'�c3z����=M���pN�n�m� ^��s1v0N�y�)/�ϲ��Rzl_��z��s$�'*k��� h��!U:[�;u��!͓4TCH�;�sa��M���#2��x���8W�56�Oh�(�%����ӡ[��g�}�`������/־t]����o:E�j@�'�"7�V|���5����R�ٍ������n1&�˰���Y��7��o�忼t�� ӓM�+I� 1�/���,.�g����`�d�J�E���x�mn_e��8M���C:@׍%|;�v�;m4\�Ttл��_� ̱�l@��2��3L�9�5ٝJ=������Jh�ZUge �:�m�B�TCŀ1�!�;��+�ϝ�����M�����#���_�'�8��x?�����������	�6�jF�䶐#���rb���tƪ���x���;a�[���S_�=��nk���3d[Ⓛ�I!�i��BG\�[5�XL DR�`1��@ӌFF�" ڎ�5Ů!c���/�bqد~�6���{΅g�x
�~{V�@L-���>APHo)�}|tHM]�ĐmLGʺ�n-N�Z�Z�0�lL$gX�Ш#�*ʞ�'	`6Y%˹[fY����
���2h�����dˤ��2j��T�`77��������_t�Z%W^��Vi!NWta��ΛE����.+խ�si1��qE~�2���TƄ]��]���U�۔$�\YO��\by�`p�iD��Js,t%8��k��v?����zύ��nV�	 1-�p��8/�j�]�Ҳ|c�9o^��DV�R-r��T-_/ra�^hP;U$0��RU0L�W�M{om��NX��{1S�u8ȅb�<)��*Ǖ����������-4��"*%���MR�^��C���OuA$16��"��L��|j�-ۥI�:�M�KWj��[�9;)��u>�t>Y*S��Y�hS^9��+NZ�Ǔ�La�	��b}.sӊue�z%L\jU��RN"{�����W�e�zŘ�Mz�-���Ζ_���6'^��E���<Âj$,��慵�'��v����������
J#���K� �a���.X���GM2�֝O ��oު,��{�d/���݁��N�� 9Y�c���!& 
R�<ښ�������n1�0	|�=G `�p�>�"����(,�ø+�5	�ž�#�G�Ճ���R��n�ń}܏^<uOq�����Z��E����z�1T('�)Y[Kќ�e�V�53�X���_A&y�����L�>Wg�Ub�����\f�������M���]�J�w�*-��T8ݎk@l>�kH�)����B����o�~��Pt� Fм؅���_1��H)En�����1�o����w����l�����U�a�n:S�o����/;��n�mt!2�~�U� Q.<�q��O���r3��K��EOQ
����0 ۆ���P`�!݆g���^0��ί
=�фo���<,oѻ�j-�2�?oln1'�`��MZqd��w�1�u�ҍ��_XvQ�h]��d�C"�� laa��M�pyE1�+���0+���.��v������\te�������7�?�r��9Y������{b,6�łm�+������\b��9h�N�&��;M�f{�ۗ}���`]�0�� �kΩ���}^�
\b�\�Y�[Rؚ��l[��'���oLZ�:��e����M܄�G�RZ`]e%j�{�n�R�zg>ih���D���A<�!����B�����qlR������HζEk�>�q���}c�v�_V`���k�zї���ϧb_,֎�]u�a����|�V���/�*�⚲Ù�D�泌uyMj,���賞H(&��z6�C���t�<'ƽ蛼dfu��� ] ��«�k�q�D�3�߰`׬΄`�����o���|�ӧd�7����z��#�+@r�Ag6t7s*6Ͱr��D���-|Gn6��6�Y�հ�ɩ�#�YW���*�ɫ��6L��S�Aؒ� ���6� �eG2��]t�PKh�����=w���=~�,.�x-�kkn7��80Fa3�����,HK-��ji�!���`�|��+�kyb.c7:�q.����?�"�*������:��T�$��&`����''a�.��U�Tx΢���[0hX���n\��~�������������LOݳ���o~�[��?��2d�{���;�m��rĂ�f ��P�9��f:�.�z81<��1W
�:V�{����.
��N�EG�"N�%{���y�"hL�1�����[	�|96�hˋ�-R���"*

�):��9�ギsH[��_��W�b�`��H�\��2>��fݥ�r-�� Y��*��|����
tC�6��ҹHHg�L�AG� g ��ɍ<P6W�[aW�rM,��k_\���W@ו�����Y��-M�T��g�"k!{��`���N���ɫ��NY�W�\�9�d��ԙ>�����(�j���Y
��q�!����缫Djl>�4�Bn��gZ[�u�W�p�0
�	�~�4+\��6A�GӖƳ�=�8ŵ���9���<����})͡Lu(u{WoK,\0�jkw�6�_�	0�Stl�t,�6�й����'�����S�>��s�,2�@vu-���R*ħ4�[�u�
Xk�
S]��-b@�K%���y+�\vo%�ڛo��@�Y}�VF*WݧKy���_�y=��El������D�1��+�6؆Л�T Ӣ�BX������|yO�Sj[?�!���q����&��e{Y�uAe�:(����ǻ�v8Be�d6�5� U�'�}�lD���[w�xCd�Ҁ�>6vNkD����R[��[�왯M�O�]	q������j�-�[�F)p��V�1���dv�47�(�ǐ��h@�q�VO"�=<x���|�ɾ�zL�@���>~�d^7�ƴ^�醒Y5Z�`^��Y�$�X$4-l���L��]f<���Y�y� sΜ����gZCd���-j�Pc���kbW���Ѩk�Y%<��Ww�����ݻ|ݺu;�|;���<z�����s��٧�S�~�`�����jt��v����0�[p1������dL��#�{F��	� 4��R�]23����;N�F��i��d�u��6c�Y!��ۊ�r�4�1'��W��0Ν[Zҋ�e�l5�30h4�!t)����g�5�{K�]+ M��"�����1��tz����XX�N�5ƣK�k�[Y���}�� �[--Q�K
LvJ�*��8g�g>9����5j����r�i�Ӝ��=����Ϧ8�L�H�-�3C�1�Ǎ�-�����|Ͳ}�9L��Mk�
�-U��xW����:�?`�a�Z���A������1�Fz6K)"�+[�qU���,�e]0����yg��e[�Ɖu*�b]ɖ;�������4�V5�i��il�{_���z�j�碅f��Y���}W�M�U�(@^��䖩�;�Wl,Z�v(o��ߑ��2���%�<�p����
]>�v��z)}A�+v���fom9���>i?#[>Ыs���*��z�\���n�˶��2�X4`��h`�����<99��Q�$����4����h7�Qɽ��K8����w恚'��N��m�I�u��G>/��xt� �B *��X��Zz��;Hy ؋�7D
��&[�ԣu0r�)����v��'��_=vώ���\Y����h�v!a�"��;zĭ(���ӂ���� ��v���mEΪ/~��A(?����R��Д}>�������Jb����������tdto޺�~���'}�>��w����B��/�r��忺��_F����HE�q�Ѧ������o<7ѐ7%q/���pb�L�Cm-���b��r/}EkLc^3����f��Qe�[$����)�¬)�1eƘZ���=���G�N^��ٌ@d� ^��/��7/�KVP(�`g���05^
�I�	��]b�:�]�&ۗ�e��H�w+-�)s&?!m���`b�K��у˩,���Uh[2�-_z$�_^C��B�)�mO���{�����vJ��ⶴ�4a��G�:u�#<C7Υ��Ki�����Jl,���hC��<�C�s���q\S�$�(<97�0����0�9	�>#ŵ2F ���c>�.�F:4L��uY��\�=��幝��lw�i�<�V>�`�����Bgx�Ȗ*q�~i>t�SYl�xW4�����c�vY�֧Y���ۅ:�T�1�.���q3[.�a9�����1�Ox�*���'�ui^� �����l��-^Y������͎R �7>9�;�C����l��K�)���1	����s	5{h&���������S���?��v�e�j����L ��^M=���:_`^m"U�Ʀ=Yh��4
@�,s�Z�o���<[�˓��bW��`Bcڷ,âUC�ڑ�����;x��=���ɣ�n����ӊ	�]��Ǯ����^�����3�f9��%�2�MrhO2t*�ǃ+Yް"��/y�GG��Z� Y� zȕ��zz��� [���(��6��-�l8����:s������s?��G����'�{���'�a1��}cAĂr��5w��MW�0���S���X�-�?��C�[����d,���9�D<�?c��E�*?��а���F���z��S���/e�� �d}bzq��l��`ad����o�M���Z�+PP�c�6:���	�B�|���hq�ln.�j�qf�r�酲z3�98�2/�$�׵S����n/�(�w���U����9��c���������-�y�+���v�r-{�Uzo[����@��%�uX���gK�=��Mj���4��C��z%B�l���;�<qk�^3��ٜhL����
;筍�nsc˝���Ǳ�,1.�F	2�{���(���5KS��C��u�	�ki\V8g�	o���!����G,.F9��4P������
|������]���)Z�׍RyE�HΎ���T/��5mNI����i�e7�t!���K@Ilk���.���)���Jq��4����7�0�|s�1�� ��M�+	�oq��˅����x",���^����^�koK�V�cޗtG��$$8��>��ֻE'��� ��.m������=�O����n0����ؖ6�]
�{ʇE0��4#�Q���\��Vc�(O�\��Is�r �u�jx	(a�T���U�����(FЩ;9z���=r�<p����~LF},��uDW��M�&���f��������ȡ����ߒm�g�)�KC�:,�Hf�tf���p	��Y�
L��}�X��uA���|i��sQ��{�>)�g�hQvl!�M�ކ���͛�g?����/~�~������FD�T&)$� ��y��-X��
��m���>>}��=��s��ԡ�|������V�	�w��e4
ój[^Z$-��1�_UA��z��b��~�.
"Mު�}I �5 k�[ /mb�K���l��C*�J��y�-I�����S�,�l�����?#�b@�e�ᬐ��4WhZ��k=s�u.��J���AuaW��Թ,1�9Ձz��s�b9}ή:� d�W�DV�U3�s������3��K9�7K��� H���ْ�wa667��Pu�ʪ����n��4�kHP�n�?Э�	����=�L��sw��_D��@�c���:D�4	0%�N��kM�@@"������R�n�k���8&�Z�v��{S���Q�p+�Cz�Kv�����+FΟN��ؒ�L��[�ךo�cб���[�l� zװ�S�*9~	�⻵�6�����7�?�}���$�r^qY���Uz��2j���鵷dt���Qy��7����WȯK�����>o�(#�� ��,M�9[:F[�@r����r<]*̙	�5Y�(��a1>���+[n}s���O��zC�����]�F���~��&�aI7�7���*��ݪ!.��mE�TB�b��L$�	"�]|�ӧ�܃�HË�;=����	)���������b���l��xI5�=x�x՗Β�YS:[ؤ�?��ŧk"o�B��lħ5�^��⳦���3��5��B��c*��t=����������_�s�w�~����k���E3>�����k�����</,dPr@���"н��=�/��K*7���_��+�����\�os��s��s9|o�f���݅s�a@58K��S���D�ț���i{�{��R�
�8a[j� 8 6P,��R�/�Mi�|�Z�8��~�љB��{�?����w�O���=���{��!��3:�V{�Z
�\�q7o�`�V0�p��՗_SB-kM?� ̺�Y���cV���]~�,z�����i��ؾBE���U9�\�+8����l`Y��ں����E���ȅR�ظ�)��EK�B���5#>wDz�޽�g���͢U�o\���1��������q�yml����;�� �����ܸ¡ f��8������[������y����߈v��v5��]Ke�kQ��/J��8�����X3�h�$��\_��g$y�`���HY���X�D����2���A ����p���ɽ��˵���Ԗ�/��R�B���D,xYGE'�K��ՃF�LPh���ɂm��bZKKp	�ȹ��o�ي|�i{o�U_����f�%=Sg�5����w�tq-
�/�?�c��[94󹔎����y��Z�
�܄%)�l���P�䰆_��om�Z��Pyw�U���>W�7��	p����k��@���N�C�y����#o�
��B��b6. �`%^����B�l8����� @�����8��� ��z*�y\H$T� �?������5�:oښ�ษ;?=r{ �_=rD�u�X�F�m'y�-�d4�5�&�������&�  �klX�'����V�pbM������EWC���%ec@��A�S�	��:5~��ż�`�Z;+���e�^%�ۆC2�`_F�y�M'���#R���J�m[ѳޫ6$W�ǜ����ܹ�v�_�y�9���Tc���с�ɓ�no�Y��y?q<t"asY1ߥS+1'�a�쾘 �Bo�m�#�A��I�¥��v��)SY���f�R0�Ǘ�o.&������n/G��l�
�=�!�|��=\�m�����NMI���`�Φ�`l��,��W8iAZ��i���Y�	>�����w��� Ӎ����H������MqН���gt� �NN���&A6��~���3�p��M���l�?z��F@����K���]��b_���E,C����{k�2��������8W0��i��\YX�gev�*Xf�*uԺ%F%yY^fP�(pٛs��G�����b��v���E���F���[�ng�*�Z8��{��[������v����o�u�y�;ц\e�tѽB��ï�q�;;kѾ4���k�������2J���E冎�W�XY.��]�'Yg�K�F�H.�\�[E�Z@�|.�>S�i������׋N�n c��3U
�K6�kmȁȘu5��7y52�T��� �;OVj��祽R!�35�Z���p6��ƅ<_�3E��Pep�9Ys'��z���2hͬe��4�^�U/�t��s]����^d��G~3З��˜=�������RQH�g:s@��Ɩ��]�_���������/I��h.�!�1��l�v
��.��kyBޥNZ,�J��&�#_��p�W�9���*�.���-��Y ��郂a�P�U8�s �����=��8����fU���p��si�L��0@��[�`7�F
R�B�'���:��(��Ι�@��o�h����(.��?r_��={�".��x���}(m/;��m�C�C^^3r]u�hd����AZ��TT�6�kg��,�ViE��U�ƹ��.?5|�V��$�d�J^�פu��������&�V��OƓ�=���./�͠I�ox��ղwI��*�����L9��Z����a\��NB�u��[��)�s����sH��M�4�lR��M�X.�A�%�5+�ixe��J��\��:����a�H��*�Y���)ɘ'x�jÂJ�E:J�4�O#@�L�$oYs!��n�B�K���B�K��d/,,!{�e���N,	G��wo�&�u$�zD�Z
UXI�+���(��Wi�������+���7O=�D���$v��-��3���ODfe��ݷ�N��Z2###�bnnn�@�w�SV2�\���TĶ�d�.Ջ���g�?E�t�? ���z�˯~�+�裟ǿ��d����=y���������g�E������u�y�������?�����@�h����W_~ŢJg��Erp���^�p�Ke��	�ėYQd.!9Pva��C>�pL�^�y^�ڸN��PХ�38��,Q̋5cؗo.�������mi,��>[��և��	
�)�~}[~�������c0ܢ�'�vw���M���2���%��ߏAȇ~(k�[,rVY5$S-�|gE޿�Љ��T��_��r5���1�ٌ���}�Ac��!������p� ���x2F����x���T������0�O�d����;\��Y"���:NN�3� ���dV����^�f���u��==v���,�\�/B�î�]\̽�2��x������gJ�M�΀`��b�,��_�-$�=�D+)1d�3���b�>�� 9����p��V[o����j�ty���{[�7')~��E���oM��-������^4��'�\b��-�']�����q[U�P?߲#Ċl擁��{��G�C[h�s�߇���)�V�l���=������{F5h��z)QHլ��"�BvVP0\ �����������ӈ�S��Ng�Jm��Ą -2X�ͤ�L�	�m 9�8�f��v�`��8yOdp�Kǀ����1
���{9~�/�d(s����rT���yḂ�%w�7��C���t3���1�����4�
���آ?o�z]]��5|���M]���3
nSW&���k�a���;�?���'��zU��.���0��d!��yS���n+��y$ݿ_���O�ٳ�,l ������y��q�R�k!f/fK�O'�W�������h:ԣ���tR�� �d0x��m1�� ����9U`����%�i|�T���,�O�M���XYj� )E���F����{�{��'��tcv
l�~o����~��S�Ht�u�Wv!����0��{dg7/mj����ا`���]���-O Q��Mc0u����S�ܼ��8�������+r��5f+ ��7.�|�0����x�oH�ei<,2��$��Eҙ�<��2��͹#�ūu��1���:?�V�n��Ty�5���s�TU�r� i���E����<SG��z\s�\������`7��F�������#��r�Aw�"���G���ϔm�?�a<�ݻ���V�40;fa�� Xu,�5j�S�_�g<ߋ�|�s��T�3�:t��uYs��,�r�R\n�kt�|���%��jc%Zv��$!���E\*1s�i.�F%���y5�e�=tM�yU��u�e�I/���@}/9���'>���L���%��	�k��4�u����`�Ǳ|`�L��{q-���٤W��_]�p-�M�0���AT�����l������礯3��g~%��שq��G��҃K�kxSt��A�Nޟ*j ^��}�OLoe������J ^8$�ƥ���t!�V#���p"k�@i�ƈjx�D]Y�/n��x�0W�K:(#c�v�yE�kt���nU�"�*�AhN�I�	ֶ�sŨuD6�p�@�>ّ�����UW�V?'F#AS�
xc��+S��j��Pq�N^\��<E9��%AN
~L[:@�� ��XR.`�v��(ɘ�)� h�Aެ	te��6��m�l1T�@�Ņ��hZqzr&< h��0j��f�P�������KA���2}�{lQ������79�1��"�^�����P����M#+��r^G� ����K���&^��`E�4�w$#l���3�ٵ��5�FQ���R��=�:h���i���g��}��� �~u.�C]�����3�
_denU��jyj8K��y=u�v'�2���#�\�.xi�������P���;�)���hk�R�z68����Г�E� 8Y��jEp)uv�:��k}D]7�,n�ZĴ����U2�lՎ
��0�)in4��qKGܿ�6�	j��e���>f=8��v.�zqf�NW)��N��%�!h�������^�� �����?$l��U��@�?�Pk�cH���.n������͓�$Η�7��q��[I�O�������l��< �.?�Oz��P��a8�˝�Zho[M�&�萑!�v�znk�aA�@������pL����de5w������y洎I�E��8�_�u�E�8�g�3v8=>9a[vF��A'��%Cp1"0w�5�䃜B]F��O�`qY�M_�)0� ��?�3ѐ��='��.�'��3��}D�qJ�$����Ҥ �Ŝ��1���=º�D�D�iS}��p�������ME:�_���D�G]��
�f�^p>����T�Kߋ ��:���t�&���Si�.i�8aFqBL�C�E��G�޶�D�������F��&����Y�noCo����o�(�9)�/�Os]�hfl~��ti���a��2KdQ��Ц(nv��#j��Nd�p Gh��z�%
�e����>�1�H�dn�⊔R�tߌ�r�cT8��F�5���4~��P-X���ԡ�Msw	��2��^g�4e���x�*�+˫��ڦ�ѩB��NOO�xԚCgKj&T�TZ�sfDG���� v������<�x���d���.��I�2I_��v���A����m���~�my��7���_'3�J��X��Ya���u��5��CQ@��U��c ^��I��C�Cy��1�*� �>� bi������y�Y?�<��P)���<�n�Lܜ��"7���酓Ħ�>���yEx��૯���B���k�����x����_��q���[@��,���vUY����`��"H��+�A8��s��LX�,sb�YU����~0����J��J�*2�8/쓛S@��9���k�5`�zZ�o40[<-�l'9����Ij[y ��p�e>ækQ���\�(��k} ���&]X��'h�>�5u��T��oWW�Y�6�L���D@9�k���ů}ɯ^��+m���m�������CvF�Y��,5bpY
�#��d���m�*������%4��l���^�9��I_��߸�!��8��\��E��*"���������O�����7�׎�^��խk��ͫ���Z����A.� X>|@'4~B`
?���3�C8x��"9]��sҎ�u6g2���*���dv�D�8�A�l�N�/_b��J����׮ɥ�M^�ʈ��F���q�"F(�j~<:��u�gIL��&�߳O9�4,�7q��_����v�����_<��ei�<��&��i@�O����ys��m}�O"k�(]�Ɖ�C��O;[��K#����ᭌ���3��z��
ծ���@���^���,b�jd]�r�<:��S��ƿ��%vs�5׬�z�jm\�xp�x�
BO������R]/�R����ef��C2���	(f��o!���6�HӐ�ដ��vəW���{��H�^��X�H�& M��X67X9̫6Sf�M׊L�lՔ������Vo�L5n��z�&�X;c3}��� z�:��r�lmm�w������ԡ'O��B��4�@k/.�ش����c�N��5��k��Zſ#=^��E����#��߲�7Y8u���]xW֘)>���"�Ҫ��s���X0d�[P�<1/X ^	7�<��-�X[�������q����
��� d/�t����}�r�u�k`A���Fv,o�@-����\x��cw���~R�
�s�1����c0t$� �=���I�蠅�30����c��Xt���G��n%�>�j�,�E � ���Tfo� Q�e�%��즱�<1���-xG��?��3�΄c�̬�]���}�o�ō@U�"���0wZ����Gb�t�̷Ξ���5H�e�4�v�V��Ո���M^gd3v����|��~|^/ν[�t��?}"q-����5��g�C_[Q*�I�.�t�3��d֯���L-���67.ǹ��ܸy�#?z��.��(����3����.�kN���}Yn�z�2�ed������n�{�{��=�ME��g���*�D��ɯ>��?�����;����#4ψ�9����b,�VL���z=M	���	΃M\��x\�2�>ٽv����!8�J`����*7�k�1m��W�ѣG�#�������#�8�N�39�qe� ���qO
���s�ÚH���P$Z6�o_kչu���1�~�������<�������z�r���~�i��y����M �	N�}]v۳ƿŇK����������Ԩ,M `�Z��vec}5Fuq㆟s�o��K]
�2��O]l�c��4�p3��Ej�-�u��}�I���F&I���iAV�oe��S=U��n7�1Rh��<i#�Ƃ1����Env�����%Y� ��rT���a���k�*���/k�S*4����o"~�ҫ&K`E�>@zjLa?U/c�c��݊�����Ssvةwq���7��p��m���~'�߹��^#k�Z�i�mV;�D�lXx�������z�Q\ #>i����L��:���N�7��u�vr��ڛ��u��|��qÁ����V�ب�L u�r�׳jU0ؖ$�I6^�������40	`����M�'�ܹCۧ��1�)r�N�J\��0mjO�U�����=�&{�b�n*vap�.Uf=�ʔ�t�����2��t}�y�;q~��S�-�P={��@�l�����Ȭ�BO��	L,Ɛ��!qݮ]+������˪�&��� �{rrDg��5!���\��6����>����y�vm�M��2�NM�]e�[�QF���[7�`�~��1�U3�u�˧e�()4��^j>�M��~�e��˙^��I\/�n>����_�[����}���ep��>����"ۇ�!����� ���.��|R���v�e6��s�T���#3����>
@ߔ޻#~��o~�k����y���h���?�����Y�1�y����⋵L��L~����?����u��om�����ޖO?��|��W�����JecŲ_$L2dS����o�o��_�����}'w��F���[u=�u�:J�GؿJ^o0�E��'��0�(���o���Zbz����zδ���:��a<> ��)drtX���Ž{z���!�c2ޛ�k��q|�	dXS6Y���cZ����ZΎ� �#8~�Ɩ\�Z��7.�3밾�in��߳
����"����GH��ן�����9�_�SM6]t����!HHR���ī��,e�Z�/Ғ�lOB�U5#Ҍ{B:��?~���m��Sy5�L�d"7�P�� �ZiG@0�\� �'*�˂)�T�'[?N���U�EPM��u�Di+��<
] @�$�<4'd���&(����7�@g�jb�{0���gZ@��Mg��-�
N��R����)"�ю��ʌ@wz:M:���9M���vg�?E�߿"k�,H p�Vn�6-q��3����7�s�h~��!s~p�dC#�`ǜ��<���
Y0�����I�i��$j�DP��ndp�1��X����Ϗ>�H~����k��V[��J�V�H� 6m�p}إ�@����"�͝�)���i�s��O���Y���9�s���H�c�"� ���-|��Yn�~O�~�6kx{B��s��q`���a��3g�ԇ�L�rU�a���j#��ڑ,]n�(6lwR;T�C�a��R/����z�(p���>ì�4���{����L�:f��#��
ӯ��R���^�	v�5S��>�a~��g`��h�:R���5�, (��W ă��%U��-y�X�����n�Im(��餒�O�Yơ���GK2��aIƪ��4�5����eu�,�)��*�4 qV��k9G0����*	`J�F2𥹧H����>�7�yv��H��O��(�{�֨&{[�^},jq,^z�,���!��J��?{�OA�B�b�B�Nǲ�l?^�]ٍ��� ��b�4�ʉ2s�`�F��L��,������7w��\pro�cC�e�Q?\�0.&�^�(j7��y띷�_}��]�q�����	��ԑ�orMG�]-�(
w��t�}R�O~�1�H�*��lUK��+je˸G"���tK>�����o���e�m�(��ȝ��R{녣��J|M��7p_�38��׃%t�*̝����͕������Y�ȅ�H,�P�};2��~{GA����zQ�7��HF��}rR��cpf�Axi����H�~d}5^�x�#�u��9ȶ���8�-dZ�R/��'�����;n��]r��KN�^����̈�DRd�\Bu�o��/�xC��.���WMn��W�q��IZ/la��VH��?z+=�y��Bolj'�_���WE�N6�SR�y���m�ti�գl	���h�U	��fڈ���0��k�F�vQS(�n��.�xYEa�?x�Ũ���}�2�#������2!��sQ���d<��p��xLP.&��4ͬ�#W�oQ�D�>��ũ��@�2���U���+�\JsS�4M��qz� �Wj�m���Z�K��� n�Q�	�^8~��6�	�x`S�u��Q�;��jl�u���� n3I֠�L�1�2[�0�{QŬzZlԁb,�h#��{�ɛo�A�L�o�O�t	�[&���y�w�Ń�"���N�N����al�u������֖����4��A|	Eh�/q���~��w䗟|,�����k��T�Zf��rl���" 1	Kf]U�z��^��^�Ƽ��� '���5n�������{���qqlv#���9P�XA1ͦ��pijm��S���.YP]iE�%�yÃAҥ�)��7�u0OYG���+-���o@X:dh��ƈth�ng�wGɯX5�j�Ǣ�x�E�-��	�=��,���Ǫ���@�+��/����}��uH�O�n��?�?�]�f1$�(-�r��u[`O/�Ou )҆�������U=�g�����n��4Uu�Ze&cU�g�Fa���m��v����تw���F(��{Q���S�ݍ�5�1�ηn���4?z�L��{"��� �im[<:�%������,�h����8�Վ���/v�z���g<Rͮ^�Jp@������������"��W�;��_�u}gC�8O�.�g(ܪX�u�<���P.Ǡw=y `��{��_�����]j���ҕ+[[�Q|�{�ߑkW���tE��
�&r�t)]��h�ڸ}���¼�32�8_��r/�R�0�][�ϸ����Ś�b74�K������y�����J����Zr}��=�A>��vSk�=����#9>�}y�Zi�w��B3%?����^�
z�x�.Q��}��K��/<��6Y�&���]�G{9Y�}$�v�Z���^��ɋ�j��Ջx�Y��=������"s�S=�R`F���L�Ib���97�^N ��Ί���a����Htz�݅�*��B8�Ktc��bx*�1<x�R�E����P����HC���hȴ&*ddv��q"ce��p������L[!��*Y�~� ���5b%�ؕ �=%JT��&�>tZɶJr�T���I�<Ε2�
�W7¼�`����i��~�����!b�߬BK䒝�����*���R�rc�������+z7�����.��M��Y`
xB+�� ���w�� ��l �v㊛�_�6. [[�r�z�me�G�˸�H��a�u����n��m�m��)�}�
`w�|����d P�+��]:�P���4��a�8�۵-,ʄ�3Q���H�C&��5���&�c-�V�U2����%�1�W���o�gf�R�}fۊ>x;O��=u��P_�y��k<�f����x�?E���=H#����p���.��@8��u%���z5�Ǧ��y4�
fM2q�g�q�B3�R��sL�m����{�w�,��N�0�M�0� z�i�����xl`�UG��i�����+�4-��5j�_�O=]w�k�4s��2�כ=7��� �*�=.�]��� ��3/t�����O�ۆ{�,<�wJu�y�x/γ��H|<�_G����}<S_q�o�Yx��V3 I��R3��'hg�s�4���{94��Wk��?��|�|�ݏ�����a� ����B�H�Jk[��3�� �Z?{�L�����>�w�y�kѭ������|����tA�|�H�1W����-9�kP����"Ѕ�s��w�M���F��.s-���q���>������-�.�(*3�`r��${�R�@:ᚮ��0����W�����c�A�U	�~�Sй�Ţpw�a1]<����/�WM����:��޵��	Z�c됯	/?H����䅳�I���8�Ⱦܻ�Dfz���_���y=�^�
5����N�G��}��̶�/�4Z!,Sgv�姟F�O~mt��vMg8
�5�GJ����;�J�4q��+�Q��.ܒ	m�N�L�t������S�:���X�<Xcv5b�'m�
�Oha�>~%�.�.���6'�bJK�M	�gX�G���~LaUz	��U���!�7N�^����t�қ+�˭�[�X�ھ\k����/ʍ������/�"뤀�FF�6��⽚�#ɫ���J�[��ɦ���m�m0�^�BP��"|�,& �lKˬ2��&���������.qP"TeЫ^�~#�kɺ	H�� ݰ|��ӱ��{,Z^́�L��(�06JYB�e�\�EԷ�zS�z��x.WiI���
`��[S�ϩf�p���)) 3lȕ7������XYU�i؞� ��̾Ϲq�j��X��7ޤn�B� h*����K���xq_]67�ER��k�G����b�3�7���{\�	9&�V2�ճ�EN;{i�m�|l��p��kqQ�vj�
��M6����^��,��� q���x�HM#E͹��?X�҂`�Wނ���J�Z�f�d�+ck�*1������b#�R�$RșȍԻ5��S+���-hQ-qK���X\���L�� ��>�<����B�l�5sasV��D�NNɔ����B;�q�։��������e�2�Z���&��u���F��צ8m���1>�6‷�a��UɌ�d�s�-�u�5��X,�w(_}����/_�չ������t{�L��r����.�Z٧� +��''gꤐ��Bjc����u���G���G����>�1�Ŷ�\J�����{
�
�I�Gaϥ�i�Y��R�!��f�b[�8�k�~�=�d�Wj�J�$��0\;g�xm�}�A�ђ�X�z�c��I��d��V:3L���.���*I'�W)�2�$��L?s�-ބO�4���������>�-czn��S���L�//>�l�ﶍ'7"ɋ������w��O��c9���7H��K�+C�	����s.�Xx�y��]�]?��ٱ�I�)���ru�`�t��'�A/<u��eSX���#Ȣ��4= Ю�)3vvv�P\�*JZcMQ!b��4�n����L9V�٪P]�(�F�J7>�}���&�l=���9=>��6�Zw2c�gd�����H�!�Hg�4���"5���L��)�T��RN&ݝ��m�����m~1Ә�!�Nn8zly��Np�]����ηܢȺ?e���0�*c#��l��:�=� ��e�&H��v������|IЖZr�?�Q-o+nW"0>���l���Q�ꫯ8ml���II�z5XD+�>�h�V�����P��TX����j���T+�`��	r	zCɔ;�شqĘ���`�6	�:k��ݻ��N�u���>�L�aC�}��E�Z�l˫�ݒ7n���s�=�e_GgB�$ ��A���|�܁h;m�ھT,U��`6��L���`3~�hỻC�06]VZ�6�Ow�:Ba^�Ӗe5���}:��m�G.�R=ys�f�zR�뵙B�Կځ1��5Oڃ����7g	}��Z���ԍliM�%�e9��~.z����Z	���lN�ˡ��3�[����l���Y勺���D�n��$h>�"$}��/��2�gIc-�������6$
g�3z�B:r$�*���W��*�(��;��3�?��I]���fL:�Y�$T8Pfc]ռ�����Ay�u�\��/���o��pƚ���ww�F�����o�{�|���p�@�D�C������ؐ}��W��{��=0>��������>��N#�����:������@��s���'t���
���6�8����df�z��7���xhҕY5�JZ�5�!F,���+
����W�~�m�'W�k��qNg��}����wuM;����2�q�G�AP���hO֍{f5+�,~�,�+���Gw��r���}^�Cp���|�Km�M�6�X�gZG	ϙ$�y&��xw�iZS��=��HZ����j|��ח}�nW�'|�:�5��T�� ���pgu3��Ӥ3-l_���H�jF	Kه���$Qts/h���8�T3.B�'nt��mi��2���ʛ�E�TN���p`X�������d`g��i���f�?�N<�₣t4�GJ�]�r����ϖl��:�c����ɐ�����
[��O������jI�la$��D��C��h���3m���]gw\x�~b������&���Ws�/GKn\=Q�����C�E{$�4���*co��77�v��$�#�H�'�}!�.^O��	�pYv��߻wO~��O	z����:������*~F7�M�1�
�ploM�L�6]�~���8C��[��8"݇��	�� �`�`��9~Y��L�L�,J�{����v�\�7�����\ c��DK���V���(��uR�|��1p؎����f� �Y|~�M�����ηwjoљ9d�fࠦ.�T�b~�Ha�T��'��p p�-��
���[�nQ������Y���,>y�D>�����?���)��Vf��?6W�>֌#>g撞�66g���.Yц2��e-\�@.2�x!Un�����ϛ�A�~�>ˌE\�H X/�ձNS�	�Ȳ4��53K��2��-���</ �P�e�$�k�s��u�lh� ��Δ���e�4���iʩD�o�֖f���z�
�/�����(�7��jK�<K�,�?���L7�\� B�L�k(u�Q�=���1��8ۙZ[�"c�d�׭Yc79�xa��V�`e��œ'O���?gCh���l��F��Z���-}�ʻ�qx9�%a:���������?8����h�e��?%��������L��d}sU�{�x�=f�P�����b��L�o�� 5BͲ���f� )���Z��T��єqQ�
�L�}��}�ZIm<3�!���O��tX�_|Fدq��Kľ�9��Tw�o=���r���Q���P���p�aͬ�?�����W[.k<�9Dq��Ӂ��Ɉ�i��9�_|��_��^u֕�A��Z���	>�����Zduj�϶Tm�5�dBEi`���:���F6W�2���[��u�=/"�vIw�.���i*U�h39��B;;����ͅ�7)|V j���"^��bC�� ��aB	�pp���e�ߗ�d�/��
�k�\+\��ѥ��S1�6����$��^Iƨo��q�B�'E��J+6��Eݮ�o H�]�������X[��\D������Y��4"i8`������ՀWĵ������:Gx���1yvJ=����{Q�ݱ>��SyA@%�O���T���n���w�^y�U�y�&��.����}J����y�W?T)}�ޕ
�PѬO�d*G�[��ݠ�f�O�
9��D�(�}�(~N|=f���
��r��Z �s[%Zz65p ��~α��u��1�H1�r���W�k�L-�C��t޸q�-Ή��*���̠{\;s1+�ϕ 4�3���
`����^�~]��o�V>����Ï(;���Z�����.;�=z<$�	},�.�1Ƽ�FC�'��'(�-�Z�n��x�ru& �N+'�lם��>t�b�+40�B�E�ݲy�Y!�Pf��E�*\D]d�,���yc�n�x�!��)�`v�:ݵ��P4��B/������hx;�i̖���s@ఝ)c�q��q7���z��H@�)��1Z�b���Z���e�
�����d2Һ�H�h��)�,�3���Y��X�]��§�����L���@�뭿MלK�>����.�2�� �X�q��8�����3�S�g2�=��8G��7Xǀ��O����f#�	�:�:���+j|Y3��Θ�(%�C\��;�2������ͫ������'����y͈���]���mw��g�u,������΄õ/��;�Y-���#)m��G˽�ON�,g`��#999������y�i���^�
�3�G�Y�S�=����g��Y]��%���x5iis��4�>�+Ǽ����/ϛ ��/�Z%J�y�y�{N��A������=}eu@��ZވRl!I|��k���M���3�ƗQ��0i��4���Z{|+8��X+Fd(V�:ʾ�	�z��y>���*m�8>��i�gA��ʦ�t�Y�Q���ݽ$p]�vw���<��c���>�irL\D�`�V��I��%���N� 8�v����C�;D����z99�ש���T����&�P�V9�c"�%{��.i:C��@ �Z�H{�P�@E[攀r��x�nnH9�p�mim+���D��������>kޗ삱iAPТ�u��^�`Ѳ�T�ia�\��<�6��,�S���i@M��~6	
�x�V[Z���k���1U�l��uMr�x`� f}M�nXԽ�; \
p�8���@os���}�[�x�.�|h�PHHb�:99`�^��G*Y��с�+6�V^Xg6Pb�7���+ ��Y�i�^2�֍_=t!h�r|�� ��l�[[G ���@����$��>�q���kh$Ӗ�/�٦�E��4�3K�^�� ��M�ʕ+qÿ?�F��?��/���fe6X�`&��������MD:H�F���G&���5���C}?g�iL���k��F���k�������&nӕ�=�5��Xd4�X@����Ӂ�3�ڢV����R/�������tК�Q֝6b`%K�w�I�[0[�[7�Fm�-�	U8�[&�𴿯ﵓ�|[���4�@�ᙂ����2>�.!=2�;x�[E?�]Ȏ`��^:W_nь�����I/2;g���y���z!�B�;���k]W��ܚ�AR`��DY撌)��~��fR�ʼj�d�dF��9� �R��&XO�p]��e�������v��r00�o��&�7������M���ЉkY��������Vѓ���<?�2�Z�):�ű}r|�9���E���.��5�@�K�A�e�� W�r��dn��� �Xsp��e�kViPh� +��J�N�Nd�C��TFÊn��p�Y\���<��i�j|��jp��P��9p�"\)�~)�m�|�m���o;�S�,i�#�'Z����>��8��^��3M+�y(�`�o`��_�~��4j���ݧ y+T������e���y7�d������(����7��怇�&�U�K�%��-2�a'�,7�"���XƃS�`CD�.�+q��Ȭ���v7H?��Yd��3c�{�cOFg�!��߷�|�h�(��\���A��Z��q�b��S�����399�gj|0�gg�r�n�+Սu���Zd��H������N���_�d��&孊]ݴ�C���%#Eeu[	�jJN�h�W���V6"�%鋰���L�1,��,���%%�oh+�k�}�&K���N��u�,M"�����}����d2&��K|޶\�~]�x�My��	Y���J�C��J�"h�2��� i���s�E a~�����ɩ��+E ��\�'���_f����bt��F���flf�l`�Y���8�5�v�%�QV�L{�"-�aj\��ÓR�5(��R�$�t	���7�ۍ�]��al8��ݸq��*��UjFs�fO�ג���x�+����ۥx�7���Vݸ~�N�kkl����Wo� d#nB^�5�ٷ�.aH� �ηmMl3-�����=r�(�)s�T�7 �9	��������L�v[Veo�0�{-\+K�<��Mǥ�yd�`�/\��2V�L҇�M����'@�t�LI��4�[�Py�[U��c�����3��Pi��� Z�8T�^^��%3���]����<��	ϫ�}���K����'�����і�me�g�=ӈr?1�8��sw��ӵL��
���x�����s12�t���oQ�3W�7��2��4ScVpX��lC6.m����h�eR
��P�7ӎ�=ί�1�['�E� �(m$Rrõ(��3��-���=�^�M�`�vt�lʡllj��¥���eg z=c�9�TΕ,�#d@)Ø�VoD	d^Ñٶ)+���0(��;U
<`jY��4~H�h +�Z_�d�e������?����!Y@	Qs�ό�%�j�i�m��+��?.x��ʖ��K�l�,��2������ƿ�׬>^S������e�8����������`��`	Hn�9�G+���<���G;������G�'-V��"V!�,c��l�"IF���"x�g������lx��L��"�3m��o1jC�@�h�	Z������kr����w:=�+��Y�F���.+K��ꂉ�0�w/F�m�yOO"xx�=�s�P��VY+MpT���
� �������{��(������cۘ`Q����|�7�i�	���� ;:A ���wf�f�Ƹ���V�-mD>K�[� /
�V��U:�բ��6J^��Hhv���o,r8OЪ&�QT4)�����"���=�#0ƦR�]�C����;�v(���ЮTSM�M��(�ᡈ1/��Ӧȷf��)���c��!x#]�%^e1��f2�qLB�
=l�����M�z^�ܑ*F�Tt�A>Zڈ�cw[�� �U;�@�2�Z �6�	��)@~��.���\�2޳���w�}'���@�z��M����dj�4\����L��=ĵqv��x��{�]��A��1G&��ĹG��.Cqڙ�|�&�K�h��0������{5!�\�UR33h{W+�[�A6,3� ��a�]~+�ڸ&ރ��U^�x�^�B�6�k�hc�향�5uܲ�lz-��R�XuX����PC�-���YcA�[nm�89�7߼u3���ީ�0� ��)��Q��Ja �ge�����4+C���f�!�������6�s;\�gv�~>'i�Xe
�W	��Z�Mb�_.��zasG�UBRF��(޽n-�����y��u�!c��!�i0�У�ȍဟŲ���o�9*hE{ࣣS�i��q��χ����� �ʀ�l_%��z��r��~��~��HM�V.��Y߸��q||��V�5��x]���?��>��7��,l��� W[�w���6=r1���LdU��R@o)�;+;)p��f�^��in�([#��P5�*I����{�@zp6�BQӛso��Z���h;Fw{k�`�hp�p7�w���t��3�j�5?f_�>�5ftc�^�ԅ����ܫ��S�u���N�%�����B��?�;����Y�e z���'.p���=4,P�C�W�d�=w���F�;qQ��{���G��� *�XWGg�>J; ڟQ���rvG�v����6u��)>L$�t��b^Mݑ�s3Ħ���p��Q�.t`�L&��.�풬��=j�P��3�~���;1u�����xx�������[0����ԭ(�<�;X��H]��Ѵ{�rb{*ϟ�����E������~���e�̻@y�l��[${�JvP,T�+I�\���#v�)X����.�	X�w�}����N-.6����F|�w�y[>���q�yE��6OOX9��=f�:}Q`5�ΐ�רv↲�6��̡:�~���G`<R�9��Ύ\����e���c$\dd6�t�x�2�d��j��R���gk[7)���Kk1�89=&#}68��r�rC���F��u���9:N���Y��(��� ����*���?xOn�~K����=���c���&��Ea��' �%+��k�v�#JP�G���[����.RZ��N�r�ˬ��R5C�{ ���:%�wh��}���t�,l�n~S���p����������![��ti�d-�=(��(>7(/�j�ZG��b������X���2$�V\;�1W��7r��2}�b�#ر��Ṷ^��
;ņ&��?�̓����Db��Z-S0��uu�Z�b�b��歒�[츩���~��'~M���<��y�@t��&4tUc���H�db&���pTf�����@w�{Ȼ����A���E�&�1��d�k����;�ַ`��Y	�jJ�W����&0�q�pw�v���_�����[����U�1�w�a�8�ʈk�>3N�|�-�*�pBu� �\gZ��i;f��,���� F�:'"D�-fd����k�Iv��iG�{|tBV{0\���5l''3�Q���tl�[\S&�R7�Nkf)mj������l:���SpH\ϵ%����h���fվ?/�Oˎ�$F�{��.�S��?�6�a1d�/�?q�[�@󢵤yj�6;���rY�l�$��i��7�0��4>�+{���C���Qk��� �6�u����4��1��M��>qd�\�G��Y��P�@ ە�-Y��c��gD���z�ɍ^�%�F�'�w��Ӎ?G�=m��� �5�]����lkx6��ۄ� �G�HA36d�<�k�C|�b���g�� �^���lʚ/�j��f�h`s������A����7�Z�3w/R�R���5�>Zoc�!1/��.�j��d�7Z����_q�d�2�G@���KZ=����e�+�Pͼ��,������#���o��o䣟��&,��4pn VX�aK�v@}-x��`��o'C�������Շ�#��b3���k,��f��1N Ux����^��P��p�"�<�ۑ�x��/]�ԥ����8v��Ӛ�Xt��*Ҧʆ'��1x���Z�	|�g����	������8���c�����9��)�����_�`�k�7����=|@�w�7d��P����/�����&�Y��`��)��;�I.�S� ���l\�L��?�x��fZ0��W���3:&���ٙ� ذ���}����>����{ڭ���Ҋؼ{\�� Y���m޿�N�.�q�0��e���A��f�������Jq�����M���߹_�V�2��\�`m@�eV�>�8��Nm��g�d��ؤY�Zg>�[�u��B1�Y6�-�Q��N�<w��3�/�u++	�Wo��J[T3��R�y	��}�2XhUS�/U�}�5���Z
����#��e���{{R��jǤK[\�ϱ`-�K+�L����2R(�����'�i�iXTX���%��;w����G6�ε�U�V��uO�x�����z���s>^���/���~����	e	� �i��Z��!����h���N���}��v7C����nMVY��*qh?���A�z�17��A�F�����2�8(-���tOӶ���Q�.i��x�@v��UP�@@�L

�P��q���6"��ײ�5ep۳��s�Q��i��✟[��$�0�s-��w���|4]����U9{��>��e�����=��f.G��=S �8��{�,�q7���K&��u����Ѻ�_G�>���г��Ш2~���5K����S��1���N4VZ�Gh'�BQ	XL:l0t?�㿹u;r�<K[|y.�-m��d����PO��	<���󈗩�A��s�Tp'.��͕���+����Z���(NP���T[��;lVXt�'�P��Y�\��f��%cM�y)޲��f��lN�
[��N��H�r�J5��׽��m�qzՋ8\��/]L�6'r�)�C�aI���&�w�����*����m�� m��ͪ�!��� ��������؁!�A;�q]�?���j����NХ�y�R���cy��m����-UO��X������7ul�T���+l
V��;����2M�}��]��O�dEƪ�� ܑ��"�����^{�f��II�
�3��i���&RW�[���"]�����#4&���ф�"��{�m��o�-7o��k�J��_��%8���'V��6YBI�7�`�QE���=��?�,^�o���@������z�h�:���-�g�̬20���ƖX�4&s��X!�Vv+�;:P�1A���4\�~M���=��!��g2�>9j1hnzֆ'�� ?R���G���k�*��eR�x>�s���Ǭ��f�˷ Ņ��������z#�x�@�X��y���v0(��\ :_�Y�zy�Uc����y�ٛнh�l25�~?.���+���K�h.]ڤ�fcc����>�18FKgܗ�I���E�N��U?�tu�J�2���|` t_>���5A��2GM����e�F�\��f�Y(dP0�]�A���0f����A�	ʐ�=�2@�,�mh����FW�?�����W_��M�d_�ڼ��e4Ӧ�3d�R�9�`�r;H-�T���=�зR3�Z��/�����`C��K�vL�I���.t��J#fWf�6h�<�H%��S^#ma<���'f�P���Uo^�{����j�2yo�4�DP�,��Lp�����42��s�;��^��X�K�.>��e<|�9���]�Y.<���Ik�.���H��]|uy���:�W/tYz����u�o��C�Z��AԶ�M��̵�iθ��VXA�c: jo�K}IճݓrT.�!';]`���?\7h�dæ���q����8�W� b��7�& S��-��D���A\��jmƐ����dv��n^��i���q�]h�`@?�?0�74�@s���Ek�0
6K3�/��S�1�.k�k<Ϝzd$M�%el,ԓ�1�g%�}�a/��7�c��>ݠC�����De��s��*1BZ��ai��B
b|�?��3-ʸ�IM64�m��X���е���,6-�5����g�ɽ�y���q|�Ѵ(sF�E������A�
�*��z���@�������w�p�fa��~��"0^т5�;���r]�i�Gۻ,F��{��e8@��Up�G:��t?��Sz��@��}����k�d{�*�6E�E(�������xh�|Ɗjhr��������'_���q�B�>}�篮]�ǽ$�k=�	dG�@}k����9c1ҀZƳ3�DкH����l6��zJed�n � =� ��q��@��7ߔw�}W>��l�1���_��������Z�W)�A3����R���6�6�>}������B��ʫ��-\|������Ǐs0c��<��]_�k��<��8l�JE���y�L9L��C&�6��R�5�M��$ߑ��Zc��X<x�S� >����ϥ���3:c���w�Ŏ���M�o�Y���lL �7�/ޗ��˓�d7�3 C�� p{���re�
���q�=��I��o�הm^+8���h�5�ox�7�17��E�����u]��/�Ɲ��[��2���� Զ\^���SM��*�������������s��h:�Ош	:�T��	��h4f����ꆸTG�M�!�*�PR��T�t7d,x�,���M�F��#��Lav��
�E}�iPF�Zó=��;�0�B��%�R�Cm��Z�3e�32�q]���X��ሞ������?o&�k���<���5�w�z��|0�+Xޗ~,��8;�.���fs���o��34^�<��/��ܗ����d���4߈������Gn����������<�
��o���닑��8�\�6��p��a⬭\����Y_�@v;�p%p����\(�r��Y��B ��D��Tb|2���SJC4yys��^���"�Њ�v������ll��q[{{�eO�\�[�v�Bd�2���*uK�י�%���b�/'�N��%%��.;�tzmk�a޲&���J�J�B�K�(���2�nD���jU�-rg���i�f|�Ӆ�6?�5KZ����Ԙ�M�J��ZeP	�i��O�L�H���<z�� P}��7�����K��	�W��Y�5���c+{�����{y��17e�M?}�ݖs��?�
ؚwn�#|�\� 	��E�S�Ҍ_�u܄:��؍�66\7�~W�V�YJ��CN����f���3�ױ�\�9��"8V5�:p�M�������@t7�G,���藿y73O����3�U��z�f>�L�o���#�x�Ոz;j�/o�߼y��[��]zq�Ĭ|C���%�{����>f��ρi��3Y�g��&c)�� �.�6���=��r�rh(��}�7x��\�L�$�	8 d���_��ċ�Js���o�>��g,^���k��o܊�}��#��@?���W_����S��ۧ�V[�q���b��L2���9,��u�'y�fs�4��*��,���hi���y[�~��mI��"ɓ����wM�ZTs�,h��?�����LR��Ǳ�E�5��zV,��ͯ��E]H ���<��e���,� �y㊼v�FP_ц,��o8e��%8�66����s�=�Hk�5����ޗy�EH���Vr��Z�ۏ_�r��y��)�����/䂓�/�8�'ت�1�eC6ԁ��믿����F6e
lH���aM|�^<�)�
�S R
�s_]��ZH��CƟ]׋9�zܺ���[5��28-^��(��Yn1[��m~�N�m>������56��9�~��@w0�	9�������V�w��ឩn8��BL��Pt���Z[��f#?Y-�|F�Ē�!3�a�9�7$�1j1��o
r����:G�̃��aftMnz#��`:�:��u�2��p�ǋ���Z|���P��Y�sl�s0o]�_՟`��M�p�����a��)���)Yԅ��]�jo3�ޭ8A��My��Hf젢��b �=�	x�.�(��ظ��Ϩe:;9��V&�1mO._~&��乼uUV6↸c�6�V�*�];���Ҋ@/9AկV)g�P��v��	���(�8��wO����<v�� &� �m�Ƣ��P(�vP���`*V+�7Ѫ
5��j�*����B������4�f*�o���6��i���iܥHۃ�z��g��.ٴ�^n��m57.m��w���W��/0|�C1X6��O�O,��'��e����as����^��
� � 0f��C��_��|�՗�����+��y�ES�,OްEJgI�T`����4�|��U���C_Ji �K�6	�Ɗ��G@������-<��u��Mvk�� %@�6�s��g�1�Z�-�ǲ��'�޹��nR���vu+������5 ��# � R�D͸� ��{���R*W5�c>tA��yK�C6����'O��x�Ppw�`����>�������w�" �S����I�	�q�o��
��9�����PuE]
Jl6���	K�Kd<���x�w��c�^�q�~�PKB�R l��\�fE��t1k0�>���d+&��ۥKs���:y��?O7)/�ϩ���T��s��5X���-X�cA�"O���un��XI�,k>���|J�Rv
�Wܗ��%`�������<�b�����r�h�2Gl0���,]�uQ>�%7%:(Ȅ~c����)ZPhK���w�/����vr����5����B��z��.�N8��RM�@~��~�;㸶`ǆ��U@��l���D���=��%�`S u��}.7'�˴�^�z6�1fw6Ӗ�.O(9�̪��p��	���l/�
�Y���`.N��3������{��̲1|ߛ�3��o�,�]�Id�yW��IXF�νm�sM�>�{ο��yo�`ݟ�>���Ԅ�^?�u��3�D�3��NE��N,����놡�������ěi� s7���E�.���I�Z�7�Z��s���s+��wU�i�n����A���e�u7c��N�
���eUz,�(,5F���pd�L�"(:���pw_���������l��֕c�r�\���ܫ���ݕuv"��^- {q�C��p�E$�/�M"��O�+S˪�l$�ɉ��e�f -��L=�x�Q���T�7��y��|������u��d�6'.�Y(�L����h �׵��(�1���B�>� r�&qq-��˴�H��j�%yj���Nxd~��]�]���M���"�4@���d�k0̞1�?��C��]t��ăr�6q��������>A`ߥ�CW|��@� �8�7�[p$Zq� ��1~��j��f��tBf-��0��{�{l͌�=�������`����Y��g�\';�u+��U1ى`����K�� E�o��:v�kk� �]�q] �]��[Ȼ�%�'��wYh7����$��O� &`��:��	�ܫۡAl��a`�=8::�`�P>�GS�_��CZPmmmRV4����H�t<y��R��:�i�T�&	�R�6ר�W?ge�F�3��5�MV�G��pj���i�9ñ�F�}�m�t�l��2�B�:,Zg-sI������uP��*c~C���2��(�d��|������[���{M�{�Z�PŦ�+n�^A.<�m]�	@��K�e��I�C�+�V�8�Ĺ��5Uc~�B��t�u��6n��d���e�(�r�	]P���}Y�H����!�`s��@�A�iE�Sj�3+���e�|Ck����Xqz �X�p��H���U�2th�T�7������攅r�m��0��׮�����ul֌x���7eeր�o�U� ���X�0'�8���3Z�1�����Z�� mٱ�nn��a��ի2��ц�����j��d���E����[��1ϲ"��X��m����`AÅO?�/��K�	t	��&�\|d�|v�[^�`R�x�ǥ������#�Lj��h���RD�#�T8R�-$3%���fq��פ�^Y�$X�@�'�.�8�]&����7`Z'�Ŭd�������ƨ{_v����A�ݩ�:
���D���pA�T(]ظ�-+뙂YѮM��)k��{F�]e+Ԍ"�dd<��!.V���$?����P�a|M�"��J<�jGZhÈT*����f�gH/�kY�
V�oY��4#S���^��^Z�d�������Tzj�x�Vdd.+OWj����>g�&����:��e�ˑ͎hI�T7�Sj���7��5�G<���^h��Y����9�fU�oz�-��΋w|/��=z(�"�����8&��_ Z0���vu��Sy���lo�7��)�3Up���_^��(8�f�C��7�}�s�ư�{�����>ӥS�x�=`�~��uJn�x��. �C��rK5xY���:t���y���z�%�Y@��}a��~PZi
X�=��u듍;���vnc��j�"8�3�2f�fm�߲Nk��n8ˏK��,����R�o��a M8����G�����"���@G��lpb�D�Mc��*�r��j-����@m�Ϡ�,J��'��YMx&$�����4�q� ���qQ6�)�H�;��Eǡ���l�? ��P��Yd��1J`#��{Y-ݘh�� ���"bj������BvM�����Al2�xmz�52���@O��7��̩�CL�lk��MW|-h�R4S��>��!Y�х��3d w��uvԎ�����m��b6 A�WE��@�mim�q�څT>XH�z�=�xu�ҥ��G��@�R���o4Fq�@5Ģ�XO�V[�E(�ZK�i�P'R��F���|����Z�_���L�1I5 ���k�f�ؚ��Y9�.r���l]nS���� ��a�/�<x���X%x�!�zϚc4_��D�����<O����s���c��_v��������?�V�Kq��ÁG*N �6��D4���7�J6�nH�=KK�a���-M��k�JO���tq�r��d��X��J�/mwp�1��:@wW�>ݕ�'��{�2��]�%��}F�ڄJ��`S���+h�'�~j�j�<�N��[��ϭƽo'.X;�Xǳ��K����gz&'�C9���u�t�q�XiIg�-m ޸�]���I[1
7��4b5[����~�K�`1/�phs�z��L��4`Y���T32�	6/�$�:nTy�C0�B;$iڰ�ң:�4�w�����U���`! #�;\���נ��:m�/J�i�nˮ��5�ŸvhP�vY�V�+:<@C�n� X���'���ݏ ��	����#y�uO�~�}Y�i��E�L�W
x봒�\��?o���,6�}|�Q�ԟ>y,�����P��/�HP��{��6��:��0���0ҫ���K=�O�!3e��9�5)˓x�Mxh<�7�`�(x}� WQ6]���6�r��SBf���U�W�^���<~�,��A��]�HE;nC6f���;F@�mw�6B�iN�W��_>����e�{��#%��C��pS�/4�9�`Zm���� cs���5�]hӵ��vT�Ϊ��E�#���h�A+����	-����.��ܐ@4�^ϗj����V$9���W�o�o�ϡ�i������A6�4%>�릖b�gZY2��RB&�w���
~�-���t���e�k}m�*]CN��0�KX��sVіvH��Ի��g��\?���:��[���u¡�n8x��(tL��.��`���е�u`-g�^��$_z.��:�ANF��wn�q��������J[��������[��K̼�;�z�/vYy�K,à�gMs�	��Ϧ^ǆ ޙ�t�l��h�����٤��͂��?��Q���J��ړu����[��N`7O��?���1\�h�h�`s�g�]�_憶�s��G<Z�&���%另��?>����!k^L���B��A�٩�7s�����`��ѫ��=�tU�����1�1:;��ç�0�|g�X��Л"{�Ȗtpk�g<ҕe\TO�Sy�l/��.�663��mv|C�B)�:`<����Bv�� ��a<��# �6�B�Z%+�]Y]���JPW$�/���D����l(m�ށ`�e��J_�vlj��?�7��{g����DU��1�?Wl�.+ՔVzo���Y����F�](8RF �I���g�\(��ئ�&h���nx�櫌D�/��a�E���֝  l�3sp��iD|Nu���psF��2>n>�;w���SZ�t�YY�������ƶ�v8��`xs0q퐢���/�H=�E_�V�A������^�4y�VPw
�r��鷵ः��q��ۑ~��0'�e�/���c2�6�|2�g�_�A�ӄ}��FB�"�;�~K�T�p�OO�\���˗ջ7uh2a�q�2�j0�Gg)0{�>�bƓ�3y�h�s����9~A���6����������脵�w�6fڑoB�1��)��WR6,�����{��i�IAA�y��f�R���M�<�%1su�Z� Y���)y���}u�����e'n���"�<�h�2�����L��uamc�E°�S�[0�G�8x�-��'������ԀV�ps8:9``]ƀ=H~�c^ә%}7��2��W��)/�2A��?|��+,���G ߍcm�Q�>��T�R���uu����G����{�k��?�(�<�sf�b�P3�Y}_kE˲а���sU���e"Ț�����^$��/.C�v��淍@y:=K$I��ʁ�(��`od��	�-���&�?��rZ��v���R��������h���߆:��?7_S�FP��q��?�m�fj�I���mFײ��E��<�o>�?dHo����V�����@��$����&�`��Z�e�����
�����4�W�5���X�w	x�>~Fxcba�9v�`S�ڸp��#8�E �Vk��É���.֬G� ����2OC�H����`�����ϫ�E�ۓ���Ǩ��  ~�ڮT����T�	�dg���x���M6a!H�-����.�S�ĩh��_���9I��giqS�w{��4�VѲ�b_{"f����A�������-L%�>��D�r����`�f����Ϭv;AK�Y�V?�4�` ��P״{Ev��������� �؈�ش��60� ��	`8h]�!���i��di_S��frz: s������k�w@�e%��EP�%��7_y�+��U�S�����R�c!�ݜ���C�=J|x��
S�	������6I�qF�#;0�olf�:*�o޼)[�[rpx��ѱ��@E���hDP�.}`�!%q�@��y�X���X��Mc\0���]�*��wp^���S��~�`�:�����do� ����Ŕh7�@(1�R���Y�4����g�,Ѿ_����zR��G�R65c#�@���TPin
	K�#3-_}J��0�ρ;�ݾ��+ڋ��V��
m\R-i���C����!��G��N�t �q��J��9�ON�\�;���#6&��ŵ�a0�x��5_�Fl �k��&�h �W^}�c��ڃ=fE��M�Q�u.��l�~�A.º~nx<�Kk��k��AY	4�8�02eu`�N@���	v=qi �E-��/��/+��4-k�6p�8�ը����-�^"6��uVI�XX��'��r4S2�;|j����-/L,,8�����#��c�g�ج	���7��dK�����2�����	���,RZZT[?ۿ�J���)�0���[�����3#�w5���Kj��Rg��w�lղ�� t����uu{̚�Pf� ��p���l+�iL��5[Z�V�$V5�8���.�:��aOH�NhWs#��g�k~��L��U�T�kw���2��z�ͦ���^��FL�ܸ1������I���	DV��;��pl�)�mB)�#eڇ|�%��\zk�Յ�m�ۣV�
�+ѵC7�zz-����l@��+Ch�����|�����s���Յ�?q#�o_�c�P���lRH2�GJ�[�U���K�{�Irׂq3���N�`,	Љ���o���i������{��@�H��������̻���&+�� ���	�twU��y͉�'2*M��ľ촜�&���\��	G�P$o����=Z�����g����f�M�����.�4�:?K ���|B�8��`]��P
Bg5V"M����n.}�ɂ�4>�~e��☁96$~A���1%��炩 � ��n3��, ���0�~�)5
."�Q�7�9���2c�-����+*� ��8EH�#xp@	$��f�]-�q���"��e
Yp�8����r+ ���{?�τ�>��-����"M^�-�������0�2��^rr<� !08}���Xu�ڳ�X��P0�>}�w/��g��
  `	)�޻w���i �<b�O
��q��*���1<[��Y���Бس��/�����a���0ѠM�ѿH_����xK\|qW����r��9	���9ҁe���Q 6��޽��9�H����~�J)/]���h�O?�4mO�1􊍏�CH�I�2W%:P|�)���nx�PT0�{��6�3�Z�0I4��S8�2�[�'�3<Р����L���/I_|�%�C���~�O��	�K��UH&�o�H�����=���#�7�ς�`e��iuV����|�L�R㟁�b)B�T��x��>&/Ź_������b��w����s���Ժ{+�>0�+k����8��`�/*isu&�B��H�i����%�~K�D�����S��DÕ�#���s;����l���s?痯1R�z�Q�W!��m�(�����;6�D�כ�8��};V#�//>M4���fJ�b?R�R8|�B��Kfx���fh�+w�c��N��/:�E�cR�03�ٝ�pW3�t8G��� �H�UP�J�ț Ҿ�,�-��x�X�����s"a�����H��ᱝ@����:�C��_�P��g�
@��=r��ɶ`7 �� r�YBB�DB��ek6OJ��+>�S7������nz�i�pn饙������v���YۉN��o#��"x��C-o�M��{J�N8��"�$5���s�䪭�{��L	@��u0f g�6 �C��=�*vh4<����]`[.{���� � M��2�/'ڗɚ�刏�I,�x��[E�"Ѣux_��c>#�f���5UY6/rK��y���T3I����ŋ�U[����h�g��b��L���	�������,����c�0*.���#|��+�'�ǼpMYᘮ^�ʞ�˗�r:�;���/^��&tqa�/"�����*�j�g�{��~1_h9�V�z���ŝp���`H߿���&�r����&��ݡ*���Nd���+	p��R�l��ķRH����x���z�����خ��Ӊ�|����c`��^�N_���	MhL���_��X�B�t-��@�؂��?x�%ʠ�P���?|��+��0�꩎���������a^�F��7�d�;J �EP%��P����s ��X� �>���/�JT��D����w�U/l>�t_D��Ed4��[��0i%�}�TQ�i�Bg�(�tm�]t����8�Y$P���r'{�l�����H�>5�T���6V@�J�+��,�l�ᗮ+_i���5�!��YaJ��B����9w֕?;��s�OX���5x5�u��l��φ��K���[.�n�sg�ɭ�l�l��O��3��/�N����sK�oB7d����M�����"�G�����K3��dF\�k�����i"�d�:H��s����ޙ��A �:����:[�uf�m ɝ�(+Ȥ�����y�:<:�W.��ŝ�]x��=Bն#�yAX�o� �[���E>Z�٫;���eR+�]c��0j���>ƻN����xz���������Q�1���'���"�0/�s`�!+8J6���dl}2z3 �}?�/�r90� oN1�
B�/�� �s��2���8�;���s�ep
��&��I���,��P7<�&7d>�����dgW)2�����p`�pR�3/�����"	>X��qE1/ak�5k�6�7A@y^�o �F����C�R���ѭ[�,	�hU���S[e��e�n����Q ��N�h1 [�T��\�����z/_�F���a��������
�>��t4�9r����U���E�E����ˀ C$�Pj��ҩ3��Hh8��^���g|������C�]J��sI��XJt[Ыܵ���sn�k]��Dv�3�f,�a4=m�csR"T�jq�_�Y����*x9X��%��-�u�]�3�Mh7�9������9�g�MT	${��\$�#Qh=�$��y���Yq��G�,b�虶aN��e���7��Um�̙GE��k������5�G;N�4�"K��8~�%��q���Z���~P^�����!��%ŵZ�17tر����R��>o����M*���Ζ���_�����o�Y��g%	�rH�bhK^C�3��A���eC�r�B��^���r`��%�~����#��Aޕ�z.Y�q�h'�9M8g<Xī�	k��q����+br��oij��',ͯ�A'�����б�t-'P��#��5ˆ�a"i݄���`�j�8��0��۴�S�u�F]�4��Rjs{��`2�G�Q�b{�e҅`�t��˽ð���wk��D,;�f��e��Z (�b�ar�Di����X����Xj�C�L��X���;P�<_8��)M.��z@���י?�D���+5t[k�d��e���mUŠ�G��Iך�F��Xg��)9%Е�<��������=�A"m�	'�t��&����%�б�SbƉ2G"��+�׋�:v2��I��c��J�D���
w�����Z���{�%���Ep( M��Xnu�DR�E>gJ���O��%J�K����/���x饲KUV	���y\�\o��E��Nʆ��]S(*��1�P������}A�����9}�°��`hy��+eh���cڼq���92�Q��f�H��hwCI�,sZ�j��{H��� ����%�?b��&�g-���,�3/JFg�^=�7�T����4ƼBg���ݒN~1�O;Nf$��ǆl=/Q�`L�H��u1U-T5�}m�������-��c3ІGմ�)�$K�
�4��d�K�>?�Vx��Q!�bNέc�0���Ї�g���K.I}��uz��w�?"�|_\�0ևNi$�.�#F�j�ƹRyU���M9��M�]��<�,cLr��K�����{'�N���S θ��U�� J������B	����)ϋc6��%�OV|R�&e��7���y��eˣ�q�2�VQEk��@cv��_g����6Ѣ��,�U���9� ����2Y\]��LO�g��LE'����n�h�t~�9�K�ȃ�i��ԫoYxzN� y�c�ۇ�w�# �uj6.�,��IgS��Tj�#|�Q�٢�
c�PI�'2g�D:}�K�a������n&(P�Jn�x#Q\m����	k�N��+�Z#��N̳+�W�bVrgs�[,oy{����������p�aŁ��9_�E-���1�X�z$� K�.�K�����b`q��>�2M���6�ߑ|f�i���y*t1g���*V2���$T�Fe���Y�`Iʫ�A��:�Kxz�� T�w.�K+�9	�!L�jJB�w͈A��GV���U�P� �1gX���@*3�G/^�ы�(:aY"RS��v./D�-VҺx1v��D�Ѝ�s�a(�)��F���}��)'���������|�M.ߊjr\�N�� �����P��9]�v��V���:r9fM\E0�\M* $$�-XZLuG��	:)C�W� ;�X�a��˼g�LL��9�*��MH�4�${Ȩ�lo��%�X��^^3�L���8���N��>i�}y/���%�z�%�7�̝n��u1
� N���k��Y1�_��dxq�њr�5�!�hh�ϣ`�a�y1b(�/�#���V6mp�U���=H�ݾs�Kc#j�����O��i	��!�[�ΫT�2����&x� ��(S��W�����)���w�na�ϔ�Oڒ�;ҟ�UC1z5"�6�w�jx�V�˕�9���Lt2����6�M��67�4w.@0����촹e��U���zP�:���8�g��&P_�3ON���?)��ط���#��icg�܂�l�q��2� 8}�`�x��q�,<�u��0��K�P#V���]�n��i>��ل�mF�5�$�@!�E�9�^��$�T3�?HF3��P���څ���n3	� 	kkR]�K���f�:3}��Z)�n�g�����?�f�h[��Il�\��S-^��i�/�� #�������;��Y����s27�H�\�GϼQ�8쇊S���=��#4����&k�n���d��2����]��f��c>��ق!�G�x��E����5-�$q ��h��W��R �VhY.��*a�sjХ�de>G��{��=�򋯸M�F����*ݹ�&]�z�nݺ�ł��'��˛��qoT7�Fu,�E�O*65V�Ix��k^�v��^���	�$'��@�0�g5>����@;~𶬌��7S��Ӫs-w�|,	-'� � ٍ5)n�&<B��k�V���y+����)\���!f�L�Yz��-��sm�@�ͼ�g�b��,��G�~��RY�Vc� 친9��ЮSd�3G�wԕ���H5�V����޲�A�HTT��,{��"*�ȇ�?�%���E��+�g_K��mk`�(m��2���Wd��?�%�)hc�`F�8��6����,��U�����a�y��z�M!Ǟe������麍z�Sp�>lί��<��䫋�o��س�
F��U�ǡ�qU�5��Gd2���2�j�"J4�V��0ۀ�Z}�%���a�'Ȧm�ݶ���u�c���ֲ7׼�~�۾�g�M�����2/nq;Ce��XX�^���d���;��Z�64=�"���(`-dZW���u�`�9���^�6E�MW1@�H����@Zv�j09H�n�ݪ	hXgG�MPD���5��P�G�a�k瑊4u�(�.e`w�5�)�4����+l�#M.Xa}���<!=��E��Gp�d�f' T�ц��ƭ�-��ܦ��V&��z9�ԧO�\AO�Q������'�V�@�d�p� �Wo��}��,���Xp�W�P��"X�*#h�v��Ҕysřj:�U�,��se궬o��i�xI8w&�&�ߦ+#R>��"������H��po�[wnҕ+��ƍ���8|6�E�k�H�w�ei�o�����	�d����0�'���vs5'�LCv���'R�u:�~��]��>G�{��
UK��6*����6#�A2\�4"[�?�6�}����6�>��XDzK�F@��3�Ϳ�(���~�)]YҒ�`怰�WyB��A˛�>�Y��K��J�J�$����@�7ZIq�E!F��A������5pB%;�E�qQ�O���Z�ˊ�D�3%]�ʥ6!5����#��|Ƞy����xⱝ��K�hp�F�[�R�tu:-7.�ð�ؐh���S���EY�|}��U<O]�)9E�p�f�e�O�Ța�ɞ1�7W]�aY?�T��~+;Td�sd5�Ak�dU�6�1�M�+U��r��,����G��\��	eo�#g��5d�n�۹�s��i���x�<�w�ڌ�}l1H�PtـO�.�����'˖�x���l�C��Xl&�T|� �)�k�c�f�]�ǼZH*T�U�{».5��ʚ�J�$�|� ���v�E���^.,F#O�;��8���-���tT����ȋv)�ӭZN@s#x�z#��]�.�;ޘ0m�2x��; �h��dp��	SXG���t)���r��i��J�-��e���]�}�ENy�6�f���ʠ�3=	�2Ie��\���MW�^f��8�D��li����Y��!�A�������z�Pv"w���ڭx;���>k��|Y�TSH.@0����xm\%!z�]�U�U���u�������/��v��n���ɨ���/��^4�q B
j��:�Q�b�+x��Z /���;tq'-��(_V�gs�F�1����`���ڵ+t�ۧ���p��i%U�0�xB2h=fP /�HAU�,%Ql�Uu��s#y�&�˗�0���+'筥�Z�Ngcc1��A��2��*���Y#��`u� Ԋ4
�mJq�q����4�Z����+a�Y�Ri���|Ʃ�����ɷU �<�����)1��ji������I=C�G�aK��̃7@��w�<q/zcs������e�JNl)���u���L=���l��;��-7\|'s6��:)�x�浆��r�VeO�/��:�K�{�{��h���_�5��G�DO�<���}��	ɜ<t]���ĠhDfI��y ���6'���q��Gx���q6vl��Hkt�I�x/���{��+���"^��b<*WEm��	qT;-\ekNz^#� N�����4����^(NkF�sɃ�ﺝt������y�~�29�Ӏ��qenˌ��/��'c��>y��S$�Q�3�+;I��Q�J8ɂ<���(���x�4���|Z'�%�(%�˫��z9����cs�:d������_��Y�fAj��*����� �4�#����c�";Bs/.JDN6�h�6a�4q���"$Ρ8���C�V�M��������ɍ�>t>;�Ϟ�����l϶$��G�gj��|yf�!D	�~h�Fٞʭ�����='=fY�ٹ��~*����8y�}���rj3QD�߄�L,M�d��)'�b�e���A�9{����_��}V �f*�%uuV7�P����&,�O&<�
�q}�LMiFR��Ѱ�ި����"���h�#-��ʄC��a��s��N��tt��x9��������	U�0��쐢ˊ1
 k�'m/� C�W�Z���)�/�����H"ֶ�5]Zu�/)��c�E?��8��4������l�D��joq9+w�.�*��v* �D�	o�n�G�h�i����߲R${�}<-s����U�X�u�����*��Y�K[�R8���~�\?���ai���Y0z.3�6#&�u.�.@>�� �Rֺ�s�3Ph�>}"����g�� cP<���`_��aØ�u�ݹs�nߺ���>D5`HI1����I=��Ū�Z��x�ZL$�$ә��ܰ�����F�Ly�`3`�0%Ϲ���ęx����)�Uy�NǑ&�"�˞߲�H���Dg�w����,u�hAR��'�!�ϳ��f�J���kl'����q�v�t��ļ�ﺝ��#i�*�/�ÛϠ�,�	V��+�sɱ��P�eX��������i6��J�n�`���0�r�PY�5|'L��"��s
�ynϨ�|8�[���Mv�j"����ǘ��xw�񎄧Z�Z�%?f]�q ����RE�mF���͂�*��.E9�@�Vf��2,%�S�B�޷~yKSM`���*R��6����?g��}�^�z��M�C��Hk(.�N��x���|ǋ�E��L!����E|~�hq��,Î��Rb��=�X��@��ytI�c+Q]�s�;N�-�z�ec.�w$�0%��6j����]�b�拼�-w���D�������^u�)�=���EHV��6չe��{�c�V�E^ �4a�nQ�8���F�h��6�>�ʳ�*5&ɋZ�ϋ�a��c�^��o��}ϕ�F
�$��f��66�=�S5��.��WT*�VY��Y��Օ[>��O�L�j��0�7SJ �5�j����-���XR�]*���gGh��iw�_F�`҆s��t%���6b�H<}xF�W�>�'17":�s�k��b>��݋י�	Vu�]�]��JJ^#�ׇ��O>Q��4?����Ũ��$갂��C���ݽW,�5���KzY����>|�>��{�=^���CZ�Y��6���b�9���T��j�y)�+c��mM�~��86���Ǭ�G&�������9���7������j@�N"c*zڹ��ǂi���t%(%�D[�6ޢ��Je_���(�Md����e��-��J�<4���[~%���;�kI�+�����n$�z�9�6�0��Q{�	`*�^
M���x�2!�}�zo�	�S�Y�=@���CK�Na��Ne�����>Z�Ie`�,�?G����N�[5�䝈6��#u��eu:+Œ�.I~�c��g-�/�a�;�ކOi�غ�x���QߓT�_R��=�@H� n�a���Eq��B����lN�ET����`Q�F�]f}F�f~4������r�f�K��K�qH:_r2��.y3��ע2�!�_a���ƚ�J���X�q�J�O�!�i:<:�����V�{�}g~�O"�!{v�g�5���c��]�^$�qS��r�I<g	Q�*EV�7���c�kN�Zפ�.��c,�]CU�����&�䌪����QI|^�}�8�<�EK�U��A�N�r
C�}�wz�-��;Q[5��*mWU2�iB��F�NZX��J	���.T��Ʉ�Gj�4#��0�nS����T���H�-����� ��w�e-��޽ �>�[��y s��� �Ч�y�&�d�����:(|�I���@>�� `q=��Du����6 EN���W}���ӭ۷�|?��������S���f���26��z��Ó���yڙ�[v�L�X�g7ԉN_\���1R��r����$ �q;.e��5�mj�3��<�-��[�M4�Gh�f�\[��u#����-�����G�x�K�b��t�S��$������8�x�Ri�:��񼁑���z&p�O~۟�ud�|K� �\d�'����XCgoQ�ش����bj��V�L(
N)�,�Z ��m��Ź<@@Y`�[i� q����d����*��r����x��Kf�W�|��(yH�R�1`A�Y�?�W�%K����µ�P2��/b���/�Çk��u3.�rHM��I�/�'}��maޱ!���uI\ȵB |X|P��������Ҧ�ב�"�q�����f���e��9�1t��U �{t��0/����p��Q�5�P��,��0�?�M$k6�&+��r�-�z19�.)dۣ`[����mb�ה%�>ʐ�܊/~��:�
��@���s���"�a��uC�8ƌ�FO٫/6J K�Պ�8� T�/��b��\��l<���%Z)�"=k�#�sp��]'����g���O���VT)YM�u<O�F��c�����3����Ǚ�/Y���DKIh[�cr�VL�R��zeͶ��Ը�dƵ�k� �
�hot��=�b��O��{�p�/�8p��(�:����_�*o����+��C���( Kk�� ���
�+�� ������k�
Ǽ~�:]�t�+�����B���H�ߌ�~���p\�:�7޸���D�vw_��s�\��:RuH�l��Xާ���Aa�۲k`ܠ���o�ľ�S����l��pN^��_X����|��E�ɟ�5�1��qZ_�(:s,z�<m�zVp��/�/�,iQ�O�C����VDT����3�������O����pF�����ѕ�yb ں�r�b�����sX��e�!?m� ����:�y�K+��� ��*c	@ �0o��}]{r�%�ʗ��A3�����A��0Q�xɛP��񬟋�'�>z�\-V�����|�۩x��wz������C���٢y��b9a�	������r|��w
��v6[�'���ǢC�P���&*�s`༝/S��l����U7�/>���E�V��M�K�@�j��n��z"�q�ğ��:/��\��X4�9��`9�����m�J0\8��{ְ�K(S�,�5��{6��޽��>�z�@�_ }�2)u>����	2��C�mhg^�;��Z,+Y��]���_=*-i��&y,�)��z��%I���	��N+[��`�t��gO�������}p�K�.2�y������;����G;ݻw�������y�W��"7���T^�"���4�\*��{`�T�f��«�j�eAn��x-q�w9�+�
���*�N�q���H�E�I�-Kǌ�(<�|�F�����~Ho��6ݾ}�����)��UT-�w�.=x�A�� F�L߼y��_�pQ@hCy^�7޸�I`ҷ��V�A-��g?\]x���	c����-S`$bJG�s�[oݡ��y���Cz�����p�+�i�JK\�|z�և|�w�}�+����9k��ۿ}���Wt���
-�d��8��j�ՙ���Nkyn�xLV�-7<�)a^�|p�F��?.���p�ث6����<��Ҽ
#s,U9��+�.�����H�O���A��@��2'I��fු%�n*���~)����+��E(M�<��ֻ8�&��l��n*���E� ��S�I4��CB��_���J /�D<,��JTr4� M�Ԏ܅n`!48w�� ���*�4�>����xpբ6������CK[������{�i�Pab��<�Y�q�O�B~4��b�L!�hl�	�n=��"�!C"])}s��d�^Ty c.�s����!O�ybL�/K^Y0�k#ZZ�.
fDZ{Zr�+��G�]�Rl�{�~���F�-HY�?���'���9bх�4��Xhʩ��׉�;�wC���n?
�����߹Lۛ#zJ%�3�I��T��n�iH���A1hhc���̳�CLLq��IEKd���O��8���J�
�@ʛ7���U����J�:?���B��7�8�xi��^�Ho�{�~������r5:��`����Fh��Ͽ�v��2N}�K�*{���/`"������	��m�=�7�����~ZNV�&�Ub��笆�yR��+�NH�DIG��"�q�:���?�}�Ax>��:�υ�����)�quM �˗��֭���?`#dg�R�W� &	�PD�c@E�=�hD'���1Ƴ���� Ǿhx����(��p� l���P��֝���q���/����iq#/c7�Nh}O��k�1��7B}���0��Ƹų�t�a�K�mM��RF�F�8) �����������N�P�Dx��JI~�<o�7�r�~E�ȉB���M�U��N.���J��w��Ѯ��͌�d�m��ͭ��d��2 c�f�:G\�����[:�?�{�o�g�����U�-�ç�hG�d������������x���s@i��z��A�4����W�;z�
�rO��GW���l �N��O����jL���G�f#)��NՍ�*T0����5�lB/vN�ɾ��ts=�។)j�a���o�Ҵ�&�|���/����=�t�DVu���Z��G�4d�����E@f^�.�ȥ��`2�+k�(N��GLh?>����p�sZZU���}���2��<�6t��Zz@!�۴Om�']�8�8�u��uQMP��h`�k����D�.0�rQ$	]�Mલ�\&i��	W߹h͵qr)�I�W�Q���e�	s$�-�s�����G2�f��z��
eۛ����8���\,�X����4C���Ǣy?PG�.l���=�$�m��g`ɞ�TR���͌�\[x�DbQ���S����~@�o��9�͉�h6k9�
�j ��O��0f%x��D���I[�;a�Q �����O~D}�/l|��]z��Y�h��Ls�@6���s��K��k���&e��G�����c�,D솫 fƅy"'�{FK�-s/�������ugr�>�j?gʇ3������?�a0&ޢ+W.�<�;��n�hN�p�e�g���s��-%�����u�|e�.��g�^�؝���@�r�x�}��}��W�ʃ��%t����H0Z��큾�3��� �O�<ao+����>�2���rL�sU]�3$��)���|���/�# �����5�����㚂q�c\u<�.8�a8�X�T|\�P�QvŠ�,��&�V% m��杵R��O�f���$�Z�;�����d�X!��#�!L���q���Q58ދB=sQ]b���j-�&ܮI�Y*�)8���7PU�P��.: e�yv�EY2*�;��*��_-��S�^��U�6��'��nCt�x��2[��n�z�o�n���|!_��@9mM�O�P�y|R���X��;�}���{h{�����X��~��IQ��?v�+�ɰ�M&Uʩ�Pb�9����X��x�-y���w7v���`'l:Ȗ����������� 3@�a�s'mʞr��75�e�����'�6�ne־�SJ�)S�t��n�l]��y�@*J�� ��>e�nU�u9��l��>ɰ�]��K��,q'�GOQ|?>7]��?3�K8ڢ�� �γ���������
�;�-�KWG5+��!c����^�D����-|Dy�d8K�7�-ԙ�'�ΕE��0���<ǳ�or�5�(�/!�Ԫ�T`�����ֹ�xc�|��W 
'���*����+�9M-D u+��~��;{�.���G��?)�����Nj�4�lA��aa��U�?7�$(�YyY����z7	���t�A[s	n��q�[@qa6�һ3<G.��I	fx	AX����x��\ES4og����d/@ߓǏ�O�ކꏸ*��>L�p�e�g�JC� �X�2 XK5?Q�`N��Y�G�vוU&�y��=[.P���[7��7����8ƣ���<0�j�y�˸G��q��-z��wX��ʕk|m��u��O����1w��%�D��|��Gq �LE�/��%��#�v�:a�ּ�� �8s*l@�`F���<� n8hXO x�G���c�:��Mq=�is��C�`[�Sؔ��O���X�N�Ϝ�}wp[-' G��x	�ԣ���s�a��ߖ8�C��'��%���m��2��ݬ}�d�$���N�z�;�g����dy#~8t^�t���u�F����sNRw�|���)9+Js�WϴG��=u�V>[kd@�H6���U�.K
	�zR��>u1|��ԝf��i���ެD�뽊�3��t�"W$����R�3�WPyQ�Է��/"Y�҇�u-���&�.|�(�<|{��%Il�*2��{�:T�:��	����x�- b�!<F���/�]�Z�PH!�3�݌�ɫ�ϫ�ƫ�Xq���c)@ ��1XA��̦"�g�C�a4����]:�Z�=H X=z�^% ��2=y��?��6I|�~>���Ϟ����]̥����k�֩pϪ�����*i7G���l� ϖ93�ș���Y��<�JQ0�jK�KI&��G�]_1d�	 ~�i�B� ����� ^�� ���U��%�?y))��W/�8�?n��/�R4�F�΅ 
���W"�����_#�l��
0�Jh1W�[ŹN׶�������}U�0���q!�:ɳ�(Ko�{w ��7ȥ��2�a��: ֑T	pt��@]S�Ï��m������F�����|hm(����@�}�)�} y>�=� &Y~O�]�+��	�ሽ̸w��@DL�Ȉׂ=���B�r�/l��ƾJ��>�A��b����{��i�����=b0������Ng�֌���ZZ�~y��g��?�C�9��|j�Ӧ��n�\�V~��%�Tڥ��ɤ@pig�{����K�<�����ZHJ�.�xìS����B �q7e�4zAj��k��o��S= 
n�0��ߊ�c��}ֶ��?a�<7<��=�ă���� 2�)��q+�/�޼~�?�����e�ǂ��<\��s�L'�xn 9F���C�����I�c� �m��'=ݫ|W���	Z�7�n�>tV�)\�\u8-��;�S&�	��0�$ ��F�(��qX �MhOo�;�IX�&�a��ڥ����:��%��eG讽Oq;,�a�m�x혭�f�&^��ۤ�9�_�<MY��˗�D�T3�e�o���?�� GM�����x�5,�#;x��l-^�v�^/�_�Z�N¼�7Û�Pa	����h9�@�*��z�W�L�5?&�em&�����L������������^_$����gR���ͭ�����K�0�!?~��"O����;��q��&�m��p����tq�"S��b�����iH��s���3�/ ��[��E� �������Q�)%��vC��Ng�݆!��S��?|Nw�z����?���>�} �GZ �?�\���ƍ��_�˯���9����|0���ч��	P#�b�=�N�E7�e�9��S�D�%�M�AW,���ax}����s����5c��� �yÅ�&�6��q9��͓@[a�Y��* ݆�^�����>{�i04�lt�j��k��*k��Ɨ��G��Ku�DPlڒ3��X�㬇�{:h��5"�����i�e��e���ǫ���'��F/�)�֜�O	 �$6�l�;ݕN�YJ���T��H|�ZoÉּ['�I�g�'��&�U��|����~���u���c��n�v�sŶ��*�.��v�yңQqw�z�	�;�=��?�6�2��w%�xLa��� +PSƫ
�L�ÀW0��gY�[�v��y�v͝ V	9Vi3��6r�2a�t jPF�x�/d��;c�t��M�{�C+%��X�����
��`�!��W��Hl�J ϗC�� ��8�
��%j��z�6 `��L�dx
�m ���e%M�����{>��*B� 2��g����#z��9��娪�v9����\f% x��N���!Ӯ��w,�)pϦ�;4L��}!��AV��ͧ���#v��o
P�
�	�.�G�<�K���t+ɠ��H@'G_F{�x�"�ی��;w؋���IB%��9���_��$�����>=~򌿻��ŀ��a��c���s��a0tF��+J,5��OPч �\2�9�]�q�i��ē�2н�y��#�^���ťJiy��$|J1p���}��	�Ĺ�0�>�o��+�����s�jC5�k��+/]����[t���Џ����7�~˅,��U������p���P-�N�i�#��F��0��%n����M:j eH�1��m�����h<����P�$��1dAC���d�QNt��`dΏ]�����Wa|�������	�\�N�Z�Mr?��N��tn�u��2G����0[1��Գ�~�l�����Y^�Ϧ���
g�]�wZ�}K3�Wgc�U��)�гʒyu�G��"�h��1]s^ο���	�O�n�VK�KT�"&L�VωYl����0�AlקB������dܮ��[���<��sg�NB*Q��"�	����(Ӛ�JU���I*�y[������������{o���kx餴�h�^
��ŝz@&y�� �:��:^��ρm���T#�8Ti��G\�K2 b4�B��J�~tS�Lz$v�f�h!�e4�k_��᭽z��<�#���p/|���{�r?��序g]x��?b��!Ӛ%�$����0�@�C��ق�P��x�\a�`�H�^E"N��g�
�\ ���=>_C���p�#��utxD����*GXRV�9鎎��:6�6��֝w��7n��H�F@4�+�������CbH��0�5Ӳ�ˀ^d��(�������k�B���2�G=�>����|��&�es�b ���t��Ws��X��
����91���C�t�
?������}���m>|J���u�0)�[���N6�l�
�w��C���7����g������0c�i��~eQ���=�WH�J舩��|��9���G���_p�`xym�3چ9b��S�/"�^��g�}F�1}��G,qv�{@������;�~��_|N�|�ǔ$g#���c)� �믿��������� �·{�=�w�������D*��"��\uP^ ��+����5ˆe��\����l`➾��T�
�UK�Qz��?����>�D���6ӣ]z���6@�wkk��]�����˺R�ꣀ�u=Y ����A������w3ks5�^a�~?[l���h^�E?��]q�w�!�[~��	AI�>+\��%}F�Y�Ϻ~I�z�k�������s���w��/&���>	��c��<�b���!n~L���ٳ�u�����Fj|W���O��W��ɛK}-��e"}"~����[UY�i'S0�����b%�r��m_=�e�'f^�Ak�B�ij�g������+=K��9B����I@[�w�=d�ûk�l�5x�1�À�3�%����M)
�����e��S�P����M	B��a�x}�od^��H���� �N݌���Z(ڋ�P��̋5�|,B�^aA�ѫ�� P ��s��k!�`�"�䙗۪l�����x|ޱ�4�l�\iQ�X_�H}[%���Y��5<+,��G) �P1rf_:R�s˕���11�ں��?y�B�8r�[����gt��=6Q���'�̱�r���ݒ���Tz��ӹ[z�G���8��!�j�.G]RdCΛ�������Z�UT3j��ġ�P��FKj�}���?x� 
�l{{����<�B
���?��>�O?�����=~��R��ױU����F��E ���1=<O�u�s��F��[��aT G.1��?�|�рC��ߺy�~�_��~�3�ٟ��KLF㴢�XM��gH�xa�!q���M�|���g�2F�7 �˗v81�����ߔ�X���K_��K/�6z��)K����X����"���#����is��J�^��s /g
�ہ7�h-�w��;;�t��e�v�rH�;��j/�+��׆�i�Ԏ�9��ИS�4c���4���m�cx�s�vgA�}��#�/�GY���$��2&N��2,q��ή&~=sf$HW\���˞_�;����z%�r8�V�S��<M��k@�Կ��8���h��J��N��$�^^,��2���>���Gfp"�	�.�����"V�	�?���	/).����BN|�A�]D��BM���qK7t��w�xw����eTט��~`��'^�:)(�r�$���$�ߖ��yۗb�U��+h�sJrW�2��'�~R���N�9�5]P�̸�Y �T"q��y(y�b����*��,be��p� �g�  �T̶���6M$�Iٌ� -ءq�4	�5��qXh������H
a10����,u���X]	�E!(�:=���(,¯x1������b%�F��f\��e�������{E= $���hP�?������b��k�9��Z�(2�����M��I��<k\k��#�c��F�ݧ{�2����]�
`�e\#����n O�oT�bp�b���"���=x���Y��ي8��*}�^J4s����kUsM~�~U��']h|4(��B�J���2�[ۦ
��$�������j��1���%��aoNG���K�O���3wv���s��߻���z��W��MN��1h˭s  ��IDAT?7"))��$.8A�$��B��)�/�1��F��D�������Q޿������ۿ���y�=��l|�A��$m��b!���޺M|�C���_��#����_�����ǮН;o�'|�e�^�d�����������`�镫��/�?�?�r[������|N�-O�i�c��`.c�5TD���:Gl�s'cjz��۬���E?n޼AW�\
��Gs�Z �@b���gt��g~����A ��Pk���x=���DK-kL ����)���7M��J9{� 9��z?�lk����-Ӿ�ú��"%���8l9��3�MZ���0����5�����k���h75[�̌����x���<!�W��%�"#=d[y/��+�_�y���i�R/��e�/o�%'o�,��~�U�O^|�2�P���i�+���aj ��.
��.V�:���T�,�g��Ŧ�-�KLt�O�|���%�����e^g���è9е�ϒ�⽝a��9�;z͸o�g���Fu��२M�ʥ�p,.�TG�V�z��D�	�ZVK�</������{��GZ^����ޯ�x����T�Z8�f4��b ��4��/����o�
���-U��b�-x�Dj��c�?z���W���qJ7�����{���05B×/����>�5@�k�Zmq����j@ӫ���d*P=��}�`����qb8�,c�	ju���o0�(�3�7��G;�_=�x�����y��7�k|�~��I��6���p�H�<IT�I����O�Ȋ�F��@>'�x��׍����]=��?����y���'=�I1��z*8�pbʵ����l۩���a:���ρ��U�NKW._eP�����B�a�ӣ)W[Ë�w6�`���ք���7��Ux���~����/��/�Q ����ӷ���� x��=��^���>��xnk�B����o�,��C�Bw��U�[l��Tܞ�tc��s�1�>�A4�@7�9nļt�>E^8n	F�������޸~��}�]�q5��Y����,���K���j��W���~��iO�<���c�
�2#��kk�O*��5� �p?���y�x^��y���s�ۯ�v���y5���ٿ�8�n���X�g��h):%������˝��.H�&�1���+�u��0��u�U]4\ʓ��ܨY��������V|��_���i���̛"hM�(��u���N|�~�]�wݜy�ٹSI�ʥ�U�m��o�jC�]�d��r�,dq��ano���m�ӳ���Y�ݥ��|�O��xBE}xa���-�N�.���M�;� ��꽮bIO�o�㚷�=Y��Z���K�(O7�NW�sN�&I���>���f�[x�K])7�=kz] �\^��b_�4h��Lu��7����/�����!��J��hЦ�Ǟ�g�S�^
���JZGG����%	-�~�s�Js7	w��K�B���o]Y�7W�Tu
���ַ�޽�<ʵ5T���?�������:{���/�=DS��w��g4of�O"�>�_6ݚ�1�/V��� ��,�O��:�&��=%�)x�;�&�XQ�I�ы��j>z���-Qn�q� ҙ���;)�E�6 ��Ϟ#�PAT}ʢB�ϓ�z��5B<*�D����N�6x��g%�=�R��}���=S�@E����>����N��	'-"��������}z	���X^� �^@&�R7߼���j �(�}��������={A<�/��?���O������v�]������O��{��M�����я����A-8���v�j��d2�6gJNge�7Do8Z3.2��{f`X����;���`|�=�����Hr�z�rL d���~0H��f�/��P���!��6�ຂ� i6H!���'�I��:l�}潟'o'9���a����B>7t3>��V�iy���9�<�g�)'��������9�Rc;ȼb�L�Bg}�GþΦ���^��S>��,�G.uەA�#��y��	n���(����8߷7x���HV����k�hDզ��w+�H\�����üF�ʁ�i���/Zy�	vt��o�ЌoJ.�G������Z��@�prV����RD��\pF3x\�xN�(;Rj��n����N���/�9Y�<W�H�B=��<���>k4�g"F��Z�o�@�� >�G��}㍛�^
`�RX�v/�>U̧�R{�8^�Vq�N������S��9kw޼y�~򓟅s�ɉx�! �
�rR1�ʥ�W;�J����F
�0���+.�D���dY���K��K�b�
 x�D`�W+��@{O�,�`�Ы��
��x�Z�NKC�=�h{�e����V�Z��']�}G�-Rë*8�2׈w����І��a.<����Q���0�]jI�;]���Xd	7�<�#Vmw���� ���M;�|����{p^�1��A
�b�����_���ǳc}b�yȓF�F�ӟ��~��O�S�xtP�67/pQ����/(�G��C�v�*�׿�?����#�����~@�����(��j��s�v�*Ws{��{W�m!�w����BҦ$�u:��q��x�<��βo[a�2���p�U��]	�"^� {��t��K��?a�Aa�����j��'Ϯ��j�?��(��p4[��AZoD�����+e���f���o�Xz��͝�A�%xB.Z�����=-�.,r�b~���Kk�o�8�}h��1����1��M�Y��/�aآ׀��cvr�{�V��=m�"�P��]�S���I�4'��ˡh}��F:����wj�� ^�� ��:��~û�{Lxkv�Ͻ�n��^�[�~�Mk���
�A������I15�=���`e3� ��}��-W�h���iHZ3�-Nj�;���3��V�c�I�kb��]��`༦o�O�ˌ���X+��sB�!��k�J7�&y��ׂ#I�H�]�-[	V�� Y@!5�v�=<C���Aų� ��0�� z@�����Oa�:z!K�y�u� �&�64Z���*h7o��0�x�$�d�-�vR����f�䝦����h(������i:��mrO�6N���9y�/��9+ڑ��]��K5�+�!��Q}�;@rn���,T1^H��*�����H�I[	nS��m	�:}����Ȫ 2 �k$�;��q�s����pMݫ��>"0���*�/���u艣A���}
�@�4&|���`nmn�dYhW�������~���#%�!��H��2��$�x���������D�	�[��O�Ps�F��Z ��v��`�
`����M���� �� +���iݭq{""��'�!�wDo\ړb�M|��Ǟ3�g����m�0_��� �h�r77&��F�e��s:<x�������@����ru+r~��5x��T�!�&� z7�yZ�-���LD���;��S�����as9�rf�o�QgO�^��h*���+?��av��k��a�jG_*E�G�}�ֺ�&N8Z������o��SNߐ�|yj�ĉ�2ΔN�
�+�o����s]s�C9<���2�ˠ�e�9��H�|����w�$�-�?��Y�is&����[)�A�5�G��a�k:.Y��g�W����Dm{x.���y6 ��a��]���9H!��� �HP���/�w��]����6t.;�3gp@5��2[C�����p�J-U.Q(�6���$��BBg�ga�c�4��k"��J	cy˸��6��F6��U�3m����RL��S��\-״��BH���a�J��%q�fǠ������Z��6]عT/^�v����6ݻ��=�u-U�r�4���x+�E @A�����,v������+�)c��$��zg����LJ�p�.��u5��!�n���nݳWr����i���,ك�M���S�z14�c[��'��!���}{{/���P���1/
���<�r�DX��j�6��Y(#.D�FE"%�GI��i�c��q���Upg|�V��S�.��M�$ynYN��$Tk�Z�ӥ�1��DB{�ݪ�Ufܐ̷L	AE�/����ۏ����@�}�VZ^rX�¤���u�ܿw��)~�ӟл�G$	���l�m����d*�j�v�5��W_}M�����책q����,��J,o�y�)5Hp�LU�D{�ȅ����e'�0�,�-� �M60bu������Ga������Q�%�+}~"�m���҅�<Ǝ�}-�MTkl�B��g��6b��&k��'TBq�-��ی:{��o\1m-��gJ�~u�v����}M8�n��_N�_�;���v|��E�׉�R��{����r�*��m��4�$���,���h��L���t6�.{S��gx���?�\����	���>�=�������o}��՟��FU�3�6�zZ�d�6*-���&p�9v�Jd箄��i�b��$��i&��G6�Mz,�6�{K&�^�)���r����:+��CNZ���Բ��$4��D�M,�HB�y�&���{,�����VM�/�8���?�G��eҟ�6/1�q�����-Y��% ╣�x���:��y\V�[=z�b��a7��m��7�<�v�>y�"��B�\iM�
�K+��������L��\��C���� /��R����s��W��\�F��>��5z��$̈́���]�6N���hĞzl�u�=,k���I�é��!`.y'<��'$�D����B�����#M@�����j����[�X�J�����7�d��ε��X&���vZe!e��s�n���?��u��ؑdԪ�9��4�c����\�k��B�I��r��+s��X�q�R04+�$�S3��b0Tu>s���분3��"m�����!������9��WT_p��fg�s\�<[��E��O��2�q��oU�*/^��1!y�� �Y+����0D���d�����G�X�B���./>x�4 �/�Ĝx6[Hyd�	�O��5P�U+�.�	-H5z[��w�_Z�_<K�����<§an���׽�1᤻�`���H�l���&��``��S����������oW<��h���&�
â�.�_�ψ�4�%u�⸾~��V�u��h>����/K]��[�=P[xZ��0�O�O1��?�-�s��j�A���yտ	|#�,�n�`��k�kK�q.FG�r*MZ��Cdz���EU��WmK���.Ne��!�'Y����ɍ��Lz:�����7|�n�_�8/� q��{���C�]������{U�S+P�
oS�RU641���-W��0e �'l[��2'y������j8�&Do�d�8)���ȡ]��^G ���t��`�2���o�M|�g ��t��I���m���=����,�����fIV���6z�L
*��ٴOF��q�-�h!�1��-1�´:.��ٌ�]��M�MY_����S�<��j��V�p���j�����^[[�D�!��{m�f[ʥ�Dܞ)�J䜫�C��\�`|��5z����o��|@'��>���d����N�3���͞�扌��Td������\���g���gn�f�=eJ����x�U�`�F<��`1�kKm������9�O�����po>X0��F'�a��+Z��T���t�d8�t�bT��Vש��ڬ4K���?xA��{�[�d��t�
@497M^.~��K��܋���M�H!�Fs�I�6�˱&����A�,>טMMn'�ܙ��߯�x�����1ˏ��5%m
���~��X�����w�Cs����.kCK�p������ ׷@'n	��/H�=��|�ɺ�����Dے���Bq��9�\�@A�	{o�_�B�a��p�޹D�ߺ���M�"#A���R704�η<�v���p�������հ�yV�"��VǕ�"I9������Z��4� ��Y��9U���R�O$�5�%�ᬯo.m��������c�fc���B�d�F�s������[T8�#r�:7��s�ó��MD�FJ�&3k������GDɦU ��4x}�}yѳ���/=����[q���w���x��G����h��g~�t����_�[E��:r._���=P?QE����Ɖ���o�2�� mj��B���m�T�����F$Y��\C@v' .����u/H��=|���8��>|��>��s���M_}���7O��-���Pd���7�t�+�>w#'�$�\ֶ��!�ԃTa�2�����sA�S�"�uUX��Mb�-�r^ �xFHp�����԰��Y�X�Q��w��;z���(&�<�L�3�5lQ�C��&e1�����36���Kz>��?vJj�4�/����B#�À�M"��]�|�{�I�aꖆ��[�W�g������b�(w[nl;%~7��Heȫ����(u�۷�"����)�~�d��e`A�w�}���=c�H�}���"'���~��_�˗{��ž�FD� /�sd*>��[7/����wF�h��8'��xU7'���k�ܲ���^�rU�G�p��A�@���5�ժJⲹ��W�^��EB?M8lX�Nec[��"�J�L�, _�����>�����9�X �!��}a��SL�3��PmrL�y�#U�h�� ��r�tW^�h"���"�a���W�G��S摢�E��^ .W�yE|ʸ�b�\əz�Fu�ا��CoUEE7��v��~��.#�f{�s��+�;%4����[5�|�z��l�J�A�hUql=Ce]MHx5�Ug�N	�ڂf᪰M~+�mQ�����o 3�DEN��3�����������\:�~�<�K���n��P|v�ar�0��t�[r7�XTߥ�hi��G*���ks+�г�y�<�h<{����f:���	_�7�S	-��:'p�r�G^\�nrB8��-��PL� � *HN����D/R5aOK�ʽo摆��uң~X�,��<�r�Aq,�[L�AA���]O�&��&,ݞ|b��~rN?QG�E'.ؠ�	o��'OX�ƅ�7����k�#�+B�J�2"���qY��"ɦ��"9��+�$����y�~�[�w� ��mf��7Q�,��|̴� �g�8�{B��b���6��񢹼T��<�n[��w��9(b9+oQ�{�R�=���｝Eز��L�|�>�����]�?���q��C)o6��vUf��q�����{����i[��d^l��-�K��joLK�6��	C�@-���RP�s��ӑ�8��5JC���}����������ፊ&D���g��pZy�Ǌt��B�l`��B���Wv�«-�R�0��hsc�F��y��tώh>I�����P���L�%�,�%yA��9�ek��e}�k�1��W8쎱��&�h]���^�?>�{����g�8Wu�|�����)���Qb��[x5�Xh?��HrB�mL��[���zs�\g~�Fڭ�c�WD�������`N:1�ǀ��Q{�뵯���{{�&|�=���+9��	�|j(�r��ܟ��.Lq�_\<��H�0.�/CK[�ʔ���AK�:>��L^�z�WN�9����A��|�y;oo�O/�p��%���dV�S�V�=�"�Hq��|A!@8�D����z��ܹ����ػ{�Cq��}��1�C�!�G�1��������\m��yg�I4eۻ�3ok�����F(
���7��{�K�acn�H�v��m�}8I�1�rpy�2S�"8�OZ����{aaz��yX���gs�i$��ݣ���",>B�@U%�8��[+=E�^�N#)�w�8�ۊ�A�usc3���')��^i���5�?�f^�ܛi �$� ����zq>�w�d$Rf����K}�/�s�yV����x��]$o�JRUjq�?��*�V����f �祝2[K^̮<�3�����)�a+������8 �q ���ܴ��˞J��4UT�0% �?� ��9����i�.N �r�𠡹˕�H�к67�x�>�n8b%	���O�l����@���TH�{����+?z��Z=����@��\�gŉ�ܯ#�W��Y�ϸH���H�|��e0zǔ��7������H��E��t�b��6��2�����z�G�Ŝm�
IV,@�R����DA�d�H��
��XU�׹Nˆ�T�s>F7�O� ���90�9�jm�����dm%�sС끷ŷ��x�(d���?���9}ҌK��l�9s
.�NTW��{���)��ċ�rUI5�Hz�M��*����v!�4wy�t|{z9�vK�MO�,` U;T��cë4&��g�����]h��-��Z��מY�'�JԠ-�c�^K�.?��'�n 4��&cy�ryu�_Za�`7�&X�I����F�O������� t��}���2�LjL� �HJC�,xM�q�{ ��*��zϩ99y+o�����8�{g}�,��}��*�颭����n�Y��:�"'�}��g�����(�_�������:�{�E�B�*e!LkrK2��I^�9:��nХ�k���^^D$#!�dX Q�I��G�ly�^��ʰ������l�̹���y
��S��*�&�̍��6��w�+����\��]�iT�7������ys/pl+�6�Z�Nl0'�`�8�vo:U����><8b���*��@	�n�x�^<��&�J❌��9�J�e}R�_W��ж#I~��/�g&m�V ���cw����,T�@�4H���yZh8RҼT�W�mt0�Fk�g���h)��(^��Z��`��>bZK��+*�DQ�ཱི$�p�G"	)�7e���"K�_������阦�c�SD]Ŕ_�%mU҅%/b,�"�9��}�Ԇ(�
�b�H����,A���O�W���x�}цk]%�F�yӄ/�?.��:.U�� 76 ��N�5~��b��06��0��}���tu�aLC62�/�%oN��aZ��;y�w'|"Y���"��rR;e3�G�y�$I�r��T~Ņ��m ��[G7@�����I���D�c��ڊ�?��E��,]{��B�;}t�`t��%����o�=��ɗK"�M��D���͞S�mx�Pt�*���������7 ],�R��%{jt�7 ��@�3/6+)lE)Ў�xu�&�l�e���j�!FKD:�&�B�u��D>���T��2,�U=c���Ҽ��b	����o�G�#΁���'O�܁�����`��"��Ǐ�����I��G�`Tf[x~ޗ.^dC�
�+t���a?|���)a�����{ɞ���4�Ѭ�$�N��>�0�� ���f���G���{7N���t�U�Yx�"�%��\S�ҋ�kp�c�Ti��<zb���(��@�X�բ0l��&����>`�.[)à�c�A�j���"	�S��t�h��Í�o0��,�`g�0�p�1�rY>xQQ���������F��)�Ig���*�|�b��� ����W�8���^_��:��k�b�\��ʌ�4�e�e'�EY���.�ް��6�a�p��K�v�W�/�rM�Zf`���*o�#b�k$�"b�6���q0���ؐ>7�J�R^��-|Χ��V�2��vrBIqny���4�����xT�C��i��aR�G�+�
�K�8im���zز���iM�.S���5���i�;;��@"�QxƐr̫�&4��/�}B�Wߡ&���^�Pe�@��^�գ:���a�T]/�����'<L'��t�h�,sq�J�~�^���Z���mQ��T�D�kS�+;HjƁ��D�/ͤ�������W��u��J}��ܓWu.�(������:}��=�&gd��jCC]�숮�������ߴ�wVŽ㞕 |���j ��m�P�g�/d߹s��{�]�0��ϕ�*MA�ܷ����'�|B�~�)K�0'lw��i�>�;Ipձ��i�Z[���kO"�M�����}����v�+G��JO�ޓg�6*A�s��8'�]�����Y�{�%=�P�$���c���b�y�^I��X����!��
aD�h(h,B\�P4z����gc�ҩ��j^^,�8?,
��tVy�rP�?�8EY77:�ro�=�>�����_C�|��
���ڳh[�`�|��<��6�oYUAQ����zёJc|Ѧh�4&�=%c�L5�&(-Ҭ�����Nڊ�{m��R��b�$�����ykթ�}� �����w��H"!�Zt,g}��ծɼ��K[�k�l�d��p�眏��|ĉ^-�O�:��g'xA��n�ư�!��L*�A2P �̉Xq^�*`L�8 ^��5���rIy�Ǌ�2_UZ5�S�h��y�%
-��Gk4j&�n��l����C��;����E'�ۜ���0~��e.)��̯Ix�5Ë���2�<���:���z�>�<��ʼ�����1���.sND��`[�u{Rƽ��Ή�����y�Pw
��jcQ���U��Z!��;2
D�.E�̳̟*�Tf;IND?F%���3Po���R������/����iXKv�9�mNgGz��f�P��a��1,��eN�+�3WO��N������B$�%'�r���� �"����sҦȑy�ߖ��K�I��fijgвP�<6��'����Z�{'�p*t��x��]��M��Dc�5�gʧ{uz�Q]��۾������Ԗa����՚�r�ta+ƒ�݂�G*5���U��t�"KXHi�C�_�����w$�
�d.�g���{��-���x��#���Ju~��?ii˖'p<+���'6�Q�Xx_fɯ�l��5�%�#�1��\��"�<��n�'-�ń�D�$�|�t+��s��ހ�;�_���|�ڳ��9�[k�%v6W���)	Y"]�/py�����%��#�e�0�"�c=���т0+B�\����1sA����{v��Ӄ��C�������g�'���>�:��k.����O�_gT���\�;�ȎC�DQsZ���ٮU~�|��imc�}�O���5Ȥ�rn����{Ϡ�֕���){�2�V�������W���_�o�1{W�y�mڀ�V��d�p�F�c��H��0����������3�7�(?|�%���ˀvƊ ����2hm�0N���xnN"(��ԕz�j�D ii-��q��_r׹��̬�7t7 ��"-˞c�I��<�����<�}�Ȳ��M�2A$v����%3&��DDfeu7HP�y)]U�ˍ�nߥX1�1f4M]��ȦȖ]ݓ`��j�T2?��s��5�g
e�A���Ǩ8���f ��޹M����w�8ny4�HLs�0�j� őa��WlQ�Lo��68�ߥ����QM%�"Cd�����}_7��ðcƞXt(�/Λ��{Q�X3`�:lS�:-Y�3�H1�:Ip.�Z�DQGb�øC9p�`A�
W�sm2ٌ U��\�O�%�N�N�;��Pb.�R]���W��О"%ZE��4�PN:(o���Wa�_Y�*i'�� ��Z9��-���G����_S�u�{��+>m*�Նo�Z��� �z� /�H��W��&�$K�1iP���E��Dc�n!���|������Saj�3���)�1��%���:m���{R�ڽ��'�M�$K6v�v�}��6�����CZޓ '�HQY�R9�q�' �ckk;n �� İ�4a�� �i�f3"���J�w�%����h/,���I)��h� �x!�K�L�,)*E�����s���O4�ZiU~�L�jo�A�b�c��:��T��-٪Z;�H A_��w�S�"0�3���Q�[즁dlm%����@#7[�����MF��o�>�!�E���,S>���~��Þ�i���Z�� Ws� �n̮�*��{�I{9�����#�uߛ'� ��^�?���L�<|D�߻O�l�"�g0z*G�u#����W^Q�/�ׅw!]`9���L�ϔ)���@�D�p~�r�Z=G�����|�cl���S�����H��{F+�Qca:��Y+��cV�K'P���y��+F�:<7�7x���ۧ�쌓� �P�f<�P��h>���EU���1��2k�o[[`x�3M�ʌ�^�U5R��0����iݐlg}*�S���9b��)�(��)xg!f��b.�M�]�u�P�)��:6H�5+���b�$�����(x��T�n�?��&4��o�Ե�D��+鶏G|�N���K ��l=�U��M���ù�-P��)L��HS���dK��r�;>k(^����e�6�ɽ�g��}<�h�
�W[�Y�x���.���[�@�S�ػB�B@�������� G��ڍ(=mP����o`��)��
���{�����&�0_���b��8�t2�kb�,�넗63��?��Ͽ�2l$ƃ��!�c�!��̀�^ķ��JJYJ��L�-,�>��o!&:`y�d�

�{�au}�����F���/ڋޑ����Y����`^�U�D��L��t�%K�M��dA�N����\qJ�'��<��j��g�bз��Z��:<�p��NZu���\��/q�!Hwz����.wW�ǎ���dmy��K닏���[�_���`o����dF_���e�f�4뤭����4����������xؚ*9~��jοf�|�| ��A
�J%�m�"�X*ݢP �Ş=$`W��R4��\�sV
�h m������E�XX�x&�Lf\q.�%�ꂋ�p�p$���M���(;�����r6����g�~D[�F+�KM���?	2x����//y�/��8�~�C�6��g�-Y+�����Dkk^f��#��}4R�N����M��ך-���R^���%�� Q�t�O�k �:	2�v
�\�?ư�ܹ�"�^�X<�g�Z�8��aӉ-��p@5��0t��r�+~��쳀]�3�[�����n�)���Ah���eڋ�S�5���;!ys��D�[H)��&�j�~������ж3����ŉ�~gg��O�*Sh�Q�<�61��]�e^g���Ů����"�=�KM�p���D�
t������]饖�Ţ��3
�"�ơ�G$lW�Y6�g�}��3t6�:t~~ѕ�1��3����,�Wm@I��_��/�g��N��U@g7u����|�˱�� �͌)Bjb˺�J{��e�Ꚉ酅���V��]n''G\$ьk� �[���{�>��>��S.qy|r�� {6�G�>�:�/^<g������梴�ܝ��(�lV�-OX�jDaS����-���4�8ϝ|�L�T���j��3/ݢF�/�� �P:������eXåP� ���:�`�O��8,a�����1sk���-�4��P��|TF�})IR�������e����uzN^�����5�s���_��튗oˊ|�ø�y�j��d���,9-��Z��ܒ+�`�h�5��"��r?�����V�+�]�׍�B{	љ���L��E�E�+[�L���^��i,,�c�1�A�")4R�RI��MEV������s)m���Ԗq�I�Dà�i֪2���g?K[%�b�v�����Ɋdp_������6�7��!`��
��0���рs�����Q.�ѡ�>G��8����&MF[4�9@��`k� �QA�2��R��(7�i(d4$pg��\�X�%	��w>%w\�ڵ )��^Cn��ֳ0�nThf�z����,����+kV�P6B�e�+Ϟ;����u։�2�T�����p�p�4�!��W�����(	w�0��wmN�&�s�*^���W�� �K`2��3�E�Uu��+=�'���4���?k��&H��ا�;p8�|��q=���Ą4L�Z��:̜�\��vW��p��!�� X�"@�u!vF��%�0,8�i��q�'�" �{h���c�b��v:xĴ&� u�9]��k&q�R�u�XLh/�v:7\� _./�F�{�����v'��&���I�R�s�=�k}$k��\�4�C_EW��S�B�5�I�4���^'I��q8�(�� �1��C&28+���ioo�A/�@`��;>GR�����ۧ�w��G~̌O�>a����`
�l��6�2�t_,�	j��'D�gVA(YU��iTwAW���[�Zt�^_>%0 S/i��M1��r�fy�T�g��?�(���(˥���t���X+'��bQN�1��Q��rs#+������t�7>Z
�_��
���o����$�z��4�H%��Dp� �5��%�q̮�1t�y��e	�7�)���N�j����JrDb���&��j-�.E���܎�B�d�b����0\�H����l)+b�6��)�L��ɔ"�KM�+#cG��9്�fpU�܈m����ZW�*��,&]Z�%o�����8�2bQ��UI[�{��ih��[���ሆՈC��7��V�\yh%�Z�J��*3d2.����=�_C�?ۼō�E��������|�O����|`�^.�^��f��X�M�U��6�O���<?�4v��� l�7jC�!,�\<R�l�%�WEE�N���k�̏�?��VR���*٩����,��
xKIXs#1��ޞU�m���"�]2 ��b�ꈖ�:0��p��5���qg`�r��z d/�4�^�@{�=J��&A��M���8L�	�QA�]t��sLԜ�pSmv���hf� ޠyL6����`��y~@r ��S:������N�O����._���2�{!��3�Lj�ȹ����-�ڂ�k�O+V�֛o��P�85�j��ĈZLPî������hh�q@�3Tt����Q4�-��77�h{k��.(�>��S��㏸-��E������p�Ӄ������=��:��[f��ˋ^E���
� ��.CP��ůY�o������%ہ**6/2 �c�QYg�jB��f��x�HdJ�	q�Z���D��Y���O��X�������qb'��J�oa������8�ҳ�k�q��h|?�����^g��n�b}M �G�Mw����F�5uŒ�?˪E�fk��,��fLA����<f7g�x���oY!���n�Ħ´�e�����'OBI&�6CS`��hj���*�^��5.�D.ȉU$Zzcx���$L�����33�Q7R��������]��V,�2o,a���D1����2J��$צa�(39Kff��J�a����2'
[4��7�X
Qʾ�y��T��2�WS��B���\k�%)�ƒ8Uj�M���Ĕ�v7����!�P�ux�F��Ē��+b����ba�[�,DFR���5f1���%��_J�
��R��Yy�1��i�Q��׺��O�#�;���4��@R���y5�1�yZZK��=������(����(;ɚ`�����`5���u٦ɛ\��fY�$o���	P�Jm<�M���K�,�s�g�����a�SQO�k;|� .���n
�}): ,�ќJT���¸O �|!�a
o����$�cй��y�X�=�64����Â;���m����Χ�"�a:�:�r�@��_o}��aM�ݬ+��ֻ}eT�=C����ӆ`�������K���4�a�znt�Ħ�8�B�R>D����� �"37I��1�nC}�b�u>�gA�B>��s��{�����7������~���� ����7r����[o-2<;b���&��C����WCH<?��%a@�Ap�J3 �ZBq�p\'���16��X�K	��$Y��'}���΄�x���f�� �1l�D��"�E�k�ψ��=V�Zrdv�V)�)�,��,W��Б,��R�׎Yw�.����[RV�Ţ�kْ�Z듻O�
r��u�rݥ,�˔��&m��U�bo��M��:�s1S�[�+'�%�E��2�ߚ�֬��V��r�oq��놆t�_�{���ٮ{��&�n7�_���i�u;���F%9Ad�
S{7�0���40�F�HE���Oe~׵5�w�ٺ�<k�YO�f�%�Ȏ(���d�$�4���$�k�c9��P�̩N�
��xbQ��<�!��6���P�	�LKe]h2�U�Lk���k�X9�1Ņc^K:�&��"](����1�l8���H �a?o����+�|vCo��E�	��7�<i3&l��\k(�b�!3��#��EhIa��#<�2�����^��@}��� {	?s�&�W�&�>hL�`�-�Z9���>R`�� �a���w����-Y�4�"A	�w&����g�_�I�ʻ�j'��/�(Qʙt��2 �.WdZ�� 6A�: |<#C/L&��Y �~'�n��w�	B�F��&b�P`V��]�������P�!�,� �x�L���m@�=
�`�"�af_�՜��U��i#��,��dzLg�ih�B���O#��jM��{�	�b��h)�D��;oY�+�yL�ا;��f�t��'��I��i5� j[0�r�)\[Y�J�"2WP���*�2W���8lĪ���s<.������=�{�V�{����O��;����K�;�ܡw(���9��\����v�T!�o�#�G?b �XJҎ��-4n9ʔ,�20�i��S� m��\�"S'����"��[�I��	%�|�Z���L��1�Έ2�����M�2}%�<�g�.U�YG�e�J2#ݧ+�ޒAP�c��vS*ZZ�kkN�4��Z�Tr.�o
��_wF��M���n�M+��	��J2@�+�\p�h)����ch����n5¼8K�5�P���	�]�\��=|=+twͭ�JE��'�2�M�;.�b�:���y;�0k�j[S��?���Y]l����Q���;��&�;HcT��+!��+�#�j<p�XXk��S���$R�ҵ\�׷q��J!P�%)���$�а�:�g�7���	�,�M-����`=���C����b�@/����nb�TᲽ����8uM|�����Dcl, inY��3CUY��0A
y�!	V4�|*?��%��� '��4��<��#g�T�����vh�1�s��'�I�F(>iO�>�S>��lO�?D�@�,
��L5Om[<?��t9���s~I�n��	�4#@(^ ��Iؤ�;mʻ�U6���8�:��&qh)Cvm�N�������֬'q��[fB��M341��6MFg5n�ƴ9?	���^��E=�E �r0������:��3�����@h{��U��숮p&�� W���2��֯�Mf��"6�"ƈ��8���1I�gm�3�;::�����_0�;b|Q���>㒜�o�fk,>|��#�w����2��e�fX;�ԊQ�l�*������L����,��A�4�"���Q�K��XfG����a�=�'���2@��_楔s��g�
\�y�)��Z�W� �Y���f��K�2Rޝ������YaS0hs܌ڇ��T�Z[ژb#1��&�	x�wY�ل�@����Z2�u��฼4w�]�v���omnv�Uܟi����D�Y~��rԉ	`VJ8a2]�$�2sR�����դ0`�;>]�6r��"{��T�4���}�A1Pfq!�Y����4�/��=A�H�"ư��T���0؄�/�E�v�FVy�Si��������7|�XB�^��e
VM^3��|���4����Zk+I���o�B��z3Z�3k��Z�um6^Y�n�5������O��ȭ68GJ�5d�k9�RƉhs��\HXI�ƴD����(<蘙\�ݐ-3n�f~7�s<�H�ٲ�.sR-��5�o +�	���K=?��$) ��V�)ݰ%�܁���
%�{v�]MnP1|I��Gtzq,�f>�%4Q?Dy;ҦPL,�:ә�FVǹ�ӻ7����7�+��[�o����f~�@���6��l�oOv��b�4����HyZ����;�&sOnp}��2(�ZE�8���?|�!V-���/(�$����u.�<�.����m�>���Wj.>�+KF��Ԗ1s^t�3���|$mP�:�>k_��K	,mB���k��9���י_���w��4�rS��u2��nw_��A���s��YF��QQ����:OA����	�ߧ1-��V��-r�&)Ex7������r�]�h���F�R���6������8�o�}��w�+_�y}w������YC0[a}v��=\�8�-Ιs)����3�1��W �z��K�5-��6,���s;�R`��7���>��s	�C� �F''^	��#�M-�w�� H�n���!��.��l�^Y?��#���j���Z`=����c��՗�AS�2N2�3d��(ǃݼ#����e�j(,aapE�J����t�k���x�#��@����8h�>vS�y߫�d<�`w����b��@��� ��tt�I^q�I�x7$�	�" /ճ�:`�$��o��M�l���fƯ�����^�v��ϧF�H�l ��(L΋Іy�=��&����D�cC��&[7hr����M�g�
��Z���x[0Ӛ����!�H�x��*)s�%��������o�L8�du�,��U�~J����m`��Q���VLw�@�k������I��k�o�bw�, De%g
�{~>��/�1��'�������}�@�.����N-�q���.���Lߺi���'�1�yAk�DW��Uc��6 ���F�#��*_� ����}1�[���������-���7���������^:�>)��m ���Ɓ�)h����"O��ﾣ�/��b�����r�P��o�P~ �lg�|{�j�5��TN�
�F�J$�d{&+B��*�Y(�]C�U��ټ��v����[}��k{O�/��Z(�w_R�ۛ�*��5��uZ�~��sd�׵~/e����� ���BA�;������^+�W�oh�77P� �ԄxP�B~lLfAl��lB�e؟89~��KP�������^R'��ӗ�^bq�ȫi�|t��'��Tb(M��{��
}�9��A8��$�s�4xj�u��/�I���KGҿ�T7@,���a0V+">��G ��N/���#�~m�E�t�5�;�l�Aq�0�ƲY�$,�h���2�jd<�.�&m�w�q���1׻���"��bI�qE�ixM�Pi�W�f�!T17�Y�����|v&0��$��?����yG��*�-*��LC�,խ&���xs��7�(�wp��O_�)�WX T\�������8�<Ao�7��]����!o�-l]/m�i�¯?��Pp:๕�kucAU�bQn�j�����>��'��?��>����vvv�Je#�l��b:���#a���z��W����𵔹Uˮi�Δ��{��nq�)�A긣�Y�l,��U��PT�⪅���Y[����"��;\L��B�F�uQyӨ�e�����iE'�F5wt�ǹйԏ v�~��o�>����j�z� 6����>����E��ӓ3.�[B#����0���*�9���Xh�6���6Z`�ֲ�H �g��Ǻ�N+��X�>kG���C�]7�x�5_]�M9��%�����ڇ��￀��XGϣ��Hb@�$O�Y&���.�tFy�,"����5��vר�c���%�4n�`��@���Q�`F]
�Xp�x	W0o���Q#��6y'%!�XT�Qr[Z`5ӫ:�䚥�L��[������a�V�s�HDMB�-9��|��m/[���j0��CLt7+t,��9cN�}��&!wmq{Ś�Ñ;H>���G3��6��Iʠ!����m��U �%���\ ����h	]#hVΉ𻙸x=�i# ދ	�ÖJ�]�T���N$S5 ҵ,�Ve�坆��ΦGt~vĕQ���L���r)�фƓ4�ا�� nkZ�k�R�eH�1\�N������vq�8@��B3��[Py��Zs�S+��\���T��k��=[��	�|����\u�P�0}��鳨�E+j��_�g���%�ψ�vQx�W������]�`�+m��Q��Yo�R�������W%''Ǒn���+�����l�JSt-��!iW6�U�J��w�>�MꌖW�h�F�ǠQ�p,�e�J�ѻp_8�yF���.	�tx]��e� �Y�z�}鑃�5��g:Z+�K�Z�E5wY�A��1{�G|��9�Gc���N �ѷ����	Y|tYX񐤠�����/}VI��4+uW�vG"aD�n���ě�Y6r�05Hw��
UV�\���
 4�c�d�[�"ɼ>���Ic�(�W�H�mnӾ��V�ū�������:����=zL��Y����,�v���$��<5/�l�
n��]~;N�ʕ0kZ4I��H /8G�IX;ޓ�`U%Wꥱ��Op��"yy�hF!g��
�X|�Wo�1J�nw�\6�h5�>�,w(yk��N��Zn�J��%� �^�k�*�e�\�1=-� 9�w���ږ ��y������l��,Z��P��FF_�C��J��UXm��z�Vy�\��\�l�����^r#׳�d��� �u��
���G��a�<��YA��XQ+7�NY^�lz�[p���A唓t{g�͈�<x�ڞsX�_3����e$�$������l��|Jtr4���.�@̱��&���|L�߹Kw�}�v�n ����'��&0�i�FɕA�sp����\A��?hϘ��7Ye��Aێ�>�D.�#[��}[���VA��\�?�y8�w5�L
6G,��2��R�i����
�:��,Epmo�Ї~D�7K����{�K�n���	˙�u���l��~h׽��r�  ����w����Á�qk6~Z���+m���e�R�ڹԲ��`�BO�)$��Ʋ�uڂì�HybV�i��b��Y��^;�̞�P��6j��@(k�#�^dՇD+mq�2=LY���sX^θ{��Hs5Y��d3|�ںk����}P�ϳ��Gx��?�?I����x�
��ވG�� |a9�u��
�Q�&kaN��4�ھYo�L�oc�w��U"�g�y����{a(y�K쮴mZ�����t�y��l�x_����{gq��˦��aQ)Ģи��J�,�Q�\&�ԕY������GGJg8�X@uᚂ��p�6���W-񴲆����\�/u�ʃu�zW�
e�]mѵڴ����:�~��
u��L�z��r�k˙�b�i�Ju�K�s�0��3�aXH�=�m �a������%�%9�fJM�߰��'�*u�a�p�U�-�'��*s$8���4%�cQ�^h� ��5Y�X1���F���+N��a��V�0��r��ổ���	�yݩP%T�Ъ�o�eO���)�|�E����s��s$�q�0�u:����/�{��Y+Je���S��Dte��ݡ�zP:"\�u#1l�@�%d@�e�a�%w>����XM�1�~9
ߗbمU�k�r6��y ��g4=�2`F9�� ��a�'[4^V�`�������υR�՜���fZ`��ژ	�㋕� �!�bJa#<=m��洘a�F���!��pHDSσv�1�\�b���s�������!���ѹ��ÂpJS�*�l)���%]���.i��]��]�r�l�V05)�G�Uu6y�����Eh����'@�8Od���,���7o�������_���/�����ի�\����璿Z�	�1�w���isc�c+��_�=P�`�M��6�NH�#Y�rr��K�,��h-+��o,�+?�M6m$B�U+�[
�@h�M�h<E �mo?:���+[	Ș�>�)�?4m(\r�w-�Fٶ2���,�o�]|- ��3p����p|�:�8ŠV�icB���=�	��w�Іw�O޽w���}.n2�8����T-P�|K)���&mC�U5U�Zi����T�5���p�G@��k��R6n3�T�U�*ԕ�����.�I��fq�,�ͼ� ��dk������;o_L�7Ԅ`;��[��V����j�B���:���D/���2��9}F�(����Jz���*�|�;�?�/���w��ކ5���E��^'�+Y�j��9�-/�$���c1�Z���-����ZBtw�k�E牭�h$$RyX���=���c.�#�1���=݊*���Z�U���ۧ���$x�ú�[:�/뭯������2�`�J��(J��2P����]���*�Y؏���Ý5&3�0߅#J�$�yhH�Yyw#�w�g6�Kcx�y����^�׈  b���L�.,И�.|^0Э��2,@
�k8g>[���1�x �I �缑�(?F����xc�&a#�@�B�+�m���0� |u���_�7�}+�?4��KBE���Ї��Tt�������x�e��b����56i>��K����&�۴��ĵ���dz�FF�ω��PG�w�����v�5�I���[�� x�U��&y!�W.B�@b�	�.`��C���5PK�V�no�]����o��7L10q�Ybs��G�|C�?�]��3v,!�Ԇ߽s�~�3�c�F�⦩4z��4�#��ՍW���j���B(��Wc�zn�� 7QJ�+��G�UW��XZ�d��]>Z�縤	Ev/��G`��*m��ڴ渮%�m�E��_���,�9G,^�o��%Ӌ)�# �_TK�d��x��]��_��~��?��?x���qܺy��{ﲥw@/��˗�-�6�S(_�~n����̈-/��Q��º�eo�*'�,��
�X5�{�V^�TwX�x֝{4��zL_���B�c���xP�Z��_���}��5���
@�SP�)¬�*hg��*(�E� �������˗/�^cV-��.)��m��`�$��{��:�ǒ���ߵ>�V����u�tU0l4�R��@�b2�a��@+�൬��!��}�a8��yd��|�`��Ċz��R�l�h�{�,�vq�q� j��m/�O���l��2�Abn7����f�!\C�6�x]J��	�\�R����"I�$e�[���=�ϱ�3�^��p�����P����5`ϕ��M�D�mJ]�*�|�Z���Z�  !�8z`���El�0�[B�eE�"h�g'��ҫ篹�0�'�d�GS����CB$�2b}ga��Z����`n���u �(^:p��$\��ᤤ�"�Y�n�Z�NV��1f�p�����ه��2TS�p��moܦ[7^���h~q��s��U�\:�wmQF��=�����8/������{U>�:�Bk�n�P*�-�{��Osh�"�YEx%��U�ޤ?��JH�.ѳg��/�����I�=���Cfq�� ^z��*��ۣ���������7��w����ɓ�ۋ'Z�+gг���!�H,�� �Smղym�m�cޟ�ϳ����ì��AL���0���W��7��?��ɳMs]�%뛮��*��&V�7=����ȋwt�>��2m{k������y�5Y�`]#���s<��׿�9�2��}�-��0�P�������D���Bb�Vq@Y{����"YG]k�>�������ً�d�<�A�I����|)��QlC���18���^#���VPF�|�)m��ҿ������wtpp���m����%k�������,78V��|E	��Z���U�h��C̶�1N��|����h��>g9�����3��}ߣ?��z׾��������j�����i��}.�V�-�E](T�ټvjP��\��*L��@UL�?�}SZ�T�tY2�"�/��ш�^6���ʷ��r/�16IB2��b�ry��9��;�<o5����;$�7����\�.֛��^��x�q�a)��K��r٘qY_��9*	��QAo�<C�2 ����z�po���E�yםlaxk?��Yr}l�;tx��" xXF,|9�&b$��<��/^ӫWb�'�͐�KB��R* �-|?OggS��^p��*��R-�|4K�4z��a�(P���w�x� \���i��FK�4�0��k:9:搋2���w ً���6i#l�[��T��~B''t�1��i��1;��Ԟ;�F��`�Jm^SE�wO���
e�TB��n���bi*�X8�Us�X����g��~�>��Cfb�P�pO$���-��oG�yH�q%��u����t3 \Xsa1�(�����O>�����? �C�g'l�/T���6�s,J�����-Ϧ,!�Zj��\�p�ߧ��gex3�(Ib:Į4�qp��a��1���Ǿ�� ���]�Pe�rvȇ��c� ]?��',�i�ql���bcÜ������k�����*�!����K7o�����K:	��^5����V��*v���ׯ�"��A��ba�G\S�U�jY2�D{>��_�֙b�l4���{��9�'�jB��m��p����ޫ���B�Ƙ��o~N���� ��g�M���A^���:V!�uWb���\�t��6�$�W='�x�@�Y` ኆ�����s�9z��hC(%�ǣ�	B/�+a�Xyϧrn�k���F���ǥ短<���z�%y,v~t����X��CB��}�������-����IX�$\Yщ�b��|:)M�񮗷St8t6_���b��bHMn^e�K.�XB��̻x��X9f��H�u������U�In�ӗq�k�ޣT��[�34�mrHJ
X���m!q����^.����Xh���z��5�Ќ*��Ғ���z�M��Μ�.3*�4Q\�B��>��u�$�W-�v���X'h~3	�=�J&a"�����G����|	�y��W���0*���9�+W7�y�D5��n� �N�żf�hЗ-q �a���o�[��~���a�z�������e-�t����6�y�lR�I=�a=ܥ퍰An�2�)*�.�F�*�])PS�[,���~r��%Q�_�`��-���G��)�[u�����N����)���
ZR��B61�@I`��=^�xA�>����� VOy�0�
,ȕj�^�W�ѽ|��-��ۿ�V�ͭM��¿a� Y�K�������f�
� ��n��-h�fG�b�yh�iC���N�.���{�V��bԸ��|����*9�bW���@�u�~�a��g��he�MH%���GϞ>��?x�����O�s�鳧\�fk{���0��wo�:d+�����_�n��vP�~�WD�P�TyzB��~��]::>�� �?��?�}I#$?��QWH[�8��L �C�F����;7vxM�Tƻ��s���oZ5d	`���#z�ރ �7�
�4�)`=�~O�)5�7��4m<.�5Q��Νw�wZ�>�s�*M(�*�X{�a-��?��3�+��x����?�3+(�GG�6'z雊�վ����Wz���������Z���Uw��]3��j�������='����u��sD�o�k��1��Ea��g��b�v�f�2OC$�ʵ��]��'�����sx�\�w6�b�N�[X8���OO�e�s�@��˵*mRiT�HL{0=��1�VB1m��3�x8�F��s�q�rؐ���~ ̯�>j/�
T^�W���� �����}bt��AwNH�����������,�iZ�{M�}���-���������+�L��)��3Oc�B�N��_��&�`Z/�d� ��m�[lqlbfJ�B���_ҫttxΓ�9 ^!Dn�X��j/2�&Z~ǋ�I.�܊G�0P�X5�W���sΗ��ϡ(����>|>���(�fƱm`��9����<#*�C�dc5nm�q ��{t|:�i8g9�Q5��ZB��t�th���^����oܓ`��r�.��\�[cLH���F�x�"ϟ��ꢗE��y�d܀L}6} K� `���<�^����L�YJ�F��sjٙ��4lv�&`�r�;�І"x���u�wߊ1Y5
���4n�A�BPQ5u�z&��	����Cr+K�Z�'� �6��meǧ����5آ��um�1�\z�,?��z �s�4R�k�)-d֟}���`m�Z��v��.�(��W�h����s�*
����<��/����"��<z��cZ�]����0ᵭyN�P���!�����T���h�J;����e?ɫ�a}�6#6��}��gS�M�%oc�\�
r
_���뇴���Q���p��ǼoHG��� pfT��yCݐ(��{��л����I��<	�mXAF(�e�bi�����m�����r��������6�e���H�dq�9�M/j˰y��*��t�Udv׃}�{C�>p�3��y���K�oD��b��m�23��+>v���/}��=`0���^�5Ԓi{��|c��t1c5P ��֒B����9O���]�aSꌿ<�jNL��}���s���,LU�1V�C�U:i�y>@��r�v�B�PW�e+���c��HO��J��s��0�)1�vp~3�첗m9����3A)gQ�}�:����>��N�W)qS�������)KE���teA9պ�&e���7�-����D���ײgm���B�A�@ �̵K�37����BF�N��V��С�:Mi ������K:<8:UB�e@�&ֈ^8JZ^!��`�O�gm�sm�
�q���|Q�h��q��J�$&$��S	�H��={y@����1�6m�I�5��!J6z��Nd��l~���K�}Ù�V����u(|�o�m����O��:�"�2-K�,�L���sܑ�E����`8\���s��P�Y|62�Zc�����6d\WA��T,H(_
vQb���F�HX�ׄ��Y��̳J�ֵE��l.�-^�e��jI���8>�ڠ/g��wq��ꦕ��������/�7%e2�f�oJf��qY�����f¯�w�U��;Yy�7�N�VnA�X���ի6��s��=Mgo� o�� e���?����ߧO>��f�Ԁ�[
T��|>eʮG�<�����<��9���h���[/���<7�u�1��<|�
��{��;wnse�d���q����m� Dj���`���ڕ�7Ϟ��l�ceϘ?�NQ�L§�ĕ�����*�0+�����3 ��yh�SV:.�/�J�r��Z���K����Vw�Ub0(i�1��/��o��o=�����( ��"<�Н�7ْ���GO�~~�0��]:��Xɸ�{��{���J���p�͂D{�ݼ�(�x�(�H�)<�B)�^���`���\ne^U���Z��0#9��ڄ�X���o:��Jo2&y~Ē�s��0?�3(�����xlL6Yi1�?p�K�F,��!�@z}nq�� q�A�\�,�eT�"���'��6��B�����c����DPxp&4Z`�-)�b�����;�l�yyK=����u���.c��5����j�¦P��r��'�G���)xd�-n��5��+�8e���s��lm��l;��8�hEl%/'�Z`���ܲ0�ZxIiw#i�D�0$g�"� �x���T���u�;Oq����+���k��չ�׺�ZR�FA6�?��{m������;mp����dz|D�wx�m 8冀E�mxJY��@� vU)�v��$�@���17~�@w���%��Ii��%�5ى4���UH}gPM�sz�|N[�����һT�m-nJ��8�� 0�h�����N�IU�Iu��R�RM��O߿�qH�2
��)�+Er�,���|�X�0u��k.[W�r�YZ��,$��)u,�v�Q�x�h��`E���,lq��e@0c׻�S/��eٰƈ�`{gg�)��+tfKv����Cڶ�t�>��M�Ƭ
+�-_�o~��0[����Z�Ɇܧu��m���6mc�/��&
Z���s_�Ly�t7�˺{�u�R��\7e��~��p��>M�c��'�0 |��9��>yB��Ｙ�����C �O��K.�~p~�m�5��y��:����Ɉ�l�h���@��[�"��;��p<�_���*�b�\2Ѕ�W8�]THkЯ-e}&P$|��~��)[{OO�Fs��o8���.>��?�3��4�pN{	q�v�s~b��AH�X�G�l�~����]�us�vo z@�=~ �c��	� d��dB��>�0��y*��J���bs���+\Չ+9O|������g�s���uV�u�	���lVk3��Lo&�<���{���Ri	�}ʯ��-�A�3wuS����'b�چ |̆*L.�ـECer��n��r����C�':}�h1�~fs"����m��[{�P#�7vo
�S��'/�#��ꗶgrl.�Z�H�٪2�8\�J�r�k|T�!���(����e�T�XV�h5��� �	9WZ(��֛ŚS�T�h�̴N.����ձ���b�W�3�+q�Uf��_t@E[��Jݛ.r٦�)j*��
�,��M�����E��%:U���a�"�����AX/8��`b��5��R{���ŭ���q2�EC~k��SB��袘F#����4�x�����9Xъ8���B �	={�����{hb�76�׃�{L��6wϻC��sfBn.f�܎�)��F]$�It��B��9J��\\ 	�֤�#GI����8��6��!B�7��W�x0i}�˕ӝe�Z[��ThS�4�0c%ѿC�U�F�������}L|��Wxpp̖����@X,uSoxSD�W���ŋM\�g��q����,vـ�B9�L�s�^˄w�"��9�mj�9�6Fי'���JeB2�Kf�E%� ����
Z|��Gn��-\����} ���4^�/��"���?��g���k�C�p�x�,���������$W��#y���t�1��Ot�Ih�o�F!lXl�*JB"�G8���١U�<�<T2F�-ŀ���S�H���XTQr����.��R+���� b\�( ][;8����g	D��wm^�$$�b������>�B	7�8qn01��Ya�����$共;|} �#�6on�0��g�~�`/����{V���8;4� ͮ�ÔE�N�x���Z|���������[;�x%�3��p�f�/&���=�h��B�񭄪�9s+/��q�a�/.E(d�f+n��=��O1SB)�tL+xʀ�U1��J�o܊EU0��V5�tm0��?Q�Ʊ�� &��R�0�����jǂ˳�h�,���g�7�+�6êhU�Y #B�?m�(o�뼊�L!��F��yM盆M%�[��|拶Q�բp��v�~�,�1�&T;���軥�e�J�Dg��4��ú;�
c�`�m�o�{ ����q����Kz��8-T6�M���c�Uʇ&]5��D/���v �A(�)+��	���3�#>��� �0񸠁�[��]v�q��H����ݨ�'����������'�h�G���A[�{4�[�h&�����,^I�Qy�^W�Z�,2z��V��TA�I�U1,�T9�J�I��M�-�a��.�t~6�x��xH�͉��1�Ԕ,�� �I�GkUa���q�◻�a+���	[u���e�|šUpk�1 ��n�۷8~�=����a�Ǝ"H|Cf9 �2�)l�ՏK�%:��wύB=�8�z;G�+�f'V
qu���ȋi�m6�?�@��jTw��}V��R�u��%�Cβ<�p6�s�o��x�	�HfÜC��o�/��i�&[�i��.�~g��{������.]Xq�(�GG�0��<?���Ã׬��Xx��hۆ��É{PJf�%K�B�*>q{g��H��
���<�d�c���Bb]%�u�����kd���/��j2��hp���6�ܸ��I	��>B�� p�xǄF�1���/��U�������lA�G'ttxD�^�&��?�0��6�*�չ�[����<S���Ρ�`͒g�1�ɺ0�z��qȺ���K����:_9KgU�(�7X\����2`���9O�Q]7�|��6[�)��y��`��.����Ӓ�*Ps� ��\YD��='ѫ5T�[�=*7�������(��t���V�d;�
[�Y>�?c�;ᵯ9�����+Xu���F/�8�pP��2,
�s�e25��࿖�鸯XX�����l�ힹEv�Ѫ1�����]���Ik,��^cVO�3~ԫ9�o��-a`h�8��ơW����n�h �ǂ�9C���<yA�N��h�M&�_�Rz��Y%���Ixm�;~k�%D |x�r���[؂
ˈp�9��a>����e����ס:
 �ĕ)5�%r��M��1@Dl@#�����g�6� �A����&v3@��X#T|9�3�5��%K^s�����mF1N�1�B0���*h]����E�����y@ ���8YX�Q�?w��:�6�>T0-9�����P<{����	֊�>��C`B|��_�`\jv96g������~�L��t�ܲ��}��	��	lI{��˶ 6��2Ua�$��T`7�|p�@�*&(l*�d�tt90Ϳ�k����i 7?d�)�<��
�8��'��;�����Y����w����� Ɗ��AE��X i���!5��}[�3�����2(��=~F_~�=}�< ��פ�v���)����<����B�jL(���M~���- n3���Xg�`���_)��X�ׯY&=��-��,�Xyɬ�M6�Nk���Wv�=�o����K.b:G܎����E_1g��s��wo��֍�Wѿ�����O�����x Ю������D�"��_��>�ʃ���e5���-�G��� onu��b�w�ʧ�5٬��>h�b�]k����;�E/RnL���-�}.�π��{������9_b�F*��i�2bMqYw�NE]f���%q���17 �
�R�	=ef	m,AL�?_J����Yi����Ȫ!}�n��(�����3�`Gp
�R��W/���Y̻�G�u����0/7�2�=����4t�B8������@�o�9��ot=|�&���VN�m���^�9-a���_^�����` F��P(�[���
B,\���4l8� {M�s�������5�J�)�䋪`��2ЕD�jP���@�M<��f���`��+ n59��lM���@E4��\Z��S ��&>���=O��ų����F �Z�ƶ��s�rrXh���G�zt��N�No>*8z�Yk�4��R���y�MB?o�A�T�n�?i����ŠZ�Ku�Ū3>�� �R�(���;�(`���o��<�p}b�>9=��1� �����?f�'�B�>}�E+�>}*�La<�N(��%��&b��WmY�,�!nR����/�����[A�{t��]ː��Y�N�*�����۳�EƊ	\���od���q���ڂo�X7���<3T�b�F��!W]{������`J,�`}�u�ݻ�y�~ �{�h�� ��c/�A����2�B�����W���t9 �MJe��ZXd$�q3<�l�r����,�*��Rir䥝Xs�S�7�`��Ł���;bf%�,��~�3�W2/%�'��kQB�����d;v�E���Pp{&�u�[1� � F��������\��x�Yx�k�ց��搅tg�z8�BZ}�ӎ��}sz�L�ח%�怽���{`\�=��2�`z�}����L��Kއ{B���QPj���d��5d<^���61�H�i�ĮZ15�.�����bhm�L�,���o����V6�q�%��:&�Q+�C���p��Vh��4��W����Y`UfŸc�1�X�&�Q�3k<iEH�c�"��U6�i���8otp��,��k�?%��ʦ۳i�D�۷Uu�Qc��b� ܱ�1�#6��4*���n.��$���#:=�rlf��$A�;C�?-�,�u�Ԃ�0�sN髈�bC�.gc�w[*�p���plr�Ц�$�ق�{�ҐA��r�:-b�,�,�\ͮ���I ��la3ӲDxŀ�Mf�xP�E��s6*@/�y��K�ނ��p��m~Fg�Se�d�I�1���B[E��
T1�>c!�K���ߌ����Gi��Q�G��/�����wp�������^E�a��k��p�n��
I6�*�ꫯ�"�����O��N�>�I�1M��<�~o�u�
+��OX��a�o�lI�	X�w<S�O�͔H�J&�۵Z]՞um4P�?�����n�}6��Wn[f+X���	={��y��8	Jd��N�����ؙp������g�x�;��&p�9����.�{�ަG�l	U��D&�d���*���+ɛ47���F,4����#L��tN�'b���Rj���v'\�\��A�l���b�-�K6X}�EG����j$�M��CVD�0P���s(��}�����]��IO���5� ��	͹���"���93���ۼ I�``�19�3�sρdt��nv䞰>ِ�����{w�tc~�9\[�k���d�۵�\-��Pfˁțӕ#��[Uy����T~�*ޫ第��r���׭v����)��E�o��|v}���q����뤮ʚ���8�&��*v��j,	̮%��u-d��^R@�t�6y�@���c�b��1I��7�̾��g�kf�G���R��Yd�EP�G7��xzˬ�4�&�i8��\�Av�'��5Q3�2�����G�a5@Z=`�^=���6�Fb���k4d��ױ源?�N��Ƌi�M%���h'�)P��/�N,��R�5<ST��xC�o�}ˍ��\���tR�
�F�	"�B;ے��؝�~Ya��r�Y���G4D��$��7���%f�\rJ���)�*-�[(}P�Km�`k�Tۃb`�8���l���Y�0��{��cSBl�\]���fT!fP�6�%�V�dQƹ%n�"f�b��&|xx@����$�!���|�%�n�����u�V;E[����������~���g+/��VZU*��X����2[֍�-�/���.lN�[�F��W��}�2�ii7yF����1-�0Z}4������m����,���A�vw9>���p߽n�q]P޲&e���ڍ���W���%�"�Ed�c9��� X�[�O�hzv�~&nx���E��܁��a� ��w8+��H���X��T��x�:�[^���ߤ�+u����'j,΍���ek�0��B˼�c.�V��8�uw�ch�O����̢K+���1R/�x)�vR�K�%*�A�4/� 5h�d}!A	��&�Nذ���j����d%��V֍��!4��n��U`�*�S�"�7m]Ew�z���u������͂j�R�d-������Y�k��>���51g���A)�*�z�п��#�bs�H����E������Ê��9�G�ZA�<FC*��F����-7�D��b�]�_��8W���
cyR�S����T:<���v$�#Ьډ'��qz}�U�K-tm��|j_����L�%�)�d22�Q�W^Rm�[o�Gb7n�`R|��2���η0d{-9�.���k�Y2N)!Ӑ:�Vګ!Hs�מ4�2�֢/���i^_0���iq&󐚋3����ׯ^p�Q����esE��l�H��"�����i�<�ëd��s�k+�q��|���l*��Q�'�a�a�Q�ߨa�\s�g;��{��)i���� fQ�$��xX�F �ۛ�o
��P��+� Q�$ Ir�ΜǢ�%^\�2z-V�#8��!lK�M�cV�7}t�FuR�Q���(?1�Qf���r�z��W�b����!��I ������>�ݽl�+���$)���������G�����ߏ���Ȕw��~�ÞK�9RF�&;�%\$�<�.�>�ߺS糫�\��D+Y�K���@P���rw��3���?������k�y��o{�y�ל�R�u+JZ��9pJ����4s�V��ҲhL�y
�9�D20A|���\B�沥M�o7���.�m{���߹~z>eN[��45�/��c���S=OA/'�v���Y�)	_e��n�,[L�\r��l+٬D������B��0x��i�x2�u�jj9�8 ��l�NO�\am@�h T�b9���|(�=��]�m^t��*r����������
W_��U^��3a���`���vY'�ݧkI�|�Y��r���H�3ɭ<K~�>v
��?s"�q���6�u���p;5:�ϸqk}1��Ni�J��lOcy�o��J�-�E��,���h۪q�fWȕ��"(��y�+�ֻ3���%o+E����������t�v�[y��5r��c��[-�Aov����^�Lu4����͌	.,����Mx�N�+����m��F��J�k�#$k��A�㙇�z&3h�^���:x���xA�'�wRc�dCg��S�df�.�-Q�98O�~_�P]
�D����n"�m4�p#�gX؜��7 ��4'�j�V� ���e��i��l �nN�4	8{c<`n�I��}��F�[�A��\��R�k�3+�r�H�qM@R��#Ģb�NHSԵ俶��i�&�J-�(V�
pM��uJ��R�j�H��f��0}�E%�w����g�~�����{�.��߹C7ۻ�ə��1:=�$�=y�����k���g�'g�bʐPذk�����2!�c���AA/E����� ��c���n��}�}��I�rQ�;����]�!�b��k�h�e�Ou�M����B+$쩖"a�!|��s���`+B��^�~B<l��w��q{��.��e ��Ҝ f��ۡ������t>_����jY{�V1, �?��V�q|���aT�<=�r>
?M҂��mB�5�hV$qWaS�G��w����M����'��N�Nj)��6��R�4�Z�Jp��P�$�খB3�u�U5a	��[��/^��0�Xk)?�U����L�g�G��fs�@d������A���w~���.�k�a�g���ʸ]��f�h)<�(��y��m�D�V�R����ϧ
��[l�Ǹ�����i��/h	����Zf�h�|��)=Un���2�/{���l��Y[��䇥&�Y�Y�u���W�竎�p��m*C-c��@��ϑ�<OAQ���z�^t���X�0Y�!��}���h�$*�A.A7@cJ�� '���[#⒎
��VA�U��TA���	�� ���-𴘻h!)XkK.�	m1-�&֕�p��(\W������Ňv����[3R*?-�J,�E�D�� �6�<�vBO��hs�� �!��cZ.6��ޠjvD����n��By�hwOj�
B��J��_�䝅�},!}����jΛG)c ���L�"�E`�h�5w'Z,L@�����jO���eY�;T-T°Q�;w�0P�{}@�t����32����z����?�g��c�ڑ\�>v�w��yx{l�k�8gV��O"U�&L���xv�]�����&����W	�9�1�Xlč΃r^Ys:t�2c�[��B�$[,n�R�t4�#ȴ��/���)��BiC�A�9������KM�B �p(7��-�\���g)��u�y  �����#�.��y���	��pɭ}ܔ���+ P�t'	�g|K꒕.�ڃ$���=Vr!�ҿ��1��r?߹ ��vPnC��!"�#p+Ò���5`^�{>c@0W��ݍ��Q�G'�+�+��������K �{�� ������_�K������<wˊ���+�%�I�(�%%�b�,���TE��<H'j�����1�ò˹#A���b���Uɚ+�������~�۲µO�{����M����牞��tQ���Z��k��������v��L���>\��G��J�{�x�ͧ�f���t78(k��\�I���a�	������ܯ���7c��i�����Ě��5Ozl��v��Avqp�3N�i�0�F�F�!I����(���:�BFBDU*u	,5�[k��P�]&-�	��+bHÂI�7�-H�8g^ 9@*8�ǣ pG� (璭Cml�dkO � n�Ah<t �F�� K7�
9���}�E���>���z6v}��	Q����Ʀ0 �S��#�4�ԾԆ(���n�����Ȗlq\=,?��#i�FXnn �����M�{�.����W�����A �a3<�9"z_f|����k�-aA7�R)o.9�6��cN�nN��x3�c}��xa�#;����ڑ4��p�-�k�N`\�*Y�u�65(Xӓ��%��
��2�(��X^H΀��Z� x�|+�p8Գ�/�_>����I��	J��A�o]b�ɭ�	_��l�ˉv)�	p�3�����0�R�����L���M��)k�s8�O�0	.b�7�V��<��Q�G�S����� x`Q��L����O���@aKGGgx/izq����ݢ'O^�� ���sI�}�k����)ͩܲ\x-�����N�<ɭ{�V��e��Àg�yyln7�VL^[��n� ��� ��Y�uEV�l1��$�פ~��ΥYۤ���%�cž�����98^����vQU���e�m����Ų������&����;�[{g��v]��/�y|K)p�#f	έ+���V�~�X.���'9�Ao�=�����]׹v��%�/���$�4r=ْ�һf���loc&�������\����=� D x�pW�XL8�`��c�׬a}��朵t��I��y
�wR޶��i�h �L ���f�B˭�-<cuX=#�n��},ѡP�[��[IB�Đ� mI�j�����r��JpQ�ҋ�8W\LB���ب��M��H��$.	l�K���
�!%e��ccÚ>Έ4v�m�{Ƹ�]��R�~aJ��"23���k_~y��x����+�J��"Y\��p t��}�+&}�чt��=�hŮ�08cY+��� f6��on�+�c|��[���g���O��Wl�������%��h��h�u���`��>�������E��|�v��fMH�BZm-K�6/I��8�F��p�:�����f"
�X�'_�a�/�ҏB�b������&��kJ�l4���_��{
�0+����K]{y�ݡ�R�R��$l��J�7�����G��R�C�w������P��?��+f6��n޼ş���l0����\v�Y R�Qb�Ú0E8��u}�<�($s���l���)?����J���'�ӟ~ �M���\���+�lA� �)_'9uT��<N9�\u�@������ݐ����op�"f��n������y�ˏ��W*NSkI�&��d�pm$����x-�-����jR�G���T�y�m?s���g�X��C�w�y�췠�c�+�IY��qzȞ����r���k���LR��fq���k��u���s�n�ۖc����)vw@�si2���3fƚx�ZwqT&�WL�+���u�K�Q�<�f�N�%� ɬ��%�k,��AYxe��~D�������*�г���B4!�7v*p �R�$r���
����@x�GL[X\䣵O���H	qb�m[
m�|5��6��gC�Z���i��$�  �.h�|�%�-E��&��������6�
JҤ�b�e��g,��1�D��]6i�B��F3R��9s2���Բ���!k�W�e^��efc~�l�r�����g��_��I ��! �dh#�V��d�D����6`�gB�78x>|�6��tiN�o�2�D�c�']k�q�e|s�g���}�Z/�b��(0����.;=�E n2�K���؆��P�J�:����c(v�.�H����"a��_���}gw�67J�`6�-�Ֆ\�]fF�l��jcrӖ����:���2���͙��k�Q>wEF���g���[�j�
��ֵľ����?aEQ�՞������9�����������B��X�&��SO��Ck�?���4XssM���h"g�o�i|�8��<�����?���[tcw���{����$��+�9�ǅ�ڀi�r�����G7�`]B�Yjs+o�ѽ~ގ�Bf�{1ȕ6;�rs�����+�k���/%�)�9̙<�rU����)��s�&�eEm�9�L$�
#@2��p1(�ܥXbNLG�� s�B�t�5 �	��ȧ��'�)ܳ�}������m�S経����u{ћӾ��Gt���;�S\�Z��hL$3�e}��ꏳ�ͼŦ|XX�ȥ�Jk�n��b�b�D�Yi|��Ќ����L`�owGl��\�@BX^� `�dkI/����͈�� F}��Մ|h�CE4P_�E(`��E����,j���wS4�����` 4b|a`k�[S�ѫ%x>�V&�.olF��f�z!�;$.Ԓ�Dl���9�(J����[Gj�b�q*	��l�Th���v ����f$�q�_n�X���Yo��^@/IyD$�E��5�{��3���uI�i�U�DQ�K�a�Bc\(g1��p)��+=�kZ��0 �/�oQ�t�q}����o��~��_�/~�vG2��@��)c��U�Ւr1�$E��3��ĨP���n��1p��X�-��1�l4�G�e``٪:Yl��vYlh�~艽��c<>uks��&�r2��SV�+e�;Qؼ�%\��Ǔ6��Z�uB���������D�D<���]0����I{�c��?��Ȕ��$�0�8+X�u��
�oA[[;��+Z�[P�M���%��~)��O�U'�ٜ��R
9Y��-%;.�{��{���NpU��嗿bk�|�LPq�7��D [W^�%�,�'����m��v0^H��g�)�qȰ��	ڌd���S^����8��ŋW��_�2Ȉ���[��[�}�`�`Cr�,p:�LW	���u��nHP��?��Ϭ�+�s�ǯ}�����e�	�t?6<4��9��\O� ��	�`j���Mڿ�M;7&B�Id�D�^γ V�8Y^��CK���*	�K���[˱�UPt�� ����\�73�~~x_
K��J����Bc}�NO(��.d��vWv��}Y���6D�}�c������!{Yё�E�{��{��g���[_Y�g9_z��]�:��$&��+5bz���Z3�ZSi�w�Xyy�$:����-�l���#�d���\l  ꡕW�y���
y~V�d\����+����*Pd@�d��B� ���x�WZ�5����xS��O(�lmQ7!2E9�#�d�0�1QϠ�hfɫ�2�;���ˢfk.�&x�vOq���I��^p����f�)-�� � KM�[K�#����]�教��"���r��h
Q1+�{4+= �2<�RK�����l�t�KsK�_�,�ج��{�>������;��O~�`�qի/8��C��ŵ!�Il#�hɆ���������$�q73˴���kaF�>Jz���}�OO�ޓD(pX��c{f�W�˼��D�ͬ�ꞙ5��D�5]&+�5'�=q����/,fQr�Y%&�G�r!#;v�"���M�\\�ă�fa �زa��r�_~��(��h`��[����$�1�VÈ��S��fu�.��w��wn�J��.#�}��R��cU�	)�]߻����rkoSn\��?�>���Q=����G�7� �B-��C&Um����z��\	m+��oU_��?Ɯ8��R]�v���[I �����<O��?�T A��@.xQF�(������#_�Z\�Xԏ/�;�"g�}����ؖ����G��?���y,x`y�,�rs�&��_<!����b��	��둽���Yno�~�k�߻L´�o�.�cy��_�W1���'AF��\x���@�h��+�V�U ��������}y�{$�\	����K�ssX���3����ơ��)WB���L����[�npu�$;h#��K�i��(J��s�p�=�|=`��лt�8��6 }��w�Ņ��`���J��)H�o�.�X��%��?Ѩo=0R�S#�s��^T�p�͜sͯm
8�n��/-��B��F_�Ssi��gM`*Ղ���D��3@�G��b �s��jMb�g���_㠶��Y���D�? Q�j�����T.�P�଀ ���M0�Z�3%M�� ��	|{�Į��l�+����!�u������R����L�D[��l�,2�|:f� ���H�a,����h�R��]��ɓb'��,�;�͕�D��9���p9�ua�kyۇgOづ'���1�Z^�PX���'�Ow�+h#��ܼ�'����/~�r���rک|�9��}��KZ���M�^��J,+lL&OX�=|�(}��?�1�T�Y5�tK
/o1�$j�从�y�zu��@��j���^����j���o[l��{(MӂY�]�<��l��j(�久��H��7�m�d�b\��Z56)��O�S�wgG��
y��%��t?`G�su�R�:]k����Y ]_K��Ef�����ΰ]�-/�c�<!���*�@��ꫯ,02OR?y!�������Z�����/(�:����
#0Z)�_�nűeׂKTZQ�d{{W�޹'?������2"跛>��o��J�5�|�ɓgi�R>|l�f��s��2�n�� ~����~�x��^���e������f\鼱�ue� :����۬0��;w�W���$���E���]4E�r���6�̳��)Z��Ǔ	}�i�":��J+L�`Dl)ў�:�v�v�,6b�|�S�O�"�Q��6�̤_���1����<F��z�׾Us�b�ݘ�0s�����o�ח�n���	Vi�le�� i*��j�64��yN��L\��@"�y����Ԟ�"?)'�.��gB��4�#�R�эx���6bٝ�F �"k���8W�b����1-KBk;X�$�PB���p���h=W�Z2�Щ�����蒳/��+\zP��K����#_��.��{���z��,�$����<z	x�@�4�t��<�&�Q.�grzx '�G2:9c���T�8��E�IG���k	���ZE��?M����N�x�27F�U��zۻ߶I�!�9����s�Y�uŋ��fY�j1M�si��Ɓnk����Jt[�a��v����dvY�*}�믿�?���?���g�}.��:�������:7x����&d`��\�՚�sVM*Wv��d��nuzEhe�9��G��K�߫���1��r�v��ўO��A��*8?Xc�D���h����`��/��)|��U�ݫ�w���~̇��D$Enmm˵k�����ԅ�x���.	�y�����YM	АAچ\K����\�S@�TjNB�";{�1w�k�$��~`�v�?��v��M��;���>{�z��N?������m�x�����?�.��^�vro�$�'ݽ�=�v��d!���?��ܽ{W6�¾n߾��dg�!�x��	K��8��ec����	ۮ�.�EV�Og�� ~�>^���x�����+H&�c�`�9���@��?��蠿���WT���om+XkB��*��sU��\?3��z�+�L���!����<�� ^麒��)H�����y�m�ռ��ͮk��˶�m�N*؋�]����I��!m�|������W�Å�Xy����m�o?�u�Sy�XqG�������!��n7�Ʃ���)[�r�?�ql*�����ۙL/�6��M�%@.�G����w�zvȕ�@�ġ�P�\yi�'@2;?���I:�յ�]���[���R���e�2��F�:�l�̪�L�[Zv),ǰ܁%�y.��D��x���P��
����T�`Q���=f����leB�2/Z��`s��V~�ab�xt*G/���1nQ�5�/]��x��m��n����6m�,ioV��o4*��v2@��-s�5�,W��ttgq�P��,��Q�chiYu�d:��/l���f�Bn0L��������Ԕ%�������|����H�/���y���Ľ^i���S��ںL��O%k�&-�ʪe�,I�����'*�W�RL]���M�!0/m�/i�g���.�?\�  r�lH�+�m�!�ţ��o����6(�$��~�XE(+�h��A���h޷^O��э�0=I ���>-�����[�5tݪg��k��x��n�dR(��q<;�;dTQ��^��M���'[��%����e�����'r366��aem��C"Ɍ��-�w��_X����3�ܹM�;kA!0�g)�m�S	�P��w�:u���ؖ��U��>��}^zc�OWK�&��*,T"�V|��Aq
�Ҥ4�� �ej׻��4Wk_�ݦ�9�d��3��`IP0<�%�Q�e����vw��d7��
O�Wk!a,�;[Aokg�=1=���Z��Ch�Tת����������ɸ�K�.>�ƌ/����uв_�x�/v���m�/���wy�3���C��~Nrn�p��:��M�G����Φ���I5(d3ݛ��^
p��<���������W����>�[�g���ѭ EzE��G�F1g1�������r�‶# a�[[���}CY�F�Y��d�z�\N'f�X���qn�}ړ A�1�2<׆`�4�� ְK�
��q���:`�n
s�e�f)��e��| c&[ii��لeDl��t2���~��c���op� �Th���1���m��ť��eS��-v���f�{Rh�-�cx;��gH���t�P$.��A���ח��9��xR��x�����Nl ��9����,���������4�������y��,�8hRڑfo�0��0��|�zlf��m�";�T-�����iȿ�m��2�}�ݟP0�mc1���C2�2f�T�+6��=���������7go�)��K��Mmu��K^���yy��JM��sժ,�L���h�'�`Y)S�3��nȝ�w�Aʀ�`�oܸ�@�-������G��/���?�LA}�؞�:�U��v����,ک��c���J�}H�~����t�������6��n�f_��wC^�|��%-��L��!�UޣﺐJ���U��o�����^��!h�
��J!��+F�`�w=�{�n��E�7d9����/@�gm@ڤ8��}���\�F�躶�Y�C��5��&�>��Q�KƮ�R�SQ}�����وd������х`���5�o���7�,.����Ûd�8��A��n���:}����6�	�@Bu ���\���[�(-+�y������"���ַ�]�*G%���ձF������l��v^B���u"���f'��V��t*�/��p�X���IY&Ğ@�lg�K&�;�J�Ij�*}���+�� Ԇ[Bhҷ�D�s���P$�%P�v.c$��щ{,��o�N,�F�E�R���Z�3����`,��Y�=���}�6 s��.qn1_JtBxyK������@����11�������R�\�\��t��N�N$��G����L�������f���BN@�Ĳf�z���WRS��+��y;��M4�Fok��Afٌ����F1R��3�M5^*�:b�Q(�n�6qK.ݺ����4��cH����0µyH��� ������i�.��lH��=�} |g��ö3g�oO�0t�l���e���A4g�¤޶��ӷ7I�n~-�Z5���J;<0I�����Z�J�c^��h�W=0Mf)�M����Xˤ�4��ͅ 7b��㥷}i�E�޴	�B����<�Sٻ�Ǖ����we��/�hTn$�
��x<K��35ã5���'d�}\O�����]_c�V�ƴ��r������j�{ݾ�α|�ˌ�*p����E�����Lb�\� H�H�O ��ȥ�ga9'N�Dνv���?d�� Z������jW�u�ҡՕi^��K� ���|llW(/�q��v��C��|�=Wh紸�^�.�phG֥{��|x~/l��ʊ}��6Ƿ�[}4W���/{����L�shx�|� �L�[M��G�
����o���V�f@Q�>C�����2��.���~V ��
%6���	�B��r�<q%o�:�S8#���C~��39;H����~?u����y_z.�	�)h�V(�u����P�\G,�0i���`	�̡�]��*�Zb`�Y��r[�\��!r�Jni�e�Ƭ���a�3�]�߬W��'��;P�Ll�;�� �z��!�_XbxЇLc'=�L�,�~:@0r���o�]��{�u�;�_��O1/�.�̌F���T�[�P�g"�,D �=0�%�W�5�P	�}�:�֣/�)pg�Q�b�s�w57�%d0S�A��K%�B,��ji�����bX����Ɨ�<���`i�%������T��M�����eڜ��6��C�@Չx/vEc�2��6���]�|��c����R�'��m�^���JVM�,6�,b������+����W/�����
�nA�VI�ѩl�6	�	�]�����rn�u�m��	ՎON�����#K�kw_q�ݲP]�[0���7�����s����_�F^�xA)������r8GZZ�?�k��e���G��y�����Q�t����q���tm����ݕ_����Nr���-�M`�Q}�0}��|�r�q��+�f�8o
�W1��Ƕ�;W�ס�_�t������%��_���!����3(�ˤ��,�d�<I��h90hS�
�Z���YZk�b^p�ǲt�w=w��\��4�=�k�IO��)�]j��e���)_�j��s��i����A�%7&���!���ׂ-EW/�P��p�.�y��ϋ�b��<]Ht\��A��%
��.��	�lls_����ߡ
�x&i.j� �%���A_�_y��7�V^��'��ah�WoD��M�X�G?����i�ؐk��r~4��4��sս�([�uݵBYA��D0k��h�:�hec�ˁ
~��/�0**��V���xH�'`9J-�dz�S9���0"d�c)�f��B[���-Ҡ3�%0:��r�������M9N ������
Y����ަl\�.��o���3�{=�r�� �
B<��8vl�.��C裸�G��E�~�c7:�\j&��Ђ̖2_s�/1؊A��1/f�ǖ��Q�4���t��͸�qL�1,�䢱���{�����	�i_�@e���Ѷ��D-N1��=:�������|�򒛞�%<������}Kg����Y�c��.��u��eի��:����^�V�ʚas�P����,����~ݘ�$�H7��w$%�VS^;��-&�]���_z�D²��}`�r>��M�/���LA�Vi�^g`�۰��{yv�򩇼��%�Z�+e+���`l� h��1�љ�|y����O{?�8A:���2�g��g����m�E &��y���za?���$!*�1�"@�5C���/_ȃ_�w��
�l2=O��M w��!X�{��b����'�r_Ϟ=��m���R��c�l�
�Vݍ��u��w�Q^����-A�X�������E�cw����0�������8�B���&�ն�V["xc^�:wiP�-��|��#�o. v~$�*_���n����L����;m��ӷ����B�;��}��|{��ge/��A8�uu��$�Z&(�9%Wʃ�s:[����/���P��W��2<zm�]7:0��	ao����.�����B�2 %=��'�CL�rz���}�4O'��l�%�����>�v����� �S2��,��8O�a�x-� ��X�2���V��`�L@T�E:'c8�����i���<儇�N�̙m0���MU�9層0P�~��pC��{O����ؕ��3i��:�A�҄Y�Mz	����o����nfo��$��`Ѥ���t���=$6Z�;*�;n�R�'�Fo0Y�`��"|T����9`�U~a��uBfu�����3�U�d�7�Q����}v���i�A��wަ��4Mθ���dK����3���cN�`��P�c�	x}C; x���9�nb#�w-^�@@�,�.=���}�̹9`��x���]6�,V�V`�Kg�m����\Y��2� !�� Zt� �	x�}`gg[�ӳ�>'���D�z�������a�A],�����u<9�dg���w6Y�_�_�J������q������W�;Ɂ\g�.�
]�������A�qW!'�����?������Ȍ��7�`	��a�<~"O�<�><�<!ql�����.�|Y A�ȡ斸�S������y�K�0�& <���Oo�Cz�����@��v�=����w�-pV����=����e�>S��2�?�Zю�ك^�ok/3�԰�]����67��g2y�Z=�ƈ+���2iex-���o��g�8$���+�A�%�}���V�م&f�N:}����M��Ë�v�Z����#��l����2��j&�����ǔ�"qҙ��6[��E��U{p��7��Z疬�:�"�2�kr0��z����/��ۖ��z:�4�^K ��M�u�Z��o���߱2�1��mٽu_n�}[��;	�<77}'����I� �鵁��SQM���Ǹ��i]=�‿c��|	F����$�
M��],���lzB&f�
x�V��	�I���\c��b8�Y-k��[���nz�/�q��\+ñ2@���J����C?��^��r?�XWܛ�˷]<�c��b�,aM�,o����� F3�^�n=�.lnm0�p��h�������t��mCh��$���+�	�B[�����ܭ۷h�������*���ߒ��6mq��B��b���P=z$�~�)�P=�5��-Ϭ�0����%�u���l15���Fc�T" ��bFOimv�ס�kY�Ev�ٍh���i�Qs`��^f'�Z����ľ���NZa��c�t���`v����g?�����<�J��bN6����z���1�7`�2�Q�l=��;Y���op�Qƽ�y�}�Ҭ�c��O
������y�^Ay�%�-B��h{���j�U^ ���a��ː
�_��_��AR��l_>����^�7���jˌN�ltHf	E��ݫ���͚E��ի
]�)�)T���^:0১� �Y���=��203��������������I�jk�˹R��}���Ӊ��&8�P�/�ZsE育L�E��>3h��t��1�
jN�ߌ�2���⶜f?�]�1���K����t0���q�G��{�vƦ�;;i�������UI�n���Aꌵ�K;]���1������$����7ݴ���Itzv��c��1��>Mxb-�GA�#4�y�+�����:��+�ǁP�>�^q���F/q���R�؜��	���k2L����ڹ\��-7������g�c����벶sS��Z:qԓB�S�7���q��[��ժ�Y�3~.�GY�]]/�����;z�6N<�2�TjN���L�ߦ�{��#���g���e9h�&#+�
mŤ�a:�^1$#-,o8��z�P���.];q@ԣ���Fw��5'��#��T��HR�faMI�Y�Uw��F
Z����;m��[�б3Q�e �U������8� �Ē�g��TvFO�Ȳ����=,J���!}w�зw�����aa���}�˞���$ek���"(� �|dx��D��6Y7�K��ؖ'G �H��ḁ��޶c���`��5xD�O��@��ʍ�TO�;:�"/ɭ<~�@٘;�S�� ��Z�Am�2�j�3�W6�����NNNy7�7��=S���Ȫ夿%9C�=���^�+�'��]j�e�8� k8��:�ݶ�'w�=��$=\M��[�q�t5��n��]O�i�@.�Zl�:R��x�;FxH�%^q��o�_h_���Wg0�2�_=�R���K�]�H�>���uK�
Xr�c	��3��t�����$�o���ɥM��<{�$�����'���/�ŋ�/^�|PUe.������^�����p[J�Za,����B*b�+�U�l��N��I^��:�,M:�VJ���\� `Hw������0/�1,�Tݖn�����Z�?Za���c��
����"����1�V2s�X[��{��u���*��߹���u�ά�(�?fP��!p��ϧ�|�%��m�;��1(�|�BM-���o�-v�p���2k�q C�;�%0�-�=aBd[�r��-J�z�@d�sd���vBf��LG2���K��I�Yғ:�l�8=F괐�k]����C�5�H:�n�Ѥ^7��~�1�+����4݀cNt��	'�ؚ��'�%$�d���졌1F��0�Y���j�J�n�Q��LS���q� 'ɴO3��&¯�zȊ�4&`��`v��"˺��x�xO�o��-����ZUM��5�!MI@���A|`���xc`����2�`џ�?�J��{���2��(պlЗ�6�-���B;��c.C��'�, _�Xg��۪%�VҠI�8.��߹s��NX6F�9���B�w�&�1}m�,�jԨ���[�罪��Q�djZ���[8�Iq���"�`��?�@�_|%|M?ST�������W��^�p}=2p����4�{wؽ�6���T`�W�����נ�d,�z1#���9��"�Li����49�i�Vi`隣+7��䭷ޖ�9X�)��-���8�-�Ӫx̐7Oh�t곿"(G[�L{���?oooH��FP���c��o�Q>����4�JT������ޮ�{h�^��-��|.�'؜^O�2��kez��7+=%Ӭ8)r�CP��{�A0$��J���(��rm}e��]�^�Un��~��}�DFh_#�ſ4�(pK;�w����
x9�6�T�zX�p�������enU8�9v|�r���U����[���y��t�Y�=��7nv��z�Y���Rǻ������HZ����M��j�M�␱���H�ŭDѩ����nr� �/Ȫ���nr���ZUmµR�'��\E�0|�Inu���,J��;A/jc皸v��%��r�_&���xҌdk�Aq�I�� V�a��^���d$��P��Q'��Z� ����I=9��dC�����`������~צ��%��i漣Y�]����i��&�o��Q�#3柵`�L\C�bتA��82�Qf1$�K�(j�0��Җ�E�O��Q�iR{�2���8���4�ܩ�T��+v���c5������}kϲ������8jb��}(�M簦60 ���z ci����#e�?4J'j�H%�f����&&��ߖ���C'���������>��o�՜�V8�.�R< &$2(G�R�H� ��ǣ[t�C^ j�\Z£�V�6V�
��9����,���	���ecZ,93���)d7��K3�/K�twV��R)E ;�P�:@�F��;ﾛ�ӌK�(��T�2��/~.?��	���}n�~d��9l9�%���ͶU@�B�{��o�+����X�C�6X��t�*XcP��(7ҽ��5Uc|妪�%	�Z2H�{���>�����1�2k4���y� �Z�BV����DX���י�DSH�Fg�rr<��g��2������?��c9:>������B;��c{F;��
^C�m��m�@w{�b>B1/ܲl�l�[)�ܕ�ׯS��Tg|��>"���3J�����Zc$��m��!�rݬ)Kc�qm�<�k�7\�4뛗^mQ���b����Q5�N��-:c�h,�K�q�Z��sҌR-���h2CW��#Si�Պl��3���^�0��(
g�y������UW����|��/��;��ɍo�+���X��˅���ïy��ZZ��}I�!��0�����@�ko2��,;�ZM�o�|���*-(	�@F
"+� #7���ֶ8��*�� n)kU���W��<H���]6C;U��q���|���dZ��t&<�������Z��`6�Ez�Y�u���tJ3iBM?�`y6?I��\B�I3:N��d�ZU �NU�0���d��ji��Y�p�߈f��-.уg��vc,�;�e7�l��D��l�.��a7Tje5�ƪ��V�悪�(n1�G�t��6���P������s)g�� 3g�8���`���/��+�w�����]q�[���J_�x_�P�7KpJ����l�$ f�f�B�3���jI��'�tړ3��A-N�~ ��̐��l&�`'>|�R�Ϟ=����/���/d{k��s��͙b&x�^a�,�g�~&~�a����OQ�~��6�޳����'��ƪ�.7P_\�v��6�ņ�v}}����,:�sA�*�;N@�r^�(�I6	Ih'gؚ�,��2���M��ݪW$��&��ܒ{	�#I	u�?��C[ ���}�����|��h�Y��q���r(܎#+'.K��l�0qK��.^�O\��et"H����xD�w��P���V�~��@�ƀ�8�>�_0n�G��4��`x8SYL
H6S[��A���8�dʲc�) (<+3�`�������޽%�o\��g��{� eɕ���}�C�����O�>�=��y/�v,B����)�����y�R$�N�2�0f9a6����w��>���wR_�{��x�HX�E�e�7|��G
�$��9&Z��<�B��j�*�}ȃẾ���u���>��خ�%ƥI?�h2��w�:
5��� ��@��gn
����Co��u���2�j�_)�m�TI,.gssC*2�)��25M�Pf;x���<We��p�ZF5.������hg�LD-'��9�I�.�Z�cѓ��7����[���<\,oQ:R�WX�������ᵭ���2d��
tI6�zݭ��_�����1M���jr-p��f��"#�f�K����x��X����~��k���Y���(�g�/0-'���΃c���C_������u1�DZ��鑻��M�R0���m��{p;j�/
��s�?�o�d��04������sj�U�NUI�hް5Ya��õ�z�a9��=o���=\�N�b7}��;��o������dV����ޏ��$�;�+�����T�,��A�e[�2�9h)��3{Xm�,�b���������/�1�%�9��(Kc����lt�� ����S��՗_R_�N�#;�.(0q��0��~�O��j�U�Z��$ޣ����r�k1�b�G&9��(��D:��&p��;�����3�_~Υ���M-�gL���n��<�8��A�N�x@t^�r%�`E�����hl�<�@nܸn�9U?y��m�}����?���]]��~�s`@� ^����t�l�!�l�l�0�9���9Ў'h�U��ݾA�,����5,.�U�eܘ���q
ƞ����3V�>�'?�I��t%��&��z1^춝-�7���"������l���[��08˫;�eMT��U����J0��;�b�u���9a��2/A�A�^��vאn ���� ������_�R���(w@;����ibf.+�W��|� wN���j�����Kh����?D��koс���:�Fpi躁��^�� pQ9e�u^o�4�
���E!��%]"�' Ƙ���rN�6���;X��A��}���t��3��K��tE��8�]f</_�`�B�cYdr}�y����/�Vg:��V�pt�[� y����5+�h.|]�W��+���??oTKl%}�LI�u�ۻIi\�0~�j��GvzvB'���S��2� �AH#��]�|J�&�K"Zp{�bXW]��0��2��d<=�^���ҧ�.��Id�� " R�^\j�zp4XO 8����4��b���S-'�E5��Z3"@T1���1yD+�[��ݔ&uLH!$�|�yx��@����jecLl����[ۛ
z�z�֢��X<����8$0�q���-��������< /҄�"���w=�C�H��caE�~�x���5��c�]��m�� � /�æ��4S���)+.����2,�ˎ?2-F���Dk��� m��jL���R�A��K���eP�v�_�ΥzL�7o�$����b���p����%�����4إa�K���=q�l�-�!�Q���ǜxߺ�-p�ΖA���Z�Y��6�C��q�L�d��ܖk��r��	�a���g/�l� �FdnݺIM$���0|��bի��)g��4J^�?8``�Ο	�)�b�����8L�����O��h�r.%W��g�2��VL���'I �;�[yU�nT2'ڽt.^�Rp͊����w�Ռ����;�[���o3C����J���k1�q�!�'��4�A
��|��>����%��f���	0�-E]!
қ�䭷ߒ_��o��������~�	����}5Yƃ�U9Ϝ�0��� Fgcy�l_^��r297猶� ~�;^�e�zk�R�Ƥ#|�v3I�����1]j ;���u�2�i��"��n�ĶF%��`x5���鵦� ,>�Lj�#Q���K�.���������=Ho�V;��4��b_���u�W[��l�%c�U���$�w��,�\���h��9f��KA���⻱�֪�d\w�􌍎x�1E���R�|��k��:�-�1���ЮR���<�L����F�7W�d�A��՛�z.8xpc�\��b�!&\��Q��.
�޹��� "�dOu�-u���i �(��Kln���-�� ]�ݲ�����\-�^����3&��R�s`�g,Q�"�V?���\Q[��R��^?�����k�nΆlnn���Ťdq,Ee����V��I�G�:�u n����П��}�"�G	l<���L&(�A��hY�����1Zh;�/���؅�7u�����?�֡�jzMgw֠1�Xr��S���$gu��:^��:(8��+楷�;����p�A;��S��������O>��ݗ_~!�^[rЊ��&G�mb���g�N1t����������\�U�I�������b��_|5���t��ݹ%��M��)�4�b+��k�hB�_V���+�����[ 1(&�}�M�������_�2�N�o?6w�� �{ſ�}�]�s{�A������zWd���R0�2]O�m�+(Ѓ
�������5�l����	V��AyK��X�ܬ:����)�uȶ��>� �''�����oߑ�߹��(L$Z�*�jG���<�y�� ���O�S�8��#4w`[�D��5�bn�Z�en^�8����!�S�$���m.k޺y�רf~������걊��~����熹~�ZD�ǜ6���v�/CY����]>?ڗݝ-ٻ��p��x"�>5���u�~� x����K{_�zXd�Xږ�F$Uf��%���e�}ܛ#D�R�`v�4��H\���d�3sȫ�ˠס�%�fN����Ƌ�n�]��ʨ^�d=����L�,�}�#��+��XL����Ҋ� ��o�W�ۜ/��DK~�W��_�6�Hp��<��cy���4N����k���2��~B{�;ތdR�������[s0�W��x���d���f2�Ne��M��nj̛dD	|�7a3,�fvQ��}���j��F��.�5�f̒R' 8-{����8G,)�"|�E�n���k>8���,� u�����qa�/��r�	,E9���ڶ,�w�`�(ڨ��M�������)����r<z)�f�K%�g�W�
�h_��f]���%�J�-�@�8�@Ts��g�{a�a"�U�@�T+6e͕i�}��n�e�+�1B#&ʦ��lcM[�����ŵ�]��?����y����K��,��~���%]��% L���<�2�6��r�H��	��6���ZU�\���?6�`v����?��ڦy�9�C���4��E5�U�],�C�׬�����O�q���ǂc pG�>��h��T�n���<�)Y�����S�������}��� ���u�ٹA���񾠟c)^e�[���,#]�?4�d�7<�n�T����&�����������s�*���a|A�	�
 ��9�"23����e��lV��+�'�`<��s|F���,���ʆ�^����?7�<���:��H�|���BX�A�v�ρi��Vi� �J��d$:ChPvjr�U�kY����U�"�xq�/H �����d��v�w�8����+}��ـ6��3&��J_�1��#�+�>�DKʦ�zi��-e�u��Oyj{(E\)p�W�C,���W3�d1�����>E��t��3g�䙱Bp�g�*�嗖ޗl
����^\��>�l|�Q�|��%s4�L���|3a��z��VF�ٙ��x��*�.(})�*�k_��W�q��p����?�g��}!�A-�GG/�E⭮�gw��3�V����Zĸ0�� e��)�w�o�%F�S���]؝�H΋#�Oe}m*õZC���ғ�«5��1�I?��>?뽛���=�7ؐ,�Go���r5���F���b�G{��F���]h��]�	h�̈́剫�v3��J����WOb�%eR�����giP?L7w_�=}.��ci�.�`���',��mDuy෢q^��`���y���H���ј�ମ "yP������b�l,�tN���.��b���4
��h���NN��|�6lm���t5&JO��/I)d�V�L��[R�c����5f�xqN
�����a��3;1H.\.�6^xa����e��(M 릕=<<�w����\�Թ��]@F�}V�x����V͍C�UY�� �����u��#�^>���P� �O��ev��_�=i]��R���f�@�)�+3�_s�EW������@������;�R��՗iWx����^�׃+ ��Pw���S$n�d'gQ�N��j�&�����~uf�V�i��h��P�r>:�޾���>��` ɢ
8�<V��Ǆ6�Y�L*=����-�V<�W\a�l昵�3c`����R%sfy����!]Sx����?����}K3P#9��!5=��IN��M�	�+L���*����WzYl;�ۿMf� at�H�b>89>��'�_�8�7vdcm��"����1������1����y��6_q��'=tR{��m�Қ��vv�odol���0���}�.�����v����l�(J����e{�T3:�������Kg]��W���Lȣߧ�L�ۭ�lX��gM�q�4�Xe�p>��|�~��cmJ��f�Z��ǄP���a���:	x6��U
;=~(�����׿��|��OR�m��?��(RC������o�?v���1�^�.���/r����|w$䁴=T{�߿%5(`�d�8h3�jʹ�*���Iy;�3��2��'b��A!����5���3cӴ��ɠ�{���r�aY�:�1��r��4}b��v�,��W!~����YO(�Gb� kt
�^:�J���TQ~e��>���I,5Sk=J����ɑ��I�z�󨍈^�k��Ҁ��t:��>����B��Wm�/�_b[�16����`F�f�B-[,i ��������'�W(ڊV �h=ڄ4H@�I���i#�������V�����̢��{1�bóg�V�ҙ���E�uH0��8��p�:%
�-�[T]>�+����E��/*�ۂ�H���h=�����K �k� �=��>�l$������Nf��gF�|�qt|��mV�«T1�����L�Wm~��Xr��u��
\t��U������X�� wc}K�?3����)�8��*��uf/^�1M��r=�<y=�A�f�c����¶��5����(k�.6gms�!w��t�aa����ʃ)P�#��4~!��?~οU0S���Dm�ll�(����b/`|��N�EO��@��Z|��|�)Qhz��u�C�-�F)��R&6\���_�ǟ|L/Wr���ӵ���w� ƺY���r1׾T�:���l+o������|Y�Cd�מkp�08�h��9m�����J��zZ$��3[U$�0��h��u�o������g!ّcg{S����دɍ�Mٻy-��8V&�����"���V=�X���m�2	��M�2�`ר�������,��j�?�Ly�/,hn�r��}^n�R\�ݢK����봿��a���[�xj�!���/��C�A�%V��iTb��y?ѫ�	��������ǟ˃���80\�*~M8�� xg�s����.[!����mIk���f����}�����^��.8��)��77f(2�JjcL�R���+��1AoDD f�kPb�0�Ҩe�V�(3��6��q�(DV��EW�B�ټux��W�+���ʓ��V����E� �|�Ih^�J���Aa=,�X�6�b�|5�[�����-!]�p"�vxO'gr�Čt}  �j��G ����d��.��h�D�K#��fi8^�շ|��{6P5u�&}�cg�$����^��mg`빼oet��fɛ'd)��,5�q���"[,)^S�ve�ɴoJ;�/���G�{��-p�1� �]�^&���L�3���� �AU?{b@��SЫҴ��9 `&҈����>n4`q �˵-K��}�d0\��T�܊(���C������f�d�%v19�Ĥװ�ҳ���o7�/�?�}S���<i�`@6#]��E	����S�=���'�{7���㧬���dl��;�	38]������!�,�?�`S��ە���q��Bp���.cR�^������8[���)�y��~���N�~���x6ѕ�Mn�Ԩԡ��	ɘ7n �zM�O�Q�	��$J��A�,~�MS+S�D����~x�EP�������6��?*��/-�����VK~Cfr�ō��g+tޗ���vy��b��_��N�SS&���H;JZ�U�V,N���i^1���Y�:�r�^�|i:�!��|�q��a��o1�\"�\K`wKn��$໓^���Y�be:�2��w �8@,��<h���~��lp�Ĉ���mZ�[:�m���_������� d���պ�	,��f���l�i�bcN�\.�Rmb�hRtӒWE�%A�p^�U�mf��ז�r�Q�;7���W������{�z�a�1�=O�x��P��il��i�ߝ�w�&�+.N�k�y���3d��A�	=g�Tu ��=Y�D�J�kq�u�Q�-��SËfV��mp�?�0`q�	iS��N��i�N�1S������31�Ȝ���R[Pw�#N��L-� ���ɸ!��;�Q����:��!� �l�D=�	��8�Ճe��76we;M�������Z��kq(�g�2��d�$�����E"\�#�or#v �,��εw �/-]�E�t�n��u��w}�e�vD�_g��m^k����Zo���"����y�[浤�|C�RÇe���ݽG�XN ����=zm͋6hr��]~�vz���]xnv��t�ʬ��&�`ZXT�d�Z�X��JHD�X6����c�bp��s�����UA�^���l}��'�'oA���3`_�33�>C�e"UA��0�R�{�o�e�7OF�|�6`���.����,mQ�ac�#`�}��R��Ԟ���;2�gg'�7�ŗ���V�;�ԥ#�o�f^���e�v�����*.��7�w�m���������0t>��}��ɜ�#�_�P�*L�47��:��=�g`K1�c�����)5�h���n���6��HH���LĐ���'?�Ãcf���i7V �����d\b��A(*�Q�-)�~�����\����t||N�&@`�SQZ�2QUy��Չܺu�l4��`���XHX� �5~�I\���6%�l9��:/p�A�vH]u�M=scN��'퓋�� ��&:]�N��:K��фK�z����	@ʓ��esrCa�a���đ��d��ň��u]F�\���D��b�t���>�:��oc��ɩ�$x�h�W�cw��K���;D{d�����kFR5-�춘�Ԋ}
�9�W�9$�2���m5ʮq�����\�>��|!o��N�\_��]��b$ޞ��1j=��MWu��{���d��[���s���f� �.�
`�S���ϲ<0"�tC��;��K���`<�"��{��̧k,�[����D
�X�&t�ˍxV����Fo�j��v�dQ�an��'.��(��Pq)Q�|������Xem:֨����D��C99|!��	��N��e��l��g��ª�]O n��-����k	�6e�d\�}LNd�"�w�Ze0(��j��i���|�|� z�۫��Z��"z%5�2~Ye����Ғ(���Af�KKk��(9rT�W�nuc�5���+���/4TXK{�I[<��;�v���(^�v�� S{AU���ȓ�-�J]Pҙ �WQ&Vm׮�D�_��U���~����9JwI&z�ѯrf�:��m��,�1V9	���~��* 
>@YS���+Z�Ulګ��7�.�O�X���w�{��}����Z[<�����}&IQ'��n2��KG�/�?������.9��A���>[s��ĵ���,�c1fǗ65��%�H�����U�
NL���v��[,��sK��E2#��ʮ�o�Vf����/��s�=��G�^>zzh�AV:�M� �s�/s��%Z���\\r��=gH��hs��^����	k߅&���yȡz� �(Q)��^����D����f�~x�w4JP�e֗L2wr94QZ�>?5�"���i��Q�
�A��fi9A�kw-(s�(Xr&�By!�F�D�=o����NU��P�i.d@ͿQɘ�hyxuo)3��(�W̹�o+�����[��_�n�q��K$@��2��Vǝ�3g{Ё߅�zs�����#P[�䪭�����H	�d��o���\�~���m]�@l��� 93 ���i�X��rzo��z�˘�o�u���r�F���	\0���@�!5�z$2n,��$��!giP������TFG2�L�����nQ �fh��iL�E�*z��B��ec�-i����%uM�A)������L���64��ّ�N�����O���C9;�pb�Nx�KqѲ��%�Jy睻����\�u�E�����%��8�)��z��(3�d9L�Ax8T]^��%���#imԫ���ۡ�up	y�К�:!�m�jl�{/N\�4��!5 �pYW�kaK-����%�G�\$���g?c��ܮ+�|ޣ���~��¹k��e���*���QF�ds�Iun��= �� �s2���ʊR(ޣ��	�a�Vx��j�Ә�/�p35�g���4�<h����8��~.�QC�nܴ]B\c���
���^���?�Ɖ�
��뻉�(<~�D~�����O�2 �B�;7�Y�L��t�1��u�ʙC]��j�j�K�%�K��������CNڞ��%?�uԌt����Hl�v�lf5177zZ1�؎F�ԧ�B���:׍��ysO~��w孷�b{A�tt|"/_������9��hͦ%~�uB�Z%��}v_�+�y�N>9�5�c���!8���QEO��6��d�b��5�UK�R��"�>$F-/��1�e{��ա^\��:N�;!P��3���p\��ׄ����1;��=2��9� 9���Hf�����i��g�K�*hpd�7�X.��Qr���a����H�F\����B�
")����x~���nc��kk��ue'��z����K��0k��gD��SR�-�b�itnk��8��������{a+�z{�<>� x ��:~���J�%PNط�Ur���kR��mYK}w��N\�\Z�5t̗�ϟ�1�x�`���e���%���]f�������z������Js.�M	v!���pL�rzt*g�'|�'09�u��t6����2"X^K�gmkK���j�f6@e��c*���}��jo��/�xp<�Ɉ`w�&�鼐Y�����9>B��}���Sy�4�ь���X��gHaBVjx�y_N�k9������L*0?(�Qͤ����Z�T�{�#�D��˫>i��,>r�}����L-ݿ�)�=!j�J9�;��&�$�c	
z�N�(�e7��F�؋���|��` ����,Zi��e 7�=���Y�f��n�m}e�}��ͬ�\0��{�V�`5�-�`��eT+'5�F`C߲��nІwwv�^q�� ���R�������5M��1$`�F�` m�o<=x)O�=K@��l����m�|����x�^���E��Oj�//��F���\?�����5�N8?�D�oc�::L��|J�3V���Qj A206�`r@bUi��`JO�H&p��G�?4��:9����
�e ���\��Vо0i�������+�0"<��+3�z1�!���C�$�`���3��_=dЄ���fjc;���m��Uŵ�E:�n�c'��I|��M[�4���$�uL�H2����JZ��#��r)u6�T�&��xЈ͓1����m�����T	�ܚ)�|�{�/晄��� �0D�ct��U�L�˙�F�;�<Z;I�Q����e�j���'ӑRC�I�ḷZ��Vt�܎H��g���r<&�k�m�v�.O;�,.L�M���Ƃɢ� 7t�t��uQ��&�y%�e�=�0J�p�"���3��VU�x�H�OY� vYevc����B�y+�KX���.����1��� �a/��b�j>�yh��}}�C�F:���Ͷ�̨�\�EШ��H�hRT6�۩I:�i�Y����r�2�ޣQz>���3֗w�sM�6t���H��ݻr���2H�\�%}aM��7���C@* S�S�n�t��9 �LZ��w��A�����l� MZO����+�VQ�K�HV�齘��:����K�]��Ƭ�(X��Q��UtyC#:]�!܍�,�,��h�o?�{��~���A�-��X���j����%��K}��6�� uLV_|���׿�}ם;w�S��#���猶��	�%&RTVC���w4���2AcBp�흝N� ��.�ł��u����lw`� �{<70V�o\�%�� �ڛ/1U� �@�[__���,��{Me�\&F������ѣGi�x���)=cK-u���.��2+�jL�"��Sl��[3�.�d��,Q	��G`N�v�^���t>��K�v}�%����D��4!PφﲊP�����>�b�`R����dh�)̇���Z^��z�I�!K�&�Ӹߟ~�9wx,S�ȉJ�P��X6Wm��S��E�g�{���F���d7M���u`�	�n��.���ij23�a���������,�G����A�'�������X�L!��� �|�15�v�}�����W���N��ʷ��#�[],�ο�r$�+�ˀ%�e#}X��d�k�;7����.�K'���0�|�G��%�5��
�Pt�檙I� r��|�R$��*��e���aP����������ܽv]Ǭ�7�?zD�jW�s����ֵY������ֱ��s����
l���jWl�*�X�?�J��Y��+����H��Y�-6�Z>�U��ܕ/E;6(ֳ��yK���]ے��>W�i:�;nQ������[b��D�.,U\f��<J��)d/��	��\�Գ��$D�%,�Ҡ���L@1M�Y�Odr~F`	��&�iRCgf���Ō��4��5��J]'�q�q@���u�[)L-��4��a�|�&��
�Q�h:Od�c[OQe���պE��=)X��r#��M�oz�r^��R��ftt��_�=Ͽ�|͖%�L��f���)\���]�w^���񱓷Y�:ѿ^�����%����[W�l� �Y�G0����Ϧ�׎��#4�Ϟ=#����O3�\+A)���Q��P ��D���d��&�<Q�>��&�e��2&H�?��E�W!��gL��U�,5�@tww�	d�4�k�	Y�A��usS�
���`�&����9�'��>��� ˱)[`�ل�3�zQ=��@��~��m[�����Z����F�*���n�7��ʕ�u�%W��g7g>�w�%�u�~�H5�����ϒ�h�Xy�=�T������}"�f��}T^���Z�Q��3��Z�
6�qxE��G�t��}N�8N0�`wq�4��X��J�mЉm�eG�P��g�/���>��x�-��������3W��N��_��
�����	�(ݍ�mwfe�C@w��\ڳDM�9��
�l�r�v�m�ʀ⛯\\�v;`臶��X�X��(�y9I�uS�Ȃ��X�q���n�Q	E�y��X��`ӕ9�/x����.�D?[m�\W�I���܊���=�%��/q��{f �s�3���
����	� I@V]FFXyy��+�O�x`܁ct�v�d��]ieAT�E:H}���:�ܬ�ʼo�?��9cgg�~�p;����03�%%
����@,꥝�m,��J�OV�@�o�(��
���x�P�Y����ܓ�wn�pԝ��5G��+�&�A����K I^[�/\��q�!E����逝t�x��RQ ߡ�"o�%����K��\�Ұ�������В����,�A\���B�(�
ǅ��AJ���І`gn��'�ei?<+HMM?:��#�і&Q���L�?&� �N�nQ�jL�}T_Z��K�@I?�r}#ށL�.{�,�T��5+l:`���x�ԝ��|�v���T�z�f������Io+�j%>��;�D-�KM�t�ܿ&���^:��ʪK��ѿ#�	���q���Z�W���7�r&D|�-������y������֭[���زC�>���o"i@-���5�U�Ҭvj���R:p~��	���yU����� Za�h���� ��;xz� }��v��V��&�쥌�9�:�L�������>�uj�O�'�����6�e
����I@�����}^������g��`P�o�Z�<�����ɹ<Kҋ�SB<j�&��d��D@��S�>T��
|p���dR��N��ĕ�ԓ��������(�������m����Jl��&��5Ps� �
[�ۚP��ŘW��N�@l� � ��U���y0������<�}��Fە�,9[�]���KJ%*ݯʾd�7_�ua֟�	������[��m��'����S��T��%r`�ԁ��}�C�J@:���#�$ץs�݅ G/���[ѡR�i]���X=C<C&蠡���Jk�uȉz �HڪzH�*�j�a�<�!z��|��=W\I�  
���i?�6k�A��QT��w��g�N�cd��UȒ�׆�7��&�}����t<7S*�nS�V��n����e4�/Vr�S�����3�3K��f����Tj:U�v��3���M;;�V)����,_Q�5�obK�2������v��c�����%�bB'��ZPVm @�R�e�Y�����!%O��\�,f�
n��I`c�E_K�i"�۫��4aF'+��l�Z�QѢ:\u���-ӄ )NS�	�̦��)�U�ݐU�_�^y��c�] � N�b�)3�Ģ&�		W!�����G_C�sx��4p(۾a���@��.�V�8v�I:6�/)�"��kM��ˬh(��jaL��g�t� P�6JuC�q��]���	��J��D+4�X�\��zr�<��\���_w�P͢,/�� ����8��Qg�4�R���-� ��`9:;��p�qΈ���b� ;�;��	��Qj�]&�!C@N%�}h8��Ǐ9�<���?���RZ!��Ĳ��Ҧ�ū"O9h�{r/$|�S��?߿A��~��`�W<�%ƚ+6}�&��� @Q�
]N�ǳ�3�3x�-�v:�T�'�|�",(�@��ލ�� OQ6U��ћΧ0�<����8Wy�y=;�q?�C'̹UAS��1�[W���TH�����?I������a����ku��q�0a�b��±�M����>� ��	ߥ��<[&dD�77����V���V�ν�~�a;�ٛ����Ɠ�ܭ�Q�
{��  ��IDATw��d3�x����!���ʊɐ:=z�D&�����G��.�]��������R�0��������U��t �;���a{g�}]W�^��'�d4�Q�$R�.�,Z�����x��@�<y&�}��<J�c��6��`n�u'���HFb剖f��R�?޿Wn��c�h�C6ye��൫;�Қ��V��-"������ظ�����N�-FXJTSbiu&e_=ɠI �[44�H�Z�wf���Ӎ=><�.0�p��	0����!+�&4�jc+eKU7\�HDN�24�b�7`N`xޠ̹�qYZ����p��"��`��+2��tSy~=��Iz-�~�&�"M(��Y��Y�T���kZ˶���wR����7a�#�;/��4�V������}߮�"W�3@��M:ie�
ؿ�o�+���������K
���r�za4ɥN��|��G�>�䌿�o�C���&I,�T%��̊�h� ��%fe��=ӤI��  n�M��Pg�5�d����^��Vw#�<#���tf W�0h�D+���gϹ�urzLi�`��\��_�����^�}�sm�Njs�x��"�L�5龁���ʑf�����������/7��C�o�n��l�SL�5�/<�(�VX\���x��0�����`��!��i��G�i�KgsT>�Ď	~cru�r�i��Mg+AT\=2i�&��z̬��H�Y��ʵ�+ۇ�������>��xҧ��r�����`��{�Yذ����+���Й�<1�����S]�����z
sk���nЪ��al��0m.d"X-�<��/���	]�I��ܢe	���*s����j�N��]d꜃>�1s��k�V����'��6����ޖ~ò��VN���R2����,�/�Ͽ��ˋ�9��jv�V�[jኁ�	�Hd)�Ik;�s�uz���X���g�j�N��WV�17����d�m�u�]ݘb�L":*�
z����p B�{�74i��]���w������H��2��GO	Y>L	���d�߁�^o�5�LҳF%l|5��4|'�Y+ k:6��\�Ä ˓�#���A�'���M�}�g��0Z#�LJ���_+�lQ�`�G*չ ����7ja	)4Q��ee�@�u�F{U��jZT|�ͻ�aqk���%�,�h��Qf��5m1�3g�}B
�r+2��^5y�@r(��_��e|Yƪ�5Zf��`�L����K������Rx�>x��z( O����O�r��XX���� ,�{�.�6�x�Z���J`�44�*�_�H��W�8K�M��>O�[�ںi�z����p���1 �����[	 OY�~�m#�W�����7c���mZ<j�={���� ]�;��P2 �����t�u�_A-�$S�%˚� �,�lˊS&Zy�]y f��W��ܔ�; �1����v:NL6�*��Pr;8���q�z��-��y4�TY�;L3�6�>Z���,@���I������c�X*8M�9��K��N�\X�sG�[I"t}s���΋��e�~���e����^��8{վ��ݹ�������>�H�fQ��̴J~�%a�h�VA�K��DQ��U�3h]�~+ڷέ �9�*nl��^)�[r��-����:�`�n�i� rr>�����C��W�Jںa�ĸ1�����M&o��
�(k���=8x&}�G��o�9ޯ8��
�G
�xo�:��}���]���Ir=/
��C�lK�{��ZR�|��Y,!^�2>�y�f��8K'�}�^�	e�ȴ(���j]m��P�&-�Z��ڀ�&J�i��!�(���cL�?]�w�[@�b�:=>�1�̲>�4����J����t=,�XA�k$;���(̛��
V%F�Rj@b��R��w��`9��JA0_����� (���~w���҇霫I�v�(J-&�
�u�h�O`.��Wp��K�׹Gv��.2�����t��zX����Xy� !����d�?ݵ.�����J�xms=��k�(ܾu��Z��%��2K;eE=�'�} �o���� ���6)E%ߔ��]H|���F��,��HZ�#�,C��`�-J�ƖM��u�͓���(=�X'~��d��Y����#��l ��g�l�@&��%�ѿ���b�3�"L<�47#��3�1� ��������0&�|IF2���'W��F�{�c�'�yR
����`��&������n�ˬ�ۀ���m~�&��9�q?�︧gűv�kc�齲���F�o{-'ᘻγ�ەl���7���%�]�,WNqQ�ӊF��`��t0q���۪o�1�$K���5�K�e��k��в����Xစ�g$_F[=�Z�F�(^�<&HnܼAr���ڂUU�U_d=v��o���	�	M4�1a29���cV=�,n{k'��WQ�@������?�Q~��N���J�W#����	� �.��b>�.y@�T/'��]g��
�1��`�����m�p�V��!z5��w����c�U��K�c��]s��Q�T�V�Nr�v�V҉Þ���e>�U;��&�s��=JƓ�<-��ØLJW��9�
����:�F-�b��2�� {���fA}���ST�Z�2��l��r(,1`��.�&Q%��K�����H�]��_N���Fe��%���l�^�9s��'v:}�-t��9Fr�����%�Z[��N�m��ANƳ�����ƪ@iY��V����<[n�̎��Ȭ�)i�[o�g���gF��0.�����:���?���C� (� @� �7 t���o�IpAǈt|���ر̄Ώ�g|~`It1{����j@I��z]���ޛGri����8��.V�uK=�ݻ����ٿ{�~�;-iZjQ�D�H�Q8yD��g��G �꠪�t)	222�Ï��>���KK��y�m<[�5Sz�-� &?C���&G�F"��k�88����h/Ok8�gs8P��+׆M�0�u�#��$
�x�>(�N ,����~���T'̼� �BS�y�Ł���Z���-j<B��n<̵Un�Y�������	��Edc:|%���,�S;�}0��D,@�b�kϵ�ZK�����JN�{���gY��^ˣ��`���}�3�wm�Y�gb^K\�ʉ���5�=G��f��V��<��<�~�����c � �ө(+ ��yS�D7r��J��F"��}�k5���v/�準'<�;����_>z�Dt��3̥�٢M(-l���� x�R �p�I?ܼ�y"����+�֝�H��O�}�)]y�
�yHe2�ae��*0z�x%��^�K.1�$��Ik@�������WPTt�P�*j�&��R�s�m����'���9���`�1�6�����4��c'��56�c�du���FR�whg��Jx@k,_6�ЉL?$���֕�g� �%U�֓N���H�Ha���`�dH�T�a����_O�U�*��	���4p�N���R�>�X��2(Ry|� s8�Şz�jؑ���� �g�^PD��f��TmhU6�w�;�������Fл׃YW����k�"�k2�~�Ɉ� ���&��d�K1��TI���W���}F׮]��kF�2���h�,\&Ę��\�淿�?}�'���u���zoDi"n���Y�r�-��s�Z�����G/~��%�;"����~�)[�����D�����l] C�X�t��%�(���/������Y�}�Q�B�e��s^��٦d>��>���8�[��~����׶/����e��Y�,��� W�����Lk�{Kh��]���~u�����,��Z�[����MvN�5�w��na~y���[ljL_�d,ڰ��+`�
JX/�c���������u�����0u�ЄO\�=�g��ƥ�5�C@t���Q���_���u��_�+�t����E��Ӊ����sŞ�g�;���Z�T��ʿuT�]Qt�Z{��).�&�Me����>4b�(> %�+��;0K�E\�����<�*t6�dM�+�Q�z�I�M�����+
!z���>�05Ќ�t{���@��&w��]��/��{I�I{��8�*��裏>��ػ�J�(�h�.	�>;��v�ƴ�Dh��*�c��oU5�h����d����*���1]���<;���R̎2��/��l��dP�0��	�!q��A3Ƣ.��������c�x�v� �#������	Ur�6�������E��".�X����<���@V=���
��X�7p4���R ��p͍�7�]�j� �%s{v��q՗���ۨ�4[ "�N&?��-$Q�Y��&y�lJϼ��&@�%`v<>��̅.�" �)�rY�?K(�0���d)���O�oBy��w�W����?�[�Hb�*WtQY�i��a��iÇ�{@��G�!�/���~�;� o.u��:�yb�'��Z(�7qaq�߇t��?ލ�;��`�a�6%
X�\��$4�'�H7 �_&>��tM����f�7��n����K�{�$���7���L�K����d�fB�
��j}�6�WA�ճ�\�Ƌ���Þ��JA���pl�8M�@�$³�A�?7
��#��bNO'�<�u�0�VP�Z�G��Ӳ��ۃ3ҝ���:�%J�a������<V�ӵ�ޔ����۞c���f���It�2k�{��x���\��[=������e���F���ˈqRh��2�؊V5��jx_(��qQ����J	v!"ߥ.��q�++�SG�!=��h"�l��7�/̛-e1�V8Ԟ<^�[����n�ڳu>�$��9�,}��/ؽJ�/���E-P|u��꺌Ӂ�uV��+žpQr_���cW�A��Л-�ʆ�"�][(�*�i �^p�0ư���3�ˠ͉� �M�;�
5��_E~���(,|β�s��z���.���3��ܤcKS�]���r�U�7^K���H6�5���@��M��Q��n D���
���%��M�
`v�� o�ʀ��s���sH^��w�{�u���NB;RC�����SO�3l?o����\z=7l�rds�m�%7f�R�j]k!�ˡ�Z�[�wj
����}'��F�,�u��E���g���E��Xe�z��X��¤��W濾H���_�����pg�:��󗬣�W�sw�uB�Nf�w7R���Y�4 Z�+p���2y~>�1�3\iN�ɵ%�A�Йίxz�J"����j�0����Ea��Ġ�����-����\�������c/�X����<\k��nGu��X5/M4������W<D�g�'��tno\n��5̅sy���b́&EoD�{O�A]����EZL����ۛߘ��$>u3��/pVw��x���$QU���,��̘k�F췾Y���g-M�B5e�b�G#0-��#}�g���rIA�@�SPj��}��D�'Z�!�676������a8Ճ�����E^��,r��}@�o�eO/��pF!G���Ν�k�ޡ�׮б�%B�Wj������f��a�;�J�bMa$ʪ��>�RG��yqh���K��^�L���͹�3��$Օh
�+�DTiS���d��=��id �X�K�ς^�N'�-Pn4I��AUK8/��U+,$�l�X7�
hX_��� bC��8�^�]v�OMw�OY�̱GWh��>��B@��nrf�2���|�Ϟ�ޠ�B�vղ��jUgT��6��h>�2#%�%�=d���,�4�s\� �|(>SN�լ�o�1e<�,&.�W��=h�^�t�>���`%^���+^kϴ�C�<�9� `�O ��'�B���?fM��׿��&�o��=o����fT�ЗS[�r�  /�&��L���C�Ҹ�uL����87K���Em�.w���*ɔ�$k}��f//�z�J��M��87����Rv�D�����P�OӲ����Ȟ�x대�(1V�ό�R���d��F������Z��XM�̋��`���,�÷v�lx�^:\��^�p�����3�}��F������B3�����Y6��.����ǈ`{NvYJ��3d�7�QH�	�pN��Y��V=��Nk��Q�v�78v�2EZ�W�W���Z����1hM(�U �'�]�����/pe���W�F��J�@����ݻ��?z´;��Ĺ��e�t�]�t>�� �q_tC�K�U,���4E�5RH����P�q�T��q^��Ĭ���ćm�ş�e.X����Y� eh=sOj.�'3BD<�	���1��`m���go�L ��a�^�4�/Q�?FM�HSZ�I3GV�aI֐��d��&���6__C� nwi�@�o�h&���D��!�U�g7XF� xح���4��| ��Ks���,!x�{�M�v�
J$�yحqRS��D��h��ǡ��δ8���e����Ŏ/���yt��Tt[@є�p�xl�� P�r�
��G�S��~�:W�a�Y-;�V��rvϟ?O��.g�T�@���ϟ�Q��z��B/�xߝ~0o��.�7NԢ���d�kk�c ��v��h �l�2�'�)P͹�"u%�Z�b��w/ɓ��D�&�x�vQ���v���?��J�y���( �ʎ��c�DYM�Ӑ��R�Rx��ͪ�e�e^Ó^y���&��L���B�F�G/K�V�cC�����Է�y MMft��6G�S��������S	^�7� Ǭ{����G��t��mJ�I�݇
�)�-��ũ!��:��*0�qb�BR�A/@���j}ŕ�N-����_q��"zt-/�����-Y
�8^ NG��|��w�s�����I �y�8C�O�ZV�4�c����uz��=y���7��P��W�^�s�Ns�r�.�痥8��K�b�L�lT���!��ښ
v����*K&cj'y�DM�@+�'�ܳ��dƿ�,��T=%��d�'�����7�֠INX������"\} ��{,�z.]ˡ�!���{gQx; ��v�{Qq��%W�������Ԅ�v`��^[��N�k�E�i8�t��ᜮW�`1��~)Z�U ��g��6� �^�}.�>����J�d�<j��	�o�L���6ˢ�3&Q�3�9��E�_�g����nL��ib�lC�WF���h��(�^��d�)փ�e/3�o��BS�/�K�Hoҳ�g1�� :V$���Jo�<�A}-�
}O�ݝ�M��`%TKMnD)��ǣ�X\�y^�2���L~\���v�s�PuCAL�2�]��c/��=�6m�G�[�*�Q �a��u��;�a[~-��&�NZ�ۯ��;vZ_���=Ay2OL��S�j\4�@����o�:�D[lH�$��aG�1Y��5���4� �����Sf8 \��{ޤW��~noT�����qɋ��������:D�99�����==X��3o�`�TЗEv<+�Ԝ�^UE,�P2v�:�:̜��ȸ�z>X��ib[�s���t��m.P���{��qN��/~!�ᬓ[�r�kk�R��=do�9i���z�+��>}*ͨ(�y/��Dj�.��J�b��*���j���dZ��r!|��\F*+�J��)�P5hEܞ��'Cd3���z=�:����B�'��^
��g�(��9��A�]*�y�,�Ĺe~��WJ���Q�|r�8��9�e��d�~��<y����0i�� 2 �x=,�k�����i� ��&��7C*M 8%WT�1��1�W`w��#���2=�2�G2�����K���1�Ib���T���_w��¸և��Kr�&EW�Y2 *���7��KM2:�Ƚ�W�pZ�u!J7�~���	���R� �,΍
gب�M�$"��Qk7��@�@�yP���`�KW�=֕�Q��ڱ�)��"j3�j ��r�ܭ��^�p5j �g�Z4��x��5�^����s=/���B	L�����3u �'7=�v3@�6b�2�Rx4]�z~��h�⚋���=���9MFduYL!o4G�l��[���M��^�?U��:&I��7%W�����9�(����ۅ{�̬Q8�u����>�����o��uIG��:����~��X{��!�9��4��{������{���RЍޗ�����I��,�x��ɜ�������M#�`�,�N��M-{�nݺI�o�b�.��cG;���<G'Ƚt�]�v������U,x��re�0��&8�B�ډ�B��zV�
�e϶�M� q\�S�[2���>�:�c#��ULv&��XMD���Y��0$u�&�sR���>l�bVF|_�D�ɕXe!�:�#��H��D��
�]
��b�{���L��-��Џ�T�<M��T4}j��)�*k�gPQϓ��#�`���4m�x�F�[�xz�S֥ۅ8z=&כ���z���Ư ~����d��@(HT�ʃug�x�41O��Td��\�g�L��f�$��)�e���1��>M�l.�Mg�Q�	}���%�3��iԚ>�Ӓ�}�Y������;�,r"���?��c���B(��	h/(��}�Zx��\`���[A Lv��LnlVK ����<��7� &�qvs0j����
.;~!����&����Z�HŶ������e��G���2r�t�ͺ��\o���8��9�j^S֊�M	�r�Ln�6"+� �s5���ٵ�͌'3�
��Rʓڨ���Lբ6�B� �S��4��Y�Օ�lx���l��޴�9��XG1_`p.-.�����מ>	�y��چ����^��Asf�O��f���l\�:���E���u>�;G�������{3B��oɣ������+4_G�{y�=�)�Gu��ܳ��Z|��^�����U�\2ʜy!ې63�bA�N��n�FB�Z<��D�e0k����v,u��8�d�/�ԣ�J'�u���F�Q�rg�|"��<��7o�_����!Q��ڸ��(|�qN6�t�B �K�0/;)6!�����"�$���c���Ee����x�]ɛ2�)���#u ���T)��.�}�#�*�832�^��K39��xJ9D���Zp���YZ��m?G��T�5	\��vK�I4L��� ��K����gn���x*E#F�jvw�U�/p��(\P!yh^d� Y��7��|0�����:ml��p���`���#���v��XW�_pE��*Z,��h��}�^qi�k;{��l�����$r�5g��f����)=g�>�7�&H�*UN�<�e�ov<�%(Ѐ*V�����܇�\�z���,DS��*x�^�ʚ���8WY�{�k��W�B×z ��##*���ь#k��Y�>����{�(-z�f|�y �����6嗡4X�IXYy�\V�U\SnL�
5�Q`��M8�����l�ժ�,��j5%�ƥ�=�l�H�t�/��x�ю�2�M���x�Q��-�tM�]8�����w����d�0'�� ��S���`(>z�����;��<��71�&z�UC"<��^��kE*Ɍ�l��������SH-O�M��>I'ϗ�n��^9�C�@�O���T�j���֝��b3u�x��赟]�N<�۸��X��k�0J>&����݌a�S�k��YJ�^Ǵa��Q�``����%�Hv�y��PDIv���p4���^�N����h)�D����V���3��{��칳�������g�"I�RXO��b��a0����hzv=^��ҽ xJ��*kd����UӸXu=Ξ@��'P����[C�/6��� -�}?�ox��"�6�3��c�IM]2���GЋ,���Wʢ8xm�p b��r�lY�P�Ͽ;�	�����O��]ڭ'T��C�`���6��
@�os*����ܰ�r/���j��F��	�e�vâ>�3e��~�cz����j�����N��^�1�n�B�&4�4�N�x=�{�>��}����T�Z6����V>��-6vȨ�J (}��}��Wl�BN����O�20�s�ܙyP�w��(	v��n����:K!�M���wm{9�G?�aZ�Os�nNհ�{��;�Q�1~�E�]ZY�'O�'��8��ia~���H��wB��,:�\�|2M�m}�����L]��:+�����[��ra�}IE>Rp��E�^V�x��?z���S�N�/?��Ο?��v��]�ᇛ��ŵ`�Z^`��)6Ϝ=˞����������������a�haqQr�Z=J��5%��L�lZ�fE'���}VF�i��:�F�O�RN߳q�������6���e�w���訏֜{�_��o��C9��:~��K4JT5�#KKNV'Z)y���Sz���#�*6��З �R���W\��0o1Y�P{�j ��_�o�o�ߩ;V��M2M�ۢXb���Ⱥ%�Y���W9uVhM�^�h.yzc?y{91�G5>�%P%`�:���+�C��F\����f��?�����v��0 n���NI*�:K�4�&I� �ͩ�%��C�#�G5+,�P��&���*#nB}U~7XF���������M�8�}|���֓
i؜��;ʂy���'�&��(��yvMO�@`�{;M,�dxx5=���?7-r�b���9[}�b]���a<����k�L_K�F_6h����
6����������m����Jy�-/-��¢��^��8��'B.�;�t��m���/��_���<~,�2u���K��NΩ��Y�gW	�m�X_�7�E۬M����S�SG�w��<��{���M=e.���*]{�*����I��}O�(	\ɜ���>�-
Ѩz	���"����jdmc��4B��J)t ���bM%!zμrqw�,(��Оf�����s��� �_Rv�V�=ǉ��Νa�<�6j�I�O�����'�`�$�Bd�&�{a:�z}�o�-K�^J3�&NU��f8J�{�;ur�=��-����usZ��$����|௳%p�������n�����X��6S��&����Y�
�o��Ҕ���J�s<?�\iM����Gc�%��u*��o�������?cN?�Z��]:q�8���>��>��#NZ�_��FV�[k��b��Ԝ�"���]|k��O�<�� #s�	AC��9]�c����6إ���:��G�r���p�\�d��7K�o-1��#L�w���D2=��mK�+���0�N�z�Q��eȋ�	�UX��)�J������]P��P6RA�����00{����؈Xu����DhF��P�����ޑ��X��U��,a&�pE�o1k13�����9���sCg����F�/��Q��w^M�L�2!!|�����g����R,ހ&�`)��������������?��S�j��*kEg3l������TH���f����'p�\oS{U����.��Y��7�����$�=�\����W���"� �������{���s煶���"jaʘ��ި����F�<�| ����z��� ߢ��j�8�^���5L��֪�P���F<��st����AA{������k.8y����i6ǭ0�~���v�!��q,�7��N_��5'�B��HM�~�:�Yt����ɏ섲3#^V���L/�e�0��O��N����"^ʱI�}�u\t]��3������"��k�a��V"�J /�+�e"�\_�1�����\��NC)M!UV9���(+l�v�q0N�������g������uM:}�$}����y��W�^���y]'r�[�H��77�~Y?7�Ԁ�Q"!��ɉ�����o���gQoo5��ǘ�X�����g��}<���1/o>�Io�.��zіa���[;\V7(5���|lUբS�
�x�����47i�a�&VVүK��$���2$��B�'�o�xV(�-�����O]�a��,L�{&�~s�|�spٿ��"���6��ѹY�t]�^/I�hYI�F�]z�<Ľ�l�A*���BIx���uϝ;ǡ��'N�> ���A�^*��?}�?�*�ݻ��|F[�����E�'��Z	`�JX�(d�=��"����-P�ҳ+�z���k��G(��B��:�A	m�Yfv�S$rQ3	�T�nߺA�ÿ�����1�>�$��= �Ln�H[Pke˅��*��N�9�u�Q�W�8i����.�M 0��8�H)\Lw Qjx��!�;���	�(����.(�?��[;;��A0�o�p�F��'����x&��/�e�����m-w�F�,!�����չ��YCȜ	<��Y���2�c�{H�l�y�a;�{���]�2��'��΅�=ҽEc�/� _�C����H`ckF�D
�J/�ThQ���Ȳ���ѝ;��?~A�^�>�OE� |vg�C�O��s����F�|�1�+���#�)�!��EDI��eG��
L�q�V�(m�o��*�^�i���k�k
�T�<�FkH^t3������*�����%�`n�d�N��w��GeX<I�v �Ͼ����%��o��n6;>?�Ҫ����xd�4Y#%��v��稇*i�1��
�|+��Hz��Rq�dY+oNC��7���N��f\kM�ٍǘ����:����݀��*oOn+�����k�4>��L��w����$�H�d�ƴd2{N�Å�7�l$|g{�=J�?����J����잤�'E�Zh�����1 �Hx[/x{1���E��U�iX{��M*�zus��������E@�Q �8��1e���2��(�d/+�!�5��r�mޖ��`߭���`$c���b�������/�ۭ�ѳ�� ��*����
r�҄Ѕ"9(�
�J3�����<�l�3fy��b���M���6�5��oݢg�k��r��+�ч�e�v�ʖVh%����~��z��Q �SZY9.�����|6 t8iؓC,%�r�o(Y*�9D"���۶�u�K9G�t��U|�l���Þw�U���A����u[�p�������O�z+�-b3|G��Giθ�3�l�8���>:Zu!�����'_�]>��}b��tjG����~t\))��i�	r�wK�0�RL��Pg�{�]@����sr*��y�w�Щ������+K�4:��؍�w�Ka�ezEp=e�����O��"��Wj����U2(^�����a�͵���S��K�K�Z�8�"�Qd��*u�g��6q�E�d�ZSș�2�����) �|#��A�8�<Μ��(���O]�4kB=�����ϲa�Lt#px9�����9�D(V=�~�dc��&��E�'�s+N�Y�Ӭ�C7��[�ʭ�| 6K�"��jp�u�e?��[��>�a!ל�;�����ޓ�����U}�vl���b������^ �LK�o�"������Px��ȗ�:�Z�Vf^���tqÅH�=��,f�0�]n�D��M~�^^�����&����~�A�\�=?��*ˡ��k�5 S�ǒ��,���+�3~}~�9�b�����y@�w�`]�w�f8�P�E6)_�m�i!�Ĵ��Iԍ��`��;C�@����=|x��u�r����[Il�ITIy�^��g��|��Is\�iL�9?�����t��.�	;���rl���o|�=ݽ}����z0&��jI��ϝ�˗.H�� ȑ�˴� x���m�`�5~}�O0 ūOQ�D��)qXN��T�ش?�Ӵy�}����z���7���*u+�Dl��嵢S����m��-��9������n����u�;�O�vWt����u�9ܑ��DD��t�"����̛�k��H��:E��U����b[�E�Q��Pi���]��9@��O��#'�ݽs������¼��5���O�~�k�.-.�3ͩ����T,[[�	(;�z|U��S9�Q<{�A��ݧ'O���j8f�/�W����'k�Z<�m	�,��d�=S��P��~�s�W=H��|IoIi���R�-^Ro�;6��離8�9Jͽ��~���0���2oL��t�.����±�G77�2�a��'2�Ao`�ҹe�۸��X�������(趣ʉ�(Oѓ�e��Rt\&�W:���XOQ��]p���$}n?07�eݾ��5�g{g��)&��a����${���U�J�%)���N�첍R��y���EO�Y����9Q �>+{/������P =ߏ�g,�2��jw���XxG�% e�s�>}�[u�Z]܌|#�p�3�O�ɓa_]�����(�� ��hcsK�/�N?\'@��U��S*��$�m2 ]&�
xdv�wēZP.ry�h��q�V�W�"&<������׮�P8Ŀ�x�n߾IOמ�\E��=�����t�"]�|���Eib��vkk��m��W�-���Q�k5�#ޞR�AZ��j�)bjd&5���-sҥę�w��"7>}�K����<x�/Y���&�(�]���v�w�>�޻;���㟳ؼ�zx�ϵv�,zB�o�u��.�M�>3�K��[���2g���r$��<���nhw8�7ns��7�|G��=ss'��1{VO�:�*-�~�	}��t&����y٭��}��5Y��AW�Zp��)Z�?�[[���9�������_�a^����YŞ^Mm��i���
uh䣊�Q�$���&�Μuf8�Ϧ*]�		�e�S$P��^�;���k�B�MT�Ά�O^��ԝ	>��D����4�"�HV�&e��d#u������W����YU
�o�k#:p�g9^y<��o�
$�8Q!��2�m���}g@z`��:bng�L��J�Ό�~���.�����/�G���E��ݱu��cV� C턷Xk �p�'
�QcN���u�����*/
�D�ڳ�K���1*�7�f^���O�I�Y�Z^zƫ-��F�̳����q���T�ܓg �`���j-���6C��HE�2��D>'�A��a!��;:�������]��`Ij��i {H�-�ݦ�w����&r��(��P�J>��W�]���k����O�������6 �;���3�3���#.�]��P���ؗNSO��<�-��=���N�z��y���˿�K8�i
��!���0���O�p�;�\
Ǎ�ɓgt��E����Ч���.�s1,��&9���?��%}��\����բ�i�̖w�5:�n��-O�3��^1��PhZ���s m������B.^��9�^��o��k6駨��8���z��O�u\n?��j��\r�`7͋;!�S��&Shb�-{5e-%�	�Jy"�&{7EU5�h�h��m�˟�������~ ��#v��\Vu �g�O~A�������3LO���y��T�1���"���j.}Z=��;a̓ܧ������(k_��Ξ=Gs�`����7�:�)0T�x��{�7q�ao7c��1E��e3����ld�֪m�&�&np����Z	�GR޶!���-*��/\
�FG+%�%sF8CV��~�T�.��_Dz��7R�i�w�Nj�L�" �2`hY)>�y|t+�	�����E0��d����u�9���a0�F��	F91F���}�ٙ(���Hkp�ٗ��U�*�7�0G����vl�bB�i�ӷ�oз�ޠ����pnѺ�7�������U�6���x>��]�{�<�]^�O����i�y3M��ͨ�[a�'왮=$<n���|�$� �z%(a�����GШ��T3�|�h- �gz��w�Y M;J���6S��5l\�r`�X\\b�k�ŘCO�z��)�܅ŅXB0N���(Ô1c�����hRx^]�Up"��t=l����y&�&���ٰ��y�"� ���o��m�Oh�+�30�w��kO�8�)���ɧkP��3�o�q�a�n�a���#fH��՗p��Y�N�ë��;��\gTo�~�:-�<�'�U�Ri�]���y�Z7�6o-5u<�GXK��v��,�T�L�ex#�����yF��"2�|���bYJۑ�M�.t�N蚁(fE�����h<�ٳ��w7��/�J��6��U��0{��Y.,����'�~��].Q��h����t�Uy�ij����91������}Ρ��y�և�ҟ���ɏ>���]�J�K�\�����VxJT���QǙ�YPf�Κa�'�U�����x��.�� ���Lt�=`]��R֥F���a(U�Iܹ۹5�@O�-`>j���`Ek���Tl��^˞����_��2ˢ��6�vo��]���<���'H&�h����j1��G^����Aћ/Rz0�@���ɞ�pu��`Na�ʛN%��E�(AM ���gk4��t�����[����[��Hf�^y�7d���Ov�P�tE�J|�n͞hr��.�������������s� �%�ߌ�m���I2o� ��)�f�Q8�x���'n�;���Nwæ4d~���w�&s;�]H����hA,pA� ����M8Z>v��}�L�f����
��'O�ĥ��&�'�d�p�k���X"�E?
�7�13���xMŵ�Qf{�v���Psu�;�H'Ng�k�{~�$Gf@���q��<&�t�VVO��è��E�D�4{��u�e��n�E��e�R���=J�))�J<C:����$�x;��qd���x��o�'�|��A��v�8Y�(wX���[���9�m�e��;�2�������u`m=�q�O4�h����f���pS����q�rZ�,5_�)�=�Fr�PI�����U�S����==y���毈�ر`�^�t��{�]�%!Z*儉�kP�����'ir�ݳg�7�0O׮]e���p͈n�����ƽM�(U^��􉕕�nQĒ�M5��EC�Z����}�_�qjTnZR��(lc�7� �ŧj���
��d�R�2�$<`quk���W��u��#�.��b�,��%�Y؜"��6�*	_J/)�< .����b�ir��Ng�zJ��^�q)~�$�X��U_D3&�s ��t|����t��Zxo��f�H�x�Iܘ��A���!!m�;�/GWGQ���>����Bc����r�t��A���{Mí��{6�g<Q$۳�����,$�[�W�%����6j�<���{~E��4���F9���-��b��Q�ϼ_g%��L��*B���f��2+٬���"O�՜s(ʌ��e�076 4K,�W����4��X*��4/ ���[�n�w��`j�4�VΤ.+���Q�����3�'\8�XԱ�c���e��c��>or<����y� �/�.Y�g��N�
��Dp����~C�֓'��z�>p��I �㒗$�a4�2~�����	ܺ��_|�.\|�6�6��`� T�0��dc)����K������y�`>�E���z߮��Α��#�ѣG��������O?eO/�����:�"uD��9Β��O�E
�+(��P�0e<��KU9-*�D�F�4���K��bzy����>c�D( Éy��8�JB04�Z�w�}��9���:��Q� QQJ^���縺l�xA�S�A;�H�w-����Ph���0��Xk��Ν��4���W�a����++�.I�^�6�.���K��zr���U���6nۦ��!{!��2u��"����Ҹ�$"V3��������ߍ���>� ��h3Ծ���'��%�(��Wa2japX]^�"[C�Tl@�R�@�K#F$�n
=���cR��3.�p2�*%nr������*�hvA��lg��|W��O˦�����D��<[�
(�(Y9P�6E4�`��a�z�ƒ����C����,�xaM�&��p�V�dZ�5mo�hg�1�l� �U�;����zo6X2�9*O+����4>Swx{�-�u����|s �s;M6&�ř��=��=�?vˁl���m�7K�2y>�{=��9f�A�X�fH�+XQ;�IP�s1<o/� �#2�I!L�� [�,�!t�BC<�xk���� ə������a-}F�[����Ik��Y��Ҋh=�V�W'��qgg��	f`�$Q--�=͉T��Ǥ$�zlms�Z��V�Lr)-���ɪ%s�"�h��fo�0�������9#[��Rh" � ����v���Z�Q�
̈́yzE)ɾ����VNP�k�z'�Geܙ�y��4i�t��ȼ����	�ާs4V���a�-�\d���$�C4T�B?B��;��L)��Y��ï~���z~�~o	�{� ��G���8�`��b�b�q�ڟ��M ��v�c�"��[	J��I @$��>��7�㱿��1G�x��=~������	��A�9�s��F�X�{�� X���#��wV�ȟ���t��Y�%��0�;
������_|��*�.ݼu���pw��aa샦����3�A"�L(>���w�Ab���*_]�5�V�	�	�#����5��z������xBw�?�,b��~@�`�/X�^,��"��I���U�aʋ NO\꽊%�C��b^RdA,)w[�,U���pw��D�u
`ao]-������P,?Kn�"B����⛰XGgs�y�b��� ��<����WrA��F���a���%�t�����V/��}�1,K���%���̞!��0��7����P>��4��v���4�M�[D	�S~��H��\z|2D77��譙߳��K[�;��&�?粰2tM��[��>����t����#e��-�l���G���-�1��I�D �{�"��ᬍ�e���b��>��4�/�)�zq��*U��8O,y,I��'��U��w���������l��
�k�йG1��2��2y�Qq0��A�ʥk��FԊ��d����z�2����s�/���
mn�0N�g^z��#p̳\�H�Ua]�F"��$&a�Gz0`�{��yz���EZ����%ޝ�EU��K{^b5��:+ �)�{M�P��B�@u�F#(pj�����%��B? Wʆ�x#�	P<�S̒lU��^j��w}�)WY+�(�h݌y׸Q��$(2�M�t�8�����L��Lgkle�q��jۤ2��� I����O=ތ=z@��t��I�\1~��A��i|κ�K��e��Q�AT����:8���B�Y�f:{�5 �4�B�9��Ā��U׺���o�C#�V�6E�e�m4�l`�"+RBX������c�V�|]�w�&�:�;��2�E!	���f������̈́#9�[����\X��Z�J5�u�5��ر%��/?	��\`baaN}J)gxaw��g�.\8��8!��������n�����'O�J�?b��[���E�u��0��?x����?ҊnĆ��.��=0#7�rU�	'��pcB��oҝk|¹xq�����:tu�otiy��}�����;����>#i���	���LV6�H���of��A�@o5���c��D����@n���G [b	�F^���A�G7b-I�"-�Þ������B���:*��sx ס��ֶg��V��f�.Q��Sk���?����
�v���feI�`�����,qLY���Q*�H�Bbk�v�(p���x`��y�LX�S2ާa3����h�3f� /8"Ն�W�o.�EL�����w\s���đʄ�D��ū$�kℚ��DO����Y�l��a�p��Ǥ��ښ���;��Lsɬ����?�ZRW�s5�+�Yh �bt�Bir)f���>��,v/�R� %o
aM��:&��u�ֲ*%��q6f=Z�'�<��l4=L��#a���4��譇yB<�1_ʳ��_A[H^�>-�����9��P���'hu�xXk���i	=��.�t���F��X���]�7�)�P��yx�� 
5{qk��İ�c����bxd�i±0(�@�b٘� }>���K�9"�]-a�<��x�S�Z�����x;P��-�l+�cOK�K7�E54�3aae�oC�G߂6�<}��G?����^i;������hm�5��o<j�A%
1w�#A�����mh�Ҡ�N�K��+WiyiE�e�^=R�m\����'�+�Ir�}E��F� ��u �%;>�M"�����:䈏��1�Ղ��;�\f����3t3 ^x����$Q$�OÚ�T�e2��x(��ʒie���={�� 9V�R氪�@�!ˣ�t�
%r]�a !k�����uZ�x����+'e���=F+����R ���ZXZ`a�9>f���ԟ�ԯ��.+/��Ak�v�'�y)�Kz���`C����O�D�4�*&�S˽��j���KF;�՚��(����UKq'^^xC'W�SZ� 4d̘�� ����FdJ�O��X�Y�h��tQ����!���<�n�ߵ��H�$��]-���k�g|J��w���ǆ� �a���֒���u<���mLí]���q�K�;��|�[X�i&&6O�;X�j�H��T_�"q�W�;�Y���^�W����@1�k��s��pت����sx�3+���|���D�:�ժgC�;����s���Y<�F�ѿi>@��H��W�Y{!��@y YxB9y��߈�fE^��F
48� h�L7ۥvж��DQw^�ހ��Er��&ӆ�>���65��½�~ n
H�o����VW�өS��j�|�XP����;�f��K��nwW�D��Q$����XQh�5��2A/f�#Z����9���|l�)n�S�cE\8v撼 <C���d����c���K���a�[�n^C}�2B���u�h�z�*q��\�S�n֍8��z;�Q�&��7�~�ɢ���$8�HҞ���W��\2��ϐ ���3����h���{�ӻ��!�G���E�T&D&>��ɅAax�!XH�G�:�e�\�XD���Lֈ3g΅�K�hp��+�KS� ɵ���8P�P�棏>����7�������� ���k7S�j�+O�`��V=�}������/���"�r�Ĵ�v � ���d��]Aӓ);�ä���zxMh��N��7hii��k�~α��b �ˋ��9x�'�A��g��	�O�4sC��k�(��.y��|�:���&������� �E���y�������3_k�J�*��6$�<��c ����k�_#���u(s�Wv[�~aܨ�q�Yb�����(�FX��7X��:N�u�k����arLG�'ҏ�������\�[�v�;eO.(
��vwG��������\#���3UP`�c-KQ�@k�%ސyASh�<�7E��W�$�7��	?r����	 ���	|��i�@��m�v�v�WO hX�p����..�hQ�#q����\����bmc��}�1h4Js�Ή�'h~n��GQ˴/t= Px|��>W�B�xP��d���ؚ�g�~��6�Y�"�<��h�W����P98��K8E(�¢j�|ؘVWOЩ���a����d^�e4�Jd�#�����X�S#M3~-;S�:AZ�H��S.֢eu�sB�����	N��^�����%�%ժ��S�f.��WT�Q�F�7�o�=CB��)�m8�B�i&_�|�p��(D��/:S[
�v�&���&k��y���|DDG�[���[{[�S���|ٯ�"���8ձ����q��wG<- ����Հ=�Q���؈N�9E'O�h��8�]^��A0�ϝ?Ǒ�s���P��V�)E�<�����;��2$	�Λ_�Qls�ץ���,��{q~`��zoؐ�t�{y��y�wn�8(�3�����W�왓t�¹p������ɿ0�G"�X���>�JkU)�Kޗ��� x'},H�ה��h'���1<� /.��<� xye��WG4@y<�Q��>\��z�<���C�E��1�Nd$�20���W�؇LwҤ*dA�r�N�|ּ`�ф�d$��s���4l�5+W�������S�E�E�Z��it��X��E�)Ot�'�JP�R*��+��1�p��������ˋ�^P�n�3�,IL�q �S���L��0e�B#	ic�����x�	�i�ˋ���9�4�yo I����͠�*JWٳT�ܴ������g�h������{�z���ġ���oK�JY � 	u��Ph����ؽ|�2}�чt��;��"��9�E�2��T�z%K�
����hep+U��3*��f\�w ē�O�� �J���Bj��!ow��=���/���[R��X��u$:t�"G�ԦG�ų�����9�0PD\�K�lp����x GCY�c���O�<�c8G���mBE�UQ��0�hRȸJF���J�JIU���S�tJS��~�t���g.o�?GV�Ij�8��jxv�%q���l� ��ޜ���3�A�.f�+[� ��Pm?>��i$��i��:���<�o~��մ���s;|������\�c�?үb��	԰�։Ǐ3���<����p�N����sF(����B���������Z(-ZN�\Y��6�E~�T-�0a�[sz�J(הF���\�K��h�C�Q��-J���9�6<Ҹ祀9A��:SUBCt��lmnq9cQ�x�$��������@�b��ٛ��1��
\��|PV�]�  nl�dJ<��q����D�����{�|�/�O��+ۈD�^�ɳ�
	�d��X��)_��n쉙D�Gt߷8����H�/�	ke7vt��+�x:�^WTV�S���X�ּ+eY�����^d�����=$Na�/΁���)H���QJ�F�ؐv�O�ގhw;\��H�Ϧ1��DpT3o40¶��/�m�H�w:$��"�ϠF�<�]6��F�fOGy�[���.�}�߼��7�OR�p�EB&,&3�&3{�2 ��6�C��{�=��������O�_����j��'L�%Tk)L+l��*���J�T<�֟�a�/��K�F+'Ņ�2@�2�%Z�����h6��f������;g"s�L��/���#�/) ��?�3^[[g.�^�\����$0{3&�Yn���saS;��
=x�0��'<?����դҺ�T���*�lT����HB��k�gu��M0:�!�F_�{���Odd_=Π�4b���g���ڄ�!���L'���@�Ϝc�����jO�»+��
0��E.�Pv��s�������Y͒���Vj��DkQ
�F���<q?�����mI�`o3��x�Ѫ�����7K�c�.�MG^���2�FTUO?cQ�䜁��"�"�An^�i�ܜ#0eo�h4� ����N�w���g_���z�Iz�_v�X�9R���>S�̑x�T�E��D�޸&�n����;�����f>d%鿽���r��g0P��%+4۪1Y1�:S��1{���	S!*�J�2 �.,�c�橄�%���eA݁z�Yi�Z��m��dN�I�[ŭ/ޡ*�����+��젴�2�>㏊��7��Ҏ�����SU�,@���Di����+c2��^�|�KS�Қ����H�)~��x|��wYmyxx�3��d���zd��6vhgK~�݂�W/���R3.��u Ԇp{�mX����"��!�ˆN�. ����$Q;Hy�q4�����F̏������iE�],���Zh?��N�Ւ��DR n!V�j9H$`U�����/�)����z�L5RO����7�U���r��HQ����6U+U?`�Ĵ�s�<ᙜ>}�5r?���u�&���S\�^�^%�l�&vZ���B��fVYK�E�W	�=���<���c�>/�%�Ie�#Ue���+T��Z��3��txl�Kjɭ��,+�NꤠVI�"�T	U�)_�r'������4S^_EWZ��޲A�S� �;	��(�<��!S��W�܎�'�ѩ�����Xc��S�*$����0�~n��,Ő�{pM�+��b��bK�:V�Je�<y����ٵ��j���l*�[�/ںQɃ����]��h�6�G�0���v��
�)�\�Q�פF�p��<��T1 ^�SxY���|�d�Z�ք�[8�`�#g�	��虶�P~�"e�(�^���.�0s*�8ǿ�����a1���`ǤF���-.�����;/%e#%��3���_��]D�U�@Z=	ON<���$$$(�����.mn�
��R�`���=,, ��&%?%�,�9�����@��j�g��D(bfÔ��R��bV#6Vlx\E���̭���F]򅨼�}��+�5�G<ǿC�B²�9��s	��jX���D�	������8�(�K^�r֒+I[�eħ�A�̢	kп쥌pP�w��+�Clc}�֟m���:�1a�L� ��D%��l��V
?�m"�����{�ہ�cD���>+��:���/��&����-Яc#2���l1���,��q��<�Z�Z�W�x�`��~2�i!�o�3���TX� �z����ܧ۷o�ݻwtOL�Ƽl�o��׈瘽�U/.��C�:�^+�.ǣݴ`��L���z�����@/]b�{��%:s�4�ϵ�fTbt���0�&��J���'��)�o)�#�ѣ'���S��z-��xx�#R3��3g�b܀�O���Ȕ�b/�f�a���)H�������.&�1���4)VH�H��ϐ��b�b9?8!j��~���E4pa~^~��#j��g��N ��ϟf/�ʱU>� 4G�烮��5�_~�΢0�0o���ZK�qZ��}�u5�L�/�p���x���!���W�����^`�s�V�7Ky��;W�H���2����){f��|���_vl��weƤs��,�Ʈ��~_��`�n3z��
�qa9X��k���\�f0С`�$gϨ�`�E�DҰ�db|�v,����y�ِs!�Z���;R��6�ٳGt坋a���$i_��Rp*yt�o������I=�>3A�8���CË�x0'ct2<��N���M�yI��C{�t��r���j6vT�v�YfHR����Z��]����:�e~�������G���ʠ?�Ba�x��y�7f��{��{���r=|V$	| �H؂7�*b�z�`� �i��B�,^��."��k�g+�P�: (&��=���o��y�͍�x�Y��ו,�pO������!���]D��J�g����\MiO�&*�f67��E3�KP3*�����M�x����~��JӔo�'� t~��=�s�븢rO�R*�c�y�c�dїb	�����C�Ew�<6��Y�D$/#�Zs��T���lo3�<";C�5���07Ϡ��^4�c�#��W}j�ؠ���ј�RxD��T5�E��`�w�c����ke�v��Y�pͤ_�tO�;cƁ����d�����jW�4ϯD�
�ح�o��ﳁ]:���S�^�gҀ���Z�g�+�Ҕ2r�y�	�^d��<�7$@���}H%��N����cF�^W{ӞL����5�,9���gO*�E�`��z�Ȣ�dg̢bR`"�Yè|6���#�)�ͪ*}�yC�"S3�Ȗ I~%�d���]���*��4����!�a8D�9K�up��GC���Y�(����1[IrQ{@K��V��`�����M@J�J��h:f{���;[��쳆� U�mȖ~�X2�x6�&����l�u�F��h�	��^�ɉ��H_�@�0�D�f'>Q�߽�@��� $��}�f�o;��JB�"b0������=�w�|]�.�2V����B��E5yx��4)IEr!J�Z�\�1��h�<6���݁�7��]�	g���$[��gy����<�~���< ��Z 7�;'�8���ޖ�0o��+Z�M�(�R�xE��5q$�I�E�#���s���s����'t��-�ӟ�D�~�-ݻ{�vGC>�F����U_kb:̫��@�h^������Vk�S�1�b}8*$Xc.^8���'N�9����$,�}���]h��5¸���S�b����^��)�(Ì����o�D���l��#Ø�H�C�wss��2K�0�^���t�g�4J�>�oVN�K�r�))�#Q�&gB������ϑ����^�(������q���ƴ��B���̋x�"]�G
�[��|y2-��mo?p���<�M�I��B^���m5���s'��Ψ�"�i�����-:A����8�תB�*��W��F�^N�w��."�����rm8
�����n�5�"�R�P� 7�y��H�2��%�lBJ��p�ˑ�Si1��(,QzI��z��H�*Bmz�i�f��
DK��6��(o6MzY�,^{8�Xr��Q��`d��vo�{ ���p�e�νk�_oy�07Z�L6b��"q�e���s�dR��a~j�wOmy�v)��X^nY�(�2S������@�P�4h��GdU_,,���v���8��R��s�kd��A~x��2-��_�wH�G .�G��Fiȉ�oCˁ�ݗQ��.���*a7~������7nܠ�׿���|CQBr�� �m,��'�ӬZ��&楘SX�sEj�i���MK �1JY��9SL�RT��w���o���%'j�[L)@�!<���x��TÁ�z$enb΂�c��b�-��y�$�^oGL��N1�v��џ�m�7����4Kq���K^IdťW��gĒS��q'�Y&�[��wX���:HўCB8��J��wi���cZ]Y�$5t/�Oɳ��3�}q��=?v��F4�LyѠ�As�Us�E:���@n����#��+���ayϳ���0�)������,R�o���^��Ȼ����fM)�E���M�H��6���y�"@&��9�B���m?m����k��{�]si���s9
Ƶ`���:uL��&����Z���|DY���Rb���$���b�zaŕ�"H,\�0����z�>i�zJ�ui�N=�f}ئ�im�r�^q��=�n/	���""Uq��&�6pZ�L���oȮB�N��<K���tj��M�^���D5��y=��𜉥愗K���(X}#4��d��ܣ��.��L�7+e!�~nx�i��0��+�}�Z�(9�zo�}x��p��m�< ���{t��� v���Ɵ[r+�� a�nJ�J'Q�HgJR{ ���6}^���? ј�l%:�j.d������>u�V���3�.�EגM7x>�
@����o�ӣ��8I�in�0��oJt����y���[��~3�^)�\27k&�6�-HP�"%UT�hl���?d^z��͟�������"��l�����8n]<o���g�_��/^jTNc�N���Q?�ykM�uR|�%@�bZ��u�G��F�l#n��~" pV?��C���ZN;:�3c��~F�-e�0O�{v**e,�7~�Yx+�[0�2�ʽO�G�Nq�i�+��%$�vt>Z,�_/� }s$���a,̑g�o���ya@�F��1{+�k�g�6*����'�^@(U�\���1$9�O��r#pO���L%,�(��Y�s錂�8e���Ļ\7�zo%I����n�ᥢJ�zӃI�S�+��K��A�n��H�S_�E�>����Y�X̀�����$����yR�c BE���5[��\tI���$5� 6��6�Pj:�é��iHY8�6�:�E��uB���lv^�	z�@�>����{f�[���Fe0�m�5��i�� �i�«�d(�}��r3e~��dp�X1���z�y+�_STqI}�#��I����:��P�l�~H2*�#��*��0�

�.^�w��G�N���b*�(Ӱ��(Nd�ܠS'O�9ן��V�7����c�?�x�Y�g.�g��?��S�q�y_%�X�֯3�R�G���*Z<�
v�oŧ��y�^����sC��4M'�Ơ<n*����8[�MN�$8�MI�	�Ք�y�"Gh{�=_S��P���ޱYo��~7k�x��AFAn �������Ȍ�ܨ�px�
(���1����x�w�[fx��t�)X):���G��M�q�\�AkW�^�*�wr΅���x抮��{2�%�HR��*�V�)�R\�2��]�K�c��3��.�(�q�Wo$�71q8N;�m�K�eh/&��O��3�W�8�גtAr�g~��M9��6�̭K�&t��P�Ϥm=�0sM�#����q�����f\���<_�T���)���uK֣�Bv>y\]~������u	슗���h�s$�{d�mW��w�:~y����d�v���Ú���}K�2Ϛ%Xu��^���^ⶇW�(�cQ}��巷� K��1����	�7p��on�����y�y�q�0
vh������.X��2��TA8r4	�qu��	 w��Ԇ�����G�hq������ ���w�@U��d�^�� �l�T�Ltv%G�%���k.�`)�������,�UG���f�I�e�Ԙܥ����h3�kJ���i�!�8U��y`�v�&�7�@�TnBN=ߍ��n�s$�����ت��d�ކ�9��"_�l�y�����6t�����+=o�`;Z{��)��FŎN�`c�gFeNȮ���^�:�k�N^28]���wN�$w�aٱ��Ng�����n����)K��p���B�t�ԫʔ�'����`�7�y��N���;�R�Z����*���dՇ���]����8?�,�R9�\Gi^���T��'��34 �����WM�����{�2~���UJ�i�;N���~[9�-�Ut�IL[��u[�5��������6.��yKK��̘����>�O�0j�Z��#�����4��4�f��hU+0�[����0 #U�i~a��\�LgϞ���W�ﾧ����(-�ja�;������޼y��>y��O���~V�.!!*�j=
�����YU��_��#,#��+�8R>����S-���7�ր�f��-DD��I��Uq��3qw=���1^�R̤� �����زL!D��	�^�$����>��|�i&�A����+�~�2�wB<���}��M���Y"���M�c���v��[�g&]��!�����X�*�;7�ޝ7Ƌ�Y��~�& { ��<=~�n��^�1�y��^�E��a�%��C�e�Z�W��Ϣ�{>y�봵��X5,�]P>��:븃Z��:�}�~�״�Ů�5H����X
��P����3�++��t˞�W��Z���Xq�$Qb�������]��7Z�������7���������hk{��34KF�.x��C��R���w�7������R���V�<q�>��s:}�4\HO�8�ʞ>$��: ��N����[wZ:ą��B.l��$��E�Q�;�������ȴ�]��Ȧ�rT%�SBu�p��gB��7׹���G��;W��+
L������L�+��￧���������#l67��%^�
�c�.��	�����X
bH	O՞�
c�+Y5ʵ(��]��@�si��T6����Hh�2C���=¶ɦc�c���$��Ć�Tu}%i�������sR]�Yb��T�A����e�s''�ٟ=ķ�e���߻����|�v�5}�������|�m�ҫC�kC��Y��>I���2��ca̵�k/y�Ι��Gnd�}�{��t���ޘwt�+>ػ��g��^�3�g��@!~�S�q����V����|�9��{l p��5���PZ@�;כ��|�x�y0��O=w�,m����z��-��Zʘj@q_uu�z��Z)b��58�M7�� @�~�4$�
Y<X���rZ�	���YVG9_�������Q�`�4���=� �����w����Ѓ���
�1��k�_K Υ�^�@��\�Zc�A�ҧ��	��}�G`o����so�i�v�W]�e �ǥ�a�����9$��i�e��(d�1ޢwL�3�M�/���M\ԉ}��a۷��w��w�zZ4
u_|��,�j�����m�`��7q:��]�WX�\�r4�j��[	\4纃�E@����Zޅ,ܿ���{"���C��h�It����{�O�		d��>����w��2�1� "3`���}~�-_p^�D6�PV�++��
�����(��Z,8l=���/C?x��xȢ', ����IKK4���g�B'������o跿�-�x��SP��̙�����&�pW�E�_���A�p�� �������7\M�2�,�����͔�6V���Q	u���E���~�%��9��~Acp����.'�mmoU��>�9L�1��.�Ɨ窕(x3�u}�3��e��JaJ�hM����OԚ��x�6�r��Tf��R����D�������phYD�Q�A.T\K���
y�{.Ȥ���
7�v�����ؖS�L*-��ٗkf9��y^unˏ�8�ĹS�B��f�Ϻ�Jx#u�?I���zZ
��|���{��v >l�/ �:@�|�|p���8���\�����ir�O�t�X�.�Ƅ3�]�=�b�M��i-a� >��ƽ�w��"J������<^^^�r֥,���9{�'¨�f��&�<��(ת��d#�q� a� N�����N%�����+W��kW���� h���W�����ɧ�h>�p|���S��J����J���}��UG�\�b{gH��<g�ck^h�����p�ǈ[�r``��^A���yI�Y���K�B���ʸ��E�^s��3�^x�����bx0�єT���k�)����z-<Rz{�����53R����������i�Rw�ٿY��$�1�-h/ZZe��>[�%�(�|�96yج�8�������������c�K��j������P�D6��ho�3�^ư�w�t��I.������i�n����Ǐ���J�n��l3eЋ���ɈΝ;K׮]�w�}�U���:'�1����ix���hL�>�1��9�/֦i-�q��N%!ʷ�ڒDIhV��m��\�_������
��/Xc��\�w����ǜt�r��$���y�?�i��% �7
}��(�%�(�+����h3���RtkI�<ǽ�3����3��Zǒ�&D_���y��G<yp�V8�H<��ju��Z��i�.��QQ�T��ݚ�7Qu�c8!qʊQ��?
�U�1O�~^{nh{"?���3��cD8ߔ&��j*{)"y���8�)ˌ~�~��^��>�wF���ߚ<�[d���U\�a�ǫ�j_���:�W�4�4 ���lΒ�9�u���i��ƒ%h b�}crI����Jzݧj�N�������螞/u�tU����h�d�KD�
`����@"rc�L��uB��@ `~��5�����܍��~��
\R� q���l������kz��*3��,h :`M�ZZW���g#0�3�,��e-tRd$h��YW��6�H��s��C�o��,3A-��Pr��$��g�?����É�'˿��@"ATT7#�- -j�׸�Z�Ӡ���������
K(�^����mwl���8�2�ϥڜgJ]]8��|Q�����3�����v>��1�hg�S���> ���b<��Ol�U,���$�%E�#�}��jP3��'�p|$�nv3�����|0 M_2~��˵��`���(��8��e繩�������s�g{0��t�fs�eZ	�P���g�ZR�ga���f��Y1+�R�����n�(����ҳ�Y�O=�+QE����
�ňT[V���}�2��>��3Fw�Mޥ����E �2۽K���/��M���g�������dL��h��Z�}m�����}�P����Jă��(�� ����ы/i{{�^�|���vwvT蚮�%~Qh����0�˃*��: �qM��>��f]�ݲk\r�2`�s�#��Wr�4���g� �O���K�"m�N]�z�;�ۥ�򈏭#!o���)��	l���%t��ڴyw��V�;mZ�;���̵H�PB����㓎�j|��3��v�_ы'g��M"D�J��c*���8�i+OжX�b�^�¸ot1�]|DA扰Y���}����cE*�Q�����Ŧ��O���q�_Y����v�u�{�< �paZ� �%~<A��6����֙��Jە�ì�Aoh{ʟ���ڶ>�t��_��A1�����>i��!rK�Id<Ω�@��� �M���HB�咭*?�-ie-P�J�Z����M���=&a�pu�T]f�P�ߛ!���T�.TXٌ�7�a]^Ya����L/����}}�^vmu��?d@�Te�gP��k`�c�q�S�9��r.Ed��A�����Z���B�)�'��!��$u��iĺݥ�~�R�o��P�w��uBG�G��`8���]./̅D��q�8��^4�m��� �\B��i���2ݿ�I+�+�NO�
t��\���|D�*�oe1!�#���0���=�EU���R��~v;,o]~6����P|i�Z��ߦi ��7�m�8A�:�����KB�.T�{eF�cr�4�����\���[�_��j7.��؟Ŏ��!(�h_�
��B`:���ʼ��M~�f���fsgX��`�S
qk�~�ɖ�����t_����rHƉ�,Yn��3���P�0/���m�_�θ��J�]tc^�a��s8o�s��i+
M2�e7���{,Ӽ��%����|���u<s�n�K�q�5� ���fl�u�rȫq��Ff�H=J���9�YC<MD>L����ʚ�Ќ1�� �c�u������cG�].�������v��O���E~���	��kZ�4��s,��h�9E�Q��@IY~��9�H
bR�-���~IȠ5�Օ�Ay����W�۝f��2K��X\��u��=z�� ֬�lL�����u��'�����T�*#�[$s��R���nCm�]��y_U�^U=<!�-3�aa��מ{ۏ�Tّ�vO�ĹX����fI>r#�u��>!�4D�9���$)"c)xQqijl�k���T9DIq��:�8�o�خڢ�V�|��(R�)Ц�c�UgW�`T�����;v�\�����;�����*͓e`�ڂ� |��gaF��U��C5�^�)����<��l43s���_�zM''G�nwܴZm�`�����˗��w(�0<��z���|�(S�,���q$r��^��޸/����ۡ�0��}Y�o�}2��[o���ӛ7�t�@ϟ��JjZõ�y�����/�@���ЬN5\��x���+�������޾ݦ�I����<�����MU"��"��uZx_���Iy�#�v����+� mb,$	��L�4p� �'S�C �}E�,�Tf����޾�o|OFs����y>m��U��}~^+�������M4c^%Ť�c{�X�va�Fcf��^慲>]�%�>`?8�e�1e�ٟp1.Ĺ����0���1�x���ȓ��������������`��~(f�<f���~�����5 4�/������8�wU=�����j� F��v�8��e`�����)�B ���Z-K��iK�\ ֓�	���3�	 ������	8�T��hH�_��Ŵ�o4�,!��-���Į/�6�=�$,�Ig�9�Q���6���������zڧ��#~�9�ˬiM�F��4���u�`�N+gv�P;��L.�1�y�C��{��z�� ��ZSlkTH�Bv��\�_�_H8�e�H�z�Z������|�.��-)�#@�X�c&�[� N�ty��&4�+�l̾�yp�>T����%?'_���E���TwŔ��>?��_�_a{_����b`Ӟ�Гc��bYN��#� И�0�j&����7�@�b;�;�*Y83�M\{d��az���yi����Ŋ��^߉R�x/s�\W�X���7�g`�ԗ��_���>q��)�?\��J�	W�V	�<t[���I�@�-���̎Z�aֺ�u�SN��w�Wݝ�<�ݭqpS��$ �B�փ:@��~.�L2,P.�]2���. ���E�^*׳Ê��{rʲ
��m3�n��ܸ��Y�:d��Y�*����Lh������:����}�������ֶ�4������L�͟��7l�2&451��y׬V�m�n�3��h����g.��%�{殍<c��'�'H�����@B!���ݣ��K�)�0��Ym��`��fE0&��G���������P��Z��cۗ��-�R�l/.�'U�/man,qM�2a�0ٟeq��%�-K��s�ه �]��leA�Z�(�q�JCK�c;�w���|n�d�[��c̨CO6�5r�
�*��"/%�nz�j�$PC��+�eI���L�U�،Uu6Ad�c��)�����"�Hdƶ���z̉�5��FD���}��QtK&�)�bi�Qf��`��Z˖���ޚ���8d`����7haq��vw�ŋ,m���l�:T��se���Y�!`�H����b�ҢY*�BQ<�`� 82�����,�J>���dxM2I���s�D9w�����[x�Uf���
Ü)�
�C@�[Ԉ�So��ao;#�r��`���� ��TV��F����	I�t	v�g\1���ޗsZDe����J������"D�v��E��#*��@�%����!ۙ�"F��܎'�=A��_C��! {0]�y=����-���f˄h&o���%3;oi��M�}���rKe�7uh�BAEJ����-�y��mI%Su���E��s�� �>�	�i�����ր�=�foM�k���*�3�@ Y Wx�����3�I�f���Ƽb�4��
�i�}��\C�R�"y�Od�H��SK&�ʠr1�E����� �A���꺗7*��n| :禋B-ndFC�ƮD6���xL-����þԉ��4�����t�i
����y#�gC2-Ql>;�a�ǬA)�f�>s�^Հ�}��m��{�] �u5�U��C���C�Z(k��?�=���V�����a��Gf����r_�m3�
v�^�{��װ����e��
��u� [
3�FLT
!���� -�BTr�	�n�Q��vz��1����IP��X��j��e��'SyX3s�{6��kl׹��d��M�'u�Lv�D��v*�`C��Ɔ����(��0��/�@:9�=���(�i-(5��<M�?��V��W���k��I:�?2x0[�秓g{�xj�Q��h�`h�/�~H=0����[Ac�+��揰�8�M�'ۮ3������N}�Q5�_������Z���r�2����1��O�`�
J�B[jvA��6��2��)$;��M�B$�QU$d�V&J�[�xI�f��)�-���iќٍ�	���
��%�jaNJ3����"����*D����آ��`B
�]}�|.М��u���ʅ	/�
Q�T��Թ���޸�_�D7?	|�v`�C��,�$�3�b5wLx�f�W3X��?��ƲU���6�������W_}�+r�^|�0�
f�+K�s�(���?���[��Z%,V=d�H!����a�+�b<h�@�y$҄L�p`1曛wiq��qy���Ï�v�2�(�k(�SYP�3e,m����9�P,���𘵺�w6�#��h8v�/��݌U�٭�/y{c}A?dќ��"��BV7�Eࡌ?� ā��u�	�!6�t�-�߻��t���A����e�H�}�O�g`� F�a�p�04�����ϱ7\%�����1[p��}(!���h���y#<�յ@^�}�FÿM�[���� ��0�l���`��l~�J���	�Wm���4�Ak$h�W	7�N)��K]��'�(T5�!�1����RPŴH�
ȼa���?K"L���?�!Hb{{�_��geb�#K�&%�Ϝ�kk瑇��b+#l�Nj�G�P�`(��7y�jUҁ�ه��AJ����ΩZ���tQ�"�'�����:�O��� !@�Ǐ����\�U�8@�&���h�݉gwM��fI�����h�E�]S}��c"̱V+��B=5E�1���=|LO�<�{��|��K��z]>�e��c�׮p���T���9�v����8����m��8�?���'24@��dr��>�������mՈ�ފ�LXU���,7�`a��_��`H|or����M
f�>�]Sc�a�!'����u�X#�.����G�i��6�v��	�u�,��4U-f�zү�ԪH��پΜv���
�1�B9�n��)h���ʙ � ;���l $��5=oX1��e^B��%�'Af��r�jՋ�sG+ؼƃG�������6
���l3fnHar-����Y v�X�0IYLx��Ef35�$�o$<J����D��ư���ӗ1ޕ�;�H��شb�X�}�H)z��(��H�|�ij[ӮcV�ܢ�������U��y.��zMȮك�욺���4+��Ǟ���X���a�����P絲�BO�>����[����̄bۄ���X�}D���ݾuzh��  n�����;e�p��Z��fY�`�-�o&9�6O"��'#~v���/�ӣG���珹� �;�����s	�(Ќ�b����0Į|0��Ij��x�g�������D�&�����}�A�~{�-߉6/����c��TӴ�������22ϸG����55)���OM����4di�6:"+��f�>�n<M-'ls��8hJ��z?t�zC�_���.����d���ݯ��۹��;�֩}���]�o�\޿�4�!��������u����e�	\�sa06/$h蓱�� ���]��E߱�ɾɵ�QeT�4y�=�i�V����4�
�Cˇ�/�"Eb���&	F�ȼgb���Q�ʱ�M{��΋�qd;�]p�8�+�'�I>���4�B�����c������,���j���.Ze����Dh�j4[][�%i��r �X������`�B� F�
�XZ<'������] CO�{��i�K�H4�����a�� K��L]�if�x�>▾����9{��N��+<aķ�n;��C�j�ò�x�.�-�-/�������.	�D����I��NrvYJ���Ӿd��༂�S��y.ޢL���6]�0�E�g���~�J���,lF^[;Š�V�nZ"�/��i��l=~W0�&m�T�&L��?�=�1����ޯ�o�=��y���O޷���ڮתt�Wajg-�ޥ�sM�.?�U�CKC�6Q��B�nx�p�mv�5`k�1��Պ2�3^��Zg�f��Y*��{�!�}z�A�U���%�x�Ƣ�)��w����H��l5H*q��T'D�^���.���2D�*���F�=avg2qiT�L&�P��G��}`�s�m�{�Q�)�r;+�L�'�X�u�2�����Qո�d�Yc�)�^�pBˉ����\E��ٶ�\��!}�f적[�[�r1��!s�۫�;��·���' _�zI[[[Y?dE�sjZRs��x�yk1I�{�U��
��&�Mf��@�j�t�a��0q��=z��-.-:�;�2�o޼a��pP	`@��wN0�8_a3S�1����;���Eק�羺���ܜ�!l��?�-d�<6��i���{(���'��Q���ǜg֧�2_VL`��К�����c_��G��:+Xeɔ!�&IHH8�;��J�\տ?F���X���S���m�~m7Ӯ�����t���ٻ�*���ҼЋ	��i6�<a�{c��E6>3Ќ�-�C�/zf���@��s\�}��&�I�G|���Ef���#_
2�5:Y�<+Z��������(�A��	�ۘ9Ҕ��t�Z;W�^�&=���pYӚ{��u7q�|.�>FXt{b�Se��T]����}<�tF �c��4f �i�܄8���&�a�@8#��0�Q@��E&���2	fv��3%y��Q���g���m�7Ѫ\����wM˥Z�? �镼�ʞ���U�C��d�wf�L�k��*���Р��4�	��yw�S� P,_j�t-��5�F�M���[]La�����j�hG5Iy�bkk+��;��?E9�r�]I��}��7t͑�>oe�!I8uFO!Kܳ��:�: �Y0�2ĹX,���;p�������"+Ř_�WlQ��2��&�9�s�>ڤ�*�ʛ��*)�ӉN�o,�6��D�KZ7/}0۟�L�'���	�{<@�TeX�L�E�zi��FCo	l����=x��q���&ﲬa:=���9����}���������1���g�#!`����<���G�k1� 5,	l-�-��U�<[D��c���9#<��q��3��48�=�p�5ͨ%��NgY���d��JX-�, 31�,L.4�PW���W�Q��X5���dE�@���≜ք���F�Mz���[D������9�;�
�74��M5>8�۲�["xѪa�]�����3I���$0B�2p����}���#.'JƜG�y1\�@�$�Kf��c<u�+�?:��;����dE��'�Y�nQ�	k�g�d�F�}Mn�0�k:�U~�{��۷\f���J r��Ʉ��V��T<��"�#�x~�� �aY�D� A�#��ˑ����68��lQ���B0�{�{X����z����B�}X:�����㥚r����j��$�2��8d���M���JOk���.���� �+Ͳ!�X%{���d�Ԅs�FE"��c-��h!r��b�_\we���s���
�()�&A����d,�����"h��I���RfTZT��������-:�x�_�/�͚7�����w���`������eƷ
 ��G�SR޾L���׬�E����,�
��<uʭ&�+R�f�L+<q�iiH�"��Wk��r��xq��1Z������@��7��ݶ��4�0Gmr;s��p�&�؁^qcJ��		��(e54 �&@'�JePd.Ff�K`�1�QJ���@�سŭ"h�$칛�F������� �`yv��03�)�ͻ���N���[�8�?�X���}�&'��B��yB0��yQ���7�{�ط���d E�7����?2�
)���Ύv���C�o���mx�*�C�3 �Du�e@��ht�W�8.P ` ݦ.~�����	����d,�H
u�Wjiu`	\�>
��>m���%��1�,��0����QQ)Rm��V�kF�쪘�>3���G�$gl����f���);�K��е(��c�S0�=d��g�1��Nd��pr��`��<R/W�Ï�fI���,�=��k��v��,`yނ�Ϯ��P�P�Y<WZ��m�;��^��LE)?URr�\ӒE�և��s[ej���d�30�j���s�bD��0�;fR ^�*`�tZ4�n9����-j��m:��� �����	#�0\��b�sþ̶fnb!E�$g�6�L2��'"-����$1�X��"DA��[-0Y-�,5��i� n�7r@`���������\��Y1�����-8���LB��-��̭Q&7�sn�i��������h�]Kf������\����J���붐��D����駟��Ćq@.���b�)���\�9�EE�!��>li	��C(�R�^V�̖\��$YzM��i<�4;ݓ.�	�D!�����E�ξ��Kt�Zḿl��v:st�T#��O�)ި��1/̅]���%%ע���| I�Gcz˅(`����d�.[ѡ�Wk�c�E"�/;�h�%���Ū�f�Y�12�A_�U���|�;�_�-��]��=�r�W������l!���g��,CmÇlUR���_���8��	=Vb��8?��Z��y,��F[NH+F�;(L�U�͘bv��$����u�?s���F/�5i}}�6֖icc�e�F�1oO�P��K�f6����򄤮4?kiffx��"=�2K3f��Rv���� �Y�n9ϵ�*tx(�IR���i��5��0��:I�&�!�tig�����h;�ɱ�,�p;f��s��ȇ�Z=*������;,�L�N�L(L?|���L_��NC_e��\-�fύe0�k%C@lLb�>�c����p,�`C�vc.9�������z��}�~ؾ u ��E"���>��d�(�!ˋ�W���L,�D�N2 ��7�Y�s�a�0�ۜma��Hd(e���̩(w��N��Lc�����WV�is�k������d }��>`,d�kϬ|�1(��S��H���|2����M߷,���e�'�i���"��h�~�}?�H�1�`�*��(�Z���3�L�L��	?V��J�ݯ��ZȞ�Z�\�e���E�8���o���hW���˦>1ⴈ�9���ř�ՠ�m�X[��w��V|V�ȥ2p�:;�/U��0XX�)H�YLC���F+�t>K�s��Ԧ�9Z_��N��n����H��`&̲2��i�3�n� �Tݨc�sd^�^��.�/Q�����n�N�����I�%	�QB�N��l�̓�D&�Zp��k:3��� 8�;�9Z\h�ڏO����)������;��םC���s<z|Sz��1�\�����V��J;���� Y52c֤Ѐ���`-�nY���MW��~��X��u2c/ϛ�RK7���|���-��ҏ�w�>HV���:eqa�"+)��,/��	�68}�ŸaA�iw���M�̱�~���/rq�1���U�p����w�:\R7��"!�!|id�?����E1O?Wr���j�=��OO^! �@4g#�@�ǚ�S��f-q�%�>�qf�3}�J)��2  W�܍�Z����,hp?0C#���.��_N��<V�mU��e�y�/S"Aʬ�elR8� 6�\��ˢ�Z�0��\���kY��$��؋h�M�N��F�E#��������>Q�/o�P�7�c>�_���\�%�0� ���eq�E�K���H+�.9л��fC
6u4��9��y&yx��Ғ�[S�~�Yy�l��l�]�����u�랛���͉h�=z����l��Ѷ����4��H�>�W�U�I&����93� ��z��6��-��=s����w:�z+�ݽ.�Ni8��(d���״7��s��S)J��O��v�
�7xh�]����k�q+�,>�7eT������n�@U�Y���&�;���+�j�+��©ߠ�vߟߦ���ɭ��xZjȎ�^�����gI��t,,��?M��ϔ,�K�'�O$3D�sھ��<$Ԉ����r	c��cXp׊����i�Fw�R�����+�L�(�|��1��Jؽ��?OX�f�������,H�Ʝ�mh���{�K �H,��� 8���g+Fd>ĩ��|�;�	���޴�+�qr	��;�sgܡdj��������#��/?�`��O��_���9�̲ ��:��T1�!3|���=��JZa��:�E}�u������UsR�ڙB^!X#�rɻ��}&�����sW��%m�8��Seg�G�Ƚ�T#���/@s����Bd���+�a"�c���#��Z̈́���h��2}�`�6�,9�;�爠���$�BN�3�g~����$Ӄ01�q.�D&=��uZ\Z��G���ң�Oiym���6�Lx�������￣���t����'4lOh����#�g����1�� hKz���l	d�:=��Dw�,ғ���͛Cz�|ǁ�=z�v�z����d�����#-I�##����ʜJ�� R1���w�}q�����wa���n�}nӸ- g��hV��2X�.�he{�U�,C1�'�X��ʹ�\r���%$m,0�J�]�F�Ά
�J�d� ��i�5���{ g��	]j��랱壌A $�\��S�w�,1����Dr����`�37�ZZ�v%��-*����q�g+~���ghj��<Y|ODb��8�Ye,�U#Zr��&�b��hi��T�Hk���r_���<�I�u�Y6�5T��f^�P� r��>DJ8O_D��-\��g��-B,�Bn��Pc���$E�x�ƚy!p��=��S���<�Pٙ�'4����J�%}[R���?ۇW`��i�/�yY�e�S�e9�e���[�g�dL��}qi|B�Y����V�+���.�&1��Z�GgK��6U��y���<Oٿ˅�.n:p�`�R�~#��B"8I�s��"%
��U&6;�����f����T�o� ֜��y��%Y��@�P��gt�I�V��hՁۍ�yx�k�ڝ&�o�gZ�	e�-/S���9�sȩ\=MR��<�ԡ���cm~N~���7t��ԙ�g �f	nY79�-,9�b����y��	fn�/O��d�(�n �Y$A&�����o\��;����m��s��rc1��2��"��F=�$�5w��'�s��n���xF>)�S`�d��S�^�75���*�#�w�g�Х���p��ʆ� �ӓQ�P��I?�����-�s)��f}c�<�GO�|�yo_<{�������lg����ޟw6!�g�_�ā��[��W���[�@dl�\���a�/���i����G��������?r�4�k|�٬=�+foIr.�(l"	P6-&�1�g�i ]M���jl�0��'�HV�Q�Z�rS�Dl���p���׶y�@�����E(2c�����99�W��f�?d=(���J���̆m������C?=!8o�y�}L�5zB��/��S�f�2KkeG[T��g;��*b���U�X�<���{�������6��{~�cX��������eo�I+R/���#��)%P�,a�0Y���Jb�\�q�&� �	�˹�?� �Q�'#괚4?ߡ���=����wP-��~�NOO�X���*�;�a�ra'P��$�a\s�M��-.ޡ���}��?���C�_\����	9p�ݠ����eJE<#�D�(3MY'�ZA���&c-Q�(>�Aj.����!�]o���}v�=~4�������3���[zv����h�@����3����3z�3%��]����4�6I˧�_�]����>��+��u&[o��������a_gϳ�0 [>c������?��������D����w�tt�E��H�V�ѣǴ0�@����i:��:oi	�T�p�sp8��G�߱,����vqa~���ۤ�/�}��o�����txx@���%`}�O�ץf��v��2�ʋ1� F0? ~`�-UY0�l;����5d���E7jT~kxض7�����!0��Y�4�R�f��ceA{v݅��xD&�z�@-�iY�A��L7rc񲴴Bk���7����m=��vo���t�sa��s�Z�����>�VffY������ٵ�h��#!М��f��jW%SΓ\��8���v��qޜR����� ƚ5�)��ؐ$��5%"0h5+a�]8���2� Q��hw�:9��&"�P��BW䮭�� #��VO�t�����Ʋyk��]^FV�!���D0t} ����в�y!Zf���"��-���Y���l��i��ە�v7hiy�MJ����,�e8�I
2�	}��1l���k�������pǑ��c�~@Ruu�D�G<��EiC�ƌ/)�����,���Kڼ�J�k��zk�޾�������.1[��6Y�a�#ո��pl��(��Et���<��y7�/���,��Y?oz������6��w�O�,pUɳl&��ͻ��c��;tgs�͘~����������-r@h�'�N'q�{�NNv����kHͶ[؍�э��ȄXkϚ���P�#�
�D0r��}�c���rlC�`��ŋgؐ��g��V�졥E#2�S����Vr��9��?L|����;�i���(�@lܬ���?X�Z��q�{���� ��c.��._��ٿMj!�$Պg,A�9v!����mq�\ r^x�x�c��3&9`oF�۰z3�E�=�ml���;�1���Wγg�#����~)n���~��.~���et1)C�hE+gB�V~V�����`|��nj�60_f��;�E���{�"s!+�3�av8��}Ga��j�rU��*3�7p��[�>�0��4_�2pE&�KH���P��Ԭ--���g+������c��i�&'qKF��,^�Qӑ�;���`"�Buq؞��q�:�������+� ϻ	�n�_Bcf�S�N��m�ڴq�.ݽ{�޼�C{���Fr�d�B4�d�0$�LQ4B�/̀,*�h�;7L������_���t��czpo��S�ۿ��գno�ޡ� $��0���5/Yqۜe{C�B���"�F��r�ؿ?�x��^���@��M���y�9U*���/����=����	�ywSN�N��W�s �K��h��:v��3_���xr�T'<p�����-|H���I�$��u�4o$�"Q�����gZ�F�)�����县�{�}�����yc8WK��+ƳP�9M�XZ�@��iC�fi� n���Y�`�7҅5��p4:��l��T�aa1
;&r	����kj-��i�:�%abO�h5K�g%�M�,~�%�!�R�`�~i�<���c.�� )�YK�b_�����\4r3C��b)�7���E�-/&.��vا�p�`4J���si���� Q�脀�����V���e~6oUY�6�x�ڧ����}����0ѬtM�S&g(���:e������l�R)L)��tk���Ո�۠�W��MN9��n��;��p�%|fVY��e�΋������+���Ӈ幝���Ւ�5$��X����rGp��	g[��"}���i<<���K�iu��D&j4P "�B���'�(��i|ܫwr@�1���$ڡo�y�@���\������K�V����;J�G*�Șa�3���y�B��V5!�R'�� תI�][a-�l5�T��2&�s�:��u�ĸ��3Z�~���*"WA����K	�����k��?P����E�ww�6��iaa��+����'���g6xb�\����s#�xYt�>U5�-@1����������@׀m���&�� 9x���7�I����@U�� �r�g�8<<� �12�
w���
����?�L�ȗL6-����MKm�`a�ܐ������W��F�q�-=��/���N�L����t"1r�et4�Y�I�-btpp��z�/���1���s�;�9}f�&o����_ۅ �J���v�Ì!�k��CɬQ�!a�|�ߕ��M��Es�M��z���
^�B�Ś�޺ZRH��a�zk5����!��[��� v����dF�'?,�E
v3܈�t�+s�����	�"��n��q�[L|БE�X���@q��\Je��k��}��gKYanW�ٵX������)�:RF�����K����t@o���&���)��JE®_\�\:a35f%��)�1-//��ߡ���#�o����=h<�MI6��6]\��'Xz/_}����\d�~ɓC���߼�C�2�����ʌ��������;4���᫚���������ZZ��g���{�������zI�^�L��ߧ��G�����/��ں{����^�~����r,��s�i�\�P�WM��2����f�힛5�w�������1�z��0�Xu�k#'.���"{���e/��k�C.���+P�;&: �n�ˀ��E�8|��V*�Z��R�lL�0��٢0����R5y��h:)�����@
���3{�i	�s,lu˽Qgb��唻�S�c���?8�}wOp�����w5����͏��E`8��&��h�e�>o^ت4�6��YӰ���4,Dd�eكf��0�Bq����M��Y��蚝w]/ӿ�m�7}-b#>��PD�ۋL�I.
.*IJ�TJ�e�~7+t�!�tr�$�����bިs�4H2j7Rz����7��Ǜ�8�p���h��2�C��Z=�	��$&�,�-�`��@��,���\�0��D݈������Iw���{<�I=w�&��
s��gܸC7i�B[4?ס^�E����=���Y27��_���6�D�cl=�З���簇��#������
=}=䷜������^�|K{�]�tb��9I��!�4+O�A.S[��>��^߫��n���D+W�����}�˞�E�rM���di�_������v���S��)u���X\\���yֲ���H�3a.���9N�(�� �����W_=�o��[vmw����O��-�م�y��>W[_[�~����K�؃�g��=(�`�O87,yЫI�|�
��p0���Ve���z�V����.���Ջ7���+��;t���;F��V�<<,M��l]��sI�G���� ��B#XP��qttD= ���^�xC� �MN=���+L��~��!��g��ݗ�
K�u\�A����D�K��QV/f�x�ȧ�D����cI�TtXĠ�� ��IN}����ߧ��c�����pҋ+��䪬z>T��|4-)�o����]���V��������DA�����&�	�}�=/�=�3�K\��
��*���he9ެ��ͳ$���M�5�"�)�M��)ۙ�z�F���c���7o���O�z3>ʨ�1�5����H
I$�.��F��6	-�,��;���&=�l�:-��S��Wމ4�Q�w�_��6�:Ògu����,R�O�,�� �����6��������M[������_XaD�é�x2q�8���~G�+8�j�h�=�͜���E�'e
��+�7] �D\��PY�5|��\�p���FL���{ȋ�Ng�����@���Q�l$�"t�(�X�y���X�\�ͺ�?%�g�*�D�C\x�W�7��:�{�a+39M�eM�f9�͘(g���nӛ�� ��	��~��7�������������%����yN6�^ ������=�k�nu�@K%��x�N (���Wb� b?���$�~�g¬�c�@1<�(f;��8������m7����߻{����JF�%`6!`a�|"Q�����r��7�N�tx �|o0 L��fK� ��)n�E�"�dN�3U����bSc�r=�����p��*��I��bC�2E��p�58�y��[d�x��8���Ԥ��;齇�s��[D���@�+��܇7�f�k�ye�ۗ	������B&?�Qk��lb�!�~��
rv��d��0�Y�kc���ӽs����S�bK��M��`_���1�DMbI[��*��ϸO��8 /����i����nDԙ�Ӄ�K�������[a����[�wE����j7u�_c��ZT�0n��6rR�46���/I�].�7]�*G��m7�b�H����k��}�m���T��z:���Ұ�^Gn'��1�IR��As�3y�b�(xeU�O�� ���{n���� X��trt���{�ѓ�7��n�ћ7oiw��&�>-�w80�+1sRQ2�n:���?~mA+k��Zh�B�����d)��+�=�I.���x;���h�ת��`���9�3;7IE�a>�]�����=�������������g4�9U����F����؁�#����t��FA�n����Cj��΂@V+2Cy x#[�K��8�E.�E�N�,�jwȮ5�ۭV�M�9���-,.0ù����#��A.!nK��=�ɵ��y3�>3=p w hWy0�
����D�!d4���$�:fa�����u>�Y)/�����챋"�`;�"��U���+�Y�L�x�ƚ"�Ȫ��}A�HP�v���2�/^���� b�3W���)�Q�Q�K�y�Z���kl�<�����++[��we����j�̠���ؔ�L�d�5�nzU�9�m<�;c�m<�ʉ�>���>�u��`�5I�x+�Q��UZЧ*�N�WYqc
㫃�}�z��Q��D�n��W�/ �%7�<�b��<�C�"�m��	�*!]��;��Ӿ��]��O��҆>��m-*Y�
�X|�^.z����bQ�{r2f��i�:�%z�p��������)�V�6Y�/�'}:�{C�ޮ��xO);�>v�b>�Jq�s߱�1"Y���Fr*@�_��	O�LŏQ�k�@ �u�՗d����S�!�(m����.�/�n_��~�����A������O?��J`I�$�]��_��
��t��S� �s�>�\�!�0�7����W��p�lS]��@���.�OU0[1����}$�Zuq�`g��@kkwhs�>�j������^�����+4��J��-�#X_Iە�2$I�_BR@E���r��@v#�F3�g�w�w�r�������>��N�-��������r�tqv>���`y��y��I`���R�f��]�A� �R��.R'T��k�B�L'd��TJ'f�߸o�( .r�q��X�L���n4�.�y���=��t3&}���e���vۍ�{aQ�����߅\\�K�+t|$�^s.y�N暈V�Z����ȟ�M���>��������!L=f`��^^�@�6�\�$���'�1K��e���>T����[þ���J���/0�=����+w��j�]_����gW�i������%0�ĩ���m�w���\��s�>\���u{�t��To�:�Ap�K�4���3��e�H� ���U��y�ҋX�����"ǣ�Q������n���%v�lыg-�S��p�"35�����7�;C�&�I�M�',q �d�8zp�S r��#��������r�w�t��o��t�-�\�N�c�fdD�x��23&�A�����:��+���>�v���fyI��n�̈|j���z<TVQ��Sbp�ELBW��<�rJ�Ԗ��M��TQ�6O�ʺwoxЕ(����i����n�R�\> h�ڭy�Ya\�Rw��k,�!~N'�䑗6�ł��Ғ�0����N�N�s��@�p8b �>�K�Qg��>��|��=�@�ga�	�h�,�Y^�D�V:+
BL||�dq�ױ���f���Oζa�n�/�#��F*����_v�m�Ŀ�T=��E ��'n��֊�O4":	l[���� Wd2]W��7�{2�`�p- �9��Ki�Z�ʍ�\g�kLܑJ�B�@�b��r��%%U��YvmS9�{�-�ݡ���~�*��-���=ku�Y�0�x:+ˇi�[|s-��,2����l�3{N���&+�{)ح�db��:�H��"��kw!ch8��p`�ъ�ɓ��7_ߣ���N�����H)1�pձ�  έ���z�fk�5�h��z�c~G�j6�dU�5G���xN�%�HrS:��M�gb� �2�4� ��B��x�A{�o�_w�����<Gn���j��j 7Y�px���}�cT�7h|�͑��69��G�G�}�_��q ������E������νU�@-.�r`�?��W�n�����E/��%��n�7�������ݾ��t� G1����a;���@��eLB=���~�$�
PGm"�g>�����'bͯ�rs�x!0	yV��矞џ��=�l��#�Lre<3�ڷ�8�^e�Ɔ
HEƐiڼX�G,!�-�\j`�r�����U�	��i[XX`�����#b����Qʹ��Ѳ�S���q2�(z=ͽ+yw��Z�Yc�9�4N���%>� /��'��F]�l���F�yfr,k	����d �ɓm����y�I�T���k�&}Ev�5�5�w�L=���yq!6��@��:�����>a	֫W���:���0v��ڧ�[� ޛn�g!lU��C@ދe�mie�kϯ��3����<g����mҰ�م}�Ũ'��ھ~m�B~j�"��x�,'M�(ۄ`����"	E ��0�$Fߦfv#TN����D��&w7���t�����ѣ5���s�6ty\~����l.�=� ��L˫��� ���� �����^�@�D�*S�{ ���������TO�@/t�C0�'��'f��	3��.&���2L�T�n�<9�3�><��-��\�X]��M2OD���n����?�C7Qd1�Vhq~�#�1Qc���v�ȁ�ɤOGG#���h6t P��>��\r�"v�tDXO�y�Ǥ�i-� ��X'�c�o���}�B�&�hͯ��nz��࿯V�SX?F@�1P1 l��Ҕq�.u�Opp�m{�b-siJ�����1m9@��?ҏ?�LϞ��TT�>�ڬ�u��TR�1ӘJ_� ��M��x)��b#�-�Bvf��r�ο��-��; 9f����	��nk�Тz��{���q��Y$�$�������7�Q����`���a�3� k�y�z��7�l50�s-�O)X1ͺ�5���R6��ܗi��Oq�LL!E!b�� ��z�Ǫ�m�����1�ǫ(F��4�944�����ZD�w���X�x0q����'�������E�e���"�捵Fg��U�+U�{(�������@]�l�Ԙ�P�e����o��zw�L9a���e����������=�{yU^�pA�NLG�q�{��r��V�I 	��X�YĮs	\��ş[t���31�s�ʀ�?&�V+�͍z��z�p���ۜc�-�&��b�l9��L���ރ��������d�J��������?�+�x�':��y!��|����c���?N�|��f�w�Y*!��ā�Z������D����f֮1����r��^��^��nI	�T'&0����'�łK���v@�4��m#���?v�؜�/}MO��-}��o�$���������O���^����v���ā�V�V�(�d���U���2��?~�ο��!�zn�7\�������Fe��XE�2��y�>��!��,�c�._zCh���-^h 9�<k��q]�t���41�)�8s��"E����o�!�T7�2 	����>W=���!���gf�����@o�lsA	�C�ђTb�TݚL,*9ㅥ�^)2��;�8 8_�i�k��H�o��B\<"�v���x��9'x-��¤ƀ}A���!_/ȋ0n������?��ޤ�<,���2^��^��χ���
�?2��EVRw�B!0�H���t9��wzZ\S�h�3�,KH"�a �'�}�\l�-�������i�sφ��I��e��:)g*��i�b��.쾋%��2��"���2c��s`���`�A'��`4�H��{����r��m�{�BPS�g_����Β �[UZE�?��K��c��#d��^��� ���e�F�i��[cv-���]��(�G�c\�^g�g'\\���$�s^�M%���L|��+!��ަDV�v��dŞq45�d�@C��XT"�$h��H�ݝ�4h}�M_|~���Z؄#���Lv�1s�o�M�봲�m�����>���*�;����a	�X�A"!~�����Fa��-���EJ��i�8cdؘG���bY�g� � �B(�`E��������)TV0p��I�W(y�l$��$J�BcLR�ؼO�k��o��|���gn?5��V��nѰA���������&�}����o�:2:�9��x��	��>��~~�	;T#)��k�<����$W}��Fǌ�=�2`�N���A .C�����c%n�]n`a�����[ZZ���yv��}t��~FQ���E���磌�K=8�� p�N�B����Fb�H2 �Z�
�?y*1�����C�QDU��E��[�ctb��_n����sH��J3��=�W8�Uf��dT��������	{����,p�󶭖�An쒱5�����v�5���� ��KX���[������h�%#C�6P�Qg uK$���pO�V8C&��e����*�I8���L��.�0������]4Y�6p�1�u����@����9v�~f�fW�����8��̦zңb��?��pD�^,4�n���'ie��Ҍp���iЩ��=���YJ����^Ό4��&�]TQk��{������o���6��'� eW�K�:�[˴�z�<��l|NK�@�rNȨrB�v���۾�ѿ�������h�]��\ �D�ZĶ4ha���U �����>Wwc�MK΃�a=�p�y85�	����Ut�� Re�<j���A�1�``�����O^��>�/��-������q�oz�>^"7Nw��g_P˝��������Z���[9.�8�.�;�ݱ>�c��޼�%�Dp��.��Q��j�>~3�X���� �5�gyy٧���d����Z?��t?0�&Q0�- 4�>���7>87�l��[�����X�И<$��z$����� 'S*h.���j��4%u�����XF�\���Dɳ)���B�r�Y�`�5�(��`��/49/]�:�N���x�1���g����M��i�G;;;~�m���I;S���f��=��Nj�0N'��L�[�/SQI�Az"1�6�j�� ���X���f��^Sa��)"f� �,	|J�^���\��]d�j���kΌ�ĮU��o��M���6_������"�̘{N���z���=E
��'얳;\6F��&M��_�[V�&���C�U��U7#�j��1v�����DR�����4�8׎�ia.��w��/���J�M����O"�ǋcwS���]X\���2��6@�����{-�$�O��@�˛>r�Fy�=�G~�F��*A_��>)�K��M��y�F,�@�����X�	O����Xy�c����\��b�I&f�"?n��xV�l���1o5;��BBq��z��K��,�������;���b���ν�����������.P�	:]���@�M<q�������g��{@�{'ttأ�)��%�V\#ՅL��y���O��ga0�`$!0Ё����{_�7�f'�ʁ[ !-ئ�;�7�2`��c�Ģ(�:��� ��-y���{��>�37�{z�i��,WY�T��ȧcMo�LSI�%YF��e��V>��2�2�݊�~2���e��f+�"�	���
8�Lь�[�dE�ő> 3���"��W������>}J���c/�����x�a��� ��p�޴E���v�<$�m\ʨQ�	e1��3Y:�{++oldj�zY^v�0�LO,W��׺F�G�X`����E?���:py�e�0]m���K�>��x�j���z�lc��w�+@�C����y����{,Q�GX���N��!��i�]�h��SC�={eY�l�ه���nK��8�f���&���(%�%�D�z��k�l�<�%n4�@$�6Ñ �V�N�Mj7Sx�6�Z�-�g֨�N�{� �i%l,�,�j-�7��M1��"��z�����4N��djs7������o����|A\�8��ϭʼ#"�i�Hz��h8�d���_H����Yb`�;�Զ
@����r���M����1Wl��\��.�^�y>%���DZ��$�;
�F���}}�>��?p�i��*����X&s0�fBK+����#z����4H=z�;�!���G]Z\B��������l�F��Ao�1�l�w!����!��a���:`sV�ʔ�h��>>��������P��~���t�^D ���|��j`��w�:O���wl�l;;u8Xms�`kM$�x"�ITYKk��Ȏ����DrQ���r)F�e��>����fϑy-p4�h�sq��+��d\0-\�<��.��3M~�����FBƅ�1񭮮җ_~I_}�%�u��Z���5�O�A�<VmG�O�<��񷠶"��p�J�r��{� �T�9˼�`K+F��-���/A�����h�_�}������|L	X+��`Q�18'yfL:��-����Y���Z�Kme9Z9�nXYr�+���,"�ƀV��[ւ���>=��V���d6���r�1��y�%��Њc����k��HLq=�f�M<���!s��������O-z��Y��w�iq��6X�#Қ\�^�Tb��͎{�q50���E�Ƃ\��T.�����C�E�F--C�� �	Z��m�Cd�-c4b�~0L]��nB>�㣞�.� )6�Ԩu$�)���:��4 �?s�P�#S�E!�[���q}�g��D�����0&p�pLp�����r�� .��8?�'+��'�&-.,1x�n��Θ�����9��%�G=�y�<X����[��9�W�_#���@�F��V�R�2�wٗ����[6p�Y������2�Ӌ ) !�����{g�����YGv�H��8�_�/����ϩ�P>�L�=/�@p�����z�� .���f��_m�]R��W�Kz��`5��(�#�g�n�x�k,a��ӑ�585�0�k��0H�!����3�tQ���$m�L�&3 �<88�T\,s@���[l����o �4*�黀�B�&��4�(��-UZ�$��ll>���#������˿1�ݲ�`�^\���,
�yKXl�s_>{�����;�������g�`:Yht��|�� ��8��n��9�N@O�s�+f3�����{�b3B�&�oϧeO=$e�z�B�}ٮ�k�nĞ��T5k��������c�ˬzjc�HD���ȩ�d!�|�A�S��M-I
M����[^k�#�?�y�BE5��[1-/����%Z[�sۏ���]WR8"ɏ�	���3E�U0���,N\\�|�䒺i�`$��hee���q:ԉ0�<��@�d	`�0�X��nĤC+�������&��uo��8`$��J�Y�b��0yc����������)��G�Wo�X��ָ�;�����+p�
�5�\s�<�$Y$Dl�w$�jS������
��n2R��9��Ȉ�C^d`���{��Ɇ���q���()�y����=|�1(���,�a�#���C���5�
����[^(���_�;�Bgi�$�I�:^Qt�@O��K��1��,o��}�i�t��S���S���\�k(���(\1�����悶���>M��E4<"�A�DS�':b�9����|�%�:� �����u�� ��Q�Y��¹ksR�M���≴��o���_��_ .����d#ͳk��$��1���v *�-c���h6[��1��ت0q�
%o�{bg$�\��]E"QP|����TSə�+�󭫎]��ٚ]z��5�}�H�$���6�`~�Ƣ����b�H`]oDa,��[���$o���_�����<����g���GH|��JVtVnUR�*f7,	���/�>��k�[f�Pa�r�*���z/"���ev��[�"�/���K�&�-�n��4����YN�îŌ%l0T�$H�CHaBX�Q{�Mw֥���bہ�.̩�M��+��0��h�����u ���X��c��2R�B:��S��8πw�l}�<�2 ������>;;ttr� �6�ܣ;�wicY���򺛄�ky�Ͷ�Eu@�ݘXM5�g�����z���|�3=���Y����f쎳B���4�i�~��5�"A�)d������I��E�i�Kq.a:�F���ǣ��6\�+��=�w@AԊ<�E�<p��hݝ�Ç��7_�a$��e�֘�e|�v�2��"��^g�~c�%��t��.�v�5�(禍�1{p�����}��}�����>_|No޼a@V
��B����I!�?�S{�>����ۤ��U�_�s�-i�q�}�����u�!n� �~��Fa
<�D`�e��	e�|pȹ8E�e�X/�-�9>��'R ^�A��0A� ��H*"X�)8-[C�������U;����[�ܹ?y�3 p:�L�ܟ~��~��/�^��5��,]`�HQ�N*������yb�~��#�������ݯ&%��k��g��d Z����U��Rē��*��mk*;�d�)Ǡc6�:X\vc�c�&3 ��_�����su���@:�@9��h�άz���] z��s�f�����3�#��e��y���5����۽y^����������dE���������I��2O�i�����lm8_\FFp��?o���Z^���MUM)�׈�I	���@��$��h<�����8�ZY�bkLf-"�Zԍ���I")�VX�o���())�$j.�\�%>y��5FTKG��En:��헴�Ǵ�ޑ���.���ˤ�,��������e�	I�� �&@���!�[�y����I��8`�� �]t�Pg~Ł� =��d2%بK��zӁ�9o�2����O��o�EQ����@���Kw>o�wB�'�nR���B�jGR���C�t���:`zĬ����z�Ǻ�/�oN�6p`�x�N�v8R-	�	�T�Jtu� 6��܃��u��ۧ�z����sDz]]�XxD���hQtv�0�}f�wg&��q���6�<^�|ɠAk�1 ��y�% $s�X6��ߐ��#6"֬��YfHP�z�-�d�r�B�`znA����F�� �7�²f�t�f���g�\SJ�]I7��qL�GC_��������o��!� <O&͐�fP!�O^�/�4f@�ii�H����D��A� ��f���2P$���!̶�c�s̠�����[��ĤV���S������ր��+��i-VY+�㡀t��咁����2�5�ÿR�5F�&�<x�g��.���&x۟�7э�]��� ��g3�YU���*ݕ�d���Z˞`zݲ��R2�v�졁b�1�L��,��Ee�o��1���v�4���Or�Y�L��w8�Z��`��P�KĀ�S�!x��v+q�V��l���"��*U� �3'd�\J=�L��4f��q��emL�Xbq:!IF/w<�q3��۩�H
��c�E������҉��zt|<`����
���1=��)}��+Zrǘ_X�(i2��k��k Ϝ?t���|�K��s�"�(
?�������?��?�矾������r�)�$�L�9-�4���́�vX��Z�s�b��b����A�N���`�M��n]��~�Q���MѮ�E�w�����}��C���z�'tptත��:2#�}����b�35����m�a��E�<�D��]__��?�0���PF��i0'�iia�����u�j���-��1�'�E��ф��օ����\xa��2��2�C��������Joi�pЃ��g����[Ե�'C-<����~tt,�s�*�h�\x��a�%~�l监����<�җ��Yg�0.��N�Hv��y��8q��d�(�w�m�p5�oY�!Y9�J0$U^1��s�G^#����������6L�G�\w�rʋ�{��Ζ�-��µk��Y�n���n�l�yU��/�ޭ�:�D�ڋ�˟L$�O���>]���\k̂�j����w�iC�EX��l�^�3�/]oz��c��2��*�Y~�3�sፋ�U|V��m�ߒ��f6"�8A���тp��-ҺS��G�B��t���6-D�t���!��5c�g��[ԙ�w�p���4�����=�g���!M�t�����n�K����ۧnwB;{���,��'��-�Ս��;�Ef4#�ť���C>-��2�<7�/���>痚To-���}�����^>����������f��������<-��1W�����uZ^[��o����x\�Gwyy�A/&�V�y��^���Mrn�����w�G��v�2@!��&�ûI�tp��[�,-t����pD��G$���s��ژȳ���q��<��c6^s{C� �}e(_�=4cx�cR$��l����i�P�������G^���X�ј�Zb��`�"�<�XC���.�6G��;���G<?*�R�V�>�4�/����r��5�h@����R
�8�;\I .���0�"��ӂ�ˆ�C̲L�p{�C�K���l33LZ�4�i,�j�9s�|����#4�ss"�hjU(wnsK+g��J4,��Y�Z��3���L�ad� H/$/
P���:���U�keLKZd+�&�(���i�%�	�C�J�v����)
�K����-a�:v�4�"[k ���4<�%j�`C���gh}��Zm�N���Jw|����c3�UǮ1���ެXL�d�<�ك���̻����b�`�k<!��Z\j����n���
_n�dB�,�yk��rq0���5�p���s��}z��]������Rf8{ΐ�؍?�����y�%8��_�1X��vw��ã�_ї_��{��KθC�x��M�$�f�gJ��8���Q^ǹ�� �Y�r�}q�������&��W�����@�~������!_���.K/�76���2�[''��ɞ+��-΋���M{o���hy�=�+m�h9=�2�8%N��ã� �>n�ưO��<=~t�޼9�~H�D�i��;�`¯���x�ە>V�(SM }�? �q�_� ���A�,�"�D6�N�� �n>Ɇ������Ip���[!0�'<� 7�P`d�9��$ה�[����=��1�Xk^�j9Lr��SkKD��gk#E`�]��a#I�����z�J.,#���@�xQZe�HmE��7�)rx$���ʭNn��	r+F\c��:���L/1i����7��Ȳ�{��$ARԾ��KWu���=ݟz��|�3�g�j��tWeuVU�2S%q'v ����c�>{� d�)�tB ����]�����n������w�$��ͻ��<�q<ϐ� Q�!UQ0�h6X�����̃���D�3�zm�����C&<B�@�}%�TA�-3k�������ٵ��	������6�V}ǘ����ST:���Z��_$���^@\V�C�������hR16�|��r)�p;6��c�����g-� [3"�Ml?4�Νe��3�U�����f���Y�b���6���f�&�v���K]����[T&�"�XY���l�@Q�A�7QV(�Oe6�v �җ���ewg�����E�N�9������;����6�69�����"mȍ������o��;ɵ�H��� z�r�d��E���H�S�(�{�`�k����::��6,�$�s�󜳬���uYXZ��>�T����/����O>���m����y�����e�����;�?��k���W�0��! ���������2�@5�UO���5��%�G�<0����g�B�{kcM��v�jR2�*J˲FVhD#�o^ˊ\̩�"�;ګ����5�j���/�$.���pvy2΁0����'rxا�ɝ�L��$S0*�᧵�����ł�Ѱ�i6;^�	gI�޺xkn��,*QP�G12f�3���۶�Z��z�o4�ƚ�����L�`BS�4�	�Rci�� ������$�F�W� ����\ 3wb#�6�R	�m���6~��_���KW�.������XJ=~$�[�� ��,cv͇�Ӂ��./-SނJp Ψ���~��t�����;^W&��5�W�c"��{$3@�t�|�	�2��L��=��(�s&�.V��JN�Ŏ��ʳ��Q���:�?t�v���lVa���1_\r��c�V۟i|���?��g���%a�~Ƀ7��P����I;�P��
�j��7���L7��B?K�:7G4�/�z,�V������,�0NǪk�������3M@���t?���55�:�F]|�P�n`�k�wR5v�nB;�H�`O���=��7��ڲ��&��ޒ���X>��Mk�e~z`�Ƭ�r��э<��ī���� v�#�b=G�x� �=&~��L���~�F�+�ӿ8P�X>ؓ� )}5N����_#�}kE������p�l���6�5! F����JX�L�$��p��y0�������)�srscI>|��|�͖�T8;ũ�"5�:�i�a[��=[;���S�f�a�G�ϥ}�<��wjcA0�����Й���&yHO()@���g�Y���J|����y�.v�5�J��d�ć��,�3Xd7]d�Ee�E&UI�A���ڧ�=�R_`aRL�ł�,k�E;$`��O�{D�2�6�[͖���[ �1!��Y4q�v������ƾ���`fQ�����r������E��A��~Ǆ����M��f���Q'�H��ц�}�`�}v�:`�Q�� K���Mw��X��Z�K<8�{[3���`뭚�a���T���&0�+�;�.��h������k�m��9�>i��%&M�3c�F�i ��A����!C���Ǝ2�y�6+�{����}��B`����3�M���1��ʟ�:�p������TDA�mr�]<{��5�Ы�~VY/�,�%��`��Zձ���Wy|�}���ؠ�\��[�{R!���X%�(�/����	x�#c鲔�1�ȁ]7x72i9p�u�we�`s��蹫 �?�RQ�1����V���O��.lm�Zj�5��ɩ֥�$�D`���ۑ}�ts2˱�s쮿#���An;�����nFwL�6��ES�[L�@R�U>u֠#>�)�
o�X�8IFd{1)���r��t�X�rM�����'��ω��۷��ڵUy��u�u��c�Ԍ���	����<PɊ�GM�c�Z�'���<.v�A�Mf�x �v&7�/�g�x[���r��-e�j)��B����C���]&�e�{���P�	b#E P�UNDyH/��U�����:Fg���V���F 9r�f4�>�)@:�°�2�J "w�N .Px���:��E�QSЅ_����2���e��b�J8�q`��Ϻ͖~�gh-��_J=<�ǭ�V>������(�s=�o(61O�pK.X�A�<7��9��N�'�x;u����rs�&�.&p���q�\	�� S��<lmo���!����&�լ0�/ ��G�! /��g��|���]�{�m�^�����u>��@�'c�.��9Յ����?+��{l*|Y��N�]�Ƽ/Dx��u�c�z�S�^uԇ�u���a��Ғ� ���+r50ު|�{)��R䏹l9�~� ��}F�mUQ���{�]HYT1��/���*�����4��s��r?��)G�zϋ1�j1:<ӿ�`���ю;d���c��MՂ��.��^w0��Z(e(^,`��Y:a��/3��z��c���q.G+wg=�
~(Z��o���Ѐ��~����!������vK�}b�a���N4ٍ��TD5p,�;��sL�4�enp�y+�STj:�������m�hOVV�w)o���ܸ����V�`
��f�L�Ќ�}��< ɾ��=���|�zu�����
�?��o�O���l��ݯ�s�%*-�r�ǉ�Ռhe�J�#��Ѓ	oMX�Eq��5F���ԣM^s���N�-?89����ƪ[�td�'2�v��x*���������Ou y��?�_C0��;�o��h6�>�Ц��t��jd���# �px�{��`��yZ����A��;��t��p���f��/�Y�M�/y��w�X��LG���!�Xp���O>��?z_�~�-�ew��銢��1�j��� 2N���P�ga����-=����Rn����<r�HG�W��Z$�(�,�N_a��s4bU<�a�Pr"�Ӭ�� �UzcE#�8a��Zn�CK��Ժ:΀�^XPv;G�U$��G�>�r]��������+�ɸ����QM�&٤�d^ j�����8�҉/΄ݷ� �j<���|��[L�arS�?�x�����<�Y���$%� ���W�ȕ������a���sk�6�iKP��-����m�P��N�5�;�]�������D�O���9kz?�o����=ܸڬkq3F�m��"#`/R=�A4��&F B�jM�v��렊X��=���p2J`�>�8xr�|�����c9��XrJ������t<��`��?>b	/VQ�I��$�����ɝw>u���^���s̗�2oY��pa��B"��UawON�����'�!Ki�v|<'��ZzXɄ�@�g����V����&)Ɋ[��|zr�V?�vuYV��eieNv�Ne0�h�f�@/�#��Y����E�R��g�Rۛ��pF�~n��P��}��8�T����+2�s��NK�}&snnn��t_��jNyІ�6�`ǈ��Bc:5?�{9�հ>C��J�,*B����Rɐ샾�@�)C�p�y�����_}&~���Y���}kd�W�e?�i�v([�O�h��T�RW������������_���Q��F-.r"��e�g2�Z=���9X����r� �����Wc�[��R#F�1KӺD�� �e���|�I�1��/������[`%�a�;0�Ś�lB��Y�呂݋�ً4g��jp-i5��(3iѿ����R�e�& "�!3� ����1>W�y@��B�x��ycY�x��^������Z��g�������
�mZRr�|��t�\�/gv/�����*����BG4�f=V%3�)��E��p����
���&ȭyk�<R5v��1�M�j9}�5�����Ϸȍei��V����J��\�����H�`�21%I��y�||����Һ�K��!�����G�J�^{��.����
a�-�r�J�|�(�`һ~�L~9fb�o��o�O��t�@���N]7A�/A�O_i�296Q�BSd���<�Ї5b�V�J���uC!�k�+�.'�M9>=�[���3�v����P�����4�0�_�r��ι�FP���=�-�AG	o���|������~����t$_~�5�����ݸqC������o��?�I����_�+��5�S`�⒭� Ȕ"V,30ce~���}��l� ��.1 �E���6��3���n���]�vڴ�B������Ǵi[\\�����~��4�X���`pQ��$��.�/��	� ��1�� �����}! dE�7'�q��Ǣ�z瀆���NQh�뚅����,=25��d��M���uX��;wޕ�7eee�@�_|)���������Ltj���V�l�����gٍq�Dt�Y�񮬬����6o� ���]�5Z�~��ɑ���"�G��ɣGL�F* �jd�z��t3@a�e��v�ε�^�K?g�6��%!��r��uY|^�0yqV�d�e�����~�l���y�4d��HCQi0,?l :�0s� ���۬���ݪ�����Wr�>���5�_�3��G�7�]�f3r�k$�KmY]�#���&��^5�
k/�%c���K�<�� X�h1�g�=��'rLu��Y[�P�lieC6n�'�7ޗNo�I1A�(~H�¥3�$��A �-wW�7��_����o���r����4Z�O��y�s��D�o�$9�LA���ŋ��t�B�7��OK3�P���</ׯ������C�6�W.��Zu��~�^�P�v�s��M�_���6aB��|���_�Z>�����cB�Ƨ��XnݾM����5�:��?~.>��h�{�ݮ챂R�/�s�ɭ#�xF�����(^]Mд���i�&�$�'��A��FӃ�Q<u��;`�u�ԉLF'_��pO&�ԲA����mD���o˃��޽�ekg��8כ�������k����`�6c r(�޺������=�y�;�,��|r�'���,)�,x^#徐Ć��y��5��k���OSސ��~Onn�&PF� ��j�~{��Ȣ����0q��-�w�n�Wh���: '��u�z�:�:�9���2\F�u�~��*����g5������e�1'�� �	��`ˀ���M�l�g�~+���Q�Uͤ !��ɪ���˪c��W�*�4���&��M�m�߶�01͘_�c��Xg��g�2T1���O��6ka�}�;#[���A.�dz.+u]���%�4�Y�T�gn�����E��ﰲ�jɊ�|ޗL��,\�z �Inܞ�+��y��՛pv�<Wbw��/\�w���ܼ���7���uM���Z~���X-�8ͦ(2
�ǩ����{���ޖ�w���esk�-(zn���&�?���22�	'50V� \��N�9�t��\_�ގNe�^YZ��ƍ5����f݊L��:h`;V����g��2��{��  �^IDATT�W��/j1,�uL�ς��|'�Ir*�Β�_]����x߁�ey����G�d� >���� ���7�,��]�j����<����H�RL�\4'C��B-kh9H$���z��E}��}�J�_Su^���
� �"��̻ ����(����~��o=}�m ����.�U�ȁء<�������F�؃{���ݻ��}��ۍk��w��h��`H�7� ]�=#T�����k�Lq��7A��M5�J�E.�7�^/�3��- O²ЉwYe���9�����<E��Ne�o\���5&#�"q`������^>��s�Gq�: �|eh��w$��g�},�|�����[�7gty?-.�J����Ŧ���T]Fh�̹�&�G'r��";�<�Ã>�s� �N�e�,���%$�犯��2[<uvY��~Qߔ��Ϛ5�g�ᵿ�X}U��bxC@���f����e�ge)�m �@0���,�Z1�G���T��2�1cv�µ���v_l+G��KZ��T����P_]���'*7�0�iA0"�f�n�X�Ȗz&G�/��E13��%Q)h6
Y��,Z؍*��Pv8I#?)5�����/��t����x[���q�)6`��̅p�t�ϫ=��K�zg�6_̚�1��}�}w�N�t ��g9:�dyyQ�E���K$2�&X�R2$�:7��A��o�,o� �dH/����LBl���7�h��R8K�K��r~�e�Ky���|p�T?ص�h�V����Q��iB��;�o�o~��[���7_��� ���'w�-���=�6��u���λwd0������%n�k�-Mς�0(��,���1>h�����Ǜ7oK߁�﾿��S9��,$%^������0����Ź���D2�Scȓ� =Rmp���G���0��|O�Z��G�����.��ڪ���`��c Ѓ���e���9�5��K����w.��e̍�1b�mK<�� [�� ��P�muuU>x�}���{��!q���z�-{����x�}0�����8�i2�#����z��Z�[����wnʻ�E9L�&�'�P��X�WN��������zR�F�}�?�A.�����
(Xu����s��04>��`>��6�5����}�y�E�l(C�s�[�V��e-�e�+�F�E��Q�z�p.��� r��$���}v����-Ҟ�:�ڱ~�1�+�gf�cU��j�B�^���[L�� �'��E�"K���F�N�C�hu^�DcsT��i5 hc�k���S����Tz��f�r���S���}ui��9������9����;������r��YY�)��%�y�M�w�uxug^�"~!-��n {��뭁`Yv���D�r���n@=��݇r�2�y���\F~3K���_3n;?o�T�����t���q�+�����/p��l"��T����m�a��h/��.��{�g!�G2 Cn
�Mܱܺ�A�.4�w��F���[.���|��eEVegw��@D�I$���_���GG�p�{A����Hy�(c5�&Ӣ��^߁1�6Lb>�@�k���������r��'�QƃEM��I��d%��4g�H�b�=����<���B�=�0��{`�~�k<w$��:��hv��ﴻ�����廻��������j\xf�;p��Qs�"��T6�!�Ǥ����!^=nث��,���U`�_s�V��cw��� ��~�� a�����s�#������8W� S=2�xӌ^4��r��[��ݽsE�_�ʟ��[�[r�L^�z��|�w���Sy����r ��k����N�؁\���M�c2�	���0A��Yܟ�t�U-��7�������������wƵ
d� �<ps�D�2�O�Z��x~��K�b$���k��[����:�6f�`����G#~-�u����Ӭ���ؿü�R|�B���6l|�
*J播`�u�*VR3����VW�v�Jv�#K�wh_��,5$L ���ld���?Ϭ��o��xC��v��Y�%�zO֮\w��:��徏��	^�4��Z�j��H��K��{�Q[~�O[n����0��N�w�)5q�6Ǿ i����&�C`?�C���Ͷ�Ě�� B�.�c��+�7�C�.�ϑ����s{�v���Yڙ�G��4��%)���(�6�ܼ3KK����M�)��P��o�¯]��g !���-����:���K�5��-��NO��m4[v ��7KW�F���+WW�4����8`���/����q7-�U�+4�q��E�s����� ���KG�S���u��Ɓþ,�\u@i��g����g�Jȗ��Ǉ;o�q�򊬬�3q�g=�/��3�v\���G�+4T2��1��M
��u����y��f�@ >�f��H��o~#�}��ܾ}��ؕ?~�g���f`p�bi�������~�z|���u3����U>C��[]��5�{��<|�H��{ �="�����d:$�H��	���=���t8�p�1N�������1z� Q�#Xj�Ż}�l�E�=L��f��S�]Xz�Za��*Pb��̪f��m��{�#%�C��CU��{e&��3�3�}�?f����v��L�_d4��c:^;�Y?�ת"
�{��Ut1��������SN6Q'�,M����M�d��M�)�V^���둚��`G֤
���(����f�Ɂ 9���%z�8%��Z)yK2�<d#VE0�$��#�����S��n��vl���5��2��n���׵�Œ���h����ƭ��`��|�͟|�����z�Z7�`)����+O��װ)�K?�̊d�"h��p�������%�1k&/�(�&�aTq�����մ�+�����Y�~�曚�=�tS �}�x���0����E�?a��)H��q �Y6hE�Ihl!G���W���g�:�6A-<��0�w�۷o���ui��d� nQ�a�>��dvQel~IL]�1Ԣ�`�x�i�k��{f�3Y��`�@�nG]N ��noﻟ~�y����,,.�4��h�`ze,�������𢎡n������>�T�+��B��lC�#?$~���1���7G^�,��E����G����_�y�&~�����7w�h `��:IU��yzݖ�U&�Ula��]�)�R)�8�
s����w�h_�߿'��R�U2����A ˀ�!���2
�>Oi!wpp@��͂ �2v�,�-s(�����9��1�I�ȇ9�.#�(���Vm/��*�gK�
����г��(��������53v��i�aT�P��ՈC��׮�-@��W�����)��D���"����~6��ɯL�e��vW�u��Y��媇Ed�������i4#6k�6d�זEv#B�2��{�$!?`p�^;j ��^_z����P9;�)�3T!s��Y^�!�˫��$B&o凞�3;�65h���uN�r��\���]��o�+�n�-�~}*��<���o��J��ZҾJ��P�9�'������PC�q���9Z�<��e4��E�5<�f�g�r��&yf|-*����E�F]���﹤Ӻ�~��U��!;XX�cуI��-б��ݻ_���/�jqQx�ﾣ֢{&PX�<�����D.��
z�'O�����q�����<�!��Ҧ�Q���%�� +`�V7����yam��H�T��3�2��o����&�MXaN]f67w�}�c�[�^�2O��.���Z��~����/�k���޵�yvǝ�2v�
5���dr�3�*q�є]υ��E�L�������Vj��N���y@m����#X��K���F�~W���yZU=��I0��C�Py,_}uW�>}�@���;���Ó�	e	C��#6r?{���|���^�؆��N!�hR��R>¸'���<L~��A�s�vv�^v�-������m�6\U�,��U	y���D��!��w�6���sC]�}�$a��]?;O�{��^~|z��Sm����(��ӮY�ݜZ�˴�;M
-|d�c�ͩ�-Y+5�̴D$&��^�M(`F�@�d9(��d���$5+,ezH'�a�lq ^��[�d=vK�E0��ιIn��1�	�3��O� ��kz��oY�_�jMFwc m�o�zG������n�3�[�wܵؕB7xv�~��U��+QV������� �✿���p�LÙ����5��W����':o͕��e�_P�7���{dYjCM�:��uVl�/�AG��n�mD �� OZh@o\����&���<��kH#����G����K�OX��ED��VYfTp���'ą�1��l"�
�kc�J�5Ʀ&�����98�;0~���ޕ��}��Z����V�2�L�b.CSNx��cow����X�u��%d�t�ǉ�y]l�^�'��J<��@etu�H9fӓvcc�,u����^b���V���I���񫏺�D}�r$��pr�ɲ�r�&*~ǟ&�Q?���֎�$=���9w�,�6M���>��I9�=�Z$���圜y���v���`�닑t⶛�F<+�\8Z$�}�_j/:�Y����������;�n��m�)�	X��.U����,M�y�X�����}�E�91�E�1�XE��OQ���ho/Ӟ�)(��zoKN>D~���m�|��7��X���E
$��׳������)�
x��E�ƒ2lf-�z����0�^�d�"�`�Ў�}�YK�͎���$B_�s�25��ݍ*��f���ވ�H*�&� {ҐvoIn��������F�I��my�ȳL%6\�R�vdj�n�K5��!�#�,.��k��H����d�K�g8���Ko�lY��\�H��I��5T]���"�p]@E5+j�E���#�B.J�p�|XZ�ܼ��N�N�zJ ���5&����m�����2�̭۷��`s���"��V.�B�F�['رn-V0���%��>��ڣ\�!>�L���Qd�ݔ!�)=��&����#@���<y�����Ɉ�z Y w0���#y�d��-�/�vvw�O2c:��}F�Ԏ�1�.�ْ�o��,A�X��'�D�9aˋ��x}px(w�~G/[�@���ɸ�y���CƂ�f`�OO��q��t���\��x�9��y���gV���s�F�磣S����L���u�"�*��劋�ɴeÜW	T�kw����O��]y�hSZ�=p���*r��5c�ª^:���,���c�_ 
N߅!�l�<|U��`c��X��z�|��|^TA�2���wނ�\]�~����s���0��y�}U��cj�Yp\�ͼe�ީ�BX3���'��� Re�3�;an�g6���3�#
I�L	�PZ8V�US���	�����,f��y����b�T��BTD�Gl[�a��յ@"�$P�E��f�G-¤�D�DcUx��/���b��+U���|�t��3��7ޒ�ޑ�׾p�b�&�!×�X��zf#ctc/i�\7�i&Z��BI�^V+^K��D����6Z���٦^���&Q𿲌D$|�W�q���y��t�=�=ݨ�薽�m��W�l˲w �CF��"�N�#x�k��?�N<"(��M)g �@i�Fc�Fj)V��{���_ݕ۷o;����H6�uq����d{{S���?@#3Z�qP�,�l����޾l��1�I�GX��{ڇ6�g��4"Qד����SPWx�h�Q)��8wXx�@����XTΣ�.��ܱ�vr��Y�8v���N�r��C��x7��ܹ>�}w챕Ƥ�&jl�!�N¿�5�f���c�r'��IhL4�޻��!E9�j�����3�D�����~�����5I'��馴��nQK����k�ly J�G�� �t���o�ɏ;�O�\~2�Ӌ8c�)���Ikn���"��7�}�F���i�9�sY��Jk��#�&.-�k�tE�s`��/���}hv�}ڲ>*|������J�h`��h���d֦�1��~���%�y��763L�
�Ɗ�����E�z��j!�Sa4��9�v��5������j��z���v��E�����T�w.��T�پ��_~�<v�*� ��j�K�P��<��x:���0Pv��6�K�2��y2�i�5x�[ �V�}x����I j��s�GFRrBA[����}�}�u��/�ؔ-�wE��k z���ت�->����
Y��ʺ��o���7ݤ����!��H/��ye�t���E��ʉ��/L�n�M�6���ie5h�� �u� 
�'V�~�Î>`�s����'�r�'f���/����S{m����k$�E��u����T'ǰ�:���5�_����p�n'��(n w����:=�z媌���������&
7<��\d�΀�"!!m<�C(��䶡o=<8v��W�/l�|g�WnY����re�^ �w,�>}*�~Of���ut�A
P�h�z��/q��{4>&K�k�>����D���
���~x�Z9��fV0ۅ�N-�ؐ&*UaO,ø�gͮ�g�5J����ޞ��<��h�K�п�\�+> ��#��� ����U�wh�����ճ4c|���9o�l�x8����3��J+��N���,V��N��VCz�yZ�-��`���yK�WD�r���M.:�Pv��j^ˬmȒV���h'˟{��<��l��ne`U��E����z�M̾����d?�vY�J��� �g����ڏV݊�=+�S䍥�ް��2-Z�@9	Tk�s��4�H�kq>0N_]�B���Px���Ӽ����"�U�ś�Tkm���{������ �m�Uv��s��Hl��~5�K�L��[���?��J��
FKre���r��� ^w��pe�7�h�����h�vP	i�ꄍ�{���\�ҋ]���܃So��lU�Ug�"�a���vn?�K6_o��h����;��a�x ���rE�84Y�B +X�^�~]�<�"�O�Ǐ���ʊP���'OeqiI>��c�NZ�y�^�)�6vYV�0ˢ<`nIZ�s�q?�b��>`>�z=y��m�����O�t�x�Ӊ�L��#l#����f�䭶�S=$ 0�}�jL$��5� `�Q����?�+ˎk�m2�Fd����s�>���=�6?����C�ZHЗ	����������7�h)yO�tǄ>�:� #!P9o�4�&�a���琶��xc�:+tbEr��Q�����m�Y��b��g���d�>؏5��SMv��2���``�Pj��.v/!h��8VB�g]x���V�7�8������-��אַ�jM��Z~z�vV;Oƀ������F>���� /�C)~��r��b����
:M����f�aM����6A`��C����;���V &�-&[��*�m�3:v�|P������`�1A�Vý�lqrTFEc�P���/�'��W(٬�������ܸ�!ۛ��޶�r�;��e��I����`����t}�XZԆ�Dr� �x��}��nѰԓN��k+0�6�|�u�Ţf�y�`�����~n?�f�u����J�QM��v���[#4<I�@<M�����/��^o�h�I&^A/������`]����ȭ[7^�w�yǍ3*���T丧��{�Djik޸���pU�~���
thc�'�=��u�V��:�Ք�~bOm�da�}$�x��4�+]��Ǽ�\~�s�*��EbU-̧a�T@`l|Z�x��W�PW�<��3����}V!���8�_� i(*V5x諰����$�jN�J �E��Kq�J�ť�+�ք@� GGQ����=m�.X��D5wo1�Z��pl���5�ݪ�:�����q��}�>��.��6C�¬}_�16)���/{���2��~Y�}Ȫ�o�6���c�4��n��3�/y�����۬{��/�㰞O�"�/�����+*V[5c��f��Y�I6p�v���/��&���'C7Ќ��]�ŅU�[X��J���8}�n�����L*���d�!�pq>�n7
�|&�
��:�˞�a�T777� 7�����=�X,���3��A�x����@p�Z�9��-2�p}��lƁ�xwvd�p,�HڡdD���YFM���nbv�w��E�����<�a��~�-wE)=�� �XX\t@C5�xh��48�����B��j���7N��w�}���T���������g���6�����o~��zwg���ԟ�}4�	+7j�9�^�B0����+��Ohʹ*�7��1���ϭJ��b ��n��{8>d����b>��~��A�+���9���]V�M�F�IH-MLգ�I	>���Q�8R�/����=Ʉ��挘O��=�E���"'�8o�?��v����@��Z]�3p�*�a�(���f���"��ЙI8�yPn8N�'cM�x��_�Ҽ$��)H7΍j~h�E���BAf~+�{����_|��z-8&[H���۳��0	+LH+o�y��PW���s�1��B����Ӷ���K&_�
\��U��Y��)0���y ����L���V$�E��a��iE��zl��	�8`�E�"�1g(M�M4�0!�E[��벴rU��r#;�n���c�y�y��]y��<�}����i��@]G�5VR��.u�I���*��;4X+K2l /�%&70\K��Ԡ�i���0���.&0?K�
����*�0�%Oe{�<}|_��F�8�9t�C��E�hx~�A��GM��ە[�����^M�!�Y�7��`��!��`���*ju�r_n7с
@zH����r�*�1�����VS�N�h��...ѱ�G�v~����ӣ���n����E��]YY���Ǹԃ7�.�VV�ؙ� 5-�����=��N����Z���̆�ڝ�	r�.�d>ai���^���g�c�Z=L��V�Y�ݪ�д�R4�V�5�ʾZ>F<�'���-r}�^�^;��p���>!5����2�2c���D��(< �����	��YV��$���{�,�*��T�[rF$�������?q����/��c]@4|1/�P�r�kǤK8^ԏ�y�ek{���1�X�4�����ޒ��c�
�_V�P ������J8���e ���~�vYI�,?�g�n�B�֜�}�6T��e��p������.:�Wyެ�I��f��d\7��t�mW/����m�5��XD��y�~l!�$�q��aB�����s�nȻ�*�k�����-�l��p���W�1���O�`��!�S̭t�����&���sM�"�����4��__H����^L
�����(Ó>'n$wЮ��X�Htr�{������=7�H�'�d,[OɃ�wy����M��{��iYX�I�M:���۩''�I2����mU���5�?dX��N�&��`Od5�P�����(��)��~wg{��he�J^��
<���� �����w��8�,��G�'�=�HTO��[{%\0�I`e%�A�c��m�Jœ�z;�Q΀��D1K(��2�ZleL��Q��W��E��'�%IP񪩺[���}�Z�H�e�TV$L���'i�&�Đ�%�7��X�l� ���,�\�l��R�"�
�jW5�N��D���z�Ȫ!�ZA��Ѯ��z�����ey��YlR�w8类`��,@*pPʐ��M�+�{�29��H�Nܱ�{P�(ӋbHQ�,f����Z�z-�-��k����m��C���
ŗ[UbPv�N��:�E�o�*�1����_�e�� ��Ip���6<��[7,6�k���ˀ�2��S��r?^v�{�^a�.o9	��_0�<�p�kH����t����u@���~'�Y8&'��M&0�g�,�ܔ�+o���-ؖ�&;�+P椢�Ƚ�\�#�ʀ���f���T�G�t�ʟ�8X]'u�M�7L��	lJ��bs�(���[�t|&�@(��:m�c�� 3f�O��a��ڜt�W��>���ߕ�+7� ��вr�^X�&o�:d-�z�헿�t|D��q�z���/����`�:��j�^exC���^��B��d�������E0/�y�5����~S�lb-������0"��e�T �eg�Q���������!h���U&�� U������br��:�Nű p����;4X�TS�l&����}�HT��^�c������&U�6r���ϣ�T�Tf�%��w���Z�`��	k��.�IeYa����m�1WD��n9�Կ���E%���ZƲ��6yp�20�~�G���/ 0a�g��T��	f,���%�:��)_H��B�
�x9�_`I�����h�l�� ��h`�������9p4�Z��X�i�	�`,m��,/��9j�jD
`%wz�}�|��y_^ќ$Hc<�<�{��PԤժ�0H�G)�^x��n/�88g��M�p�q6|?��[U�Rl_�������>B�k�0^�����`�ᶫB��޲}Z���MSn�4�>[G��a�X^>��	��%�|��zV������y�&��}fT��k�����,����q�>Qxh�#?��4�UTT%�XH��b�ǝZ���vgY�\� ���V�v:n��\L\$$2?�B���[w��h�:S��}��Wo�<�nhX0�/�[Z3ț֢��v@�]'��!�"��s�&��ܜ��y�[~��e��M7�`���[�`�F�E�.�n�u�حh�r|�Dv����������Y]�4��|^5�}�-g�в��M}��P-g>�r������5Ȕ��yy��|������>��s�Ei�\�{��T�$"8��I�#_B��"&c���u����^�	��h!	`X�M4Y���!F�c_���|ިmw�M"
	ƛ�x��Ϛ�����3]ѫ��������U]NOh!�����a�/�'c����U���$>ú��_~��r��}���GR� y�,�Gj�|�90��g�R�x WL(&������ c��`X����e.�pX�;����6�7<x���,r�[���~M��x7���&��tb�<�����N�a�ϋ_l���"�X�5�#�x���7�R�u�{�.s`�k:�L�����ŵ=����A�(�-d��������4���3�lz�R���ox�U�w���/b}��φlm�Ϧ�5�C�2^x�.���Is_�q���c�ﶟ�\�y�	�+��Y0Z�o�Sӫ��"�h�j����n����3�9��:�iZc"	*��9 ��,09$����
�D~;Q���%++We��5y�辤��j�|7��e�V�|�R�����|�ӊ?��AC�}}�ҜKKnA�\��������.^q�aR���C�nArmC�o�t���l��d��< ^Lb��y��y��қ%tTi��mK��c��?�	Z���� -���/G��- Y�� �`t���s	@�����:Y�fni���M�
�9  �l�����ƨ� �x�j *��(� C��c�Y�lX�#}�0���XQi�{gZ��A�ɦL�ʔY8EY���O>���ŧ��� ���ͧ��'O�ߗ��c���90�ߏ܋Z��W�kh5zl{-���̙�**�3ڝ��r���^�P�+��pQM=�/�i�At8/h�Q@f0d��4�����0���c����{ߍQ=� w7G �<�����wݵ�3%+�'CZ���='J��tg~W�;s�W��^�8&�.�xO��M�Ex��"5,���ԥH��ھ�s8��"qK�+������ZX\�L����]f`ˡ���l@AD�l�B�ƭ��5�k��µ���Ll`&>R`װ86�~�b,���Y��@�%�ٹX���f�S����/��eEU��D���*]��t�B�~1>L_�ժ6�ax��%��������6ME���u+Qi�3˼5�@�o�Ƀ a���{���\��eV��&bq	��8��|yy�	'�����2�	�V
h�k��O-���F�	�F�5�F��I��i9��V˷V�}Nɇ/ȑy������6A��,,-KwwN��봖C�M�A02؞����PZD9;?�ޯ��~Y�-\�Y���T���4X�Y �M�G���	����urJ ������@*V}��W�_~�5'�$Is&��FV4��M�+��'i������x�9�o�6Sܿw�%q��>y����'O��������p^y��,� |�)�=�a����Ɋ�c��v����7�x�ܹCp�~��ٖG�7�wݱ�
݈	\G�nO�0���Ɠ��xH�4�I�L�j{�Z��,�ZzrT�kq��/���H�h�oZ�h�������dmu��9q��(*����kr���~cÁ�y7�͹��5pf���dx��&nc�Ðt���#?�pU�,$&�:nl\\X��5T�CD��K���=�foi�����3��g��ie��{!���5[M�?���VU�5-��� !�5�Xt��XR��m�WH�/��gM$���9<F���2Z�$�����~��	?W�Fp���jj�i�*�ElChQ�:���|�/��}�m�&?���)?�y~E-�8X�Jx�L�7dW:�Y��.=3Rw�z<hG㸩����Ғ��=2�Y]LG�p�M`,�1�\�~P���?���wVɏ�E�,�B��p�xR'�Ex��j����mܢ��
r���wW�q�4n�EI#��E����h�23{��&��֝����k�1 3B>�f?���+��6��0��ʊ������ޜhu��6b��;r��]d��B7�H��cy��V�8�e>��fR,_�J"nW'6��hV~�A�ɓ����#~ei'�k�ɉ(�_2.�Q�x<�fL]=�֒A:>���k�駟����+���-���o��UYZ\$�I����C�/���n�����羽�C=2u� a>4��6ʣ~ƊC؟��G(�V���#-��>¹E���V3ۣ�?�D�q�����	���0�"x�Ï>�?x_�s/h�1�t�B���1jU���hp� �80����b�#��g��5egE,|n��X����,6��w\�ߒ��'����^q�*�ĴBDDZ�8�z_y,X�2QЯrD,ܢ*��o1fj���!u����Vfq��?S��������,|/�Uo��,�9��᱕�Uժ$e��*Jf@=,+]�ݪ��m��=c��m��]v�����aUҋ�緳�y	��ZL�q.����h�7?G��씤�����T�!V'��HĻ͟��ͱ4ۧҩ����}�lklO4r	�0&)���㖌����P�������?���M~$���;w�Y�@��@D��X�+����}��IP�ohf �-�M���i8G�H^��7a���*:8
��wܐ?�+2ժ�JmW6[�[���(p��b"�Z�v�:_���<z�H����̇�&|���dȬ�9Z�Yܢ/R����D�x�i�ê��Ii�&;�\�0M�ɪ�
�?��s��gfc`�����M��Ga��ܑ�7o��,}�YN�+��\0�XX� �����w�a1���eٸq]n߾�m<������5��q�4�T�Tq]�lC�m~M����K"�3w�d�������*��0#��.0��TG�]�76n�a��۹��}�ں�K����'�6K��6�7�?��ہ��)�$33I/ˊ1~�y��^�G�D�ݓ7o�~�N]��d��+Gº�Q�'���8]�H���{5�w i�u�'=�k����d',F���y�M�|x�3��2 ��ƚ�����n?Շ`ـ_8��
�O��w����e��,w���2x>��e S,n0.���!���ץU���ߗ��v�-/�^���p�������	����v��,��ǯ������l����h��a�STWs+\X�4������L9Q����q��nC����;0\��N�"�f� U{�Ħ�8~E���F��|^�1*�g��yc1�dM���'�_���&��#�{r�~B��G�Rc�ά�15���lh1�;q��C){1���|?ۆ*6��g�w�;�
��U���#�P����N�X���,�Kk�%�kWܘp,���N�@bJ�gr,�jyrX�K����O�̭*�Y}9?�:�ǆV�>է""�jeҐ�p��K�q���j���
4@�Uf-ʭ�֯�˿���N>��S�u���b� A��h�֯s�
iё���t? P���Y���'C&�~8:>�Ldo/�������>�l��A{��Me���fV����ew|��)p]YY�f5������c���b`>�$�sG�E���` x>99&XV�;�,Ξ\�<x��P �e��#{�Bf�������js25�霕�*%��^��ΥG	�`c��`��˿����Q(w�%ڬ�~y��~�>g�@�1�a�`����18^��Z�WU�f����_! /�@�j��e�]f~�����A�E��-�/��M-@�l.J��W1�U�o�����1S�e�'?(9^Ո�J�L�f��D��~�`q-���B��}���&�ӣ(>C%��5�7Yqmai���Qn�F{
C��>��`�m��v9���&D����_�t�z�S��A�1��Y[��y�Ao$Ӗj�����<���.&&�������D���|��+Wo荁��1:��Iot�@Ƒ����}�a��(��DA�,��bUT���Y4��s��m�ӌ�|�(X�+�� /��LF�<���tU������m�CR_�_0�����C�nw�}��r��7��2��j�`���D�J���2��$���S��J?��aǦ�,�j�\"̞z��z������86��]�����Ƶ�=/]��'ǧ���{�?f8{kk��,^GG��=u�52�ݎz�ι�j��t{�)�!���^�F�H������|`�������A���?I��P�F^�ܙ!�IV���������C?�|�-��RY�-ɮ\�"��ͯ��>%����8����;>�30p�pbh��L9<��������Y2��U��qϼ_�g�S�,J�9~bQ��0Z�]��{.��%_��0��Jt Uj�{� ��`Q�/�D�>�{D��]�L@��}�"a�����E��D�놾�����Uf>�@P��l
���ڬ}��AL��6k:���m��9�=��-n��/�.�f,2"�K�ɫnU��y�B��L��6���2��o����D��M�����d�Ɋ��h����$�zQ�w1�U���·�|(/�+A>�"yyE$���=>9�Cz7�����m��!�	�Շd�F�=���ce��B�W�&�����'	B�}iw����9I�Z����5�l���j�.6������	����DR�w?����Ng�M*]�y�����xWj�@&�#Vm�a��c���Ґ_-�-��ޙ�Aq�YV�޼M-<*�uFQ���]�ˬ�_����.O&/d��^�{� �TC���4{2���f��.^Áfi#:�[�\��]j~B�|�\��K.���V*&��Wj�o�V�i��,δ����x. ��hʀcU�X��GGǉ�l�ӧO�o����w���Y�ˁ^�y���I���x@���6_1��{{{d'{�5�}�-j}�3t"�?�Li^)���Ғ��� M��b86+3��_X��x�ۊ����7���[w�y���x���}��nq�l)�A�HHЗp��>�����&.Wk(Kw���{�]ke�5RUXu�l�b�����{�� )-�^W	�h<t�?�B�V��o=n�^9{������ʓ�f�P��8L����ʿ���,Z}
g%U�:�w9ÿ��)/��|��3�ri�2���5�3����m/��G��c,��<��P�CG^nO���8�<Ⓠ���6/^���37��z1zP���Gҝ��������6㯬oȍwX@�p�d��n9�{�&��롾<J�������&]d�!������EēonN��[V�P4a�]���C��H7�\������|�r�(�wy�*�2RX?��; ��T��?�帿�'�>����1Y1��M�F�U��C�7?5�.�8ʺ��a�l�.��>߰��v/�Eb��(�c �C��8p��,�/���tc���a�MӞ�Z�-́(��L��:"5��_?YV�������Y���k��no�L ��a�$ɍʹ__�e<n�4z�z� �^�� �m�`�/c8)���������'O����:�� � �`����=>�P=no[��o&,�0&֒�H4��]@$��{�k��ה�g/�2���,J}x0+���䌱�C�h�F[�x���|q�Ii{������@���>%�b��3&�u�-�)��p�5_�A�0�9]�-����c��<��D�7����M���\I�Zu޲��9��LRT_r$�5���d��;� ���̔��*C�3�˴�1�>˾���Y�󌽺����RyloB��֯��eS!�kU�f���oT�����Ü���.��:�K1�jx3)tM�N0Pf��� T3�ƪ5�Ё�V�s]��b9u ��T�;e0���M
'���l:p��;L��c�� g:��#��� �`O�N�`t�׏�c��M8IĬ���U(Ǽ-׺]��6/}p�-42�8����fW��8�%J�C9�������ED��4��@h���N�!d�=�s��?si��@�4�)�o����k���2��_S_���Fy�a��w)@L�E��l�$�Gj��9;M=�����c�`j�Lr dT�2wn���2�-RQ���aAc�m��� y iJFD�l�ED�@�ѡW�<<ܧ$���q.Ж��@����h�O�\�3ힴ�<�?$[�wkk�l0 ���0;;>j�x�7�_�����|��`��3$��m�a�� }�;��8���c4+���H��e̚w_������1�:�~����k�1�]��@V����ٯq,�{�{r��$�Ks�(��z�pe{�H�Y�mؘ,,�Z����/� ��:��LR�=��%_e��������Lә��"����_:�\��&������Bx����_j[Ad٢���L�]��iF�Q-yN���`�UL��	��p4�zS+��F@��@�ڗ^�˫n�n��P
t_��nBiq�Ci�(�J;�f�+�Z����#7�`5��LXL���� ���v��wR�9��l9i��d�2w� ^����]�1 �-��:�{����G	���w��kЃ��]�����S7��и!Fx����EH�'�I��҆G+95��lץx�􄳟��Ԋ$�ȃNf��� d��ђ�#FXڷVUH�H:�e�Q܂=���(�-�%b�[-�ӕ�^k�35N�r}1N�ʪZ6 ��*�"qD	���uVKp�p����t��������9k���M�_
7X����&ϥ�?�\���1���}�y��٣G���6b�Y-� ���/��t]HN���d`,꒩�#%BR���-��?dq�&�1���ȝױ��p�9>���.�g��2?��R̳��իW�~)�b2� �$&���C`q�n����,/��{�]E�Eo��u�B��3dG�� x��8�@�V��j$m�|3X�M����B'���*���=�^V�z�����0>/�}����� x�Jn�%�pQ˕\~��5z�| oO�E�1ԼTά�[£���O2� |Q��f�3o}��ɂ������!��Ŷd�/R�YrHO�N���
x'�|���1�u��֬��p��=��co���C(/��:��o�G��4���� �%+8P,,`����C2�Kn��� ����t�@�N�$���E)4�*e8=��&�f�=��u������xSVZC8��������p��O�$���g���n���Jo���"P*ǁT	`� X;UlQYS��� �ۨ
�ҮQ��d�qD��b����W���[��ZX��9Xb�i���7��6�nʖI���ّ@`Y�6%�}��2�[`q6��p׃a����w�V�3??�}�3��Ρ^�b  `��-FYC�^x��@���� 4�޵;��9<�є�1xV�D�GQ�b��&Dv�.��7VI�P���b� ���?�Y�v��[B�<�plmm�޾���#��u�_H�0����Lceu�-��q?_~�%���L-Ν�k8z
G���Y���L���m7���G�8--�Qn2gA���^�Os Yi ��W�Ӣ��DK�c����R-S�%�_���f.fռ�υ?/jS���/����뤩}٭*��2�b	@-'9�e86�򛋮�	+bJ`]���'2O�Djm�̊�?��N�礉�A0��op���R7Y��.3/?�7�л���N�"T��F���m8<%C2�$J�$YK�}�	)�)�~�rrt����[$xf� ����rT���v=�e��%�$@2B9C-��{J�s��#�v
ޖ�U��1(�e)X��.�ӧǇ��D�&!�u��7dF�$,q��/�;�G��t�����f�>���������+�ׯ���{)�ml��Wu_�4f�}����R^&��RY0!�K�_�-�}щzJ[�FM���밊�P�`�)����ˇ}$o�y��jg���AF����cVz�������4��	@��fSz�	�D���y���/�.���Yz��/0�h�?H.Q�,�����oXt�����W��x�VizR$ȱ�04�q=�y�ح%��	�~�0�� �'�d��B��|�ReN8��=&�c�E�U�T�{����:lR
 V�l��#Ә��y9���#(:!��;U�g5�Q�z�sQ!Z�R�ӓ}�ٮ�;w6��^c�hl���F��L�m�<q���N�q��{%���U-4��Y�E�(���gV�?�E�Ͽp�/=�n��}g���0��O~L�wV�a���u�U����.hgi�+�-��x$����!���6�~,�Xcj��?��Hn�q{r:r����t�52��tH����jy7�e�jdNc�Z=gx�ԋ�xi�c�)�}�Sh�ܤ���)�>�`oG�w�dq%�n�f��	��x簎��>�UG�D���*�$��(�I�����:3s��H���veށ^��1ðc����d�N8�D>� ���S�f0L���� ��EqE�F3e��/<���gjv\�"��` z�1��IK�ޙ�t֢ eHNÙS�-ˠ��G*��3R��d,��ɔL)ƍ�p����2� �
p�rH��eҫ���(���wr�������İ03z� ��������]��i+�U��
%A S''��望Y�x�|>�̛`�<���cϼ�q@����OsZJ=����Y0�8_�Ȑ?���26�G\0Za��pG���Z�����9VXlԽ���[X���K�	n87�qT�C��Ɉ�����*�QRUSɈ�R��Ld]6`qp|���rVVw�a�7��5�L�^�cjpA���x8�B� �k���b|�Lw]'0,�k�:�U���n��`�&�4&��q�5��.S���[�o,dl>�U �E�_�����IC0�_������^v�r>�u�/��,���gC��Ĵ�TN���k�0X��4Q{ET�D.G2Ut��T��^� �x<⃍�w�l��:@t:@�F&��;
H�p1�YF��o�-��ՠ��d����^J�(� ;I�a n��L�C� ��A�Co���! �e����N��I����ͩL�#7)�9i�^IS�Ds�b�ǵ��NE5}�j�&���6�"�fE+���M�H��t9C���T3��A�˞g��W��]ɿ������l�g-q��Ì�E����y�mV�CBK;�y��[�-�  ��zJ���
��Z|���Ufa�#PָF)T)�ۛ��zˌ�{���p��}���lo�1mH �yV �lz,����Hn]V4�RY�p�.��b,Ө�7��S��/8n����XeH��fǁ@4 �<�k���/
��a;�Z?�b����'�(M��?��;�G��Ϝ.&$;���(7����	A%d�ce�c�0`Z��ĒL�|/@=��x��Z��_��=�X�h����
�ef�Fi�$[uF�����wTӧ�g8���wh��;4�q�����Cr�kb��),���b���t���2��c�Y��*iB �̂bX�Y.HgT���V�:�r���gytE+�i�%J#ɇ�H�pu(��)�μE��(��-h"�r��!��p�V����8�$8���A&k�$�ȒO|7����7���?j�ɳ>0�we�ݔn����D�-�r�����yZ"�oF+��8���J>P}c����t�M*y�3���l�#˩KM����5b�k�����Y��9|��n��w��zc2b�N����ei-����ܴE��׀AH�p�������g�~"���/�q��?���˿�Nw��ߒ?�@��W�����Q#v��N2_J��(���G(T2��"{��L���u>��[��~�!���w��g���'���a�30�t����U&��Z���<u勦Bځ�j��|��u��ޭ�KP��uϙ��h���^k����C�揠ك�Z�uUƶ��:<^��R�T�����n�L �����7�tD�H���i��?ڸ�J0��Q�>��Z�\���qG�N�U�N���R�V�BĘ���j"/��8�=-��(Qc��v�K��Њi�ސ�P�������*j5tc76�� �y��@X5�O���Q�A7���xۏ�=o�1��E�uX
:��^f[Ϻ��J˟���T5[��϶F��D?��hW�uu������ޒp5Y�~�#�g" "��-|��#���ǲ<��\��![Q��#��W�ImU�u���gf���Iؠ�/t;m�q�����ɓ{4=G�V���Ln����9o�?��"2+^��z�/Au���}$�ܗ��.M��͚_5�9���f.K��zȘ��"o.7Q��$��,LF��9<t}|���I�����n��`�yn.2�/ ���0�{Im����Ş�d�:�#�5d�i���~%76�U��|ʄ����,/���ڊ\�~��N ^,����� �1�E��$�ԉb	�]�%��E2�Q��5�[�6Xfֺج��5z��ظA��6���)(jebCi@R�� 9��g�c�[dj�=������\��ܛ2�Y�:p0����uoy���16�Z��J�l,i��~!w��vY^��V\(�L@��4�zf�Ī��HY{�L��0Ge#͎���FlI_(�Q�/�U�k<p��2��9mr��)�W�����'(���VX"FWV����$O���5��	�]T����v��9�"A��]����y�H�J��;T���jȀ�L��v��ğZ�h���2���j����b�g���ٷd��dE�_a�GE]WR]�OR�*������[KZ�	��p$ǧ9��
%�|�a���ݰ�6i�L`�##��G0�&;S����Vc}��F�#�WW�~,�ۛrx�%''W�7��K�5Lu��h5��핍v=F�;��͘dwu�`��Gr||��k�$B�F�)�D&6�4$Rv�n[x6��@�(�E����;���%��೗��R���^�C�*w;���t<���L�}��3�R��Enܸ&~��,.,8�%�{�S�s����¢�+V��+��#R�� T�+����#GGp���
~�ڽu���Zw�������H�&h A-B�ԢtuUwUWk93�n����?�w{{���^����vWu��T:dP 矙;�D���Ȫ�*fD� �p 柛}����2��R)3x�"�r��8l��K�?tq�U?���9l�-HB�l�/���gπ��,��
�ٴ )V��/�^�(V`J��p��k��]Ox��/ ���6 �3t����7�c!� z�@=a��\�A��fhF���&�|���Ը�x���f�	�9�ϳ�4ʆ]���:F���}��{{�̟F���'V3�������^�P<ѢT s��G�楸Z]�VV���/�\��I�ĸN�7��%_�Ri�*�Eu?�8F���!=y�Bݓ^�u�.�lʚބ�6R5[����$�iI��4��0k��'�Vśp�xD�.�=����c�T~d�LҚo^,�ꋣ�ڭǂ :� F�	$�n�CX���{8C�/�r� I�E!0��@�@��ܚA	5��2H�=ek�ͩI�RY�b��b^�5�aI
gD� b%�t��*ty-��1�ԏ`��﷞��:a_M4�h�\@��pG��WF7�����'%IXu�1��pel͂��@�۠/�i��HZ�&Mq2b��T�}�7��Y��Z� w���4zÛܮӐK� �Hs7S§D��xys
<�9��Z��G8�X(%�g�>�V��*�;����3V��{��E�O�|G�������E�8��sc$�Օ�V�X�����3B�  ��Ak�=t�^mr��4����^���C���Ò��F:r�m����d82� �,�OqOy�Z�)�̉S��������皏'�#�-����F0����6�(�t�셒@�B���H{��� ���H���_5�Ǐ�;�>V��2�O��R�����Hy�I�&3�؇��;���K���o�_��_�gR3���dh�q6��s�k"�&��x��j�9k���3�>��ڊγ���Y�\54@�����j�ӥ��5Z^^��k��,�Vȗ�9l��Ad������Mk��]��������c��5�1��M��6	`�����ptm��z>�TGG}8�?��p�e�@6���:�&!J$.�\y���svk�Oo�ڽ�4�T�a1S&��"�rv4���&�V�_�/���q�w�؈��e�Tf��25�U��yA��kl����Sa?�@���| !Y=1xVCe]��~��Q�R'�m�� �N��1��}[J3�X��QF������N7�⍑98�h~77�.�� V�ڄ�V7�C��P�.{i'�P��ӟ4d��QO�g�m&,��BXj�Q�)k3�I��icr�r�6�IS���/3�����Qd`��/_n���.����򚥼�p�E��}�V��oooqyZأ۷����Z�P�j
�,{'�Gp��E_���9�0���X����T������S
�p��K]�|���M�R���:K�q�[MG0��+�EW2���by�E]Q-��������Ĺ�F�œj f4pY2-�Ӕ�F���PE�)gtmhDo�?Ft�P���JFIiړ�y^�����;l�-����y� ]]6��~��ݿ�@�_��Q%O���K/��޽w��O<y�=����5�C*v��xvM��3�A��q��#5*�!bx���U�U�+�$���7�9f4-��Rθg�]��٣Kj�+���v�X�Mr%������5#n��v�St�-Zނpi���7`<�%�ݤ�Oz?��bs�$`=��s��c��)Gb�B�a��T�W~���(��[Ҹ�4O 8����]t��
����TH�ϔaK�"Pe�"mc�_&����8��I8,A(`Ld�\	*c�DԖGKeNM�;��ߟ����{�ԤY��2�X�:��F.�F���LÓ6�1^f��i;vBI�M�0V�!��&~)���?l+�	�I����qt@C5)f1�y����fv�ѱ	y�*y���:����IU
��g��IקVs��!��%?�S�3q�����=4�Kgv���99��Cr�~$f^G��1I�<_uc#�p8Cp����kf�����J���|��^nl�R��,O�1�z���:��sH����^mn������>���U.XQ.�iU�_����=��٣�/������>��O[�<3}I�
�Q��(�pX=���)��=J�r����Z��g^���@*J4&8�}f0�R��ݹ{�n�+���*��屆x�ѫ��z��V���#kg�q_-zR���7
\�Y'�������EP���,R|�M�2	g�t�;��5��筳�Y�W-"��*����B����W�|�8��⚹�����v��}���=}������x�1��Dɩ�솑7\j,D�G�5$J)�q��v�TsV�ޖ*y�ǟ���+	j������!��NQ-\*���D�>;p��z�����E�H�3���)-<�MH���l�Uق���e���"k�w^��S<q�2��&��4��=���<�S<���pR��§)A�6��0�uBu�����ʋX<�ه-ʰs�U�y쩉��b0��ge�V�����۫�u1��F���x��D�{k��&��b��ւ�
@Ԧ�ѡ�4����P�Q�5��O��I�I�;h��#�~:�glNt�{d�]�o9�\�@ҕ�M�
�:jrk���Xm�@g��;�n�C	y�)�wMx�Ð�d�z��g�B$Ɵ"+4�ڻ)M5��A6r�ZՆG�8�)�rr�����Nd��pP����^_�]�W��K����� |]~�⋟�{
��
%�O�����T�+ �ș��:�g�g%1�>/xq��RZ�\fo,���Q�r���ޡF�ŀ�Ⴧ���#>wT(����GE-��r}C_ӪB? ,�R��'���С��ڱ.{+�!�<[���'����k�_ss�s�.��7���>����"k��ŉbj�z��6778zS�١�:f�Zcp�N��L���wL!Y$}�}f�u�����D+7Š�>�2�)�;H�Eh��iG��V��c���q{{W��}Z�_��C�l�x��҈�����;�lV�����|LVP�3C�0���Z�(0@/d���dZ��żupxL��}��~�0� u�%c�#-AG��}������/���In#J�y��$���v��8�^��x�o��^L؀tR�YR���d����
��\˂_QZI��=0��9�	왺�FV����p"��m�vZI���)�$�4�)�D�ڐ�;�uI.p�AgL�'ߑ$��yf>'H��Z^D�I�^m~�sue�2�EJg=���F�VJ0'6� �0�m9ˣFN�PW�
d��҉ Vk	hC��5h��~o�Q�p�ڭ������V�~��T
��i��1Ob��ץ��� \�7�/�S�mm�+��%�/�S���\>�ۤ��Y�s����L�n_ǸDG�!n��>�U�y^\Z������{.��lut"��jk���E�=���U/O��ʳ!�R���.\��E����m����c�K��O>���}��Ɂd{���b�D�<._k��"$��,ؠ���EϞ}�� m�>J�uE3��"�L�3���(�:����wn1��կ~)�x��q_`��u���re�����yH�(�r�}樢�:ͼ��$`8�^H�&<��P�`��TN�J�?�%ޅ�/Z��X�;�'�����9ZYY��\!�X�Y�a���p c鉊��jc�_�ttИf����	Hf�^�tٶA���,��u�����x���o��Ú:�-��)���tK7Z:�1�Λ�@�j����|�-u�bA��"�)���89o�!��7���4��c;'��Q��۬����o��٠w�y(I�aF8�������h���~����	EO�#�.S �_?v�*���K�98��r������pu�a4�8ڜE��0���r8(� ��-:�r�y|�����$.�iow�v_=��R���cZ]8J
�j%����G��x�3�05[���.���G���>�Q�ĉ\�&Q�]��2�]�j2S��������g��ΩV=���F~���\V\ΨZ��9�Q��c�Q��hꈧ���\Hdg瀞=�d.�TW��H`r2�.�]Fh҃��&�LEM��|�B�|�k�Ly/�9.���1(C�����j!�Y �C��pe���NKg~B�+K,��4���C�:������F"��W��Wg������f�=}�Z�=��!'����/�Y��-��A/���\��衺�(��$�"^h���:(
,�:�%E_BM����F��Q)s��`���\Q�va~A�/I})���!�Z������0H�{|[�fx,QB��o�e�%<�ôhqc_��H;'�4O�P֟��;�r�^}��|��-K&*���)a�oʕb ���+,��B$vՎ�t��I>[�B���G?wwv,���0�Gu:��<yB;
H6�S@Ym�e=�#������I��|�Q@>N-�B3��.�G��e�9v��2��fL��g���
x\�NOJL�s����ZV}F����S[� �*��G��2�y�'IC�mҮ��qS�T��9[�;�������N�O8BkR��m�����F^�Չ��ڀ7s4(��}�f˥F�Z���Q� �JV�3 �d�@��I SiS�B\����
K�Nl`���{t�N�J���N��=�ZM�yVm(����"q�8�]pt��(��4�#^�BDDU�A��z��� ��C}���E��?��^]
Z�o�j���A�[�UF�9f\U�Q��PMt�9z�an�a���Ji=7��8Q7tH�|xP ���]ɈG�z:S�D��`�ga|����7�z�۴U��0������4
@�R����ˑ=������Π �V���>�kuz����~N��p�� B>�f�$�$����������4,*����C󴻻��m4�Y���UТ3�+S��g�j
�bިV+@;~[hU���؆;P���0�i]B@	M�n��^��`ຸ�� �]�R3��3�=*˜��餴��<{��:���k誋�ܿ��*��M�
D���D�h�?¢Q���9�`LRM1*�0�������<�X�It9��XQ絠�����~_d�F��fC��Z��Q��].�ܯT�ǜ[�j�{��L�Z ���%�ڋ�a 4�vػ���+�M���7�n�=Ilve1�8n�	N2\�h�G��\�iO�C�iDeO r �.k<#�������^�UF*�b�W��J��q�C�(�r������3 e�.���������-.1<�S�*�
���M�=N��z�)�$��I5b�&�`t �����@�K�����L@�U˄`{Ȳ�t)���@>��z�y�IlϞ�Y��~�&1xB9�/�@�@e�b3�ؐ�k{e �}�˳]��M8;	 ��v���Q��K��}���;ʰ�d4xL�,D��|�,���RZY�ȬN#Q��ߖ���2=L1��*&��񀶶�
 Ԩvؠ\q��y̇S����t>~Zl���Ԯ���'#;��z�y�/lF��L��`eg��ս' I���P!_�n�- ���g	�aV� ����D��H��{��ȏ�޽{T(�����Rd13�V�a~n�L6s/�s���@x��7.o�P�f�pF��Y�y�XT�:Jʪ�
��@5%��`m8R�����q��?��m(+�"岶������d��ZH�k3���_��^�b,_�ؠ��׿�1����Ǭj-�'��O\��H�����x��?Bkp���?x�~���t��m~���/T29G ��TR��2�~ר	��4g[d��Q"���(1�kȎ �h�O]	n0��>{䥜pZ��e_�}j���H�c����f<���!o�{hC��n�; �]��*�Y3�߶���}}������IoW�01N��=6��F9bF��,��<��/�\��rq����3q��
û{xԠ�Â2
k�e�2�#��`(a�^���=3\V�@pxH���=�)�ʆ�)7�R���G��]�U���2���]�7Z����	��۷����d䦲�Q Y{�����X����Wۇ����C���p�Z��6����A������yA���`ws�9�7�N�B��#U�|5��	:3䉸X�rINx�LYQ�d�tH�ܤ;#��d�,W�z�|��j���Ā���7��Y��� k&��gl�h�.	�&�&�٫h3Q�=g\�^tu{�s?K��U��ΚǗDN0*2���C��"���>Z��wr)~F�ty_�:�3����/�B�4� p���o�mA�	(@�������~�Wl��4,�
��J�� ���:��r��R_���|�pmo�qeIO�_���(�� 1��C��KyQu�(�B_�A��*�`�����H(���crD��a8��;��n�y�1��E<�(�ߙw뺣��\���Z�c��������t  �T,r�Z.�ŗ�@(iH,��'nݺ�N(]`���ad_MaW׬��eV���m�ȋktv�j�IP��3ǉ
qP�gW�W1Ud���3ME@��D�:%8BQy g�*1�є�	���[�H��&�Ȁ������4�������2���^����&����ws�&��u�t�M��󁓾��+���Ԓ�֒�Z;'�8����B�������1()�L&z��<���aԡ,���������=nS��
Fye�s4�P����	�u��)Ir�Y
&%!+��EQJ��������ltyDAx2� uV�m�e�W�Q}O �y�1�o��/��7_S�~H��'�y)�$&�ڱ0[JTh-PeÐ��	��ژ��DLu�ܺ����n{�}j�	��Ju.~����A}N/77�S�٧���om����ʨ�T��|��jQ爐$&]$������l���u�bS�����Ao��j;���� b@�u�G'k�zԞ��9�<1�ӛ�Ѯ�d^���Y�E�eO2���㥇�&�o���Y:��h6��oE �#���J����|xJ��Bq��P��������U���~D�\����igo��
�K����;�׿�����K� 2��ֆ> �6[-)ڐ4|@wee�~��O�#��߾�Fm�S`�e�(dӄf5d{����aS./�x�}m�F���HvS6��}4�)���X(1���ns[&�2���J�q�ƀ����2Aq`~=snSQ��k�9�d)�Rb�y������z�8�`���|M�!~���Y��
� ���u��V9��h*X������c���*{4�<&����ǳ	��I��jr�� ƞQ�as�'Zރ�Oj��ڿTS���H��J^<����v�x\UM��~UQvp%!-�{P���'���Hf� ��'Qy�zI�3�?Y!���'�<��dN8��wʶ����A7�'�x��\�\F�q��I�?ob�i�4�V43��}��{kL�[�$��q
�+�G`�.'���=�~�5���_�$	�� n�&b�3?�	�k��Z�/)#0H��y���!�DEz�Ox�P�:�I�2g�����.�Ҏ�i��G��T�U�jttܣԫ=
U�
����}*͕�aڧ�'��������(_���Wh^���(�6妛�����n�(��B�>`o	��[���n�R������8�S��=�z�E�5���X���,U�Մ�qX�$2��l���Xmw�h�I��$Ч|�r�W7�Pg]��90�hw��67vio�@�}�9�<&��h��p~/�]7��xt�^]���1F�����&��CW ��Uc�K %*0B9��*P�p>@z &�9<�ٌPu@M��Im �)��a���wv���*��=�k5T��L�w V$_����X�|���r� Ts��NJr�zt����U���q��P��I0�r����)8Fg��9�"t.�-�)]f4�����~UnBG�D������(�Z*��N��X�b �gT�xb�ž@B�
����,dMR�g���͍�$�~�|�����p$
�+>:�F˫��SdP�օH��/�U�ڈˀ}e��]���yV(����P� ~7�ĸ^�?��X�x�������ӆW�q	��x�qAG=,�_��*�%�g�$�{I�*m������-������Ҽg?����=�Wu|�@���X��<�C�Q�����(�ܑġ����VH	�Xq��u���4�.�T����+,S�/(�6 ?M{�(.g	�W��'��Б�6�>&TT[P�j]�����Ĕ���i�qm�j�]�lH���#J�	v~aNMV���&�~�M/_l�ӧ;���Z\�C�eelq.9^�c����"�!&�9*%�,u�ub��I�8	gvZu�nR�����RJM��7���.��l��e�5��n��\�LKK�im�>ݺu_ � м<�ߥ��gtp y�C5�t��T�Y�D��F�� �1�
Gܫ�=�|�KՃw/]���!^V���o�IjI�w�A<k��Mj�u�0r ��N�1�6�\pq��VZ�T (�� m����"��9����@h* ��񊿋D5 ���]Q���s:��E������� �h�?�v�!�aT��~Q�
 ���I�u��i���#�.�K	���TI�8劼��t���-z��%S�0�\p"�Ru�R���¿T^cc�d0Db`����Z�"�v����A�镹��q�����<N4A��Or�M�q��v_�_�j5_�s�Y��y��U�@T�[^Yc����Wxߑ���7�^�7�Po׼'t� 2G�#��4�wx��~��������q̜E��8GG�I��J|�T�k��w��,C��:��BC(���oA���M���̹ڥ�M4�*<��5�c��>�aIY��
�H��R�sWT���}Ell@T�]=۷���\e�6^lѫ�m��?P�!OP� %�<q t��_��}e@3p�+�\V`IW�!a\��5	!�)�PImE��t��;�/�S6W�V���vO��x�x�D�o�m
6��w����
}��Z[]��W�,�_������}��{�U�W)��d���~��p���,�L,)]Y@��Xn��R W���&�	M�e|�Մ�;�zUM�;T=�+ 2������-r�~���]*��H�I�ͽ�1������7����2�U:T���eG3��m@�i��c�\5��j��<y����9u�4�dBGl:3���j�4NQRr�u�B-ZP�_�����񅳋���	�nW��#��7[*�u�	����(p1�0϶����4� p�y~\�l��0�p��+%�������Ʀ�ۀ��{��x��}����.*�" ���\�%�)�E�qC	���V�EG8���M�!��B�Q�Z͎Zઅf�� �o(�3��6��q�k �8XT�-���s���}���X(Cc��?�|� qP����Z'�x1�����d:�x��7'� a�
�\Dcc�9K��c���b��.�Q�b��NE�q�n}>' ���� �"�	�)�69�\DOs��U���;�(�~�}�2u� ��q�X�x�⟽��~V� ?Y-��U`�8=^�`��4J)c�&�g���CK!]��j���nl�wR3��u�^��z�N$��	���ɂ^�?��j�a�Z��?d�[F�N$T{^�g�/����Qz������˗�(Ք�q=�0���Z� ������<y���j�XY��ϓ��CL��K�
�>�����z�\��f��F�k#ϩIq�+����*��>�j������-)��ZfНN�䁚dv��K$�uhai�*kj���2y�8��=MV��h4G���]��A�'�~��&xm��mR�sL���Ȧ�xF�i�#��SW�����X���ם����GҽG?���-hǱ��re��WH@��>��5��x����5A��}�r�\>�z��1y�r��������&���A��}�(.�M3n��p��7��$��m���g@;�	="���^J*�Y7�% �[�^�|����Q
)��'���s��	���������`���Y�# 5` �+@
��
s;���˯Գ��A���$9o�~I���'G��VW+�p��<�Vk\��YҪ�l�
%�i˺�TC��7~O�@��Z���@���Y�Zy�0.���K1��7�]Ҟ�04\|��M�l4�
�n���/^R&�z����ӋR��<ӵ�1HPV�
0b�QC��b ��n|8��y �1��Erp!d>1�M� �|��}�t=�g��Fc��>Ʋ��E��㼇B�@�=,Z�Y,��x',�p����:�h�&�/�]5���\���c�6��,{�ڴ�-���#����-�8X� ����A�SϮz�=��.�ᱨ�.(j�Li B� 7Z�1�E�+�Ǐ�e��߿�Z�C::�e�C`�-��:tp�P;FŢ�2j/:�sxSo����d)x�$PQ`wy���!JK� ��q�\����Xs�Z���~�`�����l�R�|S)5z-/�ӜZկ�^P}Y���y����677i��*�im��ߺ��l^aTTR@�V�a���� ��/1��
��=R�zU��=e��=T �E�7_��\	�6ij��`ow��G�)��A=x���2�K���~J��G��*���C#t(T���Ls�y������A��?�d��^�5ߦ���Ay7L���ӳg;��]U@��ο�0mJ��"��3$,�Ɍ��0)��MjӲp_gp��X�����G���]��L�BA�S"�X���o����_�w�D��8\���h��u���J�_�� <� 8� cA	�R��$Ɍ��2�<L���*��&=���/�K�r������ Z I^R�@��&E\����y��(�y�gB��v��։SX�
X� �T�n�������]_.ȀH��t8$r;�\��hJj%#׃�9G�.�Xiבjuǵ/Dp��c��Ȓ�%��P����X�ŗ� �* �-�H��ɹH�5]	���5�13IfhXX�|
�<�l�=o.�Y�In�ZgE	\{H���8��ٳ�������rQ�}���~7�Ɋ���n��0��ݒ��͇���7ɡ0K3��Nʾ,�y�f{xM���d�dwtށ�G�粯���A��S+��j�]fL	Z�Y6��ϬX���}�}��ǜI��Uvux�a�((TR��A;�5*Wrl��RT�I�v�x����g�&V��+4����g�%ohʆ�ie�0����	�b�n��;�f�[���X��`�ێ2x�t�2
P޽�H�bN�6k	��2d��p�1�ǳ8���K��t���bM��ö�,|Izh�n��P���ɼ�;P����<s��a�j�m5q��dQ�	z�����-�s/ޢb�.-,��1Y`���}��rJ���u���u��������}�c��|�VB�j(�����
|�˖��e�_�ɉ�B��$�{�M� �j@�����\��e����Ȧ]���D�����d+��!K���3 !��� ��^���üYW?c��mJ�{��+�iQ�*�k�����e��³�(hMX�<Y	�{�����X��%��e�dJk;��-��8���!I! dY~F`��#�W�c}ږ�g?�_��)F/)
Z��j��0�~3�����,�(K�x��AHv-z�c;�U�|=Z��@']�!v�+�EϬѩ���'V_)������Tx]}�`��j��=��������t�Bg8��;D7<��ET[*M�X�{z|�7<�G�*��p�*j>�Iګpe6�서8xX=�(�$��$j��DP�I8�b$�'2�,��^��,��y�h�0���m��;�@�,}~�����8o6�<�b?��ߟ4�a��� �p��e޽�E��K�s�2�Ks�<�	�ș9zv=�S�|��U�裏9�⛯�QƢ��Ll�C���w�qчMgE2�s8	#����
 ��+�N�З\R��Ef�l��E0��~_�m����l�^����,�C�i���i�W�R������"ݾ�B�vW����!�)ЋD�^�+�!�-_(qr��ƌ��������mePq�n��UӜp@� .3,�6?W�R!�&zI�8��g�&TI�H�x@=bnq���uxo1�<�8���E�N�#)ۜJC0��o���6����
B5	u�蔧���vۧ��&=�G��7�a��Bs��v�q|7ƕ�H{]^�7�`��Y2�U��C�� �L[ wW�χ��8��Z���a7�����y�:��\K��<#� ��*[ ٩C�z π%S�$�����d���	K�[���j�^t�R��BB��x�PjX8����:�B���i}ب�/�FFrZ�}dWm�x��\>�x�㍵g5�Ȟ8M�Ur�e,�3*��}��p�����Ox�u"1S�t���|�l&�t�}�,��++���dD8*Dc�ô6�ryQ��ë��9�s���ˋ*�	Hq�R�&#�n�?=>��<�3�� U^�͍���@5���YɃ���M�E�y��h>Wm�CN����Ϧ���vQ vZ����Yڛ)�Ho��{�zT�3�l/;Oeڽ4��I���D�xr�uĉ��j�\ 
+�TV��*"w���
s,V�z��О�1�~9��?xL�<~���n��ޑ��M3$p��A�ۯ)�W����P!ȰeW�B�=�@�iO��]-�.�0:=WK��{i������"5�Whkp��Ҽ?��V��k�e�E�A>���{�� I�a/�jI�7�v�a��ݮz9�hK�'�@K8�D�b��RȩI2�>���!��ݨR�6`�$���.O:�LV���@c�`��@�e�E�S�l�j��)�@�<Yc�QT�?첱6�=�QΠT�Z������{.���I1#Rg�n�6wWkW針޶kngY�߄�;-n� �N�FE����P�c{{;�#c0�����\N8�9�
\�lo�(^?r�H*�	+x���#��$� K�c///KZM�|$�i�RFBqT���@<��gR�"��H��
#�����ʃA�Xj#hJ�QW0�aH{!����|��[|�YJ���wb���k�i�.�p��ڧQ�^�/ڽ��1L+��ť��������N��u��p�0 ��;j�x����O�6	��Ќę��Ţʷ�7����>�����2���S{�91�����?�}}S���S���;^%��6��Q�:촶�N��o����-\y�����Z�9Z[]�{�pU��n�G'�[�����!D�x�����d"wXa[�&�7��j�uB+��W�g'�d�|�VP��R)���<ULcH;9�tgo�e`Y#L�r�
�{'��ZP�s�r�����r�7���� �� ���'����� g�(�$}tS��b�c=IGdm�8�Jo�+Nyz29l��\W�ߣL�B×$�C��aD��
xw;��?�j_Yu�}��:�'O7�Ӧ�J����9r�!�]g즸���{nBK��M��:��4/��7n���*�k.ǋd��������]���s��S���a�V��r�D=?g�Jd�4���z^���}`ww��������*�I�����^Z;�̈́	l�*`6�5���ٿ��0��1`M��꒚) 1����s(�l :��H�������3�<}�8��5���Z|��u����1�k�����3�^PgYc��w�xpzS�N�Q��l��	���1=N��������M�6�b*����(�>g��b��p��/&�D�˜��~��7ݞOe�`!���V��x�Lzjߵ��#^^7�M$�=�#y��]�s�>�J��fX� ���ƖYxnN$��Sr��=Φ��)� �1��e9����qo�x"��)�U���j�	&��{D����ʾ!�ň���o����������]J�c��@xL��`�P��٬S*-:���@_ȕ8\
����yʀ��'v�B�q���Q��\���Z��@F�w��ȅ9�(�Zj������8w��S$S�2t�c�@ȘhjE�P"®�2��v3�QJ{j�����+z��[��M+ �IJJg�މ<��gF�O4�as�漝,�ܦ��4f��X���H���������WM=���k�8㒹�}^��X%-����e�w�� ~�#.:�����//B�H\�@<����/<Y瞏���p%��k@��?��!m���&7�	'�B�E5���(ZF���%���Hc��8`�m�AB1J*�y<8bc<��]k���2�Q]N�K�w|]S(��р2�\}��R�6�<x��kl�M��.�mnSM��8�g}�����樛�D�A^��R7&��:�3���&�i�k�=漝�n`���<��,4�Pɂ���C�|�)���_Ѓ��(����9c����O�xH��Z�G/^<c� {>I<��G�����2�u��-r��[y/���'������,���"9�6�a7�kZ�(�}�n�H��Ct:�B("�i�U;'hX��s��Zm�I�4���Fu��@	I^rؕ3w��t5��:�;�o�'r�Z�'�Q�Td}zjҪ���+2��4W���IS v��0{��D�C�>�l:��r�;;U����Xs����Qo>�N�wϑ�K��ܛ���a��=ɞ�IH[�����$��9]� Pa{��Z_����;�D&*?
�s^��i��&�n�E3E<-�h�k��c^���p(d�]�ͤf�A�j�gȔ�:;!�_�̂� ��0Fc�V�����Q4�_H���flqN�a�����µ�Ň�`��J�������ų{R��ۀ]���`cҶ�����5��V_��ZewG���4����L���i�	o�:/ ��<_�>L�7��?�vv�f8�Q%q�
e�������ݽ��ej� 0�Q�B5��L�|���)�K:!���U�~H�8��"֭=,�rQ�c�X�%JZ��6m��*Pi`+J���K�������'˿��� �.�=��#��.��|*��:�z_���R����5�a0d�퐳���51I0��&� �=�C�ϼ/�i�`���R��#�+\�	[5�zQ�¡�ZP��:�W�z�MYx`��4�Wt�x�Ba�n�����H�z����2�.���l�
�>�R�8n&�gU
�~o�Y�zCƺ	�I��m{M�S���g��	]�'���h����e$᧑�-�3��R����j�J�B��(j"]|����f�X%mo��9?\�{6P����v�\S�,�Ł�݌����)�H�����Ң��h���:��:W���_Q�p4`v��ńV�ک�3�4\\KCI1��E�\#��,2��0���C{ȍ��>�8@=�M�(����ᙓ�BI���@���'���IM*L����i��u6Y��|�&y��.��7m��f0*�$"��U*���L����w��#-.�*;���������h�M�ğ~�){x������Rt����#�kP
��t|�*CX�Kgi}u��%�J�<K�p�[.�9� NMP�c�jz
�-��H��!h7�Lg��A��(4Ԩݪ� *��hojDP6�-϶�V�p�������R@����V �����4W)Q���v!1_�\9ɘ��� uv��q��0��h�&�r��+�4ա��+�O�J% �h	"xc����R�R0l�mw�=`/3<�����T;n���<�o�{A��� Ey��T`��>&9L�i/��vs]f���M�&��<�u��9����+�y��{q/���%%#E��P�SĚ�I	Lz�6x2����I�<�}a@�K�Sh7'�/ ����N�ȴ�=���^ާO��
l�H��TEs�$0��X��v�����p$IlIʙ�%��n�xF�,�֋J��
�\X�X{��E��흟j/�>�u��Q_Ȁn�&B	`��3�]�Ҝ�)��ݞ�ӳ��π�XT�3ό�i�ސ������@�}ǙxŒ s�r�{@�E�p���b9"�q����q"�G�<���ß�L���h��#���{k:3�'�:b�AI�w�y�w��߿V �M���td\�D0��+P`���[ b�@��g��H��/^J���,�� �
��aDJf�w(�[j�:zUu�C��v���Q�ߚ�u��͇�q�3�נ7$N^�v}tՊ���j����C&	����=�
�����ù�"b�֓�~c!�,BMgp��vR\!j��?jrYZ���\������q�aO�pT�x��[���c/d#����\�̅@@e�������+j6�C-�B�&X�� u�T:=�:�ߤdE�.��꽹�����I����:m�q�;k�&��9��l܋�6�Φ��G߈�W6�Njg�t� Ԧe$��cߋ�w��mS.�]ĀTC1�;A�x���Y>s��ax��S"Q�k�q�v��r��aj�^�c5�^��<��C�I�6g���L�'��My&ϼ�S�%��ܕs,�Ǿa�;|̤��П�hg�9�{r�Y�j"��2�v��3�Ϥ��T{5�+���i
*"J�w��?�9����?��{��B:��1��Fφ��$�0ԜT�������?�G�t�
l6�^;�,�Jw ��ep�|j*PF��� 	�A�0��(�n�\�~�K�~�� �~��\h!͙u�t�O���o+�T���@n����q\e�����3�<9� �� 3��᪡��|6�.�9:
�ie��U� ڻH A����U��IKKEZ\T 2됗qG<XW&����y�Er��RE�Z�y�H�[V�#7K��Pg��M�=^�=�	ڐ];�ߥc�3���,�5x�b����Sz�y�@{����L.˚��e�M���C-�����]v�A�yp�t��v�Ԣ	9�|�_t�m֤��$b�^d.���,&d��h�t����﮽��w�9���}l��k�T vE �Z�	�Z3i�ܤ�����_̾�^�RL�e�D$G�Q2"�k`��K En�@���O�=|��
,Af�����q-�B������=���d����o
t�H�@h]�f`�D�&W
*���4O��8�AO��a�/sl�����d�(Bd�2�@�N�ɯv���{H�NC<��(Q�(Ύ�R%�9������kG�ྟR �H��9*�iaq��P���Zt�ύgtt�C�N�R���=*P�rZC8��rT���_��ծ�'���q㈕�VS�E�"Wd���Y<��}w������(Q\��|�+>�����o��ՎPi��X�3�Ǆg�?h�o"���/�����m?�6+b���(%��������u�i�����8��L���W�W��(����}ڞ[㵵�e�o�V�H�^M[�\�x��M�^�ct��hc�N@oLb��dFg/�8�:~�m?���ŋ���0%���5�́�;�误ߣ�?�9���w��������^�B��t�#gњh��<���ܼ�$V���?���L���}���U���(��2�EU�`��n��e7=���ϠatOgO����ii�a��tZ*���:�����i�kQ��d�n�u��n��-����ƠF'��X'�f{��[Cx9 zj@�s�P���ޣ;w���ʪs�:�~�EۛO��o����������W;���lJK2��`�\,�R��hp��L�\��3/�^���V۳Pr�����  ���P�5F�_]�}Ө7�Y�8�K3p=�ї_>��l���}�s6_`�L�p� z;��N�oΘ�N
��m?��Tf/q��vx}���±��Է�\��lg�*;9q��c��`���{6Ud���0����=�ϸW�&����D�������E�h��lW����l��u�iT���4v&��Xш�E��i�=���g�:[�m`�g|Q�۸Q���� ��^vq�L�������~N�RI�S���,����3�������a�z����O?���-�����X�k0�Yy@�����j�c~��GE�~:Z�;2v[ש��Q&�a�Z.��=�s(2�}�㴨�m3aeq��uR��;r2��������HCޥ��mZ^}H��CK+��P�'��̢I�/̓�F�W��ʸ�n?�zm����ڟ�jΈ�`�F!?V�p%qeSM�Mȥ�*r�8�$S�X��o
��})4���t�TkT����)��W�j���!}�����txXcZh(���L[��N��'"���݌
BI��-�~sڴ�c �-%6M*l�}^���٦�KR)��K&�3��=�f��q�[[��,��f�^�X�z�i������_N�vS�ڙ4OQ2��u�K�nc^~�-�;�W���&.�m|foO�|�:#�DS����w��O>�������?�r�p�`׉�^	���ቕ���ha~��}����~l��>}N�F�]��{H؂�S`�O�5h8� pʥ���:�r�c��:�L��@Z;J����r�3����2�zvE�"	���41�$�2A(�}A�Ⱥ�9Z���>����*��@(���a�#
j�9P32��n��~�J9]n���9a.��DE|�9IDj��M�6��q]���)JᒄK3�:-j��j�@��|��A/��/����6�ۯ_P*�( �W�Ud���]:��X�^k�y`�4��MEo��v�vCn�T�a�Y&�$�洬��z�<��dɦ5��BܻUӀ֦�`��f�=m��c<i�M�x��uZ��x��ҏ:W�u{w߶�ӦF}&���xx�ڡ+�A(�!A�׿�ݺuK�u�H6i����ʂW ��C5�aѺD������j���c����}�����*��1`�S: lp��v�C�6�i8���5zp�n����|�
y�զ(�����B��8�L��AH��K���8L:�U�4�7 ��� �:�Rȗ8A-tT�,*�8��dZs\=N@sF>�l�H+k���h��j��@wzw�@��mC�s�W���%��<� k�O�z���ζ�X�@	g軛�s�6�vik�J_~��vwX8�(/�9@(��C�XЪH��<1�Şp��ہ���8��vN���"��k��عf�;eL&����/M�i��"<^��8�W�����1J������ׄ��^��8N�y�s���lN�[����v�}����5#��c�B�}l�	l?����/�����Wݒ�p&n�)	��m��e�'�g��eݓ��OR��i����xgm:�8-j�V��S�+r�Ç��?�)������s���=���AyzO�idh}ꙍH'�	�X��,�ŝXy�֭u���OX�v���>'��Õ� M��^O�~v;)ë^���t*���:i���%�ߺj�dd����E5.o*7�c����������ٲ������J2Cr"�\6v��AW2+Uhqy��VoQ���Σ��|��E�����*�.����pe�)/d}�6�W����hS�LV}��lmnV�'���(V489�K�x��=2o��drr�C�AD��F7KB�@�{�ߓZ8v;��f	��7<4�{�}�i!��`8��chVxI��1񄻑0���Ž��#7��w���s��[&yo�-ɫ|�rZ�e�s��i����h"�e9�Z_p�\�aH��1>+������(g[�_���?�ݔ6	�^E)n��L�踎΁����G�������������޽{�O�1"�h�����x�F�8�m�"���m�nye�~��_��������_�������`" W`-h;;��t��R�7�վ
�� ޠR0xd�k&O�>7�־.#L֘��]u�-��/(@�����>;֒L	���e���5����U�Pr��������8��:�@^rQl��P����&2W>g�ܡ^	�x�<'��5z�j����)�|�Mǵ��S���9pH��<t����y�Y�ue��(p�&t�0��6mb�!��it����z�޶�l�e��FF(ϼ�M���FOy�"������4��e��W��a�'âE�x-����2�������w���s���j����	��˫'.���d���g�Ѡ�@�>;8ܗ�;)�cNx����������7�C�s{��V�)�s)å�E37厯���F`����CB �4�o�'��O^�"��l,*���P�E\Ѧ�t'�2����+��͕��͑���������D���DZ����]x��>@���r�j�
ж�C�7Xk���m�R���.e�K�*)����/l�������xR���E��`����:[�P���{��6A�'�w:F� \y�f_ބ�?�M��_�y����m����`�"#�1?���d�K��m��b9f[8�{�~��]�1����?�����/5_��J@�C��2b�|�*ji��'����5[-j�W�v�T����BH�}��v�-j6��V�����R�Re)��"̟rY���v���^��
f�mJk��c��x2��$������S*�D1�^9���*@٦���,���2��<���
���/[�+Q�8K�fJ�w���d�HG
Ǝ�3|�u�| �s�4{x�� ?�Xs�Z:G�4��g��0e��o�ѓ����|^�t��Nb��}Ve`?�%��3'��.ВxMI�EC�S��L3���:t2��6k1�I@�&���䞆�[�{�-~Mmnṯ���œL̀��z�����<�K>Τ���i��e���s�]v�� ^�/G%�|>O�r�~����?��?��~�3�3T��j�^�+�����s�������ɠ��˗���C�|N}�W����3H�u��l���>'q����^���EZZ�����d.����@g0 ������0��2��1���ut����M!��}ԏ���j�'��] �aN���i4)��8̹�wt
�K��E�� �н�"�\Y$@z�4���a^퀺��rԏ�T�Wicc�66����7�jiJ�\a�)�$����r͸�����r��;�Os���_���'ﾡ 9�{Ӯ���%�-^[�o*�}�~xmR�hR2�����k�NI����&}ﭧ��k� �Yr).���q�de$�좁��.�����{�1� ��{͛��� �U~$$��|�R��>�����4T�tow_<���D0W���xXX�v��m�rZ��j5�V��Vo��w��r�P)�*�rR<��!�'��(�����\Ǹщe��ʙ05���-����*�UV��A�ÊR�w�oҠ�T'�U��S%Q����JD*1v�L0%�+
K
G^�s:1ϕj"�U�r��nw@;;G
��ѓ'/hkg�vڔ�e�P,QN^�JC��\)��F���S	e���ܧoX�q�H8�Q����MJ��&���>&�Y'��~�q��&p�����>�o�dc�묙�I������)���Ki�v�K'g�*f�r����Y��g�P��Ӿw)�0�Ѿ�6���8���u_������{���5?OKR����Ug�hL�2n��J� ������_��������>�;�I��:�?�pi�i
-v|u9��.�-�,�����*@V��B�;;T;:d�qړJd����Bh��)T���ՏQTa���T�t��2ݺ�D++�X�\^$ϼ4@hWVO����2t"�.�p��������Ɛ�hii����*U7էC��-+�����}�r�j�w��㶨�o���bU�t�Q�9�@�a�
��1u 1Ń2G7�����NV�~=�zt�>���h{k�^m���a� p��{C.}�b��4'灯+da�\]�����&��M( .�e����*I}���8��-j6�����q�32q����I�w��$�G|5{Z?�;��A���,�5���Hh(9�t��N2"�ŹZI�1��=[�ƼwC<��C|IǙ�>9��v����s�P�}Bs��� �U'��ڒ��I��f�	T�imR��pf���w�������7s�My]�~f�s0`�"I����>�Yn'���\�yL���(��]�  �Q�/C��Ϯ�a�5@y�����7��g���}Ĵ9�w�hV�;�F���3�KwT.a���%��?c �����o���S�����1�V(˖9$���Մ�C�y��n_�՛t��a���\��xA�\��uk��1���b�}u�HZk0�2��K��̈́
����:5��~�.��F���pЦv��&��^�Hzj5�j���y��5T��V�a_+[�89⅖� jrw�
D�}��%)�ի]���c��N���F��t��!�
�ڇ�q�jΰ3�ޢ=  ��&�����0��k�f����V$��?��:������L^;�B������`���Nx�g��&�I�Y=�g��'�g��\'��=��M|�q��vM����I�R������]�z��P��&5�oWIhq������v���<��v"�ifqa{s�������/,,0��?�/����;whee���<��ͣ[R4�k0.k�Rf��G����2�����ӗ_�����f)���)P����+9�����l5hw�������F�n-ѭ�%Z_[b,
Z=�� z��.�� XsE6 lO�I��t��8�P�T�;��� =��f����e���@q"`8ĝ6
nTy ��1�'��� �)�
b�$)�驕�������
�S�ݤ��=�~����a��V�>�laN��ާ$�!���ti/��!Ư��si�gx�n��m��-�+7�Ӏ!>�AD3�޸���F�4Л�������Ծm�Mί���E�uo�$`~�v�����E�M�]�n��v�w�7��Okv��2���+�1���9Z#+��� Gއ8����/��#����u��/����19��$		�a���sR[.��o���677)P�V$fS,&�~���!��XR��C�vm9
�v����!�+л�4OKs
�B���h!��>�$E+����UQ���E P���m�1k���J��ͺ:a��^���2��u��n��@6˞9)}��h�	'��3���@u0p��R��a���Q�����=���*� ?��>�˫>�pF�v�y	�$1�Mib��%�Z��a�q#'�ʖw3��l'���:�h8�Wg]m�����'x�����>�k�9�cg{{�QQ��d@�)�`OT���>L{��/潿
04|�[�8���*���5�%^߳R��Ɵ�kj��	�.o���'��5����t�v���h;��"��$�h�5�n�������]����۷�ѣG�����{�)��]�#p&�k7��#./:̮l���~I��s�2����Q��C�~_@���šq2���@�N��X���C;;�(��.���w��w���"-̕��EJ��QyM�.B7�x��:���� �ק^��<\T6+�+TT =����$���t���j6i� ;1O�E v�)8��A:����IZoH�f��jm�F2����إ��*��k�@��E$
|�1~(�ǫ#]��K)�X�s(*�e�n�pm"�k}86�G�v�/��x�6r��@�c�{�v�>�J�0���u��r�)	�4iq�В���@���O`������f���e��B\w�6^�$���\�����e���i�Ft�ŉ.��Z��L�iS�fg��\w�D���$[y�y�����(�P_0*�	��������`*�vK��ıg�����J�*`R8�8u����B�ӟ�T����
}��W���g
�*����0��2E���p�L _գV%s����
���@�Ks��T�r
�s�u55N&}���W X�W/��u�(J�mNc�I�Dn����Q6y�S�s����e���n�˴���g��S?;tTo�A����!���h�����h�M��,��+��LYP}Dq�r��2�Y' �rm�{�6W�壄���kC���1!�����%y�����NO�M����	&�̫�	��I����5�o�L�(�r�0줤!������߫n7iR��β8x�s�����fxI��,`o��7c�[ؖY$�~Ͷ������l�y�����1�m4�=� �~��Lax_�|��cf@�J�1�tE�Ҧ^g�Cx�s���2	W
���R��o�<�~�ㄵ��=����S`|W H��̴�Q^ ^���z���d[��z�S���2��-*�[���UJ9*���'�o��n:�R&�2�"�}d�\-�a�t�׍. _\�aO0@e��a`�a�,��(��ZD@���B5@�b��6����~����
���A�jG-j����y���S/����(��.�,���j	.��ƀ��5¥	�K� ;.<fj�b�<��:��nt$����w��{�� c��&.�7� ���	��BCX���D�&����f�3���=y^���'�iړҗ���Ή��`>�6'z�0ю-�b�&�l�i�K���}�{�'��L��ټ�q�lo����8���o��6������|���c�����Y�}�1.�N��c�4u��{���Nr ��p��E"q٫��E��,��e�Y�<m�I�c�w��I>�x��z��f�+��S��}`�cHJC1	�V8p0v��h޴	֑�$~�'� O�srՈ���o~Mk�k�ɧ�п���J��_����Q�Q�X}����7V@_�`倡�����Q�^��S��U@7G���Y�) \��JI�.rꕥb)˚�8F.��LIdHLK1PwGʷ�����p�(�s��9�����������ԶZp�m���{pX�Z�ɟ7ի���c��_�Ϫ���4u���? )R�2 N;����
�� ���#�����HjfefJB��F�!��8F1s�:�"�q{�<�Τ�ȗ�n&���F�Q<�Vb	y���$k�~�׌�����p8�FĿgoF�0�;&�H�>�P�X��Z�c����=ˎ��Xߛ���q�$]�iFr�� ��� 7�8��f>��Y���=��N2��@���s籾d�Q�������.i�}Ϝ[R3�Z҄7k�=B���+�x�@�}��i��-�d{�'�9�;Lk��}�yƥ����ݬ;���4��e��ΟN޳��v���a�c���#��K��8i��s�ۮӞ�{�>�=N�x����mE���v^m�c��ڟO[�ǟ���ѾOM�)g��7�)a
[�ý��G�q	 ]� ?�IL�saG�es��-�d����PVư�'�+f���U`�e�B���V��/Wis����Q��P@�MR5M
T }B|�XljC�t=���m{T�{�Q 6�@d�XP�7�~fձ2�/�)�Q���|l$ҡ�ZZm��!�\�>�R��[���7`o���P��0�N{��i�. o�o���s��v�� ���<
����5�b�R]��e��(�#Յ�W�8#pȯplL(uP����bc�a�4�.�u%G�4Z�ķ9�ƌ�3�v���l��u��"�04f�7S<S	{����ӟ�����1�o��{���Jb�!O@q�r^�L�`N�q qh���t������$oƤ�����糶iǜ�6m�;+0�֟�$ug� <H�}I�̓�O��֧I�K��i�g|l���,-��Jo68�����"ʤ�ФEפ��̟�]��eҳ?�X�iI�7�_��&�7	�ƷMZ�7;{���*.9f/���	������Ç�������>����ָ@ى�RL��.��Mn0� Y�Td����J��}��W�������_��^�xAǍ�n����}%��@-�'4��4k��(Ǡ�'02m����O�Jg���@k�1����'$�{.�W`W���N@/1������W�k�{����GYdh���S�-��f(WD��{t�ܯ�2.#<�L]��nݼ�����ѱ@i$J?�s(aW9����%o��t�Cc�7���̾��V��'淓�>y�*Q����ɏ���O3P0# &?���Y�zz��%���0����'y!��Ib�_0�Fx|�>�R����bVpj��a��4y���6�^�ƭ�D2	L���@{�睔�B��i���f�����4�j��4!O:73��88��0�}'����d܋z�vڸ��Ljvf}|Iz�籇�5<ů�9椅���$[uU���j�S�g:�,������q6t�ko�c/nsp,SL�A�D^�_�����O�\px1�È�+��v%�7jz�l�h1bx:g�Ǡ<z���K��oY�����C�����I��a����R, ����r�n���v������^ѴI
D�XA������/��k@~��	� �XՀ������3V$sC'-�h�:����$Dd��w_���В@�q��wi<�z1V
76�X)H��6Z.R����=�o'�i�������K#�$/¤#9c�m >Jd�]KZQ�Ș^f�����&��#[���0`0+Ú��&������:��7i�@F��0#�4�}���:u�ͮ{�g$�p�f��YYY�NeUm3rd���T��wtNy�CC��Z�S��� ��;�Z���Ҕ�W4ֱ<s�up����i��W���� �T����@j*ι��"Q������O�����ߩ����#��N�:�﷞{�r����:�A���� ����ܽ�eW9X��������3Kp����*蹁��8����	�C�@�غ�����wf���ƍ����l��p����t��M������Tu4� �8B������>�������w�ꫯ�=}���9���#�T㰊"�/΃sQ ���d�;5�f_q8�[���{ع�4Ad������7 �F	�#"��*����c=[���.�����S�t7�8�?��V���jڋ,�I#E�lߊ�G>���@o�`pGP0�	��jog�*h�꧛��|��Їb�������E;:��W �t6E,����mP�G���g��ܻ�Z+O��jc������ޏFv�^5̱,�.?[e�Z�}�\�^�j�����i�t_6��u�o������ɟ�#M��f^8=�l�3y���k���T�[�Tn|F�\���q��j?���fi��|�Jt�O��)�������c��G�O�aA����>��s�V��`�
�?�?�0}��g��m����P!�
?�����G��� �aA@E���ۏ~����
�;�����wN���iZ����Ժ/��YY:~�.���E,(�`��-�Z� ���_!��t�<]^<����9+��Z."+G�`�ʺΩ�\�[���OY\.��- ݋?f��;/W7���}7��|% '���ŮԀ��Z�"�e�Ҡ�o8g���D�n+�9��k`�_�D�UA�v>d�%��v,Ut/���\�y];�}҈w���S�I���Ȉ b
,�""����{}*�����]���b�6�*NA�H�2����i>Z?;X=�D�oՃ �N-fu�mW�����0�)��^ePAO�O�~�/+ā1���Z�.���Au{N?8�,>�}r�,7�{��Hg�;�vV����o,�'�|RNH{/��W�w���4/\LYui�j�.����(���3�	+���3���͛�����/�H_~�e��[,l�>���������y�o{���6�B=�����Pf������f'��kb�,�_�����ں���GM���(���/<��3te���~S�d��I�RA�x�b�:���5��\��`�\󠯵��6+6�L	� k҆�1v��7vo�\�z��.K醭�Ry~Ӆ�״Ɲ����ꨌ#P;݀��hHZ��sd�5�ٞ�hc�";Յ4�إ}��\Yw�VQg�� ܾ��9vt� �V}꽨ʠ�*C+�������A�1��2�]h�8��#�����Z�+Df���EWQ�坂�j��~�����i�E��ϖ���(>]�"��h*�ֵX�V�*-�!"��Vy��Ӟ�;��#�$���ծc�S�����y��M��e���(߸� ���A]4�Uq1e�C�0K^>���y��}�][x������G�������J~<�;��|�����M�� �����-�۫����Q|?H��������/��7��Iw�|c�2c��G}������@�u���ʎ< ��Uq(��$x6w�>�9���5��t��=���3�Vl�W�y Da��͙����`[J�)ʻq׆����N� /��wsH�Ik�7S���ZBCx4zX����4 ����W�Uw՘R���k̏�9�]�K�4�n��tp�%�m�J�Vd����0��)���a��]@��:h�	����n~�En�o�t��f��س^_�sżDC��^��H�蟆p
��ȴ�H_Bk������t����=2��H�i�]�vd,E�Mɋ�i0�CA��Jwhǿ˅���s] O+�g�WN�Z"��bJ�:�ء#?1>؃E��:jj�����4}�8%�q�~s�����,�Ye����
�9~�S�Ҟxd*g,�M�c�KM�_��I�G�)���:�秘�h�Z���A��e�uFu�Kȇڝ�-�Ծ�Y�M��2��{��A���6�>��+.�k-��G��M�b�vT��=�S�U�R�������t�q����)X\�+���B4�K��7�_.�����t�ܼ8U�W�_���+�1Q`W�Te8�ʁ�o��c|��O����u�}�v�w�~����}�`o��p����-�%fg	�:��z���k+�q�tXWت,�V�W���;�Y��c�ӕ-ƺN���Y:6�"E��Fx��]��h �Gy`�W���9fX��:If��P������-J7�׳�M�) �ym������L
W�N)��%a�>�rm�,� �{�-��b,�Рx��{^d���?�QY����w�Q;.��o���1GC?wMC�c�=>[e���o��(�-��|�lk�.@;i>�Se�y�
1mv�젔��~�
vcz��4t�ӪZ�liXJ}nPȠ E˩��iԩ>"�!�x��\}qU@Pn�i\��V��\��X����'�P�5���T�l��T���-���2���^��K��p��}�ՠ2�ԶLNBih�7�O���q�Ͽ�z�N(O�R���h��>�Yu�*��`x�zl?Q_"��w V>t��D��q� ���.�,�.?`u��ꭷ~i.�׆���V3�C�j�~ܮ�w��+�ʌq��ƛ��7߲
���>M�O�ͽ���[�o�<������ݻ�?~�.����	���o��b���l� *~��;l��./z�_a۲_JGF�����{<Z�_<Q�˲ʍ>������s�]AZ2�w.E��3��E�ݭXɿ贽��rC�,Ė�,���\+���)�<���+�O�9��j�d����]^sI��d yZ^��n�"�����6o��\��N��::֎F��>�v�1vļ?��$��c�,M�V��Q :�&�{�&��<E㫀����N���2
�y��
-�H��\�}'���2��_������r|U�-0�u����v,�N���*T~+�]:+etT���e�}�Qeu(SơAY�Ȍr��WtS��|\DC���@.�udZY'd`U6
����<��#��gl]F�= @D��
o@���ơuC9�y0t���C��!Ρm,͖lR&�S�j�³�n�e �B��vzz����5�y%&�R�ˍB˯��u@mtdo�-g{�s,��6c���uO=S{ua��r�0���a��Й��=g>�>�?[�R��,ʤ�	����y�Z���mn��F��[�������_���� �8��Jv0��vT"*{��n�ӟ�dۘ�<zlG�B	�_<O�?��ӳSk�ggO�Shэ�]ga�1J}�?sn���9�/~\�P��y��V��n���j����[�uӻ�Eh�s��B&�J7~du������}�� lW[e�iD
	L�Vp�c�Ū{@I���Ə9��@|$o;2��!d���ti����U��j|]�W,(s�m��\�R˲����v�rJ� g��<;e�t�3�W�EP�� �*����6P2�|c'V=��^v��1��R�f��+#�b� �W��4��Ҩ�Y��)P��+;@���vE��l��m͟og8Ls4D H��@S��%��Θ@��+�!��"�~oz}j����N�@�ӧO�3\C'�m_�8H�V]Nչʙ���4�4(��u�&����~����9�r�gŽ�;���e���hzz�m_1Y:���T�req�C�M#\G�pɣ�r��d��`��Yd� \��)��{��P6�CP�a���� �8m)e>�6"��י���E�Bu-���k�2��������N�@�z4x[̳kʆ��
�
�.	����\�8 [��sG�6�N��D��يX���+���Jo��c:F����/�oo����y���z�z��c�] ^�s�NN�\> Y�s���1��׿� �I="�yϞ�����
!��O%�cg3��3@�M]��TS���*@��Q���=g	��e9��@�����iEŔ��G�U5;/�)yvpF0��a��V�yr_�Vm�3ɞok@�0q�=�&-W�m�z��H-��e5�tv_��eNs�l0�A �A�����رE���v��Q:��ҍ?2�,���S�S��w__q���T;RvR-��w�L�u�4�>N�Ȍ��Oc���u��P����a�Ȅ逅��G���,��S�V=ЯL�bޙf��"[;2'�+ ����DTQ�
"�W�yf�g#��_�G�La�n�T�~�d�#+�+P^l�81� ���;y�0�=�'2g�i1�q��N�b�(���ې/�>�3����A$e���X_h)��/�e��NԾ ��8`�A(�x`�u��lk �~+�AZ��"�A���*$���?u�����������9X�5�����	�ST��>\��S]����@�����e���C��ε��s���Up��Ƙ���G?���o~�~�k��M�9P�(JW���]^���b�������V����ѣG�ᣇ���.=x� �ЃfN��A�%нmk�������񾾟��5��ȷ;Լw��.�rn
�8aeM�
�sa�	�F`�+~I٧�.�| ~�.S��|����m`*�=��G�GuJ��N�;�Fo�;��ܨ��Q���_�T�!�DJ��e]_����1 eV�ߠ��6JCI��Ni]�? �z�[����Ѕ�G���%o�ԕ��q�'�,݃��"�9�o|4�v�|׎�.��S��P?{n���љ�9tH'n�ӧE��b�b�t�v�Z��Qp�;vD����X�|/���g��JV�'��%;�V �~p��ɯ|���w��!ʕ�P�]� �!�#Ǚ-��� ��� ��Q�z�����s��E!�$�!�Sk @�A��6� ��������I�f{c���Du)�ؔy�'s�%�����Պ!R8p'[�Вaܶ�Z�$��TeO| C0��#��ղ�͕Q��x���mg.����ʂ`i� �e��#��}��#�Jw ����Z\�	�q-��*A���_�@���	�V�c;�ߙg�~��ܶgfI|劫���SvBP���+wi�
^F�կ�,+s��Z����DVX�� ^;�bÅ�u���8�C����޿?ݽ�m���>|h����g/��F9	$�[\L��3ծ�ŀ��Ֆ��p*q�D�_����7;�˵��LA9W�Hf|�[Gv-����L�Nf�y,W���{B�80���G�GŐ�S�C<��g����Mq�H�psF������M&�'�U\,��yV���������
;����72���u:?�^��?�I/�I�6�ݨF�`L�7o�\;�͈��s*�: vC�l��:F��'�՝(T S�r�ME-�yU�a�y��i��S�`_ k֟&����J�:}�����:5�S����T}iFJ��6�U�����2�:���\�tZ���f�����N�)R*�(��:x�z�vY�E��,�#��(jv�H�g,��.�Im?���.b~�i���6���T>�]�w\7��({�s�g�h��NA4�P�ѥ���aУ����?_�����6�:���,^�� ����꠼�u"�8�-#�:�ʟ�1$�vm��&F�i�kx��!�Zզ�ښ�7F,�bL}v>�L&Y?/��pa �޽�v�ۭ[��c��O�lW�nv���?��.�؍#f�C>5�##90(����KCN�Mé>� ��2��3
�܁aޫ�2��X!�0�2��5/�΂�1�#���/�����҅@Y+�M7�6�� ܋FG�������([���n.�"����.̉��(͆�k�%9�������Ӌ���yv��2C1O���ےg̣��*o�e\ˉ2����l�|�gB뾲��=?�j�sajs�8^��y���u�A+�Y���s��GƗ����b����n
@C�`l�[϶�I�C�_nT���7�}ߍ!�L��"�h�f"���n�v�s4 ���2�#��׬p�`�/�Ǽ���1�?٥���}7    IEND�B`�PK
     #{dZ
��
  
  /   images/edf2d60f-7dc2-4972-a04c-2a93629ecddc.png�PNG

   IHDR   d   \   ���  0�iCCPICC Profile  x��||eE���6�ѫt�q�"�����ٰD�ݐd�b	!v��X@��)�p��)"ME��   �4AiR��=sg��E?����d�y�3��)�s$���?��j�̙�p�{���{�U]�d4�[?�l�?�`~KWWG������K���f+���Yo����$iX�_10�����K.�O��ĳ���~��a,�;D�t��ONo�xz�[A��[m��L��}��[�x�$Y�<M���>����4����93f$�j�H2s��9C���1�.�}n��9za���$Y<{�u�s�A���M
<�t�_��˴.&2�[���5����jG���3�l�4I�4m��t`���j�)�r~SgSOSvP��Ń�v��d��ɊdZҕ�D$~wK��S������Ġ�#iM&�u�df2����p2�$�$MhW�L�_F�ׁdF2'��YR�/�k��Չ��r�\�qc�m�ޛ��Y8x�Bzm�7����Y�-д�j�܁ZIOB��ۜ��yN��DlKH/����m0���GIrŃI���m�N�5�I��� ��)�J������}��c�Ӓ��ɵ�m�ɓɫ��6l� vmا�І3�mx��Qk��FMuب�F=1�2z���^6��1��sƘ'�n6v��+��s�wԸV�x��+�v�MV^��C�LX�;�<Va��+�:c�?�ֹ�]���~�z����r�s�Zk��������:��;n�3��r����^����F_�jö��с�������M��l��n���U[��|��ÿ�:~��p֖[m��k[_���_���/l{IӬ�k�����_�{��؅�$q������M���]�W�o���v<p�c�vf�eom}t�?v^y򖻴�~��]�w����ԍ�Zw[�}i����O���5{��k�7.��ߞ�w��o���i3�ۗ�<r���5�?<�ws7�w����w^p�	��?h�%KY��Ӿ��a�������1�;������=i��ǝr�i��?�QgN8���{�J�-����w~r��=?]o��^y��W������_��uO]���ˡ_�r�6��~�;�y�λ����;�������#��x�����#�y�u�������ze��w}m�7&������/�k��O|�����+r��FCF�+�(�����Q�:b��g�d���؃ǭ7�ƕ�]���˫�\9w��W;b�#�8nͥk]����ܾ���y��6�xõ6�������N���[�_}�1���7Mh�r�V3�^���_>{�˚nn����W^H��>�be��Z_ob����m��l��v�y�������#'��z��������/������i���mʜ�'t]�۽ݯ��<m���>k�c���^���#�|�[+���{�����2�7c���}���Y��p����z��s���7�2��M6-�~��u�В%w�Y�.��M߽�g��U��-����=��uܢ���N�����W�|�)�8��Ӯ:�򥗞�������:��������?���;���pя�d��.>���?��l��_:�/_���+>����>���+׬{���m�y}�7�~S�/�n^�Co9�֓o;��K��׿��]�}�Χ��]o���=����^������c>��}���[��џ�q�c<��'N��O.xj����������-����0���/�~y��Vze�W��{�ͯ����7�\�֩����;�y��O�����}�ׇ��G���s+Ƹ�8�w��7��t�1��=4��13Ǽ9��q���c��+o��?W���|�3V;q��8}�ֺb�׹g���{q���0z��7�z�6�}�6;i��[�Q}�o}i���&4m��VS��{��_>|�S�~����-_�7}<{�����Vz%��]s������� wl�i�׾�2o�᭧N�q�5;�v�<��ή��/v~uJ���]'�vY��=/M3}����{�C�Z��+���o���o�=��}��������h��Cg�w���Ͼ{�Ss_������¶E�/�u����伃�:�C����}��U���HvT�ѻ3�{{�q���/=��o9��<r�ӧ<w��t��K_?��}�g�w���|���������.���+.�/I.���-���?\z�e�_~�G_y�U��섟�v���\t�����;���Gn|�g������۷|p[��;���f���ٝ;����޻�}��{g�7�������z谇������)<�������)����=�����f�_v}v�粿6>��c_x�����ˏ���Wn{����������eo,󊷮���8�����{o�k�k8���Ώg|BH�#�Q�Zä��>����G�ї�i�_{Ӹ�ƽ���+O_e�U^��n�+W�`���8g�׺t�k׹m���{j��o�𕍧l2ӥ�ݴ�3��_ܪq�/�;��	�my�Vm��6o�^Ӷ�k�e����Dv6�D\-oU��G�3�o۽�����q�N�k-3&�z����~��&��>���j:v�\2�GSo�z�{tτ�I�����{�f���Z��M�%�=�o�އ������xp��}���¬7�>��ٛ�i��㼮��0|Ă��-������A���Ρ㿣�����_|�)G.?���?�c�[����'���y�?8y�)�N=�CO�����8�ǜy�Yǝ}�9���sO>��ϼ���~r�E�_|�%�������K{��.?��<�#~v�Ϗ���kN����~�ˮ����n����~y�����<s��r�w������ѿwW����Y��U�w������s����`����������cW?~�����'�j��'���g��ˑ��ܑ=���^�ދ'�t�����W��ο?������k���[;������9�ݥ�-�׍����?|�߯|�������@��,/NH�I|ŊǮZ�b�����iW��+V�~`Ұ��R���k�L�R�H`�k��$[�̱Z�Ks����#u��xS���������k���^�������ֹw����%�������������8-I�w/3������u=���������x�ۿ?���D�̞l�����񊜡�!�*n�Ff�����+x�G�����D���W���������M��Fo�����������oC��*_��'���c��㎡�m�W��#g �N��޷S��a�! �~ �%��C����x�-��|��_ �y	�v7����x��k�"�|�x٘.;�LaAB���}�A�U�����߭+Aֱ4�m!�'�,P3��T�jK�$�����o��Ѝ�7"����T>ukjA>���AYƀ[ǀ�	��ݴ��P7�N7W/z� �b��!�)U���a��&��u6~���EX����,w�����\Ɠ˰i�
�>w%Mu2hQ�IԞ�m2�N�Q���c���\��bȌdD��q���C�&���Az���>$d����fh�Z�b'�E�t|
�RY�,��b��O�!�/��Mg�5��d�!e�l4�W�1�� �L��6n������>��m�b��;��bNV䝽�Z�V*��zZ�ۻz�vW[�g.�=���?{h����C��V{��g.���^X����9�xcejw���)-#��Z0x�Fc������mR���a��I��jf��j;�\u�SOoom�k�h��6Nj���hٳ���>erG[ߤ�ξ�޶.�Ib���]}����,�0@紎��:Ǝ��}�m]�������+�-ݓ�z�ڧ��vO�l��[mܣ�{h�`u(�Ng�/���Tm�7{�p碹��f�2_W_�]mw�]��S�~�/[z��ڱ߬�'���������ґw��	�M�α���I���hEMe�1i�ښ��������)e�i�L�����ѾWۤ�ީ}{�eiZmܳ���2�}R�Ծ�i�}�`�����>uJ_�Ԟ���m��2�'�1����uuOݙ��T�W��Um��6�b���$Q���,Ψ8�pV�������ϝQ�O�����jY�5V�;q�#Bkc�mʤҹ+S'��uOo��d�g}8�i��Ď��]��vȏνmJ�ە�̧���ٺ?�����K;Χo"k�����H��،���:�w�L]-�������6��Rm�����	��p��k�,�"�L��9���ٹ��cROU{Oj�m�ۙN�������ᔂ4���;���j�}{��t���4���9z�z{���#�d��?%���Lh.G��ִ��Jصt�iըZ��U�j���W�qaRU����������-h+#2�87D�T�cV����,즾�����j\+�8��S����L?�_�j�Y�������L�BTL�^}?Jf�?���p�I	�RS�q������LrN{QZ
ڨU
-�,-�XlY�τ��b!��V,R�u%�1�h�Q��`�6�,
�hS�F�L!����j
�\WEZӜa�d\a��D�bG]��JM#XeRZ^��,CGQvv�cVK3EJ�3Йb�*jFI��d��-8i3F��3�i;5(�Q����c,/LM&!U�Pf��5��iU�t�q��5h���	��KuZ���Ը}��:C=3��A��8G��X�)���`�M�dL3��2RfF�5���� 7\;�2uSK!�
�35�SЩ'�-��Ȥa��4�%e������[2�:lR����T+R,����QA	6��rM�8�-�Z2^��u�F��D>CrM�� 1h��+g
[3���� ��c���`�����
�B�aԤN��1i�5 ��5%l�!U,�����f+I�pY:UV��d� ��դ"��<�F��0���T�=B���!j eR
,�F���{��	3]�������p�#�f�/��4�?��i	��df�r�Ff�C�Х,�±l�ќvTG��ʔa�s�⢟
|&�8f�_G�-�8(!�+Ν|N���T��e�Y��zAI2C�%�R`���Ra��L�YO�-�Q"�����5�
WUnk�~눌<#����-�#���hF4^[=Aڮ���;���a*�
�:I3�	�1��f8Ha��PcɡV�hI3�	�K�`���5Bࡄ���i��S�:l�,Y!]8)r�&K`CV�s ���s�!pv�,*�Q��u�%�D�Z���
SB� �Pl\B�©t3Q#~(+2����QT%ie%Ep�����#l� ���@�G����d�ď�
S��}�r*BQ���� ?����/��
D��f�m��%�zA*�?ً�[��2�ѐ�!$�D�u�WLs��-Ij�S�Ȁ"J�&ͬ'`&������	ieRWpFJհ�����B
���l5i#l<p�?1��#�o����#����J�T�RS#��'�/�LeU@&�P)��
�X�!�:�� %�����" �
��Vb��� ݳ^B˥d�8)X�X�65��I��Z�YA�pv��*�d`I3�	I�FXNQܲ$I2��U�b��.K@�*��ȰT�9 "+�T� PJ�u��̀���t.�L@�K���@�Ҵ� ~�9Mr6\~�5��+
lp,����G��'��%���� T`+*�Z$�4��Ф��$.�ȫN&�*
8�#I��	,����}ુȰTdZ�Ì�� ?L¸�[) ɐ��3�(�a�A�ip��H��V*��
�#�z�iد%���� ��R%YCLt ��}	EH�KX&tWQ�$k�Px�	��cA$�L� �Z+S�5�X��d}�!��H�*ʖd:1��=5h�C�ʓA�,@�%�Nё�$�iF����y�`����#V��ɴK�$TkNY�.�X�~U����q 萉#��h>"w���d��"�rJt	�Z�{t��.;"u�jO���T���D�O��FV *�O�dn�#r����B3 �G�)�"'�$@��1%P��3P�! Q�?2�
��"[�O��Td��$�p\;�H��c}G�Gxأ�Saj�'�*f�
�;J�� ����<��Y��)���s��C��!�#(�A��p
����O�FA��%4(��T^�0Q\p��ymyJ��@3:�C��ʃEǌJ#�H�3\��#K&�*�C@�@y
'գ���Q%G���8��)
�K)��UȺ��z��@|��$G�]�隴X�)�c�9���@M�;�D�bl����J�Q����ݒ�N��z�Y� �ȝ�)Յ!��jt�J:�s����z���\�=��
�s��-�ʪ�u��u�Ɋ�%^.
P�Ȑ��@��lV�����U��H��p`V�e��`;Bs��3𫄨1�#"2Uѡz�bUIǸTJ�p�*��%�B�.t�.q�# KE6�(S�(1
et��=FM  Cu�ѐ�QF�� [��������n�j���e%�h0TEN�(��D���YIϸXDRE�<E��Ty�2����ĵ~j����"��k�	�"ѓ��֨p����V����'���)J�kTጂ]jɹ"=�m���ziY�X�pv��:HB�O����/z�Ց��= ���L&$t=!��,�$ǝ+J��{��JW�A��4z�Ւ����A5U�Ȋ�@�&c�Z[u�j)m��RJx/�\�&�^�J���*c!�z��)8i�s�ΩgY=9�$l�l��-vEO�"}EOV 
M  `p�)6ygh>�-z���j+�"3C5-J���P(z�2�)$������2����Kَ�)��D��IO�!������J:DM���<�㔩�yq����Kf�'�������sB�M�`�TV���q�"Gٔfg
��z
Esڒ��3�T�D�<��D��R ?��`$0�����)�d1h�N�e%S��*,H�!6F�KE��6c��kF�T�@Z��3m�꧌j�+{*WA�/��d^su� z��DI�HP�x�rZ��1��P��)K�fܧ��=�)��`C����S�xͨ	�,,%�ZP��8�%b��kF��� ٰ!�jh�=��)��EO�dT�F��~��
�=m�׌�`d\t����J�����4��;�g9���&ݠ}����9���ST��T�E\��8J���x���	R�j���S�'��9/S�BT�4Uށ°>R8z��#1Q�M��(
�ҡ0��)��%̦BO��ω?!9���f���D��y�25S	JNp��r놀!���􌫥�/H�!g�l��	��l���bOh_��+#��1�>�p�Ӗ�٢'e�F�����&+5�)�\^<a�G�r�)�t��bN����B�|J'��\O�Y�����s����X��R���ckj�ag*�իk\-�a]���UޓM�)�R�ؓ1`	R`� �zJ,=W-�ᣭ�5j���r����!z�ꨆ�
�p�`�[)Be���%X3�>� �E=�`���`�4�)��Ien�/�)'�����ߎ�'��ͫ�����!+ˌ+j�)yj�|�C*�a��J�m���TIz��ω4.����gA(�@�
HA>�#�R·��������2ʧ�����e��%���IQ$Ж�
�T?�{ҩ�2L=b���)3�a�4�O�VA�S���gr����N�V�9%e:���}ҜY^z���&<<�����ƞT����fd����5aj9�Tߓ\@�Οsz�F=���Ti�X\&�G#�D�
�)��bX�*��Q�T�2Iq��f���W@ϲK�'qV���3��Sv�S�d���&H���R�$Rh�%�6J��1�v@1�H��(Y"� 41�Y3�Tf�ժ����֖�c�t�$us
�;(]���������ra�R��0K�4e�o�& `���=w������Cʖ��B2*�K�J@�6�Q,�e:��u�A��(_&]Od����C�=�~�Ƣɭ�T�9�aا���~�Cܧ!�F^�Bu��~�qBR#���=�$�2�xi�+�SOBoZ�c�'��8�JC�:z
zʃ���o�������2Y\���M�ϻ;ip���৮��,�_8��v����V?{e�ذ�pe�U��Sm^��4���Xm�	g]m�7#z���fd���.�[m�"(k�A���DS�=m��F�"a�yZH_׬y�Ϛ7ܷs����K�������4V���y��S�,�$)J.I�u������:$����AqG���#/�3.")�P�D��I�+%���N��4���s���
G�	N�@{T�s�tBrOr�kQ�J1����s^ʋdn~�����
�bD�Vѣ=ת�ԅ'��V���xΖjp�j`&6_��*��Z������"���ka'Y�*nf�"�"0:��VpOJ@��D���/-!�[9���9��y^F����[%�Q �bgN���
Z���I���\Ⓔ�`)���)=�w�6�.<���� :�|\I7Y�٠T�I	[�I��+�N�X����ړ8,��"E�o|7x���D�|�*?�j���y��X$j�K?���ڦ�T ��lVӅ�ub�7D7И�$���f<�p�p�g�y23~9\J!�s��µ
�$�=��S�R�x�SʜA�p2�d"��#1i.������nk��ʲ|\K��/�.�z��T�oSЅ��
�ΜB���B+s�c���ɒWZ��߬ĺI�s^����z�/!g�w���*I7hB7�p��(�V�a�He��F��ש�k�0]�y��m>?�N��4s�3��k	F���.ʵ���y��qG���V!1H���ޜ��W9���Q+F�{iSF`,�y/Xn0^x������x9�/�ca��=���n�:�vG�cR��0׹�g�:�
Я }���0t�����$l"�֑����l�6��e��4��5S�,r7��Z�7D�L�)�dΫ�a$>�d*�'�]�mf-B��L�3�M��.=��/c�K�&+H�ϋ��x^�_�r�&����l7'�<�t�U'j��f���%��$+t{>��M3o��OrxaO^f��r��d e�I��k�BԊ���$�?OJr0�7Y��t�/Ge��h�yU~+��;Ox�б�e� �I��#@��ņ�lP�p�Z��D������o5�ҁ޺q �Q:^2/�?A'�����ij�>��0A�#��:��n;�1m:'S�f�(����"g�	��Xa�] ��q�EC��	`�	�؏_o�����If�m"�k���aTު�WO($}�$'�.��-��3���������8�u�3H�K�B��a�o���/���ɃLM�g,wQ��4~�Ț�' �q�g�P��R+�R�Y|B ò�/����@�ԏ���U2���LN"��2�!L�j�w S�!�x�͡�k� ���]�yE^|u��e�daoPz�=�.>��$P���nd����=����l` 8�,�Fn���G�v2���x^�q�IN7��@��|�:����d�ې->g��'�I��Har��a-�Rxs�Vi<o�a�+�d�H���[`�z��-H�M����c136gl�'�"����[��`-�����#�!P��=��x�����_$���Ъ����pd_ގ![�Bk��"���iV�<dV�E�0�
�ړByA��>�GC2l��ܜ�{��E�s8�c؈ិ�0��O���!����GC��k���M
?n�04��K�PoZ����f��H*>y��`�ګ'��29�,�y���/eY�J!9%�~o�P�	�H��i��e�-0�A�0�)��4��F���JA$���Y�0T^���#��~�Aw"��,�E"S������p�I�V@�A�HLe�-0�x#�=�@�H��+"��4�_����$�3������37)������r��P����W��7b,�y�J��.�n ��[`�6`9څ�d�������i*����,ƍ:���d:�Zd1|�����0BF��y#�A�-����@���SD!)�*(y�D�`��FP����@*�㱈F�-9�)����*�Ǎ�4�)��$f���>�C]�����y���)�T��h�~����j�L鲤�!1�T��k�8)a��"���y���. �O�мJ*��]H���-0����"􄳠����-0��"����SD#�"���ҝQ��"bZNx��J��""��r���R7�������z'&`!AS��z#��r���	��� #��/���,N�
=��~��s�Ҳ�MK�d�0���Cf�WK*$�� #���jH�}�L�/�Kd�0���AKp���31ր�AjH:{�[`���*{B�r��R�0��a<�3_��HB
~op�*�@�e<o�a$��F�,'1���X1i�L)
^���[`L�y�	Rz�̥����'Œ�����,"��x�R���I�"����t ���T���LF#I~i<��`,�C�0p�<,�"��Y�k��;��6Hﱲ�Fҧ�M ����RF#��&�Oh�$}3�?��a�jø��ae��?n�0ha\"�{�#���g2b���1-H�nR�5D�V�C7(�_}���E�0�B� �����qHE#)��k�\�Ӵ�ۙ�-0��)�@�l^�r��Ak_@%!�c�`�*bEϗ�'e��L�����n�R�|�PT�����0h�60���E�M��ME�V�����+�:��-0��}�I�;�4��51�b�� ��5D覥�U��a��7��>��e�����>��ɂ�`��1�B���Kc{Ni��g*bzt��>e��L�:��F�"�*�~\A���Qݽ����Wi�㨈a�-~oT,���|�FQ�xeȥ������Q�� j>�(����,bE�H��sR�1��;�Y`>�S����(x#���>��ی۵>�@zg�7R�V�|#�Q�t�,I��cU�0вP��Y e�A��a �{U�wiC�JE�H�K��}8Pp+���#����>	�rU�>���t�0��B�V�sR��L�y��r�kH�L���mSGC�"�����ߟ��Fõ����z����!u�0:+�6�����I1�~H�z��`��T1��;<�Sa�_���#����T��9Ĝ����u�0�2_/!��S��a4� (*Vx����5D��t`0�q6Sޟ�a�ǽ�k,� ǥ��D���xՀ�Ɋ���"��{>��d*���U8ވa0��,Aѧu�?��a0����3�� ���[t�0�By��]�$=/�y#��)T�U��G�
�at�0`�M�&?��K�9o�0�"�IMR�:�,1��>k�;�wC��"��/T�PBC�܌�>���8P��k��	��� S�����G6��1�h���n��Ve|2àU���7_��{)a�à5�=M�DњW�+���*�ޢ�L��u�DC���Az������0�����k�`��M�0Ԛ^���'��x�DC��Гh�a���k��Z}�0t��OAy��Y�0����!p, ��#��a�+���+�7CUO���a�*}ܐ���5h1��ų�����F��̃S8
���{�4�CX/�C~
X��C&b0��y@=V����a�|B,Sa\j
&b�T�wW�N^�4��Fc���npaǀL���a�P(}8!���-0}����@�#$=��5&1���VNJ���31�=���N��!rx�c"�C(�������5G12;�i�1�p��ڲg���..J�ڕ���z��Ga����0`�a�t[=o�Y�-0�!ǔy�,�P=�l�7b��1 �I�5�וm�0��(/t��>I_��ㅍ(����R-�J����0H+C�e�{��l�.�y����=��Ґ��`�٢��RӰy�_}0���FC��s!�����6b�!�����	�[`K_n�7ρB�l��x�EC��}������Nů7b�d�+D���c���0�*�ab@5/_��?o���	�Dz�˼��xc�K7�
����'m�0��f �T�����:��o� MW���0���P��ǥo2��1���p�A|p<���gB7��AJ؈a���8����89����a��o���{:�H��F9o�a,=D����@��g��ۻh-��ņV�R�x�;I����Qť�   	pHYs  %  %IR$�   �eXIfII*     (           >       F   i�    N       %     %      �    �  �    �  ��    x       ASCII   Screenshot��W(  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:exif="http://ns.adobe.com/exif/1.0/">
         <exif:PixelYDimension>650</exif:PixelYDimension>
         <exif:PixelXDimension>700</exif:PixelXDimension>
         <exif:UserComment>Screenshot</exif:UserComment>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
��^  KpIDATx���`$ՙ'����R+gi��&g&�`f`6`c���:���mvo�|�ݳ���wo�^�6N��g^lLf"�09'M�F�,�:�c�}����[�+�H����ߗ^9:�9�OM���h�r	C�CH�R�����ۇ�8�o��}�0���-ͼ�cd�k���i��&�j�M>�]��9��U'�l��k~�O�����\O�k�tMn,��o��|E�tm�#�����{F�چz!��0�K#���3��z�����˙�����@MM<^/�w8&��	���_��۷al�~��NCQt�� ����ÛG���]��5i��z:�4��g��EMq���~h��L$ͅ1'&����ɵd��6��F�;d1Ҽ ���&��6	��2��9Blb^X������bw؉��Xm��A^�l6�M1�+������J&�^Zd>7�������щ����Ĝ9�q�M7c��[PRR��y������%v|��k�d�V����as��kN�9u����ؽ���S@��E�K�$Ȃ�\ē��f��1�,��ɹ�,�ɽ��x�ӡ;���j�bLs�Ԃ˵4�\W7R�Tr]�"�uE���՘s��?g"+�Q�`���%UY&�E�$��'�K\a��j��1#�>w
��ۍ�o-�G� �6m����H� />�S����/��l�m9�T�h�D)��[>�<[n�Ѐ���߾���9���]�d4Q_,5�0�Xv��,��t%	�[3�̉X���3�D����.�9�H���d].7�|��x�NYYb�	x�{�#C��K�D[����d$M-�R-��!D�����޳uj�����d2�PD��$&Q�u�����U�I:� �ڃ֖�8|h?��QYU/�$�Ӌ����.����P7��t�ۑ$�L!�� ��8Q��h"�!D&�q��&��ߟ����ibtcs]�1�zU\d�eG�M0LuBjA�2�9�A���ql޲	�|\�Ԃ��ZYh���&�s��y��Ҥ&�4�8��N&(,,DWw�Ҧ�sl��$1��j�-:�d5 ��J�L���ki�#m�K�$��|��n^�P�a8��9�7��$�u���'��cx�����������K��/��ȅ��W������!8i2�P��tÖ�
ޒX�t?���O�ɿ�����fr���t���LB�5}�X'������J+� �\VV���v���btt����t�4q�2��U�7��s)�#A6jdd�t}J�(�X6G8ߦM	ٱ����Ò�,��jJ1Y�16��`�D9�f���v�G �x�w�������_0�!���Eb"o����D��
���~�8�~�1��G��C�wC��/�-�4a��xk��]��d�L.Q�	X����g4����>�ٳ�a߾w0w�|�k8v� "�A��Ί�
R�q��.���7���Qt�t��ŋ	�N��yH2بA��P]Z���F���@$:NӉ!Rk�d#Y�Yc�K,&�%F�<�׺�K5+{i*i��H��&ڍ>���o` �O�������;��_�[N`|�f'&jg݅���P���a��ͧ_¬�r�\?��Fl�}D&�iYD�K���x<��~w߽���Ŧ[�ct�O>��	'�(�W�a�,^y�����)��P� h��PW]��[oF��"�T�p�d'I���X���T��$��O�Q^�KVލ��^�◿�_z3g6�g�>,vi�qN]�\���oY�C7W.��m
tD6�y4�Ĺs�q���p�Vcނ�4y]TI2��h9*떙5,��+��"���������tQ�j���3J��M;�k�
��y�QI���Kx�ӟ@�{{��A00��|?�z:qaf%._� C�WT��h�ҏg~�C��B@o�8�K�u�����[�s�"x�S����;ha��_E��
EP]U;�q��w������:�:��L�*���Ԩ�
:�P]]�J	�W����L�#Lz�a�ϒ�'�k��mҠ�j��{�,���pzJQ���+��#�N;�\�$�1���}�8$F(��Dd�1��74�Å�� �z-1A�����8?.��mIsk'a Uc�����#�����:��膗��H䬠,��4�H$b�f-���J�tD��v�0����-�E�G3#��Rn�n�:!A���:<n�ǎ<�܊OZϼ@Wp��l2!������W����Ul-�AS�\o;�w,�ªU��r�r�ܱ��Cx�?�3��**�De���[h����+A̜u#9�!�L]�*���sq�-˱d�BLL����o(���h8�C�N�h��V��A�L"�7�>��ȑ�ػo>t����=U*r	��%�d�"�\0�/�6�	�:�Y���Sذ8�D�P4�q����w12�����ĭ�����&���ߟ�w3�%C�����7��J��mDqQ�b�{	>�n��ل���c:!�nRA���F�~�e	��4�@�w�t��*"�� !L*.AYV��}��@a�,\<��8ّ��Z@�t*�O%�tG.�2��$_e�5��C�/�P�aE,�|�����w���]�ÈzI�c�����_e³�*�O�Ot��"8pa��H܅��Q�rj*䝊������8�w�yC�Ы��Nj+���z��=@�W�@Of7�A�tn |IА��zaQ��qr�Zp��aBaaB.�!y��������Z�b����������t��#���E�rz�vZP<W�^�1�{��Z�B�|��[d�yΚMg���r������#J0���N�5֓7�Ep"4z	y�z��׋(� sRx�c��\$Q>�?v���a���~];�:���F��;ɉ�##Ev���#�Kk��R���+p�����"[�$�8	�������M^y�u�	&#��vkH���qňP6t�����h�1b��2^FXSQ�T��uV53�h�/���2F=߳T1�7���O>��O��y'&�#��Xei�H�=҆������+�N����b��$)N�l��%�����_�a�t�&%�_>�$-�ӮP��H���#��C=���ǏǬ�FBX�ţ��V��vm�=��;p��e���D;� �z��Q�M�a�\�O��W�`nZ�T҆I\]���v�/�ֻ���0~����Oz�$*,c*))��Z6�����v����p��?ooo����2r�*�o�j��ǅ��Z�O|b5]Ї�����o_%���:N�Ñ$�~��8^~�{���/(��cl�(�ÈE/���֑�� 
j���_ �֋_��=�!i���N�yb���B�j׮]N�źu����O^y!-�E�����a"؏�t	�z��9���/Boo/�`�|[YIH?�g{�PDv:u	���r9��jK��1��~۶��$�@?����0N��Z��M�D��tΙ;�-m�,Lco�1Ì{���b��
�$���]fА�'����
��ɠ��G?��\ ��y���0>r��8�4ҽ��p�}xo�.<���tCW�#�sP�uu"�0�ц���`<8������C�K����NR#&^�p1��G��K2&&h,�v	\:x�&��s!Mv$�b`p�W;$�=:2�c'��sr�e7�b��)��6SU�!iqn����P�7]JB�/���fϞI��6Iue��M싆����C�7_F������^I(4B��'q����:�}��C�����}7���L�0��5�/j ԓ@�8����@7~��[x��G1f�g����PW���96���-����90�z4�d���g?���v��ߍ��R����0��ٮ1a8ڛ"��H
1]d�=M0-�(��b缆A"3��_yo������\L8 Q�n3�ORTۢE��|��HQf���mZF�B�*�j'C�����,&IK�I�1��h�=����6r!�v��o�q��0��؀�K�ר�#JNZ2���S���n�/!K���19�x=d���G�0����!�qh�nۈ�[�������@ƻP��=���n�aU�&��ʵ�@3A�n9�~	Op�N*���넿�0d�%D�oKR,����$?h��Aǂ�q��R�y�8E/��0ӳ��Jq4�"#b�I\�A��k!�%W*�l`4���Q�>�N�q�O�	v���	R9)�h6�<���V��\�PUR���9�� �|��Y<�O��8�\�rK�.�A�D�%$˨���H^OR��#�>G�

$���3Fb�PPp?#�f��3��0�o�
�'�AFV�IZ�HZ*02 ��ǣ�2�ff"�����e��#�o�+@��p�EL(�Q0s0B�Y��P6�Y�|~���
��uDv��3��İB�417�yg-�9��,���8q�-�Z�G�$�oہ{?tFF���ì�F���C����w�d���YMr�����m���}dƓr�Y�:]�$��P�./J5�4-8Cq�̦�=+�H���EJ94'��k�ߏ�w��&(�㐳�1qXL�_�Ȝnd��rZL	��X�K�f'�9+Su-q����p�%L�Be�F_�(�L��	�e¹u�-��G�{r�����~���7�>'r��;$k��߹sפE��
I7�8�:5ne�f�6d�����PO{{!&|�X��E�b,�.'�M��5�̠�j")���FEE)i��ǒ������W���VY$:^az�Lr<%{a�+ޒY��o3��YHz�Mh�`(�Jf3r�ny�̱��r9S-�-ƶ�|wFcϿ�[,_���|B\~�<y�mZ��^���P��Y�f�Jp���^���qX���B������Z�q��[q�����q��y**+��9$!A��8��2BwCh�Y�H$JnD>-1�D}}#D�j���N̝[�ٳ�����}dd ���$!D�=z3���b26Q<��h?R�+l��ZYAY`ZT�ry����t�4��o���3�俖+-�D`s��	�lp.�9�L�4lww7~�_�D�صk��'jlx�-&\�O�y��on�BUU�^Y���O��k���m��� �#GN�ܙ�x������.�_7ِR|�����+��O|��{��z�en:߇�7�C���������^�}�߉#�.�5�h��:/a�ڛ���y	�\� �������Jd �8��A/w�Y���b�a��E���5��q�FDB	|�[?'(=(�C��M��b� >(��>����[�lC�(q܀H���ƥ��?g��?�D��y<��!K*��JJʈxݓ�g}����y4v��=� �i|�[ߐ��_����%u�J����Al޼�{ �h����g?{�Ф��ي�s]8x�(�)�{�)���W]�N\�($�އ�9�dÓf��2Y��,�S�.�<\�����cF�G��oE�LU~1H����AӬ�9sF<���z�ق����a�౰����&��!u^��\.�@K����R"V9��iS�X�$����?�.��@݌jtvt��|f�r� g*'�cƆG��?�����H��'�G�h�{����n�F?�+V,�|�),^܀��Z�msá8v�܆�!���?Üye����ի]p�#���5�9��c��b��NvfqĈ�>G��rf��c62RL/F,E�RC��v$Ȇd��"T0��+V-%|'O��²��<�WIB�$��!̝�`0[�d�_��R��+��~\ ��?�iU�U�VBJ�ÌQ�*�ͨCOwO6>e�S�f���O���䌆��o�#��+�7��}�qtgU�~�t^���?���/AN�Ȩ��_�+b�a	6zq�����A�`''I?)�"$ ��r|,���>�����G9qy��É6l=p���!�	rzbI�I�T��f�͸QR��T�,���EY�nz�chj�-P��|���4.�\�TBd�& ��eT2���*B�aOZ��d�lF6#��2�L(PB����8!&�D$&�U�TJ�LJU�����$I��#M�H�T5�=3
Ő8P�b��4!�	����_sd�$�Nc%��CM�l<���c��l���|bp�M��*���r0w�3���u+�z'�Þ��0�	��i9�5^���PJD�k�u���Y�N�����8~���L�^���{O�t���p��FI�E}�PJf�_��gאȟ �C6�����h�*a	ai��;f���Cd�����1�k�^�-�.$UG(��	�����мT.�w�V1�UY�?x�gx�嗰h�2ڵ⏰b_���!��e�4ѓ�f�Dpy����K���5�`s��G��@I,�����c"ƺ�+�.�J�XU�q���H��2x��(�f�d�H�'V��0�Ī���+��Sd�+��4����@}��uם�կ~��{\������^��3g���9,�w/a�|�7��u����<�0�Z�?wn�eZ�ڱ}����o�,���m�$�榛HuTc���8�YB�J�Tb.�eC�a�͸i91��!�^i1%R}ǒ@�s��̙��h���<���n��8������բ�j�o@��f���%NEj�S�y�Hdg�dW�!�2JJ��#�s�e������;�O����{QWX/F?J\�&�=}��Ս��b�݋oB��G��N/�#]; �ʕ�0J�*B��x�m������s]]��#�W;zq�|+V,[��{ޑ��3��͇�o�M:?�y�ˈ����{.����XI����s>3|qm6/א�"��X��E�I:WU�L���P�z/-�f���'��/G@!A,8���*��W͐��]��V�����I��N��C��*�kH;�hi�N�'������XNNWE599�	��� ɱ�@?nZ�s-Awp]��n�6'L(�G����	����I*�.���.4&����`�%Е����H��+��2�@�Q,��W�+~�@��?;�\Ur��EQ[C��Eg�^B`$���N�¯�#����|7FN#��% #&���a�5��,!��D�1��_�����]�/'bQ,XP�ϑc�Y�m��Ҋ@���Y�����f�Ό>��o��l�{oECX���aR�9��C=X��&T�G:2҉���d�ٹ#L�����mJ8�a1K}*e��w��w��a�������!O��"iR4M>�X�@u�W��P�t2����x<�D�r嫢i�I1�e�q`��1}6 �����52�^'W6��I��b��a���P�߆�p��G�Ϲ���eD���,�S����A�L#=Sa��)Ve��E(&���8d��Ԛ�}�0����N������jlUl�U��׹������?��Ж��D�hb�]�u\g4H^��`�������=�L��Η*qM�l�A���1�PP	,�O�p�^,��$m
���X�P+1���j��2��/2�_��X�);RNR�C��s PW�\�d$�0��8�E�<�p�i��.rR,0�%ml�t��\� U0�Qb���_;�\�"(�ID�G�P:�"�.p����j֠��y:� �� �\M�t�q���$�T_Gd��꓀���@��o��v2��K/���u���	�3�NVu��Y�U�f���T�f��r^��=*1����|�� R��p���g�����k��X:8o��jdt������Ғ2��ő7{,G�	�RbA'U� �>���|Mo�%����zc�ar�cXdɷ��"-^�EK�#m�Y5P���e�Fa�ȘyB�_4�}\&��`�K����a>�.Da�]�.��j�a���٥�)M����X��q���*�w��RU�R4f� �`��@�W���{�\�Iꍛ[�[z����5�O�n��cHɡ}+ϒ{���8VY,%Ʉ���0�FR"�\Ĝ���8*�cb��ǧ��Z/��/-) ��u_~��V�S�'ƛ	��+Bk[+:�Z%�$*��tY�xJ�)_ϦY*ʨ���� 8�2z��~$F�ə�c��#�9w1J�f���2�n,F%�=�W�2�+�a�d��$���/�"��%r(�f�N��lv�z�!ǃ!c�0.��<ې@�1:_�#��G�٪\�9K"��X���e^�"��jb�$oD�'	�y�4�;w^��e�ܸr-��f�_��☬����(!{�^7���] �l"$XPINq���ɴ��hX����J�W��N�6��[f����4��!*ʐr�1�Џ�U��8�=�"D*���)��bf�B�ߋ1L�1$�Tz7t|��O�#�@�q�9��A���%��5!�]��yaB���yiI1�ܾ�h��yWB|M��-�*�����%��O�p5i�
8?�^�׾��k��׾%���,^TE��I�O'IKf2���`x_�ei��p{%Eˈ��US7u�s�e��.���U��Ćڔ8H�T���A�)f��K���p�]w�C���H8��	�E�f��SEa������ả����8h	�I�EN+�=���6,GkG��G�t2KH"�,��-r@+�b�+�N�zP�z�;��q��'?���%������O~����&���ҪF1���@b��"*/�e�������0���4�X�~K��Y�nz&��;��Z*�;�l)d�Yl�ը��v��y'3CE|-+�@�u;�0/dhh���lP�3z\��)YCb?V�MT/r�#F�w�9��J���2D���,)�� U�����5��U�_�B[���������C��N��t���	��q��)|��-b�I���x�Vi--Y��e.U&�j��(D'*˚����K�ʱ�
j3�34�l�?�srr4p���vx�%1�:[�Ǫ�C	��Aѭ*o�����J�~F=�^mCy��x� �]�������N?\0�*:R���rZԸ$�	��<Y�	�*2޲�r�bG��X�c5��v{�	����uNr�
��$�áR�^A}w&�mFF���*JTنL�in���I4����d��Y� "D'�F4�֢��W�N#B���n�r��-�nSqs[�;�+� ����0,�F�9�N�q�[J���g��](ɩ�� �4e���v� ��z�r�m�P{A�G�𕗷�	�#�fj�mqI���z(.,�?��?L�j�����~��|O�eWx��13r:����@�",'עB�u�(//#�ߧT�Q��"�����RYJ9Y�#lw%�g�N��b��
qD�7@?���h46�B�U����Q�AUSM&T!�a#(=6gc��'?Iި�&��SO=M�	7spQ���''�G��dUU�,zeE���K�Jǁ�Wi�vz�W;�$���Ӊ?��{Bc,[�H|6��I9��h�4���� uKKJN�{8v�8�z�OE�b�>�-[nC�c���<l�r;�.Y�����P8H�GcË�g���E�rK��ԓmJ��DR�CW^:7!�Jα�p�]�M�L:�!2D\�M�$1�7�c�C��'q���ɿ(�q��k�GiC�p� -��-`R$������ڽ�֮G5������Ie�`ɒ�95BaM�z]Rm����_#��7�3g.��)�ಲb)H�yg�89�o�������;Հ��[�@�~x�1{R���^xY8��L8��)՗��ӎLft���%y����{'�ؗDl�@I~�L�C5qj�����b&1�@b�4Ӄ�6�I�(q"���8<���������
R=nr�����e̓�������|��R�#8F�GA��t�.�����U�b��eU5:Daa�3�
�p��E�����|�/�H�c,@yE����K-�V��^�d>��N�Z�W������K!g��+XI)���m�X�5����:<��+V���+��~,�z�ˁ�����"'"]ji�b=1���=eP� �6̨"I�G<�(o�87�~ȩ�R�R[����P�[��.�,]Kg�:��x�q������%���'22�)�pI�왍�=g!'q{�D�l6��D�Z>w������!� �6mB=-��[�pE����E8{�"9v�.d����iZ�jn[�����ā�~AH{��sN"IH�e�H�������Ce-���뎌�����.���^$UfH%<�_N"���	�0Zd�%0T&"'��&0��M������{as�g�pm$-K��������pf`>�ZU�������e���p�G�%�S��J?Z/������o�l.,��V�f_�@C�>�^�<��W_�f��VM`����NS�5�G3��%����AQ%E������K�-:Ht��Y2�Ip��
�WjY�=���_n�B�~����cpd^�W�>��F�qB���%��/K��&����;���,��Sc��O	�cO]��D�\c�PU#��p��F�<2qs`lLj�8�_�+�׽ع�E����1�C6�ɘ!=A��)�Ԥۭ���Κ5G�e6����ĩ�P�.����G&ŋ�A�����j��4��eX�&&��ă�(N�:���:R!~���L*��E��Q-��JK����:����4�TR;��~�2j4�Y(^�+�Wp��ed�����+a����@S}�\�@��ɪ�IPVC��u�RY��V@1�K�ݞ.���H��j�^<X�t*�
0>�.�����@1b�ʚ*��^8�)QWYg�P�' ��@$�~����8p� �ܼ�&�$�v�8��ç���8��n�$��2�������r�ƙM�;g.�}/9���a�=xo�ArRu�f��p�8��ܙH7w$��*X��a|��'�>�0��x$����������������6���I�$U�`� ��*?��.$��f1L�b	�li�;�Y�)d�WCU�H	�J>D�����W�������m�ް��Em�y��| 5u��ZՄ�t\~��M%`t��=y�%�:ttH�����j��J45�Ĺ��QJ����'��MX��<|����øk�f�#����� ��8Kq:1�&8`)�	Ҧ�4�1���>��T���s}��7bd,H�{J����,X(X:->�����@��NH/O���`p�.DHu�zF���	D9�;Z��ȸYJdneuP����M�T�1�:Cŀ<ı3�"�WKp؎p�<�#,^���G��S]B��Bb�H��f��uS$���zX��?�я4�7��Aeﮭ[1:6��g�����I��K(����T�>,[�R�u�z[�q]#.SH���ά�ؼy=�!cR����_>'�]q��_zƖX�����$����w0k�l"t'Ξ9/�q������j{;ټW���휉m;��i��Y[p�63�	l�8�X����+4�6-���h�څϪ=S��.-]*~2AY�y2Z�c�?g]
����م��qt�;���68�b(����r�7�*�fb�I'�K���-��]�8y����f��]g�4�t����dl4ǃ�#=�'�ғ�NMТ\�j?Vs���¹�W�p��1�-�ua��	SVX;��C&v�9�sO|E�\,!��i]]��(y�##R9J����5k7:F�����۞��(� �,���R�����a�s,�v0���JHN�2��؊a&ht�ȏ��F#](�oæʅ�u�΋���y�>��UIa.�ҟJ$9n�av�1�Ș��x���p;]KAB�r�T�C��zE�L��듽����{ț7�!�5���hP�V�Ъ���q�D�uU��b�t�(��9����w���QՅ%�YYY!D�9r��7#����>	����<U����vd���D�L`�}O���`��Ĳ�!j�<C�AZ�f��GA������PM*������dn�B�,��3�C�I�a1g�:]n����9���c��l�:G�_����`)M<4���W!Q ���6�.�׿�l��ےƺ<ϗ'F6�?��������.D�����e�~���%����z��W-���x�����[CMe	y�����O��5�Iu�4d$Ԭr�bqP���eZ2��d�����Y��L���D���g��:�3���8��A�٤�ϟ?�
�H2|^��pVHZ݇��&z����a��'/�Nr�l�镗ߒ� �pIk�s�1��\�
^H�F3i��I>���\ʹsV%�Q|�#OHΩ�'X|����%�S\�Ųe��VMH5�Ma�2���8|p�Tn�m����Gٹ�f��$X5z&������Gqd��3��P��6�u�I��s���6�#�+���a9B�j���p��G}D��N����	S5*i�"��,�Ҳ�̪�n��
�"�?�(y�V�/G���GU��%��f*�\��!�DL&2Ke$�R�T$M.�W5uV�ݎ��FQ�l��NN�i���5FMk#��89��$-FC��s��w�K��[y���Ծ���*n��x�e|���K�n�QU'����� ҉)��FDG����8�r������v���8a���9[���#�����*� v�J�:�h���4�S7ΨȯST/<Oj�mZ�M$�{Qij�����_e�]�S\G��^)�͜��eIy�� 3dc�7^� ����*�f��+�/2!�'>�U�qg�%Z��m����j�zQB9���o���%KnƢ������h=�؆�b��P�D�IU$"a����b��%ȯ�C7�p��8�B�ю�D�܉@��OY,�2z��N�@;�j�Jٳ���V=w�l���;T{�fv�z�����8-e���
��3�����Q���%��v^e����Z�  ���#���A9�VKuڴK��Sl�a�m�h�QT�G;�R���\yO�e��[����k��i��5Cܬ_0PX�)�JZy�ru+�1�mA/:�����z��m�X �7^݋���œ�B0�.t��8%kRlR"�I�Yee96l��x��x����5��;s"�vs����j�LOJ�N�YfUaIqy���g�R:n�z��#�D-2�+��Y[�p��?*5�.��ٳQ��������/3��jjŊ�Y9#�EDj�����$�
�(.�Q��%H\M��s�[��\ЗO���Er�
�:XzY��82AS�3�'Q8�p��{�/��;Ϗ�8�ҕ�|=ٌ�^ŒM�dS��q`�B54��`
��R�:��~�}�&�9CT���OU��0P���Y�\��"p����w���6��+hooSצ�̚]�ʪRL���m8,�Z]UB�w)y�R�,������{d�*��l*Xm����ʊ�E����5k)I�B�~I�ڕTvD��m��:-&�!����Qf]�0!r�V��C^��;CE�yH�7o�c+FQJN�m��9:
G�'#!F��\w��	�ebt�Dܶ�6	��댞2����
����=��i*E2�D�yg =]M�m���H:����Q��Tf�x1�������a�O��'FڸF"���Vy)d㶆�
a��D���H��%�v�s:2Re�.��}ߒq�us#�̾�D%�n�G/�ٳ�n�}��1��������@?�ށ'���S+�`Ig�� 3Wra���c͚u���~@\WiMmp��m���p:����Y5�m3�&j�^��t��8��ؠ�p"�7�Q(ʋ�*��^�A��|�W��u@��T�;�"�����Lᑿo�*{ECC䋄�"1�[�$�-b-�ch�
<%�2���*��d���'"���͕�Yu���H�.���ג�@�	T�4�_�C��8}b!��W�X1h;�1cVn�SPJ�������������_?�����k|�+��\~D\ZP�']�s��E3�,�?���*�������uv��bC�=,�#�Bv�$���T�iڼP�.Bf���<2��.	<Fm���DXt/5$����d"�K�^�f��L�Q}\�M�����h�8�k�23k�������?
#D��C}PPR%�����_�r�;��d��`���5�.� s���p�޽����;�]]�8z��,FUumXm�Oj���n���lΕ�zV*��*&���'4������^>�GU*��w��"��W��ыK
���d�̮�f�)�~O��Io38��_���'$^�v�z,[ވ��&bj��nm��%�e�g6��
L��!p>N��B�?H�X��!0��$R����q��A��ғn�|�����ޱ�~�íwm����y$ac=A���O:��Ｙ����:�o;�-s�/TTTJ+3_c�%سw��ղ�'���eAZMj�\8w���9H�B%� ��Ϋ��w]���~ �-^��+�����3��\Ux�CT1�{��A� �f��"&C�@U��ݦ�k7�!d�HEkk����fTa������;w���|�'&��ev��)a�������T�+�	�;��3N����D��J�rz^��N�-`�ʹa{��	�%d��r��S�N�f1���.�SU''pD�7p�&�(9��l��Uh�=�١� ���; ]�LX.��-Bb�Q�Qz&G�6�C��PX �����aƏR�+�%D)3�
��FQ�UX�f-����3���v�;���/퐮�;���O��T�,C(+��`~�+]��q3y��k%kC~�6�\���jdWne�䖔M�|4�i��f����zH�68���+��1��g������i&Jv�l�bR�_�(��/�
	U����@��`���*Ll.�:Iǉ�'���N�TČ�A�jS�ld�z԰��*�r.ڤP��hR�?�6Nn�xI�@�X0>��b�4��ۿ{�>�G0�*�p99����6o�ϣ�C�y�I���Nt���yn.��;��'��X���<E�^m3�j?yr9�l�R�{w�Tr�bnQ����T? ���}&OR�,���w�s��8{n"t\r�vD�6�W�m�Q�Cǎ�{i�Θ/�Z�-LI�N?�E*Ͳ������b��ǫT��)O(����k��&3�/}�sʶL�^���v�r�]'&��b�<T��Rʴ�uw]"�\�-΃�IP6e�I�?7�py\�q���` �Ѿ B#i���{����Io�]�QA��]�����p�q�1�I�G=>>&!�Y��5�ﾌ�-]$)5��
%o�|�-��q��݊C$T*�����o���`�DG�Nb-g�P��ZET-�j�bF�;g>B�4N����+K��U+�e˝�ͳ/���
�ݺ5ՄL��`��w��t7޺ ��>�"�9M6�LH���T�f��č�>�pF\z���Fw�ID���	�D����!����onc;�?��8��S��R��XM��sڮ^śomG2Dw�&�I�j٪qtv!3$T[W�d(j�$l�HϤ)u�w��:��9UUY�L��/-�(V�H��`*��^��S�PQ^���Ohl�A���]��o�a��<i���Ν;	�52��d��+!��4�0�6t����f�Kg
�3C-�^2iD�"؜�,�����xYLv8HN+��n�a)-T.\hF�<�L��4�����_��7������"F�4��I*))��u�Τ9�E𶱒���F�ԡ6il���J���1N6�ad�m�4�*;}�}���\��O��sԛ#�3���/~VuPq��n�>;�fX�'R�)QΡ��r 
Q�H('��*3��p�EK�����b�^QY������N|*N�ٰg��h��I�H���D�#N���Mf�E�.f�a6�Og��Dh�#+19'jY���ϧ�`KE[^�Z7�����s8�.h�����5�^岱��0�3sfLZ|%1��4�L��N%�J(M��f�s�����*.b����m�{G�?0$���8����<y�ۂ��`Ui ���&?A���$|��8I�_C��_���d9%Z�jT�K��gU�E�����rɦ��l��@�ϓF}M�+}�&���t�p�tt��P�W|��`vL�$����i�>gZ�U����;e_���!y��S^V!-��"_�:$aɂ��fP�%�hIњ�0��S�J��3I����b�)�NA��6ֳJd_�H$Sb�TP�!<X�M1,�S����svJ���ڍ�����MY��q���QB-]��B-:��^S%��)L}ϒ0k�/��jjJD���@/�� &m��9�Y!�X�{�i|�-����v)n�֓�qjD7[5٘��x�y8�a1�I���u��L�Ϡ�)��nm`���Mkk���F{!.�R���ÜK���:(��$6�T�����R�<JByi�`�Ò�\і(1�U)�!�y˭�Y����"\m;#�t3���������5TN�M
�8���f��5.M�i�;�"jϦiרǬ^G�Ү��?wdmX:���u����t��d@�q�k��tH㖛*���KѰ����8��ωj��m��~��Tg8m��ᆧ`��ކ�Ko�~�~��꥘b;�7V-��eL}�ڤ��I,ޙ.@ެ^[,�i�K��{�|^�C세���644H��C�|U+��X�_x������diͩ6���~���*��-�]f�>5i�j�, �܅]%�d[�J'>|����|�y��ię���_%.X�¢Z��n�t���a�-��|�:�Gc�Mq?]������#��R��b�x�\�{Xb���^ģG�����~��!��w���%<N�^m�*sl�y?.I:��m�$��K����.��m�2�|\]�3�k���z�ER|4w����$,W2A�,M)2�֬��������p�p��~�gd�G�a�4�ۂ{~A��YL��H��rK#�^�əL��g_M�LV�쟮�s�,���%��Oh+*��C6 kQO�ao�T�M7.����>47sΘ*n�ʑHx���p��i�؊4f5VaFm-��Zۺ3c�����͇�v����濭����z��>���%CR�������/�]`�������x����c��Ո!��1*��$(9�Ƀ�2?�F�Rdl�I�!
�Zn��6U�������=r�n?�ܶ�`�s�����p��EYިɢyf�˅W^{C���DD*U>���Jmɒ��z�=� ���� �y�̜р�� ���_���et|.a�qM�x��-x�9�o�����3��4�ņT{H% ��#���d��*ĸe���g�����ARSE(̋��2��11NVO]�H�$I�J����9�#!���������� �V.Ǯ������<}��/A���UN�'F��S����|s'����N�!1�D�?��b���ͅk�����=�Ҙ>ș;Nk�L1��4��5o���pyi���.Y�ُ�������+����#���� �����2�'a�oM�$�$�A�I���n?q	W�1��K��+/|8��Y�tn\�J���P��p��0~���s�|�����rU|�x*B6�im/�.M��Ȏ��%m��W��s�U�=n��XJ�����1	m�a׼��5	F�;a�cd�5���(>��EE�4��:N����NFJ=t>�V,�����Ȉѵ���#al߾K*�9��;~�fQ2�N�x���n^n�x�cx�7U�mJ��;�܅�̝;O�;�ѥ�����G�I>S��5j��JL��Z��ً�k`E-�*��u���dL#p����ӵ�
ZPӰ2�I�5��{��u��e?C���mx2�k�LB`9��Fv��YXp�b�ryyuu1n�y~��_���#rI���oo'iIJ(��3�*H�Qa�3پcy�}�% K�@�Vݽ��J����&8)'3Q,�ɍ��JҟCcӹ|O��� ������[PS_��{�q��PTֈ��7��7kq�h9�*�����H�ӎ�a��l�qm@�z�˝��l��9��~T�S?G�#�h�|���|W�<��#�н��W�����ho���,Ē���5x�+_%�u��{�P��W@cN�}�$=�茴�7���c��ΈO%�Tۣ�3�wn$M�f�����y�w`֬�G-Da�b�b��m�G�Q5cO�p[0؍��]�t�Y�FW�!x�i���^�f�qz�7�M��l�I����!tv֢��/�'��$$hs��~Q�)~bN3bQC����
�/�#�$?�sot���#�J�I�����aB8w~�l��s�~�B��*��.>�;�,��p��X��R8>���Ã۶c��S��Cw`�,Á]���U����h�&I�trc�}����X��;ë/��C��H��T�j������s��:>��G�KU<W��3�ٙ�V�-�Ϸ���KR��*�jϛ���$q���x�<}�+ϱ.>xln7`��HD��C����oB@΃��ܭ�:��n�r���X�t9��`�S��6*�j�иO��`?ұ	�iUߌ��b��:�BK��ԉCxm�)$U�j��t�?ݡ�%�&�cqW��w�6�5�k�q�q�����G�xfyVdYm,O�B��se�e��[�vb�O������U�����+_���%1Ư~����i?y�9����;���DW4��c��N��+�)��wa�����E�PXЎ����S�v�[���r";}Uh�K�I�T\#YO7�0�_� �\C�k�feJ?� ����z�O�zj�8�����w��]���kK/����}��~��gp�d���k*�'?�ֳ����&N�vD��+8�G��f=*N=K�[ye�-Ö�yU���k��Ų �T"�r�T��{n�w�{��T5��~� �4u,S�ט�Y.r��?����O|^�Zk���O�d��ԝ[��?�>���x�i����Q��D�*gm�/�lq��n�>�l���̮H��@zRm�Y�U���X��r;���s�ܨ����~ߺ����:���FҬTZc�u���Y����s��{%7l؀G}��Ͽ��S���-[�`��[�o�>?v�|���u������	��I���+�����#���B��5&d;=Qb���
5��|������rPP7����e�f���P�[������3[��o�Tè-����f%|.�[���>��bi�6� ��k榧yxޘ���sfϖ����C�O#�9|>    IEND�B`�PK 
     #{dZ�5,*Q Q                  cirkitFile.jsonPK 
     #{dZ                        HQ jsons/PK 
     #{dZR�1FPt  Pt               lQ jsons/user_defined.jsonPK 
     #{dZ                        �� images/PK 
     #{dZ�&�y`  y`  /             � images/8c2f1315-cf23-4ba8-a920-becb97f13280.pngPK 
     #{dZ�����  �  /             �& images/6fc4b800-efc3-4a5d-827d-9566cfd108b3.pngPK 
     #{dZ�?���� �� /             9 images/ae82c023-d9d4-4942-aa8d-ab2ae3c53d73.pngPK 
     #{dZ�S��*  �*  /             �� images/cbf7ad0e-0f08-44f8-98a9-dcbe92af212f.pngPK 
     #{dZ�+s`(  `(  /              images/8a1d81a5-79d4-450c-9f72-108cd2673013.pngPK 
     #{dZ��/��  �  /             �6 images/aacc0029-e57d-4614-a443-d9bee65b5175.pngPK 
     #{dZ�1��� �� /             �B images/1d90a712-93d7-4555-ae10-1782f839eba3.pngPK 
     #{dZ��S�  S�  /             ]� images/e5551f5a-2fb7-4493-9527-57db21faeaae.pngPK 
     #{dZ?�>�oH  oH  /             �� images/a038ca8d-f9eb-4e93-ad0b-b831193aa106.pngPK 
     #{dZ-s;�.@  .@  /             �0 images/3e0a96b2-ef1c-4fb2-8b57-d71cbe1f3744.pngPK 
     #{dZ3��C� � /             4q images/cff7cff8-0125-49f3-ae91-9e6ccc0a4cc7.pngPK 
     #{dZ��� �� /             �' images/7b19d218-2217-455d-9a43-b73a208c2c5c.pngPK 
     #{dZF�i~�  �  /             �� images/85e66502-362d-4a26-afcd-97fbc4859675.pngPK 
     #{dZ�  ��  /             �� images/b13518ba-21c5-4f60-a735-1d8041d11d7b.pngPK 
     #{dZt��n� n� /             �� images/c750f18a-9432-41e6-a6ed-179e28bc29f6.pngPK 
     #{dZH��`�b  �b  /             J�* images/3f9b3f3f-db41-4a6d-b13c-7e86a7741a7b.pngPK 
     #{dZ��_mE E /             u9+ images/28139415-969f-45d3-9930-3634e76076d7.pngPK 
     #{dZ
��
  
  /             H3 images/edf2d60f-7dc2-4972-a04c-2a93629ecddc.pngPK      u  ^�3   